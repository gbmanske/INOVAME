//Benchmark atmr_intb_466_0.125

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n293_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n321_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n351_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n422_, men_men_n423_, men_men_n424_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  AOI220     o035(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n57_), .Y(ori_ori_n58_));
  INV        o036(.A(ori_ori_n55_), .Y(ori_ori_n59_));
  OAI220     o037(.A0(x02), .A1(ori_ori_n59_), .B0(ori_ori_n58_), .B1(ori_ori_n56_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n61_));
  OAI210     o039(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n61_), .Y(ori_ori_n62_));
  AOI220     o040(.A0(ori_ori_n62_), .A1(ori_ori_n55_), .B0(ori_ori_n60_), .B1(ori_ori_n31_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(x05), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n57_), .B(ori_ori_n23_), .Y(ori_ori_n65_));
  NA2        o043(.A(x09), .B(x05), .Y(ori_ori_n66_));
  NA2        o044(.A(x10), .B(x06), .Y(ori_ori_n67_));
  NA3        o045(.A(ori_ori_n67_), .B(ori_ori_n66_), .C(ori_ori_n28_), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n57_), .B(ori_ori_n41_), .Y(ori_ori_n69_));
  OAI210     o047(.A0(ori_ori_n68_), .A1(ori_ori_n65_), .B0(x03), .Y(ori_ori_n70_));
  NOi31      o048(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n72_));
  NO2        o050(.A(x08), .B(x01), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n73_), .A1(ori_ori_n72_), .B0(ori_ori_n35_), .Y(ori_ori_n74_));
  NA2        o052(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n74_), .B(x02), .Y(ori_ori_n76_));
  AN2        o054(.A(ori_ori_n76_), .B(ori_ori_n70_), .Y(ori_ori_n77_));
  INV        o055(.A(ori_ori_n74_), .Y(ori_ori_n78_));
  NA2        o056(.A(x11), .B(x00), .Y(ori_ori_n79_));
  NO2        o057(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n80_));
  NOi21      o058(.An(ori_ori_n79_), .B(ori_ori_n80_), .Y(ori_ori_n81_));
  NOi21      o059(.An(x01), .B(x10), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n83_));
  NO3        o061(.A(ori_ori_n83_), .B(ori_ori_n82_), .C(x06), .Y(ori_ori_n84_));
  NA2        o062(.A(ori_ori_n84_), .B(ori_ori_n27_), .Y(ori_ori_n85_));
  OAI210     o063(.A0(ori_ori_n334_), .A1(x07), .B0(ori_ori_n85_), .Y(ori_ori_n86_));
  NO3        o064(.A(ori_ori_n86_), .B(ori_ori_n77_), .C(ori_ori_n64_), .Y(ori01));
  INV        o065(.A(x12), .Y(ori_ori_n88_));
  INV        o066(.A(x13), .Y(ori_ori_n89_));
  NA2        o067(.A(ori_ori_n82_), .B(ori_ori_n28_), .Y(ori_ori_n90_));
  NO2        o068(.A(x10), .B(x01), .Y(ori_ori_n91_));
  NO2        o069(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NA2        o071(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n96_));
  INV        o074(.A(x13), .Y(ori_ori_n97_));
  NO2        o075(.A(ori_ori_n97_), .B(x05), .Y(ori_ori_n98_));
  NA2        o076(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n100_));
  NA2        o078(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n104_));
  NA3        o082(.A(ori_ori_n104_), .B(ori_ori_n103_), .C(x13), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n106_));
  NOi31      o084(.An(ori_ori_n105_), .B(ori_ori_n106_), .C(ori_ori_n102_), .Y(ori_ori_n107_));
  NO3        o085(.A(ori_ori_n107_), .B(x06), .C(x03), .Y(ori_ori_n108_));
  INV        o086(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NA2        o087(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n110_));
  OAI210     o088(.A0(ori_ori_n73_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n111_), .B(ori_ori_n110_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n114_));
  AOI210     o092(.A0(ori_ori_n114_), .A1(ori_ori_n49_), .B0(ori_ori_n113_), .Y(ori_ori_n115_));
  AN2        o093(.A(ori_ori_n115_), .B(ori_ori_n112_), .Y(ori_ori_n116_));
  NO2        o094(.A(x09), .B(x05), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n117_), .B(ori_ori_n47_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n93_), .B(ori_ori_n49_), .Y(ori_ori_n119_));
  NA2        o097(.A(x09), .B(x00), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n95_), .B(ori_ori_n120_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n119_), .B(ori_ori_n116_), .Y(ori_ori_n122_));
  NO2        o100(.A(x03), .B(x02), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n74_), .B(ori_ori_n89_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(ori_ori_n123_), .Y(ori_ori_n125_));
  OA210      o103(.A0(ori_ori_n122_), .A1(x11), .B0(ori_ori_n125_), .Y(ori_ori_n126_));
  OAI210     o104(.A0(ori_ori_n109_), .A1(ori_ori_n23_), .B0(ori_ori_n126_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n93_), .B(ori_ori_n40_), .Y(ori_ori_n128_));
  NOi21      o106(.An(x01), .B(x13), .Y(ori_ori_n129_));
  INV        o107(.A(ori_ori_n129_), .Y(ori_ori_n130_));
  NO2        o108(.A(ori_ori_n128_), .B(ori_ori_n41_), .Y(ori_ori_n131_));
  NO2        o109(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n89_), .B(x01), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n133_), .B(x08), .Y(ori_ori_n134_));
  NO2        o112(.A(ori_ori_n132_), .B(ori_ori_n48_), .Y(ori_ori_n135_));
  AOI210     o113(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n136_));
  OAI210     o114(.A0(ori_ori_n135_), .A1(ori_ori_n131_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  NA2        o115(.A(x10), .B(x05), .Y(ori_ori_n138_));
  INV        o116(.A(ori_ori_n25_), .Y(ori_ori_n139_));
  AN2        o117(.A(ori_ori_n67_), .B(ori_ori_n66_), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n83_), .B(x06), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n142_), .B(ori_ori_n139_), .Y(ori_ori_n143_));
  NOi21      o121(.An(x09), .B(x00), .Y(ori_ori_n144_));
  NO3        o122(.A(ori_ori_n72_), .B(ori_ori_n144_), .C(ori_ori_n47_), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n145_), .B(ori_ori_n101_), .Y(ori_ori_n146_));
  NA2        o124(.A(x06), .B(x05), .Y(ori_ori_n147_));
  OAI210     o125(.A0(ori_ori_n147_), .A1(ori_ori_n35_), .B0(ori_ori_n88_), .Y(ori_ori_n148_));
  AOI210     o126(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n148_), .Y(ori_ori_n149_));
  NA2        o127(.A(ori_ori_n149_), .B(ori_ori_n146_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n89_), .B(x12), .Y(ori_ori_n151_));
  AOI210     o129(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n151_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n153_), .B(x02), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n152_), .B(ori_ori_n150_), .Y(ori_ori_n155_));
  NA3        o133(.A(ori_ori_n155_), .B(ori_ori_n143_), .C(ori_ori_n137_), .Y(ori_ori_n156_));
  AOI210     o134(.A0(ori_ori_n127_), .A1(ori_ori_n88_), .B0(ori_ori_n156_), .Y(ori_ori_n157_));
  INV        o135(.A(ori_ori_n68_), .Y(ori_ori_n158_));
  NA2        o136(.A(ori_ori_n158_), .B(ori_ori_n112_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n100_), .B(x06), .Y(ori_ori_n160_));
  INV        o138(.A(ori_ori_n160_), .Y(ori_ori_n161_));
  AOI210     o139(.A0(ori_ori_n161_), .A1(ori_ori_n159_), .B0(x12), .Y(ori_ori_n162_));
  INV        o140(.A(ori_ori_n71_), .Y(ori_ori_n163_));
  NO2        o141(.A(x05), .B(ori_ori_n50_), .Y(ori_ori_n164_));
  OAI210     o142(.A0(ori_ori_n164_), .A1(ori_ori_n130_), .B0(ori_ori_n53_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n165_), .B(ori_ori_n163_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n82_), .B(x06), .Y(ori_ori_n167_));
  AOI210     o145(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n168_));
  NO3        o146(.A(ori_ori_n168_), .B(ori_ori_n167_), .C(ori_ori_n41_), .Y(ori_ori_n169_));
  NA2        o147(.A(ori_ori_n169_), .B(x02), .Y(ori_ori_n170_));
  AOI210     o148(.A0(ori_ori_n170_), .A1(ori_ori_n166_), .B0(ori_ori_n23_), .Y(ori_ori_n171_));
  OAI210     o149(.A0(ori_ori_n162_), .A1(ori_ori_n53_), .B0(ori_ori_n171_), .Y(ori_ori_n172_));
  INV        o150(.A(ori_ori_n114_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n71_), .B(ori_ori_n174_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n176_));
  NOi21      o154(.An(x13), .B(x04), .Y(ori_ori_n177_));
  NO3        o155(.A(ori_ori_n177_), .B(ori_ori_n71_), .C(ori_ori_n144_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n178_), .B(x05), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n179_), .B(ori_ori_n176_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n175_), .B(ori_ori_n180_), .Y(ori_ori_n181_));
  INV        o159(.A(ori_ori_n80_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n182_), .B(x12), .Y(ori_ori_n183_));
  NA2        o161(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n185_));
  AOI210     o163(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n186_), .B(ori_ori_n41_), .Y(ori_ori_n187_));
  INV        o165(.A(ori_ori_n187_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n189_), .B(x03), .Y(ori_ori_n190_));
  OR2        o168(.A(ori_ori_n190_), .B(ori_ori_n188_), .Y(ori_ori_n191_));
  NA2        o169(.A(x13), .B(ori_ori_n88_), .Y(ori_ori_n192_));
  NA3        o170(.A(ori_ori_n192_), .B(ori_ori_n148_), .C(ori_ori_n81_), .Y(ori_ori_n193_));
  OAI210     o171(.A0(ori_ori_n191_), .A1(ori_ori_n184_), .B0(ori_ori_n193_), .Y(ori_ori_n194_));
  AOI210     o172(.A0(ori_ori_n183_), .A1(ori_ori_n181_), .B0(ori_ori_n194_), .Y(ori_ori_n195_));
  AOI210     o173(.A0(ori_ori_n195_), .A1(ori_ori_n172_), .B0(x07), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n66_), .B(ori_ori_n29_), .Y(ori_ori_n197_));
  NOi31      o175(.An(ori_ori_n110_), .B(ori_ori_n177_), .C(ori_ori_n144_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n198_), .B(ori_ori_n197_), .Y(ori_ori_n199_));
  OAI210     o177(.A0(ori_ori_n71_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n200_));
  INV        o178(.A(ori_ori_n200_), .Y(ori_ori_n201_));
  NO2        o179(.A(x12), .B(x02), .Y(ori_ori_n202_));
  INV        o180(.A(ori_ori_n202_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n203_), .B(ori_ori_n182_), .Y(ori_ori_n204_));
  OA210      o182(.A0(ori_ori_n201_), .A1(ori_ori_n199_), .B0(ori_ori_n204_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(x01), .Y(ori_ori_n207_));
  INV        o185(.A(ori_ori_n207_), .Y(ori_ori_n208_));
  AOI210     o186(.A0(ori_ori_n208_), .A1(ori_ori_n105_), .B0(ori_ori_n29_), .Y(ori_ori_n209_));
  NA2        o187(.A(ori_ori_n89_), .B(x04), .Y(ori_ori_n210_));
  NO3        o188(.A(ori_ori_n79_), .B(x12), .C(x03), .Y(ori_ori_n211_));
  NA2        o189(.A(ori_ori_n209_), .B(ori_ori_n211_), .Y(ori_ori_n212_));
  NOi21      o190(.An(ori_ori_n197_), .B(ori_ori_n167_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n214_));
  NA2        o192(.A(ori_ori_n213_), .B(ori_ori_n214_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n216_));
  NO3        o194(.A(ori_ori_n216_), .B(ori_ori_n168_), .C(ori_ori_n141_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n184_), .B(ori_ori_n28_), .Y(ori_ori_n218_));
  OAI210     o196(.A0(ori_ori_n217_), .A1(ori_ori_n173_), .B0(ori_ori_n218_), .Y(ori_ori_n219_));
  NA3        o197(.A(ori_ori_n219_), .B(ori_ori_n215_), .C(ori_ori_n212_), .Y(ori_ori_n220_));
  NO3        o198(.A(ori_ori_n220_), .B(ori_ori_n205_), .C(ori_ori_n196_), .Y(ori_ori_n221_));
  OAI210     o199(.A0(ori_ori_n157_), .A1(ori_ori_n57_), .B0(ori_ori_n221_), .Y(ori02));
  AOI210     o200(.A0(ori_ori_n110_), .A1(ori_ori_n74_), .B0(ori_ori_n103_), .Y(ori_ori_n223_));
  BUFFER     o201(.A(ori_ori_n178_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n224_), .B(ori_ori_n32_), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n225_), .A1(ori_ori_n223_), .B0(ori_ori_n138_), .Y(ori_ori_n226_));
  INV        o204(.A(ori_ori_n138_), .Y(ori_ori_n227_));
  AOI210     o205(.A0(ori_ori_n96_), .A1(ori_ori_n75_), .B0(ori_ori_n168_), .Y(ori_ori_n228_));
  OAI220     o206(.A0(ori_ori_n228_), .A1(ori_ori_n89_), .B0(ori_ori_n74_), .B1(ori_ori_n50_), .Y(ori_ori_n229_));
  AOI220     o207(.A0(ori_ori_n229_), .A1(ori_ori_n227_), .B0(ori_ori_n124_), .B1(ori_ori_n123_), .Y(ori_ori_n230_));
  AOI210     o208(.A0(ori_ori_n230_), .A1(ori_ori_n226_), .B0(ori_ori_n48_), .Y(ori_ori_n231_));
  NAi21      o209(.An(ori_ori_n179_), .B(ori_ori_n175_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n189_), .B(ori_ori_n47_), .Y(ori_ori_n233_));
  NA2        o211(.A(ori_ori_n233_), .B(ori_ori_n232_), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n235_));
  AOI210     o213(.A0(ori_ori_n337_), .A1(ori_ori_n111_), .B0(ori_ori_n235_), .Y(ori_ori_n236_));
  NA2        o214(.A(ori_ori_n236_), .B(ori_ori_n83_), .Y(ori_ori_n237_));
  INV        o215(.A(ori_ori_n123_), .Y(ori_ori_n238_));
  OAI210     o216(.A0(ori_ori_n238_), .A1(ori_ori_n102_), .B0(ori_ori_n90_), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n239_), .B(x13), .Y(ori_ori_n240_));
  NA3        o218(.A(ori_ori_n240_), .B(ori_ori_n237_), .C(ori_ori_n234_), .Y(ori_ori_n241_));
  NO2        o219(.A(ori_ori_n241_), .B(ori_ori_n231_), .Y(ori_ori_n242_));
  NA2        o220(.A(ori_ori_n113_), .B(x03), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n35_), .B(ori_ori_n36_), .Y(ori_ori_n244_));
  AOI220     o222(.A0(ori_ori_n244_), .A1(ori_ori_n336_), .B0(ori_ori_n153_), .B1(x08), .Y(ori_ori_n245_));
  OAI210     o223(.A0(ori_ori_n245_), .A1(ori_ori_n216_), .B0(ori_ori_n243_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(ori_ori_n91_), .Y(ori_ori_n247_));
  OAI220     o225(.A0(ori_ori_n210_), .A1(x09), .B0(ori_ori_n103_), .B1(ori_ori_n28_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n248_), .B(ori_ori_n92_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n210_), .B(ori_ori_n88_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n88_), .B(ori_ori_n41_), .Y(ori_ori_n251_));
  NA3        o229(.A(ori_ori_n251_), .B(ori_ori_n250_), .C(ori_ori_n102_), .Y(ori_ori_n252_));
  NA4        o230(.A(ori_ori_n252_), .B(ori_ori_n249_), .C(ori_ori_n247_), .D(ori_ori_n48_), .Y(ori_ori_n253_));
  INV        o231(.A(ori_ori_n153_), .Y(ori_ori_n254_));
  NO2        o232(.A(ori_ori_n134_), .B(ori_ori_n40_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n256_));
  OAI220     o234(.A0(ori_ori_n256_), .A1(ori_ori_n255_), .B0(ori_ori_n254_), .B1(ori_ori_n55_), .Y(ori_ori_n257_));
  NA2        o235(.A(ori_ori_n257_), .B(x02), .Y(ori_ori_n258_));
  INV        o236(.A(ori_ori_n185_), .Y(ori_ori_n259_));
  NA2        o237(.A(ori_ori_n151_), .B(x04), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n151_), .B(ori_ori_n132_), .C(ori_ori_n51_), .Y(ori_ori_n261_));
  OAI210     o239(.A0(ori_ori_n120_), .A1(ori_ori_n36_), .B0(ori_ori_n88_), .Y(ori_ori_n262_));
  OAI210     o240(.A0(ori_ori_n262_), .A1(ori_ori_n145_), .B0(ori_ori_n261_), .Y(ori_ori_n263_));
  NA3        o241(.A(ori_ori_n263_), .B(ori_ori_n258_), .C(x06), .Y(ori_ori_n264_));
  NO3        o242(.A(ori_ori_n216_), .B(ori_ori_n100_), .C(x08), .Y(ori_ori_n265_));
  INV        o243(.A(ori_ori_n265_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n267_));
  NO3        o245(.A(ori_ori_n95_), .B(ori_ori_n101_), .C(ori_ori_n38_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n261_), .A1(ori_ori_n267_), .B0(ori_ori_n268_), .Y(ori_ori_n269_));
  OAI210     o247(.A0(ori_ori_n266_), .A1(ori_ori_n28_), .B0(ori_ori_n269_), .Y(ori_ori_n270_));
  AN2        o248(.A(ori_ori_n270_), .B(x04), .Y(ori_ori_n271_));
  AOI210     o249(.A0(ori_ori_n264_), .A1(ori_ori_n253_), .B0(ori_ori_n271_), .Y(ori_ori_n272_));
  OAI210     o250(.A0(ori_ori_n242_), .A1(x12), .B0(ori_ori_n272_), .Y(ori03));
  OR2        o251(.A(ori_ori_n42_), .B(ori_ori_n174_), .Y(ori_ori_n274_));
  AOI210     o252(.A0(ori_ori_n124_), .A1(ori_ori_n88_), .B0(ori_ori_n274_), .Y(ori_ori_n275_));
  AO210      o253(.A0(ori_ori_n259_), .A1(ori_ori_n75_), .B0(ori_ori_n260_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n151_), .B(ori_ori_n123_), .Y(ori_ori_n277_));
  NA3        o255(.A(ori_ori_n277_), .B(ori_ori_n276_), .C(ori_ori_n154_), .Y(ori_ori_n278_));
  OAI210     o256(.A0(ori_ori_n278_), .A1(ori_ori_n275_), .B0(x05), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n274_), .B(x05), .Y(ori_ori_n280_));
  AOI210     o258(.A0(ori_ori_n111_), .A1(ori_ori_n163_), .B0(ori_ori_n280_), .Y(ori_ori_n281_));
  INV        o259(.A(ori_ori_n98_), .Y(ori_ori_n282_));
  NO2        o260(.A(ori_ori_n282_), .B(ori_ori_n55_), .Y(ori_ori_n283_));
  OAI210     o261(.A0(ori_ori_n283_), .A1(ori_ori_n281_), .B0(ori_ori_n88_), .Y(ori_ori_n284_));
  AOI210     o262(.A0(ori_ori_n118_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n285_));
  NO2        o263(.A(ori_ori_n121_), .B(x13), .Y(ori_ori_n286_));
  OAI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n285_), .B0(x04), .Y(ori_ori_n287_));
  NO3        o265(.A(ori_ori_n251_), .B(ori_ori_n74_), .C(ori_ori_n55_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n88_), .B(ori_ori_n118_), .Y(ori_ori_n289_));
  OA210      o267(.A0(ori_ori_n134_), .A1(x12), .B0(ori_ori_n106_), .Y(ori_ori_n290_));
  NO3        o268(.A(ori_ori_n290_), .B(ori_ori_n289_), .C(ori_ori_n288_), .Y(ori_ori_n291_));
  NA4        o269(.A(ori_ori_n291_), .B(ori_ori_n287_), .C(ori_ori_n284_), .D(ori_ori_n279_), .Y(ori04));
  NO2        o270(.A(ori_ori_n78_), .B(ori_ori_n39_), .Y(ori_ori_n293_));
  XO2        o271(.A(ori_ori_n293_), .B(ori_ori_n192_), .Y(ori05));
  AOI210     o272(.A0(ori_ori_n66_), .A1(ori_ori_n51_), .B0(ori_ori_n160_), .Y(ori_ori_n295_));
  AOI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n235_), .B0(ori_ori_n25_), .Y(ori_ori_n296_));
  AOI210     o274(.A0(x06), .A1(x03), .B0(ori_ori_n24_), .Y(ori_ori_n297_));
  OAI210     o275(.A0(ori_ori_n297_), .A1(ori_ori_n296_), .B0(ori_ori_n88_), .Y(ori_ori_n298_));
  NA2        o276(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n300_));
  NA2        o278(.A(ori_ori_n197_), .B(x03), .Y(ori_ori_n301_));
  OAI210     o279(.A0(ori_ori_n301_), .A1(ori_ori_n300_), .B0(ori_ori_n299_), .Y(ori_ori_n302_));
  OAI210     o280(.A0(ori_ori_n26_), .A1(ori_ori_n88_), .B0(x07), .Y(ori_ori_n303_));
  AOI210     o281(.A0(ori_ori_n302_), .A1(x06), .B0(ori_ori_n303_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n23_), .B(x00), .Y(ori_ori_n305_));
  OAI210     o283(.A0(ori_ori_n335_), .A1(ori_ori_n305_), .B0(ori_ori_n88_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n33_), .B(ori_ori_n88_), .Y(ori_ori_n307_));
  AOI210     o285(.A0(ori_ori_n307_), .A1(ori_ori_n80_), .B0(x07), .Y(ori_ori_n308_));
  AOI220     o286(.A0(ori_ori_n308_), .A1(ori_ori_n306_), .B0(ori_ori_n304_), .B1(ori_ori_n298_), .Y(ori_ori_n309_));
  AOI210     o287(.A0(ori_ori_n260_), .A1(ori_ori_n94_), .B0(ori_ori_n202_), .Y(ori_ori_n310_));
  NOi21      o288(.An(ori_ori_n243_), .B(ori_ori_n106_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n311_), .B(ori_ori_n203_), .Y(ori_ori_n312_));
  AOI210     o290(.A0(ori_ori_n192_), .A1(ori_ori_n47_), .B0(x04), .Y(ori_ori_n313_));
  NO4        o291(.A(ori_ori_n313_), .B(ori_ori_n312_), .C(ori_ori_n310_), .D(x08), .Y(ori_ori_n314_));
  NO2        o292(.A(ori_ori_n103_), .B(ori_ori_n28_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n315_), .B(ori_ori_n207_), .Y(ori_ori_n316_));
  NA3        o294(.A(ori_ori_n254_), .B(ori_ori_n99_), .C(x12), .Y(ori_ori_n317_));
  NA2        o295(.A(ori_ori_n317_), .B(x08), .Y(ori_ori_n318_));
  INV        o296(.A(ori_ori_n318_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n314_), .B(ori_ori_n319_), .Y(ori_ori_n320_));
  NA3        o298(.A(ori_ori_n316_), .B(ori_ori_n311_), .C(ori_ori_n250_), .Y(ori_ori_n321_));
  INV        o299(.A(x14), .Y(ori_ori_n322_));
  NO3        o300(.A(ori_ori_n133_), .B(ori_ori_n69_), .C(ori_ori_n53_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n323_), .B(ori_ori_n322_), .Y(ori_ori_n324_));
  NA2        o302(.A(ori_ori_n324_), .B(ori_ori_n321_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n307_), .B(ori_ori_n57_), .Y(ori_ori_n326_));
  NOi21      o304(.An(ori_ori_n210_), .B(ori_ori_n121_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n328_));
  OAI210     o306(.A0(ori_ori_n328_), .A1(ori_ori_n327_), .B0(ori_ori_n88_), .Y(ori_ori_n329_));
  OAI210     o307(.A0(ori_ori_n326_), .A1(ori_ori_n79_), .B0(ori_ori_n329_), .Y(ori_ori_n330_));
  NO4        o308(.A(ori_ori_n330_), .B(ori_ori_n325_), .C(ori_ori_n320_), .D(ori_ori_n309_), .Y(ori06));
  INV        o309(.A(ori_ori_n81_), .Y(ori_ori_n334_));
  INV        o310(.A(ori_ori_n184_), .Y(ori_ori_n335_));
  INV        o311(.A(x13), .Y(ori_ori_n336_));
  INV        o312(.A(x13), .Y(ori_ori_n337_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NO2        m030(.A(x09), .B(x07), .Y(mai_mai_n53_));
  OAI210     m031(.A0(mai_mai_n53_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n54_));
  NOi21      m032(.An(x01), .B(x09), .Y(mai_mai_n55_));
  INV        m033(.A(x00), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n51_), .B(mai_mai_n56_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(x09), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m037(.A(x07), .Y(mai_mai_n60_));
  INV        m038(.A(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n62_), .B(mai_mai_n24_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(mai_mai_n61_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n31_), .Y(mai_mai_n65_));
  AOI210     m043(.A0(mai_mai_n65_), .A1(mai_mai_n54_), .B0(x05), .Y(mai_mai_n66_));
  NA2        m044(.A(x09), .B(x05), .Y(mai_mai_n67_));
  NA2        m045(.A(x10), .B(x06), .Y(mai_mai_n68_));
  NA2        m046(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  OAI210     m047(.A0(mai_mai_n69_), .A1(x11), .B0(x03), .Y(mai_mai_n70_));
  NOi31      m048(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n71_));
  NO2        m049(.A(mai_mai_n379_), .B(mai_mai_n24_), .Y(mai_mai_n72_));
  NO2        m050(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n48_), .B(mai_mai_n74_), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n76_));
  NO2        m054(.A(x08), .B(x01), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n77_), .A1(mai_mai_n76_), .B0(mai_mai_n35_), .Y(mai_mai_n78_));
  NA2        m056(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n79_));
  NO3        m057(.A(mai_mai_n78_), .B(mai_mai_n75_), .C(mai_mai_n72_), .Y(mai_mai_n80_));
  AN2        m058(.A(mai_mai_n80_), .B(mai_mai_n70_), .Y(mai_mai_n81_));
  INV        m059(.A(mai_mai_n78_), .Y(mai_mai_n82_));
  NO2        m060(.A(x06), .B(x05), .Y(mai_mai_n83_));
  NA2        m061(.A(x11), .B(x00), .Y(mai_mai_n84_));
  NO2        m062(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n85_));
  NOi21      m063(.An(mai_mai_n84_), .B(mai_mai_n85_), .Y(mai_mai_n86_));
  AOI210     m064(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n86_), .Y(mai_mai_n87_));
  NOi21      m065(.An(x01), .B(x10), .Y(mai_mai_n88_));
  NO2        m066(.A(mai_mai_n29_), .B(mai_mai_n56_), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n88_), .C(x06), .Y(mai_mai_n90_));
  NA2        m068(.A(mai_mai_n90_), .B(mai_mai_n27_), .Y(mai_mai_n91_));
  OAI210     m069(.A0(mai_mai_n87_), .A1(x07), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NO3        m070(.A(mai_mai_n92_), .B(mai_mai_n81_), .C(mai_mai_n66_), .Y(mai01));
  INV        m071(.A(x12), .Y(mai_mai_n94_));
  INV        m072(.A(x13), .Y(mai_mai_n95_));
  NA2        m073(.A(x08), .B(x04), .Y(mai_mai_n96_));
  NA2        m074(.A(x04), .B(mai_mai_n83_), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n88_), .B(mai_mai_n28_), .Y(mai_mai_n98_));
  NO2        m076(.A(x10), .B(x01), .Y(mai_mai_n99_));
  NO2        m077(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NA2        m079(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n102_));
  NO3        m080(.A(mai_mai_n102_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n385_), .Y(mai_mai_n104_));
  AOI210     m082(.A0(mai_mai_n104_), .A1(mai_mai_n97_), .B0(mai_mai_n95_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n55_), .B(x05), .Y(mai_mai_n106_));
  NOi21      m084(.An(mai_mai_n106_), .B(mai_mai_n57_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n108_));
  NA3        m086(.A(x13), .B(mai_mai_n108_), .C(x06), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n107_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n77_), .B(x13), .Y(mai_mai_n111_));
  NA2        m089(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(x05), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n35_), .B(mai_mai_n56_), .Y(mai_mai_n114_));
  AOI210     m092(.A0(mai_mai_n35_), .A1(x08), .B0(mai_mai_n107_), .Y(mai_mai_n115_));
  AOI210     m093(.A0(mai_mai_n115_), .A1(mai_mai_n111_), .B0(mai_mai_n68_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n117_));
  NA2        m095(.A(x10), .B(mai_mai_n56_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n59_), .B(x05), .Y(mai_mai_n121_));
  NO3        m099(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n122_));
  NO4        m100(.A(mai_mai_n122_), .B(mai_mai_n116_), .C(mai_mai_n110_), .D(mai_mai_n105_), .Y(mai_mai_n123_));
  NA2        m101(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n124_));
  OAI210     m102(.A0(mai_mai_n77_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n126_));
  NO2        m104(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n128_));
  AOI210     m106(.A0(mai_mai_n128_), .A1(mai_mai_n49_), .B0(mai_mai_n127_), .Y(mai_mai_n129_));
  AN2        m107(.A(mai_mai_n129_), .B(mai_mai_n126_), .Y(mai_mai_n130_));
  NO2        m108(.A(x09), .B(x05), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(mai_mai_n47_), .Y(mai_mai_n132_));
  AOI210     m110(.A0(mai_mai_n132_), .A1(mai_mai_n101_), .B0(mai_mai_n49_), .Y(mai_mai_n133_));
  NA2        m111(.A(x09), .B(x00), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n106_), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NA2        m113(.A(mai_mai_n71_), .B(mai_mai_n51_), .Y(mai_mai_n136_));
  AOI210     m114(.A0(mai_mai_n136_), .A1(mai_mai_n135_), .B0(mai_mai_n128_), .Y(mai_mai_n137_));
  NO3        m115(.A(mai_mai_n137_), .B(mai_mai_n133_), .C(mai_mai_n130_), .Y(mai_mai_n138_));
  NO2        m116(.A(x03), .B(x02), .Y(mai_mai_n139_));
  NA2        m117(.A(mai_mai_n78_), .B(mai_mai_n95_), .Y(mai_mai_n140_));
  OAI210     m118(.A0(mai_mai_n140_), .A1(mai_mai_n107_), .B0(mai_mai_n139_), .Y(mai_mai_n141_));
  OA210      m119(.A0(mai_mai_n138_), .A1(x11), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  OAI210     m120(.A0(mai_mai_n123_), .A1(mai_mai_n23_), .B0(mai_mai_n142_), .Y(mai_mai_n143_));
  NAi21      m121(.An(x06), .B(x10), .Y(mai_mai_n144_));
  NOi21      m122(.An(x01), .B(x13), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n95_), .B(x01), .Y(mai_mai_n147_));
  AOI210     m125(.A0(x09), .A1(mai_mai_n146_), .B0(mai_mai_n48_), .Y(mai_mai_n148_));
  AOI210     m126(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n148_), .A1(mai_mai_n145_), .B0(mai_mai_n149_), .Y(mai_mai_n150_));
  NA2        m128(.A(x04), .B(x02), .Y(mai_mai_n151_));
  NA2        m129(.A(x10), .B(x05), .Y(mai_mai_n152_));
  NO2        m130(.A(x09), .B(x01), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n106_), .B(x08), .Y(mai_mai_n154_));
  NAi21      m132(.An(mai_mai_n151_), .B(mai_mai_n383_), .Y(mai_mai_n155_));
  INV        m133(.A(mai_mai_n25_), .Y(mai_mai_n156_));
  NAi21      m134(.An(x13), .B(x00), .Y(mai_mai_n157_));
  AOI210     m135(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  AN2        m136(.A(x04), .B(mai_mai_n158_), .Y(mai_mai_n159_));
  BUFFER     m137(.A(mai_mai_n67_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n89_), .B(x06), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n157_), .B(mai_mai_n36_), .Y(mai_mai_n162_));
  INV        m140(.A(mai_mai_n162_), .Y(mai_mai_n163_));
  OAI210     m141(.A0(mai_mai_n161_), .A1(mai_mai_n160_), .B0(mai_mai_n163_), .Y(mai_mai_n164_));
  OAI210     m142(.A0(mai_mai_n164_), .A1(mai_mai_n159_), .B0(mai_mai_n156_), .Y(mai_mai_n165_));
  NOi21      m143(.An(x09), .B(x00), .Y(mai_mai_n166_));
  NA2        m144(.A(x06), .B(x05), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n95_), .B(x12), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n88_), .B(mai_mai_n51_), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n169_), .B(x12), .Y(mai_mai_n172_));
  NA4        m150(.A(mai_mai_n172_), .B(mai_mai_n165_), .C(mai_mai_n155_), .D(mai_mai_n150_), .Y(mai_mai_n173_));
  AOI210     m151(.A0(mai_mai_n143_), .A1(mai_mai_n94_), .B0(mai_mai_n173_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n28_), .B(mai_mai_n126_), .Y(mai_mai_n175_));
  NA2        m153(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n176_));
  NA2        m154(.A(mai_mai_n176_), .B(mai_mai_n125_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n382_), .B(mai_mai_n177_), .Y(mai_mai_n178_));
  AOI210     m156(.A0(mai_mai_n178_), .A1(mai_mai_n175_), .B0(x12), .Y(mai_mai_n179_));
  INV        m157(.A(mai_mai_n71_), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n88_), .B(x06), .Y(mai_mai_n181_));
  AOI210     m159(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n182_));
  NO3        m160(.A(mai_mai_n182_), .B(mai_mai_n181_), .C(mai_mai_n41_), .Y(mai_mai_n183_));
  NA4        m161(.A(mai_mai_n144_), .B(mai_mai_n55_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n184_));
  NA2        m162(.A(mai_mai_n184_), .B(mai_mai_n128_), .Y(mai_mai_n185_));
  OAI210     m163(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(x02), .Y(mai_mai_n186_));
  AOI210     m164(.A0(mai_mai_n186_), .A1(mai_mai_n56_), .B0(mai_mai_n23_), .Y(mai_mai_n187_));
  OAI210     m165(.A0(mai_mai_n179_), .A1(mai_mai_n56_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  INV        m166(.A(mai_mai_n128_), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n190_));
  OAI210     m168(.A0(mai_mai_n73_), .A1(mai_mai_n36_), .B0(x04), .Y(mai_mai_n191_));
  NO2        m169(.A(mai_mai_n95_), .B(x03), .Y(mai_mai_n192_));
  INV        m170(.A(mai_mai_n144_), .Y(mai_mai_n193_));
  NOi21      m171(.An(x13), .B(x04), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n193_), .B(mai_mai_n56_), .Y(mai_mai_n195_));
  OAI210     m173(.A0(mai_mai_n380_), .A1(mai_mai_n189_), .B0(mai_mai_n195_), .Y(mai_mai_n196_));
  INV        m174(.A(mai_mai_n85_), .Y(mai_mai_n197_));
  NO2        m175(.A(mai_mai_n197_), .B(x12), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n200_));
  INV        m178(.A(mai_mai_n158_), .Y(mai_mai_n201_));
  AOI210     m179(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n202_));
  NO2        m180(.A(x06), .B(x00), .Y(mai_mai_n203_));
  NA2        m181(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n204_));
  NA2        m182(.A(mai_mai_n204_), .B(x03), .Y(mai_mai_n205_));
  OA210      m183(.A0(mai_mai_n205_), .A1(mai_mai_n203_), .B0(mai_mai_n201_), .Y(mai_mai_n206_));
  NA2        m184(.A(x13), .B(mai_mai_n94_), .Y(mai_mai_n207_));
  NA3        m185(.A(mai_mai_n207_), .B(x12), .C(mai_mai_n86_), .Y(mai_mai_n208_));
  OAI210     m186(.A0(mai_mai_n206_), .A1(mai_mai_n199_), .B0(mai_mai_n208_), .Y(mai_mai_n209_));
  AOI210     m187(.A0(mai_mai_n198_), .A1(mai_mai_n196_), .B0(mai_mai_n209_), .Y(mai_mai_n210_));
  AOI210     m188(.A0(mai_mai_n210_), .A1(mai_mai_n188_), .B0(x07), .Y(mai_mai_n211_));
  NA2        m189(.A(mai_mai_n67_), .B(mai_mai_n29_), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n194_), .B(mai_mai_n166_), .Y(mai_mai_n213_));
  AOI210     m191(.A0(mai_mai_n213_), .A1(mai_mai_n136_), .B0(mai_mai_n212_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n95_), .B(x06), .Y(mai_mai_n215_));
  INV        m193(.A(mai_mai_n215_), .Y(mai_mai_n216_));
  NO2        m194(.A(x08), .B(x05), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n217_), .B(mai_mai_n202_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n218_), .B(mai_mai_n216_), .Y(mai_mai_n219_));
  NO2        m197(.A(x12), .B(x02), .Y(mai_mai_n220_));
  INV        m198(.A(mai_mai_n220_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n221_), .B(mai_mai_n197_), .Y(mai_mai_n222_));
  OA210      m200(.A0(mai_mai_n219_), .A1(mai_mai_n214_), .B0(mai_mai_n222_), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n224_), .B(x01), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n95_), .B(x04), .Y(mai_mai_n226_));
  NO3        m204(.A(mai_mai_n84_), .B(x12), .C(x03), .Y(mai_mai_n227_));
  OAI210     m205(.A0(x13), .A1(mai_mai_n77_), .B0(mai_mai_n227_), .Y(mai_mai_n228_));
  AOI210     m206(.A0(mai_mai_n170_), .A1(mai_mai_n167_), .B0(mai_mai_n96_), .Y(mai_mai_n229_));
  NOi21      m207(.An(mai_mai_n212_), .B(mai_mai_n181_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n231_));
  OAI210     m209(.A0(mai_mai_n230_), .A1(mai_mai_n229_), .B0(mai_mai_n231_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n57_), .B(x05), .Y(mai_mai_n233_));
  NO3        m211(.A(mai_mai_n233_), .B(mai_mai_n182_), .C(mai_mai_n161_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n199_), .B(mai_mai_n28_), .Y(mai_mai_n235_));
  OAI210     m213(.A0(mai_mai_n234_), .A1(mai_mai_n189_), .B0(mai_mai_n235_), .Y(mai_mai_n236_));
  NA3        m214(.A(mai_mai_n236_), .B(mai_mai_n232_), .C(mai_mai_n228_), .Y(mai_mai_n237_));
  NO3        m215(.A(mai_mai_n237_), .B(mai_mai_n223_), .C(mai_mai_n211_), .Y(mai_mai_n238_));
  OAI210     m216(.A0(mai_mai_n174_), .A1(mai_mai_n60_), .B0(mai_mai_n238_), .Y(mai02));
  NO2        m217(.A(mai_mai_n95_), .B(mai_mai_n35_), .Y(mai_mai_n240_));
  NA3        m218(.A(mai_mai_n240_), .B(x10), .C(mai_mai_n55_), .Y(mai_mai_n241_));
  OAI210     m219(.A0(x01), .A1(mai_mai_n32_), .B0(mai_mai_n241_), .Y(mai_mai_n242_));
  NA2        m220(.A(mai_mai_n242_), .B(mai_mai_n152_), .Y(mai_mai_n243_));
  INV        m221(.A(mai_mai_n152_), .Y(mai_mai_n244_));
  AOI210     m222(.A0(mai_mai_n108_), .A1(mai_mai_n79_), .B0(mai_mai_n182_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n245_), .B(mai_mai_n95_), .Y(mai_mai_n246_));
  AOI220     m224(.A0(mai_mai_n246_), .A1(mai_mai_n244_), .B0(mai_mai_n140_), .B1(mai_mai_n139_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n247_), .A1(mai_mai_n243_), .B0(mai_mai_n48_), .Y(mai_mai_n248_));
  NO2        m226(.A(x05), .B(x02), .Y(mai_mai_n249_));
  OAI210     m227(.A0(mai_mai_n177_), .A1(mai_mai_n166_), .B0(mai_mai_n249_), .Y(mai_mai_n250_));
  AOI220     m228(.A0(mai_mai_n217_), .A1(mai_mai_n57_), .B0(mai_mai_n55_), .B1(mai_mai_n36_), .Y(mai_mai_n251_));
  NOi21      m229(.An(mai_mai_n240_), .B(mai_mai_n251_), .Y(mai_mai_n252_));
  AOI210     m230(.A0(mai_mai_n194_), .A1(mai_mai_n73_), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  AOI210     m231(.A0(mai_mai_n253_), .A1(mai_mai_n250_), .B0(mai_mai_n128_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n204_), .B(mai_mai_n47_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n255_), .B(mai_mai_n192_), .Y(mai_mai_n256_));
  AN2        m234(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n257_));
  NA2        m235(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n258_));
  OA210      m236(.A0(mai_mai_n258_), .A1(x08), .B0(mai_mai_n132_), .Y(mai_mai_n259_));
  AOI210     m237(.A0(mai_mai_n259_), .A1(mai_mai_n125_), .B0(x06), .Y(mai_mai_n260_));
  OAI210     m238(.A0(mai_mai_n260_), .A1(mai_mai_n257_), .B0(mai_mai_n89_), .Y(mai_mai_n261_));
  NA3        m239(.A(mai_mai_n88_), .B(mai_mai_n76_), .C(mai_mai_n42_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n262_), .B(x04), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n218_), .B(mai_mai_n98_), .Y(mai_mai_n264_));
  AOI210     m242(.A0(mai_mai_n264_), .A1(x13), .B0(mai_mai_n263_), .Y(mai_mai_n265_));
  NA3        m243(.A(mai_mai_n265_), .B(mai_mai_n261_), .C(mai_mai_n256_), .Y(mai_mai_n266_));
  NO3        m244(.A(mai_mai_n266_), .B(mai_mai_n254_), .C(mai_mai_n248_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n127_), .B(x03), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n157_), .Y(mai_mai_n269_));
  AOI220     m247(.A0(x08), .A1(mai_mai_n269_), .B0(mai_mai_n171_), .B1(x08), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n233_), .B0(mai_mai_n268_), .Y(mai_mai_n271_));
  NA2        m249(.A(mai_mai_n271_), .B(mai_mai_n99_), .Y(mai_mai_n272_));
  NA2        m250(.A(mai_mai_n151_), .B(mai_mai_n147_), .Y(mai_mai_n273_));
  AN2        m251(.A(mai_mai_n273_), .B(mai_mai_n154_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n120_), .B(mai_mai_n28_), .Y(mai_mai_n275_));
  OAI210     m253(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n100_), .Y(mai_mai_n276_));
  NA2        m254(.A(mai_mai_n226_), .B(mai_mai_n94_), .Y(mai_mai_n277_));
  NA2        m255(.A(mai_mai_n94_), .B(mai_mai_n41_), .Y(mai_mai_n278_));
  NA3        m256(.A(mai_mai_n278_), .B(mai_mai_n277_), .C(mai_mai_n119_), .Y(mai_mai_n279_));
  NA4        m257(.A(mai_mai_n279_), .B(mai_mai_n276_), .C(mai_mai_n272_), .D(mai_mai_n48_), .Y(mai_mai_n280_));
  INV        m258(.A(mai_mai_n171_), .Y(mai_mai_n281_));
  OAI220     m259(.A0(mai_mai_n381_), .A1(mai_mai_n31_), .B0(mai_mai_n281_), .B1(mai_mai_n58_), .Y(mai_mai_n282_));
  NA2        m260(.A(mai_mai_n282_), .B(x02), .Y(mai_mai_n283_));
  INV        m261(.A(mai_mai_n200_), .Y(mai_mai_n284_));
  NA2        m262(.A(mai_mai_n168_), .B(x04), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n285_), .B(mai_mai_n284_), .Y(mai_mai_n286_));
  NO2        m264(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n287_));
  OAI210     m265(.A0(mai_mai_n287_), .A1(mai_mai_n286_), .B0(mai_mai_n89_), .Y(mai_mai_n288_));
  NO3        m266(.A(mai_mai_n168_), .B(mai_mai_n146_), .C(mai_mai_n52_), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n134_), .A1(mai_mai_n36_), .B0(mai_mai_n94_), .Y(mai_mai_n290_));
  NA2        m268(.A(mai_mai_n290_), .B(mai_mai_n289_), .Y(mai_mai_n291_));
  NA4        m269(.A(mai_mai_n291_), .B(mai_mai_n288_), .C(mai_mai_n283_), .D(x06), .Y(mai_mai_n292_));
  NA2        m270(.A(x09), .B(x03), .Y(mai_mai_n293_));
  OAI220     m271(.A0(mai_mai_n293_), .A1(mai_mai_n118_), .B0(mai_mai_n176_), .B1(mai_mai_n62_), .Y(mai_mai_n294_));
  OAI220     m272(.A0(mai_mai_n147_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n295_));
  NO3        m273(.A(mai_mai_n233_), .B(mai_mai_n117_), .C(x08), .Y(mai_mai_n296_));
  AOI210     m274(.A0(mai_mai_n295_), .A1(mai_mai_n189_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  NO3        m275(.A(mai_mai_n106_), .B(mai_mai_n118_), .C(mai_mai_n38_), .Y(mai_mai_n298_));
  INV        m276(.A(mai_mai_n298_), .Y(mai_mai_n299_));
  OAI210     m277(.A0(mai_mai_n297_), .A1(mai_mai_n28_), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  AO220      m278(.A0(mai_mai_n300_), .A1(x04), .B0(mai_mai_n294_), .B1(x05), .Y(mai_mai_n301_));
  AOI210     m279(.A0(mai_mai_n292_), .A1(mai_mai_n280_), .B0(mai_mai_n301_), .Y(mai_mai_n302_));
  OAI210     m280(.A0(mai_mai_n267_), .A1(x12), .B0(mai_mai_n302_), .Y(mai03));
  OR2        m281(.A(mai_mai_n42_), .B(mai_mai_n190_), .Y(mai_mai_n304_));
  AOI210     m282(.A0(mai_mai_n140_), .A1(mai_mai_n94_), .B0(mai_mai_n304_), .Y(mai_mai_n305_));
  OAI210     m283(.A0(mai_mai_n384_), .A1(mai_mai_n305_), .B0(x05), .Y(mai_mai_n306_));
  NA2        m284(.A(mai_mai_n304_), .B(x05), .Y(mai_mai_n307_));
  AOI210     m285(.A0(mai_mai_n125_), .A1(mai_mai_n180_), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  AOI210     m286(.A0(mai_mai_n192_), .A1(x08), .B0(mai_mai_n113_), .Y(mai_mai_n309_));
  OAI220     m287(.A0(mai_mai_n309_), .A1(mai_mai_n58_), .B0(mai_mai_n258_), .B1(mai_mai_n251_), .Y(mai_mai_n310_));
  OAI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n308_), .B0(mai_mai_n94_), .Y(mai_mai_n311_));
  AOI210     m289(.A0(mai_mai_n132_), .A1(mai_mai_n59_), .B0(mai_mai_n38_), .Y(mai_mai_n312_));
  NO2        m290(.A(mai_mai_n153_), .B(mai_mai_n121_), .Y(mai_mai_n313_));
  OAI220     m291(.A0(mai_mai_n313_), .A1(mai_mai_n37_), .B0(mai_mai_n135_), .B1(x13), .Y(mai_mai_n314_));
  OAI210     m292(.A0(mai_mai_n314_), .A1(mai_mai_n312_), .B0(x04), .Y(mai_mai_n315_));
  NO3        m293(.A(mai_mai_n278_), .B(mai_mai_n78_), .C(mai_mai_n58_), .Y(mai_mai_n316_));
  AOI210     m294(.A0(mai_mai_n163_), .A1(mai_mai_n94_), .B0(mai_mai_n132_), .Y(mai_mai_n317_));
  AN2        m295(.A(x12), .B(mai_mai_n121_), .Y(mai_mai_n318_));
  NO3        m296(.A(mai_mai_n318_), .B(mai_mai_n317_), .C(mai_mai_n316_), .Y(mai_mai_n319_));
  NA4        m297(.A(mai_mai_n319_), .B(mai_mai_n315_), .C(mai_mai_n311_), .D(mai_mai_n306_), .Y(mai04));
  NO2        m298(.A(mai_mai_n82_), .B(mai_mai_n39_), .Y(mai_mai_n321_));
  XO2        m299(.A(mai_mai_n321_), .B(mai_mai_n207_), .Y(mai05));
  NO2        m300(.A(x06), .B(mai_mai_n25_), .Y(mai_mai_n323_));
  NA3        m301(.A(mai_mai_n128_), .B(mai_mai_n120_), .C(mai_mai_n31_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n324_), .B(mai_mai_n24_), .Y(mai_mai_n325_));
  OAI210     m303(.A0(mai_mai_n325_), .A1(mai_mai_n323_), .B0(mai_mai_n94_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n26_), .A1(mai_mai_n94_), .B0(x07), .Y(mai_mai_n327_));
  INV        m305(.A(mai_mai_n327_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n145_), .B(x05), .Y(mai_mai_n329_));
  NA3        m307(.A(mai_mai_n329_), .B(mai_mai_n203_), .C(mai_mai_n197_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n331_));
  OAI210     m309(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n332_));
  OR3        m310(.A(mai_mai_n332_), .B(mai_mai_n331_), .C(mai_mai_n44_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n333_), .B(mai_mai_n330_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n334_), .B(mai_mai_n94_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n33_), .B(mai_mai_n94_), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n85_), .B0(x07), .Y(mai_mai_n337_));
  AOI220     m315(.A0(mai_mai_n337_), .A1(mai_mai_n335_), .B0(mai_mai_n328_), .B1(mai_mai_n326_), .Y(mai_mai_n338_));
  OR2        m316(.A(mai_mai_n224_), .B(mai_mai_n221_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n331_), .A1(x07), .B0(mai_mai_n127_), .Y(mai_mai_n340_));
  OR2        m318(.A(mai_mai_n340_), .B(x03), .Y(mai_mai_n341_));
  NO2        m319(.A(x07), .B(x11), .Y(mai_mai_n342_));
  NO3        m320(.A(mai_mai_n342_), .B(mai_mai_n131_), .C(mai_mai_n28_), .Y(mai_mai_n343_));
  AOI220     m321(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(mai_mai_n339_), .B1(mai_mai_n47_), .Y(mai_mai_n344_));
  NA2        m322(.A(mai_mai_n344_), .B(mai_mai_n95_), .Y(mai_mai_n345_));
  AOI210     m323(.A0(mai_mai_n285_), .A1(mai_mai_n102_), .B0(mai_mai_n220_), .Y(mai_mai_n346_));
  NOi21      m324(.An(mai_mai_n268_), .B(mai_mai_n121_), .Y(mai_mai_n347_));
  NO2        m325(.A(mai_mai_n347_), .B(mai_mai_n221_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n207_), .A1(mai_mai_n47_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NO4        m328(.A(mai_mai_n350_), .B(mai_mai_n348_), .C(mai_mai_n346_), .D(x08), .Y(mai_mai_n351_));
  NA2        m329(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n352_));
  NO2        m330(.A(mai_mai_n352_), .B(x03), .Y(mai_mai_n353_));
  NO2        m331(.A(x13), .B(x12), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n120_), .B(mai_mai_n28_), .Y(mai_mai_n355_));
  NO2        m333(.A(mai_mai_n355_), .B(mai_mai_n225_), .Y(mai_mai_n356_));
  OR3        m334(.A(mai_mai_n356_), .B(x12), .C(x03), .Y(mai_mai_n357_));
  NA3        m335(.A(mai_mai_n281_), .B(mai_mai_n114_), .C(x12), .Y(mai_mai_n358_));
  AO210      m336(.A0(mai_mai_n281_), .A1(mai_mai_n114_), .B0(mai_mai_n207_), .Y(mai_mai_n359_));
  NA4        m337(.A(mai_mai_n359_), .B(mai_mai_n358_), .C(mai_mai_n357_), .D(x08), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n354_), .A1(mai_mai_n353_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  AOI210     m339(.A0(mai_mai_n351_), .A1(mai_mai_n345_), .B0(mai_mai_n361_), .Y(mai_mai_n362_));
  INV        m340(.A(x07), .Y(mai_mai_n363_));
  OAI220     m341(.A0(mai_mai_n363_), .A1(x02), .B0(mai_mai_n131_), .B1(mai_mai_n43_), .Y(mai_mai_n364_));
  OAI210     m342(.A0(mai_mai_n364_), .A1(x11), .B0(mai_mai_n162_), .Y(mai_mai_n365_));
  NA3        m343(.A(mai_mai_n356_), .B(mai_mai_n347_), .C(mai_mai_n277_), .Y(mai_mai_n366_));
  INV        m344(.A(x14), .Y(mai_mai_n367_));
  NO3        m345(.A(mai_mai_n268_), .B(mai_mai_n98_), .C(x11), .Y(mai_mai_n368_));
  NO2        m346(.A(mai_mai_n368_), .B(mai_mai_n367_), .Y(mai_mai_n369_));
  NA3        m347(.A(mai_mai_n369_), .B(mai_mai_n366_), .C(mai_mai_n365_), .Y(mai_mai_n370_));
  AOI210     m348(.A0(mai_mai_n336_), .A1(mai_mai_n60_), .B0(mai_mai_n355_), .Y(mai_mai_n371_));
  NOi21      m349(.An(mai_mai_n226_), .B(mai_mai_n135_), .Y(mai_mai_n372_));
  NO2        m350(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n373_));
  OAI210     m351(.A0(mai_mai_n373_), .A1(mai_mai_n372_), .B0(mai_mai_n94_), .Y(mai_mai_n374_));
  OAI210     m352(.A0(mai_mai_n371_), .A1(mai_mai_n84_), .B0(mai_mai_n374_), .Y(mai_mai_n375_));
  NO4        m353(.A(mai_mai_n375_), .B(mai_mai_n370_), .C(mai_mai_n362_), .D(mai_mai_n338_), .Y(mai06));
  INV        m354(.A(x07), .Y(mai_mai_n379_));
  INV        m355(.A(mai_mai_n192_), .Y(mai_mai_n380_));
  INV        m356(.A(x05), .Y(mai_mai_n381_));
  INV        m357(.A(x05), .Y(mai_mai_n382_));
  INV        m358(.A(x11), .Y(mai_mai_n383_));
  INV        m359(.A(mai_mai_n285_), .Y(mai_mai_n384_));
  INV        m360(.A(mai_mai_n67_), .Y(mai_mai_n385_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO2        u027(.A(men_men_n49_), .B(x11), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  INV        u030(.A(men_men_n52_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  INV        u039(.A(men_men_n59_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  OAI210     u042(.A0(men_men_n64_), .A1(men_men_n62_), .B0(men_men_n60_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n59_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  INV        u050(.A(men_men_n72_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n74_));
  OAI210     u052(.A0(men_men_n73_), .A1(x07), .B0(x03), .Y(men_men_n75_));
  NOi31      u053(.An(x08), .B(x04), .C(x00), .Y(men_men_n76_));
  NO2        u054(.A(x10), .B(x09), .Y(men_men_n77_));
  NO2        u055(.A(x09), .B(men_men_n41_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n78_), .B(men_men_n36_), .Y(men_men_n79_));
  OAI210     u057(.A0(men_men_n78_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n80_));
  AOI210     u058(.A0(men_men_n79_), .A1(men_men_n48_), .B0(men_men_n80_), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n36_), .B(x00), .Y(men_men_n82_));
  NO2        u060(.A(x08), .B(x01), .Y(men_men_n83_));
  OAI210     u061(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n35_), .Y(men_men_n84_));
  NO2        u062(.A(men_men_n84_), .B(men_men_n81_), .Y(men_men_n85_));
  AN2        u063(.A(men_men_n85_), .B(men_men_n75_), .Y(men_men_n86_));
  INV        u064(.A(men_men_n84_), .Y(men_men_n87_));
  NO2        u065(.A(x06), .B(x05), .Y(men_men_n88_));
  NA2        u066(.A(x11), .B(x00), .Y(men_men_n89_));
  NO2        u067(.A(x11), .B(men_men_n47_), .Y(men_men_n90_));
  NOi21      u068(.An(men_men_n89_), .B(men_men_n90_), .Y(men_men_n91_));
  NOi21      u069(.An(x01), .B(x10), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n93_));
  NO3        u071(.A(men_men_n93_), .B(men_men_n92_), .C(x06), .Y(men_men_n94_));
  NA2        u072(.A(men_men_n94_), .B(men_men_n27_), .Y(men_men_n95_));
  OAI210     u073(.A0(men_men_n422_), .A1(x07), .B0(men_men_n95_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n86_), .C(men_men_n69_), .Y(men01));
  INV        u075(.A(x12), .Y(men_men_n98_));
  INV        u076(.A(x13), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n88_), .B(x01), .Y(men_men_n100_));
  NA2        u078(.A(men_men_n100_), .B(men_men_n70_), .Y(men_men_n101_));
  NA2        u079(.A(x08), .B(x04), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n102_), .B(men_men_n57_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n103_), .B(men_men_n101_), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n92_), .B(men_men_n28_), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n105_), .B(men_men_n71_), .Y(men_men_n106_));
  NO2        u084(.A(x10), .B(x01), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n29_), .B(x00), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NA2        u087(.A(x04), .B(men_men_n28_), .Y(men_men_n110_));
  NO3        u088(.A(men_men_n110_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n111_));
  AOI210     u089(.A0(men_men_n111_), .A1(men_men_n109_), .B0(men_men_n106_), .Y(men_men_n112_));
  AOI210     u090(.A0(men_men_n112_), .A1(men_men_n104_), .B0(men_men_n99_), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n56_), .B(x05), .Y(men_men_n114_));
  NOi21      u092(.An(men_men_n114_), .B(men_men_n58_), .Y(men_men_n115_));
  NO2        u093(.A(men_men_n99_), .B(men_men_n36_), .Y(men_men_n116_));
  NA3        u094(.A(men_men_n116_), .B(men_men_n423_), .C(x06), .Y(men_men_n117_));
  INV        u095(.A(men_men_n117_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n83_), .B(x13), .Y(men_men_n119_));
  NA2        u097(.A(x09), .B(men_men_n35_), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NA2        u099(.A(x13), .B(men_men_n35_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(x05), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n123_), .B(men_men_n121_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n125_));
  AOI210     u103(.A0(men_men_n57_), .A1(men_men_n79_), .B0(men_men_n115_), .Y(men_men_n126_));
  AOI210     u104(.A0(men_men_n126_), .A1(men_men_n124_), .B0(men_men_n72_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n128_));
  NA2        u106(.A(x10), .B(men_men_n57_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n129_), .B(men_men_n128_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n51_), .B(x05), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n36_), .B(x04), .Y(men_men_n132_));
  NA3        u110(.A(men_men_n132_), .B(men_men_n131_), .C(x13), .Y(men_men_n133_));
  NO3        u111(.A(men_men_n125_), .B(men_men_n78_), .C(men_men_n36_), .Y(men_men_n134_));
  NO2        u112(.A(men_men_n60_), .B(x05), .Y(men_men_n135_));
  NOi41      u113(.An(men_men_n133_), .B(men_men_n135_), .C(men_men_n134_), .D(men_men_n130_), .Y(men_men_n136_));
  NO3        u114(.A(men_men_n136_), .B(x06), .C(x03), .Y(men_men_n137_));
  NO4        u115(.A(men_men_n137_), .B(men_men_n127_), .C(men_men_n118_), .D(men_men_n113_), .Y(men_men_n138_));
  NA2        u116(.A(x13), .B(men_men_n36_), .Y(men_men_n139_));
  OAI210     u117(.A0(men_men_n83_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n140_));
  INV        u118(.A(men_men_n139_), .Y(men_men_n141_));
  NO2        u119(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n142_));
  OA210      u120(.A0(x00), .A1(men_men_n77_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u121(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n29_), .B(x06), .Y(men_men_n145_));
  AN2        u123(.A(men_men_n143_), .B(men_men_n141_), .Y(men_men_n146_));
  NO2        u124(.A(x09), .B(x05), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n147_), .B(men_men_n47_), .Y(men_men_n148_));
  AOI210     u126(.A0(men_men_n148_), .A1(men_men_n109_), .B0(men_men_n49_), .Y(men_men_n149_));
  NA2        u127(.A(x09), .B(x00), .Y(men_men_n150_));
  NA2        u128(.A(men_men_n114_), .B(men_men_n150_), .Y(men_men_n151_));
  NO3        u129(.A(men_men_n424_), .B(men_men_n149_), .C(men_men_n146_), .Y(men_men_n152_));
  NO2        u130(.A(x03), .B(x02), .Y(men_men_n153_));
  NA2        u131(.A(men_men_n84_), .B(men_men_n99_), .Y(men_men_n154_));
  OAI210     u132(.A0(men_men_n154_), .A1(men_men_n115_), .B0(men_men_n153_), .Y(men_men_n155_));
  OA210      u133(.A0(men_men_n152_), .A1(x11), .B0(men_men_n155_), .Y(men_men_n156_));
  OAI210     u134(.A0(men_men_n138_), .A1(men_men_n23_), .B0(men_men_n156_), .Y(men_men_n157_));
  NA2        u135(.A(men_men_n109_), .B(men_men_n40_), .Y(men_men_n158_));
  NAi21      u136(.An(x06), .B(x10), .Y(men_men_n159_));
  NOi21      u137(.An(x01), .B(x13), .Y(men_men_n160_));
  NA2        u138(.A(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  OR2        u139(.A(men_men_n161_), .B(x08), .Y(men_men_n162_));
  AOI210     u140(.A0(men_men_n162_), .A1(men_men_n158_), .B0(men_men_n41_), .Y(men_men_n163_));
  NO2        u141(.A(men_men_n29_), .B(x03), .Y(men_men_n164_));
  NA2        u142(.A(men_men_n99_), .B(x01), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n165_), .B(x08), .Y(men_men_n166_));
  OAI210     u144(.A0(x05), .A1(men_men_n166_), .B0(men_men_n51_), .Y(men_men_n167_));
  AOI210     u145(.A0(men_men_n167_), .A1(men_men_n164_), .B0(men_men_n48_), .Y(men_men_n168_));
  AOI210     u146(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n169_));
  OAI210     u147(.A0(men_men_n168_), .A1(men_men_n163_), .B0(men_men_n169_), .Y(men_men_n170_));
  NA2        u148(.A(x04), .B(x02), .Y(men_men_n171_));
  NA2        u149(.A(x10), .B(x05), .Y(men_men_n172_));
  NA2        u150(.A(x09), .B(x06), .Y(men_men_n173_));
  NO2        u151(.A(x09), .B(x01), .Y(men_men_n174_));
  NO3        u152(.A(men_men_n174_), .B(men_men_n107_), .C(men_men_n31_), .Y(men_men_n175_));
  NA2        u153(.A(men_men_n175_), .B(x00), .Y(men_men_n176_));
  NO2        u154(.A(men_men_n114_), .B(x08), .Y(men_men_n177_));
  NA3        u155(.A(men_men_n160_), .B(men_men_n159_), .C(men_men_n51_), .Y(men_men_n178_));
  NA2        u156(.A(men_men_n92_), .B(x05), .Y(men_men_n179_));
  OAI210     u157(.A0(men_men_n179_), .A1(men_men_n116_), .B0(men_men_n178_), .Y(men_men_n180_));
  AOI210     u158(.A0(men_men_n177_), .A1(x06), .B0(men_men_n180_), .Y(men_men_n181_));
  OAI210     u159(.A0(men_men_n181_), .A1(x11), .B0(men_men_n176_), .Y(men_men_n182_));
  NAi21      u160(.An(men_men_n171_), .B(men_men_n182_), .Y(men_men_n183_));
  INV        u161(.A(men_men_n25_), .Y(men_men_n184_));
  NAi21      u162(.An(x13), .B(x00), .Y(men_men_n185_));
  AOI210     u163(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n185_), .Y(men_men_n186_));
  AOI220     u164(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n187_));
  OAI210     u165(.A0(men_men_n172_), .A1(men_men_n35_), .B0(men_men_n187_), .Y(men_men_n188_));
  AN2        u166(.A(men_men_n188_), .B(men_men_n186_), .Y(men_men_n189_));
  NO2        u167(.A(men_men_n185_), .B(men_men_n36_), .Y(men_men_n190_));
  INV        u168(.A(men_men_n190_), .Y(men_men_n191_));
  OAI210     u169(.A0(men_men_n191_), .A1(men_men_n173_), .B0(men_men_n72_), .Y(men_men_n192_));
  OAI210     u170(.A0(men_men_n192_), .A1(men_men_n189_), .B0(men_men_n184_), .Y(men_men_n193_));
  NOi21      u171(.An(x09), .B(x00), .Y(men_men_n194_));
  NO3        u172(.A(men_men_n82_), .B(men_men_n194_), .C(men_men_n47_), .Y(men_men_n195_));
  NA2        u173(.A(men_men_n195_), .B(men_men_n129_), .Y(men_men_n196_));
  NA2        u174(.A(x10), .B(x08), .Y(men_men_n197_));
  INV        u175(.A(men_men_n197_), .Y(men_men_n198_));
  NA2        u176(.A(x06), .B(x05), .Y(men_men_n199_));
  OAI210     u177(.A0(men_men_n199_), .A1(men_men_n35_), .B0(men_men_n98_), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n198_), .A1(men_men_n58_), .B0(men_men_n200_), .Y(men_men_n201_));
  NA2        u179(.A(men_men_n201_), .B(men_men_n196_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n99_), .B(x12), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n203_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n92_), .B(men_men_n51_), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n206_));
  NA2        u184(.A(men_men_n206_), .B(x02), .Y(men_men_n207_));
  NO2        u185(.A(men_men_n207_), .B(men_men_n205_), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n204_), .A1(men_men_n202_), .B0(men_men_n208_), .Y(men_men_n209_));
  NA4        u187(.A(men_men_n209_), .B(men_men_n193_), .C(men_men_n183_), .D(men_men_n170_), .Y(men_men_n210_));
  AOI210     u188(.A0(men_men_n157_), .A1(men_men_n98_), .B0(men_men_n210_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n212_));
  NA2        u190(.A(men_men_n212_), .B(men_men_n140_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n128_), .B(x06), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n214_), .A1(men_men_n213_), .B0(men_men_n215_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n216_), .B(x12), .Y(men_men_n217_));
  INV        u195(.A(men_men_n76_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n161_), .B(men_men_n57_), .Y(men_men_n219_));
  INV        u197(.A(men_men_n219_), .Y(men_men_n220_));
  NA2        u198(.A(men_men_n159_), .B(x02), .Y(men_men_n221_));
  AOI210     u199(.A0(men_men_n221_), .A1(men_men_n220_), .B0(men_men_n23_), .Y(men_men_n222_));
  OAI210     u200(.A0(men_men_n217_), .A1(men_men_n57_), .B0(men_men_n222_), .Y(men_men_n223_));
  INV        u201(.A(men_men_n145_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n51_), .B(x03), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n78_), .A1(men_men_n36_), .B0(men_men_n120_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n99_), .B(x03), .Y(men_men_n227_));
  AOI220     u205(.A0(men_men_n227_), .A1(men_men_n226_), .B0(men_men_n76_), .B1(men_men_n225_), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n32_), .B(x06), .Y(men_men_n229_));
  INV        u207(.A(men_men_n159_), .Y(men_men_n230_));
  NOi21      u208(.An(x13), .B(x04), .Y(men_men_n231_));
  NO3        u209(.A(men_men_n231_), .B(men_men_n76_), .C(men_men_n194_), .Y(men_men_n232_));
  NO2        u210(.A(men_men_n232_), .B(x05), .Y(men_men_n233_));
  AOI220     u211(.A0(men_men_n233_), .A1(men_men_n229_), .B0(men_men_n230_), .B1(men_men_n57_), .Y(men_men_n234_));
  OAI210     u212(.A0(men_men_n228_), .A1(men_men_n224_), .B0(men_men_n234_), .Y(men_men_n235_));
  INV        u213(.A(men_men_n90_), .Y(men_men_n236_));
  NO2        u214(.A(men_men_n236_), .B(x12), .Y(men_men_n237_));
  NA2        u215(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n238_));
  NO2        u216(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n239_));
  OAI210     u217(.A0(men_men_n239_), .A1(men_men_n188_), .B0(men_men_n186_), .Y(men_men_n240_));
  OAI210     u218(.A0(men_men_n102_), .A1(men_men_n150_), .B0(men_men_n72_), .Y(men_men_n241_));
  INV        u219(.A(men_men_n241_), .Y(men_men_n242_));
  INV        u220(.A(x03), .Y(men_men_n243_));
  OA210      u221(.A0(men_men_n243_), .A1(men_men_n242_), .B0(men_men_n240_), .Y(men_men_n244_));
  NA2        u222(.A(x13), .B(men_men_n98_), .Y(men_men_n245_));
  NA3        u223(.A(men_men_n245_), .B(men_men_n200_), .C(men_men_n91_), .Y(men_men_n246_));
  OAI210     u224(.A0(men_men_n244_), .A1(men_men_n238_), .B0(men_men_n246_), .Y(men_men_n247_));
  AOI210     u225(.A0(men_men_n237_), .A1(men_men_n235_), .B0(men_men_n247_), .Y(men_men_n248_));
  AOI210     u226(.A0(men_men_n248_), .A1(men_men_n223_), .B0(x07), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n99_), .B(x06), .Y(men_men_n251_));
  NO2        u229(.A(x08), .B(x05), .Y(men_men_n252_));
  NO2        u230(.A(x12), .B(x02), .Y(men_men_n253_));
  INV        u231(.A(men_men_n253_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n254_), .B(men_men_n236_), .Y(men_men_n255_));
  OA210      u233(.A0(x13), .A1(men_men_n76_), .B0(men_men_n255_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n257_));
  NO2        u235(.A(men_men_n257_), .B(x01), .Y(men_men_n258_));
  NOi21      u236(.An(men_men_n83_), .B(men_men_n120_), .Y(men_men_n259_));
  NO2        u237(.A(men_men_n259_), .B(men_men_n258_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n260_), .A1(men_men_n133_), .B0(men_men_n29_), .Y(men_men_n261_));
  NA2        u239(.A(men_men_n251_), .B(men_men_n226_), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n99_), .B(x04), .Y(men_men_n263_));
  NA2        u241(.A(men_men_n263_), .B(men_men_n28_), .Y(men_men_n264_));
  OAI210     u242(.A0(men_men_n264_), .A1(men_men_n119_), .B0(men_men_n262_), .Y(men_men_n265_));
  NO3        u243(.A(men_men_n89_), .B(x12), .C(x03), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n265_), .A1(men_men_n261_), .B0(men_men_n266_), .Y(men_men_n267_));
  AOI210     u245(.A0(men_men_n205_), .A1(men_men_n199_), .B0(men_men_n102_), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n25_), .B(x00), .Y(men_men_n269_));
  NA2        u247(.A(men_men_n268_), .B(men_men_n269_), .Y(men_men_n270_));
  NA2        u248(.A(men_men_n270_), .B(men_men_n267_), .Y(men_men_n271_));
  NO3        u249(.A(men_men_n271_), .B(men_men_n256_), .C(men_men_n249_), .Y(men_men_n272_));
  OAI210     u250(.A0(men_men_n211_), .A1(men_men_n61_), .B0(men_men_n272_), .Y(men02));
  AOI210     u251(.A0(men_men_n139_), .A1(men_men_n84_), .B0(men_men_n131_), .Y(men_men_n274_));
  NOi21      u252(.An(men_men_n232_), .B(men_men_n174_), .Y(men_men_n275_));
  NA3        u253(.A(x13), .B(men_men_n198_), .C(men_men_n56_), .Y(men_men_n276_));
  OAI210     u254(.A0(men_men_n275_), .A1(men_men_n32_), .B0(men_men_n276_), .Y(men_men_n277_));
  OAI210     u255(.A0(men_men_n277_), .A1(men_men_n274_), .B0(men_men_n172_), .Y(men_men_n278_));
  INV        u256(.A(men_men_n172_), .Y(men_men_n279_));
  NO2        u257(.A(men_men_n84_), .B(men_men_n51_), .Y(men_men_n280_));
  AOI220     u258(.A0(men_men_n280_), .A1(men_men_n279_), .B0(men_men_n154_), .B1(men_men_n153_), .Y(men_men_n281_));
  AOI210     u259(.A0(men_men_n281_), .A1(men_men_n278_), .B0(men_men_n48_), .Y(men_men_n282_));
  NO2        u260(.A(x05), .B(x02), .Y(men_men_n283_));
  OAI210     u261(.A0(men_men_n213_), .A1(men_men_n194_), .B0(men_men_n283_), .Y(men_men_n284_));
  AOI220     u262(.A0(men_men_n252_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n285_));
  NOi21      u263(.An(x13), .B(men_men_n285_), .Y(men_men_n286_));
  AOI210     u264(.A0(men_men_n231_), .A1(men_men_n78_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI210     u265(.A0(men_men_n287_), .A1(men_men_n284_), .B0(men_men_n145_), .Y(men_men_n288_));
  NAi21      u266(.An(men_men_n233_), .B(men_men_n228_), .Y(men_men_n289_));
  NO2        u267(.A(x10), .B(men_men_n47_), .Y(men_men_n290_));
  NA2        u268(.A(men_men_n290_), .B(men_men_n289_), .Y(men_men_n291_));
  AN2        u269(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n292_));
  OAI210     u270(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n293_));
  NA2        u271(.A(x13), .B(men_men_n28_), .Y(men_men_n294_));
  BUFFER     u272(.A(men_men_n148_), .Y(men_men_n295_));
  AOI210     u273(.A0(men_men_n295_), .A1(men_men_n140_), .B0(men_men_n293_), .Y(men_men_n296_));
  OAI210     u274(.A0(men_men_n296_), .A1(men_men_n292_), .B0(men_men_n93_), .Y(men_men_n297_));
  NA3        u275(.A(men_men_n93_), .B(men_men_n83_), .C(men_men_n225_), .Y(men_men_n298_));
  NA3        u276(.A(men_men_n92_), .B(men_men_n82_), .C(men_men_n42_), .Y(men_men_n299_));
  AOI210     u277(.A0(men_men_n299_), .A1(men_men_n298_), .B0(x04), .Y(men_men_n300_));
  INV        u278(.A(men_men_n153_), .Y(men_men_n301_));
  NO2        u279(.A(men_men_n301_), .B(men_men_n130_), .Y(men_men_n302_));
  AOI210     u280(.A0(men_men_n302_), .A1(x13), .B0(men_men_n300_), .Y(men_men_n303_));
  NA3        u281(.A(men_men_n303_), .B(men_men_n297_), .C(men_men_n291_), .Y(men_men_n304_));
  NO3        u282(.A(men_men_n304_), .B(men_men_n288_), .C(men_men_n282_), .Y(men_men_n305_));
  NA2        u283(.A(men_men_n144_), .B(x03), .Y(men_men_n306_));
  OAI210     u284(.A0(men_men_n185_), .A1(men_men_n51_), .B0(men_men_n306_), .Y(men_men_n307_));
  NA2        u285(.A(men_men_n307_), .B(men_men_n107_), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n56_), .A1(men_men_n177_), .B0(men_men_n108_), .Y(men_men_n309_));
  NA2        u287(.A(men_men_n263_), .B(men_men_n98_), .Y(men_men_n310_));
  NA2        u288(.A(men_men_n98_), .B(men_men_n41_), .Y(men_men_n311_));
  NA3        u289(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n130_), .Y(men_men_n312_));
  NA4        u290(.A(men_men_n312_), .B(men_men_n309_), .C(men_men_n308_), .D(men_men_n48_), .Y(men_men_n313_));
  INV        u291(.A(men_men_n206_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n32_), .B(x05), .Y(men_men_n315_));
  INV        u293(.A(men_men_n315_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n316_), .B(x02), .Y(men_men_n317_));
  NA2        u295(.A(men_men_n203_), .B(x04), .Y(men_men_n318_));
  NO2        u296(.A(men_men_n318_), .B(men_men_n36_), .Y(men_men_n319_));
  NO3        u297(.A(men_men_n187_), .B(x13), .C(men_men_n31_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n320_), .A1(men_men_n319_), .B0(men_men_n93_), .Y(men_men_n321_));
  NO3        u299(.A(men_men_n203_), .B(men_men_n164_), .C(men_men_n52_), .Y(men_men_n322_));
  OAI210     u300(.A0(x12), .A1(men_men_n195_), .B0(men_men_n322_), .Y(men_men_n323_));
  NA4        u301(.A(men_men_n323_), .B(men_men_n321_), .C(men_men_n317_), .D(x06), .Y(men_men_n324_));
  INV        u302(.A(x03), .Y(men_men_n325_));
  OAI220     u303(.A0(men_men_n325_), .A1(men_men_n129_), .B0(men_men_n212_), .B1(men_men_n63_), .Y(men_men_n326_));
  NO2        u304(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n322_), .B(men_men_n327_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n145_), .A1(men_men_n28_), .B0(men_men_n328_), .Y(men_men_n329_));
  AO220      u307(.A0(men_men_n329_), .A1(x04), .B0(men_men_n326_), .B1(x05), .Y(men_men_n330_));
  AOI210     u308(.A0(men_men_n324_), .A1(men_men_n313_), .B0(men_men_n330_), .Y(men_men_n331_));
  OAI210     u309(.A0(men_men_n305_), .A1(x12), .B0(men_men_n331_), .Y(men03));
  OR2        u310(.A(men_men_n42_), .B(men_men_n225_), .Y(men_men_n333_));
  AOI210     u311(.A0(men_men_n154_), .A1(men_men_n98_), .B0(men_men_n333_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n203_), .B(men_men_n153_), .Y(men_men_n335_));
  NA2        u313(.A(men_men_n335_), .B(men_men_n207_), .Y(men_men_n336_));
  OAI210     u314(.A0(men_men_n336_), .A1(men_men_n334_), .B0(x05), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n333_), .B(x05), .Y(men_men_n338_));
  AOI210     u316(.A0(men_men_n140_), .A1(men_men_n218_), .B0(men_men_n338_), .Y(men_men_n339_));
  AOI210     u317(.A0(men_men_n227_), .A1(men_men_n79_), .B0(men_men_n123_), .Y(men_men_n340_));
  OAI220     u318(.A0(men_men_n340_), .A1(men_men_n59_), .B0(men_men_n294_), .B1(men_men_n285_), .Y(men_men_n341_));
  OAI210     u319(.A0(men_men_n341_), .A1(men_men_n339_), .B0(men_men_n98_), .Y(men_men_n342_));
  AOI210     u320(.A0(men_men_n148_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n343_));
  NO2        u321(.A(men_men_n174_), .B(men_men_n135_), .Y(men_men_n344_));
  OAI220     u322(.A0(men_men_n344_), .A1(men_men_n37_), .B0(men_men_n151_), .B1(x13), .Y(men_men_n345_));
  OAI210     u323(.A0(men_men_n345_), .A1(men_men_n343_), .B0(x04), .Y(men_men_n346_));
  AOI210     u324(.A0(men_men_n191_), .A1(men_men_n98_), .B0(men_men_n148_), .Y(men_men_n347_));
  OA210      u325(.A0(men_men_n166_), .A1(x12), .B0(men_men_n135_), .Y(men_men_n348_));
  NO2        u326(.A(men_men_n348_), .B(men_men_n347_), .Y(men_men_n349_));
  NA4        u327(.A(men_men_n349_), .B(men_men_n346_), .C(men_men_n342_), .D(men_men_n337_), .Y(men04));
  NO2        u328(.A(men_men_n87_), .B(men_men_n39_), .Y(men_men_n351_));
  XO2        u329(.A(men_men_n351_), .B(men_men_n245_), .Y(men05));
  AOI210     u330(.A0(men_men_n71_), .A1(men_men_n52_), .B0(men_men_n215_), .Y(men_men_n353_));
  NO2        u331(.A(men_men_n353_), .B(men_men_n25_), .Y(men_men_n354_));
  AOI210     u332(.A0(men_men_n230_), .A1(men_men_n57_), .B0(men_men_n88_), .Y(men_men_n355_));
  NO2        u333(.A(men_men_n355_), .B(men_men_n24_), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n356_), .A1(men_men_n354_), .B0(men_men_n98_), .Y(men_men_n357_));
  NA2        u335(.A(x11), .B(men_men_n31_), .Y(men_men_n358_));
  NA2        u336(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n359_));
  NA2        u337(.A(men_men_n250_), .B(x03), .Y(men_men_n360_));
  OAI220     u338(.A0(men_men_n360_), .A1(men_men_n359_), .B0(men_men_n358_), .B1(men_men_n80_), .Y(men_men_n361_));
  OAI210     u339(.A0(men_men_n26_), .A1(men_men_n98_), .B0(x07), .Y(men_men_n362_));
  AOI210     u340(.A0(men_men_n361_), .A1(x06), .B0(men_men_n362_), .Y(men_men_n363_));
  AOI220     u341(.A0(men_men_n80_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n364_));
  NO3        u342(.A(men_men_n364_), .B(men_men_n23_), .C(x00), .Y(men_men_n365_));
  NA2        u343(.A(men_men_n70_), .B(x02), .Y(men_men_n366_));
  AOI210     u344(.A0(men_men_n366_), .A1(men_men_n360_), .B0(men_men_n251_), .Y(men_men_n367_));
  OR2        u345(.A(men_men_n367_), .B(men_men_n238_), .Y(men_men_n368_));
  NO2        u346(.A(men_men_n23_), .B(x10), .Y(men_men_n369_));
  OAI210     u347(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n370_));
  OR3        u348(.A(men_men_n370_), .B(men_men_n369_), .C(men_men_n44_), .Y(men_men_n371_));
  NA2        u349(.A(men_men_n371_), .B(men_men_n368_), .Y(men_men_n372_));
  OAI210     u350(.A0(men_men_n372_), .A1(men_men_n365_), .B0(men_men_n98_), .Y(men_men_n373_));
  AOI210     u351(.A0(x12), .A1(men_men_n90_), .B0(x07), .Y(men_men_n374_));
  AOI220     u352(.A0(men_men_n374_), .A1(men_men_n373_), .B0(men_men_n363_), .B1(men_men_n357_), .Y(men_men_n375_));
  NA3        u353(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n376_));
  AO210      u354(.A0(men_men_n376_), .A1(men_men_n257_), .B0(men_men_n254_), .Y(men_men_n377_));
  AOI210     u355(.A0(men_men_n369_), .A1(men_men_n74_), .B0(men_men_n144_), .Y(men_men_n378_));
  OR2        u356(.A(men_men_n378_), .B(x03), .Y(men_men_n379_));
  NA2        u357(.A(men_men_n327_), .B(men_men_n61_), .Y(men_men_n380_));
  NO2        u358(.A(men_men_n380_), .B(x11), .Y(men_men_n381_));
  NO3        u359(.A(men_men_n381_), .B(men_men_n147_), .C(men_men_n28_), .Y(men_men_n382_));
  AOI220     u360(.A0(men_men_n382_), .A1(men_men_n379_), .B0(men_men_n377_), .B1(men_men_n47_), .Y(men_men_n383_));
  NO4        u361(.A(men_men_n311_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n384_));
  OAI210     u362(.A0(men_men_n384_), .A1(men_men_n383_), .B0(men_men_n99_), .Y(men_men_n385_));
  AOI210     u363(.A0(men_men_n318_), .A1(men_men_n110_), .B0(men_men_n253_), .Y(men_men_n386_));
  NOi21      u364(.An(men_men_n306_), .B(men_men_n135_), .Y(men_men_n387_));
  NO2        u365(.A(men_men_n386_), .B(x08), .Y(men_men_n388_));
  AOI210     u366(.A0(men_men_n369_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n389_));
  NA2        u367(.A(x09), .B(men_men_n41_), .Y(men_men_n390_));
  OAI220     u368(.A0(men_men_n390_), .A1(men_men_n389_), .B0(men_men_n358_), .B1(men_men_n66_), .Y(men_men_n391_));
  NO2        u369(.A(x13), .B(x12), .Y(men_men_n392_));
  NO2        u370(.A(men_men_n131_), .B(men_men_n28_), .Y(men_men_n393_));
  NO2        u371(.A(men_men_n393_), .B(men_men_n258_), .Y(men_men_n394_));
  OR3        u372(.A(men_men_n394_), .B(x12), .C(x03), .Y(men_men_n395_));
  NA3        u373(.A(men_men_n314_), .B(men_men_n125_), .C(x12), .Y(men_men_n396_));
  AO210      u374(.A0(men_men_n314_), .A1(men_men_n125_), .B0(men_men_n245_), .Y(men_men_n397_));
  NA4        u375(.A(men_men_n397_), .B(men_men_n396_), .C(men_men_n395_), .D(x08), .Y(men_men_n398_));
  AOI210     u376(.A0(men_men_n392_), .A1(men_men_n391_), .B0(men_men_n398_), .Y(men_men_n399_));
  AOI210     u377(.A0(men_men_n388_), .A1(men_men_n385_), .B0(men_men_n399_), .Y(men_men_n400_));
  OAI210     u378(.A0(men_men_n380_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n279_), .B(x07), .Y(men_men_n402_));
  OAI220     u380(.A0(men_men_n402_), .A1(men_men_n359_), .B0(men_men_n147_), .B1(men_men_n43_), .Y(men_men_n403_));
  OAI210     u381(.A0(men_men_n403_), .A1(men_men_n401_), .B0(men_men_n190_), .Y(men_men_n404_));
  NA3        u382(.A(men_men_n394_), .B(men_men_n387_), .C(men_men_n310_), .Y(men_men_n405_));
  INV        u383(.A(x14), .Y(men_men_n406_));
  NO3        u384(.A(men_men_n306_), .B(men_men_n105_), .C(x11), .Y(men_men_n407_));
  NO3        u385(.A(men_men_n165_), .B(men_men_n74_), .C(men_men_n57_), .Y(men_men_n408_));
  NO3        u386(.A(men_men_n376_), .B(men_men_n311_), .C(men_men_n185_), .Y(men_men_n409_));
  NO4        u387(.A(men_men_n409_), .B(men_men_n408_), .C(men_men_n407_), .D(men_men_n406_), .Y(men_men_n410_));
  NA3        u388(.A(men_men_n410_), .B(men_men_n405_), .C(men_men_n404_), .Y(men_men_n411_));
  AOI220     u389(.A0(x12), .A1(men_men_n61_), .B0(men_men_n393_), .B1(men_men_n164_), .Y(men_men_n412_));
  NOi21      u390(.An(men_men_n263_), .B(men_men_n151_), .Y(men_men_n413_));
  NO3        u391(.A(men_men_n128_), .B(men_men_n24_), .C(x06), .Y(men_men_n414_));
  AOI210     u392(.A0(men_men_n269_), .A1(men_men_n230_), .B0(men_men_n414_), .Y(men_men_n415_));
  OAI210     u393(.A0(men_men_n44_), .A1(x04), .B0(men_men_n415_), .Y(men_men_n416_));
  OAI210     u394(.A0(men_men_n416_), .A1(men_men_n413_), .B0(men_men_n98_), .Y(men_men_n417_));
  OAI210     u395(.A0(men_men_n412_), .A1(men_men_n89_), .B0(men_men_n417_), .Y(men_men_n418_));
  NO4        u396(.A(men_men_n418_), .B(men_men_n411_), .C(men_men_n400_), .D(men_men_n375_), .Y(men06));
  INV        u397(.A(men_men_n91_), .Y(men_men_n422_));
  INV        u398(.A(x02), .Y(men_men_n423_));
  INV        u399(.A(men_men_n145_), .Y(men_men_n424_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule