//Benchmark atmr_9sym_175_0.25

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NOi21      m013(.An(i_8_), .B(i_6_), .Y(mai_mai_n24_));
  INV        m014(.A(mai_mai_n20_), .Y(mai_mai_n25_));
  INV        m015(.A(i_2_), .Y(mai_mai_n26_));
  NOi21      m016(.An(i_5_), .B(i_0_), .Y(mai_mai_n27_));
  NOi21      m017(.An(i_6_), .B(i_8_), .Y(mai_mai_n28_));
  NOi21      m018(.An(i_7_), .B(i_1_), .Y(mai_mai_n29_));
  NOi21      m019(.An(i_5_), .B(i_6_), .Y(mai_mai_n30_));
  AOI220     m020(.A0(mai_mai_n30_), .A1(mai_mai_n29_), .B0(mai_mai_n28_), .B1(mai_mai_n27_), .Y(mai_mai_n31_));
  NO3        m021(.A(mai_mai_n31_), .B(mai_mai_n26_), .C(i_4_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_0_), .B(i_4_), .Y(mai_mai_n33_));
  XO2        m023(.A(i_1_), .B(i_3_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_7_), .B(i_5_), .Y(mai_mai_n35_));
  AN3        m025(.A(mai_mai_n35_), .B(mai_mai_n34_), .C(mai_mai_n33_), .Y(mai_mai_n36_));
  INV        m026(.A(i_1_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_3_), .B(i_0_), .Y(mai_mai_n38_));
  NO2        m028(.A(mai_mai_n36_), .B(mai_mai_n32_), .Y(mai_mai_n39_));
  INV        m029(.A(i_8_), .Y(mai_mai_n40_));
  NOi21      m030(.An(i_4_), .B(i_0_), .Y(mai_mai_n41_));
  NA2        m031(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_2_), .B(i_8_), .Y(mai_mai_n43_));
  NOi31      m033(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n44_));
  NA2        m034(.A(mai_mai_n44_), .B(i_0_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_4_), .B(i_3_), .Y(mai_mai_n46_));
  NOi21      m036(.An(i_1_), .B(i_4_), .Y(mai_mai_n47_));
  OAI210     m037(.A0(mai_mai_n47_), .A1(mai_mai_n46_), .B0(mai_mai_n43_), .Y(mai_mai_n48_));
  NA2        m038(.A(mai_mai_n48_), .B(mai_mai_n45_), .Y(mai_mai_n49_));
  AN2        m039(.A(i_8_), .B(i_7_), .Y(mai_mai_n50_));
  NA2        m040(.A(mai_mai_n50_), .B(mai_mai_n12_), .Y(mai_mai_n51_));
  NOi21      m041(.An(i_8_), .B(i_7_), .Y(mai_mai_n52_));
  NA3        m042(.A(mai_mai_n52_), .B(mai_mai_n46_), .C(i_6_), .Y(mai_mai_n53_));
  OAI210     m043(.A0(mai_mai_n51_), .A1(mai_mai_n42_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  AOI220     m044(.A0(mai_mai_n54_), .A1(mai_mai_n26_), .B0(mai_mai_n49_), .B1(mai_mai_n30_), .Y(mai_mai_n55_));
  NA3        m045(.A(mai_mai_n55_), .B(mai_mai_n39_), .C(mai_mai_n25_), .Y(mai_mai_n56_));
  NA2        m046(.A(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NO3        m047(.A(mai_mai_n57_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n58_));
  NA2        m048(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n59_));
  AOI220     m049(.A0(mai_mai_n38_), .A1(i_1_), .B0(mai_mai_n34_), .B1(i_2_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_1_), .B(i_2_), .Y(mai_mai_n61_));
  NO2        m051(.A(mai_mai_n60_), .B(mai_mai_n59_), .Y(mai_mai_n62_));
  OAI210     m052(.A0(mai_mai_n62_), .A1(mai_mai_n58_), .B0(mai_mai_n14_), .Y(mai_mai_n63_));
  NOi32      m053(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n64_));
  NA2        m054(.A(mai_mai_n64_), .B(i_3_), .Y(mai_mai_n65_));
  NA3        m055(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n66_));
  NA2        m056(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NO2        m057(.A(i_0_), .B(i_4_), .Y(mai_mai_n68_));
  NA2        m058(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  NA2        m059(.A(mai_mai_n69_), .B(mai_mai_n63_), .Y(mai_mai_n70_));
  NAi21      m060(.An(i_3_), .B(i_6_), .Y(mai_mai_n71_));
  NO3        m061(.A(mai_mai_n71_), .B(i_0_), .C(mai_mai_n40_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n28_), .B(mai_mai_n27_), .Y(mai_mai_n73_));
  NOi21      m063(.An(i_7_), .B(i_8_), .Y(mai_mai_n74_));
  NA2        m064(.A(mai_mai_n74_), .B(mai_mai_n12_), .Y(mai_mai_n75_));
  OAI210     m065(.A0(mai_mai_n75_), .A1(mai_mai_n11_), .B0(mai_mai_n73_), .Y(mai_mai_n76_));
  OAI210     m066(.A0(mai_mai_n76_), .A1(mai_mai_n72_), .B0(mai_mai_n61_), .Y(mai_mai_n77_));
  AOI220     m067(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n18_), .B1(mai_mai_n26_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n79_));
  NO2        m069(.A(mai_mai_n79_), .B(mai_mai_n78_), .Y(mai_mai_n80_));
  INV        m070(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NA3        m071(.A(mai_mai_n52_), .B(mai_mai_n26_), .C(i_3_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n37_), .B(i_6_), .Y(mai_mai_n83_));
  AOI210     m073(.A0(mai_mai_n83_), .A1(mai_mai_n22_), .B0(mai_mai_n82_), .Y(mai_mai_n84_));
  NAi21      m074(.An(i_6_), .B(i_0_), .Y(mai_mai_n85_));
  NA3        m075(.A(mai_mai_n47_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n86_));
  NOi21      m076(.An(i_4_), .B(i_6_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_5_), .B(i_3_), .Y(mai_mai_n88_));
  NA3        m078(.A(mai_mai_n88_), .B(mai_mai_n61_), .C(mai_mai_n87_), .Y(mai_mai_n89_));
  OAI210     m079(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n61_), .B(mai_mai_n28_), .Y(mai_mai_n91_));
  NOi21      m081(.An(mai_mai_n35_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  NO3        m082(.A(mai_mai_n92_), .B(mai_mai_n90_), .C(mai_mai_n84_), .Y(mai_mai_n93_));
  NOi21      m083(.An(i_6_), .B(i_1_), .Y(mai_mai_n94_));
  AOI220     m084(.A0(mai_mai_n94_), .A1(i_7_), .B0(mai_mai_n24_), .B1(i_5_), .Y(mai_mai_n95_));
  NOi31      m085(.An(mai_mai_n41_), .B(mai_mai_n95_), .C(i_2_), .Y(mai_mai_n96_));
  AOI220     m086(.A0(mai_mai_n74_), .A1(mai_mai_n14_), .B0(mai_mai_n87_), .B1(mai_mai_n23_), .Y(mai_mai_n97_));
  NOi31      m087(.An(mai_mai_n38_), .B(mai_mai_n97_), .C(mai_mai_n26_), .Y(mai_mai_n98_));
  NO2        m088(.A(mai_mai_n98_), .B(mai_mai_n96_), .Y(mai_mai_n99_));
  NA4        m089(.A(mai_mai_n99_), .B(mai_mai_n93_), .C(mai_mai_n81_), .D(mai_mai_n77_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n43_), .B(mai_mai_n15_), .Y(mai_mai_n101_));
  NOi31      m091(.An(i_6_), .B(i_1_), .C(i_8_), .Y(mai_mai_n102_));
  NOi31      m092(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n103_));
  OAI210     m093(.A0(mai_mai_n103_), .A1(mai_mai_n102_), .B0(i_7_), .Y(mai_mai_n104_));
  NA3        m094(.A(mai_mai_n28_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n105_));
  NA4        m095(.A(mai_mai_n105_), .B(mai_mai_n104_), .C(mai_mai_n101_), .D(mai_mai_n91_), .Y(mai_mai_n106_));
  NA2        m096(.A(mai_mai_n106_), .B(mai_mai_n33_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n52_), .B(mai_mai_n44_), .C(i_6_), .Y(mai_mai_n108_));
  INV        m098(.A(mai_mai_n108_), .Y(mai_mai_n109_));
  NA3        m099(.A(mai_mai_n41_), .B(mai_mai_n35_), .C(mai_mai_n18_), .Y(mai_mai_n110_));
  NOi32      m100(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(mai_mai_n111_));
  NA2        m101(.A(mai_mai_n111_), .B(mai_mai_n102_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n112_), .B(mai_mai_n110_), .Y(mai_mai_n113_));
  NA4        m103(.A(mai_mai_n44_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n114_));
  NA4        m104(.A(mai_mai_n47_), .B(mai_mai_n30_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n115_));
  NA2        m105(.A(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NO3        m106(.A(mai_mai_n116_), .B(mai_mai_n113_), .C(mai_mai_n109_), .Y(mai_mai_n117_));
  NO2        m107(.A(mai_mai_n101_), .B(mai_mai_n83_), .Y(mai_mai_n118_));
  INV        m108(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  NA4        m109(.A(mai_mai_n88_), .B(mai_mai_n50_), .C(mai_mai_n37_), .D(mai_mai_n21_), .Y(mai_mai_n120_));
  NOi31      m110(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n121_));
  OAI210     m111(.A0(mai_mai_n111_), .A1(mai_mai_n64_), .B0(mai_mai_n121_), .Y(mai_mai_n122_));
  NA2        m112(.A(mai_mai_n122_), .B(mai_mai_n120_), .Y(mai_mai_n123_));
  INV        m113(.A(mai_mai_n123_), .Y(mai_mai_n124_));
  NA4        m114(.A(mai_mai_n124_), .B(mai_mai_n119_), .C(mai_mai_n117_), .D(mai_mai_n107_), .Y(mai_mai_n125_));
  OR4        m115(.A(mai_mai_n125_), .B(mai_mai_n100_), .C(mai_mai_n70_), .D(mai_mai_n56_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  INV        u002(.A(i_5_), .Y(men_men_n13_));
  NOi21      u003(.An(i_3_), .B(i_7_), .Y(men_men_n14_));
  INV        u004(.A(i_0_), .Y(men_men_n15_));
  NOi21      u005(.An(i_1_), .B(i_3_), .Y(men_men_n16_));
  INV        u006(.A(i_4_), .Y(men_men_n17_));
  NA2        u007(.A(i_0_), .B(men_men_n17_), .Y(men_men_n18_));
  INV        u008(.A(i_7_), .Y(men_men_n19_));
  NA3        u009(.A(i_6_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n20_));
  NOi21      u010(.An(i_8_), .B(i_6_), .Y(men_men_n21_));
  NOi21      u011(.An(i_1_), .B(i_8_), .Y(men_men_n22_));
  AOI220     u012(.A0(men_men_n22_), .A1(i_2_), .B0(men_men_n21_), .B1(i_5_), .Y(men_men_n23_));
  AOI210     u013(.A0(men_men_n23_), .A1(men_men_n20_), .B0(men_men_n18_), .Y(men_men_n24_));
  NA2        u014(.A(men_men_n24_), .B(men_men_n11_), .Y(men_men_n25_));
  NA2        u015(.A(i_0_), .B(men_men_n13_), .Y(men_men_n26_));
  NA2        u016(.A(men_men_n15_), .B(i_5_), .Y(men_men_n27_));
  NO2        u017(.A(i_2_), .B(i_4_), .Y(men_men_n28_));
  NA3        u018(.A(men_men_n28_), .B(i_6_), .C(i_8_), .Y(men_men_n29_));
  AOI210     u019(.A0(men_men_n27_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n30_));
  INV        u020(.A(i_2_), .Y(men_men_n31_));
  NOi21      u021(.An(i_5_), .B(i_0_), .Y(men_men_n32_));
  NOi21      u022(.An(i_6_), .B(i_8_), .Y(men_men_n33_));
  NOi21      u023(.An(i_7_), .B(i_1_), .Y(men_men_n34_));
  NOi21      u024(.An(i_0_), .B(i_4_), .Y(men_men_n35_));
  INV        u025(.A(i_1_), .Y(men_men_n36_));
  NOi21      u026(.An(i_3_), .B(i_0_), .Y(men_men_n37_));
  NA2        u027(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NA3        u028(.A(i_6_), .B(men_men_n13_), .C(i_7_), .Y(men_men_n39_));
  AOI210     u029(.A0(men_men_n39_), .A1(men_men_n20_), .B0(men_men_n38_), .Y(men_men_n40_));
  NO2        u030(.A(men_men_n40_), .B(men_men_n30_), .Y(men_men_n41_));
  INV        u031(.A(i_8_), .Y(men_men_n42_));
  NA2        u032(.A(i_1_), .B(men_men_n11_), .Y(men_men_n43_));
  NO4        u033(.A(men_men_n43_), .B(men_men_n26_), .C(i_2_), .D(men_men_n42_), .Y(men_men_n44_));
  NOi21      u034(.An(i_4_), .B(i_0_), .Y(men_men_n45_));
  AOI210     u035(.A0(men_men_n45_), .A1(men_men_n21_), .B0(men_men_n14_), .Y(men_men_n46_));
  NA2        u036(.A(i_1_), .B(men_men_n13_), .Y(men_men_n47_));
  NOi21      u037(.An(i_2_), .B(i_8_), .Y(men_men_n48_));
  NO3        u038(.A(men_men_n48_), .B(men_men_n45_), .C(men_men_n35_), .Y(men_men_n49_));
  NO3        u039(.A(men_men_n49_), .B(men_men_n47_), .C(men_men_n46_), .Y(men_men_n50_));
  NO2        u040(.A(men_men_n50_), .B(men_men_n44_), .Y(men_men_n51_));
  NOi31      u041(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n52_));
  NOi21      u042(.An(i_4_), .B(i_3_), .Y(men_men_n53_));
  NOi21      u043(.An(i_1_), .B(i_4_), .Y(men_men_n54_));
  AN2        u044(.A(i_8_), .B(i_7_), .Y(men_men_n55_));
  NOi21      u045(.An(i_8_), .B(i_7_), .Y(men_men_n56_));
  NA3        u046(.A(men_men_n51_), .B(men_men_n41_), .C(men_men_n25_), .Y(men_men_n57_));
  NA2        u047(.A(i_8_), .B(i_7_), .Y(men_men_n58_));
  NOi21      u048(.An(i_1_), .B(i_2_), .Y(men_men_n59_));
  NA3        u049(.A(men_men_n59_), .B(men_men_n45_), .C(i_6_), .Y(men_men_n60_));
  INV        u050(.A(men_men_n60_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(men_men_n13_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n56_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n63_));
  NA3        u053(.A(men_men_n22_), .B(i_0_), .C(men_men_n13_), .Y(men_men_n64_));
  NA2        u054(.A(men_men_n64_), .B(men_men_n63_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(men_men_n53_), .Y(men_men_n66_));
  NA2        u056(.A(men_men_n66_), .B(men_men_n62_), .Y(men_men_n67_));
  NAi21      u057(.An(i_3_), .B(i_6_), .Y(men_men_n68_));
  NOi21      u058(.An(i_7_), .B(i_8_), .Y(men_men_n69_));
  NOi31      u059(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n70_));
  AOI210     u060(.A0(men_men_n69_), .A1(men_men_n12_), .B0(men_men_n70_), .Y(men_men_n71_));
  NO2        u061(.A(men_men_n71_), .B(men_men_n11_), .Y(men_men_n72_));
  NA2        u062(.A(men_men_n72_), .B(men_men_n59_), .Y(men_men_n73_));
  NA3        u063(.A(men_men_n21_), .B(i_2_), .C(men_men_n13_), .Y(men_men_n74_));
  AOI210     u064(.A0(men_men_n18_), .A1(men_men_n43_), .B0(men_men_n74_), .Y(men_men_n75_));
  OAI210     u065(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n76_));
  NA3        u066(.A(men_men_n58_), .B(men_men_n16_), .C(men_men_n15_), .Y(men_men_n77_));
  NO2        u067(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NO2        u068(.A(men_men_n78_), .B(men_men_n75_), .Y(men_men_n79_));
  NA3        u069(.A(men_men_n56_), .B(men_men_n31_), .C(i_3_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n36_), .B(i_6_), .Y(men_men_n81_));
  AOI210     u071(.A0(men_men_n81_), .A1(men_men_n18_), .B0(men_men_n80_), .Y(men_men_n82_));
  NOi21      u072(.An(i_2_), .B(i_1_), .Y(men_men_n83_));
  AN3        u073(.A(men_men_n69_), .B(men_men_n83_), .C(men_men_n45_), .Y(men_men_n84_));
  NAi21      u074(.An(i_6_), .B(i_0_), .Y(men_men_n85_));
  NOi21      u075(.An(i_4_), .B(i_6_), .Y(men_men_n86_));
  NO2        u076(.A(men_men_n84_), .B(men_men_n82_), .Y(men_men_n87_));
  NA2        u077(.A(men_men_n56_), .B(men_men_n12_), .Y(men_men_n88_));
  NA2        u078(.A(men_men_n33_), .B(men_men_n13_), .Y(men_men_n89_));
  NOi21      u079(.An(i_3_), .B(i_1_), .Y(men_men_n90_));
  NA2        u080(.A(men_men_n90_), .B(i_4_), .Y(men_men_n91_));
  AOI210     u081(.A0(men_men_n89_), .A1(men_men_n88_), .B0(men_men_n91_), .Y(men_men_n92_));
  INV        u082(.A(men_men_n92_), .Y(men_men_n93_));
  NA4        u083(.A(men_men_n93_), .B(men_men_n87_), .C(men_men_n79_), .D(men_men_n73_), .Y(men_men_n94_));
  NA2        u084(.A(men_men_n53_), .B(men_men_n34_), .Y(men_men_n95_));
  AOI210     u085(.A0(men_men_n95_), .A1(men_men_n63_), .B0(men_men_n27_), .Y(men_men_n96_));
  NA4        u086(.A(men_men_n55_), .B(men_men_n83_), .C(men_men_n15_), .D(men_men_n12_), .Y(men_men_n97_));
  NAi31      u087(.An(men_men_n85_), .B(men_men_n69_), .C(men_men_n83_), .Y(men_men_n98_));
  NA3        u088(.A(men_men_n56_), .B(men_men_n52_), .C(i_6_), .Y(men_men_n99_));
  NA3        u089(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n100_));
  NOi21      u090(.An(i_0_), .B(i_2_), .Y(men_men_n101_));
  NA3        u091(.A(men_men_n101_), .B(men_men_n34_), .C(men_men_n86_), .Y(men_men_n102_));
  NA3        u092(.A(men_men_n101_), .B(men_men_n53_), .C(men_men_n33_), .Y(men_men_n103_));
  NA2        u093(.A(men_men_n103_), .B(men_men_n102_), .Y(men_men_n104_));
  NA4        u094(.A(men_men_n52_), .B(i_6_), .C(men_men_n13_), .D(i_7_), .Y(men_men_n105_));
  NA4        u095(.A(men_men_n54_), .B(men_men_n37_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n106_));
  NA2        u096(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NO4        u097(.A(men_men_n107_), .B(men_men_n104_), .C(men_men_n100_), .D(men_men_n96_), .Y(men_men_n108_));
  NOi21      u098(.An(i_5_), .B(i_2_), .Y(men_men_n109_));
  AOI220     u099(.A0(men_men_n109_), .A1(men_men_n69_), .B0(men_men_n55_), .B1(men_men_n28_), .Y(men_men_n110_));
  NO2        u100(.A(men_men_n110_), .B(men_men_n81_), .Y(men_men_n111_));
  NO4        u101(.A(i_2_), .B(men_men_n17_), .C(men_men_n11_), .D(men_men_n13_), .Y(men_men_n112_));
  NA2        u102(.A(i_2_), .B(i_4_), .Y(men_men_n113_));
  AOI210     u103(.A0(men_men_n85_), .A1(men_men_n68_), .B0(men_men_n113_), .Y(men_men_n114_));
  NO2        u104(.A(i_8_), .B(i_7_), .Y(men_men_n115_));
  OA210      u105(.A0(men_men_n114_), .A1(men_men_n112_), .B0(men_men_n115_), .Y(men_men_n116_));
  NA4        u106(.A(men_men_n90_), .B(i_0_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n117_));
  NO2        u107(.A(men_men_n117_), .B(i_4_), .Y(men_men_n118_));
  NO3        u108(.A(men_men_n118_), .B(men_men_n116_), .C(men_men_n111_), .Y(men_men_n119_));
  NA2        u109(.A(men_men_n69_), .B(men_men_n12_), .Y(men_men_n120_));
  NA3        u110(.A(i_2_), .B(i_1_), .C(men_men_n13_), .Y(men_men_n121_));
  NA2        u111(.A(men_men_n45_), .B(i_3_), .Y(men_men_n122_));
  AOI210     u112(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n120_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n101_), .B(men_men_n56_), .C(men_men_n86_), .Y(men_men_n124_));
  OAI210     u114(.A0(men_men_n80_), .A1(men_men_n27_), .B0(men_men_n124_), .Y(men_men_n125_));
  NA3        u115(.A(men_men_n70_), .B(men_men_n90_), .C(i_0_), .Y(men_men_n126_));
  NA3        u116(.A(men_men_n48_), .B(men_men_n32_), .C(men_men_n14_), .Y(men_men_n127_));
  NA2        u117(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO3        u118(.A(men_men_n128_), .B(men_men_n125_), .C(men_men_n123_), .Y(men_men_n129_));
  NA3        u119(.A(men_men_n129_), .B(men_men_n119_), .C(men_men_n108_), .Y(men_men_n130_));
  OR4        u120(.A(men_men_n130_), .B(men_men_n94_), .C(men_men_n67_), .D(men_men_n57_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule