library verilog;
use verilog.vl_types.all;
entity tb_somatorio is
end tb_somatorio;
