library verilog;
use verilog.vl_types.all;
entity decodificador2x4_vlg_sample_tst is
    port(
        e0              : in     vl_logic;
        e1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end decodificador2x4_vlg_sample_tst;
