library verilog;
use verilog.vl_types.all;
entity ex3_7 is
    port(
        A               : in     vl_logic_vector(3 downto 0);
        S               : out    vl_logic_vector(3 downto 0)
    );
end ex3_7;
