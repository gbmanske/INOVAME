//Benchmark atmr_alu4_1266_0.0625

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n137_, ori_ori_n138_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n640_, ori_ori_n641_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NO2        o034(.A(i_1_), .B(i_6_), .Y(ori_ori_n57_));
  NA2        o035(.A(i_8_), .B(i_7_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n57_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n60_));
  NAi21      o038(.An(i_2_), .B(i_7_), .Y(ori_ori_n61_));
  INV        o039(.A(i_1_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NA3        o041(.A(ori_ori_n63_), .B(ori_ori_n61_), .C(ori_ori_n31_), .Y(ori_ori_n64_));
  NA2        o042(.A(i_1_), .B(i_10_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(i_6_), .Y(ori_ori_n66_));
  NAi31      o044(.An(ori_ori_n66_), .B(ori_ori_n64_), .C(ori_ori_n60_), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n69_));
  NA2        o047(.A(i_1_), .B(i_6_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n70_), .B(ori_ori_n25_), .Y(ori_ori_n71_));
  INV        o049(.A(i_0_), .Y(ori_ori_n72_));
  NAi21      o050(.An(i_5_), .B(i_10_), .Y(ori_ori_n73_));
  NA2        o051(.A(i_5_), .B(i_9_), .Y(ori_ori_n74_));
  AOI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n73_), .B0(ori_ori_n72_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n71_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n69_), .A1(ori_ori_n68_), .B0(ori_ori_n76_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n77_), .A1(ori_ori_n67_), .B0(i_0_), .Y(ori_ori_n78_));
  NA2        o056(.A(i_12_), .B(i_5_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_2_), .B(i_8_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(ori_ori_n57_), .Y(ori_ori_n81_));
  NO2        o059(.A(i_3_), .B(i_9_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_7_), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n82_), .B(ori_ori_n62_), .Y(ori_ori_n84_));
  INV        o062(.A(i_6_), .Y(ori_ori_n85_));
  NO2        o063(.A(i_2_), .B(i_7_), .Y(ori_ori_n86_));
  INV        o064(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  OAI210     o065(.A0(ori_ori_n84_), .A1(ori_ori_n81_), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  NAi21      o066(.An(i_6_), .B(i_10_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_6_), .B(i_9_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n62_), .Y(ori_ori_n91_));
  NA2        o069(.A(i_2_), .B(i_6_), .Y(ori_ori_n92_));
  NO3        o070(.A(ori_ori_n92_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(ori_ori_n91_), .Y(ori_ori_n94_));
  AOI210     o072(.A0(ori_ori_n94_), .A1(ori_ori_n88_), .B0(ori_ori_n79_), .Y(ori_ori_n95_));
  AN3        o073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n96_));
  NAi21      o074(.An(i_6_), .B(i_11_), .Y(ori_ori_n97_));
  NO2        o075(.A(i_5_), .B(i_8_), .Y(ori_ori_n98_));
  NOi21      o076(.An(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  AOI220     o077(.A0(ori_ori_n99_), .A1(ori_ori_n61_), .B0(ori_ori_n96_), .B1(ori_ori_n32_), .Y(ori_ori_n100_));
  INV        o078(.A(i_7_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n46_), .B(ori_ori_n101_), .Y(ori_ori_n102_));
  NO2        o080(.A(i_0_), .B(i_5_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n103_), .B(ori_ori_n85_), .Y(ori_ori_n104_));
  NA2        o082(.A(i_12_), .B(i_3_), .Y(ori_ori_n105_));
  INV        o083(.A(ori_ori_n105_), .Y(ori_ori_n106_));
  NA3        o084(.A(ori_ori_n106_), .B(ori_ori_n104_), .C(ori_ori_n102_), .Y(ori_ori_n107_));
  NAi21      o085(.An(i_7_), .B(i_11_), .Y(ori_ori_n108_));
  AN2        o086(.A(i_2_), .B(i_10_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n109_), .B(i_7_), .Y(ori_ori_n110_));
  OR2        o088(.A(ori_ori_n79_), .B(ori_ori_n57_), .Y(ori_ori_n111_));
  NO2        o089(.A(i_8_), .B(ori_ori_n101_), .Y(ori_ori_n112_));
  NO3        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .C(ori_ori_n110_), .Y(ori_ori_n113_));
  NA2        o091(.A(i_12_), .B(i_7_), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n62_), .B(ori_ori_n26_), .Y(ori_ori_n115_));
  NA2        o093(.A(i_11_), .B(i_12_), .Y(ori_ori_n116_));
  INV        o094(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n117_), .B(ori_ori_n113_), .Y(ori_ori_n118_));
  NA3        o096(.A(ori_ori_n118_), .B(ori_ori_n107_), .C(ori_ori_n100_), .Y(ori_ori_n119_));
  NOi21      o097(.An(i_1_), .B(i_5_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(i_11_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n101_), .B(ori_ori_n37_), .Y(ori_ori_n122_));
  NA2        o100(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(ori_ori_n122_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n124_), .B(ori_ori_n46_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n90_), .B(ori_ori_n89_), .Y(ori_ori_n126_));
  NAi21      o104(.An(i_3_), .B(i_8_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(ori_ori_n61_), .Y(ori_ori_n128_));
  NOi31      o106(.An(ori_ori_n128_), .B(ori_ori_n126_), .C(ori_ori_n125_), .Y(ori_ori_n129_));
  NO2        o107(.A(i_1_), .B(ori_ori_n85_), .Y(ori_ori_n130_));
  NO2        o108(.A(i_6_), .B(i_5_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n131_), .B(i_3_), .Y(ori_ori_n132_));
  AO210      o110(.A0(ori_ori_n132_), .A1(ori_ori_n47_), .B0(ori_ori_n130_), .Y(ori_ori_n133_));
  OAI220     o111(.A0(ori_ori_n133_), .A1(ori_ori_n108_), .B0(ori_ori_n129_), .B1(ori_ori_n121_), .Y(ori_ori_n134_));
  NO3        o112(.A(ori_ori_n134_), .B(ori_ori_n119_), .C(ori_ori_n95_), .Y(ori_ori_n135_));
  NA3        o113(.A(ori_ori_n135_), .B(ori_ori_n78_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o114(.A(ori_ori_n62_), .B(ori_ori_n37_), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n641_), .B(ori_ori_n137_), .Y(ori_ori_n138_));
  NA4        o116(.A(ori_ori_n138_), .B(ori_ori_n76_), .C(ori_ori_n68_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o117(.A(i_8_), .B(i_7_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n140_), .B(i_6_), .Y(ori_ori_n141_));
  NO2        o119(.A(i_12_), .B(i_13_), .Y(ori_ori_n142_));
  NAi21      o120(.An(i_5_), .B(i_11_), .Y(ori_ori_n143_));
  NO2        o121(.A(i_0_), .B(i_1_), .Y(ori_ori_n144_));
  NA2        o122(.A(i_2_), .B(i_3_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n145_), .B(i_4_), .Y(ori_ori_n146_));
  AN2        o124(.A(ori_ori_n142_), .B(ori_ori_n82_), .Y(ori_ori_n147_));
  NA2        o125(.A(i_1_), .B(i_5_), .Y(ori_ori_n148_));
  OR2        o126(.A(i_0_), .B(i_1_), .Y(ori_ori_n149_));
  NO3        o127(.A(ori_ori_n149_), .B(ori_ori_n79_), .C(i_13_), .Y(ori_ori_n150_));
  NAi32      o128(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n151_));
  NAi21      o129(.An(ori_ori_n151_), .B(ori_ori_n150_), .Y(ori_ori_n152_));
  NOi21      o130(.An(i_4_), .B(i_10_), .Y(ori_ori_n153_));
  NOi21      o131(.An(i_4_), .B(i_9_), .Y(ori_ori_n154_));
  NOi21      o132(.An(i_11_), .B(i_13_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n72_), .B(ori_ori_n62_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n158_));
  NO2        o136(.A(i_2_), .B(i_1_), .Y(ori_ori_n159_));
  NAi21      o137(.An(i_4_), .B(i_12_), .Y(ori_ori_n160_));
  INV        o138(.A(i_8_), .Y(ori_ori_n161_));
  NO2        o139(.A(i_3_), .B(i_8_), .Y(ori_ori_n162_));
  NO3        o140(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n103_), .B(ori_ori_n57_), .Y(ori_ori_n164_));
  NO2        o142(.A(i_13_), .B(i_9_), .Y(ori_ori_n165_));
  NAi21      o143(.An(i_12_), .B(i_3_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n167_));
  NAi21      o145(.An(i_12_), .B(i_7_), .Y(ori_ori_n168_));
  NA3        o146(.A(i_13_), .B(ori_ori_n161_), .C(i_10_), .Y(ori_ori_n169_));
  NA2        o147(.A(i_0_), .B(i_5_), .Y(ori_ori_n170_));
  NAi31      o148(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n72_), .B(ori_ori_n26_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n46_), .B(ori_ori_n62_), .Y(ori_ori_n174_));
  INV        o152(.A(i_13_), .Y(ori_ori_n175_));
  NO2        o153(.A(i_12_), .B(ori_ori_n175_), .Y(ori_ori_n176_));
  NO2        o154(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n177_));
  OR2        o155(.A(i_8_), .B(i_7_), .Y(ori_ori_n178_));
  INV        o156(.A(i_12_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n44_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NO3        o158(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n181_));
  NA2        o159(.A(i_2_), .B(i_1_), .Y(ori_ori_n182_));
  NO3        o160(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n183_));
  NAi21      o161(.An(i_4_), .B(i_3_), .Y(ori_ori_n184_));
  NO2        o162(.A(i_0_), .B(i_6_), .Y(ori_ori_n185_));
  NOi41      o163(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n186_));
  NO2        o164(.A(i_11_), .B(ori_ori_n175_), .Y(ori_ori_n187_));
  NOi21      o165(.An(i_1_), .B(i_6_), .Y(ori_ori_n188_));
  NAi21      o166(.An(i_3_), .B(i_7_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n179_), .B(i_9_), .Y(ori_ori_n190_));
  OR4        o168(.A(ori_ori_n190_), .B(ori_ori_n189_), .C(ori_ori_n188_), .D(ori_ori_n158_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n192_));
  NA2        o170(.A(i_3_), .B(i_9_), .Y(ori_ori_n193_));
  NAi21      o171(.An(i_7_), .B(i_10_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n194_), .B(ori_ori_n193_), .Y(ori_ori_n195_));
  NA3        o173(.A(ori_ori_n195_), .B(ori_ori_n192_), .C(ori_ori_n63_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n196_), .B(ori_ori_n191_), .Y(ori_ori_n197_));
  INV        o175(.A(ori_ori_n141_), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n179_), .B(i_13_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(ori_ori_n74_), .Y(ori_ori_n200_));
  AOI220     o178(.A0(ori_ori_n200_), .A1(ori_ori_n198_), .B0(ori_ori_n197_), .B1(ori_ori_n187_), .Y(ori_ori_n201_));
  NA2        o179(.A(i_12_), .B(i_6_), .Y(ori_ori_n202_));
  OR2        o180(.A(i_13_), .B(i_9_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n184_), .B(i_2_), .Y(ori_ori_n204_));
  NA2        o182(.A(ori_ori_n187_), .B(i_9_), .Y(ori_ori_n205_));
  NO3        o183(.A(i_11_), .B(ori_ori_n175_), .C(ori_ori_n25_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n189_), .B(i_8_), .Y(ori_ori_n207_));
  NO3        o185(.A(i_12_), .B(ori_ori_n175_), .C(ori_ori_n37_), .Y(ori_ori_n208_));
  NO2        o186(.A(i_2_), .B(ori_ori_n101_), .Y(ori_ori_n209_));
  AN2        o187(.A(i_3_), .B(i_10_), .Y(ori_ori_n210_));
  NO2        o188(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n212_));
  NO3        o190(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n213_));
  NO2        o191(.A(i_2_), .B(i_3_), .Y(ori_ori_n214_));
  OR2        o192(.A(i_0_), .B(i_5_), .Y(ori_ori_n215_));
  NO2        o193(.A(i_12_), .B(i_10_), .Y(ori_ori_n216_));
  NOi21      o194(.An(i_5_), .B(i_0_), .Y(ori_ori_n217_));
  NO2        o195(.A(i_1_), .B(i_7_), .Y(ori_ori_n218_));
  NOi21      o196(.An(ori_ori_n148_), .B(ori_ori_n104_), .Y(ori_ori_n219_));
  NOi32      o197(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n220_));
  INV        o198(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n151_), .B(ori_ori_n149_), .Y(ori_ori_n222_));
  NOi32      o200(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n223_));
  NAi21      o201(.An(i_6_), .B(i_1_), .Y(ori_ori_n224_));
  NO2        o202(.A(i_1_), .B(ori_ori_n101_), .Y(ori_ori_n225_));
  NAi21      o203(.An(i_3_), .B(i_4_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(i_9_), .Y(ori_ori_n227_));
  AN2        o205(.A(i_6_), .B(i_7_), .Y(ori_ori_n228_));
  OAI210     o206(.A0(ori_ori_n228_), .A1(ori_ori_n225_), .B0(ori_ori_n227_), .Y(ori_ori_n229_));
  NA2        o207(.A(i_2_), .B(i_7_), .Y(ori_ori_n230_));
  NO2        o208(.A(ori_ori_n226_), .B(i_10_), .Y(ori_ori_n231_));
  NA3        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .C(ori_ori_n185_), .Y(ori_ori_n232_));
  AOI210     o210(.A0(ori_ori_n232_), .A1(ori_ori_n229_), .B0(ori_ori_n158_), .Y(ori_ori_n233_));
  AOI210     o211(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n234_), .A1(ori_ori_n159_), .B0(ori_ori_n231_), .Y(ori_ori_n235_));
  AOI220     o213(.A0(ori_ori_n231_), .A1(ori_ori_n218_), .B0(ori_ori_n181_), .B1(ori_ori_n159_), .Y(ori_ori_n236_));
  AOI210     o214(.A0(ori_ori_n236_), .A1(ori_ori_n235_), .B0(i_5_), .Y(ori_ori_n237_));
  NO3        o215(.A(ori_ori_n237_), .B(ori_ori_n233_), .C(ori_ori_n222_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n238_), .B(ori_ori_n221_), .Y(ori_ori_n239_));
  AN2        o217(.A(i_12_), .B(i_5_), .Y(ori_ori_n240_));
  NO2        o218(.A(i_11_), .B(i_6_), .Y(ori_ori_n241_));
  NO2        o219(.A(i_5_), .B(i_10_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n243_));
  NO3        o221(.A(ori_ori_n85_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n244_));
  NO2        o222(.A(i_11_), .B(i_12_), .Y(ori_ori_n245_));
  NAi21      o223(.An(i_13_), .B(i_0_), .Y(ori_ori_n246_));
  NO3        o224(.A(i_1_), .B(i_12_), .C(ori_ori_n85_), .Y(ori_ori_n247_));
  NO2        o225(.A(i_0_), .B(i_11_), .Y(ori_ori_n248_));
  AN2        o226(.A(i_1_), .B(i_6_), .Y(ori_ori_n249_));
  NOi21      o227(.An(i_2_), .B(i_12_), .Y(ori_ori_n250_));
  NAi21      o228(.An(i_9_), .B(i_4_), .Y(ori_ori_n251_));
  OR2        o229(.A(i_13_), .B(i_10_), .Y(ori_ori_n252_));
  NO3        o230(.A(ori_ori_n252_), .B(ori_ori_n116_), .C(ori_ori_n251_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n101_), .B(ori_ori_n25_), .Y(ori_ori_n254_));
  NA2        o232(.A(ori_ori_n208_), .B(ori_ori_n254_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n255_), .B(ori_ori_n219_), .Y(ori_ori_n256_));
  INV        o234(.A(ori_ori_n256_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n257_), .B(ori_ori_n26_), .Y(ori_ori_n258_));
  NA2        o236(.A(ori_ori_n161_), .B(i_10_), .Y(ori_ori_n259_));
  NA3        o237(.A(ori_ori_n192_), .B(ori_ori_n63_), .C(i_2_), .Y(ori_ori_n260_));
  NO2        o238(.A(ori_ori_n260_), .B(ori_ori_n259_), .Y(ori_ori_n261_));
  INV        o239(.A(ori_ori_n261_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n205_), .Y(ori_ori_n263_));
  NO3        o241(.A(ori_ori_n263_), .B(ori_ori_n258_), .C(ori_ori_n239_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n72_), .B(i_13_), .Y(ori_ori_n265_));
  NO2        o243(.A(i_10_), .B(i_9_), .Y(ori_ori_n266_));
  NAi21      o244(.An(i_12_), .B(i_8_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n267_), .B(i_3_), .Y(ori_ori_n268_));
  NO3        o246(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n269_));
  NA2        o247(.A(ori_ori_n202_), .B(ori_ori_n97_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(ori_ori_n269_), .Y(ori_ori_n271_));
  NA2        o249(.A(i_8_), .B(i_9_), .Y(ori_ori_n272_));
  AOI210     o250(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n273_));
  OR2        o251(.A(ori_ori_n273_), .B(ori_ori_n272_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n208_), .B(ori_ori_n164_), .Y(ori_ori_n275_));
  NO2        o253(.A(ori_ori_n275_), .B(ori_ori_n274_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n187_), .B(ori_ori_n211_), .Y(ori_ori_n277_));
  NO3        o255(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n278_));
  INV        o256(.A(ori_ori_n278_), .Y(ori_ori_n279_));
  NA3        o257(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n280_));
  NA4        o258(.A(ori_ori_n143_), .B(ori_ori_n115_), .C(ori_ori_n79_), .D(ori_ori_n23_), .Y(ori_ori_n281_));
  OAI220     o259(.A0(ori_ori_n281_), .A1(ori_ori_n280_), .B0(ori_ori_n279_), .B1(ori_ori_n277_), .Y(ori_ori_n282_));
  NO2        o260(.A(ori_ori_n282_), .B(ori_ori_n276_), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n96_), .B(i_13_), .Y(ori_ori_n284_));
  NO2        o262(.A(i_11_), .B(i_1_), .Y(ori_ori_n285_));
  NOi21      o263(.An(i_2_), .B(i_7_), .Y(ori_ori_n286_));
  NO2        o264(.A(i_6_), .B(i_10_), .Y(ori_ori_n287_));
  NA3        o265(.A(ori_ori_n186_), .B(ori_ori_n155_), .C(ori_ori_n131_), .Y(ori_ori_n288_));
  NA2        o266(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n289_));
  NO2        o267(.A(ori_ori_n149_), .B(i_3_), .Y(ori_ori_n290_));
  NAi31      o268(.An(ori_ori_n289_), .B(ori_ori_n290_), .C(ori_ori_n176_), .Y(ori_ori_n291_));
  NA3        o269(.A(ori_ori_n243_), .B(ori_ori_n157_), .C(ori_ori_n146_), .Y(ori_ori_n292_));
  NA3        o270(.A(ori_ori_n292_), .B(ori_ori_n291_), .C(ori_ori_n288_), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n293_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n278_), .B(ori_ori_n242_), .Y(ori_ori_n295_));
  NAi21      o273(.An(ori_ori_n169_), .B(ori_ori_n245_), .Y(ori_ori_n296_));
  NA2        o274(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n213_), .B(ori_ori_n181_), .Y(ori_ori_n298_));
  OAI220     o276(.A0(ori_ori_n298_), .A1(ori_ori_n260_), .B0(ori_ori_n297_), .B1(ori_ori_n284_), .Y(ori_ori_n299_));
  INV        o277(.A(ori_ori_n299_), .Y(ori_ori_n300_));
  NA3        o278(.A(ori_ori_n300_), .B(ori_ori_n294_), .C(ori_ori_n283_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n240_), .B(ori_ori_n175_), .Y(ori_ori_n302_));
  NA2        o280(.A(ori_ori_n228_), .B(ori_ori_n223_), .Y(ori_ori_n303_));
  OR2        o281(.A(ori_ori_n302_), .B(ori_ori_n303_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n305_));
  AOI210     o283(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n253_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n306_), .B(ori_ori_n304_), .Y(ori_ori_n307_));
  NO2        o285(.A(i_12_), .B(ori_ori_n161_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n309_), .B(i_6_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n149_), .B(i_5_), .Y(ori_ori_n311_));
  NA3        o289(.A(ori_ori_n170_), .B(ori_ori_n70_), .C(ori_ori_n44_), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n208_), .B(ori_ori_n83_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n312_), .B(ori_ori_n313_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n174_), .B(ori_ori_n173_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n266_), .B(ori_ori_n172_), .Y(ori_ori_n316_));
  NO2        o294(.A(ori_ori_n315_), .B(ori_ori_n316_), .Y(ori_ori_n317_));
  AOI210     o295(.A0(ori_ori_n224_), .A1(ori_ori_n46_), .B0(ori_ori_n225_), .Y(ori_ori_n318_));
  NA2        o296(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n319_));
  NA3        o297(.A(ori_ori_n308_), .B(ori_ori_n206_), .C(ori_ori_n319_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n318_), .B(ori_ori_n320_), .Y(ori_ori_n321_));
  NO3        o299(.A(ori_ori_n321_), .B(ori_ori_n317_), .C(ori_ori_n314_), .Y(ori_ori_n322_));
  NO3        o300(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n252_), .B(i_1_), .Y(ori_ori_n324_));
  NOi31      o302(.An(ori_ori_n324_), .B(ori_ori_n270_), .C(ori_ori_n72_), .Y(ori_ori_n325_));
  NOi21      o303(.An(i_10_), .B(i_6_), .Y(ori_ori_n326_));
  NO2        o304(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n114_), .B(ori_ori_n23_), .Y(ori_ori_n328_));
  NO2        o306(.A(i_12_), .B(ori_ori_n85_), .Y(ori_ori_n329_));
  OR2        o307(.A(i_2_), .B(i_5_), .Y(ori_ori_n330_));
  OR2        o308(.A(ori_ori_n330_), .B(ori_ori_n249_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n230_), .B(ori_ori_n185_), .Y(ori_ori_n332_));
  AOI210     o310(.A0(ori_ori_n332_), .A1(ori_ori_n331_), .B0(ori_ori_n296_), .Y(ori_ori_n333_));
  INV        o311(.A(ori_ori_n333_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n334_), .B(ori_ori_n322_), .Y(ori_ori_n335_));
  NO3        o313(.A(ori_ori_n335_), .B(ori_ori_n307_), .C(ori_ori_n301_), .Y(ori_ori_n336_));
  NA3        o314(.A(ori_ori_n336_), .B(ori_ori_n264_), .C(ori_ori_n201_), .Y(ori7));
  NO2        o315(.A(ori_ori_n92_), .B(ori_ori_n54_), .Y(ori_ori_n338_));
  NA2        o316(.A(ori_ori_n287_), .B(ori_ori_n83_), .Y(ori_ori_n339_));
  NA2        o317(.A(i_11_), .B(ori_ori_n161_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n142_), .B(ori_ori_n340_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n339_), .Y(ori_ori_n342_));
  NA3        o320(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n343_));
  NO2        o321(.A(ori_ori_n179_), .B(i_4_), .Y(ori_ori_n344_));
  NA2        o322(.A(ori_ori_n344_), .B(i_8_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n105_), .B(ori_ori_n343_), .Y(ori_ori_n346_));
  NA2        o324(.A(i_2_), .B(ori_ori_n85_), .Y(ori_ori_n347_));
  OAI210     o325(.A0(ori_ori_n86_), .A1(ori_ori_n162_), .B0(ori_ori_n163_), .Y(ori_ori_n348_));
  NO2        o326(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n349_));
  NA2        o327(.A(i_4_), .B(i_8_), .Y(ori_ori_n350_));
  AOI210     o328(.A0(ori_ori_n350_), .A1(ori_ori_n210_), .B0(ori_ori_n349_), .Y(ori_ori_n351_));
  OAI220     o329(.A0(ori_ori_n351_), .A1(ori_ori_n347_), .B0(ori_ori_n348_), .B1(i_13_), .Y(ori_ori_n352_));
  NO4        o330(.A(ori_ori_n352_), .B(ori_ori_n346_), .C(ori_ori_n342_), .D(ori_ori_n338_), .Y(ori_ori_n353_));
  AOI210     o331(.A0(ori_ori_n127_), .A1(ori_ori_n61_), .B0(i_10_), .Y(ori_ori_n354_));
  AOI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n179_), .B0(ori_ori_n153_), .Y(ori_ori_n355_));
  OR2        o333(.A(i_6_), .B(i_10_), .Y(ori_ori_n356_));
  OR3        o334(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n357_));
  OR2        o335(.A(ori_ori_n355_), .B(ori_ori_n203_), .Y(ori_ori_n358_));
  AOI210     o336(.A0(ori_ori_n358_), .A1(ori_ori_n353_), .B0(ori_ori_n62_), .Y(ori_ori_n359_));
  NOi21      o337(.An(i_11_), .B(i_7_), .Y(ori_ori_n360_));
  AO210      o338(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n361_), .B(ori_ori_n360_), .Y(ori_ori_n362_));
  NA2        o340(.A(ori_ori_n362_), .B(ori_ori_n165_), .Y(ori_ori_n363_));
  NA3        o341(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n363_), .B(ori_ori_n62_), .Y(ori_ori_n365_));
  OR2        o343(.A(ori_ori_n236_), .B(ori_ori_n41_), .Y(ori_ori_n366_));
  NO3        o344(.A(ori_ori_n194_), .B(ori_ori_n166_), .C(ori_ori_n340_), .Y(ori_ori_n367_));
  OAI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n176_), .B0(ori_ori_n62_), .Y(ori_ori_n368_));
  OR2        o346(.A(ori_ori_n166_), .B(ori_ori_n108_), .Y(ori_ori_n369_));
  NO2        o347(.A(i_1_), .B(i_12_), .Y(ori_ori_n370_));
  NA3        o348(.A(ori_ori_n370_), .B(ori_ori_n109_), .C(ori_ori_n24_), .Y(ori_ori_n371_));
  BUFFER     o349(.A(ori_ori_n371_), .Y(ori_ori_n372_));
  NA3        o350(.A(ori_ori_n372_), .B(ori_ori_n368_), .C(ori_ori_n366_), .Y(ori_ori_n373_));
  OAI210     o351(.A0(ori_ori_n373_), .A1(ori_ori_n365_), .B0(i_6_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n364_), .B(ori_ori_n108_), .Y(ori_ori_n375_));
  NA2        o353(.A(ori_ori_n375_), .B(ori_ori_n329_), .Y(ori_ori_n376_));
  NO2        o354(.A(i_6_), .B(i_11_), .Y(ori_ori_n377_));
  NA2        o355(.A(ori_ori_n376_), .B(ori_ori_n271_), .Y(ori_ori_n378_));
  NO3        o356(.A(ori_ori_n356_), .B(ori_ori_n178_), .C(ori_ori_n23_), .Y(ori_ori_n379_));
  AOI210     o357(.A0(i_1_), .A1(ori_ori_n195_), .B0(ori_ori_n379_), .Y(ori_ori_n380_));
  NO2        o358(.A(ori_ori_n380_), .B(ori_ori_n44_), .Y(ori_ori_n381_));
  INV        o359(.A(i_2_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n137_), .B(i_9_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n383_), .B(ori_ori_n382_), .Y(ori_ori_n385_));
  AOI210     o363(.A0(ori_ori_n285_), .A1(ori_ori_n254_), .B0(ori_ori_n183_), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n386_), .B(ori_ori_n347_), .Y(ori_ori_n387_));
  NO2        o365(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n388_));
  OR2        o366(.A(ori_ori_n387_), .B(ori_ori_n385_), .Y(ori_ori_n389_));
  NO3        o367(.A(ori_ori_n389_), .B(ori_ori_n381_), .C(ori_ori_n378_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n179_), .B(ori_ori_n101_), .Y(ori_ori_n391_));
  NO2        o369(.A(ori_ori_n391_), .B(ori_ori_n360_), .Y(ori_ori_n392_));
  NA2        o370(.A(ori_ori_n392_), .B(i_1_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n393_), .B(ori_ori_n357_), .Y(ori_ori_n394_));
  NO2        o372(.A(ori_ori_n251_), .B(ori_ori_n85_), .Y(ori_ori_n395_));
  NA2        o373(.A(ori_ori_n394_), .B(ori_ori_n46_), .Y(ori_ori_n396_));
  NA2        o374(.A(i_3_), .B(ori_ori_n161_), .Y(ori_ori_n397_));
  NO2        o375(.A(ori_ori_n397_), .B(ori_ori_n114_), .Y(ori_ori_n398_));
  AN2        o376(.A(ori_ori_n398_), .B(ori_ori_n310_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n178_), .B(ori_ori_n44_), .Y(ori_ori_n400_));
  NO3        o378(.A(ori_ori_n400_), .B(ori_ori_n212_), .C(ori_ori_n180_), .Y(ori_ori_n401_));
  NO2        o379(.A(ori_ori_n116_), .B(ori_ori_n37_), .Y(ori_ori_n402_));
  NO2        o380(.A(ori_ori_n402_), .B(i_6_), .Y(ori_ori_n403_));
  NO2        o381(.A(ori_ori_n85_), .B(i_9_), .Y(ori_ori_n404_));
  NO2        o382(.A(ori_ori_n404_), .B(ori_ori_n62_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n405_), .B(ori_ori_n370_), .Y(ori_ori_n406_));
  NO4        o384(.A(ori_ori_n406_), .B(ori_ori_n403_), .C(ori_ori_n401_), .D(i_4_), .Y(ori_ori_n407_));
  NA2        o385(.A(i_1_), .B(i_3_), .Y(ori_ori_n408_));
  NO2        o386(.A(ori_ori_n272_), .B(ori_ori_n92_), .Y(ori_ori_n409_));
  AOI210     o387(.A0(ori_ori_n400_), .A1(ori_ori_n326_), .B0(ori_ori_n409_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n410_), .B(ori_ori_n408_), .Y(ori_ori_n411_));
  NO3        o389(.A(ori_ori_n411_), .B(ori_ori_n407_), .C(ori_ori_n399_), .Y(ori_ori_n412_));
  NA4        o390(.A(ori_ori_n412_), .B(ori_ori_n396_), .C(ori_ori_n390_), .D(ori_ori_n374_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n228_), .B(ori_ori_n227_), .Y(ori_ori_n414_));
  INV        o392(.A(ori_ori_n414_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(i_1_), .Y(ori_ori_n416_));
  AOI210     o394(.A0(ori_ori_n202_), .A1(ori_ori_n97_), .B0(i_1_), .Y(ori_ori_n417_));
  NO2        o395(.A(ori_ori_n226_), .B(i_2_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n418_), .B(ori_ori_n417_), .Y(ori_ori_n419_));
  AOI210     o397(.A0(ori_ori_n419_), .A1(ori_ori_n416_), .B0(i_13_), .Y(ori_ori_n420_));
  OR2        o398(.A(i_11_), .B(i_7_), .Y(ori_ori_n421_));
  NO2        o399(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n422_));
  NO2        o400(.A(ori_ori_n286_), .B(ori_ori_n24_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n423_), .B(ori_ori_n395_), .Y(ori_ori_n424_));
  OAI220     o402(.A0(ori_ori_n424_), .A1(ori_ori_n41_), .B0(ori_ori_n640_), .B1(ori_ori_n92_), .Y(ori_ori_n425_));
  INV        o403(.A(ori_ori_n425_), .Y(ori_ori_n426_));
  NA2        o404(.A(ori_ori_n241_), .B(ori_ori_n384_), .Y(ori_ori_n427_));
  NO2        o405(.A(ori_ori_n427_), .B(ori_ori_n184_), .Y(ori_ori_n428_));
  AOI210     o406(.A0(ori_ori_n267_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n429_));
  NOi31      o407(.An(ori_ori_n429_), .B(ori_ori_n339_), .C(ori_ori_n44_), .Y(ori_ori_n430_));
  NA2        o408(.A(ori_ori_n126_), .B(i_13_), .Y(ori_ori_n431_));
  NO2        o409(.A(ori_ori_n431_), .B(ori_ori_n417_), .Y(ori_ori_n432_));
  NA2        o410(.A(ori_ori_n26_), .B(ori_ori_n161_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n433_), .B(i_7_), .Y(ori_ori_n434_));
  AOI220     o412(.A0(ori_ori_n241_), .A1(ori_ori_n384_), .B0(ori_ori_n91_), .B1(ori_ori_n102_), .Y(ori_ori_n435_));
  NO2        o413(.A(ori_ori_n435_), .B(ori_ori_n345_), .Y(ori_ori_n436_));
  NO4        o414(.A(ori_ori_n436_), .B(ori_ori_n432_), .C(ori_ori_n430_), .D(ori_ori_n428_), .Y(ori_ori_n437_));
  OR2        o415(.A(i_11_), .B(i_6_), .Y(ori_ori_n438_));
  NA3        o416(.A(ori_ori_n344_), .B(ori_ori_n433_), .C(i_7_), .Y(ori_ori_n439_));
  NO2        o417(.A(ori_ori_n439_), .B(ori_ori_n438_), .Y(ori_ori_n440_));
  NA3        o418(.A(ori_ori_n250_), .B(ori_ori_n349_), .C(ori_ori_n97_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n377_), .B(i_13_), .Y(ori_ori_n442_));
  NAi21      o420(.An(i_11_), .B(i_12_), .Y(ori_ori_n443_));
  NOi41      o421(.An(ori_ori_n110_), .B(ori_ori_n443_), .C(i_13_), .D(ori_ori_n85_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n444_), .B(ori_ori_n46_), .Y(ori_ori_n445_));
  NA3        o423(.A(ori_ori_n445_), .B(ori_ori_n442_), .C(ori_ori_n441_), .Y(ori_ori_n446_));
  OAI210     o424(.A0(ori_ori_n446_), .A1(ori_ori_n440_), .B0(ori_ori_n62_), .Y(ori_ori_n447_));
  NO2        o425(.A(i_2_), .B(i_12_), .Y(ori_ori_n448_));
  NA2        o426(.A(ori_ori_n225_), .B(ori_ori_n448_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n227_), .B(ori_ori_n225_), .Y(ori_ori_n450_));
  NA2        o428(.A(ori_ori_n450_), .B(ori_ori_n449_), .Y(ori_ori_n451_));
  NA3        o429(.A(ori_ori_n451_), .B(ori_ori_n45_), .C(ori_ori_n175_), .Y(ori_ori_n452_));
  NA4        o430(.A(ori_ori_n452_), .B(ori_ori_n447_), .C(ori_ori_n437_), .D(ori_ori_n426_), .Y(ori_ori_n453_));
  OR4        o431(.A(ori_ori_n453_), .B(ori_ori_n420_), .C(ori_ori_n413_), .D(ori_ori_n359_), .Y(ori5));
  NA2        o432(.A(ori_ori_n392_), .B(ori_ori_n204_), .Y(ori_ori_n455_));
  AN2        o433(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n456_));
  NA3        o434(.A(ori_ori_n456_), .B(ori_ori_n448_), .C(ori_ori_n108_), .Y(ori_ori_n457_));
  NO2        o435(.A(ori_ori_n345_), .B(i_11_), .Y(ori_ori_n458_));
  NA2        o436(.A(ori_ori_n86_), .B(ori_ori_n458_), .Y(ori_ori_n459_));
  NA3        o437(.A(ori_ori_n459_), .B(ori_ori_n457_), .C(ori_ori_n455_), .Y(ori_ori_n460_));
  NO3        o438(.A(i_11_), .B(ori_ori_n179_), .C(i_13_), .Y(ori_ori_n461_));
  NO2        o439(.A(ori_ori_n123_), .B(ori_ori_n23_), .Y(ori_ori_n462_));
  NA2        o440(.A(i_12_), .B(i_8_), .Y(ori_ori_n463_));
  OAI210     o441(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n463_), .Y(ori_ori_n464_));
  INV        o442(.A(ori_ori_n266_), .Y(ori_ori_n465_));
  AOI220     o443(.A0(ori_ori_n214_), .A1(ori_ori_n328_), .B0(ori_ori_n464_), .B1(ori_ori_n462_), .Y(ori_ori_n466_));
  INV        o444(.A(ori_ori_n466_), .Y(ori_ori_n467_));
  NO2        o445(.A(ori_ori_n467_), .B(ori_ori_n460_), .Y(ori_ori_n468_));
  INV        o446(.A(ori_ori_n155_), .Y(ori_ori_n469_));
  INV        o447(.A(ori_ori_n186_), .Y(ori_ori_n470_));
  OAI210     o448(.A0(ori_ori_n418_), .A1(ori_ori_n268_), .B0(ori_ori_n110_), .Y(ori_ori_n471_));
  AOI210     o449(.A0(ori_ori_n471_), .A1(ori_ori_n470_), .B0(ori_ori_n469_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n272_), .B(ori_ori_n26_), .Y(ori_ori_n473_));
  NO2        o451(.A(ori_ori_n473_), .B(ori_ori_n254_), .Y(ori_ori_n474_));
  NA2        o452(.A(ori_ori_n474_), .B(i_2_), .Y(ori_ori_n475_));
  INV        o453(.A(ori_ori_n475_), .Y(ori_ori_n476_));
  AOI210     o454(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n252_), .Y(ori_ori_n477_));
  AOI210     o455(.A0(ori_ori_n477_), .A1(ori_ori_n476_), .B0(ori_ori_n472_), .Y(ori_ori_n478_));
  NO2        o456(.A(ori_ori_n160_), .B(ori_ori_n124_), .Y(ori_ori_n479_));
  OAI210     o457(.A0(ori_ori_n479_), .A1(ori_ori_n462_), .B0(i_2_), .Y(ori_ori_n480_));
  INV        o458(.A(ori_ori_n156_), .Y(ori_ori_n481_));
  NO3        o459(.A(ori_ori_n361_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n482_));
  AOI210     o460(.A0(ori_ori_n481_), .A1(ori_ori_n86_), .B0(ori_ori_n482_), .Y(ori_ori_n483_));
  AOI210     o461(.A0(ori_ori_n483_), .A1(ori_ori_n480_), .B0(ori_ori_n161_), .Y(ori_ori_n484_));
  OA210      o462(.A0(ori_ori_n362_), .A1(ori_ori_n125_), .B0(i_13_), .Y(ori_ori_n485_));
  NA2        o463(.A(ori_ori_n147_), .B(ori_ori_n340_), .Y(ori_ori_n486_));
  NO2        o464(.A(ori_ori_n486_), .B(ori_ori_n230_), .Y(ori_ori_n487_));
  AOI210     o465(.A0(ori_ori_n166_), .A1(ori_ori_n145_), .B0(ori_ori_n305_), .Y(ori_ori_n488_));
  OAI210     o466(.A0(ori_ori_n488_), .A1(ori_ori_n176_), .B0(ori_ori_n254_), .Y(ori_ori_n489_));
  NO2        o467(.A(ori_ori_n102_), .B(ori_ori_n44_), .Y(ori_ori_n490_));
  INV        o468(.A(ori_ori_n209_), .Y(ori_ori_n491_));
  NA4        o469(.A(ori_ori_n491_), .B(ori_ori_n210_), .C(ori_ori_n123_), .D(ori_ori_n42_), .Y(ori_ori_n492_));
  OAI210     o470(.A0(ori_ori_n492_), .A1(ori_ori_n490_), .B0(ori_ori_n489_), .Y(ori_ori_n493_));
  NO4        o471(.A(ori_ori_n493_), .B(ori_ori_n487_), .C(ori_ori_n485_), .D(ori_ori_n484_), .Y(ori_ori_n494_));
  NA2        o472(.A(ori_ori_n328_), .B(ori_ori_n28_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n461_), .B(ori_ori_n207_), .Y(ori_ori_n496_));
  NA2        o474(.A(ori_ori_n496_), .B(ori_ori_n495_), .Y(ori_ori_n497_));
  NO2        o475(.A(ori_ori_n61_), .B(i_12_), .Y(ori_ori_n498_));
  NO2        o476(.A(ori_ori_n498_), .B(ori_ori_n125_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n499_), .B(ori_ori_n340_), .Y(ori_ori_n500_));
  AOI220     o478(.A0(ori_ori_n500_), .A1(ori_ori_n36_), .B0(ori_ori_n497_), .B1(ori_ori_n46_), .Y(ori_ori_n501_));
  NA4        o479(.A(ori_ori_n501_), .B(ori_ori_n494_), .C(ori_ori_n478_), .D(ori_ori_n468_), .Y(ori6));
  NO2        o480(.A(ori_ori_n171_), .B(ori_ori_n289_), .Y(ori_ori_n503_));
  INV        o481(.A(ori_ori_n217_), .Y(ori_ori_n504_));
  OR2        o482(.A(ori_ori_n504_), .B(i_12_), .Y(ori_ori_n505_));
  NA2        o483(.A(ori_ori_n329_), .B(ori_ori_n62_), .Y(ori_ori_n506_));
  INV        o484(.A(ori_ori_n506_), .Y(ori_ori_n507_));
  NA2        o485(.A(ori_ori_n507_), .B(ori_ori_n72_), .Y(ori_ori_n508_));
  INV        o486(.A(ori_ori_n216_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n74_), .B(ori_ori_n130_), .Y(ori_ori_n510_));
  INV        o488(.A(ori_ori_n123_), .Y(ori_ori_n511_));
  NA2        o489(.A(ori_ori_n511_), .B(ori_ori_n46_), .Y(ori_ori_n512_));
  AOI210     o490(.A0(ori_ori_n512_), .A1(ori_ori_n510_), .B0(ori_ori_n509_), .Y(ori_ori_n513_));
  NO2        o491(.A(ori_ori_n188_), .B(i_9_), .Y(ori_ori_n514_));
  NA2        o492(.A(ori_ori_n514_), .B(ori_ori_n498_), .Y(ori_ori_n515_));
  AOI210     o493(.A0(ori_ori_n515_), .A1(ori_ori_n303_), .B0(ori_ori_n158_), .Y(ori_ori_n516_));
  NAi32      o494(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n438_), .B(ori_ori_n517_), .Y(ori_ori_n518_));
  OR3        o496(.A(ori_ori_n518_), .B(ori_ori_n516_), .C(ori_ori_n513_), .Y(ori_ori_n519_));
  NO2        o497(.A(ori_ori_n421_), .B(i_2_), .Y(ori_ori_n520_));
  NA2        o498(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n521_));
  NO2        o499(.A(ori_ori_n521_), .B(ori_ori_n249_), .Y(ori_ori_n522_));
  NA2        o500(.A(ori_ori_n522_), .B(ori_ori_n520_), .Y(ori_ori_n523_));
  BUFFER     o501(.A(ori_ori_n362_), .Y(ori_ori_n524_));
  NA3        o502(.A(ori_ori_n524_), .B(ori_ori_n144_), .C(ori_ori_n68_), .Y(ori_ori_n525_));
  AO210      o503(.A0(ori_ori_n295_), .A1(ori_ori_n465_), .B0(ori_ori_n36_), .Y(ori_ori_n526_));
  NA3        o504(.A(ori_ori_n526_), .B(ori_ori_n525_), .C(ori_ori_n523_), .Y(ori_ori_n527_));
  NO2        o505(.A(i_6_), .B(i_11_), .Y(ori_ori_n528_));
  AOI220     o506(.A0(ori_ori_n528_), .A1(ori_ori_n323_), .B0(ori_ori_n503_), .B1(ori_ori_n434_), .Y(ori_ori_n529_));
  NA3        o507(.A(ori_ori_n230_), .B(ori_ori_n181_), .C(ori_ori_n144_), .Y(ori_ori_n530_));
  NA2        o508(.A(ori_ori_n244_), .B(ori_ori_n69_), .Y(ori_ori_n531_));
  NA4        o509(.A(ori_ori_n531_), .B(ori_ori_n530_), .C(ori_ori_n529_), .D(ori_ori_n348_), .Y(ori_ori_n532_));
  NA2        o510(.A(ori_ori_n268_), .B(ori_ori_n266_), .Y(ori_ori_n533_));
  NO2        o511(.A(ori_ori_n356_), .B(ori_ori_n102_), .Y(ori_ori_n534_));
  OAI210     o512(.A0(ori_ori_n534_), .A1(ori_ori_n111_), .B0(ori_ori_n248_), .Y(ori_ori_n535_));
  INV        o513(.A(ori_ori_n331_), .Y(ori_ori_n536_));
  NA3        o514(.A(ori_ori_n536_), .B(ori_ori_n216_), .C(i_7_), .Y(ori_ori_n537_));
  NA3        o515(.A(ori_ori_n537_), .B(ori_ori_n535_), .C(ori_ori_n533_), .Y(ori_ori_n538_));
  NO4        o516(.A(ori_ori_n538_), .B(ori_ori_n532_), .C(ori_ori_n527_), .D(ori_ori_n519_), .Y(ori_ori_n539_));
  NA4        o517(.A(ori_ori_n539_), .B(ori_ori_n508_), .C(ori_ori_n505_), .D(ori_ori_n238_), .Y(ori3));
  NA2        o518(.A(i_12_), .B(i_10_), .Y(ori_ori_n541_));
  NO2        o519(.A(i_11_), .B(ori_ori_n179_), .Y(ori_ori_n542_));
  NA3        o520(.A(ori_ori_n530_), .B(ori_ori_n348_), .C(ori_ori_n229_), .Y(ori_ori_n543_));
  NA2        o521(.A(ori_ori_n543_), .B(ori_ori_n40_), .Y(ori_ori_n544_));
  NOi21      o522(.An(ori_ori_n96_), .B(ori_ori_n474_), .Y(ori_ori_n545_));
  NO3        o523(.A(ori_ori_n369_), .B(ori_ori_n272_), .C(ori_ori_n130_), .Y(ori_ori_n546_));
  AN2        o524(.A(ori_ori_n270_), .B(ori_ori_n55_), .Y(ori_ori_n547_));
  NO3        o525(.A(ori_ori_n547_), .B(ori_ori_n546_), .C(ori_ori_n545_), .Y(ori_ori_n548_));
  AOI210     o526(.A0(ori_ori_n548_), .A1(ori_ori_n544_), .B0(ori_ori_n48_), .Y(ori_ori_n549_));
  NO4        o527(.A(ori_ori_n234_), .B(ori_ori_n240_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n550_));
  NA2        o528(.A(ori_ori_n158_), .B(ori_ori_n326_), .Y(ori_ori_n551_));
  NOi31      o529(.An(ori_ori_n551_), .B(ori_ori_n550_), .C(ori_ori_n39_), .Y(ori_ori_n552_));
  NO2        o530(.A(ori_ori_n552_), .B(ori_ori_n62_), .Y(ori_ori_n553_));
  NOi21      o531(.An(i_5_), .B(i_9_), .Y(ori_ori_n554_));
  NA2        o532(.A(ori_ori_n554_), .B(ori_ori_n265_), .Y(ori_ori_n555_));
  BUFFER     o533(.A(ori_ori_n202_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n556_), .B(ori_ori_n285_), .Y(ori_ori_n557_));
  NO2        o535(.A(ori_ori_n557_), .B(ori_ori_n555_), .Y(ori_ori_n558_));
  NO3        o536(.A(ori_ori_n558_), .B(ori_ori_n553_), .C(ori_ori_n549_), .Y(ori_ori_n559_));
  NA2        o537(.A(ori_ori_n327_), .B(i_0_), .Y(ori_ori_n560_));
  NO4        o538(.A(ori_ori_n330_), .B(ori_ori_n168_), .C(ori_ori_n252_), .D(ori_ori_n249_), .Y(ori_ori_n561_));
  NA2        o539(.A(ori_ori_n561_), .B(i_11_), .Y(ori_ori_n562_));
  NA2        o540(.A(ori_ori_n461_), .B(ori_ori_n217_), .Y(ori_ori_n563_));
  AOI210     o541(.A0(ori_ori_n287_), .A1(ori_ori_n86_), .B0(ori_ori_n57_), .Y(ori_ori_n564_));
  NO2        o542(.A(ori_ori_n564_), .B(ori_ori_n563_), .Y(ori_ori_n565_));
  NO2        o543(.A(ori_ori_n190_), .B(ori_ori_n148_), .Y(ori_ori_n566_));
  NA2        o544(.A(i_0_), .B(i_10_), .Y(ori_ori_n567_));
  INV        o545(.A(ori_ori_n309_), .Y(ori_ori_n568_));
  NO4        o546(.A(ori_ori_n114_), .B(ori_ori_n57_), .C(ori_ori_n397_), .D(i_5_), .Y(ori_ori_n569_));
  AO220      o547(.A0(ori_ori_n569_), .A1(ori_ori_n568_), .B0(ori_ori_n566_), .B1(i_6_), .Y(ori_ori_n570_));
  NO2        o548(.A(ori_ori_n570_), .B(ori_ori_n565_), .Y(ori_ori_n571_));
  NA2        o549(.A(ori_ori_n571_), .B(ori_ori_n562_), .Y(ori_ori_n572_));
  NO2        o550(.A(ori_ori_n103_), .B(ori_ori_n37_), .Y(ori_ori_n573_));
  NA2        o551(.A(i_11_), .B(i_9_), .Y(ori_ori_n574_));
  NO3        o552(.A(i_12_), .B(ori_ori_n574_), .C(ori_ori_n347_), .Y(ori_ori_n575_));
  AN2        o553(.A(ori_ori_n575_), .B(ori_ori_n573_), .Y(ori_ori_n576_));
  NA2        o554(.A(ori_ori_n243_), .B(ori_ori_n157_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n577_), .B(ori_ori_n152_), .Y(ori_ori_n578_));
  NO2        o556(.A(ori_ori_n574_), .B(ori_ori_n72_), .Y(ori_ori_n579_));
  INV        o557(.A(ori_ori_n247_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n580_), .B(ori_ori_n555_), .Y(ori_ori_n581_));
  NO3        o559(.A(ori_ori_n581_), .B(ori_ori_n578_), .C(ori_ori_n576_), .Y(ori_ori_n582_));
  NA2        o560(.A(ori_ori_n388_), .B(ori_ori_n120_), .Y(ori_ori_n583_));
  NO2        o561(.A(i_6_), .B(ori_ori_n583_), .Y(ori_ori_n584_));
  NA2        o562(.A(ori_ori_n155_), .B(ori_ori_n103_), .Y(ori_ori_n585_));
  INV        o563(.A(ori_ori_n584_), .Y(ori_ori_n586_));
  INV        o564(.A(ori_ori_n215_), .Y(ori_ori_n587_));
  NA2        o565(.A(ori_ori_n586_), .B(ori_ori_n582_), .Y(ori_ori_n588_));
  NO2        o566(.A(ori_ori_n541_), .B(ori_ori_n214_), .Y(ori_ori_n589_));
  NA2        o567(.A(ori_ori_n589_), .B(ori_ori_n579_), .Y(ori_ori_n590_));
  NA2        o568(.A(ori_ori_n423_), .B(ori_ori_n311_), .Y(ori_ori_n591_));
  NAi21      o569(.An(i_9_), .B(i_5_), .Y(ori_ori_n592_));
  NO2        o570(.A(ori_ori_n592_), .B(ori_ori_n246_), .Y(ori_ori_n593_));
  NA2        o571(.A(ori_ori_n593_), .B(ori_ori_n362_), .Y(ori_ori_n594_));
  OAI220     o572(.A0(ori_ori_n594_), .A1(ori_ori_n85_), .B0(ori_ori_n591_), .B1(ori_ori_n156_), .Y(ori_ori_n595_));
  NO2        o573(.A(ori_ori_n595_), .B(ori_ori_n307_), .Y(ori_ori_n596_));
  NA2        o574(.A(ori_ori_n596_), .B(ori_ori_n590_), .Y(ori_ori_n597_));
  NO3        o575(.A(ori_ori_n597_), .B(ori_ori_n588_), .C(ori_ori_n572_), .Y(ori_ori_n598_));
  AOI210     o576(.A0(ori_ori_n506_), .A1(ori_ori_n414_), .B0(ori_ori_n585_), .Y(ori_ori_n599_));
  INV        o577(.A(ori_ori_n599_), .Y(ori_ori_n600_));
  OAI210     o578(.A0(ori_ori_n185_), .A1(i_9_), .B0(ori_ori_n177_), .Y(ori_ori_n601_));
  AOI210     o579(.A0(ori_ori_n601_), .A1(ori_ori_n560_), .B0(ori_ori_n148_), .Y(ori_ori_n602_));
  INV        o580(.A(ori_ori_n602_), .Y(ori_ori_n603_));
  NA2        o581(.A(ori_ori_n603_), .B(ori_ori_n600_), .Y(ori_ori_n604_));
  NO3        o582(.A(ori_ori_n567_), .B(ori_ori_n554_), .C(ori_ori_n160_), .Y(ori_ori_n605_));
  AOI220     o583(.A0(ori_ori_n605_), .A1(i_11_), .B0(ori_ori_n325_), .B1(ori_ori_n74_), .Y(ori_ori_n606_));
  NO3        o584(.A(ori_ori_n167_), .B(ori_ori_n240_), .C(i_0_), .Y(ori_ori_n607_));
  OAI210     o585(.A0(ori_ori_n607_), .A1(ori_ori_n75_), .B0(i_13_), .Y(ori_ori_n608_));
  NA2        o586(.A(ori_ori_n608_), .B(ori_ori_n606_), .Y(ori_ori_n609_));
  NA3        o587(.A(ori_ori_n242_), .B(ori_ori_n155_), .C(ori_ori_n154_), .Y(ori_ori_n610_));
  INV        o588(.A(ori_ori_n610_), .Y(ori_ori_n611_));
  NO3        o589(.A(ori_ori_n574_), .B(ori_ori_n170_), .C(ori_ori_n160_), .Y(ori_ori_n612_));
  NO2        o590(.A(ori_ori_n612_), .B(ori_ori_n611_), .Y(ori_ori_n613_));
  NA2        o591(.A(ori_ori_n613_), .B(ori_ori_n288_), .Y(ori_ori_n614_));
  NO2        o592(.A(ori_ori_n85_), .B(i_5_), .Y(ori_ori_n615_));
  NA3        o593(.A(ori_ori_n542_), .B(ori_ori_n109_), .C(ori_ori_n123_), .Y(ori_ori_n616_));
  INV        o594(.A(ori_ori_n616_), .Y(ori_ori_n617_));
  NA2        o595(.A(ori_ori_n617_), .B(ori_ori_n615_), .Y(ori_ori_n618_));
  NAi21      o596(.An(ori_ori_n183_), .B(ori_ori_n184_), .Y(ori_ori_n619_));
  NO4        o597(.A(ori_ori_n182_), .B(ori_ori_n167_), .C(i_0_), .D(i_12_), .Y(ori_ori_n620_));
  NA2        o598(.A(ori_ori_n620_), .B(ori_ori_n619_), .Y(ori_ori_n621_));
  NA2        o599(.A(ori_ori_n621_), .B(ori_ori_n618_), .Y(ori_ori_n622_));
  NO4        o600(.A(ori_ori_n622_), .B(ori_ori_n614_), .C(ori_ori_n609_), .D(ori_ori_n604_), .Y(ori_ori_n623_));
  NA2        o601(.A(ori_ori_n520_), .B(ori_ori_n37_), .Y(ori_ori_n624_));
  NA2        o602(.A(ori_ori_n624_), .B(ori_ori_n355_), .Y(ori_ori_n625_));
  NA2        o603(.A(ori_ori_n625_), .B(ori_ori_n165_), .Y(ori_ori_n626_));
  NAi31      o604(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n627_));
  AOI210     o605(.A0(ori_ori_n116_), .A1(ori_ori_n69_), .B0(ori_ori_n627_), .Y(ori_ori_n628_));
  AOI210     o606(.A0(ori_ori_n628_), .A1(ori_ori_n48_), .B0(ori_ori_n561_), .Y(ori_ori_n629_));
  AOI210     o607(.A0(ori_ori_n629_), .A1(ori_ori_n626_), .B0(ori_ori_n72_), .Y(ori_ori_n630_));
  INV        o608(.A(ori_ori_n237_), .Y(ori_ori_n631_));
  NO2        o609(.A(ori_ori_n631_), .B(ori_ori_n469_), .Y(ori_ori_n632_));
  NO3        o610(.A(ori_ori_n58_), .B(ori_ori_n57_), .C(i_4_), .Y(ori_ori_n633_));
  OAI210     o611(.A0(ori_ori_n587_), .A1(ori_ori_n211_), .B0(ori_ori_n633_), .Y(ori_ori_n634_));
  NO2        o612(.A(ori_ori_n634_), .B(ori_ori_n443_), .Y(ori_ori_n635_));
  NO3        o613(.A(ori_ori_n635_), .B(ori_ori_n632_), .C(ori_ori_n630_), .Y(ori_ori_n636_));
  NA4        o614(.A(ori_ori_n636_), .B(ori_ori_n623_), .C(ori_ori_n598_), .D(ori_ori_n559_), .Y(ori4));
  INV        o615(.A(ori_ori_n422_), .Y(ori_ori_n640_));
  INV        o616(.A(i_6_), .Y(ori_ori_n641_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m0020(.A(mai_mai_n35_), .Y(mai1));
  INV        m0021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m0022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m0023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m0024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m0025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m0026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m0027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  OAI210     m0028(.A0(mai_mai_n50_), .A1(i_3_), .B0(mai_mai_n48_), .Y(mai_mai_n51_));
  AOI210     m0029(.A0(mai_mai_n51_), .A1(mai_mai_n47_), .B0(mai_mai_n46_), .Y(mai_mai_n52_));
  NA2        m0030(.A(i_0_), .B(i_2_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_7_), .B(i_9_), .Y(mai_mai_n54_));
  NA2        m0032(.A(mai_mai_n52_), .B(mai_mai_n45_), .Y(mai_mai_n55_));
  NA3        m0033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n56_));
  NO2        m0034(.A(i_1_), .B(i_6_), .Y(mai_mai_n57_));
  NA2        m0035(.A(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  OAI210     m0036(.A0(mai_mai_n58_), .A1(mai_mai_n57_), .B0(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m0037(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n60_));
  NAi21      m0038(.An(i_2_), .B(i_7_), .Y(mai_mai_n61_));
  INV        m0039(.A(i_1_), .Y(mai_mai_n62_));
  NA2        m0040(.A(mai_mai_n62_), .B(i_6_), .Y(mai_mai_n63_));
  NA3        m0041(.A(mai_mai_n63_), .B(mai_mai_n61_), .C(mai_mai_n31_), .Y(mai_mai_n64_));
  NA2        m0042(.A(i_1_), .B(i_10_), .Y(mai_mai_n65_));
  NO2        m0043(.A(mai_mai_n65_), .B(i_6_), .Y(mai_mai_n66_));
  NAi31      m0044(.An(mai_mai_n66_), .B(mai_mai_n64_), .C(mai_mai_n60_), .Y(mai_mai_n67_));
  NA2        m0045(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n68_));
  AOI210     m0046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n69_));
  NA2        m0047(.A(i_1_), .B(i_6_), .Y(mai_mai_n70_));
  NO2        m0048(.A(mai_mai_n70_), .B(mai_mai_n25_), .Y(mai_mai_n71_));
  INV        m0049(.A(i_0_), .Y(mai_mai_n72_));
  NAi21      m0050(.An(i_5_), .B(i_10_), .Y(mai_mai_n73_));
  NA2        m0051(.A(i_5_), .B(i_9_), .Y(mai_mai_n74_));
  AOI210     m0052(.A0(mai_mai_n74_), .A1(mai_mai_n73_), .B0(mai_mai_n72_), .Y(mai_mai_n75_));
  NO2        m0053(.A(mai_mai_n75_), .B(mai_mai_n71_), .Y(mai_mai_n76_));
  OAI210     m0054(.A0(mai_mai_n69_), .A1(mai_mai_n68_), .B0(mai_mai_n76_), .Y(mai_mai_n77_));
  OAI210     m0055(.A0(mai_mai_n77_), .A1(mai_mai_n67_), .B0(i_0_), .Y(mai_mai_n78_));
  NA2        m0056(.A(i_12_), .B(i_5_), .Y(mai_mai_n79_));
  NA2        m0057(.A(i_2_), .B(i_8_), .Y(mai_mai_n80_));
  NO2        m0058(.A(i_3_), .B(i_9_), .Y(mai_mai_n81_));
  NO2        m0059(.A(i_3_), .B(i_7_), .Y(mai_mai_n82_));
  INV        m0060(.A(i_6_), .Y(mai_mai_n83_));
  OR4        m0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n84_));
  INV        m0062(.A(mai_mai_n84_), .Y(mai_mai_n85_));
  NO2        m0063(.A(i_2_), .B(i_7_), .Y(mai_mai_n86_));
  NAi21      m0064(.An(i_6_), .B(i_10_), .Y(mai_mai_n87_));
  NA2        m0065(.A(i_6_), .B(i_9_), .Y(mai_mai_n88_));
  AOI210     m0066(.A0(mai_mai_n88_), .A1(mai_mai_n87_), .B0(mai_mai_n62_), .Y(mai_mai_n89_));
  NA2        m0067(.A(i_2_), .B(i_6_), .Y(mai_mai_n90_));
  INV        m0068(.A(mai_mai_n89_), .Y(mai_mai_n91_));
  NO2        m0069(.A(mai_mai_n91_), .B(mai_mai_n79_), .Y(mai_mai_n92_));
  AN3        m0070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n93_));
  NAi21      m0071(.An(i_6_), .B(i_11_), .Y(mai_mai_n94_));
  NO2        m0072(.A(i_5_), .B(i_8_), .Y(mai_mai_n95_));
  NOi21      m0073(.An(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  AOI220     m0074(.A0(mai_mai_n96_), .A1(mai_mai_n61_), .B0(mai_mai_n93_), .B1(mai_mai_n32_), .Y(mai_mai_n97_));
  INV        m0075(.A(i_7_), .Y(mai_mai_n98_));
  NA2        m0076(.A(mai_mai_n46_), .B(mai_mai_n98_), .Y(mai_mai_n99_));
  NO2        m0077(.A(i_0_), .B(i_5_), .Y(mai_mai_n100_));
  NO2        m0078(.A(mai_mai_n100_), .B(mai_mai_n83_), .Y(mai_mai_n101_));
  NA2        m0079(.A(i_12_), .B(i_3_), .Y(mai_mai_n102_));
  INV        m0080(.A(mai_mai_n102_), .Y(mai_mai_n103_));
  NA3        m0081(.A(mai_mai_n103_), .B(mai_mai_n101_), .C(mai_mai_n99_), .Y(mai_mai_n104_));
  NAi21      m0082(.An(i_7_), .B(i_11_), .Y(mai_mai_n105_));
  NO3        m0083(.A(mai_mai_n105_), .B(mai_mai_n87_), .C(mai_mai_n53_), .Y(mai_mai_n106_));
  AN2        m0084(.A(i_2_), .B(i_10_), .Y(mai_mai_n107_));
  NO2        m0085(.A(mai_mai_n107_), .B(i_7_), .Y(mai_mai_n108_));
  OR2        m0086(.A(mai_mai_n79_), .B(mai_mai_n57_), .Y(mai_mai_n109_));
  NO2        m0087(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n110_));
  NO3        m0088(.A(mai_mai_n110_), .B(mai_mai_n109_), .C(mai_mai_n108_), .Y(mai_mai_n111_));
  NA2        m0089(.A(i_12_), .B(i_7_), .Y(mai_mai_n112_));
  NO2        m0090(.A(mai_mai_n62_), .B(mai_mai_n26_), .Y(mai_mai_n113_));
  NA2        m0091(.A(mai_mai_n113_), .B(i_0_), .Y(mai_mai_n114_));
  NA2        m0092(.A(i_11_), .B(i_12_), .Y(mai_mai_n115_));
  OAI210     m0093(.A0(mai_mai_n114_), .A1(mai_mai_n112_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m0094(.A(mai_mai_n116_), .B(mai_mai_n111_), .Y(mai_mai_n117_));
  NAi41      m0095(.An(mai_mai_n106_), .B(mai_mai_n117_), .C(mai_mai_n104_), .D(mai_mai_n97_), .Y(mai_mai_n118_));
  NOi21      m0096(.An(i_1_), .B(i_5_), .Y(mai_mai_n119_));
  NA2        m0097(.A(mai_mai_n119_), .B(i_11_), .Y(mai_mai_n120_));
  NA2        m0098(.A(mai_mai_n98_), .B(mai_mai_n37_), .Y(mai_mai_n121_));
  NA2        m0099(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n122_));
  NA2        m0100(.A(mai_mai_n122_), .B(mai_mai_n121_), .Y(mai_mai_n123_));
  NO2        m0101(.A(mai_mai_n123_), .B(mai_mai_n46_), .Y(mai_mai_n124_));
  NA2        m0102(.A(mai_mai_n88_), .B(mai_mai_n87_), .Y(mai_mai_n125_));
  NAi21      m0103(.An(i_3_), .B(i_8_), .Y(mai_mai_n126_));
  NA2        m0104(.A(mai_mai_n126_), .B(mai_mai_n61_), .Y(mai_mai_n127_));
  NOi31      m0105(.An(mai_mai_n127_), .B(mai_mai_n125_), .C(mai_mai_n124_), .Y(mai_mai_n128_));
  NO2        m0106(.A(i_1_), .B(mai_mai_n83_), .Y(mai_mai_n129_));
  NO2        m0107(.A(i_6_), .B(i_5_), .Y(mai_mai_n130_));
  NA2        m0108(.A(mai_mai_n130_), .B(i_3_), .Y(mai_mai_n131_));
  AO210      m0109(.A0(mai_mai_n131_), .A1(mai_mai_n47_), .B0(mai_mai_n129_), .Y(mai_mai_n132_));
  OAI220     m0110(.A0(mai_mai_n132_), .A1(mai_mai_n105_), .B0(mai_mai_n128_), .B1(mai_mai_n120_), .Y(mai_mai_n133_));
  NO3        m0111(.A(mai_mai_n133_), .B(mai_mai_n118_), .C(mai_mai_n92_), .Y(mai_mai_n134_));
  NA3        m0112(.A(mai_mai_n134_), .B(mai_mai_n78_), .C(mai_mai_n55_), .Y(mai2));
  NO2        m0113(.A(mai_mai_n62_), .B(mai_mai_n37_), .Y(mai_mai_n136_));
  NA2        m0114(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n137_));
  NA2        m0115(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n138_));
  NA4        m0116(.A(mai_mai_n138_), .B(mai_mai_n76_), .C(mai_mai_n68_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0117(.A(i_8_), .B(i_7_), .Y(mai_mai_n140_));
  NA2        m0118(.A(mai_mai_n140_), .B(i_6_), .Y(mai_mai_n141_));
  NO2        m0119(.A(i_12_), .B(i_13_), .Y(mai_mai_n142_));
  NAi21      m0120(.An(i_5_), .B(i_11_), .Y(mai_mai_n143_));
  NOi21      m0121(.An(mai_mai_n142_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  NO2        m0122(.A(i_0_), .B(i_1_), .Y(mai_mai_n145_));
  NA2        m0123(.A(i_2_), .B(i_3_), .Y(mai_mai_n146_));
  NO2        m0124(.A(mai_mai_n146_), .B(i_4_), .Y(mai_mai_n147_));
  NA3        m0125(.A(mai_mai_n147_), .B(mai_mai_n145_), .C(mai_mai_n144_), .Y(mai_mai_n148_));
  AN2        m0126(.A(mai_mai_n142_), .B(mai_mai_n81_), .Y(mai_mai_n149_));
  NO2        m0127(.A(mai_mai_n149_), .B(mai_mai_n27_), .Y(mai_mai_n150_));
  NA2        m0128(.A(i_1_), .B(i_5_), .Y(mai_mai_n151_));
  NO2        m0129(.A(mai_mai_n72_), .B(mai_mai_n46_), .Y(mai_mai_n152_));
  NA2        m0130(.A(mai_mai_n152_), .B(mai_mai_n36_), .Y(mai_mai_n153_));
  NO3        m0131(.A(mai_mai_n153_), .B(mai_mai_n151_), .C(mai_mai_n150_), .Y(mai_mai_n154_));
  OR2        m0132(.A(i_0_), .B(i_1_), .Y(mai_mai_n155_));
  NO3        m0133(.A(mai_mai_n155_), .B(mai_mai_n79_), .C(i_13_), .Y(mai_mai_n156_));
  NAi32      m0134(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n157_));
  NAi21      m0135(.An(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  NOi21      m0136(.An(i_4_), .B(i_10_), .Y(mai_mai_n159_));
  NA2        m0137(.A(mai_mai_n159_), .B(mai_mai_n40_), .Y(mai_mai_n160_));
  NO2        m0138(.A(i_3_), .B(i_5_), .Y(mai_mai_n161_));
  NO3        m0139(.A(mai_mai_n72_), .B(i_2_), .C(i_1_), .Y(mai_mai_n162_));
  NA2        m0140(.A(mai_mai_n162_), .B(mai_mai_n161_), .Y(mai_mai_n163_));
  OAI210     m0141(.A0(mai_mai_n163_), .A1(mai_mai_n160_), .B0(mai_mai_n158_), .Y(mai_mai_n164_));
  NO2        m0142(.A(mai_mai_n164_), .B(mai_mai_n154_), .Y(mai_mai_n165_));
  AOI210     m0143(.A0(mai_mai_n165_), .A1(mai_mai_n148_), .B0(mai_mai_n141_), .Y(mai_mai_n166_));
  NA2        m0144(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n167_));
  NOi21      m0145(.An(i_4_), .B(i_9_), .Y(mai_mai_n168_));
  NOi21      m0146(.An(i_11_), .B(i_13_), .Y(mai_mai_n169_));
  NA2        m0147(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  OR2        m0148(.A(mai_mai_n170_), .B(mai_mai_n167_), .Y(mai_mai_n171_));
  NO2        m0149(.A(i_4_), .B(i_5_), .Y(mai_mai_n172_));
  NAi21      m0150(.An(i_12_), .B(i_11_), .Y(mai_mai_n173_));
  NO2        m0151(.A(mai_mai_n173_), .B(i_13_), .Y(mai_mai_n174_));
  NA3        m0152(.A(mai_mai_n174_), .B(mai_mai_n172_), .C(mai_mai_n81_), .Y(mai_mai_n175_));
  AOI210     m0153(.A0(mai_mai_n175_), .A1(mai_mai_n171_), .B0(mai_mai_n1046_), .Y(mai_mai_n176_));
  NO2        m0154(.A(mai_mai_n72_), .B(mai_mai_n62_), .Y(mai_mai_n177_));
  NA2        m0155(.A(mai_mai_n177_), .B(mai_mai_n46_), .Y(mai_mai_n178_));
  NA2        m0156(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n179_));
  NAi31      m0157(.An(mai_mai_n179_), .B(mai_mai_n149_), .C(i_11_), .Y(mai_mai_n180_));
  NA2        m0158(.A(i_3_), .B(i_5_), .Y(mai_mai_n181_));
  OR2        m0159(.A(mai_mai_n181_), .B(mai_mai_n170_), .Y(mai_mai_n182_));
  AOI210     m0160(.A0(mai_mai_n182_), .A1(mai_mai_n180_), .B0(mai_mai_n178_), .Y(mai_mai_n183_));
  NO2        m0161(.A(mai_mai_n72_), .B(i_5_), .Y(mai_mai_n184_));
  NO2        m0162(.A(i_13_), .B(i_10_), .Y(mai_mai_n185_));
  NA3        m0163(.A(mai_mai_n185_), .B(mai_mai_n184_), .C(mai_mai_n44_), .Y(mai_mai_n186_));
  NO2        m0164(.A(i_2_), .B(i_1_), .Y(mai_mai_n187_));
  NA2        m0165(.A(mai_mai_n187_), .B(i_3_), .Y(mai_mai_n188_));
  NAi21      m0166(.An(i_4_), .B(i_12_), .Y(mai_mai_n189_));
  NO4        m0167(.A(mai_mai_n189_), .B(mai_mai_n188_), .C(mai_mai_n186_), .D(mai_mai_n25_), .Y(mai_mai_n190_));
  NO3        m0168(.A(mai_mai_n190_), .B(mai_mai_n183_), .C(mai_mai_n176_), .Y(mai_mai_n191_));
  INV        m0169(.A(i_8_), .Y(mai_mai_n192_));
  NO2        m0170(.A(mai_mai_n192_), .B(i_7_), .Y(mai_mai_n193_));
  NA2        m0171(.A(mai_mai_n193_), .B(i_6_), .Y(mai_mai_n194_));
  NO3        m0172(.A(i_3_), .B(mai_mai_n83_), .C(mai_mai_n48_), .Y(mai_mai_n195_));
  NA2        m0173(.A(mai_mai_n195_), .B(mai_mai_n110_), .Y(mai_mai_n196_));
  NO3        m0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n197_));
  NA3        m0175(.A(mai_mai_n197_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n198_));
  NO3        m0176(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n199_));
  OAI210     m0177(.A0(mai_mai_n93_), .A1(i_12_), .B0(mai_mai_n199_), .Y(mai_mai_n200_));
  AOI210     m0178(.A0(mai_mai_n200_), .A1(mai_mai_n198_), .B0(mai_mai_n196_), .Y(mai_mai_n201_));
  NO2        m0179(.A(i_3_), .B(i_8_), .Y(mai_mai_n202_));
  NO3        m0180(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n203_));
  NA3        m0181(.A(mai_mai_n203_), .B(mai_mai_n202_), .C(mai_mai_n40_), .Y(mai_mai_n204_));
  NO2        m0182(.A(i_13_), .B(i_9_), .Y(mai_mai_n205_));
  NA3        m0183(.A(mai_mai_n205_), .B(i_6_), .C(mai_mai_n192_), .Y(mai_mai_n206_));
  NAi21      m0184(.An(i_12_), .B(i_3_), .Y(mai_mai_n207_));
  NO2        m0185(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n208_));
  NO3        m0186(.A(i_0_), .B(i_2_), .C(mai_mai_n62_), .Y(mai_mai_n209_));
  NA3        m0187(.A(mai_mai_n209_), .B(mai_mai_n208_), .C(i_10_), .Y(mai_mai_n210_));
  OAI220     m0188(.A0(mai_mai_n210_), .A1(mai_mai_n206_), .B0(mai_mai_n57_), .B1(mai_mai_n204_), .Y(mai_mai_n211_));
  AOI210     m0189(.A0(mai_mai_n211_), .A1(i_7_), .B0(mai_mai_n201_), .Y(mai_mai_n212_));
  OAI220     m0190(.A0(mai_mai_n212_), .A1(i_4_), .B0(mai_mai_n194_), .B1(mai_mai_n191_), .Y(mai_mai_n213_));
  NAi21      m0191(.An(i_12_), .B(i_7_), .Y(mai_mai_n214_));
  NA3        m0192(.A(i_13_), .B(mai_mai_n192_), .C(i_10_), .Y(mai_mai_n215_));
  NO2        m0193(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n216_));
  NA2        m0194(.A(i_0_), .B(i_5_), .Y(mai_mai_n217_));
  OAI220     m0195(.A0(mai_mai_n83_), .A1(mai_mai_n188_), .B0(mai_mai_n178_), .B1(mai_mai_n131_), .Y(mai_mai_n218_));
  NAi31      m0196(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n219_));
  NO2        m0197(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n220_));
  NO2        m0198(.A(mai_mai_n46_), .B(mai_mai_n62_), .Y(mai_mai_n221_));
  NA3        m0199(.A(mai_mai_n221_), .B(i_0_), .C(mai_mai_n220_), .Y(mai_mai_n222_));
  INV        m0200(.A(i_13_), .Y(mai_mai_n223_));
  NO2        m0201(.A(i_12_), .B(mai_mai_n223_), .Y(mai_mai_n224_));
  NA3        m0202(.A(mai_mai_n224_), .B(mai_mai_n197_), .C(mai_mai_n195_), .Y(mai_mai_n225_));
  OAI210     m0203(.A0(mai_mai_n222_), .A1(mai_mai_n219_), .B0(mai_mai_n225_), .Y(mai_mai_n226_));
  AOI220     m0204(.A0(mai_mai_n226_), .A1(mai_mai_n140_), .B0(mai_mai_n218_), .B1(mai_mai_n216_), .Y(mai_mai_n227_));
  NO2        m0205(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n228_));
  NO2        m0206(.A(mai_mai_n181_), .B(i_4_), .Y(mai_mai_n229_));
  NA2        m0207(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n230_));
  OR2        m0208(.A(i_8_), .B(i_7_), .Y(mai_mai_n231_));
  NO2        m0209(.A(mai_mai_n231_), .B(mai_mai_n83_), .Y(mai_mai_n232_));
  NO2        m0210(.A(mai_mai_n53_), .B(i_1_), .Y(mai_mai_n233_));
  NA2        m0211(.A(mai_mai_n233_), .B(mai_mai_n232_), .Y(mai_mai_n234_));
  INV        m0212(.A(i_12_), .Y(mai_mai_n235_));
  NO3        m0213(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n236_));
  NA2        m0214(.A(i_2_), .B(i_1_), .Y(mai_mai_n237_));
  NO2        m0215(.A(mai_mai_n234_), .B(mai_mai_n230_), .Y(mai_mai_n238_));
  NO3        m0216(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n239_));
  NAi21      m0217(.An(i_4_), .B(i_3_), .Y(mai_mai_n240_));
  NO2        m0218(.A(mai_mai_n240_), .B(mai_mai_n74_), .Y(mai_mai_n241_));
  NO2        m0219(.A(i_0_), .B(i_6_), .Y(mai_mai_n242_));
  NOi41      m0220(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n243_));
  NA2        m0221(.A(mai_mai_n243_), .B(mai_mai_n242_), .Y(mai_mai_n244_));
  NO2        m0222(.A(mai_mai_n237_), .B(mai_mai_n181_), .Y(mai_mai_n245_));
  NAi21      m0223(.An(mai_mai_n244_), .B(mai_mai_n245_), .Y(mai_mai_n246_));
  INV        m0224(.A(mai_mai_n246_), .Y(mai_mai_n247_));
  AOI220     m0225(.A0(mai_mai_n247_), .A1(mai_mai_n40_), .B0(mai_mai_n238_), .B1(mai_mai_n205_), .Y(mai_mai_n248_));
  NO2        m0226(.A(i_11_), .B(mai_mai_n223_), .Y(mai_mai_n249_));
  NOi21      m0227(.An(i_1_), .B(i_6_), .Y(mai_mai_n250_));
  NAi21      m0228(.An(i_3_), .B(i_7_), .Y(mai_mai_n251_));
  NO2        m0229(.A(mai_mai_n48_), .B(mai_mai_n25_), .Y(mai_mai_n252_));
  NO2        m0230(.A(i_12_), .B(i_3_), .Y(mai_mai_n253_));
  NA2        m0231(.A(mai_mai_n72_), .B(i_5_), .Y(mai_mai_n254_));
  NA3        m0232(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n255_));
  INV        m0233(.A(mai_mai_n141_), .Y(mai_mai_n256_));
  NA2        m0234(.A(mai_mai_n235_), .B(i_13_), .Y(mai_mai_n257_));
  NO2        m0235(.A(mai_mai_n257_), .B(mai_mai_n74_), .Y(mai_mai_n258_));
  NA2        m0236(.A(mai_mai_n258_), .B(mai_mai_n256_), .Y(mai_mai_n259_));
  NO2        m0237(.A(mai_mai_n231_), .B(mai_mai_n37_), .Y(mai_mai_n260_));
  NA2        m0238(.A(i_12_), .B(i_6_), .Y(mai_mai_n261_));
  OR2        m0239(.A(i_13_), .B(i_9_), .Y(mai_mai_n262_));
  NO3        m0240(.A(mai_mai_n262_), .B(mai_mai_n261_), .C(mai_mai_n48_), .Y(mai_mai_n263_));
  NO2        m0241(.A(mai_mai_n240_), .B(i_2_), .Y(mai_mai_n264_));
  NA3        m0242(.A(mai_mai_n264_), .B(mai_mai_n263_), .C(mai_mai_n44_), .Y(mai_mai_n265_));
  NA2        m0243(.A(mai_mai_n249_), .B(i_9_), .Y(mai_mai_n266_));
  NA3        m0244(.A(mai_mai_n254_), .B(mai_mai_n155_), .C(mai_mai_n63_), .Y(mai_mai_n267_));
  OAI210     m0245(.A0(mai_mai_n267_), .A1(mai_mai_n266_), .B0(mai_mai_n265_), .Y(mai_mai_n268_));
  NA2        m0246(.A(mai_mai_n152_), .B(mai_mai_n62_), .Y(mai_mai_n269_));
  NO3        m0247(.A(i_11_), .B(mai_mai_n223_), .C(mai_mai_n25_), .Y(mai_mai_n270_));
  NO2        m0248(.A(mai_mai_n251_), .B(i_8_), .Y(mai_mai_n271_));
  NO2        m0249(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n272_));
  NA3        m0250(.A(mai_mai_n272_), .B(mai_mai_n271_), .C(mai_mai_n270_), .Y(mai_mai_n273_));
  NO3        m0251(.A(mai_mai_n26_), .B(mai_mai_n83_), .C(i_5_), .Y(mai_mai_n274_));
  NA3        m0252(.A(mai_mai_n274_), .B(mai_mai_n260_), .C(mai_mai_n224_), .Y(mai_mai_n275_));
  AOI210     m0253(.A0(mai_mai_n275_), .A1(mai_mai_n273_), .B0(mai_mai_n269_), .Y(mai_mai_n276_));
  AOI210     m0254(.A0(mai_mai_n268_), .A1(mai_mai_n260_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  NA4        m0255(.A(mai_mai_n277_), .B(mai_mai_n259_), .C(mai_mai_n248_), .D(mai_mai_n227_), .Y(mai_mai_n278_));
  NO3        m0256(.A(i_12_), .B(mai_mai_n223_), .C(mai_mai_n37_), .Y(mai_mai_n279_));
  INV        m0257(.A(mai_mai_n279_), .Y(mai_mai_n280_));
  NA2        m0258(.A(i_8_), .B(mai_mai_n98_), .Y(mai_mai_n281_));
  NO3        m0259(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n282_));
  AOI220     m0260(.A0(mai_mai_n282_), .A1(mai_mai_n195_), .B0(mai_mai_n161_), .B1(mai_mai_n233_), .Y(mai_mai_n283_));
  NO2        m0261(.A(mai_mai_n283_), .B(mai_mai_n281_), .Y(mai_mai_n284_));
  NO2        m0262(.A(mai_mai_n237_), .B(i_0_), .Y(mai_mai_n285_));
  AOI220     m0263(.A0(mai_mai_n285_), .A1(mai_mai_n193_), .B0(i_1_), .B1(mai_mai_n140_), .Y(mai_mai_n286_));
  NA2        m0264(.A(mai_mai_n272_), .B(mai_mai_n26_), .Y(mai_mai_n287_));
  NO2        m0265(.A(mai_mai_n287_), .B(mai_mai_n286_), .Y(mai_mai_n288_));
  NA2        m0266(.A(i_0_), .B(i_1_), .Y(mai_mai_n289_));
  NO2        m0267(.A(mai_mai_n289_), .B(i_2_), .Y(mai_mai_n290_));
  NO2        m0268(.A(mai_mai_n58_), .B(i_6_), .Y(mai_mai_n291_));
  NA3        m0269(.A(mai_mai_n291_), .B(mai_mai_n290_), .C(mai_mai_n161_), .Y(mai_mai_n292_));
  OAI210     m0270(.A0(mai_mai_n163_), .A1(mai_mai_n141_), .B0(mai_mai_n292_), .Y(mai_mai_n293_));
  NO3        m0271(.A(mai_mai_n293_), .B(mai_mai_n288_), .C(mai_mai_n284_), .Y(mai_mai_n294_));
  NO2        m0272(.A(i_3_), .B(i_10_), .Y(mai_mai_n295_));
  NA3        m0273(.A(mai_mai_n295_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n296_));
  NO2        m0274(.A(i_2_), .B(mai_mai_n98_), .Y(mai_mai_n297_));
  NA2        m0275(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n298_));
  NO2        m0276(.A(mai_mai_n298_), .B(i_8_), .Y(mai_mai_n299_));
  NA3        m0277(.A(mai_mai_n217_), .B(mai_mai_n299_), .C(mai_mai_n297_), .Y(mai_mai_n300_));
  AN2        m0278(.A(i_3_), .B(i_10_), .Y(mai_mai_n301_));
  NA4        m0279(.A(mai_mai_n301_), .B(mai_mai_n197_), .C(mai_mai_n174_), .D(mai_mai_n172_), .Y(mai_mai_n302_));
  NO2        m0280(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n303_));
  NO2        m0281(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n304_));
  OR2        m0282(.A(mai_mai_n300_), .B(mai_mai_n296_), .Y(mai_mai_n305_));
  OAI220     m0283(.A0(mai_mai_n305_), .A1(i_6_), .B0(mai_mai_n294_), .B1(mai_mai_n280_), .Y(mai_mai_n306_));
  NO4        m0284(.A(mai_mai_n306_), .B(mai_mai_n278_), .C(mai_mai_n213_), .D(mai_mai_n166_), .Y(mai_mai_n307_));
  NO3        m0285(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n308_));
  NO2        m0286(.A(mai_mai_n58_), .B(mai_mai_n83_), .Y(mai_mai_n309_));
  NA2        m0287(.A(mai_mai_n285_), .B(mai_mai_n309_), .Y(mai_mai_n310_));
  NO3        m0288(.A(i_6_), .B(mai_mai_n192_), .C(i_7_), .Y(mai_mai_n311_));
  NA2        m0289(.A(mai_mai_n311_), .B(mai_mai_n197_), .Y(mai_mai_n312_));
  AOI210     m0290(.A0(mai_mai_n312_), .A1(mai_mai_n310_), .B0(mai_mai_n167_), .Y(mai_mai_n313_));
  NO2        m0291(.A(i_2_), .B(i_3_), .Y(mai_mai_n314_));
  OR2        m0292(.A(i_0_), .B(i_5_), .Y(mai_mai_n315_));
  NA2        m0293(.A(mai_mai_n217_), .B(mai_mai_n315_), .Y(mai_mai_n316_));
  NA4        m0294(.A(mai_mai_n316_), .B(mai_mai_n232_), .C(mai_mai_n314_), .D(i_1_), .Y(mai_mai_n317_));
  NA3        m0295(.A(mai_mai_n285_), .B(mai_mai_n161_), .C(mai_mai_n110_), .Y(mai_mai_n318_));
  NAi21      m0296(.An(i_8_), .B(i_7_), .Y(mai_mai_n319_));
  NO2        m0297(.A(mai_mai_n319_), .B(i_6_), .Y(mai_mai_n320_));
  NO2        m0298(.A(mai_mai_n155_), .B(mai_mai_n46_), .Y(mai_mai_n321_));
  NA3        m0299(.A(mai_mai_n321_), .B(mai_mai_n320_), .C(mai_mai_n161_), .Y(mai_mai_n322_));
  NA3        m0300(.A(mai_mai_n322_), .B(mai_mai_n318_), .C(mai_mai_n317_), .Y(mai_mai_n323_));
  OAI210     m0301(.A0(mai_mai_n323_), .A1(mai_mai_n313_), .B0(i_4_), .Y(mai_mai_n324_));
  NO2        m0302(.A(i_12_), .B(i_10_), .Y(mai_mai_n325_));
  NOi21      m0303(.An(i_5_), .B(i_0_), .Y(mai_mai_n326_));
  NO3        m0304(.A(mai_mai_n298_), .B(mai_mai_n326_), .C(mai_mai_n126_), .Y(mai_mai_n327_));
  NA4        m0305(.A(mai_mai_n82_), .B(mai_mai_n36_), .C(mai_mai_n83_), .D(i_8_), .Y(mai_mai_n328_));
  NA2        m0306(.A(mai_mai_n327_), .B(mai_mai_n325_), .Y(mai_mai_n329_));
  NO2        m0307(.A(i_6_), .B(i_8_), .Y(mai_mai_n330_));
  NOi21      m0308(.An(i_0_), .B(i_2_), .Y(mai_mai_n331_));
  AN2        m0309(.A(mai_mai_n331_), .B(mai_mai_n330_), .Y(mai_mai_n332_));
  NO2        m0310(.A(i_1_), .B(i_7_), .Y(mai_mai_n333_));
  AO220      m0311(.A0(mai_mai_n333_), .A1(mai_mai_n332_), .B0(mai_mai_n320_), .B1(mai_mai_n233_), .Y(mai_mai_n334_));
  NA3        m0312(.A(mai_mai_n334_), .B(i_4_), .C(i_5_), .Y(mai_mai_n335_));
  NA3        m0313(.A(mai_mai_n335_), .B(mai_mai_n329_), .C(mai_mai_n324_), .Y(mai_mai_n336_));
  NO3        m0314(.A(mai_mai_n231_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n337_));
  NO3        m0315(.A(mai_mai_n319_), .B(i_2_), .C(i_1_), .Y(mai_mai_n338_));
  OAI210     m0316(.A0(mai_mai_n338_), .A1(mai_mai_n337_), .B0(i_6_), .Y(mai_mai_n339_));
  NA3        m0317(.A(mai_mai_n250_), .B(mai_mai_n297_), .C(mai_mai_n192_), .Y(mai_mai_n340_));
  AOI210     m0318(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(mai_mai_n316_), .Y(mai_mai_n341_));
  NO2        m0319(.A(mai_mai_n100_), .B(mai_mai_n122_), .Y(mai_mai_n342_));
  OAI210     m0320(.A0(mai_mai_n342_), .A1(mai_mai_n341_), .B0(i_3_), .Y(mai_mai_n343_));
  INV        m0321(.A(mai_mai_n82_), .Y(mai_mai_n344_));
  NO2        m0322(.A(mai_mai_n289_), .B(mai_mai_n80_), .Y(mai_mai_n345_));
  NA2        m0323(.A(mai_mai_n345_), .B(mai_mai_n130_), .Y(mai_mai_n346_));
  NO2        m0324(.A(mai_mai_n90_), .B(mai_mai_n192_), .Y(mai_mai_n347_));
  NA3        m0325(.A(mai_mai_n217_), .B(mai_mai_n347_), .C(mai_mai_n62_), .Y(mai_mai_n348_));
  AOI210     m0326(.A0(mai_mai_n348_), .A1(mai_mai_n346_), .B0(mai_mai_n344_), .Y(mai_mai_n349_));
  NO2        m0327(.A(mai_mai_n192_), .B(i_9_), .Y(mai_mai_n350_));
  NA2        m0328(.A(mai_mai_n350_), .B(mai_mai_n155_), .Y(mai_mai_n351_));
  NO2        m0329(.A(mai_mai_n351_), .B(mai_mai_n46_), .Y(mai_mai_n352_));
  NO3        m0330(.A(mai_mai_n352_), .B(mai_mai_n349_), .C(mai_mai_n288_), .Y(mai_mai_n353_));
  AOI210     m0331(.A0(mai_mai_n353_), .A1(mai_mai_n343_), .B0(mai_mai_n160_), .Y(mai_mai_n354_));
  AOI210     m0332(.A0(mai_mai_n336_), .A1(mai_mai_n308_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NOi32      m0333(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n356_));
  INV        m0334(.A(mai_mai_n356_), .Y(mai_mai_n357_));
  NAi21      m0335(.An(i_0_), .B(i_6_), .Y(mai_mai_n358_));
  NAi21      m0336(.An(i_1_), .B(i_5_), .Y(mai_mai_n359_));
  NA2        m0337(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n360_));
  NA2        m0338(.A(mai_mai_n360_), .B(mai_mai_n25_), .Y(mai_mai_n361_));
  OAI210     m0339(.A0(mai_mai_n361_), .A1(mai_mai_n157_), .B0(mai_mai_n244_), .Y(mai_mai_n362_));
  NAi41      m0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n363_));
  OAI220     m0341(.A0(mai_mai_n363_), .A1(mai_mai_n359_), .B0(mai_mai_n219_), .B1(mai_mai_n157_), .Y(mai_mai_n364_));
  AOI210     m0342(.A0(mai_mai_n363_), .A1(mai_mai_n157_), .B0(mai_mai_n155_), .Y(mai_mai_n365_));
  NOi32      m0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n366_));
  NAi21      m0344(.An(i_6_), .B(i_1_), .Y(mai_mai_n367_));
  NA3        m0345(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(mai_mai_n46_), .Y(mai_mai_n368_));
  NO2        m0346(.A(mai_mai_n368_), .B(i_0_), .Y(mai_mai_n369_));
  OR3        m0347(.A(mai_mai_n369_), .B(mai_mai_n365_), .C(mai_mai_n364_), .Y(mai_mai_n370_));
  NO2        m0348(.A(i_1_), .B(mai_mai_n98_), .Y(mai_mai_n371_));
  NAi21      m0349(.An(i_3_), .B(i_4_), .Y(mai_mai_n372_));
  AN2        m0350(.A(i_6_), .B(i_7_), .Y(mai_mai_n373_));
  NA2        m0351(.A(i_2_), .B(i_7_), .Y(mai_mai_n374_));
  NO2        m0352(.A(mai_mai_n372_), .B(i_10_), .Y(mai_mai_n375_));
  AOI210     m0353(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n376_));
  OAI210     m0354(.A0(mai_mai_n376_), .A1(mai_mai_n187_), .B0(mai_mai_n375_), .Y(mai_mai_n377_));
  AOI220     m0355(.A0(mai_mai_n375_), .A1(mai_mai_n333_), .B0(mai_mai_n236_), .B1(mai_mai_n187_), .Y(mai_mai_n378_));
  AOI210     m0356(.A0(mai_mai_n378_), .A1(mai_mai_n377_), .B0(i_5_), .Y(mai_mai_n379_));
  NO3        m0357(.A(mai_mai_n379_), .B(mai_mai_n370_), .C(mai_mai_n362_), .Y(mai_mai_n380_));
  NO2        m0358(.A(mai_mai_n380_), .B(mai_mai_n357_), .Y(mai_mai_n381_));
  NO2        m0359(.A(mai_mai_n58_), .B(mai_mai_n25_), .Y(mai_mai_n382_));
  AN2        m0360(.A(i_12_), .B(i_5_), .Y(mai_mai_n383_));
  NO2        m0361(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n384_));
  NA2        m0362(.A(mai_mai_n384_), .B(mai_mai_n383_), .Y(mai_mai_n385_));
  NO2        m0363(.A(i_11_), .B(i_6_), .Y(mai_mai_n386_));
  NA3        m0364(.A(mai_mai_n386_), .B(mai_mai_n321_), .C(mai_mai_n223_), .Y(mai_mai_n387_));
  NO2        m0365(.A(mai_mai_n387_), .B(mai_mai_n385_), .Y(mai_mai_n388_));
  NO2        m0366(.A(mai_mai_n240_), .B(i_5_), .Y(mai_mai_n389_));
  NO2        m0367(.A(i_5_), .B(i_10_), .Y(mai_mai_n390_));
  AOI220     m0368(.A0(mai_mai_n390_), .A1(mai_mai_n264_), .B0(mai_mai_n389_), .B1(mai_mai_n197_), .Y(mai_mai_n391_));
  NA2        m0369(.A(mai_mai_n142_), .B(mai_mai_n45_), .Y(mai_mai_n392_));
  NO2        m0370(.A(mai_mai_n392_), .B(mai_mai_n391_), .Y(mai_mai_n393_));
  OAI210     m0371(.A0(mai_mai_n393_), .A1(mai_mai_n388_), .B0(mai_mai_n382_), .Y(mai_mai_n394_));
  NO2        m0372(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n395_));
  NO2        m0373(.A(mai_mai_n148_), .B(mai_mai_n83_), .Y(mai_mai_n396_));
  OAI210     m0374(.A0(mai_mai_n396_), .A1(mai_mai_n388_), .B0(mai_mai_n395_), .Y(mai_mai_n397_));
  NO3        m0375(.A(mai_mai_n83_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n398_));
  NO2        m0376(.A(i_11_), .B(i_12_), .Y(mai_mai_n399_));
  NA2        m0377(.A(mai_mai_n390_), .B(mai_mai_n235_), .Y(mai_mai_n400_));
  NA3        m0378(.A(mai_mai_n110_), .B(i_4_), .C(i_11_), .Y(mai_mai_n401_));
  OAI220     m0379(.A0(mai_mai_n401_), .A1(mai_mai_n219_), .B0(mai_mai_n400_), .B1(mai_mai_n328_), .Y(mai_mai_n402_));
  NAi21      m0380(.An(i_13_), .B(i_0_), .Y(mai_mai_n403_));
  NO2        m0381(.A(mai_mai_n403_), .B(mai_mai_n237_), .Y(mai_mai_n404_));
  NA2        m0382(.A(mai_mai_n402_), .B(mai_mai_n404_), .Y(mai_mai_n405_));
  NA3        m0383(.A(mai_mai_n405_), .B(mai_mai_n397_), .C(mai_mai_n394_), .Y(mai_mai_n406_));
  NO2        m0384(.A(i_0_), .B(i_11_), .Y(mai_mai_n407_));
  AN2        m0385(.A(i_1_), .B(i_6_), .Y(mai_mai_n408_));
  NOi21      m0386(.An(i_2_), .B(i_12_), .Y(mai_mai_n409_));
  NA2        m0387(.A(mai_mai_n409_), .B(mai_mai_n408_), .Y(mai_mai_n410_));
  INV        m0388(.A(mai_mai_n410_), .Y(mai_mai_n411_));
  NA2        m0389(.A(mai_mai_n140_), .B(i_9_), .Y(mai_mai_n412_));
  NO2        m0390(.A(mai_mai_n412_), .B(i_4_), .Y(mai_mai_n413_));
  NA2        m0391(.A(mai_mai_n411_), .B(mai_mai_n413_), .Y(mai_mai_n414_));
  OR2        m0392(.A(i_13_), .B(i_10_), .Y(mai_mai_n415_));
  NO2        m0393(.A(mai_mai_n170_), .B(mai_mai_n121_), .Y(mai_mai_n416_));
  OR2        m0394(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n417_));
  NO2        m0395(.A(mai_mai_n98_), .B(mai_mai_n25_), .Y(mai_mai_n418_));
  NA2        m0396(.A(mai_mai_n272_), .B(mai_mai_n209_), .Y(mai_mai_n419_));
  NO2        m0397(.A(mai_mai_n419_), .B(mai_mai_n417_), .Y(mai_mai_n420_));
  INV        m0398(.A(mai_mai_n420_), .Y(mai_mai_n421_));
  AOI210     m0399(.A0(mai_mai_n421_), .A1(mai_mai_n414_), .B0(mai_mai_n26_), .Y(mai_mai_n422_));
  NA2        m0400(.A(mai_mai_n318_), .B(mai_mai_n317_), .Y(mai_mai_n423_));
  AOI220     m0401(.A0(mai_mai_n291_), .A1(mai_mai_n282_), .B0(mai_mai_n285_), .B1(mai_mai_n309_), .Y(mai_mai_n424_));
  NO2        m0402(.A(mai_mai_n424_), .B(mai_mai_n167_), .Y(mai_mai_n425_));
  NO2        m0403(.A(mai_mai_n181_), .B(mai_mai_n83_), .Y(mai_mai_n426_));
  AOI220     m0404(.A0(mai_mai_n426_), .A1(mai_mai_n290_), .B0(mai_mai_n274_), .B1(mai_mai_n209_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n427_), .B(mai_mai_n281_), .Y(mai_mai_n428_));
  NO3        m0406(.A(mai_mai_n428_), .B(mai_mai_n425_), .C(mai_mai_n423_), .Y(mai_mai_n429_));
  NA2        m0407(.A(mai_mai_n195_), .B(mai_mai_n93_), .Y(mai_mai_n430_));
  NA3        m0408(.A(mai_mai_n321_), .B(mai_mai_n161_), .C(mai_mai_n83_), .Y(mai_mai_n431_));
  AOI210     m0409(.A0(mai_mai_n431_), .A1(mai_mai_n430_), .B0(mai_mai_n319_), .Y(mai_mai_n432_));
  NA2        m0410(.A(mai_mai_n291_), .B(mai_mai_n233_), .Y(mai_mai_n433_));
  NO2        m0411(.A(mai_mai_n433_), .B(mai_mai_n181_), .Y(mai_mai_n434_));
  NO2        m0412(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n435_));
  NA3        m0413(.A(mai_mai_n333_), .B(mai_mai_n332_), .C(mai_mai_n435_), .Y(mai_mai_n436_));
  NA2        m0414(.A(mai_mai_n311_), .B(mai_mai_n316_), .Y(mai_mai_n437_));
  OAI210     m0415(.A0(mai_mai_n437_), .A1(mai_mai_n188_), .B0(mai_mai_n436_), .Y(mai_mai_n438_));
  NO3        m0416(.A(mai_mai_n438_), .B(mai_mai_n434_), .C(mai_mai_n432_), .Y(mai_mai_n439_));
  AOI210     m0417(.A0(mai_mai_n439_), .A1(mai_mai_n429_), .B0(mai_mai_n266_), .Y(mai_mai_n440_));
  NO4        m0418(.A(mai_mai_n440_), .B(mai_mai_n422_), .C(mai_mai_n406_), .D(mai_mai_n381_), .Y(mai_mai_n441_));
  NO2        m0419(.A(mai_mai_n62_), .B(i_4_), .Y(mai_mai_n442_));
  NO2        m0420(.A(mai_mai_n72_), .B(i_13_), .Y(mai_mai_n443_));
  NA3        m0421(.A(mai_mai_n443_), .B(mai_mai_n442_), .C(i_2_), .Y(mai_mai_n444_));
  NO2        m0422(.A(i_10_), .B(i_9_), .Y(mai_mai_n445_));
  NAi21      m0423(.An(i_12_), .B(i_8_), .Y(mai_mai_n446_));
  NO2        m0424(.A(mai_mai_n446_), .B(i_3_), .Y(mai_mai_n447_));
  NA2        m0425(.A(mai_mai_n447_), .B(mai_mai_n445_), .Y(mai_mai_n448_));
  NO2        m0426(.A(mai_mai_n46_), .B(i_4_), .Y(mai_mai_n449_));
  NA2        m0427(.A(mai_mai_n449_), .B(mai_mai_n101_), .Y(mai_mai_n450_));
  OAI220     m0428(.A0(mai_mai_n450_), .A1(mai_mai_n204_), .B0(mai_mai_n448_), .B1(mai_mai_n444_), .Y(mai_mai_n451_));
  NA2        m0429(.A(mai_mai_n304_), .B(i_0_), .Y(mai_mai_n452_));
  NO3        m0430(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n453_));
  NA2        m0431(.A(mai_mai_n261_), .B(mai_mai_n94_), .Y(mai_mai_n454_));
  NA2        m0432(.A(mai_mai_n454_), .B(mai_mai_n453_), .Y(mai_mai_n455_));
  NA2        m0433(.A(i_8_), .B(i_9_), .Y(mai_mai_n456_));
  NO2        m0434(.A(mai_mai_n455_), .B(mai_mai_n452_), .Y(mai_mai_n457_));
  NA2        m0435(.A(mai_mai_n249_), .B(mai_mai_n303_), .Y(mai_mai_n458_));
  NO3        m0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n459_));
  AOI210     m0437(.A0(mai_mai_n253_), .A1(mai_mai_n187_), .B0(mai_mai_n459_), .Y(mai_mai_n460_));
  NA3        m0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n461_));
  NA4        m0439(.A(mai_mai_n143_), .B(mai_mai_n113_), .C(mai_mai_n79_), .D(mai_mai_n23_), .Y(mai_mai_n462_));
  OAI220     m0440(.A0(mai_mai_n462_), .A1(mai_mai_n461_), .B0(mai_mai_n460_), .B1(mai_mai_n458_), .Y(mai_mai_n463_));
  NO3        m0441(.A(mai_mai_n463_), .B(mai_mai_n457_), .C(mai_mai_n451_), .Y(mai_mai_n464_));
  OR2        m0442(.A(mai_mai_n289_), .B(mai_mai_n206_), .Y(mai_mai_n465_));
  OA210      m0443(.A0(mai_mai_n351_), .A1(mai_mai_n98_), .B0(mai_mai_n292_), .Y(mai_mai_n466_));
  OA220      m0444(.A0(mai_mai_n466_), .A1(mai_mai_n160_), .B0(mai_mai_n465_), .B1(mai_mai_n230_), .Y(mai_mai_n467_));
  NA2        m0445(.A(mai_mai_n93_), .B(i_13_), .Y(mai_mai_n468_));
  NA2        m0446(.A(mai_mai_n426_), .B(mai_mai_n382_), .Y(mai_mai_n469_));
  NO2        m0447(.A(i_2_), .B(i_13_), .Y(mai_mai_n470_));
  NA3        m0448(.A(mai_mai_n470_), .B(mai_mai_n159_), .C(mai_mai_n96_), .Y(mai_mai_n471_));
  OAI220     m0449(.A0(mai_mai_n471_), .A1(mai_mai_n235_), .B0(mai_mai_n469_), .B1(mai_mai_n468_), .Y(mai_mai_n472_));
  NO3        m0450(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n473_));
  NO2        m0451(.A(i_6_), .B(i_7_), .Y(mai_mai_n474_));
  NA2        m0452(.A(mai_mai_n474_), .B(mai_mai_n473_), .Y(mai_mai_n475_));
  NO2        m0453(.A(i_11_), .B(i_1_), .Y(mai_mai_n476_));
  OR2        m0454(.A(i_11_), .B(i_8_), .Y(mai_mai_n477_));
  NOi21      m0455(.An(i_2_), .B(i_7_), .Y(mai_mai_n478_));
  NAi31      m0456(.An(mai_mai_n477_), .B(mai_mai_n478_), .C(i_0_), .Y(mai_mai_n479_));
  NO2        m0457(.A(mai_mai_n415_), .B(i_6_), .Y(mai_mai_n480_));
  NA3        m0458(.A(mai_mai_n480_), .B(mai_mai_n442_), .C(mai_mai_n74_), .Y(mai_mai_n481_));
  NO2        m0459(.A(mai_mai_n481_), .B(mai_mai_n479_), .Y(mai_mai_n482_));
  NO2        m0460(.A(i_3_), .B(mai_mai_n192_), .Y(mai_mai_n483_));
  NO2        m0461(.A(i_6_), .B(i_10_), .Y(mai_mai_n484_));
  NA4        m0462(.A(mai_mai_n484_), .B(mai_mai_n308_), .C(mai_mai_n483_), .D(mai_mai_n235_), .Y(mai_mai_n485_));
  NO2        m0463(.A(mai_mai_n485_), .B(mai_mai_n153_), .Y(mai_mai_n486_));
  NA2        m0464(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n487_));
  NO2        m0465(.A(mai_mai_n155_), .B(i_3_), .Y(mai_mai_n488_));
  NAi31      m0466(.An(mai_mai_n487_), .B(mai_mai_n488_), .C(mai_mai_n224_), .Y(mai_mai_n489_));
  NA3        m0467(.A(mai_mai_n395_), .B(mai_mai_n177_), .C(mai_mai_n147_), .Y(mai_mai_n490_));
  NA2        m0468(.A(mai_mai_n490_), .B(mai_mai_n489_), .Y(mai_mai_n491_));
  NO4        m0469(.A(mai_mai_n491_), .B(mai_mai_n486_), .C(mai_mai_n482_), .D(mai_mai_n472_), .Y(mai_mai_n492_));
  NA2        m0470(.A(mai_mai_n453_), .B(mai_mai_n383_), .Y(mai_mai_n493_));
  NA2        m0471(.A(mai_mai_n459_), .B(mai_mai_n390_), .Y(mai_mai_n494_));
  OAI220     m0472(.A0(mai_mai_n494_), .A1(mai_mai_n222_), .B0(mai_mai_n493_), .B1(mai_mai_n56_), .Y(mai_mai_n495_));
  NAi21      m0473(.An(mai_mai_n215_), .B(mai_mai_n399_), .Y(mai_mai_n496_));
  NA2        m0474(.A(mai_mai_n333_), .B(mai_mai_n217_), .Y(mai_mai_n497_));
  NO2        m0475(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n498_));
  NO2        m0476(.A(i_0_), .B(mai_mai_n83_), .Y(mai_mai_n499_));
  NA3        m0477(.A(mai_mai_n499_), .B(mai_mai_n498_), .C(mai_mai_n140_), .Y(mai_mai_n500_));
  OR3        m0478(.A(mai_mai_n298_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n501_));
  OAI220     m0479(.A0(mai_mai_n501_), .A1(mai_mai_n500_), .B0(mai_mai_n497_), .B1(mai_mai_n496_), .Y(mai_mai_n502_));
  NA4        m0480(.A(mai_mai_n301_), .B(mai_mai_n221_), .C(mai_mai_n72_), .D(mai_mai_n235_), .Y(mai_mai_n503_));
  NO2        m0481(.A(mai_mai_n503_), .B(mai_mai_n475_), .Y(mai_mai_n504_));
  NO3        m0482(.A(mai_mai_n504_), .B(mai_mai_n502_), .C(mai_mai_n495_), .Y(mai_mai_n505_));
  NA4        m0483(.A(mai_mai_n505_), .B(mai_mai_n492_), .C(mai_mai_n467_), .D(mai_mai_n464_), .Y(mai_mai_n506_));
  NA2        m0484(.A(mai_mai_n301_), .B(mai_mai_n174_), .Y(mai_mai_n507_));
  OAI210     m0485(.A0(mai_mai_n296_), .A1(mai_mai_n179_), .B0(mai_mai_n507_), .Y(mai_mai_n508_));
  AN2        m0486(.A(mai_mai_n282_), .B(mai_mai_n232_), .Y(mai_mai_n509_));
  NA2        m0487(.A(mai_mai_n509_), .B(mai_mai_n508_), .Y(mai_mai_n510_));
  NA2        m0488(.A(mai_mai_n120_), .B(mai_mai_n109_), .Y(mai_mai_n511_));
  AN2        m0489(.A(mai_mai_n511_), .B(mai_mai_n453_), .Y(mai_mai_n512_));
  NA2        m0490(.A(mai_mai_n308_), .B(mai_mai_n162_), .Y(mai_mai_n513_));
  OAI210     m0491(.A0(mai_mai_n513_), .A1(mai_mai_n230_), .B0(mai_mai_n302_), .Y(mai_mai_n514_));
  AOI220     m0492(.A0(mai_mai_n514_), .A1(mai_mai_n320_), .B0(mai_mai_n512_), .B1(mai_mai_n304_), .Y(mai_mai_n515_));
  NA4        m0493(.A(mai_mai_n443_), .B(mai_mai_n442_), .C(mai_mai_n202_), .D(i_2_), .Y(mai_mai_n516_));
  INV        m0494(.A(mai_mai_n516_), .Y(mai_mai_n517_));
  NA2        m0495(.A(mai_mai_n356_), .B(mai_mai_n72_), .Y(mai_mai_n518_));
  NA2        m0496(.A(mai_mai_n373_), .B(mai_mai_n366_), .Y(mai_mai_n519_));
  NO2        m0497(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n520_));
  NA2        m0498(.A(mai_mai_n39_), .B(i_13_), .Y(mai_mai_n521_));
  INV        m0499(.A(mai_mai_n521_), .Y(mai_mai_n522_));
  AOI210     m0500(.A0(mai_mai_n517_), .A1(mai_mai_n203_), .B0(mai_mai_n522_), .Y(mai_mai_n523_));
  NA2        m0501(.A(mai_mai_n254_), .B(mai_mai_n63_), .Y(mai_mai_n524_));
  OAI210     m0502(.A0(i_8_), .A1(mai_mai_n524_), .B0(mai_mai_n132_), .Y(mai_mai_n525_));
  NO2        m0503(.A(i_7_), .B(mai_mai_n198_), .Y(mai_mai_n526_));
  OR2        m0504(.A(mai_mai_n181_), .B(i_4_), .Y(mai_mai_n527_));
  NO2        m0505(.A(mai_mai_n527_), .B(mai_mai_n83_), .Y(mai_mai_n528_));
  AOI220     m0506(.A0(mai_mai_n528_), .A1(mai_mai_n526_), .B0(mai_mai_n525_), .B1(mai_mai_n416_), .Y(mai_mai_n529_));
  NA4        m0507(.A(mai_mai_n529_), .B(mai_mai_n523_), .C(mai_mai_n515_), .D(mai_mai_n510_), .Y(mai_mai_n530_));
  NA2        m0508(.A(mai_mai_n389_), .B(mai_mai_n290_), .Y(mai_mai_n531_));
  NA2        m0509(.A(mai_mai_n385_), .B(mai_mai_n531_), .Y(mai_mai_n532_));
  NA2        m0510(.A(mai_mai_n1047_), .B(mai_mai_n223_), .Y(mai_mai_n533_));
  NA2        m0511(.A(mai_mai_n484_), .B(mai_mai_n27_), .Y(mai_mai_n534_));
  NO2        m0512(.A(mai_mai_n534_), .B(mai_mai_n533_), .Y(mai_mai_n535_));
  NOi31      m0513(.An(mai_mai_n311_), .B(mai_mai_n415_), .C(mai_mai_n38_), .Y(mai_mai_n536_));
  OAI210     m0514(.A0(mai_mai_n536_), .A1(mai_mai_n535_), .B0(mai_mai_n532_), .Y(mai_mai_n537_));
  NO2        m0515(.A(i_8_), .B(i_7_), .Y(mai_mai_n538_));
  OAI210     m0516(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n539_));
  NA2        m0517(.A(mai_mai_n539_), .B(mai_mai_n221_), .Y(mai_mai_n540_));
  OAI220     m0518(.A0(mai_mai_n46_), .A1(mai_mai_n527_), .B0(mai_mai_n540_), .B1(mai_mai_n240_), .Y(mai_mai_n541_));
  NA2        m0519(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n542_));
  NO2        m0520(.A(mai_mai_n542_), .B(i_6_), .Y(mai_mai_n543_));
  NA3        m0521(.A(mai_mai_n543_), .B(mai_mai_n541_), .C(mai_mai_n538_), .Y(mai_mai_n544_));
  AOI220     m0522(.A0(mai_mai_n426_), .A1(mai_mai_n321_), .B0(mai_mai_n245_), .B1(mai_mai_n242_), .Y(mai_mai_n545_));
  OAI220     m0523(.A0(mai_mai_n545_), .A1(mai_mai_n257_), .B0(mai_mai_n468_), .B1(mai_mai_n131_), .Y(mai_mai_n546_));
  NA2        m0524(.A(mai_mai_n546_), .B(mai_mai_n260_), .Y(mai_mai_n547_));
  NOi31      m0525(.An(mai_mai_n285_), .B(mai_mai_n296_), .C(mai_mai_n179_), .Y(mai_mai_n548_));
  NA3        m0526(.A(mai_mai_n301_), .B(mai_mai_n172_), .C(mai_mai_n93_), .Y(mai_mai_n549_));
  NO2        m0527(.A(mai_mai_n220_), .B(mai_mai_n44_), .Y(mai_mai_n550_));
  NO2        m0528(.A(mai_mai_n155_), .B(i_5_), .Y(mai_mai_n551_));
  NA2        m0529(.A(mai_mai_n551_), .B(mai_mai_n314_), .Y(mai_mai_n552_));
  OAI210     m0530(.A0(mai_mai_n552_), .A1(mai_mai_n550_), .B0(mai_mai_n549_), .Y(mai_mai_n553_));
  OAI210     m0531(.A0(mai_mai_n553_), .A1(mai_mai_n548_), .B0(mai_mai_n459_), .Y(mai_mai_n554_));
  NA4        m0532(.A(mai_mai_n554_), .B(mai_mai_n547_), .C(mai_mai_n544_), .D(mai_mai_n537_), .Y(mai_mai_n555_));
  NA2        m0533(.A(mai_mai_n279_), .B(mai_mai_n82_), .Y(mai_mai_n556_));
  NO2        m0534(.A(mai_mai_n346_), .B(mai_mai_n556_), .Y(mai_mai_n557_));
  NA2        m0535(.A(mai_mai_n291_), .B(mai_mai_n282_), .Y(mai_mai_n558_));
  NO2        m0536(.A(mai_mai_n558_), .B(mai_mai_n171_), .Y(mai_mai_n559_));
  NA2        m0537(.A(i_0_), .B(mai_mai_n48_), .Y(mai_mai_n560_));
  NO2        m0538(.A(mai_mai_n559_), .B(mai_mai_n557_), .Y(mai_mai_n561_));
  NO4        m0539(.A(mai_mai_n250_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n562_));
  NO3        m0540(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n563_));
  NO2        m0541(.A(mai_mai_n231_), .B(mai_mai_n36_), .Y(mai_mai_n564_));
  AN2        m0542(.A(mai_mai_n564_), .B(mai_mai_n563_), .Y(mai_mai_n565_));
  OA210      m0543(.A0(mai_mai_n565_), .A1(mai_mai_n562_), .B0(mai_mai_n356_), .Y(mai_mai_n566_));
  NO2        m0544(.A(mai_mai_n415_), .B(i_1_), .Y(mai_mai_n567_));
  NOi31      m0545(.An(mai_mai_n567_), .B(mai_mai_n454_), .C(mai_mai_n72_), .Y(mai_mai_n568_));
  AN4        m0546(.A(mai_mai_n568_), .B(mai_mai_n413_), .C(mai_mai_n498_), .D(i_2_), .Y(mai_mai_n569_));
  NO2        m0547(.A(mai_mai_n424_), .B(mai_mai_n175_), .Y(mai_mai_n570_));
  NO3        m0548(.A(mai_mai_n570_), .B(mai_mai_n569_), .C(mai_mai_n566_), .Y(mai_mai_n571_));
  NOi21      m0549(.An(i_10_), .B(i_6_), .Y(mai_mai_n572_));
  NO2        m0550(.A(mai_mai_n83_), .B(mai_mai_n25_), .Y(mai_mai_n573_));
  AOI220     m0551(.A0(mai_mai_n279_), .A1(mai_mai_n573_), .B0(mai_mai_n270_), .B1(mai_mai_n572_), .Y(mai_mai_n574_));
  NO2        m0552(.A(mai_mai_n574_), .B(mai_mai_n452_), .Y(mai_mai_n575_));
  NO2        m0553(.A(mai_mai_n112_), .B(mai_mai_n23_), .Y(mai_mai_n576_));
  NA2        m0554(.A(mai_mai_n311_), .B(mai_mai_n162_), .Y(mai_mai_n577_));
  AOI220     m0555(.A0(mai_mai_n577_), .A1(mai_mai_n433_), .B0(mai_mai_n182_), .B1(mai_mai_n180_), .Y(mai_mai_n578_));
  NOi21      m0556(.An(mai_mai_n144_), .B(mai_mai_n328_), .Y(mai_mai_n579_));
  NO3        m0557(.A(mai_mai_n579_), .B(mai_mai_n578_), .C(mai_mai_n575_), .Y(mai_mai_n580_));
  NO2        m0558(.A(mai_mai_n518_), .B(mai_mai_n378_), .Y(mai_mai_n581_));
  INV        m0559(.A(mai_mai_n314_), .Y(mai_mai_n582_));
  NO2        m0560(.A(i_12_), .B(mai_mai_n83_), .Y(mai_mai_n583_));
  NA3        m0561(.A(mai_mai_n583_), .B(mai_mai_n270_), .C(mai_mai_n560_), .Y(mai_mai_n584_));
  NA3        m0562(.A(mai_mai_n386_), .B(mai_mai_n279_), .C(mai_mai_n217_), .Y(mai_mai_n585_));
  AOI210     m0563(.A0(mai_mai_n585_), .A1(mai_mai_n584_), .B0(mai_mai_n582_), .Y(mai_mai_n586_));
  NO3        m0564(.A(i_4_), .B(mai_mai_n339_), .C(mai_mai_n296_), .Y(mai_mai_n587_));
  NO3        m0565(.A(mai_mai_n587_), .B(mai_mai_n586_), .C(mai_mai_n581_), .Y(mai_mai_n588_));
  NA4        m0566(.A(mai_mai_n588_), .B(mai_mai_n580_), .C(mai_mai_n571_), .D(mai_mai_n561_), .Y(mai_mai_n589_));
  NO4        m0567(.A(mai_mai_n589_), .B(mai_mai_n555_), .C(mai_mai_n530_), .D(mai_mai_n506_), .Y(mai_mai_n590_));
  NA4        m0568(.A(mai_mai_n590_), .B(mai_mai_n441_), .C(mai_mai_n355_), .D(mai_mai_n307_), .Y(mai7));
  NO2        m0569(.A(mai_mai_n90_), .B(mai_mai_n54_), .Y(mai_mai_n592_));
  NO2        m0570(.A(mai_mai_n105_), .B(mai_mai_n87_), .Y(mai_mai_n593_));
  NA2        m0571(.A(mai_mai_n384_), .B(mai_mai_n593_), .Y(mai_mai_n594_));
  NA2        m0572(.A(i_11_), .B(mai_mai_n192_), .Y(mai_mai_n595_));
  INV        m0573(.A(mai_mai_n594_), .Y(mai_mai_n596_));
  NA3        m0574(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n597_));
  NO2        m0575(.A(mai_mai_n235_), .B(i_4_), .Y(mai_mai_n598_));
  NA2        m0576(.A(mai_mai_n598_), .B(i_8_), .Y(mai_mai_n599_));
  NO2        m0577(.A(mai_mai_n102_), .B(mai_mai_n597_), .Y(mai_mai_n600_));
  NA2        m0578(.A(i_2_), .B(mai_mai_n83_), .Y(mai_mai_n601_));
  OAI210     m0579(.A0(mai_mai_n86_), .A1(mai_mai_n202_), .B0(mai_mai_n203_), .Y(mai_mai_n602_));
  NO2        m0580(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n603_));
  NA2        m0581(.A(i_4_), .B(i_8_), .Y(mai_mai_n604_));
  AOI210     m0582(.A0(mai_mai_n604_), .A1(mai_mai_n301_), .B0(mai_mai_n603_), .Y(mai_mai_n605_));
  OAI220     m0583(.A0(mai_mai_n605_), .A1(mai_mai_n601_), .B0(mai_mai_n602_), .B1(i_13_), .Y(mai_mai_n606_));
  NO4        m0584(.A(mai_mai_n606_), .B(mai_mai_n600_), .C(mai_mai_n596_), .D(mai_mai_n592_), .Y(mai_mai_n607_));
  AOI210     m0585(.A0(mai_mai_n126_), .A1(mai_mai_n61_), .B0(i_10_), .Y(mai_mai_n608_));
  AOI210     m0586(.A0(mai_mai_n608_), .A1(mai_mai_n235_), .B0(mai_mai_n159_), .Y(mai_mai_n609_));
  OR2        m0587(.A(i_6_), .B(i_10_), .Y(mai_mai_n610_));
  NO2        m0588(.A(mai_mai_n610_), .B(mai_mai_n23_), .Y(mai_mai_n611_));
  OR3        m0589(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n612_));
  NO3        m0590(.A(mai_mai_n612_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n613_));
  INV        m0591(.A(mai_mai_n199_), .Y(mai_mai_n614_));
  NO2        m0592(.A(mai_mai_n613_), .B(mai_mai_n611_), .Y(mai_mai_n615_));
  OA220      m0593(.A0(mai_mai_n615_), .A1(mai_mai_n582_), .B0(mai_mai_n609_), .B1(mai_mai_n262_), .Y(mai_mai_n616_));
  AOI210     m0594(.A0(mai_mai_n616_), .A1(mai_mai_n607_), .B0(mai_mai_n62_), .Y(mai_mai_n617_));
  NOi21      m0595(.An(i_11_), .B(i_7_), .Y(mai_mai_n618_));
  AO210      m0596(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n619_));
  NO2        m0597(.A(mai_mai_n619_), .B(mai_mai_n618_), .Y(mai_mai_n620_));
  NA2        m0598(.A(mai_mai_n620_), .B(mai_mai_n205_), .Y(mai_mai_n621_));
  NA3        m0599(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n622_));
  NAi31      m0600(.An(mai_mai_n622_), .B(mai_mai_n214_), .C(i_11_), .Y(mai_mai_n623_));
  AOI210     m0601(.A0(mai_mai_n623_), .A1(mai_mai_n621_), .B0(mai_mai_n62_), .Y(mai_mai_n624_));
  NA2        m0602(.A(mai_mai_n85_), .B(mai_mai_n62_), .Y(mai_mai_n625_));
  AO210      m0603(.A0(mai_mai_n625_), .A1(mai_mai_n378_), .B0(mai_mai_n41_), .Y(mai_mai_n626_));
  NA2        m0604(.A(mai_mai_n224_), .B(mai_mai_n62_), .Y(mai_mai_n627_));
  NA2        m0605(.A(mai_mai_n409_), .B(mai_mai_n31_), .Y(mai_mai_n628_));
  OR2        m0606(.A(mai_mai_n207_), .B(mai_mai_n105_), .Y(mai_mai_n629_));
  NA2        m0607(.A(mai_mai_n629_), .B(mai_mai_n628_), .Y(mai_mai_n630_));
  NO2        m0608(.A(mai_mai_n62_), .B(i_9_), .Y(mai_mai_n631_));
  NO2        m0609(.A(mai_mai_n631_), .B(i_4_), .Y(mai_mai_n632_));
  NA2        m0610(.A(mai_mai_n632_), .B(mai_mai_n630_), .Y(mai_mai_n633_));
  NO2        m0611(.A(i_1_), .B(i_12_), .Y(mai_mai_n634_));
  NA3        m0612(.A(mai_mai_n633_), .B(mai_mai_n627_), .C(mai_mai_n626_), .Y(mai_mai_n635_));
  OAI210     m0613(.A0(mai_mai_n635_), .A1(mai_mai_n624_), .B0(i_6_), .Y(mai_mai_n636_));
  NO2        m0614(.A(mai_mai_n235_), .B(mai_mai_n83_), .Y(mai_mai_n637_));
  NO2        m0615(.A(mai_mai_n637_), .B(i_11_), .Y(mai_mai_n638_));
  INV        m0616(.A(mai_mai_n455_), .Y(mai_mai_n639_));
  NO4        m0617(.A(mai_mai_n214_), .B(mai_mai_n126_), .C(i_13_), .D(mai_mai_n83_), .Y(mai_mai_n640_));
  NA2        m0618(.A(mai_mai_n640_), .B(mai_mai_n631_), .Y(mai_mai_n641_));
  NA2        m0619(.A(mai_mai_n235_), .B(i_6_), .Y(mai_mai_n642_));
  NO3        m0620(.A(mai_mai_n610_), .B(mai_mai_n231_), .C(mai_mai_n23_), .Y(mai_mai_n643_));
  INV        m0621(.A(mai_mai_n641_), .Y(mai_mai_n644_));
  NA3        m0622(.A(mai_mai_n538_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n645_));
  NA2        m0623(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n646_));
  NA3        m0624(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n647_));
  NO2        m0625(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n648_));
  NA3        m0626(.A(mai_mai_n648_), .B(mai_mai_n261_), .C(mai_mai_n44_), .Y(mai_mai_n649_));
  OAI220     m0627(.A0(mai_mai_n649_), .A1(mai_mai_n647_), .B0(mai_mai_n646_), .B1(mai_mai_n1045_), .Y(mai_mai_n650_));
  NA3        m0628(.A(mai_mai_n631_), .B(mai_mai_n314_), .C(i_6_), .Y(mai_mai_n651_));
  NO2        m0629(.A(mai_mai_n651_), .B(mai_mai_n23_), .Y(mai_mai_n652_));
  AOI210     m0630(.A0(mai_mai_n476_), .A1(mai_mai_n418_), .B0(mai_mai_n239_), .Y(mai_mai_n653_));
  NO2        m0631(.A(mai_mai_n653_), .B(mai_mai_n601_), .Y(mai_mai_n654_));
  NAi21      m0632(.An(mai_mai_n645_), .B(mai_mai_n89_), .Y(mai_mai_n655_));
  NA2        m0633(.A(mai_mai_n648_), .B(mai_mai_n261_), .Y(mai_mai_n656_));
  NO2        m0634(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n657_), .B(mai_mai_n24_), .Y(mai_mai_n658_));
  OAI210     m0636(.A0(mai_mai_n658_), .A1(mai_mai_n656_), .B0(mai_mai_n655_), .Y(mai_mai_n659_));
  OR4        m0637(.A(mai_mai_n659_), .B(mai_mai_n654_), .C(mai_mai_n652_), .D(mai_mai_n650_), .Y(mai_mai_n660_));
  NO3        m0638(.A(mai_mai_n660_), .B(mai_mai_n644_), .C(mai_mai_n639_), .Y(mai_mai_n661_));
  NO2        m0639(.A(mai_mai_n235_), .B(mai_mai_n98_), .Y(mai_mai_n662_));
  NO2        m0640(.A(mai_mai_n662_), .B(mai_mai_n618_), .Y(mai_mai_n663_));
  NA2        m0641(.A(mai_mai_n663_), .B(i_1_), .Y(mai_mai_n664_));
  NO2        m0642(.A(mai_mai_n664_), .B(mai_mai_n612_), .Y(mai_mai_n665_));
  NA2        m0643(.A(mai_mai_n665_), .B(mai_mai_n46_), .Y(mai_mai_n666_));
  NO2        m0644(.A(mai_mai_n115_), .B(mai_mai_n37_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n83_), .B(i_9_), .Y(mai_mai_n668_));
  NO2        m0646(.A(mai_mai_n668_), .B(mai_mai_n62_), .Y(mai_mai_n669_));
  NA2        m0647(.A(i_1_), .B(i_3_), .Y(mai_mai_n670_));
  NA3        m0648(.A(mai_mai_n666_), .B(mai_mai_n661_), .C(mai_mai_n636_), .Y(mai_mai_n671_));
  NO3        m0649(.A(mai_mai_n477_), .B(i_3_), .C(i_7_), .Y(mai_mai_n672_));
  NOi21      m0650(.An(mai_mai_n672_), .B(i_10_), .Y(mai_mai_n673_));
  OA210      m0651(.A0(mai_mai_n673_), .A1(mai_mai_n243_), .B0(mai_mai_n83_), .Y(mai_mai_n674_));
  NA3        m0652(.A(mai_mai_n484_), .B(mai_mai_n520_), .C(mai_mai_n46_), .Y(mai_mai_n675_));
  NO3        m0653(.A(mai_mai_n478_), .B(mai_mai_n604_), .C(mai_mai_n83_), .Y(mai_mai_n676_));
  NA2        m0654(.A(mai_mai_n676_), .B(mai_mai_n25_), .Y(mai_mai_n677_));
  NA3        m0655(.A(mai_mai_n159_), .B(mai_mai_n82_), .C(mai_mai_n83_), .Y(mai_mai_n678_));
  NA3        m0656(.A(mai_mai_n678_), .B(mai_mai_n677_), .C(mai_mai_n675_), .Y(mai_mai_n679_));
  OAI210     m0657(.A0(mai_mai_n679_), .A1(mai_mai_n674_), .B0(i_1_), .Y(mai_mai_n680_));
  AOI210     m0658(.A0(mai_mai_n261_), .A1(mai_mai_n94_), .B0(i_1_), .Y(mai_mai_n681_));
  NO2        m0659(.A(mai_mai_n372_), .B(i_2_), .Y(mai_mai_n682_));
  NA2        m0660(.A(mai_mai_n682_), .B(mai_mai_n681_), .Y(mai_mai_n683_));
  OAI210     m0661(.A0(mai_mai_n651_), .A1(mai_mai_n446_), .B0(mai_mai_n683_), .Y(mai_mai_n684_));
  INV        m0662(.A(mai_mai_n684_), .Y(mai_mai_n685_));
  AOI210     m0663(.A0(mai_mai_n685_), .A1(mai_mai_n680_), .B0(i_13_), .Y(mai_mai_n686_));
  OR2        m0664(.A(i_11_), .B(i_7_), .Y(mai_mai_n687_));
  NA3        m0665(.A(mai_mai_n687_), .B(mai_mai_n103_), .C(mai_mai_n136_), .Y(mai_mai_n688_));
  AOI220     m0666(.A0(mai_mai_n470_), .A1(mai_mai_n159_), .B0(mai_mai_n449_), .B1(mai_mai_n136_), .Y(mai_mai_n689_));
  OAI210     m0667(.A0(mai_mai_n689_), .A1(mai_mai_n44_), .B0(mai_mai_n688_), .Y(mai_mai_n690_));
  AOI210     m0668(.A0(mai_mai_n647_), .A1(mai_mai_n54_), .B0(i_12_), .Y(mai_mai_n691_));
  NA2        m0669(.A(mai_mai_n243_), .B(mai_mai_n129_), .Y(mai_mai_n692_));
  OAI220     m0670(.A0(mai_mai_n692_), .A1(mai_mai_n41_), .B0(mai_mai_n1044_), .B1(mai_mai_n90_), .Y(mai_mai_n693_));
  AOI210     m0671(.A0(mai_mai_n690_), .A1(mai_mai_n330_), .B0(mai_mai_n693_), .Y(mai_mai_n694_));
  NA2        m0672(.A(mai_mai_n112_), .B(mai_mai_n105_), .Y(mai_mai_n695_));
  AOI220     m0673(.A0(mai_mai_n695_), .A1(mai_mai_n71_), .B0(mai_mai_n386_), .B1(mai_mai_n648_), .Y(mai_mai_n696_));
  NO2        m0674(.A(mai_mai_n696_), .B(mai_mai_n240_), .Y(mai_mai_n697_));
  AOI210     m0675(.A0(mai_mai_n446_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n698_));
  NA2        m0676(.A(mai_mai_n125_), .B(i_13_), .Y(mai_mai_n699_));
  NO2        m0677(.A(mai_mai_n647_), .B(mai_mai_n112_), .Y(mai_mai_n700_));
  INV        m0678(.A(mai_mai_n700_), .Y(mai_mai_n701_));
  OAI220     m0679(.A0(mai_mai_n701_), .A1(mai_mai_n70_), .B0(mai_mai_n699_), .B1(mai_mai_n681_), .Y(mai_mai_n702_));
  NO3        m0680(.A(mai_mai_n70_), .B(mai_mai_n32_), .C(mai_mai_n98_), .Y(mai_mai_n703_));
  NA2        m0681(.A(mai_mai_n26_), .B(mai_mai_n192_), .Y(mai_mai_n704_));
  NA2        m0682(.A(mai_mai_n704_), .B(i_7_), .Y(mai_mai_n705_));
  NO3        m0683(.A(mai_mai_n478_), .B(mai_mai_n235_), .C(mai_mai_n83_), .Y(mai_mai_n706_));
  AOI210     m0684(.A0(mai_mai_n706_), .A1(mai_mai_n705_), .B0(mai_mai_n703_), .Y(mai_mai_n707_));
  NA2        m0685(.A(mai_mai_n89_), .B(mai_mai_n99_), .Y(mai_mai_n708_));
  OAI220     m0686(.A0(mai_mai_n708_), .A1(mai_mai_n599_), .B0(mai_mai_n707_), .B1(mai_mai_n614_), .Y(mai_mai_n709_));
  NO3        m0687(.A(mai_mai_n709_), .B(mai_mai_n702_), .C(mai_mai_n697_), .Y(mai_mai_n710_));
  OR2        m0688(.A(i_11_), .B(i_6_), .Y(mai_mai_n711_));
  NA3        m0689(.A(mai_mai_n598_), .B(mai_mai_n704_), .C(i_7_), .Y(mai_mai_n712_));
  AOI210     m0690(.A0(mai_mai_n712_), .A1(mai_mai_n701_), .B0(mai_mai_n711_), .Y(mai_mai_n713_));
  NA3        m0691(.A(mai_mai_n409_), .B(mai_mai_n603_), .C(mai_mai_n94_), .Y(mai_mai_n714_));
  NA2        m0692(.A(mai_mai_n638_), .B(i_13_), .Y(mai_mai_n715_));
  NA2        m0693(.A(mai_mai_n99_), .B(mai_mai_n704_), .Y(mai_mai_n716_));
  NAi21      m0694(.An(i_11_), .B(i_12_), .Y(mai_mai_n717_));
  NOi41      m0695(.An(mai_mai_n108_), .B(mai_mai_n717_), .C(i_13_), .D(mai_mai_n83_), .Y(mai_mai_n718_));
  NO3        m0696(.A(mai_mai_n478_), .B(mai_mai_n583_), .C(mai_mai_n604_), .Y(mai_mai_n719_));
  AOI220     m0697(.A0(mai_mai_n719_), .A1(mai_mai_n308_), .B0(mai_mai_n718_), .B1(mai_mai_n716_), .Y(mai_mai_n720_));
  NA3        m0698(.A(mai_mai_n720_), .B(mai_mai_n715_), .C(mai_mai_n714_), .Y(mai_mai_n721_));
  OAI210     m0699(.A0(mai_mai_n721_), .A1(mai_mai_n713_), .B0(mai_mai_n62_), .Y(mai_mai_n722_));
  NO2        m0700(.A(i_2_), .B(i_12_), .Y(mai_mai_n723_));
  NA2        m0701(.A(mai_mai_n371_), .B(mai_mai_n723_), .Y(mai_mai_n724_));
  NA2        m0702(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n725_));
  NO3        m0703(.A(mai_mai_n725_), .B(mai_mai_n384_), .C(mai_mai_n598_), .Y(mai_mai_n726_));
  NA2        m0704(.A(mai_mai_n726_), .B(mai_mai_n371_), .Y(mai_mai_n727_));
  NO2        m0705(.A(mai_mai_n126_), .B(i_2_), .Y(mai_mai_n728_));
  NA2        m0706(.A(mai_mai_n728_), .B(mai_mai_n634_), .Y(mai_mai_n729_));
  NA3        m0707(.A(mai_mai_n729_), .B(mai_mai_n727_), .C(mai_mai_n724_), .Y(mai_mai_n730_));
  NA3        m0708(.A(mai_mai_n730_), .B(mai_mai_n45_), .C(mai_mai_n223_), .Y(mai_mai_n731_));
  NA4        m0709(.A(mai_mai_n731_), .B(mai_mai_n722_), .C(mai_mai_n710_), .D(mai_mai_n694_), .Y(mai_mai_n732_));
  OR4        m0710(.A(mai_mai_n732_), .B(mai_mai_n686_), .C(mai_mai_n671_), .D(mai_mai_n617_), .Y(mai5));
  AOI210     m0711(.A0(mai_mai_n663_), .A1(mai_mai_n264_), .B0(mai_mai_n416_), .Y(mai_mai_n734_));
  AN2        m0712(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n735_));
  NA3        m0713(.A(mai_mai_n735_), .B(mai_mai_n723_), .C(mai_mai_n105_), .Y(mai_mai_n736_));
  NO2        m0714(.A(mai_mai_n599_), .B(i_11_), .Y(mai_mai_n737_));
  OAI210     m0715(.A0(mai_mai_n603_), .A1(mai_mai_n86_), .B0(mai_mai_n737_), .Y(mai_mai_n738_));
  NA3        m0716(.A(mai_mai_n738_), .B(mai_mai_n736_), .C(mai_mai_n734_), .Y(mai_mai_n739_));
  NO3        m0717(.A(i_11_), .B(mai_mai_n235_), .C(i_13_), .Y(mai_mai_n740_));
  NO2        m0718(.A(mai_mai_n122_), .B(mai_mai_n23_), .Y(mai_mai_n741_));
  NA2        m0719(.A(i_12_), .B(i_8_), .Y(mai_mai_n742_));
  OAI210     m0720(.A0(mai_mai_n46_), .A1(i_3_), .B0(mai_mai_n742_), .Y(mai_mai_n743_));
  INV        m0721(.A(mai_mai_n445_), .Y(mai_mai_n744_));
  AOI220     m0722(.A0(mai_mai_n314_), .A1(mai_mai_n576_), .B0(mai_mai_n743_), .B1(mai_mai_n741_), .Y(mai_mai_n745_));
  INV        m0723(.A(mai_mai_n745_), .Y(mai_mai_n746_));
  NO2        m0724(.A(mai_mai_n746_), .B(mai_mai_n739_), .Y(mai_mai_n747_));
  INV        m0725(.A(mai_mai_n169_), .Y(mai_mai_n748_));
  INV        m0726(.A(mai_mai_n243_), .Y(mai_mai_n749_));
  OAI210     m0727(.A0(mai_mai_n682_), .A1(mai_mai_n447_), .B0(mai_mai_n108_), .Y(mai_mai_n750_));
  AOI210     m0728(.A0(mai_mai_n750_), .A1(mai_mai_n749_), .B0(mai_mai_n748_), .Y(mai_mai_n751_));
  NO2        m0729(.A(mai_mai_n456_), .B(mai_mai_n26_), .Y(mai_mai_n752_));
  NO2        m0730(.A(mai_mai_n752_), .B(mai_mai_n418_), .Y(mai_mai_n753_));
  NA2        m0731(.A(mai_mai_n753_), .B(i_2_), .Y(mai_mai_n754_));
  INV        m0732(.A(mai_mai_n754_), .Y(mai_mai_n755_));
  AOI210     m0733(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n415_), .Y(mai_mai_n756_));
  AOI210     m0734(.A0(mai_mai_n756_), .A1(mai_mai_n755_), .B0(mai_mai_n751_), .Y(mai_mai_n757_));
  NO2        m0735(.A(mai_mai_n189_), .B(mai_mai_n123_), .Y(mai_mai_n758_));
  OAI210     m0736(.A0(mai_mai_n758_), .A1(mai_mai_n741_), .B0(i_2_), .Y(mai_mai_n759_));
  INV        m0737(.A(mai_mai_n170_), .Y(mai_mai_n760_));
  NO3        m0738(.A(mai_mai_n619_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n761_));
  AOI210     m0739(.A0(mai_mai_n760_), .A1(mai_mai_n86_), .B0(mai_mai_n761_), .Y(mai_mai_n762_));
  AOI210     m0740(.A0(mai_mai_n762_), .A1(mai_mai_n759_), .B0(mai_mai_n192_), .Y(mai_mai_n763_));
  OA210      m0741(.A0(mai_mai_n620_), .A1(mai_mai_n124_), .B0(i_13_), .Y(mai_mai_n764_));
  NA2        m0742(.A(mai_mai_n199_), .B(mai_mai_n202_), .Y(mai_mai_n765_));
  NA2        m0743(.A(mai_mai_n149_), .B(mai_mai_n595_), .Y(mai_mai_n766_));
  AOI210     m0744(.A0(mai_mai_n766_), .A1(mai_mai_n765_), .B0(mai_mai_n374_), .Y(mai_mai_n767_));
  AOI210     m0745(.A0(mai_mai_n207_), .A1(mai_mai_n146_), .B0(mai_mai_n520_), .Y(mai_mai_n768_));
  OAI210     m0746(.A0(mai_mai_n768_), .A1(mai_mai_n224_), .B0(mai_mai_n418_), .Y(mai_mai_n769_));
  NO2        m0747(.A(mai_mai_n99_), .B(mai_mai_n44_), .Y(mai_mai_n770_));
  INV        m0748(.A(mai_mai_n297_), .Y(mai_mai_n771_));
  NA4        m0749(.A(mai_mai_n771_), .B(mai_mai_n301_), .C(mai_mai_n122_), .D(mai_mai_n42_), .Y(mai_mai_n772_));
  OAI210     m0750(.A0(mai_mai_n772_), .A1(mai_mai_n770_), .B0(mai_mai_n769_), .Y(mai_mai_n773_));
  NO4        m0751(.A(mai_mai_n773_), .B(mai_mai_n767_), .C(mai_mai_n764_), .D(mai_mai_n763_), .Y(mai_mai_n774_));
  NA2        m0752(.A(mai_mai_n576_), .B(mai_mai_n28_), .Y(mai_mai_n775_));
  NA2        m0753(.A(mai_mai_n740_), .B(mai_mai_n271_), .Y(mai_mai_n776_));
  NA2        m0754(.A(mai_mai_n776_), .B(mai_mai_n775_), .Y(mai_mai_n777_));
  NO2        m0755(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n778_));
  NO2        m0756(.A(mai_mai_n778_), .B(mai_mai_n124_), .Y(mai_mai_n779_));
  NO2        m0757(.A(mai_mai_n779_), .B(mai_mai_n595_), .Y(mai_mai_n780_));
  AOI220     m0758(.A0(mai_mai_n780_), .A1(mai_mai_n36_), .B0(mai_mai_n777_), .B1(mai_mai_n46_), .Y(mai_mai_n781_));
  NA4        m0759(.A(mai_mai_n781_), .B(mai_mai_n774_), .C(mai_mai_n757_), .D(mai_mai_n747_), .Y(mai6));
  NO3        m0760(.A(mai_mai_n252_), .B(mai_mai_n303_), .C(i_1_), .Y(mai_mai_n783_));
  NO2        m0761(.A(mai_mai_n184_), .B(mai_mai_n137_), .Y(mai_mai_n784_));
  OAI210     m0762(.A0(mai_mai_n784_), .A1(mai_mai_n783_), .B0(mai_mai_n728_), .Y(mai_mai_n785_));
  NA4        m0763(.A(mai_mai_n390_), .B(mai_mai_n483_), .C(mai_mai_n70_), .D(mai_mai_n98_), .Y(mai_mai_n786_));
  INV        m0764(.A(mai_mai_n786_), .Y(mai_mai_n787_));
  NO2        m0765(.A(i_11_), .B(i_9_), .Y(mai_mai_n788_));
  NO2        m0766(.A(mai_mai_n787_), .B(mai_mai_n326_), .Y(mai_mai_n789_));
  AO210      m0767(.A0(mai_mai_n789_), .A1(mai_mai_n785_), .B0(i_12_), .Y(mai_mai_n790_));
  NA2        m0768(.A(mai_mai_n375_), .B(mai_mai_n333_), .Y(mai_mai_n791_));
  NA2        m0769(.A(mai_mai_n583_), .B(mai_mai_n62_), .Y(mai_mai_n792_));
  NA2        m0770(.A(mai_mai_n673_), .B(mai_mai_n70_), .Y(mai_mai_n793_));
  BUFFER     m0771(.A(mai_mai_n625_), .Y(mai_mai_n794_));
  NA4        m0772(.A(mai_mai_n794_), .B(mai_mai_n793_), .C(mai_mai_n792_), .D(mai_mai_n791_), .Y(mai_mai_n795_));
  INV        m0773(.A(mai_mai_n196_), .Y(mai_mai_n796_));
  AOI220     m0774(.A0(mai_mai_n796_), .A1(mai_mai_n788_), .B0(mai_mai_n795_), .B1(mai_mai_n72_), .Y(mai_mai_n797_));
  INV        m0775(.A(mai_mai_n325_), .Y(mai_mai_n798_));
  NA2        m0776(.A(mai_mai_n74_), .B(mai_mai_n129_), .Y(mai_mai_n799_));
  INV        m0777(.A(mai_mai_n122_), .Y(mai_mai_n800_));
  NA2        m0778(.A(mai_mai_n800_), .B(mai_mai_n46_), .Y(mai_mai_n801_));
  AOI210     m0779(.A0(mai_mai_n801_), .A1(mai_mai_n799_), .B0(mai_mai_n798_), .Y(mai_mai_n802_));
  NO2        m0780(.A(mai_mai_n250_), .B(i_9_), .Y(mai_mai_n803_));
  NA2        m0781(.A(mai_mai_n803_), .B(mai_mai_n778_), .Y(mai_mai_n804_));
  AOI210     m0782(.A0(mai_mai_n804_), .A1(mai_mai_n519_), .B0(mai_mai_n184_), .Y(mai_mai_n805_));
  NO2        m0783(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n806_));
  NA3        m0784(.A(mai_mai_n806_), .B(mai_mai_n474_), .C(mai_mai_n390_), .Y(mai_mai_n807_));
  NAi32      m0785(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n808_));
  AOI210     m0786(.A0(mai_mai_n711_), .A1(mai_mai_n84_), .B0(mai_mai_n808_), .Y(mai_mai_n809_));
  OAI210     m0787(.A0(mai_mai_n672_), .A1(mai_mai_n564_), .B0(mai_mai_n563_), .Y(mai_mai_n810_));
  NAi31      m0788(.An(mai_mai_n809_), .B(mai_mai_n810_), .C(mai_mai_n807_), .Y(mai_mai_n811_));
  OR3        m0789(.A(mai_mai_n811_), .B(mai_mai_n805_), .C(mai_mai_n802_), .Y(mai_mai_n812_));
  NO2        m0790(.A(mai_mai_n687_), .B(i_2_), .Y(mai_mai_n813_));
  NA2        m0791(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n814_));
  OAI210     m0792(.A0(mai_mai_n814_), .A1(mai_mai_n408_), .B0(mai_mai_n361_), .Y(mai_mai_n815_));
  NA2        m0793(.A(mai_mai_n815_), .B(mai_mai_n813_), .Y(mai_mai_n816_));
  AO210      m0794(.A0(mai_mai_n360_), .A1(mai_mai_n350_), .B0(mai_mai_n398_), .Y(mai_mai_n817_));
  NA3        m0795(.A(mai_mai_n817_), .B(mai_mai_n253_), .C(i_7_), .Y(mai_mai_n818_));
  OR2        m0796(.A(mai_mai_n620_), .B(mai_mai_n447_), .Y(mai_mai_n819_));
  NA3        m0797(.A(mai_mai_n819_), .B(mai_mai_n145_), .C(mai_mai_n68_), .Y(mai_mai_n820_));
  AO210      m0798(.A0(mai_mai_n494_), .A1(mai_mai_n744_), .B0(mai_mai_n36_), .Y(mai_mai_n821_));
  NA4        m0799(.A(mai_mai_n821_), .B(mai_mai_n820_), .C(mai_mai_n818_), .D(mai_mai_n816_), .Y(mai_mai_n822_));
  OAI210     m0800(.A0(mai_mai_n637_), .A1(i_11_), .B0(mai_mai_n84_), .Y(mai_mai_n823_));
  NA2        m0801(.A(mai_mai_n823_), .B(mai_mai_n563_), .Y(mai_mai_n824_));
  OAI210     m0802(.A0(mai_mai_n398_), .A1(mai_mai_n203_), .B0(mai_mai_n69_), .Y(mai_mai_n825_));
  NA3        m0803(.A(mai_mai_n825_), .B(mai_mai_n824_), .C(mai_mai_n602_), .Y(mai_mai_n826_));
  AO210      m0804(.A0(mai_mai_n520_), .A1(mai_mai_n46_), .B0(mai_mai_n85_), .Y(mai_mai_n827_));
  NA3        m0805(.A(mai_mai_n827_), .B(mai_mai_n484_), .C(mai_mai_n217_), .Y(mai_mai_n828_));
  AOI210     m0806(.A0(mai_mai_n447_), .A1(mai_mai_n445_), .B0(mai_mai_n562_), .Y(mai_mai_n829_));
  NA2        m0807(.A(mai_mai_n109_), .B(mai_mai_n407_), .Y(mai_mai_n830_));
  NA2        m0808(.A(mai_mai_n242_), .B(mai_mai_n46_), .Y(mai_mai_n831_));
  NA3        m0809(.A(mai_mai_n830_), .B(mai_mai_n829_), .C(mai_mai_n828_), .Y(mai_mai_n832_));
  NO4        m0810(.A(mai_mai_n832_), .B(mai_mai_n826_), .C(mai_mai_n822_), .D(mai_mai_n812_), .Y(mai_mai_n833_));
  NA4        m0811(.A(mai_mai_n833_), .B(mai_mai_n797_), .C(mai_mai_n790_), .D(mai_mai_n380_), .Y(mai3));
  NA2        m0812(.A(i_6_), .B(i_7_), .Y(mai_mai_n835_));
  NO2        m0813(.A(mai_mai_n835_), .B(i_0_), .Y(mai_mai_n836_));
  NO2        m0814(.A(i_11_), .B(mai_mai_n235_), .Y(mai_mai_n837_));
  OAI210     m0815(.A0(mai_mai_n836_), .A1(mai_mai_n285_), .B0(mai_mai_n837_), .Y(mai_mai_n838_));
  NO2        m0816(.A(mai_mai_n838_), .B(mai_mai_n192_), .Y(mai_mai_n839_));
  NO3        m0817(.A(mai_mai_n452_), .B(mai_mai_n87_), .C(mai_mai_n44_), .Y(mai_mai_n840_));
  OA210      m0818(.A0(mai_mai_n840_), .A1(mai_mai_n839_), .B0(mai_mai_n172_), .Y(mai_mai_n841_));
  NA2        m0819(.A(mai_mai_n409_), .B(mai_mai_n45_), .Y(mai_mai_n842_));
  NO4        m0820(.A(mai_mai_n376_), .B(mai_mai_n383_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n843_));
  NA2        m0821(.A(mai_mai_n184_), .B(mai_mai_n572_), .Y(mai_mai_n844_));
  NOi31      m0822(.An(mai_mai_n844_), .B(mai_mai_n843_), .C(mai_mai_n39_), .Y(mai_mai_n845_));
  NA2        m0823(.A(mai_mai_n698_), .B(mai_mai_n668_), .Y(mai_mai_n846_));
  NA2        m0824(.A(mai_mai_n331_), .B(mai_mai_n435_), .Y(mai_mai_n847_));
  OAI220     m0825(.A0(mai_mai_n847_), .A1(mai_mai_n846_), .B0(mai_mai_n845_), .B1(mai_mai_n62_), .Y(mai_mai_n848_));
  NOi21      m0826(.An(i_5_), .B(i_9_), .Y(mai_mai_n849_));
  NA2        m0827(.A(mai_mai_n849_), .B(mai_mai_n443_), .Y(mai_mai_n850_));
  AOI210     m0828(.A0(mai_mai_n261_), .A1(mai_mai_n476_), .B0(mai_mai_n676_), .Y(mai_mai_n851_));
  NO3        m0829(.A(mai_mai_n412_), .B(mai_mai_n261_), .C(mai_mai_n72_), .Y(mai_mai_n852_));
  NO2        m0830(.A(mai_mai_n173_), .B(mai_mai_n146_), .Y(mai_mai_n853_));
  AOI210     m0831(.A0(mai_mai_n853_), .A1(mai_mai_n242_), .B0(mai_mai_n852_), .Y(mai_mai_n854_));
  OAI220     m0832(.A0(mai_mai_n854_), .A1(mai_mai_n179_), .B0(mai_mai_n851_), .B1(mai_mai_n850_), .Y(mai_mai_n855_));
  NO3        m0833(.A(mai_mai_n855_), .B(mai_mai_n848_), .C(mai_mai_n841_), .Y(mai_mai_n856_));
  NA2        m0834(.A(mai_mai_n184_), .B(mai_mai_n24_), .Y(mai_mai_n857_));
  NO2        m0835(.A(mai_mai_n667_), .B(mai_mai_n593_), .Y(mai_mai_n858_));
  NO2        m0836(.A(mai_mai_n858_), .B(mai_mai_n857_), .Y(mai_mai_n859_));
  NA2        m0837(.A(mai_mai_n308_), .B(mai_mai_n127_), .Y(mai_mai_n860_));
  NAi21      m0838(.An(mai_mai_n160_), .B(mai_mai_n435_), .Y(mai_mai_n861_));
  OAI220     m0839(.A0(mai_mai_n861_), .A1(mai_mai_n831_), .B0(mai_mai_n860_), .B1(mai_mai_n400_), .Y(mai_mai_n862_));
  NO2        m0840(.A(mai_mai_n862_), .B(mai_mai_n859_), .Y(mai_mai_n863_));
  NO2        m0841(.A(mai_mai_n390_), .B(mai_mai_n289_), .Y(mai_mai_n864_));
  NA2        m0842(.A(mai_mai_n864_), .B(mai_mai_n700_), .Y(mai_mai_n865_));
  NA2        m0843(.A(mai_mai_n573_), .B(i_0_), .Y(mai_mai_n866_));
  NO3        m0844(.A(mai_mai_n866_), .B(mai_mai_n385_), .C(mai_mai_n86_), .Y(mai_mai_n867_));
  INV        m0845(.A(mai_mai_n867_), .Y(mai_mai_n868_));
  AN2        m0846(.A(mai_mai_n93_), .B(mai_mai_n241_), .Y(mai_mai_n869_));
  NA2        m0847(.A(mai_mai_n740_), .B(mai_mai_n326_), .Y(mai_mai_n870_));
  INV        m0848(.A(mai_mai_n57_), .Y(mai_mai_n871_));
  OAI220     m0849(.A0(mai_mai_n871_), .A1(mai_mai_n870_), .B0(mai_mai_n658_), .B1(mai_mai_n540_), .Y(mai_mai_n872_));
  NA2        m0850(.A(i_0_), .B(i_10_), .Y(mai_mai_n873_));
  AOI220     m0851(.A0(mai_mai_n331_), .A1(mai_mai_n95_), .B0(mai_mai_n184_), .B1(mai_mai_n82_), .Y(mai_mai_n874_));
  NA2        m0852(.A(mai_mai_n567_), .B(i_4_), .Y(mai_mai_n875_));
  NA2        m0853(.A(mai_mai_n187_), .B(mai_mai_n202_), .Y(mai_mai_n876_));
  OAI220     m0854(.A0(mai_mai_n876_), .A1(mai_mai_n870_), .B0(mai_mai_n875_), .B1(mai_mai_n874_), .Y(mai_mai_n877_));
  NO3        m0855(.A(mai_mai_n877_), .B(mai_mai_n872_), .C(mai_mai_n869_), .Y(mai_mai_n878_));
  NA4        m0856(.A(mai_mai_n878_), .B(mai_mai_n868_), .C(mai_mai_n865_), .D(mai_mai_n863_), .Y(mai_mai_n879_));
  NA2        m0857(.A(i_11_), .B(i_9_), .Y(mai_mai_n880_));
  NO2        m0858(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n881_));
  NA2        m0859(.A(mai_mai_n395_), .B(mai_mai_n177_), .Y(mai_mai_n882_));
  NA2        m0860(.A(mai_mai_n882_), .B(mai_mai_n158_), .Y(mai_mai_n883_));
  NO2        m0861(.A(mai_mai_n880_), .B(mai_mai_n72_), .Y(mai_mai_n884_));
  NO2        m0862(.A(mai_mai_n173_), .B(i_0_), .Y(mai_mai_n885_));
  INV        m0863(.A(mai_mai_n885_), .Y(mai_mai_n886_));
  NA2        m0864(.A(mai_mai_n474_), .B(mai_mai_n229_), .Y(mai_mai_n887_));
  NA2        m0865(.A(mai_mai_n373_), .B(i_4_), .Y(mai_mai_n888_));
  OAI220     m0866(.A0(mai_mai_n888_), .A1(mai_mai_n850_), .B0(mai_mai_n887_), .B1(mai_mai_n886_), .Y(mai_mai_n889_));
  NO2        m0867(.A(mai_mai_n889_), .B(mai_mai_n883_), .Y(mai_mai_n890_));
  NA2        m0868(.A(mai_mai_n657_), .B(mai_mai_n119_), .Y(mai_mai_n891_));
  NO2        m0869(.A(i_6_), .B(mai_mai_n891_), .Y(mai_mai_n892_));
  AOI210     m0870(.A0(mai_mai_n446_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n893_));
  NA2        m0871(.A(mai_mai_n169_), .B(mai_mai_n100_), .Y(mai_mai_n894_));
  NOi32      m0872(.An(mai_mai_n893_), .Bn(mai_mai_n187_), .C(mai_mai_n894_), .Y(mai_mai_n895_));
  AOI210     m0873(.A0(mai_mai_n603_), .A1(mai_mai_n326_), .B0(mai_mai_n241_), .Y(mai_mai_n896_));
  NO2        m0874(.A(mai_mai_n896_), .B(mai_mai_n842_), .Y(mai_mai_n897_));
  NO3        m0875(.A(mai_mai_n897_), .B(mai_mai_n895_), .C(mai_mai_n892_), .Y(mai_mai_n898_));
  NOi21      m0876(.An(i_7_), .B(i_5_), .Y(mai_mai_n899_));
  NOi31      m0877(.An(mai_mai_n899_), .B(i_0_), .C(mai_mai_n717_), .Y(mai_mai_n900_));
  NA3        m0878(.A(mai_mai_n900_), .B(mai_mai_n384_), .C(i_6_), .Y(mai_mai_n901_));
  OA210      m0879(.A0(mai_mai_n894_), .A1(mai_mai_n519_), .B0(mai_mai_n901_), .Y(mai_mai_n902_));
  NO3        m0880(.A(mai_mai_n403_), .B(mai_mai_n363_), .C(mai_mai_n359_), .Y(mai_mai_n903_));
  NO2        m0881(.A(mai_mai_n255_), .B(mai_mai_n315_), .Y(mai_mai_n904_));
  INV        m0882(.A(mai_mai_n717_), .Y(mai_mai_n905_));
  AOI210     m0883(.A0(mai_mai_n905_), .A1(mai_mai_n904_), .B0(mai_mai_n903_), .Y(mai_mai_n906_));
  NA4        m0884(.A(mai_mai_n906_), .B(mai_mai_n902_), .C(mai_mai_n898_), .D(mai_mai_n890_), .Y(mai_mai_n907_));
  NO2        m0885(.A(mai_mai_n857_), .B(mai_mai_n237_), .Y(mai_mai_n908_));
  AN2        m0886(.A(mai_mai_n330_), .B(mai_mai_n326_), .Y(mai_mai_n909_));
  AO220      m0887(.A0(mai_mai_n909_), .A1(mai_mai_n853_), .B0(mai_mai_n345_), .B1(mai_mai_n27_), .Y(mai_mai_n910_));
  OAI210     m0888(.A0(mai_mai_n910_), .A1(mai_mai_n908_), .B0(i_10_), .Y(mai_mai_n911_));
  OA210      m0889(.A0(mai_mai_n474_), .A1(mai_mai_n221_), .B0(mai_mai_n473_), .Y(mai_mai_n912_));
  NA3        m0890(.A(mai_mai_n473_), .B(mai_mai_n409_), .C(mai_mai_n45_), .Y(mai_mai_n913_));
  OAI210     m0891(.A0(mai_mai_n861_), .A1(i_6_), .B0(mai_mai_n913_), .Y(mai_mai_n914_));
  NA2        m0892(.A(mai_mai_n884_), .B(mai_mai_n301_), .Y(mai_mai_n915_));
  NA2        m0893(.A(mai_mai_n186_), .B(mai_mai_n915_), .Y(mai_mai_n916_));
  AOI220     m0894(.A0(mai_mai_n916_), .A1(mai_mai_n474_), .B0(mai_mai_n914_), .B1(mai_mai_n72_), .Y(mai_mai_n917_));
  NA3        m0895(.A(mai_mai_n814_), .B(mai_mai_n382_), .C(mai_mai_n637_), .Y(mai_mai_n918_));
  NA2        m0896(.A(mai_mai_n90_), .B(mai_mai_n44_), .Y(mai_mai_n919_));
  NO2        m0897(.A(mai_mai_n74_), .B(mai_mai_n742_), .Y(mai_mai_n920_));
  AOI220     m0898(.A0(mai_mai_n920_), .A1(mai_mai_n919_), .B0(mai_mai_n172_), .B1(mai_mai_n593_), .Y(mai_mai_n921_));
  AOI210     m0899(.A0(mai_mai_n921_), .A1(mai_mai_n918_), .B0(mai_mai_n47_), .Y(mai_mai_n922_));
  NO3        m0900(.A(i_5_), .B(mai_mai_n358_), .C(mai_mai_n24_), .Y(mai_mai_n923_));
  INV        m0901(.A(mai_mai_n923_), .Y(mai_mai_n924_));
  NAi21      m0902(.An(i_9_), .B(i_5_), .Y(mai_mai_n925_));
  NO2        m0903(.A(mai_mai_n597_), .B(mai_mai_n102_), .Y(mai_mai_n926_));
  NA2        m0904(.A(mai_mai_n926_), .B(i_0_), .Y(mai_mai_n927_));
  OAI220     m0905(.A0(mai_mai_n927_), .A1(mai_mai_n83_), .B0(mai_mai_n924_), .B1(mai_mai_n170_), .Y(mai_mai_n928_));
  NO2        m0906(.A(mai_mai_n928_), .B(mai_mai_n922_), .Y(mai_mai_n929_));
  NA3        m0907(.A(mai_mai_n929_), .B(mai_mai_n917_), .C(mai_mai_n911_), .Y(mai_mai_n930_));
  NO3        m0908(.A(mai_mai_n930_), .B(mai_mai_n907_), .C(mai_mai_n879_), .Y(mai_mai_n931_));
  NO2        m0909(.A(i_0_), .B(mai_mai_n717_), .Y(mai_mai_n932_));
  NA2        m0910(.A(mai_mai_n72_), .B(mai_mai_n44_), .Y(mai_mai_n933_));
  NA2        m0911(.A(mai_mai_n873_), .B(mai_mai_n933_), .Y(mai_mai_n934_));
  NO3        m0912(.A(mai_mai_n102_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n935_));
  AO220      m0913(.A0(mai_mai_n935_), .A1(mai_mai_n934_), .B0(mai_mai_n932_), .B1(mai_mai_n172_), .Y(mai_mai_n936_));
  NO2        m0914(.A(mai_mai_n792_), .B(mai_mai_n894_), .Y(mai_mai_n937_));
  AOI210     m0915(.A0(mai_mai_n936_), .A1(mai_mai_n347_), .B0(mai_mai_n937_), .Y(mai_mai_n938_));
  NA2        m0916(.A(mai_mai_n728_), .B(mai_mai_n144_), .Y(mai_mai_n939_));
  INV        m0917(.A(mai_mai_n939_), .Y(mai_mai_n940_));
  NA3        m0918(.A(mai_mai_n940_), .B(mai_mai_n668_), .C(mai_mai_n72_), .Y(mai_mai_n941_));
  NO2        m0919(.A(mai_mai_n810_), .B(mai_mai_n403_), .Y(mai_mai_n942_));
  NA3        m0920(.A(mai_mai_n836_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n943_));
  NA2        m0921(.A(mai_mai_n837_), .B(i_9_), .Y(mai_mai_n944_));
  AOI210     m0922(.A0(mai_mai_n943_), .A1(mai_mai_n500_), .B0(mai_mai_n944_), .Y(mai_mai_n945_));
  OAI210     m0923(.A0(mai_mai_n242_), .A1(i_9_), .B0(mai_mai_n228_), .Y(mai_mai_n946_));
  AOI210     m0924(.A0(mai_mai_n946_), .A1(mai_mai_n866_), .B0(mai_mai_n151_), .Y(mai_mai_n947_));
  NO3        m0925(.A(mai_mai_n947_), .B(mai_mai_n945_), .C(mai_mai_n942_), .Y(mai_mai_n948_));
  NA3        m0926(.A(mai_mai_n948_), .B(mai_mai_n941_), .C(mai_mai_n938_), .Y(mai_mai_n949_));
  NA2        m0927(.A(mai_mai_n909_), .B(mai_mai_n374_), .Y(mai_mai_n950_));
  AOI210     m0928(.A0(mai_mai_n296_), .A1(mai_mai_n160_), .B0(mai_mai_n950_), .Y(mai_mai_n951_));
  NA3        m0929(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n952_));
  NA2        m0930(.A(mai_mai_n881_), .B(mai_mai_n488_), .Y(mai_mai_n953_));
  AOI210     m0931(.A0(mai_mai_n952_), .A1(mai_mai_n160_), .B0(mai_mai_n953_), .Y(mai_mai_n954_));
  NO2        m0932(.A(mai_mai_n954_), .B(mai_mai_n951_), .Y(mai_mai_n955_));
  NO3        m0933(.A(mai_mai_n873_), .B(mai_mai_n849_), .C(mai_mai_n189_), .Y(mai_mai_n956_));
  AOI220     m0934(.A0(mai_mai_n956_), .A1(i_11_), .B0(mai_mai_n568_), .B1(mai_mai_n74_), .Y(mai_mai_n957_));
  NO3        m0935(.A(mai_mai_n208_), .B(mai_mai_n383_), .C(i_0_), .Y(mai_mai_n958_));
  OAI210     m0936(.A0(mai_mai_n958_), .A1(mai_mai_n75_), .B0(i_13_), .Y(mai_mai_n959_));
  INV        m0937(.A(mai_mai_n217_), .Y(mai_mai_n960_));
  OAI220     m0938(.A0(mai_mai_n533_), .A1(mai_mai_n137_), .B0(mai_mai_n642_), .B1(mai_mai_n614_), .Y(mai_mai_n961_));
  NA3        m0939(.A(mai_mai_n961_), .B(i_7_), .C(mai_mai_n960_), .Y(mai_mai_n962_));
  NA4        m0940(.A(mai_mai_n962_), .B(mai_mai_n959_), .C(mai_mai_n957_), .D(mai_mai_n955_), .Y(mai_mai_n963_));
  NO2        m0941(.A(mai_mai_n240_), .B(mai_mai_n90_), .Y(mai_mai_n964_));
  AOI210     m0942(.A0(mai_mai_n964_), .A1(mai_mai_n932_), .B0(mai_mai_n106_), .Y(mai_mai_n965_));
  AOI220     m0943(.A0(mai_mai_n899_), .A1(mai_mai_n488_), .B0(mai_mai_n836_), .B1(mai_mai_n161_), .Y(mai_mai_n966_));
  NA2        m0944(.A(mai_mai_n350_), .B(mai_mai_n174_), .Y(mai_mai_n967_));
  OA220      m0945(.A0(mai_mai_n967_), .A1(mai_mai_n966_), .B0(mai_mai_n965_), .B1(i_5_), .Y(mai_mai_n968_));
  AOI210     m0946(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n173_), .Y(mai_mai_n969_));
  NA2        m0947(.A(mai_mai_n969_), .B(mai_mai_n912_), .Y(mai_mai_n970_));
  NA3        m0948(.A(mai_mai_n611_), .B(mai_mai_n184_), .C(mai_mai_n82_), .Y(mai_mai_n971_));
  NA2        m0949(.A(mai_mai_n971_), .B(mai_mai_n549_), .Y(mai_mai_n972_));
  NO3        m0950(.A(mai_mai_n842_), .B(mai_mai_n54_), .C(mai_mai_n48_), .Y(mai_mai_n973_));
  NA2        m0951(.A(mai_mai_n493_), .B(mai_mai_n471_), .Y(mai_mai_n974_));
  NO3        m0952(.A(mai_mai_n974_), .B(mai_mai_n973_), .C(mai_mai_n972_), .Y(mai_mai_n975_));
  NA3        m0953(.A(mai_mai_n390_), .B(mai_mai_n169_), .C(mai_mai_n168_), .Y(mai_mai_n976_));
  NA3        m0954(.A(mai_mai_n881_), .B(mai_mai_n285_), .C(mai_mai_n228_), .Y(mai_mai_n977_));
  NA2        m0955(.A(mai_mai_n977_), .B(mai_mai_n976_), .Y(mai_mai_n978_));
  NA3        m0956(.A(mai_mai_n390_), .B(mai_mai_n332_), .C(mai_mai_n220_), .Y(mai_mai_n979_));
  OAI210     m0957(.A0(mai_mai_n844_), .A1(mai_mai_n645_), .B0(mai_mai_n979_), .Y(mai_mai_n980_));
  NOi31      m0958(.An(mai_mai_n389_), .B(mai_mai_n933_), .C(mai_mai_n237_), .Y(mai_mai_n981_));
  NO3        m0959(.A(mai_mai_n880_), .B(mai_mai_n217_), .C(mai_mai_n189_), .Y(mai_mai_n982_));
  NO4        m0960(.A(mai_mai_n982_), .B(mai_mai_n981_), .C(mai_mai_n980_), .D(mai_mai_n978_), .Y(mai_mai_n983_));
  NA4        m0961(.A(mai_mai_n983_), .B(mai_mai_n975_), .C(mai_mai_n970_), .D(mai_mai_n968_), .Y(mai_mai_n984_));
  INV        m0962(.A(mai_mai_n613_), .Y(mai_mai_n985_));
  NO3        m0963(.A(mai_mai_n985_), .B(mai_mai_n560_), .C(mai_mai_n344_), .Y(mai_mai_n986_));
  INV        m0964(.A(mai_mai_n986_), .Y(mai_mai_n987_));
  NA3        m0965(.A(mai_mai_n301_), .B(i_5_), .C(mai_mai_n192_), .Y(mai_mai_n988_));
  NA2        m0966(.A(mai_mai_n988_), .B(mai_mai_n240_), .Y(mai_mai_n989_));
  NO4        m0967(.A(mai_mai_n237_), .B(mai_mai_n208_), .C(i_0_), .D(i_12_), .Y(mai_mai_n990_));
  AOI220     m0968(.A0(mai_mai_n990_), .A1(mai_mai_n989_), .B0(mai_mai_n787_), .B1(mai_mai_n174_), .Y(mai_mai_n991_));
  AN2        m0969(.A(mai_mai_n873_), .B(mai_mai_n151_), .Y(mai_mai_n992_));
  NO4        m0970(.A(mai_mai_n992_), .B(i_12_), .C(mai_mai_n645_), .D(mai_mai_n129_), .Y(mai_mai_n993_));
  NA2        m0971(.A(mai_mai_n993_), .B(mai_mai_n217_), .Y(mai_mai_n994_));
  NA3        m0972(.A(mai_mai_n95_), .B(mai_mai_n572_), .C(i_11_), .Y(mai_mai_n995_));
  NO2        m0973(.A(mai_mai_n995_), .B(mai_mai_n153_), .Y(mai_mai_n996_));
  NA2        m0974(.A(mai_mai_n899_), .B(mai_mai_n470_), .Y(mai_mai_n997_));
  OAI220     m0975(.A0(i_7_), .A1(mai_mai_n988_), .B0(mai_mai_n997_), .B1(mai_mai_n669_), .Y(mai_mai_n998_));
  AOI210     m0976(.A0(mai_mai_n998_), .A1(mai_mai_n885_), .B0(mai_mai_n996_), .Y(mai_mai_n999_));
  NA4        m0977(.A(mai_mai_n999_), .B(mai_mai_n994_), .C(mai_mai_n991_), .D(mai_mai_n987_), .Y(mai_mai_n1000_));
  NO4        m0978(.A(mai_mai_n1000_), .B(mai_mai_n984_), .C(mai_mai_n963_), .D(mai_mai_n949_), .Y(mai_mai_n1001_));
  OAI210     m0979(.A0(mai_mai_n813_), .A1(mai_mai_n806_), .B0(mai_mai_n37_), .Y(mai_mai_n1002_));
  NA3        m0980(.A(mai_mai_n893_), .B(mai_mai_n371_), .C(i_5_), .Y(mai_mai_n1003_));
  NA3        m0981(.A(mai_mai_n1003_), .B(mai_mai_n1002_), .C(mai_mai_n609_), .Y(mai_mai_n1004_));
  NA2        m0982(.A(mai_mai_n1004_), .B(mai_mai_n205_), .Y(mai_mai_n1005_));
  NA2        m0983(.A(mai_mai_n185_), .B(mai_mai_n187_), .Y(mai_mai_n1006_));
  AO210      m0984(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n1006_), .Y(mai_mai_n1007_));
  OAI210     m0985(.A0(mai_mai_n613_), .A1(mai_mai_n611_), .B0(mai_mai_n314_), .Y(mai_mai_n1008_));
  INV        m0986(.A(mai_mai_n643_), .Y(mai_mai_n1009_));
  NA3        m0987(.A(mai_mai_n1009_), .B(mai_mai_n1008_), .C(mai_mai_n1007_), .Y(mai_mai_n1010_));
  NO2        m0988(.A(mai_mai_n461_), .B(mai_mai_n261_), .Y(mai_mai_n1011_));
  NO4        m0989(.A(mai_mai_n231_), .B(mai_mai_n143_), .C(mai_mai_n670_), .D(mai_mai_n37_), .Y(mai_mai_n1012_));
  NO2        m0990(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .Y(mai_mai_n1013_));
  OAI210     m0991(.A0(mai_mai_n995_), .A1(mai_mai_n146_), .B0(mai_mai_n1013_), .Y(mai_mai_n1014_));
  AOI210     m0992(.A0(mai_mai_n1010_), .A1(mai_mai_n48_), .B0(mai_mai_n1014_), .Y(mai_mai_n1015_));
  AOI210     m0993(.A0(mai_mai_n1015_), .A1(mai_mai_n1005_), .B0(mai_mai_n72_), .Y(mai_mai_n1016_));
  NO2        m0994(.A(mai_mai_n565_), .B(mai_mai_n379_), .Y(mai_mai_n1017_));
  NO2        m0995(.A(mai_mai_n1017_), .B(mai_mai_n748_), .Y(mai_mai_n1018_));
  INV        m0996(.A(mai_mai_n75_), .Y(mai_mai_n1019_));
  AOI210     m0997(.A0(mai_mai_n969_), .A1(mai_mai_n881_), .B0(mai_mai_n900_), .Y(mai_mai_n1020_));
  AOI210     m0998(.A0(mai_mai_n1020_), .A1(mai_mai_n1019_), .B0(mai_mai_n670_), .Y(mai_mai_n1021_));
  NA2        m0999(.A(mai_mai_n255_), .B(mai_mai_n56_), .Y(mai_mai_n1022_));
  AOI220     m1000(.A0(mai_mai_n1022_), .A1(mai_mai_n75_), .B0(mai_mai_n345_), .B1(mai_mai_n252_), .Y(mai_mai_n1023_));
  NO2        m1001(.A(mai_mai_n1023_), .B(mai_mai_n235_), .Y(mai_mai_n1024_));
  NA3        m1002(.A(mai_mai_n93_), .B(mai_mai_n303_), .C(mai_mai_n31_), .Y(mai_mai_n1025_));
  INV        m1003(.A(mai_mai_n1025_), .Y(mai_mai_n1026_));
  NO3        m1004(.A(mai_mai_n1026_), .B(mai_mai_n1024_), .C(mai_mai_n1021_), .Y(mai_mai_n1027_));
  OAI210     m1005(.A0(mai_mai_n263_), .A1(mai_mai_n156_), .B0(mai_mai_n86_), .Y(mai_mai_n1028_));
  NA3        m1006(.A(mai_mai_n752_), .B(mai_mai_n285_), .C(mai_mai_n79_), .Y(mai_mai_n1029_));
  AOI210     m1007(.A0(mai_mai_n1029_), .A1(mai_mai_n1028_), .B0(i_11_), .Y(mai_mai_n1030_));
  OAI210     m1008(.A0(mai_mai_n1048_), .A1(mai_mai_n893_), .B0(mai_mai_n205_), .Y(mai_mai_n1031_));
  NA2        m1009(.A(mai_mai_n162_), .B(i_5_), .Y(mai_mai_n1032_));
  AOI210     m1010(.A0(mai_mai_n1031_), .A1(mai_mai_n765_), .B0(mai_mai_n1032_), .Y(mai_mai_n1033_));
  NO4        m1011(.A(mai_mai_n925_), .B(mai_mai_n477_), .C(mai_mai_n251_), .D(mai_mai_n250_), .Y(mai_mai_n1034_));
  NO2        m1012(.A(mai_mai_n1034_), .B(mai_mai_n562_), .Y(mai_mai_n1035_));
  NO2        m1013(.A(mai_mai_n809_), .B(mai_mai_n364_), .Y(mai_mai_n1036_));
  AOI210     m1014(.A0(mai_mai_n1036_), .A1(mai_mai_n1035_), .B0(mai_mai_n41_), .Y(mai_mai_n1037_));
  NO3        m1015(.A(mai_mai_n1037_), .B(mai_mai_n1033_), .C(mai_mai_n1030_), .Y(mai_mai_n1038_));
  OAI210     m1016(.A0(mai_mai_n1027_), .A1(i_4_), .B0(mai_mai_n1038_), .Y(mai_mai_n1039_));
  NO3        m1017(.A(mai_mai_n1039_), .B(mai_mai_n1018_), .C(mai_mai_n1016_), .Y(mai_mai_n1040_));
  NA4        m1018(.A(mai_mai_n1040_), .B(mai_mai_n1001_), .C(mai_mai_n931_), .D(mai_mai_n856_), .Y(mai4));
  INV        m1019(.A(mai_mai_n691_), .Y(mai_mai_n1044_));
  INV        m1020(.A(i_2_), .Y(mai_mai_n1045_));
  INV        m1021(.A(i_1_), .Y(mai_mai_n1046_));
  INV        m1022(.A(i_12_), .Y(mai_mai_n1047_));
  INV        m1023(.A(i_12_), .Y(mai_mai_n1048_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  NA2        u0028(.A(i_0_), .B(i_2_), .Y(men_men_n51_));
  NA2        u0029(.A(i_7_), .B(i_9_), .Y(men_men_n52_));
  NO2        u0030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NA3        u0031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n54_));
  NO2        u0032(.A(i_1_), .B(i_6_), .Y(men_men_n55_));
  NA2        u0033(.A(i_8_), .B(i_7_), .Y(men_men_n56_));
  INV        u0034(.A(men_men_n54_), .Y(men_men_n57_));
  NA2        u0035(.A(men_men_n57_), .B(i_12_), .Y(men_men_n58_));
  NAi21      u0036(.An(i_2_), .B(i_7_), .Y(men_men_n59_));
  INV        u0037(.A(i_1_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_6_), .Y(men_men_n61_));
  NA3        u0039(.A(men_men_n61_), .B(men_men_n59_), .C(men_men_n31_), .Y(men_men_n62_));
  NA2        u0040(.A(men_men_n62_), .B(men_men_n58_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n50_), .B(i_2_), .Y(men_men_n64_));
  AOI210     u0042(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_6_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(men_men_n25_), .Y(men_men_n67_));
  INV        u0045(.A(i_0_), .Y(men_men_n68_));
  NAi21      u0046(.An(i_5_), .B(i_10_), .Y(men_men_n69_));
  NA2        u0047(.A(i_5_), .B(i_9_), .Y(men_men_n70_));
  AOI210     u0048(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n68_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n67_), .Y(men_men_n72_));
  OAI210     u0050(.A0(men_men_n65_), .A1(men_men_n64_), .B0(men_men_n72_), .Y(men_men_n73_));
  OAI210     u0051(.A0(men_men_n73_), .A1(men_men_n63_), .B0(i_0_), .Y(men_men_n74_));
  NA2        u0052(.A(i_12_), .B(i_5_), .Y(men_men_n75_));
  NA2        u0053(.A(i_2_), .B(i_8_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n55_), .Y(men_men_n77_));
  NO2        u0055(.A(i_3_), .B(i_9_), .Y(men_men_n78_));
  NO2        u0056(.A(i_3_), .B(i_7_), .Y(men_men_n79_));
  NO3        u0057(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n60_), .Y(men_men_n80_));
  INV        u0058(.A(i_6_), .Y(men_men_n81_));
  OR4        u0059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n82_));
  INV        u0060(.A(men_men_n82_), .Y(men_men_n83_));
  NO2        u0061(.A(i_2_), .B(i_7_), .Y(men_men_n84_));
  AOI210     u0062(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n84_), .Y(men_men_n85_));
  OAI210     u0063(.A0(men_men_n80_), .A1(men_men_n77_), .B0(men_men_n85_), .Y(men_men_n86_));
  NAi21      u0064(.An(i_6_), .B(i_10_), .Y(men_men_n87_));
  NA2        u0065(.A(i_6_), .B(i_9_), .Y(men_men_n88_));
  AOI210     u0066(.A0(men_men_n88_), .A1(men_men_n87_), .B0(men_men_n60_), .Y(men_men_n89_));
  NA2        u0067(.A(i_2_), .B(i_6_), .Y(men_men_n90_));
  NO3        u0068(.A(men_men_n90_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n91_));
  NO2        u0069(.A(men_men_n91_), .B(men_men_n89_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n92_), .A1(men_men_n86_), .B0(men_men_n75_), .Y(men_men_n93_));
  AN3        u0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n94_));
  NAi21      u0072(.An(i_6_), .B(i_11_), .Y(men_men_n95_));
  NO2        u0073(.A(i_5_), .B(i_8_), .Y(men_men_n96_));
  NOi21      u0074(.An(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  AOI220     u0075(.A0(men_men_n97_), .A1(men_men_n59_), .B0(men_men_n94_), .B1(men_men_n32_), .Y(men_men_n98_));
  INV        u0076(.A(i_7_), .Y(men_men_n99_));
  NA2        u0077(.A(men_men_n46_), .B(men_men_n99_), .Y(men_men_n100_));
  NO2        u0078(.A(i_0_), .B(i_5_), .Y(men_men_n101_));
  NO2        u0079(.A(men_men_n101_), .B(men_men_n81_), .Y(men_men_n102_));
  NA2        u0080(.A(i_12_), .B(i_3_), .Y(men_men_n103_));
  INV        u0081(.A(men_men_n103_), .Y(men_men_n104_));
  NA3        u0082(.A(men_men_n104_), .B(men_men_n102_), .C(men_men_n100_), .Y(men_men_n105_));
  NAi21      u0083(.An(i_7_), .B(i_11_), .Y(men_men_n106_));
  NO3        u0084(.A(men_men_n106_), .B(men_men_n87_), .C(men_men_n51_), .Y(men_men_n107_));
  AN2        u0085(.A(i_2_), .B(i_10_), .Y(men_men_n108_));
  NO2        u0086(.A(men_men_n108_), .B(i_7_), .Y(men_men_n109_));
  OR2        u0087(.A(men_men_n75_), .B(men_men_n55_), .Y(men_men_n110_));
  NO2        u0088(.A(i_8_), .B(men_men_n99_), .Y(men_men_n111_));
  NO3        u0089(.A(men_men_n111_), .B(men_men_n110_), .C(men_men_n109_), .Y(men_men_n112_));
  NA2        u0090(.A(i_12_), .B(i_7_), .Y(men_men_n113_));
  NO2        u0091(.A(men_men_n60_), .B(men_men_n26_), .Y(men_men_n114_));
  NA2        u0092(.A(men_men_n114_), .B(i_0_), .Y(men_men_n115_));
  NA2        u0093(.A(i_11_), .B(i_12_), .Y(men_men_n116_));
  OAI210     u0094(.A0(men_men_n115_), .A1(men_men_n113_), .B0(men_men_n116_), .Y(men_men_n117_));
  NO2        u0095(.A(men_men_n117_), .B(men_men_n112_), .Y(men_men_n118_));
  NAi41      u0096(.An(men_men_n107_), .B(men_men_n118_), .C(men_men_n105_), .D(men_men_n98_), .Y(men_men_n119_));
  NOi21      u0097(.An(i_1_), .B(i_5_), .Y(men_men_n120_));
  NA2        u0098(.A(men_men_n120_), .B(i_11_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n99_), .B(men_men_n37_), .Y(men_men_n122_));
  NA2        u0100(.A(i_7_), .B(men_men_n25_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n123_), .B(men_men_n122_), .Y(men_men_n124_));
  NO2        u0102(.A(men_men_n124_), .B(men_men_n46_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n88_), .B(men_men_n87_), .Y(men_men_n126_));
  NAi21      u0104(.An(i_3_), .B(i_8_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n127_), .B(men_men_n59_), .Y(men_men_n128_));
  NOi21      u0106(.An(men_men_n128_), .B(men_men_n126_), .Y(men_men_n129_));
  NO2        u0107(.A(i_1_), .B(men_men_n81_), .Y(men_men_n130_));
  NO2        u0108(.A(i_6_), .B(i_5_), .Y(men_men_n131_));
  NA2        u0109(.A(men_men_n131_), .B(i_3_), .Y(men_men_n132_));
  AO210      u0110(.A0(men_men_n132_), .A1(men_men_n47_), .B0(men_men_n130_), .Y(men_men_n133_));
  OAI220     u0111(.A0(men_men_n133_), .A1(men_men_n106_), .B0(men_men_n129_), .B1(men_men_n121_), .Y(men_men_n134_));
  NO3        u0112(.A(men_men_n134_), .B(men_men_n119_), .C(men_men_n93_), .Y(men_men_n135_));
  NA2        u0113(.A(men_men_n135_), .B(men_men_n74_), .Y(men2));
  NO2        u0114(.A(men_men_n60_), .B(men_men_n37_), .Y(men_men_n137_));
  NA2        u0115(.A(i_6_), .B(men_men_n25_), .Y(men_men_n138_));
  NA2        u0116(.A(men_men_n138_), .B(men_men_n137_), .Y(men_men_n139_));
  NA4        u0117(.A(men_men_n139_), .B(men_men_n72_), .C(men_men_n64_), .D(men_men_n30_), .Y(men0));
  AN2        u0118(.A(i_8_), .B(i_7_), .Y(men_men_n141_));
  NA2        u0119(.A(men_men_n141_), .B(i_6_), .Y(men_men_n142_));
  NO2        u0120(.A(i_12_), .B(i_13_), .Y(men_men_n143_));
  NAi21      u0121(.An(i_5_), .B(i_11_), .Y(men_men_n144_));
  NOi21      u0122(.An(men_men_n143_), .B(men_men_n144_), .Y(men_men_n145_));
  NO2        u0123(.A(i_0_), .B(i_1_), .Y(men_men_n146_));
  NA2        u0124(.A(i_2_), .B(i_3_), .Y(men_men_n147_));
  NO2        u0125(.A(men_men_n147_), .B(i_4_), .Y(men_men_n148_));
  NA3        u0126(.A(men_men_n148_), .B(men_men_n146_), .C(men_men_n145_), .Y(men_men_n149_));
  OR2        u0127(.A(men_men_n149_), .B(men_men_n25_), .Y(men_men_n150_));
  AN2        u0128(.A(men_men_n143_), .B(men_men_n78_), .Y(men_men_n151_));
  NO2        u0129(.A(men_men_n151_), .B(men_men_n27_), .Y(men_men_n152_));
  NA2        u0130(.A(i_1_), .B(i_5_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n68_), .B(men_men_n46_), .Y(men_men_n154_));
  NA2        u0132(.A(men_men_n154_), .B(men_men_n36_), .Y(men_men_n155_));
  NO3        u0133(.A(men_men_n155_), .B(men_men_n153_), .C(men_men_n152_), .Y(men_men_n156_));
  OR2        u0134(.A(i_0_), .B(i_1_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n75_), .C(i_13_), .Y(men_men_n158_));
  NAi32      u0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n159_));
  NAi21      u0137(.An(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  NOi21      u0138(.An(i_4_), .B(i_10_), .Y(men_men_n161_));
  NA2        u0139(.A(men_men_n161_), .B(men_men_n39_), .Y(men_men_n162_));
  NO2        u0140(.A(i_3_), .B(i_5_), .Y(men_men_n163_));
  NO3        u0141(.A(men_men_n68_), .B(i_2_), .C(i_1_), .Y(men_men_n164_));
  NA2        u0142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OAI210     u0143(.A0(men_men_n165_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n166_));
  NO2        u0144(.A(men_men_n166_), .B(men_men_n156_), .Y(men_men_n167_));
  AOI210     u0145(.A0(men_men_n167_), .A1(men_men_n150_), .B0(men_men_n142_), .Y(men_men_n168_));
  NA3        u0146(.A(men_men_n68_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n169_));
  NOi21      u0147(.An(i_4_), .B(i_9_), .Y(men_men_n170_));
  NOi21      u0148(.An(i_11_), .B(i_13_), .Y(men_men_n171_));
  NA2        u0149(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  NO2        u0150(.A(i_4_), .B(i_5_), .Y(men_men_n173_));
  NAi21      u0151(.An(i_12_), .B(i_11_), .Y(men_men_n174_));
  NO2        u0152(.A(men_men_n174_), .B(i_13_), .Y(men_men_n175_));
  NA3        u0153(.A(men_men_n175_), .B(men_men_n173_), .C(men_men_n78_), .Y(men_men_n176_));
  AOI210     u0154(.A0(men_men_n176_), .A1(men_men_n172_), .B0(men_men_n169_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n68_), .B(men_men_n60_), .Y(men_men_n178_));
  NA2        u0156(.A(men_men_n178_), .B(men_men_n46_), .Y(men_men_n179_));
  NA2        u0157(.A(men_men_n36_), .B(i_5_), .Y(men_men_n180_));
  NAi31      u0158(.An(men_men_n180_), .B(men_men_n151_), .C(i_11_), .Y(men_men_n181_));
  NA2        u0159(.A(i_3_), .B(i_5_), .Y(men_men_n182_));
  OR2        u0160(.A(men_men_n182_), .B(men_men_n172_), .Y(men_men_n183_));
  AOI210     u0161(.A0(men_men_n183_), .A1(men_men_n181_), .B0(men_men_n179_), .Y(men_men_n184_));
  NO2        u0162(.A(men_men_n68_), .B(i_5_), .Y(men_men_n185_));
  NO2        u0163(.A(i_13_), .B(i_10_), .Y(men_men_n186_));
  NA3        u0164(.A(men_men_n186_), .B(men_men_n185_), .C(men_men_n44_), .Y(men_men_n187_));
  NO2        u0165(.A(i_2_), .B(i_1_), .Y(men_men_n188_));
  NA2        u0166(.A(men_men_n188_), .B(i_3_), .Y(men_men_n189_));
  NAi21      u0167(.An(i_4_), .B(i_12_), .Y(men_men_n190_));
  NO4        u0168(.A(men_men_n190_), .B(men_men_n189_), .C(men_men_n187_), .D(men_men_n25_), .Y(men_men_n191_));
  NO3        u0169(.A(men_men_n191_), .B(men_men_n184_), .C(men_men_n177_), .Y(men_men_n192_));
  INV        u0170(.A(i_8_), .Y(men_men_n193_));
  NO2        u0171(.A(men_men_n193_), .B(i_7_), .Y(men_men_n194_));
  NA2        u0172(.A(men_men_n194_), .B(i_6_), .Y(men_men_n195_));
  NO3        u0173(.A(i_3_), .B(men_men_n81_), .C(men_men_n48_), .Y(men_men_n196_));
  NA2        u0174(.A(men_men_n196_), .B(men_men_n111_), .Y(men_men_n197_));
  NO3        u0175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n198_));
  NA3        u0176(.A(men_men_n198_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n199_));
  NO3        u0177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n200_));
  OAI210     u0178(.A0(men_men_n94_), .A1(i_12_), .B0(men_men_n200_), .Y(men_men_n201_));
  AOI210     u0179(.A0(men_men_n201_), .A1(men_men_n199_), .B0(men_men_n197_), .Y(men_men_n202_));
  NO2        u0180(.A(i_3_), .B(i_8_), .Y(men_men_n203_));
  NO3        u0181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n204_));
  NA3        u0182(.A(men_men_n204_), .B(men_men_n203_), .C(men_men_n39_), .Y(men_men_n205_));
  NO2        u0183(.A(men_men_n101_), .B(men_men_n55_), .Y(men_men_n206_));
  NO2        u0184(.A(i_13_), .B(i_9_), .Y(men_men_n207_));
  NAi21      u0185(.An(i_12_), .B(i_3_), .Y(men_men_n208_));
  NO2        u0186(.A(men_men_n44_), .B(i_5_), .Y(men_men_n209_));
  NO3        u0187(.A(i_0_), .B(i_2_), .C(men_men_n60_), .Y(men_men_n210_));
  NA2        u0188(.A(men_men_n210_), .B(i_10_), .Y(men_men_n211_));
  OAI220     u0189(.A0(men_men_n211_), .A1(men_men_n208_), .B0(men_men_n101_), .B1(men_men_n205_), .Y(men_men_n212_));
  AOI210     u0190(.A0(men_men_n212_), .A1(i_7_), .B0(men_men_n202_), .Y(men_men_n213_));
  OAI220     u0191(.A0(men_men_n213_), .A1(i_4_), .B0(men_men_n195_), .B1(men_men_n192_), .Y(men_men_n214_));
  NAi21      u0192(.An(i_12_), .B(i_7_), .Y(men_men_n215_));
  NA3        u0193(.A(i_13_), .B(men_men_n193_), .C(i_10_), .Y(men_men_n216_));
  NO2        u0194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NA2        u0195(.A(i_0_), .B(i_5_), .Y(men_men_n218_));
  NA2        u0196(.A(men_men_n218_), .B(men_men_n102_), .Y(men_men_n219_));
  OAI220     u0197(.A0(men_men_n219_), .A1(men_men_n189_), .B0(men_men_n179_), .B1(men_men_n132_), .Y(men_men_n220_));
  NAi31      u0198(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n221_));
  NO2        u0199(.A(men_men_n36_), .B(i_13_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n68_), .B(men_men_n26_), .Y(men_men_n223_));
  NO2        u0201(.A(men_men_n46_), .B(men_men_n60_), .Y(men_men_n224_));
  NA3        u0202(.A(men_men_n224_), .B(men_men_n223_), .C(men_men_n222_), .Y(men_men_n225_));
  INV        u0203(.A(i_13_), .Y(men_men_n226_));
  NO2        u0204(.A(i_12_), .B(men_men_n226_), .Y(men_men_n227_));
  NA3        u0205(.A(men_men_n227_), .B(men_men_n198_), .C(men_men_n196_), .Y(men_men_n228_));
  OAI210     u0206(.A0(men_men_n225_), .A1(men_men_n221_), .B0(men_men_n228_), .Y(men_men_n229_));
  AOI220     u0207(.A0(men_men_n229_), .A1(men_men_n141_), .B0(men_men_n220_), .B1(men_men_n217_), .Y(men_men_n230_));
  NO2        u0208(.A(i_12_), .B(men_men_n37_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n182_), .B(i_4_), .Y(men_men_n232_));
  NA2        u0210(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  OR2        u0211(.A(i_8_), .B(i_7_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n234_), .B(men_men_n81_), .Y(men_men_n235_));
  NO2        u0213(.A(men_men_n51_), .B(i_1_), .Y(men_men_n236_));
  NA2        u0214(.A(men_men_n236_), .B(men_men_n235_), .Y(men_men_n237_));
  INV        u0215(.A(i_12_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n44_), .B(men_men_n238_), .Y(men_men_n239_));
  NO3        u0217(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n240_));
  NA2        u0218(.A(i_2_), .B(i_1_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n237_), .B(men_men_n233_), .Y(men_men_n242_));
  NO3        u0220(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n243_));
  NAi21      u0221(.An(i_4_), .B(i_3_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n244_), .B(men_men_n70_), .Y(men_men_n245_));
  NO2        u0223(.A(i_0_), .B(i_6_), .Y(men_men_n246_));
  NOi41      u0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n247_));
  NA2        u0225(.A(men_men_n247_), .B(men_men_n246_), .Y(men_men_n248_));
  NO2        u0226(.A(men_men_n241_), .B(men_men_n182_), .Y(men_men_n249_));
  NAi21      u0227(.An(men_men_n248_), .B(men_men_n249_), .Y(men_men_n250_));
  INV        u0228(.A(men_men_n250_), .Y(men_men_n251_));
  AOI220     u0229(.A0(men_men_n251_), .A1(men_men_n39_), .B0(men_men_n242_), .B1(men_men_n207_), .Y(men_men_n252_));
  NO2        u0230(.A(i_11_), .B(men_men_n226_), .Y(men_men_n253_));
  NOi21      u0231(.An(i_1_), .B(i_6_), .Y(men_men_n254_));
  NAi21      u0232(.An(i_3_), .B(i_7_), .Y(men_men_n255_));
  NA2        u0233(.A(men_men_n238_), .B(i_9_), .Y(men_men_n256_));
  OR4        u0234(.A(men_men_n256_), .B(men_men_n255_), .C(men_men_n254_), .D(men_men_n185_), .Y(men_men_n257_));
  NO2        u0235(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n258_));
  NO2        u0236(.A(i_12_), .B(i_3_), .Y(men_men_n259_));
  NA2        u0237(.A(men_men_n68_), .B(i_5_), .Y(men_men_n260_));
  NA2        u0238(.A(i_3_), .B(i_9_), .Y(men_men_n261_));
  NAi21      u0239(.An(i_7_), .B(i_10_), .Y(men_men_n262_));
  NO2        u0240(.A(men_men_n262_), .B(men_men_n261_), .Y(men_men_n263_));
  NA3        u0241(.A(men_men_n263_), .B(men_men_n260_), .C(men_men_n61_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n264_), .B(men_men_n257_), .Y(men_men_n265_));
  NA3        u0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n266_));
  NA2        u0244(.A(men_men_n238_), .B(i_13_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n265_), .B(men_men_n253_), .Y(men_men_n268_));
  NO2        u0246(.A(men_men_n234_), .B(men_men_n37_), .Y(men_men_n269_));
  NA2        u0247(.A(i_12_), .B(i_6_), .Y(men_men_n270_));
  OR2        u0248(.A(i_13_), .B(i_9_), .Y(men_men_n271_));
  NO3        u0249(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n48_), .Y(men_men_n272_));
  NO2        u0250(.A(men_men_n244_), .B(i_2_), .Y(men_men_n273_));
  NA3        u0251(.A(men_men_n273_), .B(men_men_n272_), .C(men_men_n44_), .Y(men_men_n274_));
  NA2        u0252(.A(men_men_n253_), .B(i_9_), .Y(men_men_n275_));
  OAI210     u0253(.A0(men_men_n68_), .A1(men_men_n275_), .B0(men_men_n274_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n154_), .B(men_men_n60_), .Y(men_men_n277_));
  NO3        u0255(.A(i_11_), .B(men_men_n226_), .C(men_men_n25_), .Y(men_men_n278_));
  NO2        u0256(.A(men_men_n255_), .B(i_8_), .Y(men_men_n279_));
  NO2        u0257(.A(i_6_), .B(men_men_n48_), .Y(men_men_n280_));
  NA3        u0258(.A(men_men_n280_), .B(men_men_n279_), .C(men_men_n278_), .Y(men_men_n281_));
  NO3        u0259(.A(men_men_n26_), .B(men_men_n81_), .C(i_5_), .Y(men_men_n282_));
  NA3        u0260(.A(men_men_n282_), .B(men_men_n269_), .C(men_men_n227_), .Y(men_men_n283_));
  AOI210     u0261(.A0(men_men_n283_), .A1(men_men_n281_), .B0(men_men_n277_), .Y(men_men_n284_));
  AOI210     u0262(.A0(men_men_n276_), .A1(men_men_n269_), .B0(men_men_n284_), .Y(men_men_n285_));
  NA4        u0263(.A(men_men_n285_), .B(men_men_n268_), .C(men_men_n252_), .D(men_men_n230_), .Y(men_men_n286_));
  NO3        u0264(.A(i_12_), .B(men_men_n226_), .C(men_men_n37_), .Y(men_men_n287_));
  INV        u0265(.A(men_men_n287_), .Y(men_men_n288_));
  NA2        u0266(.A(i_8_), .B(men_men_n99_), .Y(men_men_n289_));
  NOi21      u0267(.An(men_men_n163_), .B(men_men_n81_), .Y(men_men_n290_));
  NO3        u0268(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n291_));
  AOI220     u0269(.A0(men_men_n291_), .A1(men_men_n196_), .B0(men_men_n290_), .B1(men_men_n236_), .Y(men_men_n292_));
  NO2        u0270(.A(men_men_n292_), .B(men_men_n289_), .Y(men_men_n293_));
  NO3        u0271(.A(i_0_), .B(i_2_), .C(men_men_n60_), .Y(men_men_n294_));
  NO2        u0272(.A(men_men_n241_), .B(i_0_), .Y(men_men_n295_));
  AOI220     u0273(.A0(men_men_n295_), .A1(men_men_n194_), .B0(men_men_n294_), .B1(men_men_n141_), .Y(men_men_n296_));
  NA2        u0274(.A(men_men_n280_), .B(men_men_n26_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n297_), .B(men_men_n296_), .Y(men_men_n298_));
  NA2        u0276(.A(i_0_), .B(i_1_), .Y(men_men_n299_));
  NO2        u0277(.A(men_men_n299_), .B(i_2_), .Y(men_men_n300_));
  NO2        u0278(.A(men_men_n56_), .B(i_6_), .Y(men_men_n301_));
  NA3        u0279(.A(men_men_n301_), .B(men_men_n300_), .C(men_men_n163_), .Y(men_men_n302_));
  OAI210     u0280(.A0(men_men_n165_), .A1(men_men_n142_), .B0(men_men_n302_), .Y(men_men_n303_));
  NO3        u0281(.A(men_men_n303_), .B(men_men_n298_), .C(men_men_n293_), .Y(men_men_n304_));
  NO2        u0282(.A(i_3_), .B(i_10_), .Y(men_men_n305_));
  NA3        u0283(.A(men_men_n305_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n306_));
  NO2        u0284(.A(i_2_), .B(men_men_n99_), .Y(men_men_n307_));
  NOi21      u0285(.An(men_men_n218_), .B(men_men_n101_), .Y(men_men_n308_));
  NA3        u0286(.A(men_men_n308_), .B(i_1_), .C(men_men_n307_), .Y(men_men_n309_));
  AN2        u0287(.A(i_3_), .B(i_10_), .Y(men_men_n310_));
  NA4        u0288(.A(men_men_n310_), .B(men_men_n198_), .C(men_men_n175_), .D(men_men_n173_), .Y(men_men_n311_));
  NO2        u0289(.A(i_5_), .B(men_men_n37_), .Y(men_men_n312_));
  NO2        u0290(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n313_));
  OR2        u0291(.A(men_men_n309_), .B(men_men_n306_), .Y(men_men_n314_));
  OAI220     u0292(.A0(men_men_n314_), .A1(i_6_), .B0(men_men_n304_), .B1(men_men_n288_), .Y(men_men_n315_));
  NO4        u0293(.A(men_men_n315_), .B(men_men_n286_), .C(men_men_n214_), .D(men_men_n168_), .Y(men_men_n316_));
  NO3        u0294(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n317_));
  NO2        u0295(.A(men_men_n56_), .B(men_men_n81_), .Y(men_men_n318_));
  NA2        u0296(.A(men_men_n295_), .B(men_men_n318_), .Y(men_men_n319_));
  NO3        u0297(.A(i_6_), .B(men_men_n193_), .C(i_7_), .Y(men_men_n320_));
  NA2        u0298(.A(men_men_n320_), .B(men_men_n198_), .Y(men_men_n321_));
  AOI210     u0299(.A0(men_men_n321_), .A1(men_men_n319_), .B0(i_5_), .Y(men_men_n322_));
  NO2        u0300(.A(i_2_), .B(i_3_), .Y(men_men_n323_));
  OR2        u0301(.A(i_0_), .B(i_5_), .Y(men_men_n324_));
  NA2        u0302(.A(men_men_n218_), .B(men_men_n324_), .Y(men_men_n325_));
  NA4        u0303(.A(men_men_n325_), .B(men_men_n235_), .C(men_men_n323_), .D(i_1_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n295_), .B(men_men_n290_), .C(men_men_n111_), .Y(men_men_n327_));
  NAi21      u0305(.An(i_8_), .B(i_7_), .Y(men_men_n328_));
  NO2        u0306(.A(men_men_n157_), .B(men_men_n46_), .Y(men_men_n329_));
  NA3        u0307(.A(men_men_n329_), .B(i_7_), .C(men_men_n163_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n330_), .B(men_men_n327_), .C(men_men_n326_), .Y(men_men_n331_));
  OAI210     u0309(.A0(men_men_n331_), .A1(men_men_n322_), .B0(i_4_), .Y(men_men_n332_));
  NO2        u0310(.A(i_12_), .B(i_10_), .Y(men_men_n333_));
  NOi21      u0311(.An(i_5_), .B(i_0_), .Y(men_men_n334_));
  AOI210     u0312(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n99_), .Y(men_men_n335_));
  NO4        u0313(.A(men_men_n335_), .B(i_4_), .C(men_men_n334_), .D(men_men_n127_), .Y(men_men_n336_));
  NA4        u0314(.A(men_men_n79_), .B(men_men_n36_), .C(men_men_n81_), .D(i_8_), .Y(men_men_n337_));
  NA2        u0315(.A(men_men_n336_), .B(men_men_n333_), .Y(men_men_n338_));
  NO2        u0316(.A(i_6_), .B(i_8_), .Y(men_men_n339_));
  NOi21      u0317(.An(i_0_), .B(i_2_), .Y(men_men_n340_));
  AN2        u0318(.A(men_men_n340_), .B(men_men_n339_), .Y(men_men_n341_));
  NO2        u0319(.A(i_1_), .B(i_7_), .Y(men_men_n342_));
  NA3        u0320(.A(men_men_n339_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n343_));
  NA3        u0321(.A(men_men_n343_), .B(men_men_n338_), .C(men_men_n332_), .Y(men_men_n344_));
  NO3        u0322(.A(men_men_n234_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n345_));
  NO3        u0323(.A(men_men_n328_), .B(i_2_), .C(i_1_), .Y(men_men_n346_));
  OAI210     u0324(.A0(men_men_n346_), .A1(men_men_n345_), .B0(i_6_), .Y(men_men_n347_));
  NA3        u0325(.A(men_men_n254_), .B(men_men_n307_), .C(men_men_n193_), .Y(men_men_n348_));
  AOI210     u0326(.A0(men_men_n348_), .A1(men_men_n347_), .B0(men_men_n325_), .Y(men_men_n349_));
  NOi21      u0327(.An(men_men_n153_), .B(men_men_n102_), .Y(men_men_n350_));
  NO2        u0328(.A(men_men_n350_), .B(men_men_n123_), .Y(men_men_n351_));
  OAI210     u0329(.A0(men_men_n351_), .A1(men_men_n349_), .B0(i_3_), .Y(men_men_n352_));
  INV        u0330(.A(men_men_n79_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n299_), .B(men_men_n76_), .Y(men_men_n354_));
  NA2        u0332(.A(men_men_n354_), .B(men_men_n131_), .Y(men_men_n355_));
  NO2        u0333(.A(men_men_n90_), .B(men_men_n193_), .Y(men_men_n356_));
  NA3        u0334(.A(men_men_n308_), .B(men_men_n356_), .C(men_men_n60_), .Y(men_men_n357_));
  AOI210     u0335(.A0(men_men_n357_), .A1(men_men_n355_), .B0(men_men_n353_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n193_), .B(i_9_), .Y(men_men_n359_));
  NA3        u0337(.A(men_men_n359_), .B(men_men_n206_), .C(men_men_n157_), .Y(men_men_n360_));
  NO2        u0338(.A(men_men_n360_), .B(men_men_n46_), .Y(men_men_n361_));
  NO3        u0339(.A(men_men_n361_), .B(men_men_n358_), .C(men_men_n298_), .Y(men_men_n362_));
  AOI210     u0340(.A0(men_men_n362_), .A1(men_men_n352_), .B0(men_men_n162_), .Y(men_men_n363_));
  AOI210     u0341(.A0(men_men_n344_), .A1(men_men_n317_), .B0(men_men_n363_), .Y(men_men_n364_));
  NOi32      u0342(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n365_));
  INV        u0343(.A(men_men_n365_), .Y(men_men_n366_));
  NAi21      u0344(.An(i_0_), .B(i_6_), .Y(men_men_n367_));
  NAi21      u0345(.An(i_1_), .B(i_5_), .Y(men_men_n368_));
  NA2        u0346(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n369_));
  NA2        u0347(.A(men_men_n369_), .B(men_men_n25_), .Y(men_men_n370_));
  OAI210     u0348(.A0(men_men_n370_), .A1(men_men_n159_), .B0(men_men_n248_), .Y(men_men_n371_));
  NAi41      u0349(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n372_));
  OAI220     u0350(.A0(men_men_n372_), .A1(men_men_n368_), .B0(men_men_n221_), .B1(men_men_n159_), .Y(men_men_n373_));
  AOI210     u0351(.A0(men_men_n372_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n374_));
  NOi32      u0352(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n375_));
  NAi21      u0353(.An(i_6_), .B(i_1_), .Y(men_men_n376_));
  NA3        u0354(.A(men_men_n376_), .B(men_men_n375_), .C(men_men_n46_), .Y(men_men_n377_));
  NO2        u0355(.A(men_men_n377_), .B(i_0_), .Y(men_men_n378_));
  OR3        u0356(.A(men_men_n378_), .B(men_men_n374_), .C(men_men_n373_), .Y(men_men_n379_));
  NO2        u0357(.A(i_1_), .B(men_men_n99_), .Y(men_men_n380_));
  NAi21      u0358(.An(i_3_), .B(i_4_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n381_), .B(i_9_), .Y(men_men_n382_));
  AN2        u0360(.A(i_6_), .B(i_7_), .Y(men_men_n383_));
  OAI210     u0361(.A0(men_men_n383_), .A1(men_men_n380_), .B0(men_men_n382_), .Y(men_men_n384_));
  NA2        u0362(.A(i_2_), .B(i_7_), .Y(men_men_n385_));
  NO2        u0363(.A(men_men_n381_), .B(i_10_), .Y(men_men_n386_));
  NA3        u0364(.A(men_men_n386_), .B(men_men_n385_), .C(men_men_n246_), .Y(men_men_n387_));
  AOI210     u0365(.A0(men_men_n387_), .A1(men_men_n384_), .B0(men_men_n185_), .Y(men_men_n388_));
  AOI210     u0366(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n389_));
  AOI220     u0367(.A0(men_men_n386_), .A1(men_men_n342_), .B0(men_men_n240_), .B1(men_men_n188_), .Y(men_men_n390_));
  NO3        u0368(.A(men_men_n388_), .B(men_men_n379_), .C(men_men_n371_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n391_), .B(men_men_n366_), .Y(men_men_n392_));
  NO2        u0370(.A(men_men_n56_), .B(men_men_n25_), .Y(men_men_n393_));
  AN2        u0371(.A(i_12_), .B(i_5_), .Y(men_men_n394_));
  NO2        u0372(.A(i_4_), .B(men_men_n26_), .Y(men_men_n395_));
  NA2        u0373(.A(men_men_n395_), .B(men_men_n394_), .Y(men_men_n396_));
  NO2        u0374(.A(i_11_), .B(i_6_), .Y(men_men_n397_));
  NA3        u0375(.A(men_men_n397_), .B(men_men_n329_), .C(men_men_n226_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n398_), .B(men_men_n396_), .Y(men_men_n399_));
  NO2        u0377(.A(men_men_n244_), .B(i_5_), .Y(men_men_n400_));
  NO2        u0378(.A(i_5_), .B(i_10_), .Y(men_men_n401_));
  NA2        u0379(.A(men_men_n143_), .B(men_men_n45_), .Y(men_men_n402_));
  NO2        u0380(.A(men_men_n402_), .B(men_men_n244_), .Y(men_men_n403_));
  OAI210     u0381(.A0(men_men_n403_), .A1(men_men_n399_), .B0(men_men_n393_), .Y(men_men_n404_));
  NO2        u0382(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n405_));
  NO2        u0383(.A(men_men_n149_), .B(men_men_n81_), .Y(men_men_n406_));
  OAI210     u0384(.A0(men_men_n406_), .A1(men_men_n399_), .B0(men_men_n405_), .Y(men_men_n407_));
  NO3        u0385(.A(men_men_n81_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n408_));
  NO2        u0386(.A(i_3_), .B(men_men_n99_), .Y(men_men_n409_));
  NO2        u0387(.A(i_11_), .B(i_12_), .Y(men_men_n410_));
  NA2        u0388(.A(men_men_n401_), .B(men_men_n238_), .Y(men_men_n411_));
  NA3        u0389(.A(men_men_n111_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n412_));
  OAI220     u0390(.A0(men_men_n412_), .A1(men_men_n221_), .B0(men_men_n411_), .B1(men_men_n337_), .Y(men_men_n413_));
  NAi21      u0391(.An(i_13_), .B(i_0_), .Y(men_men_n414_));
  NO2        u0392(.A(men_men_n414_), .B(men_men_n241_), .Y(men_men_n415_));
  NA2        u0393(.A(men_men_n413_), .B(men_men_n415_), .Y(men_men_n416_));
  NA3        u0394(.A(men_men_n416_), .B(men_men_n407_), .C(men_men_n404_), .Y(men_men_n417_));
  NA2        u0395(.A(men_men_n44_), .B(men_men_n226_), .Y(men_men_n418_));
  NO3        u0396(.A(i_1_), .B(i_12_), .C(men_men_n81_), .Y(men_men_n419_));
  NO2        u0397(.A(i_0_), .B(i_11_), .Y(men_men_n420_));
  NOi21      u0398(.An(i_2_), .B(i_12_), .Y(men_men_n421_));
  NA2        u0399(.A(men_men_n421_), .B(i_6_), .Y(men_men_n422_));
  NO2        u0400(.A(men_men_n422_), .B(men_men_n1114_), .Y(men_men_n423_));
  NA2        u0401(.A(men_men_n141_), .B(i_9_), .Y(men_men_n424_));
  NO2        u0402(.A(men_men_n424_), .B(i_4_), .Y(men_men_n425_));
  NA2        u0403(.A(men_men_n423_), .B(men_men_n425_), .Y(men_men_n426_));
  NAi21      u0404(.An(i_9_), .B(i_4_), .Y(men_men_n427_));
  OR2        u0405(.A(i_13_), .B(i_10_), .Y(men_men_n428_));
  NO3        u0406(.A(men_men_n428_), .B(men_men_n116_), .C(men_men_n427_), .Y(men_men_n429_));
  NO2        u0407(.A(men_men_n172_), .B(men_men_n122_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n99_), .B(men_men_n25_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n287_), .B(men_men_n431_), .Y(men_men_n432_));
  NA2        u0410(.A(men_men_n280_), .B(men_men_n210_), .Y(men_men_n433_));
  OAI220     u0411(.A0(men_men_n433_), .A1(men_men_n216_), .B0(men_men_n432_), .B1(men_men_n350_), .Y(men_men_n434_));
  INV        u0412(.A(men_men_n434_), .Y(men_men_n435_));
  AOI210     u0413(.A0(men_men_n435_), .A1(men_men_n426_), .B0(men_men_n26_), .Y(men_men_n436_));
  NA2        u0414(.A(men_men_n327_), .B(men_men_n326_), .Y(men_men_n437_));
  AOI220     u0415(.A0(men_men_n301_), .A1(men_men_n291_), .B0(men_men_n295_), .B1(men_men_n318_), .Y(men_men_n438_));
  NO2        u0416(.A(men_men_n438_), .B(i_5_), .Y(men_men_n439_));
  NO2        u0417(.A(men_men_n182_), .B(men_men_n81_), .Y(men_men_n440_));
  AOI220     u0418(.A0(men_men_n440_), .A1(men_men_n300_), .B0(men_men_n282_), .B1(men_men_n210_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n441_), .B(men_men_n289_), .Y(men_men_n442_));
  NO3        u0420(.A(men_men_n442_), .B(men_men_n439_), .C(men_men_n437_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n196_), .B(men_men_n94_), .Y(men_men_n444_));
  NA3        u0422(.A(men_men_n329_), .B(men_men_n163_), .C(men_men_n81_), .Y(men_men_n445_));
  AOI210     u0423(.A0(men_men_n445_), .A1(men_men_n444_), .B0(men_men_n328_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n193_), .B(i_10_), .Y(men_men_n447_));
  NA3        u0425(.A(men_men_n260_), .B(men_men_n61_), .C(i_2_), .Y(men_men_n448_));
  NA2        u0426(.A(men_men_n301_), .B(men_men_n236_), .Y(men_men_n449_));
  OAI220     u0427(.A0(men_men_n449_), .A1(men_men_n182_), .B0(men_men_n448_), .B1(men_men_n447_), .Y(men_men_n450_));
  NO2        u0428(.A(i_3_), .B(men_men_n48_), .Y(men_men_n451_));
  NA3        u0429(.A(men_men_n342_), .B(men_men_n341_), .C(men_men_n451_), .Y(men_men_n452_));
  NA2        u0430(.A(men_men_n320_), .B(men_men_n325_), .Y(men_men_n453_));
  OAI210     u0431(.A0(men_men_n453_), .A1(men_men_n189_), .B0(men_men_n452_), .Y(men_men_n454_));
  NO3        u0432(.A(men_men_n454_), .B(men_men_n450_), .C(men_men_n446_), .Y(men_men_n455_));
  AOI210     u0433(.A0(men_men_n455_), .A1(men_men_n443_), .B0(men_men_n275_), .Y(men_men_n456_));
  NO4        u0434(.A(men_men_n456_), .B(men_men_n436_), .C(men_men_n417_), .D(men_men_n392_), .Y(men_men_n457_));
  NO2        u0435(.A(men_men_n60_), .B(i_4_), .Y(men_men_n458_));
  NO2        u0436(.A(men_men_n68_), .B(i_13_), .Y(men_men_n459_));
  NA3        u0437(.A(men_men_n459_), .B(men_men_n458_), .C(i_2_), .Y(men_men_n460_));
  NO2        u0438(.A(i_10_), .B(i_9_), .Y(men_men_n461_));
  NAi21      u0439(.An(i_12_), .B(i_8_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n462_), .B(i_3_), .Y(men_men_n463_));
  NA2        u0441(.A(men_men_n463_), .B(men_men_n461_), .Y(men_men_n464_));
  NA2        u0442(.A(i_2_), .B(men_men_n102_), .Y(men_men_n465_));
  OAI220     u0443(.A0(men_men_n465_), .A1(men_men_n205_), .B0(men_men_n464_), .B1(men_men_n460_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n313_), .B(i_0_), .Y(men_men_n467_));
  NO3        u0445(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n468_));
  NA2        u0446(.A(men_men_n270_), .B(men_men_n95_), .Y(men_men_n469_));
  NA2        u0447(.A(men_men_n469_), .B(men_men_n468_), .Y(men_men_n470_));
  NA2        u0448(.A(i_8_), .B(i_9_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n287_), .B(men_men_n206_), .Y(men_men_n472_));
  OAI220     u0450(.A0(men_men_n472_), .A1(men_men_n471_), .B0(men_men_n470_), .B1(men_men_n467_), .Y(men_men_n473_));
  NO3        u0451(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n474_));
  NA3        u0452(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n473_), .B(men_men_n466_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n300_), .B(men_men_n106_), .Y(men_men_n477_));
  OA210      u0455(.A0(men_men_n360_), .A1(men_men_n99_), .B0(men_men_n302_), .Y(men_men_n478_));
  OA220      u0456(.A0(men_men_n478_), .A1(men_men_n162_), .B0(men_men_n477_), .B1(men_men_n233_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n94_), .B(i_13_), .Y(men_men_n480_));
  NA2        u0458(.A(men_men_n440_), .B(men_men_n393_), .Y(men_men_n481_));
  NO2        u0459(.A(i_2_), .B(i_13_), .Y(men_men_n482_));
  NO2        u0460(.A(men_men_n481_), .B(men_men_n480_), .Y(men_men_n483_));
  NO3        u0461(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n484_));
  NO2        u0462(.A(i_6_), .B(i_7_), .Y(men_men_n485_));
  NA2        u0463(.A(men_men_n485_), .B(men_men_n484_), .Y(men_men_n486_));
  NO2        u0464(.A(i_11_), .B(i_1_), .Y(men_men_n487_));
  OR2        u0465(.A(i_11_), .B(i_8_), .Y(men_men_n488_));
  NOi21      u0466(.An(i_2_), .B(i_7_), .Y(men_men_n489_));
  NAi31      u0467(.An(men_men_n488_), .B(men_men_n489_), .C(men_men_n1115_), .Y(men_men_n490_));
  NO2        u0468(.A(men_men_n428_), .B(i_6_), .Y(men_men_n491_));
  NA3        u0469(.A(men_men_n491_), .B(men_men_n458_), .C(men_men_n70_), .Y(men_men_n492_));
  NO2        u0470(.A(men_men_n492_), .B(men_men_n490_), .Y(men_men_n493_));
  NO2        u0471(.A(i_3_), .B(men_men_n193_), .Y(men_men_n494_));
  NO2        u0472(.A(i_6_), .B(i_10_), .Y(men_men_n495_));
  NA4        u0473(.A(men_men_n495_), .B(men_men_n317_), .C(men_men_n494_), .D(men_men_n238_), .Y(men_men_n496_));
  NO2        u0474(.A(men_men_n496_), .B(men_men_n155_), .Y(men_men_n497_));
  NA3        u0475(.A(men_men_n247_), .B(men_men_n171_), .C(men_men_n131_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n499_));
  NO2        u0477(.A(men_men_n157_), .B(i_3_), .Y(men_men_n500_));
  NA3        u0478(.A(men_men_n405_), .B(men_men_n178_), .C(men_men_n148_), .Y(men_men_n501_));
  NA2        u0479(.A(men_men_n501_), .B(men_men_n498_), .Y(men_men_n502_));
  NO4        u0480(.A(men_men_n502_), .B(men_men_n497_), .C(men_men_n493_), .D(men_men_n483_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n468_), .B(men_men_n394_), .Y(men_men_n504_));
  NA2        u0482(.A(men_men_n474_), .B(men_men_n401_), .Y(men_men_n505_));
  OAI220     u0483(.A0(men_men_n505_), .A1(men_men_n225_), .B0(men_men_n504_), .B1(men_men_n54_), .Y(men_men_n506_));
  NAi21      u0484(.An(men_men_n216_), .B(men_men_n410_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n342_), .B(men_men_n218_), .Y(men_men_n508_));
  NO2        u0486(.A(men_men_n26_), .B(i_5_), .Y(men_men_n509_));
  NO2        u0487(.A(i_0_), .B(men_men_n81_), .Y(men_men_n510_));
  NA3        u0488(.A(men_men_n510_), .B(men_men_n509_), .C(men_men_n141_), .Y(men_men_n511_));
  OR3        u0489(.A(i_4_), .B(men_men_n38_), .C(men_men_n46_), .Y(men_men_n512_));
  OAI220     u0490(.A0(men_men_n512_), .A1(men_men_n511_), .B0(men_men_n508_), .B1(men_men_n507_), .Y(men_men_n513_));
  NA2        u0491(.A(men_men_n27_), .B(i_10_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n317_), .B(men_men_n240_), .Y(men_men_n515_));
  OAI220     u0493(.A0(men_men_n515_), .A1(men_men_n448_), .B0(men_men_n514_), .B1(men_men_n480_), .Y(men_men_n516_));
  NA4        u0494(.A(men_men_n310_), .B(men_men_n224_), .C(men_men_n68_), .D(men_men_n238_), .Y(men_men_n517_));
  NO2        u0495(.A(men_men_n517_), .B(men_men_n486_), .Y(men_men_n518_));
  NO4        u0496(.A(men_men_n518_), .B(men_men_n516_), .C(men_men_n513_), .D(men_men_n506_), .Y(men_men_n519_));
  NA4        u0497(.A(men_men_n519_), .B(men_men_n503_), .C(men_men_n479_), .D(men_men_n476_), .Y(men_men_n520_));
  NA3        u0498(.A(men_men_n310_), .B(men_men_n175_), .C(men_men_n173_), .Y(men_men_n521_));
  OAI210     u0499(.A0(men_men_n306_), .A1(men_men_n180_), .B0(men_men_n521_), .Y(men_men_n522_));
  AN2        u0500(.A(men_men_n291_), .B(men_men_n235_), .Y(men_men_n523_));
  NA2        u0501(.A(men_men_n523_), .B(men_men_n522_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n121_), .B(men_men_n110_), .Y(men_men_n525_));
  AO220      u0503(.A0(men_men_n525_), .A1(men_men_n468_), .B0(men_men_n429_), .B1(i_6_), .Y(men_men_n526_));
  NA2        u0504(.A(men_men_n317_), .B(men_men_n164_), .Y(men_men_n527_));
  OAI210     u0505(.A0(men_men_n527_), .A1(men_men_n233_), .B0(men_men_n311_), .Y(men_men_n528_));
  AOI220     u0506(.A0(men_men_n528_), .A1(i_7_), .B0(men_men_n526_), .B1(men_men_n313_), .Y(men_men_n529_));
  NA4        u0507(.A(men_men_n459_), .B(men_men_n458_), .C(men_men_n203_), .D(i_2_), .Y(men_men_n530_));
  INV        u0508(.A(men_men_n530_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n394_), .B(men_men_n226_), .Y(men_men_n532_));
  NA2        u0510(.A(men_men_n365_), .B(men_men_n68_), .Y(men_men_n533_));
  NA2        u0511(.A(men_men_n383_), .B(men_men_n375_), .Y(men_men_n534_));
  AO210      u0512(.A0(men_men_n533_), .A1(men_men_n532_), .B0(men_men_n534_), .Y(men_men_n535_));
  NO2        u0513(.A(men_men_n36_), .B(i_8_), .Y(men_men_n536_));
  NAi41      u0514(.An(men_men_n533_), .B(men_men_n495_), .C(men_men_n536_), .D(men_men_n46_), .Y(men_men_n537_));
  INV        u0515(.A(men_men_n429_), .Y(men_men_n538_));
  NA3        u0516(.A(men_men_n538_), .B(men_men_n537_), .C(men_men_n535_), .Y(men_men_n539_));
  AOI210     u0517(.A0(men_men_n531_), .A1(men_men_n204_), .B0(men_men_n539_), .Y(men_men_n540_));
  OAI210     u0518(.A0(i_8_), .A1(men_men_n60_), .B0(men_men_n133_), .Y(men_men_n541_));
  AOI210     u0519(.A0(men_men_n194_), .A1(i_9_), .B0(men_men_n269_), .Y(men_men_n542_));
  NO2        u0520(.A(men_men_n542_), .B(men_men_n199_), .Y(men_men_n543_));
  NO2        u0521(.A(men_men_n182_), .B(men_men_n81_), .Y(men_men_n544_));
  AOI220     u0522(.A0(men_men_n544_), .A1(men_men_n543_), .B0(men_men_n541_), .B1(men_men_n430_), .Y(men_men_n545_));
  NA4        u0523(.A(men_men_n545_), .B(men_men_n540_), .C(men_men_n529_), .D(men_men_n524_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n400_), .B(men_men_n300_), .Y(men_men_n547_));
  OAI210     u0525(.A0(men_men_n396_), .A1(men_men_n169_), .B0(men_men_n547_), .Y(men_men_n548_));
  NO2        u0526(.A(i_12_), .B(men_men_n193_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n549_), .B(men_men_n226_), .Y(men_men_n550_));
  NO3        u0528(.A(i_10_), .B(men_men_n550_), .C(men_men_n477_), .Y(men_men_n551_));
  NOi31      u0529(.An(men_men_n320_), .B(men_men_n428_), .C(men_men_n38_), .Y(men_men_n552_));
  OAI210     u0530(.A0(men_men_n552_), .A1(men_men_n551_), .B0(men_men_n548_), .Y(men_men_n553_));
  NO2        u0531(.A(i_8_), .B(i_7_), .Y(men_men_n554_));
  OAI210     u0532(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n555_));
  NA2        u0533(.A(men_men_n555_), .B(men_men_n224_), .Y(men_men_n556_));
  AOI220     u0534(.A0(men_men_n329_), .A1(men_men_n39_), .B0(men_men_n236_), .B1(men_men_n207_), .Y(men_men_n557_));
  OAI220     u0535(.A0(men_men_n557_), .A1(men_men_n182_), .B0(men_men_n556_), .B1(men_men_n244_), .Y(men_men_n558_));
  NA2        u0536(.A(men_men_n44_), .B(i_10_), .Y(men_men_n559_));
  NO2        u0537(.A(men_men_n559_), .B(i_6_), .Y(men_men_n560_));
  NA3        u0538(.A(men_men_n560_), .B(men_men_n558_), .C(men_men_n554_), .Y(men_men_n561_));
  AOI220     u0539(.A0(men_men_n440_), .A1(men_men_n329_), .B0(men_men_n249_), .B1(men_men_n246_), .Y(men_men_n562_));
  OAI220     u0540(.A0(men_men_n562_), .A1(men_men_n267_), .B0(men_men_n480_), .B1(men_men_n132_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n563_), .B(men_men_n269_), .Y(men_men_n564_));
  NOi31      u0542(.An(men_men_n295_), .B(men_men_n306_), .C(men_men_n180_), .Y(men_men_n565_));
  NA3        u0543(.A(men_men_n310_), .B(men_men_n173_), .C(men_men_n94_), .Y(men_men_n566_));
  NO2        u0544(.A(men_men_n222_), .B(men_men_n44_), .Y(men_men_n567_));
  NO2        u0545(.A(men_men_n157_), .B(i_5_), .Y(men_men_n568_));
  NA3        u0546(.A(men_men_n568_), .B(men_men_n418_), .C(men_men_n323_), .Y(men_men_n569_));
  OAI210     u0547(.A0(men_men_n569_), .A1(men_men_n567_), .B0(men_men_n566_), .Y(men_men_n570_));
  OAI210     u0548(.A0(men_men_n570_), .A1(men_men_n565_), .B0(men_men_n474_), .Y(men_men_n571_));
  NA4        u0549(.A(men_men_n571_), .B(men_men_n564_), .C(men_men_n561_), .D(men_men_n553_), .Y(men_men_n572_));
  NA3        u0550(.A(men_men_n218_), .B(men_men_n66_), .C(men_men_n44_), .Y(men_men_n573_));
  NA2        u0551(.A(men_men_n287_), .B(men_men_n79_), .Y(men_men_n574_));
  AOI210     u0552(.A0(men_men_n573_), .A1(men_men_n355_), .B0(men_men_n574_), .Y(men_men_n575_));
  NA2        u0553(.A(men_men_n301_), .B(men_men_n291_), .Y(men_men_n576_));
  NO2        u0554(.A(men_men_n576_), .B(men_men_n172_), .Y(men_men_n577_));
  NA2        u0555(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n578_));
  NA2        u0556(.A(men_men_n461_), .B(men_men_n222_), .Y(men_men_n579_));
  NO2        u0557(.A(men_men_n578_), .B(men_men_n579_), .Y(men_men_n580_));
  AOI210     u0558(.A0(men_men_n376_), .A1(men_men_n46_), .B0(men_men_n380_), .Y(men_men_n581_));
  NA2        u0559(.A(i_0_), .B(men_men_n48_), .Y(men_men_n582_));
  NA3        u0560(.A(men_men_n549_), .B(men_men_n278_), .C(men_men_n582_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n581_), .B(men_men_n583_), .Y(men_men_n584_));
  NO4        u0562(.A(men_men_n584_), .B(men_men_n580_), .C(men_men_n577_), .D(men_men_n575_), .Y(men_men_n585_));
  NO4        u0563(.A(men_men_n254_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n586_));
  NO3        u0564(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n234_), .B(men_men_n36_), .Y(men_men_n588_));
  AN2        u0566(.A(men_men_n588_), .B(men_men_n587_), .Y(men_men_n589_));
  OA210      u0567(.A0(men_men_n589_), .A1(men_men_n586_), .B0(men_men_n365_), .Y(men_men_n590_));
  NO2        u0568(.A(men_men_n428_), .B(i_1_), .Y(men_men_n591_));
  NOi31      u0569(.An(men_men_n591_), .B(men_men_n469_), .C(men_men_n68_), .Y(men_men_n592_));
  AN4        u0570(.A(men_men_n592_), .B(men_men_n425_), .C(men_men_n509_), .D(i_2_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n438_), .B(men_men_n176_), .Y(men_men_n594_));
  NO3        u0572(.A(men_men_n594_), .B(men_men_n593_), .C(men_men_n590_), .Y(men_men_n595_));
  NOi21      u0573(.An(i_10_), .B(i_6_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n81_), .B(men_men_n25_), .Y(men_men_n597_));
  AOI220     u0575(.A0(men_men_n287_), .A1(men_men_n597_), .B0(men_men_n278_), .B1(men_men_n596_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n598_), .B(men_men_n467_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n113_), .B(men_men_n23_), .Y(men_men_n600_));
  NA2        u0578(.A(men_men_n320_), .B(men_men_n164_), .Y(men_men_n601_));
  AOI220     u0579(.A0(men_men_n601_), .A1(men_men_n449_), .B0(men_men_n183_), .B1(men_men_n181_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n198_), .B(men_men_n37_), .Y(men_men_n603_));
  NOi31      u0581(.An(men_men_n145_), .B(men_men_n603_), .C(men_men_n337_), .Y(men_men_n604_));
  NO3        u0582(.A(men_men_n604_), .B(men_men_n602_), .C(men_men_n599_), .Y(men_men_n605_));
  NO2        u0583(.A(men_men_n533_), .B(men_men_n390_), .Y(men_men_n606_));
  INV        u0584(.A(men_men_n323_), .Y(men_men_n607_));
  NO2        u0585(.A(i_12_), .B(men_men_n81_), .Y(men_men_n608_));
  NA3        u0586(.A(men_men_n608_), .B(men_men_n278_), .C(men_men_n582_), .Y(men_men_n609_));
  NA3        u0587(.A(men_men_n397_), .B(men_men_n287_), .C(men_men_n218_), .Y(men_men_n610_));
  AOI210     u0588(.A0(men_men_n610_), .A1(men_men_n609_), .B0(men_men_n607_), .Y(men_men_n611_));
  NA2        u0589(.A(men_men_n173_), .B(i_0_), .Y(men_men_n612_));
  NO3        u0590(.A(men_men_n612_), .B(men_men_n347_), .C(men_men_n306_), .Y(men_men_n613_));
  OR2        u0591(.A(i_2_), .B(i_5_), .Y(men_men_n614_));
  OR2        u0592(.A(men_men_n614_), .B(i_6_), .Y(men_men_n615_));
  AOI210     u0593(.A0(men_men_n385_), .A1(men_men_n246_), .B0(men_men_n198_), .Y(men_men_n616_));
  AOI210     u0594(.A0(men_men_n616_), .A1(men_men_n615_), .B0(men_men_n507_), .Y(men_men_n617_));
  NO4        u0595(.A(men_men_n617_), .B(men_men_n613_), .C(men_men_n611_), .D(men_men_n606_), .Y(men_men_n618_));
  NA4        u0596(.A(men_men_n618_), .B(men_men_n605_), .C(men_men_n595_), .D(men_men_n585_), .Y(men_men_n619_));
  NO4        u0597(.A(men_men_n619_), .B(men_men_n572_), .C(men_men_n546_), .D(men_men_n520_), .Y(men_men_n620_));
  NA4        u0598(.A(men_men_n620_), .B(men_men_n457_), .C(men_men_n364_), .D(men_men_n316_), .Y(men7));
  NO2        u0599(.A(men_men_n106_), .B(men_men_n87_), .Y(men_men_n622_));
  NA2        u0600(.A(men_men_n395_), .B(men_men_n622_), .Y(men_men_n623_));
  NA2        u0601(.A(men_men_n495_), .B(men_men_n79_), .Y(men_men_n624_));
  NA2        u0602(.A(i_11_), .B(men_men_n193_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n143_), .B(men_men_n625_), .Y(men_men_n626_));
  OAI210     u0604(.A0(men_men_n626_), .A1(men_men_n624_), .B0(men_men_n623_), .Y(men_men_n627_));
  NA3        u0605(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n628_));
  NO2        u0606(.A(men_men_n238_), .B(i_4_), .Y(men_men_n629_));
  NA2        u0607(.A(men_men_n629_), .B(i_8_), .Y(men_men_n630_));
  NA2        u0608(.A(i_2_), .B(men_men_n81_), .Y(men_men_n631_));
  OAI210     u0609(.A0(men_men_n84_), .A1(men_men_n203_), .B0(men_men_n204_), .Y(men_men_n632_));
  NO2        u0610(.A(i_7_), .B(men_men_n37_), .Y(men_men_n633_));
  NA2        u0611(.A(i_4_), .B(i_8_), .Y(men_men_n634_));
  INV        u0612(.A(men_men_n627_), .Y(men_men_n635_));
  INV        u0613(.A(men_men_n161_), .Y(men_men_n636_));
  OR2        u0614(.A(i_6_), .B(i_10_), .Y(men_men_n637_));
  NO2        u0615(.A(men_men_n637_), .B(men_men_n23_), .Y(men_men_n638_));
  OR3        u0616(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n639_));
  NO3        u0617(.A(men_men_n639_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n640_));
  INV        u0618(.A(men_men_n200_), .Y(men_men_n641_));
  NO2        u0619(.A(men_men_n640_), .B(men_men_n638_), .Y(men_men_n642_));
  OA220      u0620(.A0(men_men_n642_), .A1(men_men_n607_), .B0(men_men_n636_), .B1(men_men_n271_), .Y(men_men_n643_));
  AOI210     u0621(.A0(men_men_n643_), .A1(men_men_n635_), .B0(men_men_n60_), .Y(men_men_n644_));
  NOi21      u0622(.An(i_11_), .B(i_7_), .Y(men_men_n645_));
  AO210      u0623(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n646_), .B(men_men_n645_), .Y(men_men_n647_));
  NA2        u0625(.A(men_men_n647_), .B(men_men_n207_), .Y(men_men_n648_));
  NA3        u0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n649_));
  NAi31      u0627(.An(men_men_n649_), .B(men_men_n215_), .C(i_11_), .Y(men_men_n650_));
  AOI210     u0628(.A0(men_men_n650_), .A1(men_men_n648_), .B0(men_men_n60_), .Y(men_men_n651_));
  NA2        u0629(.A(men_men_n83_), .B(men_men_n60_), .Y(men_men_n652_));
  AO210      u0630(.A0(men_men_n652_), .A1(men_men_n390_), .B0(men_men_n40_), .Y(men_men_n653_));
  NO3        u0631(.A(men_men_n262_), .B(men_men_n208_), .C(men_men_n625_), .Y(men_men_n654_));
  OAI210     u0632(.A0(men_men_n654_), .A1(men_men_n227_), .B0(men_men_n60_), .Y(men_men_n655_));
  NA2        u0633(.A(men_men_n421_), .B(men_men_n31_), .Y(men_men_n656_));
  OR2        u0634(.A(men_men_n208_), .B(men_men_n106_), .Y(men_men_n657_));
  NA2        u0635(.A(men_men_n657_), .B(men_men_n656_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n60_), .B(i_9_), .Y(men_men_n659_));
  NO2        u0637(.A(men_men_n659_), .B(i_4_), .Y(men_men_n660_));
  NA2        u0638(.A(men_men_n660_), .B(men_men_n658_), .Y(men_men_n661_));
  NO2        u0639(.A(i_1_), .B(i_12_), .Y(men_men_n662_));
  NA3        u0640(.A(men_men_n662_), .B(men_men_n108_), .C(men_men_n24_), .Y(men_men_n663_));
  NA4        u0641(.A(men_men_n663_), .B(men_men_n661_), .C(men_men_n655_), .D(men_men_n653_), .Y(men_men_n664_));
  OAI210     u0642(.A0(men_men_n664_), .A1(men_men_n651_), .B0(i_6_), .Y(men_men_n665_));
  NO2        u0643(.A(men_men_n649_), .B(men_men_n106_), .Y(men_men_n666_));
  NA2        u0644(.A(men_men_n666_), .B(men_men_n608_), .Y(men_men_n667_));
  NO2        u0645(.A(i_6_), .B(i_11_), .Y(men_men_n668_));
  NA3        u0646(.A(men_men_n667_), .B(men_men_n538_), .C(men_men_n470_), .Y(men_men_n669_));
  NO4        u0647(.A(men_men_n215_), .B(men_men_n127_), .C(i_13_), .D(men_men_n81_), .Y(men_men_n670_));
  NA2        u0648(.A(men_men_n670_), .B(men_men_n659_), .Y(men_men_n671_));
  NO3        u0649(.A(men_men_n637_), .B(men_men_n234_), .C(men_men_n23_), .Y(men_men_n672_));
  AOI210     u0650(.A0(i_1_), .A1(men_men_n263_), .B0(men_men_n672_), .Y(men_men_n673_));
  OAI210     u0651(.A0(men_men_n673_), .A1(men_men_n44_), .B0(men_men_n671_), .Y(men_men_n674_));
  NA3        u0652(.A(men_men_n554_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n137_), .B(i_9_), .Y(men_men_n676_));
  NA3        u0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n677_));
  NO2        u0655(.A(men_men_n46_), .B(i_1_), .Y(men_men_n678_));
  NA3        u0656(.A(men_men_n678_), .B(men_men_n270_), .C(men_men_n44_), .Y(men_men_n679_));
  OAI220     u0657(.A0(men_men_n679_), .A1(men_men_n677_), .B0(men_men_n676_), .B1(men_men_n1113_), .Y(men_men_n680_));
  NA3        u0658(.A(men_men_n659_), .B(men_men_n323_), .C(i_6_), .Y(men_men_n681_));
  NO2        u0659(.A(men_men_n681_), .B(men_men_n23_), .Y(men_men_n682_));
  AOI210     u0660(.A0(men_men_n487_), .A1(men_men_n431_), .B0(men_men_n243_), .Y(men_men_n683_));
  NO2        u0661(.A(men_men_n683_), .B(men_men_n631_), .Y(men_men_n684_));
  NAi21      u0662(.An(men_men_n675_), .B(men_men_n89_), .Y(men_men_n685_));
  NA2        u0663(.A(men_men_n678_), .B(men_men_n270_), .Y(men_men_n686_));
  NO2        u0664(.A(i_11_), .B(men_men_n37_), .Y(men_men_n687_));
  NA2        u0665(.A(men_men_n687_), .B(men_men_n24_), .Y(men_men_n688_));
  OAI210     u0666(.A0(men_men_n688_), .A1(men_men_n686_), .B0(men_men_n685_), .Y(men_men_n689_));
  OR4        u0667(.A(men_men_n689_), .B(men_men_n684_), .C(men_men_n682_), .D(men_men_n680_), .Y(men_men_n690_));
  NO3        u0668(.A(men_men_n690_), .B(men_men_n674_), .C(men_men_n669_), .Y(men_men_n691_));
  NO2        u0669(.A(men_men_n238_), .B(men_men_n99_), .Y(men_men_n692_));
  NO2        u0670(.A(men_men_n692_), .B(men_men_n645_), .Y(men_men_n693_));
  NA2        u0671(.A(men_men_n693_), .B(i_1_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n694_), .B(men_men_n639_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n427_), .B(men_men_n81_), .Y(men_men_n696_));
  NA2        u0674(.A(men_men_n695_), .B(men_men_n46_), .Y(men_men_n697_));
  NA2        u0675(.A(i_3_), .B(men_men_n193_), .Y(men_men_n698_));
  AOI210     u0676(.A0(men_men_n261_), .A1(men_men_n698_), .B0(men_men_n113_), .Y(men_men_n699_));
  AN2        u0677(.A(men_men_n699_), .B(men_men_n560_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n234_), .B(men_men_n44_), .Y(men_men_n701_));
  NO3        u0679(.A(men_men_n701_), .B(men_men_n313_), .C(men_men_n239_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n116_), .B(men_men_n37_), .Y(men_men_n703_));
  NO2        u0681(.A(men_men_n703_), .B(i_6_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n81_), .B(i_9_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(men_men_n60_), .Y(men_men_n706_));
  NO2        u0684(.A(men_men_n706_), .B(men_men_n662_), .Y(men_men_n707_));
  NO4        u0685(.A(men_men_n707_), .B(men_men_n704_), .C(men_men_n702_), .D(i_4_), .Y(men_men_n708_));
  NA2        u0686(.A(i_1_), .B(i_3_), .Y(men_men_n709_));
  NO2        u0687(.A(men_men_n471_), .B(men_men_n90_), .Y(men_men_n710_));
  AOI210     u0688(.A0(men_men_n701_), .A1(men_men_n596_), .B0(men_men_n710_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n711_), .B(men_men_n709_), .Y(men_men_n712_));
  NO3        u0690(.A(men_men_n712_), .B(men_men_n708_), .C(men_men_n700_), .Y(men_men_n713_));
  NA4        u0691(.A(men_men_n713_), .B(men_men_n697_), .C(men_men_n691_), .D(men_men_n665_), .Y(men_men_n714_));
  NO3        u0692(.A(men_men_n488_), .B(i_3_), .C(i_7_), .Y(men_men_n715_));
  NOi21      u0693(.An(men_men_n715_), .B(i_10_), .Y(men_men_n716_));
  OA210      u0694(.A0(men_men_n716_), .A1(men_men_n247_), .B0(men_men_n81_), .Y(men_men_n717_));
  NA2        u0695(.A(men_men_n383_), .B(men_men_n382_), .Y(men_men_n718_));
  NA3        u0696(.A(men_men_n495_), .B(men_men_n536_), .C(men_men_n46_), .Y(men_men_n719_));
  NO3        u0697(.A(men_men_n489_), .B(men_men_n634_), .C(men_men_n81_), .Y(men_men_n720_));
  NA2        u0698(.A(men_men_n720_), .B(men_men_n25_), .Y(men_men_n721_));
  NA3        u0699(.A(men_men_n161_), .B(men_men_n79_), .C(men_men_n81_), .Y(men_men_n722_));
  NA4        u0700(.A(men_men_n722_), .B(men_men_n721_), .C(men_men_n719_), .D(men_men_n718_), .Y(men_men_n723_));
  OAI210     u0701(.A0(men_men_n723_), .A1(men_men_n717_), .B0(i_1_), .Y(men_men_n724_));
  AOI210     u0702(.A0(men_men_n270_), .A1(men_men_n95_), .B0(i_1_), .Y(men_men_n725_));
  NO2        u0703(.A(men_men_n381_), .B(i_2_), .Y(men_men_n726_));
  NA2        u0704(.A(men_men_n726_), .B(men_men_n725_), .Y(men_men_n727_));
  OAI210     u0705(.A0(men_men_n681_), .A1(men_men_n462_), .B0(men_men_n727_), .Y(men_men_n728_));
  INV        u0706(.A(men_men_n728_), .Y(men_men_n729_));
  AOI210     u0707(.A0(men_men_n729_), .A1(men_men_n724_), .B0(i_13_), .Y(men_men_n730_));
  OR2        u0708(.A(i_11_), .B(i_7_), .Y(men_men_n731_));
  NA3        u0709(.A(men_men_n731_), .B(men_men_n104_), .C(men_men_n137_), .Y(men_men_n732_));
  AOI220     u0710(.A0(men_men_n482_), .A1(men_men_n161_), .B0(i_2_), .B1(men_men_n137_), .Y(men_men_n733_));
  OAI210     u0711(.A0(men_men_n733_), .A1(men_men_n44_), .B0(men_men_n732_), .Y(men_men_n734_));
  AOI210     u0712(.A0(men_men_n677_), .A1(men_men_n52_), .B0(i_12_), .Y(men_men_n735_));
  INV        u0713(.A(men_men_n735_), .Y(men_men_n736_));
  NO2        u0714(.A(men_men_n489_), .B(men_men_n24_), .Y(men_men_n737_));
  AOI220     u0715(.A0(men_men_n737_), .A1(men_men_n696_), .B0(men_men_n247_), .B1(men_men_n130_), .Y(men_men_n738_));
  OAI220     u0716(.A0(men_men_n738_), .A1(men_men_n40_), .B0(men_men_n736_), .B1(men_men_n90_), .Y(men_men_n739_));
  AOI210     u0717(.A0(men_men_n734_), .A1(men_men_n339_), .B0(men_men_n739_), .Y(men_men_n740_));
  NA2        u0718(.A(men_men_n113_), .B(men_men_n106_), .Y(men_men_n741_));
  AOI220     u0719(.A0(men_men_n741_), .A1(men_men_n67_), .B0(men_men_n397_), .B1(men_men_n678_), .Y(men_men_n742_));
  NO2        u0720(.A(men_men_n742_), .B(men_men_n244_), .Y(men_men_n743_));
  AOI210     u0721(.A0(men_men_n462_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n744_));
  NOi31      u0722(.An(men_men_n744_), .B(men_men_n624_), .C(men_men_n44_), .Y(men_men_n745_));
  NA2        u0723(.A(men_men_n126_), .B(i_13_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n677_), .B(men_men_n113_), .Y(men_men_n747_));
  INV        u0725(.A(men_men_n747_), .Y(men_men_n748_));
  OAI220     u0726(.A0(men_men_n748_), .A1(men_men_n66_), .B0(men_men_n746_), .B1(men_men_n725_), .Y(men_men_n749_));
  NO3        u0727(.A(men_men_n66_), .B(men_men_n32_), .C(men_men_n99_), .Y(men_men_n750_));
  NA2        u0728(.A(men_men_n26_), .B(men_men_n193_), .Y(men_men_n751_));
  NA2        u0729(.A(men_men_n751_), .B(i_7_), .Y(men_men_n752_));
  NO3        u0730(.A(men_men_n489_), .B(men_men_n238_), .C(men_men_n81_), .Y(men_men_n753_));
  AOI210     u0731(.A0(men_men_n753_), .A1(men_men_n752_), .B0(men_men_n750_), .Y(men_men_n754_));
  AOI220     u0732(.A0(men_men_n397_), .A1(men_men_n678_), .B0(men_men_n89_), .B1(men_men_n100_), .Y(men_men_n755_));
  OAI220     u0733(.A0(men_men_n755_), .A1(men_men_n630_), .B0(men_men_n754_), .B1(men_men_n641_), .Y(men_men_n756_));
  NO4        u0734(.A(men_men_n756_), .B(men_men_n749_), .C(men_men_n745_), .D(men_men_n743_), .Y(men_men_n757_));
  OR2        u0735(.A(i_11_), .B(i_6_), .Y(men_men_n758_));
  NA3        u0736(.A(men_men_n629_), .B(men_men_n751_), .C(i_7_), .Y(men_men_n759_));
  AOI210     u0737(.A0(men_men_n759_), .A1(men_men_n748_), .B0(men_men_n758_), .Y(men_men_n760_));
  NA3        u0738(.A(men_men_n421_), .B(men_men_n633_), .C(men_men_n95_), .Y(men_men_n761_));
  NA2        u0739(.A(men_men_n668_), .B(i_13_), .Y(men_men_n762_));
  NA2        u0740(.A(men_men_n100_), .B(men_men_n751_), .Y(men_men_n763_));
  NAi21      u0741(.An(i_11_), .B(i_12_), .Y(men_men_n764_));
  NOi41      u0742(.An(men_men_n109_), .B(men_men_n764_), .C(i_13_), .D(men_men_n81_), .Y(men_men_n765_));
  NO3        u0743(.A(men_men_n489_), .B(men_men_n608_), .C(men_men_n634_), .Y(men_men_n766_));
  AOI220     u0744(.A0(men_men_n766_), .A1(men_men_n317_), .B0(men_men_n765_), .B1(men_men_n763_), .Y(men_men_n767_));
  NA3        u0745(.A(men_men_n767_), .B(men_men_n762_), .C(men_men_n761_), .Y(men_men_n768_));
  OAI210     u0746(.A0(men_men_n768_), .A1(men_men_n760_), .B0(men_men_n60_), .Y(men_men_n769_));
  NO2        u0747(.A(i_2_), .B(i_12_), .Y(men_men_n770_));
  NA2        u0748(.A(men_men_n380_), .B(men_men_n770_), .Y(men_men_n771_));
  NA2        u0749(.A(i_8_), .B(men_men_n25_), .Y(men_men_n772_));
  NO3        u0750(.A(men_men_n772_), .B(men_men_n395_), .C(men_men_n629_), .Y(men_men_n773_));
  OAI210     u0751(.A0(men_men_n773_), .A1(men_men_n382_), .B0(men_men_n380_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n127_), .B(i_2_), .Y(men_men_n775_));
  NA2        u0753(.A(men_men_n775_), .B(men_men_n662_), .Y(men_men_n776_));
  NA3        u0754(.A(men_men_n776_), .B(men_men_n774_), .C(men_men_n771_), .Y(men_men_n777_));
  NA3        u0755(.A(men_men_n777_), .B(men_men_n45_), .C(men_men_n226_), .Y(men_men_n778_));
  NA4        u0756(.A(men_men_n778_), .B(men_men_n769_), .C(men_men_n757_), .D(men_men_n740_), .Y(men_men_n779_));
  OR4        u0757(.A(men_men_n779_), .B(men_men_n730_), .C(men_men_n714_), .D(men_men_n644_), .Y(men5));
  AOI210     u0758(.A0(men_men_n693_), .A1(men_men_n273_), .B0(men_men_n430_), .Y(men_men_n781_));
  NO2        u0759(.A(men_men_n630_), .B(i_11_), .Y(men_men_n782_));
  OAI210     u0760(.A0(men_men_n633_), .A1(men_men_n84_), .B0(men_men_n782_), .Y(men_men_n783_));
  NA3        u0761(.A(men_men_n783_), .B(men_men_n781_), .C(men_men_n538_), .Y(men_men_n784_));
  NO3        u0762(.A(i_11_), .B(men_men_n238_), .C(i_13_), .Y(men_men_n785_));
  NO2        u0763(.A(men_men_n123_), .B(men_men_n23_), .Y(men_men_n786_));
  NA2        u0764(.A(i_12_), .B(i_8_), .Y(men_men_n787_));
  OAI210     u0765(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n787_), .Y(men_men_n788_));
  INV        u0766(.A(men_men_n461_), .Y(men_men_n789_));
  AOI220     u0767(.A0(men_men_n323_), .A1(men_men_n600_), .B0(men_men_n788_), .B1(men_men_n786_), .Y(men_men_n790_));
  INV        u0768(.A(men_men_n790_), .Y(men_men_n791_));
  NO2        u0769(.A(men_men_n791_), .B(men_men_n784_), .Y(men_men_n792_));
  INV        u0770(.A(men_men_n171_), .Y(men_men_n793_));
  INV        u0771(.A(men_men_n247_), .Y(men_men_n794_));
  OAI210     u0772(.A0(men_men_n726_), .A1(men_men_n463_), .B0(men_men_n109_), .Y(men_men_n795_));
  AOI210     u0773(.A0(men_men_n795_), .A1(men_men_n794_), .B0(men_men_n793_), .Y(men_men_n796_));
  NO2        u0774(.A(men_men_n471_), .B(men_men_n26_), .Y(men_men_n797_));
  NO2        u0775(.A(men_men_n797_), .B(men_men_n431_), .Y(men_men_n798_));
  NA2        u0776(.A(men_men_n798_), .B(i_2_), .Y(men_men_n799_));
  INV        u0777(.A(men_men_n799_), .Y(men_men_n800_));
  AOI210     u0778(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n428_), .Y(men_men_n801_));
  AOI210     u0779(.A0(men_men_n801_), .A1(men_men_n800_), .B0(men_men_n796_), .Y(men_men_n802_));
  NO2        u0780(.A(men_men_n190_), .B(men_men_n124_), .Y(men_men_n803_));
  OAI210     u0781(.A0(men_men_n803_), .A1(men_men_n786_), .B0(i_2_), .Y(men_men_n804_));
  INV        u0782(.A(men_men_n172_), .Y(men_men_n805_));
  NA2        u0783(.A(men_men_n805_), .B(men_men_n84_), .Y(men_men_n806_));
  AOI210     u0784(.A0(men_men_n806_), .A1(men_men_n804_), .B0(men_men_n193_), .Y(men_men_n807_));
  OA210      u0785(.A0(men_men_n647_), .A1(men_men_n125_), .B0(i_13_), .Y(men_men_n808_));
  NA2        u0786(.A(men_men_n200_), .B(men_men_n203_), .Y(men_men_n809_));
  NA2        u0787(.A(men_men_n151_), .B(men_men_n625_), .Y(men_men_n810_));
  AOI210     u0788(.A0(men_men_n810_), .A1(men_men_n809_), .B0(men_men_n385_), .Y(men_men_n811_));
  AOI210     u0789(.A0(men_men_n208_), .A1(men_men_n147_), .B0(men_men_n536_), .Y(men_men_n812_));
  OAI210     u0790(.A0(men_men_n812_), .A1(men_men_n227_), .B0(men_men_n431_), .Y(men_men_n813_));
  NO2        u0791(.A(men_men_n100_), .B(men_men_n44_), .Y(men_men_n814_));
  INV        u0792(.A(men_men_n307_), .Y(men_men_n815_));
  NA4        u0793(.A(men_men_n815_), .B(men_men_n310_), .C(men_men_n123_), .D(men_men_n42_), .Y(men_men_n816_));
  OAI210     u0794(.A0(men_men_n816_), .A1(men_men_n814_), .B0(men_men_n813_), .Y(men_men_n817_));
  NO4        u0795(.A(men_men_n817_), .B(men_men_n811_), .C(men_men_n808_), .D(men_men_n807_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n600_), .B(men_men_n28_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n785_), .B(men_men_n279_), .Y(men_men_n820_));
  NA2        u0798(.A(men_men_n820_), .B(men_men_n819_), .Y(men_men_n821_));
  NO2        u0799(.A(men_men_n59_), .B(i_12_), .Y(men_men_n822_));
  NO2        u0800(.A(men_men_n822_), .B(men_men_n125_), .Y(men_men_n823_));
  NO2        u0801(.A(men_men_n823_), .B(men_men_n625_), .Y(men_men_n824_));
  AOI220     u0802(.A0(men_men_n824_), .A1(men_men_n36_), .B0(men_men_n821_), .B1(men_men_n46_), .Y(men_men_n825_));
  NA4        u0803(.A(men_men_n825_), .B(men_men_n818_), .C(men_men_n802_), .D(men_men_n792_), .Y(men6));
  NO3        u0804(.A(men_men_n258_), .B(men_men_n312_), .C(i_1_), .Y(men_men_n827_));
  NO2        u0805(.A(men_men_n185_), .B(men_men_n138_), .Y(men_men_n828_));
  OAI210     u0806(.A0(men_men_n828_), .A1(men_men_n827_), .B0(men_men_n775_), .Y(men_men_n829_));
  NA4        u0807(.A(men_men_n401_), .B(men_men_n494_), .C(men_men_n66_), .D(men_men_n99_), .Y(men_men_n830_));
  INV        u0808(.A(men_men_n830_), .Y(men_men_n831_));
  NO2        u0809(.A(men_men_n221_), .B(men_men_n499_), .Y(men_men_n832_));
  NO2        u0810(.A(i_11_), .B(i_9_), .Y(men_men_n833_));
  NO3        u0811(.A(men_men_n832_), .B(men_men_n831_), .C(men_men_n334_), .Y(men_men_n834_));
  AO210      u0812(.A0(men_men_n834_), .A1(men_men_n829_), .B0(i_12_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n386_), .B(men_men_n342_), .Y(men_men_n836_));
  NA2        u0814(.A(men_men_n608_), .B(men_men_n60_), .Y(men_men_n837_));
  NA2        u0815(.A(men_men_n716_), .B(men_men_n66_), .Y(men_men_n838_));
  NA4        u0816(.A(men_men_n652_), .B(men_men_n838_), .C(men_men_n837_), .D(men_men_n836_), .Y(men_men_n839_));
  INV        u0817(.A(men_men_n197_), .Y(men_men_n840_));
  AOI220     u0818(.A0(men_men_n840_), .A1(men_men_n833_), .B0(men_men_n839_), .B1(men_men_n68_), .Y(men_men_n841_));
  INV        u0819(.A(men_men_n333_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n70_), .B(men_men_n130_), .Y(men_men_n843_));
  INV        u0821(.A(men_men_n123_), .Y(men_men_n844_));
  NA2        u0822(.A(men_men_n844_), .B(men_men_n46_), .Y(men_men_n845_));
  AOI210     u0823(.A0(men_men_n845_), .A1(men_men_n843_), .B0(men_men_n842_), .Y(men_men_n846_));
  NO2        u0824(.A(men_men_n32_), .B(i_11_), .Y(men_men_n847_));
  NA3        u0825(.A(men_men_n847_), .B(men_men_n485_), .C(men_men_n401_), .Y(men_men_n848_));
  NAi32      u0826(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n849_));
  AOI210     u0827(.A0(men_men_n758_), .A1(men_men_n82_), .B0(men_men_n849_), .Y(men_men_n850_));
  OAI210     u0828(.A0(men_men_n715_), .A1(men_men_n588_), .B0(men_men_n587_), .Y(men_men_n851_));
  NAi31      u0829(.An(men_men_n850_), .B(men_men_n851_), .C(men_men_n848_), .Y(men_men_n852_));
  OR2        u0830(.A(men_men_n852_), .B(men_men_n846_), .Y(men_men_n853_));
  AO220      u0831(.A0(men_men_n369_), .A1(men_men_n359_), .B0(men_men_n408_), .B1(men_men_n625_), .Y(men_men_n854_));
  NA3        u0832(.A(men_men_n854_), .B(men_men_n259_), .C(i_7_), .Y(men_men_n855_));
  OR2        u0833(.A(men_men_n647_), .B(men_men_n463_), .Y(men_men_n856_));
  NA3        u0834(.A(men_men_n856_), .B(men_men_n146_), .C(men_men_n64_), .Y(men_men_n857_));
  AO210      u0835(.A0(men_men_n505_), .A1(men_men_n789_), .B0(men_men_n36_), .Y(men_men_n858_));
  NA3        u0836(.A(men_men_n858_), .B(men_men_n857_), .C(men_men_n855_), .Y(men_men_n859_));
  OAI210     u0837(.A0(i_6_), .A1(i_11_), .B0(men_men_n82_), .Y(men_men_n860_));
  AOI220     u0838(.A0(men_men_n860_), .A1(men_men_n587_), .B0(men_men_n832_), .B1(men_men_n752_), .Y(men_men_n861_));
  NA3        u0839(.A(men_men_n385_), .B(men_men_n240_), .C(men_men_n146_), .Y(men_men_n862_));
  OAI210     u0840(.A0(men_men_n408_), .A1(men_men_n204_), .B0(men_men_n65_), .Y(men_men_n863_));
  NA4        u0841(.A(men_men_n863_), .B(men_men_n862_), .C(men_men_n861_), .D(men_men_n632_), .Y(men_men_n864_));
  AO210      u0842(.A0(men_men_n536_), .A1(men_men_n46_), .B0(men_men_n83_), .Y(men_men_n865_));
  NA3        u0843(.A(men_men_n865_), .B(men_men_n495_), .C(men_men_n218_), .Y(men_men_n866_));
  AOI210     u0844(.A0(men_men_n463_), .A1(men_men_n461_), .B0(men_men_n586_), .Y(men_men_n867_));
  NO2        u0845(.A(men_men_n637_), .B(men_men_n100_), .Y(men_men_n868_));
  OAI210     u0846(.A0(men_men_n868_), .A1(men_men_n110_), .B0(men_men_n420_), .Y(men_men_n869_));
  NA2        u0847(.A(men_men_n246_), .B(men_men_n46_), .Y(men_men_n870_));
  NA2        u0848(.A(men_men_n870_), .B(men_men_n615_), .Y(men_men_n871_));
  NA3        u0849(.A(men_men_n871_), .B(men_men_n333_), .C(i_7_), .Y(men_men_n872_));
  NA4        u0850(.A(men_men_n872_), .B(men_men_n869_), .C(men_men_n867_), .D(men_men_n866_), .Y(men_men_n873_));
  NO4        u0851(.A(men_men_n873_), .B(men_men_n864_), .C(men_men_n859_), .D(men_men_n853_), .Y(men_men_n874_));
  NA4        u0852(.A(men_men_n874_), .B(men_men_n841_), .C(men_men_n835_), .D(men_men_n391_), .Y(men3));
  NA2        u0853(.A(i_12_), .B(i_10_), .Y(men_men_n876_));
  NA2        u0854(.A(i_6_), .B(i_7_), .Y(men_men_n877_));
  NO2        u0855(.A(men_men_n877_), .B(i_0_), .Y(men_men_n878_));
  NO2        u0856(.A(i_11_), .B(men_men_n238_), .Y(men_men_n879_));
  OAI210     u0857(.A0(men_men_n878_), .A1(men_men_n295_), .B0(men_men_n879_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n880_), .B(men_men_n193_), .Y(men_men_n881_));
  NO3        u0859(.A(men_men_n467_), .B(men_men_n87_), .C(men_men_n44_), .Y(men_men_n882_));
  OA210      u0860(.A0(men_men_n882_), .A1(men_men_n881_), .B0(men_men_n173_), .Y(men_men_n883_));
  NA3        u0861(.A(men_men_n862_), .B(men_men_n632_), .C(men_men_n384_), .Y(men_men_n884_));
  NA2        u0862(.A(men_men_n884_), .B(men_men_n39_), .Y(men_men_n885_));
  NOi21      u0863(.An(men_men_n94_), .B(men_men_n798_), .Y(men_men_n886_));
  NO3        u0864(.A(men_men_n657_), .B(men_men_n471_), .C(men_men_n130_), .Y(men_men_n887_));
  NA2        u0865(.A(men_men_n421_), .B(men_men_n45_), .Y(men_men_n888_));
  AN2        u0866(.A(men_men_n469_), .B(men_men_n53_), .Y(men_men_n889_));
  NO3        u0867(.A(men_men_n889_), .B(men_men_n887_), .C(men_men_n886_), .Y(men_men_n890_));
  AOI210     u0868(.A0(men_men_n890_), .A1(men_men_n885_), .B0(men_men_n48_), .Y(men_men_n891_));
  NO4        u0869(.A(men_men_n389_), .B(men_men_n394_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n892_));
  NA2        u0870(.A(men_men_n185_), .B(men_men_n596_), .Y(men_men_n893_));
  NOi21      u0871(.An(men_men_n893_), .B(men_men_n892_), .Y(men_men_n894_));
  NA2        u0872(.A(men_men_n744_), .B(men_men_n705_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n340_), .B(men_men_n451_), .Y(men_men_n896_));
  OAI220     u0874(.A0(men_men_n896_), .A1(men_men_n895_), .B0(men_men_n894_), .B1(men_men_n60_), .Y(men_men_n897_));
  NOi21      u0875(.An(i_5_), .B(i_9_), .Y(men_men_n898_));
  NA2        u0876(.A(men_men_n898_), .B(men_men_n459_), .Y(men_men_n899_));
  AOI210     u0877(.A0(men_men_n270_), .A1(men_men_n487_), .B0(men_men_n720_), .Y(men_men_n900_));
  NO3        u0878(.A(men_men_n424_), .B(men_men_n270_), .C(men_men_n68_), .Y(men_men_n901_));
  NO2        u0879(.A(men_men_n174_), .B(men_men_n147_), .Y(men_men_n902_));
  AOI210     u0880(.A0(men_men_n902_), .A1(men_men_n246_), .B0(men_men_n901_), .Y(men_men_n903_));
  OAI220     u0881(.A0(men_men_n903_), .A1(men_men_n180_), .B0(men_men_n900_), .B1(men_men_n899_), .Y(men_men_n904_));
  NO4        u0882(.A(men_men_n904_), .B(men_men_n897_), .C(men_men_n891_), .D(men_men_n883_), .Y(men_men_n905_));
  NOi21      u0883(.An(i_0_), .B(i_10_), .Y(men_men_n906_));
  NA2        u0884(.A(men_men_n185_), .B(men_men_n24_), .Y(men_men_n907_));
  NO2        u0885(.A(men_men_n703_), .B(men_men_n622_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n908_), .B(men_men_n907_), .Y(men_men_n909_));
  NA2        u0887(.A(men_men_n317_), .B(men_men_n128_), .Y(men_men_n910_));
  NAi21      u0888(.An(men_men_n162_), .B(men_men_n451_), .Y(men_men_n911_));
  OAI220     u0889(.A0(men_men_n911_), .A1(men_men_n870_), .B0(men_men_n910_), .B1(men_men_n411_), .Y(men_men_n912_));
  NO2        u0890(.A(men_men_n912_), .B(men_men_n909_), .Y(men_men_n913_));
  NO2        u0891(.A(men_men_n401_), .B(men_men_n299_), .Y(men_men_n914_));
  NA2        u0892(.A(men_men_n914_), .B(men_men_n747_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n597_), .B(i_0_), .Y(men_men_n916_));
  NO3        u0894(.A(men_men_n916_), .B(men_men_n396_), .C(men_men_n84_), .Y(men_men_n917_));
  NO4        u0895(.A(men_men_n614_), .B(men_men_n215_), .C(men_men_n428_), .D(i_6_), .Y(men_men_n918_));
  AOI210     u0896(.A0(men_men_n918_), .A1(i_11_), .B0(men_men_n917_), .Y(men_men_n919_));
  INV        u0897(.A(men_men_n485_), .Y(men_men_n920_));
  AN2        u0898(.A(men_men_n94_), .B(men_men_n245_), .Y(men_men_n921_));
  NA2        u0899(.A(men_men_n785_), .B(men_men_n334_), .Y(men_men_n922_));
  AOI210     u0900(.A0(men_men_n495_), .A1(men_men_n84_), .B0(men_men_n55_), .Y(men_men_n923_));
  OAI220     u0901(.A0(men_men_n923_), .A1(men_men_n922_), .B0(men_men_n688_), .B1(men_men_n556_), .Y(men_men_n924_));
  NO2        u0902(.A(men_men_n256_), .B(men_men_n153_), .Y(men_men_n925_));
  NA2        u0903(.A(i_0_), .B(i_10_), .Y(men_men_n926_));
  OAI210     u0904(.A0(men_men_n926_), .A1(men_men_n81_), .B0(men_men_n559_), .Y(men_men_n927_));
  NO4        u0905(.A(men_men_n113_), .B(men_men_n55_), .C(men_men_n698_), .D(i_5_), .Y(men_men_n928_));
  AO220      u0906(.A0(men_men_n928_), .A1(men_men_n927_), .B0(men_men_n925_), .B1(i_6_), .Y(men_men_n929_));
  AOI220     u0907(.A0(men_men_n340_), .A1(men_men_n96_), .B0(men_men_n185_), .B1(men_men_n79_), .Y(men_men_n930_));
  NA2        u0908(.A(men_men_n591_), .B(i_4_), .Y(men_men_n931_));
  NA2        u0909(.A(men_men_n188_), .B(men_men_n203_), .Y(men_men_n932_));
  OAI220     u0910(.A0(men_men_n932_), .A1(men_men_n922_), .B0(men_men_n931_), .B1(men_men_n930_), .Y(men_men_n933_));
  NO4        u0911(.A(men_men_n933_), .B(men_men_n929_), .C(men_men_n924_), .D(men_men_n921_), .Y(men_men_n934_));
  NA4        u0912(.A(men_men_n934_), .B(men_men_n919_), .C(men_men_n915_), .D(men_men_n913_), .Y(men_men_n935_));
  NO2        u0913(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n936_));
  NA2        u0914(.A(i_11_), .B(i_9_), .Y(men_men_n937_));
  NO3        u0915(.A(i_12_), .B(men_men_n937_), .C(men_men_n631_), .Y(men_men_n938_));
  AO220      u0916(.A0(men_men_n938_), .A1(men_men_n936_), .B0(men_men_n272_), .B1(men_men_n83_), .Y(men_men_n939_));
  NO2        u0917(.A(men_men_n48_), .B(i_7_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n405_), .B(men_men_n178_), .Y(men_men_n941_));
  NA2        u0919(.A(men_men_n941_), .B(men_men_n160_), .Y(men_men_n942_));
  NO2        u0920(.A(men_men_n937_), .B(men_men_n68_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n174_), .B(i_0_), .Y(men_men_n944_));
  INV        u0922(.A(men_men_n944_), .Y(men_men_n945_));
  NA2        u0923(.A(men_men_n485_), .B(men_men_n232_), .Y(men_men_n946_));
  AOI210     u0924(.A0(men_men_n383_), .A1(men_men_n41_), .B0(men_men_n419_), .Y(men_men_n947_));
  OAI220     u0925(.A0(men_men_n947_), .A1(men_men_n899_), .B0(men_men_n946_), .B1(men_men_n945_), .Y(men_men_n948_));
  NO3        u0926(.A(men_men_n948_), .B(men_men_n942_), .C(men_men_n939_), .Y(men_men_n949_));
  NA2        u0927(.A(men_men_n687_), .B(men_men_n120_), .Y(men_men_n950_));
  NO2        u0928(.A(i_6_), .B(men_men_n950_), .Y(men_men_n951_));
  AOI210     u0929(.A0(men_men_n462_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n952_));
  NA2        u0930(.A(men_men_n171_), .B(men_men_n101_), .Y(men_men_n953_));
  NOi32      u0931(.An(men_men_n952_), .Bn(men_men_n188_), .C(men_men_n953_), .Y(men_men_n954_));
  AOI210     u0932(.A0(men_men_n633_), .A1(men_men_n334_), .B0(men_men_n245_), .Y(men_men_n955_));
  NO2        u0933(.A(men_men_n955_), .B(men_men_n888_), .Y(men_men_n956_));
  NO3        u0934(.A(men_men_n956_), .B(men_men_n954_), .C(men_men_n951_), .Y(men_men_n957_));
  NOi21      u0935(.An(i_7_), .B(i_5_), .Y(men_men_n958_));
  NOi31      u0936(.An(men_men_n958_), .B(men_men_n906_), .C(men_men_n764_), .Y(men_men_n959_));
  NA3        u0937(.A(men_men_n959_), .B(men_men_n395_), .C(i_6_), .Y(men_men_n960_));
  OA210      u0938(.A0(men_men_n953_), .A1(men_men_n534_), .B0(men_men_n960_), .Y(men_men_n961_));
  NO3        u0939(.A(men_men_n414_), .B(men_men_n372_), .C(men_men_n368_), .Y(men_men_n962_));
  NO2        u0940(.A(men_men_n266_), .B(men_men_n324_), .Y(men_men_n963_));
  NO2        u0941(.A(men_men_n764_), .B(men_men_n261_), .Y(men_men_n964_));
  AOI210     u0942(.A0(men_men_n964_), .A1(men_men_n963_), .B0(men_men_n962_), .Y(men_men_n965_));
  NA4        u0943(.A(men_men_n965_), .B(men_men_n961_), .C(men_men_n957_), .D(men_men_n949_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n907_), .B(men_men_n241_), .Y(men_men_n967_));
  AN2        u0945(.A(men_men_n339_), .B(men_men_n334_), .Y(men_men_n968_));
  AO220      u0946(.A0(men_men_n968_), .A1(men_men_n902_), .B0(men_men_n354_), .B1(men_men_n27_), .Y(men_men_n969_));
  OAI210     u0947(.A0(men_men_n969_), .A1(men_men_n967_), .B0(i_10_), .Y(men_men_n970_));
  INV        u0948(.A(men_men_n876_), .Y(men_men_n971_));
  OA210      u0949(.A0(men_men_n485_), .A1(men_men_n224_), .B0(men_men_n484_), .Y(men_men_n972_));
  OAI210     u0950(.A0(men_men_n972_), .A1(men_men_n971_), .B0(men_men_n943_), .Y(men_men_n973_));
  NA3        u0951(.A(men_men_n484_), .B(men_men_n421_), .C(men_men_n45_), .Y(men_men_n974_));
  OAI210     u0952(.A0(men_men_n911_), .A1(men_men_n920_), .B0(men_men_n974_), .Y(men_men_n975_));
  NO2        u0953(.A(men_men_n259_), .B(men_men_n46_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n943_), .B(men_men_n310_), .Y(men_men_n977_));
  OAI210     u0955(.A0(men_men_n976_), .A1(men_men_n187_), .B0(men_men_n977_), .Y(men_men_n978_));
  AOI220     u0956(.A0(men_men_n978_), .A1(men_men_n485_), .B0(men_men_n975_), .B1(men_men_n68_), .Y(men_men_n979_));
  NA3        u0957(.A(i_5_), .B(men_men_n393_), .C(i_6_), .Y(men_men_n980_));
  NA2        u0958(.A(men_men_n90_), .B(men_men_n44_), .Y(men_men_n981_));
  NO2        u0959(.A(men_men_n70_), .B(men_men_n787_), .Y(men_men_n982_));
  AOI220     u0960(.A0(men_men_n982_), .A1(men_men_n981_), .B0(men_men_n173_), .B1(men_men_n622_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n983_), .A1(men_men_n980_), .B0(men_men_n47_), .Y(men_men_n984_));
  NO3        u0962(.A(men_men_n614_), .B(men_men_n367_), .C(men_men_n24_), .Y(men_men_n985_));
  AOI210     u0963(.A0(men_men_n737_), .A1(men_men_n568_), .B0(men_men_n985_), .Y(men_men_n986_));
  NAi21      u0964(.An(i_9_), .B(i_5_), .Y(men_men_n987_));
  NO2        u0965(.A(men_men_n987_), .B(men_men_n414_), .Y(men_men_n988_));
  NO2        u0966(.A(men_men_n628_), .B(men_men_n103_), .Y(men_men_n989_));
  AOI220     u0967(.A0(men_men_n989_), .A1(i_0_), .B0(men_men_n988_), .B1(men_men_n647_), .Y(men_men_n990_));
  OAI220     u0968(.A0(men_men_n990_), .A1(men_men_n81_), .B0(men_men_n986_), .B1(men_men_n172_), .Y(men_men_n991_));
  NO3        u0969(.A(men_men_n991_), .B(men_men_n984_), .C(men_men_n539_), .Y(men_men_n992_));
  NA4        u0970(.A(men_men_n992_), .B(men_men_n979_), .C(men_men_n973_), .D(men_men_n970_), .Y(men_men_n993_));
  NO3        u0971(.A(men_men_n993_), .B(men_men_n966_), .C(men_men_n935_), .Y(men_men_n994_));
  NO2        u0972(.A(men_men_n906_), .B(men_men_n764_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n68_), .B(men_men_n44_), .Y(men_men_n996_));
  NO3        u0974(.A(men_men_n103_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n997_));
  AO220      u0975(.A0(men_men_n997_), .A1(men_men_n44_), .B0(men_men_n995_), .B1(men_men_n173_), .Y(men_men_n998_));
  AOI210     u0976(.A0(men_men_n837_), .A1(men_men_n718_), .B0(men_men_n953_), .Y(men_men_n999_));
  AOI210     u0977(.A0(men_men_n998_), .A1(men_men_n356_), .B0(men_men_n999_), .Y(men_men_n1000_));
  NA2        u0978(.A(men_men_n775_), .B(men_men_n145_), .Y(men_men_n1001_));
  INV        u0979(.A(men_men_n1001_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n1002_), .B(men_men_n705_), .C(men_men_n68_), .Y(men_men_n1003_));
  NO2        u0981(.A(men_men_n851_), .B(men_men_n414_), .Y(men_men_n1004_));
  NA3        u0982(.A(men_men_n878_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n879_), .B(i_9_), .Y(men_men_n1006_));
  AOI210     u0984(.A0(men_men_n1005_), .A1(men_men_n511_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  OAI210     u0985(.A0(men_men_n246_), .A1(i_9_), .B0(men_men_n231_), .Y(men_men_n1008_));
  AOI210     u0986(.A0(men_men_n1008_), .A1(men_men_n916_), .B0(men_men_n153_), .Y(men_men_n1009_));
  NO3        u0987(.A(men_men_n1009_), .B(men_men_n1007_), .C(men_men_n1004_), .Y(men_men_n1010_));
  NA3        u0988(.A(men_men_n1010_), .B(men_men_n1003_), .C(men_men_n1000_), .Y(men_men_n1011_));
  NA2        u0989(.A(men_men_n968_), .B(men_men_n385_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n306_), .A1(men_men_n162_), .B0(men_men_n1012_), .Y(men_men_n1013_));
  NA3        u0991(.A(men_men_n39_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n1014_));
  NA2        u0992(.A(men_men_n940_), .B(men_men_n500_), .Y(men_men_n1015_));
  AOI210     u0993(.A0(men_men_n1014_), .A1(men_men_n162_), .B0(men_men_n1015_), .Y(men_men_n1016_));
  NO2        u0994(.A(men_men_n1016_), .B(men_men_n1013_), .Y(men_men_n1017_));
  NA2        u0995(.A(men_men_n592_), .B(men_men_n70_), .Y(men_men_n1018_));
  NO3        u0996(.A(men_men_n209_), .B(men_men_n394_), .C(i_0_), .Y(men_men_n1019_));
  OAI210     u0997(.A0(men_men_n1019_), .A1(men_men_n71_), .B0(i_13_), .Y(men_men_n1020_));
  INV        u0998(.A(men_men_n218_), .Y(men_men_n1021_));
  OAI220     u0999(.A0(men_men_n550_), .A1(men_men_n138_), .B0(i_12_), .B1(men_men_n641_), .Y(men_men_n1022_));
  NA3        u1000(.A(men_men_n1022_), .B(men_men_n409_), .C(men_men_n1021_), .Y(men_men_n1023_));
  NA4        u1001(.A(men_men_n1023_), .B(men_men_n1020_), .C(men_men_n1018_), .D(men_men_n1017_), .Y(men_men_n1024_));
  NO2        u1002(.A(men_men_n244_), .B(men_men_n90_), .Y(men_men_n1025_));
  AOI210     u1003(.A0(men_men_n1025_), .A1(men_men_n995_), .B0(men_men_n107_), .Y(men_men_n1026_));
  AOI220     u1004(.A0(men_men_n958_), .A1(men_men_n500_), .B0(men_men_n878_), .B1(men_men_n163_), .Y(men_men_n1027_));
  NA2        u1005(.A(men_men_n359_), .B(men_men_n175_), .Y(men_men_n1028_));
  OA220      u1006(.A0(men_men_n1028_), .A1(men_men_n1027_), .B0(men_men_n1026_), .B1(i_5_), .Y(men_men_n1029_));
  AOI210     u1007(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n174_), .Y(men_men_n1030_));
  NA2        u1008(.A(men_men_n1030_), .B(men_men_n972_), .Y(men_men_n1031_));
  NA3        u1009(.A(men_men_n638_), .B(men_men_n185_), .C(men_men_n79_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n1032_), .B(men_men_n566_), .Y(men_men_n1033_));
  NO3        u1011(.A(men_men_n888_), .B(men_men_n52_), .C(men_men_n48_), .Y(men_men_n1034_));
  NA2        u1012(.A(men_men_n504_), .B(men_men_n498_), .Y(men_men_n1035_));
  NO3        u1013(.A(men_men_n1035_), .B(men_men_n1034_), .C(men_men_n1033_), .Y(men_men_n1036_));
  NA3        u1014(.A(men_men_n940_), .B(men_men_n295_), .C(men_men_n231_), .Y(men_men_n1037_));
  INV        u1015(.A(men_men_n1037_), .Y(men_men_n1038_));
  NA3        u1016(.A(men_men_n401_), .B(men_men_n341_), .C(men_men_n222_), .Y(men_men_n1039_));
  OAI210     u1017(.A0(men_men_n893_), .A1(men_men_n675_), .B0(men_men_n1039_), .Y(men_men_n1040_));
  NOi31      u1018(.An(men_men_n400_), .B(men_men_n996_), .C(men_men_n241_), .Y(men_men_n1041_));
  NO3        u1019(.A(men_men_n1041_), .B(men_men_n1040_), .C(men_men_n1038_), .Y(men_men_n1042_));
  NA4        u1020(.A(men_men_n1042_), .B(men_men_n1036_), .C(men_men_n1031_), .D(men_men_n1029_), .Y(men_men_n1043_));
  INV        u1021(.A(men_men_n640_), .Y(men_men_n1044_));
  NO3        u1022(.A(men_men_n1044_), .B(men_men_n582_), .C(men_men_n353_), .Y(men_men_n1045_));
  NO2        u1023(.A(men_men_n81_), .B(i_5_), .Y(men_men_n1046_));
  NA3        u1024(.A(men_men_n879_), .B(men_men_n108_), .C(men_men_n123_), .Y(men_men_n1047_));
  INV        u1025(.A(men_men_n1047_), .Y(men_men_n1048_));
  AOI210     u1026(.A0(men_men_n1048_), .A1(men_men_n1046_), .B0(men_men_n1045_), .Y(men_men_n1049_));
  NA3        u1027(.A(men_men_n310_), .B(i_5_), .C(men_men_n193_), .Y(men_men_n1050_));
  NO4        u1028(.A(men_men_n241_), .B(men_men_n209_), .C(i_0_), .D(i_12_), .Y(men_men_n1051_));
  AOI220     u1029(.A0(men_men_n1051_), .A1(i_10_), .B0(men_men_n831_), .B1(men_men_n175_), .Y(men_men_n1052_));
  AN2        u1030(.A(men_men_n926_), .B(men_men_n153_), .Y(men_men_n1053_));
  NO4        u1031(.A(men_men_n1053_), .B(i_12_), .C(men_men_n675_), .D(men_men_n130_), .Y(men_men_n1054_));
  NA2        u1032(.A(men_men_n1054_), .B(men_men_n218_), .Y(men_men_n1055_));
  NA3        u1033(.A(men_men_n96_), .B(men_men_n596_), .C(i_11_), .Y(men_men_n1056_));
  NO2        u1034(.A(men_men_n1056_), .B(men_men_n155_), .Y(men_men_n1057_));
  NA2        u1035(.A(men_men_n958_), .B(men_men_n482_), .Y(men_men_n1058_));
  NA2        u1036(.A(men_men_n61_), .B(men_men_n99_), .Y(men_men_n1059_));
  OAI220     u1037(.A0(men_men_n1059_), .A1(men_men_n1050_), .B0(men_men_n1058_), .B1(men_men_n706_), .Y(men_men_n1060_));
  AOI210     u1038(.A0(men_men_n1060_), .A1(men_men_n944_), .B0(men_men_n1057_), .Y(men_men_n1061_));
  NA4        u1039(.A(men_men_n1061_), .B(men_men_n1055_), .C(men_men_n1052_), .D(men_men_n1049_), .Y(men_men_n1062_));
  NO4        u1040(.A(men_men_n1062_), .B(men_men_n1043_), .C(men_men_n1024_), .D(men_men_n1011_), .Y(men_men_n1063_));
  NA2        u1041(.A(men_men_n847_), .B(men_men_n37_), .Y(men_men_n1064_));
  NA3        u1042(.A(men_men_n952_), .B(men_men_n380_), .C(i_5_), .Y(men_men_n1065_));
  NA3        u1043(.A(men_men_n1065_), .B(men_men_n1064_), .C(men_men_n636_), .Y(men_men_n1066_));
  NA2        u1044(.A(men_men_n1066_), .B(men_men_n207_), .Y(men_men_n1067_));
  AN2        u1045(.A(men_men_n731_), .B(men_men_n381_), .Y(men_men_n1068_));
  NA2        u1046(.A(men_men_n186_), .B(men_men_n188_), .Y(men_men_n1069_));
  AO210      u1047(.A0(men_men_n1068_), .A1(men_men_n33_), .B0(men_men_n1069_), .Y(men_men_n1070_));
  OAI210     u1048(.A0(men_men_n640_), .A1(men_men_n638_), .B0(men_men_n323_), .Y(men_men_n1071_));
  NAi31      u1049(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1072_));
  AOI210     u1050(.A0(men_men_n116_), .A1(men_men_n65_), .B0(men_men_n1072_), .Y(men_men_n1073_));
  NO2        u1051(.A(men_men_n1073_), .B(men_men_n672_), .Y(men_men_n1074_));
  NA3        u1052(.A(men_men_n1074_), .B(men_men_n1071_), .C(men_men_n1070_), .Y(men_men_n1075_));
  NO2        u1053(.A(men_men_n475_), .B(men_men_n270_), .Y(men_men_n1076_));
  NO4        u1054(.A(men_men_n234_), .B(men_men_n144_), .C(men_men_n709_), .D(men_men_n37_), .Y(men_men_n1077_));
  NO3        u1055(.A(men_men_n1077_), .B(men_men_n1076_), .C(men_men_n918_), .Y(men_men_n1078_));
  OAI210     u1056(.A0(men_men_n1056_), .A1(men_men_n147_), .B0(men_men_n1078_), .Y(men_men_n1079_));
  AOI210     u1057(.A0(men_men_n1075_), .A1(men_men_n48_), .B0(men_men_n1079_), .Y(men_men_n1080_));
  AOI210     u1058(.A0(men_men_n1080_), .A1(men_men_n1067_), .B0(men_men_n68_), .Y(men_men_n1081_));
  NO2        u1059(.A(men_men_n1116_), .B(men_men_n793_), .Y(men_men_n1082_));
  OAI210     u1060(.A0(men_men_n75_), .A1(men_men_n52_), .B0(men_men_n106_), .Y(men_men_n1083_));
  NA2        u1061(.A(men_men_n1083_), .B(men_men_n71_), .Y(men_men_n1084_));
  AOI210     u1062(.A0(men_men_n1030_), .A1(men_men_n940_), .B0(men_men_n959_), .Y(men_men_n1085_));
  AOI210     u1063(.A0(men_men_n1085_), .A1(men_men_n1084_), .B0(men_men_n709_), .Y(men_men_n1086_));
  NA2        u1064(.A(men_men_n266_), .B(men_men_n54_), .Y(men_men_n1087_));
  AOI220     u1065(.A0(men_men_n1087_), .A1(men_men_n71_), .B0(men_men_n354_), .B1(men_men_n258_), .Y(men_men_n1088_));
  NO2        u1066(.A(men_men_n1088_), .B(men_men_n238_), .Y(men_men_n1089_));
  NA3        u1067(.A(men_men_n94_), .B(men_men_n312_), .C(men_men_n31_), .Y(men_men_n1090_));
  INV        u1068(.A(men_men_n1090_), .Y(men_men_n1091_));
  NO3        u1069(.A(men_men_n1091_), .B(men_men_n1089_), .C(men_men_n1086_), .Y(men_men_n1092_));
  OAI210     u1070(.A0(men_men_n272_), .A1(men_men_n158_), .B0(men_men_n84_), .Y(men_men_n1093_));
  NA3        u1071(.A(men_men_n797_), .B(men_men_n295_), .C(men_men_n75_), .Y(men_men_n1094_));
  AOI210     u1072(.A0(men_men_n1094_), .A1(men_men_n1093_), .B0(i_11_), .Y(men_men_n1095_));
  NA2        u1073(.A(men_men_n634_), .B(men_men_n215_), .Y(men_men_n1096_));
  OAI210     u1074(.A0(men_men_n1096_), .A1(men_men_n952_), .B0(men_men_n207_), .Y(men_men_n1097_));
  NA2        u1075(.A(men_men_n164_), .B(i_5_), .Y(men_men_n1098_));
  AOI210     u1076(.A0(men_men_n1097_), .A1(men_men_n809_), .B0(men_men_n1098_), .Y(men_men_n1099_));
  NO3        u1077(.A(men_men_n56_), .B(men_men_n55_), .C(i_4_), .Y(men_men_n1100_));
  OAI210     u1078(.A0(men_men_n963_), .A1(men_men_n312_), .B0(men_men_n1100_), .Y(men_men_n1101_));
  NO2        u1079(.A(men_men_n1101_), .B(men_men_n764_), .Y(men_men_n1102_));
  NO4        u1080(.A(men_men_n987_), .B(men_men_n488_), .C(men_men_n255_), .D(men_men_n254_), .Y(men_men_n1103_));
  NO2        u1081(.A(men_men_n1103_), .B(men_men_n586_), .Y(men_men_n1104_));
  NO2        u1082(.A(men_men_n850_), .B(men_men_n373_), .Y(men_men_n1105_));
  AOI210     u1083(.A0(men_men_n1105_), .A1(men_men_n1104_), .B0(men_men_n40_), .Y(men_men_n1106_));
  NO4        u1084(.A(men_men_n1106_), .B(men_men_n1102_), .C(men_men_n1099_), .D(men_men_n1095_), .Y(men_men_n1107_));
  OAI210     u1085(.A0(men_men_n1092_), .A1(i_4_), .B0(men_men_n1107_), .Y(men_men_n1108_));
  NO3        u1086(.A(men_men_n1108_), .B(men_men_n1082_), .C(men_men_n1081_), .Y(men_men_n1109_));
  NA4        u1087(.A(men_men_n1109_), .B(men_men_n1063_), .C(men_men_n994_), .D(men_men_n905_), .Y(men4));
  INV        u1088(.A(i_2_), .Y(men_men_n1113_));
  INV        u1089(.A(i_5_), .Y(men_men_n1114_));
  INV        u1090(.A(i_3_), .Y(men_men_n1115_));
  INV        u1091(.A(men_men_n589_), .Y(men_men_n1116_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule