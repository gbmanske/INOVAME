library verilog;
use verilog.vl_types.all;
entity tb_absolutesum is
end tb_absolutesum;
