library verilog;
use verilog.vl_types.all;
entity mult_vlg_vec_tst is
end mult_vlg_vec_tst;
