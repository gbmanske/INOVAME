library verilog;
use verilog.vl_types.all;
entity tb_signed_sum4inputs is
end tb_signed_sum4inputs;
