//Benchmark atmr_9sym_175_0.5

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m00(.A(i_6_), .Y(mai_mai_n11_));
  INV        m01(.A(i_5_), .Y(mai_mai_n12_));
  NOi21      m02(.An(i_3_), .B(i_7_), .Y(mai_mai_n13_));
  INV        m03(.A(i_0_), .Y(mai_mai_n14_));
  NOi21      m04(.An(i_1_), .B(i_3_), .Y(mai_mai_n15_));
  INV        m05(.A(i_7_), .Y(mai_mai_n16_));
  NA3        m06(.A(i_6_), .B(i_5_), .C(mai_mai_n16_), .Y(mai_mai_n17_));
  NA2        m07(.A(mai_mai_n14_), .B(i_5_), .Y(mai_mai_n18_));
  INV        m08(.A(i_2_), .Y(mai_mai_n19_));
  NOi21      m09(.An(i_5_), .B(i_0_), .Y(mai_mai_n20_));
  NOi21      m10(.An(i_6_), .B(i_8_), .Y(mai_mai_n21_));
  NOi21      m11(.An(i_7_), .B(i_1_), .Y(mai_mai_n22_));
  NOi21      m12(.An(i_5_), .B(i_6_), .Y(mai_mai_n23_));
  AOI220     m13(.A0(mai_mai_n23_), .A1(mai_mai_n22_), .B0(mai_mai_n21_), .B1(mai_mai_n20_), .Y(mai_mai_n24_));
  NO3        m14(.A(mai_mai_n24_), .B(mai_mai_n19_), .C(i_4_), .Y(mai_mai_n25_));
  NOi21      m15(.An(i_0_), .B(i_4_), .Y(mai_mai_n26_));
  XO2        m16(.A(i_1_), .B(i_3_), .Y(mai_mai_n27_));
  NOi21      m17(.An(i_7_), .B(i_5_), .Y(mai_mai_n28_));
  AN3        m18(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .Y(mai_mai_n29_));
  INV        m19(.A(i_1_), .Y(mai_mai_n30_));
  NOi21      m20(.An(i_3_), .B(i_0_), .Y(mai_mai_n31_));
  NA2        m21(.A(mai_mai_n31_), .B(mai_mai_n30_), .Y(mai_mai_n32_));
  NA3        m22(.A(i_6_), .B(mai_mai_n12_), .C(i_7_), .Y(mai_mai_n33_));
  AOI210     m23(.A0(mai_mai_n33_), .A1(mai_mai_n17_), .B0(mai_mai_n32_), .Y(mai_mai_n34_));
  NO3        m24(.A(mai_mai_n34_), .B(mai_mai_n29_), .C(mai_mai_n25_), .Y(mai_mai_n35_));
  INV        m25(.A(i_8_), .Y(mai_mai_n36_));
  NOi21      m26(.An(i_4_), .B(i_0_), .Y(mai_mai_n37_));
  NA2        m27(.A(i_1_), .B(mai_mai_n12_), .Y(mai_mai_n38_));
  NOi21      m28(.An(i_2_), .B(i_8_), .Y(mai_mai_n39_));
  NOi31      m29(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n40_));
  NA2        m30(.A(mai_mai_n40_), .B(i_0_), .Y(mai_mai_n41_));
  NOi21      m31(.An(i_4_), .B(i_3_), .Y(mai_mai_n42_));
  NOi21      m32(.An(i_1_), .B(i_4_), .Y(mai_mai_n43_));
  OAI210     m33(.A0(mai_mai_n43_), .A1(mai_mai_n42_), .B0(mai_mai_n39_), .Y(mai_mai_n44_));
  NA2        m34(.A(mai_mai_n44_), .B(mai_mai_n41_), .Y(mai_mai_n45_));
  AN2        m35(.A(i_8_), .B(i_7_), .Y(mai_mai_n46_));
  NA2        m36(.A(mai_mai_n46_), .B(mai_mai_n11_), .Y(mai_mai_n47_));
  NOi21      m37(.An(i_8_), .B(i_7_), .Y(mai_mai_n48_));
  NA3        m38(.A(mai_mai_n48_), .B(mai_mai_n42_), .C(i_6_), .Y(mai_mai_n49_));
  OAI210     m39(.A0(mai_mai_n47_), .A1(mai_mai_n38_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  AOI220     m40(.A0(mai_mai_n50_), .A1(mai_mai_n19_), .B0(mai_mai_n45_), .B1(mai_mai_n23_), .Y(mai_mai_n51_));
  NA2        m41(.A(mai_mai_n51_), .B(mai_mai_n35_), .Y(mai_mai_n52_));
  NA2        m42(.A(i_8_), .B(mai_mai_n16_), .Y(mai_mai_n53_));
  AOI220     m43(.A0(mai_mai_n31_), .A1(i_1_), .B0(mai_mai_n27_), .B1(i_2_), .Y(mai_mai_n54_));
  NOi21      m44(.An(i_1_), .B(i_2_), .Y(mai_mai_n55_));
  NO2        m45(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n56_));
  NA2        m46(.A(mai_mai_n56_), .B(mai_mai_n12_), .Y(mai_mai_n57_));
  NA3        m47(.A(mai_mai_n48_), .B(i_2_), .C(mai_mai_n11_), .Y(mai_mai_n58_));
  INV        m48(.A(mai_mai_n57_), .Y(mai_mai_n59_));
  NAi21      m49(.An(i_3_), .B(i_6_), .Y(mai_mai_n60_));
  NO3        m50(.A(mai_mai_n60_), .B(i_0_), .C(mai_mai_n36_), .Y(mai_mai_n61_));
  NA2        m51(.A(mai_mai_n21_), .B(mai_mai_n20_), .Y(mai_mai_n62_));
  NOi21      m52(.An(i_7_), .B(i_8_), .Y(mai_mai_n63_));
  INV        m53(.A(mai_mai_n62_), .Y(mai_mai_n64_));
  OAI210     m54(.A0(mai_mai_n64_), .A1(mai_mai_n61_), .B0(mai_mai_n55_), .Y(mai_mai_n65_));
  NA3        m55(.A(mai_mai_n48_), .B(mai_mai_n19_), .C(i_3_), .Y(mai_mai_n66_));
  NAi21      m56(.An(i_6_), .B(i_0_), .Y(mai_mai_n67_));
  NA3        m57(.A(mai_mai_n43_), .B(i_5_), .C(mai_mai_n16_), .Y(mai_mai_n68_));
  NOi21      m58(.An(i_4_), .B(i_6_), .Y(mai_mai_n69_));
  NOi21      m59(.An(i_5_), .B(i_3_), .Y(mai_mai_n70_));
  NA3        m60(.A(mai_mai_n70_), .B(mai_mai_n55_), .C(mai_mai_n69_), .Y(mai_mai_n71_));
  OAI210     m61(.A0(mai_mai_n68_), .A1(mai_mai_n67_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  NA2        m62(.A(mai_mai_n55_), .B(mai_mai_n21_), .Y(mai_mai_n73_));
  NOi21      m63(.An(mai_mai_n28_), .B(mai_mai_n73_), .Y(mai_mai_n74_));
  NO2        m64(.A(mai_mai_n74_), .B(mai_mai_n72_), .Y(mai_mai_n75_));
  NA2        m65(.A(mai_mai_n75_), .B(mai_mai_n65_), .Y(mai_mai_n76_));
  NOi31      m66(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n77_));
  NA2        m67(.A(mai_mai_n77_), .B(i_7_), .Y(mai_mai_n78_));
  NA2        m68(.A(mai_mai_n78_), .B(mai_mai_n73_), .Y(mai_mai_n79_));
  NA2        m69(.A(mai_mai_n79_), .B(mai_mai_n26_), .Y(mai_mai_n80_));
  NA2        m70(.A(mai_mai_n42_), .B(mai_mai_n22_), .Y(mai_mai_n81_));
  AOI210     m71(.A0(mai_mai_n81_), .A1(mai_mai_n58_), .B0(mai_mai_n18_), .Y(mai_mai_n82_));
  NA3        m72(.A(mai_mai_n48_), .B(mai_mai_n40_), .C(i_6_), .Y(mai_mai_n83_));
  INV        m73(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  NOi21      m74(.An(i_0_), .B(i_2_), .Y(mai_mai_n85_));
  NA3        m75(.A(mai_mai_n85_), .B(mai_mai_n22_), .C(mai_mai_n69_), .Y(mai_mai_n86_));
  NA3        m76(.A(mai_mai_n37_), .B(mai_mai_n28_), .C(mai_mai_n15_), .Y(mai_mai_n87_));
  NA3        m77(.A(mai_mai_n85_), .B(mai_mai_n42_), .C(mai_mai_n21_), .Y(mai_mai_n88_));
  NA3        m78(.A(mai_mai_n88_), .B(mai_mai_n87_), .C(mai_mai_n86_), .Y(mai_mai_n89_));
  NA4        m79(.A(mai_mai_n40_), .B(i_6_), .C(mai_mai_n12_), .D(i_7_), .Y(mai_mai_n90_));
  NA4        m80(.A(mai_mai_n43_), .B(mai_mai_n23_), .C(mai_mai_n14_), .D(i_8_), .Y(mai_mai_n91_));
  NA2        m81(.A(mai_mai_n91_), .B(mai_mai_n90_), .Y(mai_mai_n92_));
  NO4        m82(.A(mai_mai_n92_), .B(mai_mai_n89_), .C(mai_mai_n84_), .D(mai_mai_n82_), .Y(mai_mai_n93_));
  NA2        m83(.A(mai_mai_n63_), .B(mai_mai_n11_), .Y(mai_mai_n94_));
  NA3        m84(.A(i_2_), .B(i_1_), .C(mai_mai_n12_), .Y(mai_mai_n95_));
  NA2        m85(.A(mai_mai_n37_), .B(i_3_), .Y(mai_mai_n96_));
  AOI210     m86(.A0(mai_mai_n96_), .A1(mai_mai_n95_), .B0(mai_mai_n94_), .Y(mai_mai_n97_));
  NA3        m87(.A(mai_mai_n85_), .B(mai_mai_n48_), .C(mai_mai_n69_), .Y(mai_mai_n98_));
  OAI210     m88(.A0(mai_mai_n66_), .A1(mai_mai_n18_), .B0(mai_mai_n98_), .Y(mai_mai_n99_));
  NA3        m89(.A(mai_mai_n39_), .B(mai_mai_n20_), .C(mai_mai_n13_), .Y(mai_mai_n100_));
  INV        m90(.A(mai_mai_n100_), .Y(mai_mai_n101_));
  NO3        m91(.A(mai_mai_n101_), .B(mai_mai_n99_), .C(mai_mai_n97_), .Y(mai_mai_n102_));
  NA3        m92(.A(mai_mai_n102_), .B(mai_mai_n93_), .C(mai_mai_n80_), .Y(mai_mai_n103_));
  OR4        m93(.A(mai_mai_n103_), .B(mai_mai_n76_), .C(mai_mai_n59_), .D(mai_mai_n52_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NA3        u013(.A(i_6_), .B(i_5_), .C(men_men_n23_), .Y(men_men_n24_));
  NOi21      u014(.An(i_8_), .B(i_6_), .Y(men_men_n25_));
  NOi21      u015(.An(i_1_), .B(i_8_), .Y(men_men_n26_));
  AOI220     u016(.A0(men_men_n26_), .A1(i_2_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n22_), .Y(men_men_n28_));
  AOI210     u018(.A0(men_men_n28_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n29_));
  NA2        u019(.A(i_0_), .B(men_men_n14_), .Y(men_men_n30_));
  NA2        u020(.A(men_men_n17_), .B(i_5_), .Y(men_men_n31_));
  NO2        u021(.A(i_2_), .B(i_4_), .Y(men_men_n32_));
  NA3        u022(.A(men_men_n32_), .B(i_6_), .C(i_8_), .Y(men_men_n33_));
  AOI210     u023(.A0(men_men_n31_), .A1(men_men_n30_), .B0(men_men_n33_), .Y(men_men_n34_));
  INV        u024(.A(i_2_), .Y(men_men_n35_));
  NOi21      u025(.An(i_6_), .B(i_8_), .Y(men_men_n36_));
  NOi21      u026(.An(i_0_), .B(i_4_), .Y(men_men_n37_));
  INV        u027(.A(i_1_), .Y(men_men_n38_));
  NOi21      u028(.An(i_3_), .B(i_0_), .Y(men_men_n39_));
  INV        u029(.A(men_men_n34_), .Y(men_men_n40_));
  INV        u030(.A(i_8_), .Y(men_men_n41_));
  NA2        u031(.A(i_1_), .B(men_men_n11_), .Y(men_men_n42_));
  NO4        u032(.A(men_men_n42_), .B(men_men_n30_), .C(i_2_), .D(men_men_n41_), .Y(men_men_n43_));
  NOi21      u033(.An(i_4_), .B(i_0_), .Y(men_men_n44_));
  AOI210     u034(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n15_), .Y(men_men_n45_));
  NA2        u035(.A(i_1_), .B(men_men_n14_), .Y(men_men_n46_));
  NOi21      u036(.An(i_2_), .B(i_8_), .Y(men_men_n47_));
  NO3        u037(.A(men_men_n47_), .B(men_men_n44_), .C(men_men_n37_), .Y(men_men_n48_));
  NO3        u038(.A(men_men_n48_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n49_));
  NO2        u039(.A(men_men_n49_), .B(men_men_n43_), .Y(men_men_n50_));
  NOi21      u040(.An(i_4_), .B(i_3_), .Y(men_men_n51_));
  NOi21      u041(.An(i_1_), .B(i_4_), .Y(men_men_n52_));
  AN2        u042(.A(i_8_), .B(i_7_), .Y(men_men_n53_));
  NOi21      u043(.An(i_8_), .B(i_7_), .Y(men_men_n54_));
  NA3        u044(.A(men_men_n50_), .B(men_men_n40_), .C(men_men_n29_), .Y(men_men_n55_));
  NA2        u045(.A(i_8_), .B(i_7_), .Y(men_men_n56_));
  NO3        u046(.A(men_men_n56_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n57_));
  NOi21      u047(.An(i_1_), .B(i_2_), .Y(men_men_n58_));
  NA3        u048(.A(men_men_n58_), .B(men_men_n44_), .C(i_6_), .Y(men_men_n59_));
  INV        u049(.A(men_men_n59_), .Y(men_men_n60_));
  OAI210     u050(.A0(men_men_n60_), .A1(men_men_n57_), .B0(men_men_n14_), .Y(men_men_n61_));
  NA3        u051(.A(men_men_n54_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n26_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n63_));
  NA2        u053(.A(men_men_n63_), .B(men_men_n62_), .Y(men_men_n64_));
  NOi32      u054(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(i_3_), .Y(men_men_n66_));
  NA3        u056(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n67_));
  NA2        u057(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n68_));
  NO2        u058(.A(i_0_), .B(i_4_), .Y(men_men_n69_));
  AOI220     u059(.A0(men_men_n69_), .A1(men_men_n68_), .B0(men_men_n64_), .B1(men_men_n51_), .Y(men_men_n70_));
  NA2        u060(.A(men_men_n70_), .B(men_men_n61_), .Y(men_men_n71_));
  NAi21      u061(.An(i_3_), .B(i_6_), .Y(men_men_n72_));
  NOi21      u062(.An(i_7_), .B(i_8_), .Y(men_men_n73_));
  NOi31      u063(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n74_));
  AOI210     u064(.A0(men_men_n73_), .A1(men_men_n12_), .B0(men_men_n74_), .Y(men_men_n75_));
  NO2        u065(.A(men_men_n75_), .B(men_men_n11_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n76_), .B(men_men_n58_), .Y(men_men_n77_));
  NA3        u067(.A(men_men_n25_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n78_));
  AOI210     u068(.A0(men_men_n22_), .A1(men_men_n42_), .B0(men_men_n78_), .Y(men_men_n79_));
  AOI220     u069(.A0(men_men_n39_), .A1(men_men_n38_), .B0(men_men_n18_), .B1(men_men_n35_), .Y(men_men_n80_));
  NA3        u070(.A(men_men_n21_), .B(i_5_), .C(i_7_), .Y(men_men_n81_));
  OAI210     u071(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n82_));
  NA3        u072(.A(men_men_n56_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n83_));
  OAI220     u073(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n84_));
  NO2        u074(.A(men_men_n84_), .B(men_men_n79_), .Y(men_men_n85_));
  NA3        u075(.A(men_men_n54_), .B(men_men_n35_), .C(i_3_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n38_), .B(i_6_), .Y(men_men_n87_));
  AOI210     u077(.A0(men_men_n87_), .A1(men_men_n22_), .B0(men_men_n86_), .Y(men_men_n88_));
  NOi21      u078(.An(i_2_), .B(i_1_), .Y(men_men_n89_));
  AN3        u079(.A(men_men_n73_), .B(men_men_n89_), .C(men_men_n44_), .Y(men_men_n90_));
  NAi21      u080(.An(i_6_), .B(i_0_), .Y(men_men_n91_));
  NOi21      u081(.An(i_4_), .B(i_6_), .Y(men_men_n92_));
  NOi21      u082(.An(i_5_), .B(i_3_), .Y(men_men_n93_));
  NO2        u083(.A(men_men_n90_), .B(men_men_n88_), .Y(men_men_n94_));
  NOi21      u084(.An(i_6_), .B(i_1_), .Y(men_men_n95_));
  AOI220     u085(.A0(men_men_n95_), .A1(i_7_), .B0(men_men_n25_), .B1(i_5_), .Y(men_men_n96_));
  NOi31      u086(.An(men_men_n44_), .B(men_men_n96_), .C(i_2_), .Y(men_men_n97_));
  NA2        u087(.A(men_men_n54_), .B(men_men_n12_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n36_), .B(men_men_n14_), .Y(men_men_n99_));
  NOi21      u089(.An(i_3_), .B(i_1_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n100_), .B(i_4_), .Y(men_men_n101_));
  AOI210     u091(.A0(men_men_n99_), .A1(men_men_n98_), .B0(men_men_n101_), .Y(men_men_n102_));
  AOI220     u092(.A0(men_men_n73_), .A1(men_men_n14_), .B0(men_men_n92_), .B1(men_men_n23_), .Y(men_men_n103_));
  NOi31      u093(.An(men_men_n39_), .B(men_men_n103_), .C(men_men_n35_), .Y(men_men_n104_));
  NO3        u094(.A(men_men_n104_), .B(men_men_n102_), .C(men_men_n97_), .Y(men_men_n105_));
  NA4        u095(.A(men_men_n105_), .B(men_men_n94_), .C(men_men_n85_), .D(men_men_n77_), .Y(men_men_n106_));
  NA2        u096(.A(men_men_n47_), .B(men_men_n15_), .Y(men_men_n107_));
  NOi31      u097(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n108_));
  NA2        u098(.A(men_men_n108_), .B(i_7_), .Y(men_men_n109_));
  NA3        u099(.A(men_men_n36_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n110_));
  NA3        u100(.A(men_men_n110_), .B(men_men_n109_), .C(men_men_n107_), .Y(men_men_n111_));
  NA2        u101(.A(men_men_n111_), .B(men_men_n37_), .Y(men_men_n112_));
  NA4        u102(.A(men_men_n53_), .B(men_men_n89_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n113_));
  NAi31      u103(.An(men_men_n91_), .B(men_men_n73_), .C(men_men_n89_), .Y(men_men_n114_));
  NA2        u104(.A(men_men_n114_), .B(men_men_n113_), .Y(men_men_n115_));
  NOi32      u105(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n116_), .B(men_men_n108_), .Y(men_men_n117_));
  INV        u107(.A(men_men_n117_), .Y(men_men_n118_));
  NA4        u108(.A(men_men_n52_), .B(men_men_n39_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n119_));
  INV        u109(.A(men_men_n119_), .Y(men_men_n120_));
  NO3        u110(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n115_), .Y(men_men_n121_));
  NOi21      u111(.An(i_5_), .B(i_2_), .Y(men_men_n122_));
  AOI220     u112(.A0(men_men_n122_), .A1(men_men_n73_), .B0(men_men_n53_), .B1(men_men_n32_), .Y(men_men_n123_));
  AOI210     u113(.A0(men_men_n123_), .A1(men_men_n107_), .B0(men_men_n87_), .Y(men_men_n124_));
  NO4        u114(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n125_));
  NA2        u115(.A(i_2_), .B(i_4_), .Y(men_men_n126_));
  AOI210     u116(.A0(men_men_n91_), .A1(men_men_n72_), .B0(men_men_n126_), .Y(men_men_n127_));
  NO2        u117(.A(i_8_), .B(i_7_), .Y(men_men_n128_));
  OA210      u118(.A0(men_men_n127_), .A1(men_men_n125_), .B0(men_men_n128_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n100_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n130_));
  NO2        u120(.A(men_men_n130_), .B(i_4_), .Y(men_men_n131_));
  NO3        u121(.A(men_men_n131_), .B(men_men_n129_), .C(men_men_n124_), .Y(men_men_n132_));
  NA4        u122(.A(men_men_n93_), .B(men_men_n53_), .C(men_men_n38_), .D(men_men_n21_), .Y(men_men_n133_));
  NA3        u123(.A(men_men_n74_), .B(men_men_n100_), .C(i_0_), .Y(men_men_n134_));
  NOi31      u124(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n135_));
  OAI210     u125(.A0(men_men_n116_), .A1(men_men_n65_), .B0(men_men_n135_), .Y(men_men_n136_));
  NA3        u126(.A(men_men_n136_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n137_));
  INV        u127(.A(men_men_n137_), .Y(men_men_n138_));
  NA4        u128(.A(men_men_n138_), .B(men_men_n132_), .C(men_men_n121_), .D(men_men_n112_), .Y(men_men_n139_));
  OR4        u129(.A(men_men_n139_), .B(men_men_n106_), .C(men_men_n71_), .D(men_men_n55_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule