//Benchmark atmr_9sym_175_0.25

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_1_), .B(i_8_), .Y(mai_mai_n25_));
  NA2        m015(.A(mai_mai_n25_), .B(i_2_), .Y(mai_mai_n26_));
  AOI210     m016(.A0(mai_mai_n26_), .A1(mai_mai_n24_), .B0(mai_mai_n22_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n28_));
  NA2        m018(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n29_));
  INV        m019(.A(i_2_), .Y(mai_mai_n30_));
  NOi21      m020(.An(i_5_), .B(i_0_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_6_), .B(i_8_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_7_), .B(i_1_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_5_), .B(i_6_), .Y(mai_mai_n34_));
  AOI220     m024(.A0(mai_mai_n34_), .A1(mai_mai_n33_), .B0(mai_mai_n32_), .B1(mai_mai_n31_), .Y(mai_mai_n35_));
  NO3        m025(.A(mai_mai_n35_), .B(mai_mai_n30_), .C(i_4_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_0_), .B(i_4_), .Y(mai_mai_n37_));
  XO2        m027(.A(i_1_), .B(i_3_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_7_), .B(i_5_), .Y(mai_mai_n39_));
  AN3        m029(.A(mai_mai_n39_), .B(mai_mai_n38_), .C(mai_mai_n37_), .Y(mai_mai_n40_));
  INV        m030(.A(i_1_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_3_), .B(i_0_), .Y(mai_mai_n42_));
  NA2        m032(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA3        m033(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n44_));
  AOI210     m034(.A0(mai_mai_n44_), .A1(mai_mai_n24_), .B0(mai_mai_n43_), .Y(mai_mai_n45_));
  NO3        m035(.A(mai_mai_n45_), .B(mai_mai_n40_), .C(mai_mai_n36_), .Y(mai_mai_n46_));
  NOi21      m036(.An(i_4_), .B(i_0_), .Y(mai_mai_n47_));
  NA2        m037(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n48_));
  NOi21      m038(.An(i_2_), .B(i_8_), .Y(mai_mai_n49_));
  NOi31      m039(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n50_));
  NA2        m040(.A(mai_mai_n50_), .B(i_0_), .Y(mai_mai_n51_));
  NOi21      m041(.An(i_4_), .B(i_3_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_1_), .B(i_4_), .Y(mai_mai_n53_));
  OAI210     m043(.A0(mai_mai_n53_), .A1(mai_mai_n52_), .B0(mai_mai_n49_), .Y(mai_mai_n54_));
  NA2        m044(.A(mai_mai_n54_), .B(mai_mai_n51_), .Y(mai_mai_n55_));
  AN2        m045(.A(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  NA2        m046(.A(mai_mai_n56_), .B(mai_mai_n12_), .Y(mai_mai_n57_));
  NOi21      m047(.An(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  NA3        m048(.A(mai_mai_n58_), .B(mai_mai_n52_), .C(i_6_), .Y(mai_mai_n59_));
  OAI210     m049(.A0(mai_mai_n57_), .A1(mai_mai_n48_), .B0(mai_mai_n59_), .Y(mai_mai_n60_));
  AOI220     m050(.A0(mai_mai_n60_), .A1(mai_mai_n30_), .B0(mai_mai_n55_), .B1(mai_mai_n34_), .Y(mai_mai_n61_));
  NA3        m051(.A(mai_mai_n61_), .B(mai_mai_n46_), .C(mai_mai_n28_), .Y(mai_mai_n62_));
  NA2        m052(.A(i_8_), .B(i_7_), .Y(mai_mai_n63_));
  NO3        m053(.A(mai_mai_n63_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n64_));
  NA2        m054(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n65_));
  AOI220     m055(.A0(mai_mai_n42_), .A1(i_1_), .B0(mai_mai_n38_), .B1(i_2_), .Y(mai_mai_n66_));
  NOi21      m056(.An(i_1_), .B(i_2_), .Y(mai_mai_n67_));
  NO2        m057(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n68_));
  OAI210     m058(.A0(mai_mai_n68_), .A1(mai_mai_n64_), .B0(mai_mai_n14_), .Y(mai_mai_n69_));
  NA3        m059(.A(mai_mai_n58_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n70_));
  NA3        m060(.A(mai_mai_n25_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n71_));
  NA2        m061(.A(mai_mai_n71_), .B(mai_mai_n70_), .Y(mai_mai_n72_));
  NA2        m062(.A(mai_mai_n72_), .B(mai_mai_n52_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n73_), .B(mai_mai_n69_), .Y(mai_mai_n74_));
  NA2        m064(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n75_));
  NOi21      m065(.An(i_7_), .B(i_8_), .Y(mai_mai_n76_));
  NA2        m066(.A(mai_mai_n76_), .B(mai_mai_n12_), .Y(mai_mai_n77_));
  OAI210     m067(.A0(mai_mai_n77_), .A1(mai_mai_n11_), .B0(mai_mai_n75_), .Y(mai_mai_n78_));
  NA2        m068(.A(mai_mai_n78_), .B(mai_mai_n67_), .Y(mai_mai_n79_));
  AOI220     m069(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n18_), .B1(mai_mai_n30_), .Y(mai_mai_n80_));
  NA3        m070(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n81_));
  NO2        m071(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  INV        m072(.A(mai_mai_n82_), .Y(mai_mai_n83_));
  NA3        m073(.A(mai_mai_n58_), .B(mai_mai_n30_), .C(i_3_), .Y(mai_mai_n84_));
  NO2        m074(.A(mai_mai_n22_), .B(mai_mai_n84_), .Y(mai_mai_n85_));
  NAi21      m075(.An(i_6_), .B(i_0_), .Y(mai_mai_n86_));
  NA3        m076(.A(mai_mai_n53_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_4_), .B(i_6_), .Y(mai_mai_n88_));
  NOi21      m078(.An(i_5_), .B(i_3_), .Y(mai_mai_n89_));
  NA3        m079(.A(mai_mai_n89_), .B(mai_mai_n67_), .C(mai_mai_n88_), .Y(mai_mai_n90_));
  OAI210     m080(.A0(mai_mai_n87_), .A1(mai_mai_n86_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  NA2        m081(.A(mai_mai_n67_), .B(mai_mai_n32_), .Y(mai_mai_n92_));
  NOi21      m082(.An(mai_mai_n39_), .B(mai_mai_n92_), .Y(mai_mai_n93_));
  NO3        m083(.A(mai_mai_n93_), .B(mai_mai_n91_), .C(mai_mai_n85_), .Y(mai_mai_n94_));
  NA2        m084(.A(mai_mai_n58_), .B(mai_mai_n12_), .Y(mai_mai_n95_));
  NA2        m085(.A(mai_mai_n32_), .B(mai_mai_n14_), .Y(mai_mai_n96_));
  NOi21      m086(.An(i_3_), .B(i_1_), .Y(mai_mai_n97_));
  NA2        m087(.A(mai_mai_n97_), .B(i_4_), .Y(mai_mai_n98_));
  AOI210     m088(.A0(mai_mai_n96_), .A1(mai_mai_n95_), .B0(mai_mai_n98_), .Y(mai_mai_n99_));
  INV        m089(.A(mai_mai_n99_), .Y(mai_mai_n100_));
  NA4        m090(.A(mai_mai_n100_), .B(mai_mai_n94_), .C(mai_mai_n83_), .D(mai_mai_n79_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n49_), .B(mai_mai_n15_), .Y(mai_mai_n102_));
  NA2        m092(.A(mai_mai_n102_), .B(mai_mai_n92_), .Y(mai_mai_n103_));
  NA2        m093(.A(mai_mai_n103_), .B(mai_mai_n37_), .Y(mai_mai_n104_));
  NA2        m094(.A(mai_mai_n52_), .B(mai_mai_n33_), .Y(mai_mai_n105_));
  AOI210     m095(.A0(mai_mai_n105_), .A1(mai_mai_n70_), .B0(mai_mai_n29_), .Y(mai_mai_n106_));
  NA3        m096(.A(mai_mai_n58_), .B(mai_mai_n50_), .C(i_6_), .Y(mai_mai_n107_));
  INV        m097(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NOi21      m098(.An(i_0_), .B(i_2_), .Y(mai_mai_n109_));
  NA3        m099(.A(mai_mai_n109_), .B(mai_mai_n33_), .C(mai_mai_n88_), .Y(mai_mai_n110_));
  NA3        m100(.A(mai_mai_n47_), .B(mai_mai_n39_), .C(mai_mai_n18_), .Y(mai_mai_n111_));
  NA3        m101(.A(mai_mai_n109_), .B(mai_mai_n52_), .C(mai_mai_n32_), .Y(mai_mai_n112_));
  NA3        m102(.A(mai_mai_n112_), .B(mai_mai_n111_), .C(mai_mai_n110_), .Y(mai_mai_n113_));
  NA4        m103(.A(mai_mai_n50_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n114_));
  INV        m104(.A(mai_mai_n114_), .Y(mai_mai_n115_));
  NO4        m105(.A(mai_mai_n115_), .B(mai_mai_n113_), .C(mai_mai_n108_), .D(mai_mai_n106_), .Y(mai_mai_n116_));
  NA2        m106(.A(mai_mai_n76_), .B(mai_mai_n12_), .Y(mai_mai_n117_));
  NA3        m107(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n118_));
  NA2        m108(.A(mai_mai_n47_), .B(i_3_), .Y(mai_mai_n119_));
  AOI210     m109(.A0(mai_mai_n119_), .A1(mai_mai_n118_), .B0(mai_mai_n117_), .Y(mai_mai_n120_));
  NO2        m110(.A(mai_mai_n84_), .B(mai_mai_n29_), .Y(mai_mai_n121_));
  NA4        m111(.A(mai_mai_n89_), .B(mai_mai_n56_), .C(mai_mai_n41_), .D(mai_mai_n21_), .Y(mai_mai_n122_));
  NA3        m112(.A(mai_mai_n49_), .B(mai_mai_n31_), .C(mai_mai_n15_), .Y(mai_mai_n123_));
  NA2        m113(.A(mai_mai_n123_), .B(mai_mai_n122_), .Y(mai_mai_n124_));
  NO3        m114(.A(mai_mai_n124_), .B(mai_mai_n121_), .C(mai_mai_n120_), .Y(mai_mai_n125_));
  NA3        m115(.A(mai_mai_n125_), .B(mai_mai_n116_), .C(mai_mai_n104_), .Y(mai_mai_n126_));
  OR4        m116(.A(mai_mai_n126_), .B(mai_mai_n101_), .C(mai_mai_n74_), .D(mai_mai_n62_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  INV        u002(.A(i_5_), .Y(men_men_n13_));
  NOi21      u003(.An(i_3_), .B(i_7_), .Y(men_men_n14_));
  INV        u004(.A(i_0_), .Y(men_men_n15_));
  NOi21      u005(.An(i_1_), .B(i_3_), .Y(men_men_n16_));
  INV        u006(.A(i_4_), .Y(men_men_n17_));
  NA2        u007(.A(i_0_), .B(men_men_n17_), .Y(men_men_n18_));
  INV        u008(.A(i_7_), .Y(men_men_n19_));
  NA3        u009(.A(i_6_), .B(i_5_), .C(men_men_n19_), .Y(men_men_n20_));
  NOi21      u010(.An(i_8_), .B(i_6_), .Y(men_men_n21_));
  NA2        u011(.A(men_men_n21_), .B(i_5_), .Y(men_men_n22_));
  AOI210     u012(.A0(men_men_n22_), .A1(men_men_n20_), .B0(men_men_n18_), .Y(men_men_n23_));
  NA2        u013(.A(men_men_n23_), .B(men_men_n11_), .Y(men_men_n24_));
  NA2        u014(.A(i_0_), .B(men_men_n13_), .Y(men_men_n25_));
  NA2        u015(.A(men_men_n15_), .B(i_5_), .Y(men_men_n26_));
  NO2        u016(.A(i_2_), .B(i_4_), .Y(men_men_n27_));
  NA3        u017(.A(men_men_n27_), .B(i_6_), .C(i_8_), .Y(men_men_n28_));
  AOI210     u018(.A0(men_men_n26_), .A1(men_men_n25_), .B0(men_men_n28_), .Y(men_men_n29_));
  INV        u019(.A(i_2_), .Y(men_men_n30_));
  NOi21      u020(.An(i_6_), .B(i_8_), .Y(men_men_n31_));
  NOi21      u021(.An(i_5_), .B(i_6_), .Y(men_men_n32_));
  NOi21      u022(.An(i_0_), .B(i_4_), .Y(men_men_n33_));
  INV        u023(.A(i_1_), .Y(men_men_n34_));
  NOi21      u024(.An(i_3_), .B(i_0_), .Y(men_men_n35_));
  INV        u025(.A(men_men_n29_), .Y(men_men_n36_));
  INV        u026(.A(i_8_), .Y(men_men_n37_));
  NA2        u027(.A(i_1_), .B(men_men_n11_), .Y(men_men_n38_));
  NO4        u028(.A(men_men_n38_), .B(men_men_n25_), .C(i_2_), .D(men_men_n37_), .Y(men_men_n39_));
  NOi21      u029(.An(i_4_), .B(i_0_), .Y(men_men_n40_));
  AOI210     u030(.A0(men_men_n40_), .A1(men_men_n21_), .B0(men_men_n14_), .Y(men_men_n41_));
  NA2        u031(.A(i_1_), .B(men_men_n13_), .Y(men_men_n42_));
  NOi21      u032(.An(i_2_), .B(i_8_), .Y(men_men_n43_));
  NO3        u033(.A(men_men_n43_), .B(men_men_n40_), .C(men_men_n33_), .Y(men_men_n44_));
  NO3        u034(.A(men_men_n44_), .B(men_men_n42_), .C(men_men_n41_), .Y(men_men_n45_));
  NO2        u035(.A(men_men_n45_), .B(men_men_n39_), .Y(men_men_n46_));
  NOi21      u036(.An(i_1_), .B(i_4_), .Y(men_men_n47_));
  AN2        u037(.A(i_8_), .B(i_7_), .Y(men_men_n48_));
  NOi21      u038(.An(i_8_), .B(i_7_), .Y(men_men_n49_));
  NA3        u039(.A(men_men_n46_), .B(men_men_n36_), .C(men_men_n24_), .Y(men_men_n50_));
  NA2        u040(.A(i_8_), .B(i_7_), .Y(men_men_n51_));
  NOi21      u041(.An(i_1_), .B(i_2_), .Y(men_men_n52_));
  NA3        u042(.A(men_men_n52_), .B(men_men_n40_), .C(i_6_), .Y(men_men_n53_));
  INV        u043(.A(men_men_n53_), .Y(men_men_n54_));
  NA2        u044(.A(men_men_n54_), .B(men_men_n13_), .Y(men_men_n55_));
  NOi32      u045(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n56_));
  NA2        u046(.A(men_men_n56_), .B(i_3_), .Y(men_men_n57_));
  NA3        u047(.A(men_men_n16_), .B(i_2_), .C(i_6_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(men_men_n57_), .Y(men_men_n59_));
  NO2        u049(.A(i_0_), .B(i_4_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(men_men_n59_), .Y(men_men_n61_));
  NA2        u051(.A(men_men_n61_), .B(men_men_n55_), .Y(men_men_n62_));
  NAi21      u052(.An(i_3_), .B(i_6_), .Y(men_men_n63_));
  NO3        u053(.A(men_men_n63_), .B(i_0_), .C(men_men_n37_), .Y(men_men_n64_));
  NOi21      u054(.An(i_7_), .B(i_8_), .Y(men_men_n65_));
  NOi31      u055(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n66_));
  AOI210     u056(.A0(men_men_n65_), .A1(men_men_n12_), .B0(men_men_n66_), .Y(men_men_n67_));
  NO2        u057(.A(men_men_n67_), .B(men_men_n11_), .Y(men_men_n68_));
  OAI210     u058(.A0(men_men_n68_), .A1(men_men_n64_), .B0(men_men_n52_), .Y(men_men_n69_));
  NA3        u059(.A(men_men_n21_), .B(i_2_), .C(men_men_n13_), .Y(men_men_n70_));
  AOI210     u060(.A0(men_men_n18_), .A1(men_men_n38_), .B0(men_men_n70_), .Y(men_men_n71_));
  OAI210     u061(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n72_));
  NA3        u062(.A(men_men_n51_), .B(men_men_n16_), .C(men_men_n15_), .Y(men_men_n73_));
  NO2        u063(.A(men_men_n73_), .B(men_men_n72_), .Y(men_men_n74_));
  NO2        u064(.A(men_men_n74_), .B(men_men_n71_), .Y(men_men_n75_));
  NA3        u065(.A(men_men_n49_), .B(men_men_n30_), .C(i_3_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n34_), .B(i_6_), .Y(men_men_n77_));
  AOI210     u067(.A0(men_men_n77_), .A1(men_men_n18_), .B0(men_men_n76_), .Y(men_men_n78_));
  NOi21      u068(.An(i_2_), .B(i_1_), .Y(men_men_n79_));
  AN3        u069(.A(men_men_n65_), .B(men_men_n79_), .C(men_men_n40_), .Y(men_men_n80_));
  NAi21      u070(.An(i_6_), .B(i_0_), .Y(men_men_n81_));
  NOi21      u071(.An(i_4_), .B(i_6_), .Y(men_men_n82_));
  NA2        u072(.A(men_men_n52_), .B(men_men_n31_), .Y(men_men_n83_));
  NO2        u073(.A(men_men_n80_), .B(men_men_n78_), .Y(men_men_n84_));
  NOi21      u074(.An(i_6_), .B(i_1_), .Y(men_men_n85_));
  AOI220     u075(.A0(men_men_n85_), .A1(i_7_), .B0(men_men_n21_), .B1(i_5_), .Y(men_men_n86_));
  NOi31      u076(.An(men_men_n40_), .B(men_men_n86_), .C(i_2_), .Y(men_men_n87_));
  NOi21      u077(.An(i_3_), .B(i_1_), .Y(men_men_n88_));
  AOI220     u078(.A0(men_men_n65_), .A1(men_men_n13_), .B0(men_men_n82_), .B1(men_men_n19_), .Y(men_men_n89_));
  NOi31      u079(.An(men_men_n35_), .B(men_men_n89_), .C(men_men_n30_), .Y(men_men_n90_));
  NO2        u080(.A(men_men_n90_), .B(men_men_n87_), .Y(men_men_n91_));
  NA4        u081(.A(men_men_n91_), .B(men_men_n84_), .C(men_men_n75_), .D(men_men_n69_), .Y(men_men_n92_));
  NA2        u082(.A(men_men_n43_), .B(men_men_n14_), .Y(men_men_n93_));
  NOi31      u083(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n94_));
  NOi31      u084(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n95_));
  OAI210     u085(.A0(men_men_n95_), .A1(men_men_n94_), .B0(i_7_), .Y(men_men_n96_));
  NA3        u086(.A(men_men_n31_), .B(i_2_), .C(men_men_n13_), .Y(men_men_n97_));
  NA4        u087(.A(men_men_n97_), .B(men_men_n96_), .C(men_men_n93_), .D(men_men_n83_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n98_), .B(men_men_n33_), .Y(men_men_n99_));
  NA4        u089(.A(men_men_n48_), .B(men_men_n79_), .C(men_men_n15_), .D(men_men_n12_), .Y(men_men_n100_));
  NAi31      u090(.An(men_men_n81_), .B(men_men_n65_), .C(men_men_n79_), .Y(men_men_n101_));
  NA2        u091(.A(men_men_n101_), .B(men_men_n100_), .Y(men_men_n102_));
  NOi21      u092(.An(i_0_), .B(i_2_), .Y(men_men_n103_));
  NOi32      u093(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n104_), .B(men_men_n94_), .Y(men_men_n105_));
  INV        u095(.A(men_men_n105_), .Y(men_men_n106_));
  NA4        u096(.A(men_men_n47_), .B(men_men_n32_), .C(men_men_n15_), .D(i_8_), .Y(men_men_n107_));
  NA4        u097(.A(men_men_n47_), .B(men_men_n35_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n108_));
  NA2        u098(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO3        u099(.A(men_men_n109_), .B(men_men_n106_), .C(men_men_n102_), .Y(men_men_n110_));
  NOi21      u100(.An(i_5_), .B(i_2_), .Y(men_men_n111_));
  AOI220     u101(.A0(men_men_n111_), .A1(men_men_n65_), .B0(men_men_n48_), .B1(men_men_n27_), .Y(men_men_n112_));
  AOI210     u102(.A0(men_men_n112_), .A1(men_men_n93_), .B0(men_men_n77_), .Y(men_men_n113_));
  NO4        u103(.A(i_2_), .B(men_men_n17_), .C(men_men_n11_), .D(men_men_n13_), .Y(men_men_n114_));
  NA2        u104(.A(i_2_), .B(i_4_), .Y(men_men_n115_));
  AOI210     u105(.A0(men_men_n81_), .A1(men_men_n63_), .B0(men_men_n115_), .Y(men_men_n116_));
  NO2        u106(.A(i_8_), .B(i_7_), .Y(men_men_n117_));
  OA210      u107(.A0(men_men_n116_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  NA4        u108(.A(men_men_n88_), .B(i_0_), .C(i_5_), .D(men_men_n19_), .Y(men_men_n119_));
  NO2        u109(.A(men_men_n119_), .B(i_4_), .Y(men_men_n120_));
  NO3        u110(.A(men_men_n120_), .B(men_men_n118_), .C(men_men_n113_), .Y(men_men_n121_));
  NA3        u111(.A(men_men_n103_), .B(men_men_n49_), .C(men_men_n82_), .Y(men_men_n122_));
  INV        u112(.A(men_men_n122_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n66_), .B(men_men_n88_), .C(i_0_), .Y(men_men_n124_));
  NOi31      u114(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n125_));
  OAI210     u115(.A0(men_men_n104_), .A1(men_men_n56_), .B0(men_men_n125_), .Y(men_men_n126_));
  NA2        u116(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n127_));
  NO2        u117(.A(men_men_n127_), .B(men_men_n123_), .Y(men_men_n128_));
  NA4        u118(.A(men_men_n128_), .B(men_men_n121_), .C(men_men_n110_), .D(men_men_n99_), .Y(men_men_n129_));
  OR4        u119(.A(men_men_n129_), .B(men_men_n92_), .C(men_men_n62_), .D(men_men_n50_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule