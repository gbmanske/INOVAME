//Benchmark atmr_intb_466_0.5

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n136_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n226_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n375_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n445_, men_men_n446_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NO2        o017(.A(ori_ori_n39_), .B(ori_ori_n34_), .Y(ori00));
  INV        o018(.A(x01), .Y(ori_ori_n41_));
  INV        o019(.A(x06), .Y(ori_ori_n42_));
  NA2        o020(.A(ori_ori_n42_), .B(ori_ori_n28_), .Y(ori_ori_n43_));
  INV        o021(.A(x09), .Y(ori_ori_n44_));
  NO2        o022(.A(x10), .B(x02), .Y(ori_ori_n45_));
  INV        o023(.A(x00), .Y(ori_ori_n46_));
  NO2        o024(.A(ori_ori_n44_), .B(ori_ori_n46_), .Y(ori_ori_n47_));
  INV        o025(.A(ori_ori_n47_), .Y(ori_ori_n48_));
  NA2        o026(.A(x09), .B(ori_ori_n46_), .Y(ori_ori_n49_));
  INV        o027(.A(x07), .Y(ori_ori_n50_));
  NA2        o028(.A(x10), .B(ori_ori_n24_), .Y(ori_ori_n51_));
  NO2        o029(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n50_), .B(ori_ori_n42_), .Y(ori_ori_n53_));
  OAI210     o031(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n53_), .Y(ori_ori_n54_));
  AOI220     o032(.A0(ori_ori_n54_), .A1(ori_ori_n48_), .B0(ori_ori_n52_), .B1(ori_ori_n31_), .Y(ori_ori_n55_));
  NO2        o033(.A(ori_ori_n55_), .B(x05), .Y(ori_ori_n56_));
  NO2        o034(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(x08), .B(x01), .Y(ori_ori_n58_));
  OAI210     o036(.A0(ori_ori_n58_), .A1(ori_ori_n57_), .B0(ori_ori_n35_), .Y(ori_ori_n59_));
  INV        o037(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  NA2        o038(.A(x11), .B(x00), .Y(ori_ori_n61_));
  NO2        o039(.A(x11), .B(ori_ori_n41_), .Y(ori_ori_n62_));
  NOi21      o040(.An(ori_ori_n61_), .B(ori_ori_n62_), .Y(ori_ori_n63_));
  INV        o041(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NOi21      o042(.An(x01), .B(x10), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n29_), .B(ori_ori_n46_), .Y(ori_ori_n66_));
  NO3        o044(.A(ori_ori_n66_), .B(ori_ori_n65_), .C(x06), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n67_), .B(ori_ori_n27_), .Y(ori_ori_n68_));
  OAI210     o046(.A0(ori_ori_n64_), .A1(x07), .B0(ori_ori_n68_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n56_), .Y(ori01));
  INV        o048(.A(x12), .Y(ori_ori_n71_));
  INV        o049(.A(x13), .Y(ori_ori_n72_));
  NO2        o050(.A(x10), .B(x01), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  NA2        o053(.A(ori_ori_n29_), .B(ori_ori_n41_), .Y(ori_ori_n76_));
  NA2        o054(.A(x10), .B(ori_ori_n46_), .Y(ori_ori_n77_));
  NA2        o055(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n78_));
  NA2        o056(.A(ori_ori_n44_), .B(x05), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n49_), .B(x05), .Y(ori_ori_n80_));
  NO2        o058(.A(x09), .B(x05), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n81_), .B(ori_ori_n41_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n75_), .B(ori_ori_n43_), .Y(ori_ori_n83_));
  INV        o061(.A(ori_ori_n83_), .Y(ori_ori_n84_));
  NO2        o062(.A(x03), .B(x02), .Y(ori_ori_n85_));
  OR2        o063(.A(ori_ori_n84_), .B(x11), .Y(ori_ori_n86_));
  INV        o064(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n88_));
  NA2        o066(.A(x01), .B(ori_ori_n77_), .Y(ori_ori_n89_));
  INV        o067(.A(x06), .Y(ori_ori_n90_));
  NA2        o068(.A(ori_ori_n90_), .B(ori_ori_n71_), .Y(ori_ori_n91_));
  AOI210     o069(.A0(x10), .A1(ori_ori_n47_), .B0(ori_ori_n91_), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n92_), .B(ori_ori_n89_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n72_), .B(x12), .Y(ori_ori_n94_));
  NA2        o072(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n96_), .B(x02), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n95_), .B(ori_ori_n93_), .Y(ori_ori_n98_));
  INV        o076(.A(ori_ori_n98_), .Y(ori_ori_n99_));
  AOI210     o077(.A0(ori_ori_n87_), .A1(ori_ori_n71_), .B0(ori_ori_n99_), .Y(ori_ori_n100_));
  NA2        o078(.A(ori_ori_n23_), .B(ori_ori_n41_), .Y(ori_ori_n101_));
  NA2        o079(.A(x13), .B(ori_ori_n71_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n91_), .B(ori_ori_n63_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n103_), .B(x07), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n65_), .B(ori_ori_n105_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n101_), .B(ori_ori_n28_), .Y(ori_ori_n107_));
  OAI210     o085(.A0(ori_ori_n66_), .A1(x06), .B0(ori_ori_n107_), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n108_), .B(ori_ori_n106_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n109_), .B(ori_ori_n104_), .Y(ori_ori_n110_));
  OAI210     o088(.A0(ori_ori_n100_), .A1(ori_ori_n50_), .B0(ori_ori_n110_), .Y(ori02));
  INV        o089(.A(ori_ori_n85_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n112_), .B(ori_ori_n78_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n113_), .B(x13), .Y(ori_ori_n114_));
  NA2        o092(.A(x05), .B(ori_ori_n73_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n79_), .B(ori_ori_n28_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n116_), .B(ori_ori_n74_), .Y(ori_ori_n117_));
  NA3        o095(.A(x12), .B(x12), .C(ori_ori_n78_), .Y(ori_ori_n118_));
  NA4        o096(.A(ori_ori_n118_), .B(ori_ori_n117_), .C(ori_ori_n115_), .D(ori_ori_n42_), .Y(ori_ori_n119_));
  INV        o097(.A(ori_ori_n96_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n121_));
  OAI210     o099(.A0(ori_ori_n120_), .A1(ori_ori_n48_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n122_), .B(x02), .Y(ori_ori_n123_));
  NO3        o101(.A(ori_ori_n94_), .B(ori_ori_n88_), .C(ori_ori_n45_), .Y(ori_ori_n124_));
  INV        o102(.A(ori_ori_n124_), .Y(ori_ori_n125_));
  NA3        o103(.A(ori_ori_n125_), .B(ori_ori_n123_), .C(x06), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n126_), .B(ori_ori_n119_), .Y(ori_ori_n127_));
  OAI210     o105(.A0(ori_ori_n114_), .A1(x12), .B0(ori_ori_n127_), .Y(ori03));
  NA2        o106(.A(ori_ori_n94_), .B(ori_ori_n85_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(ori_ori_n97_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(x05), .Y(ori_ori_n131_));
  NO2        o109(.A(ori_ori_n71_), .B(ori_ori_n82_), .Y(ori_ori_n132_));
  AN2        o110(.A(x12), .B(ori_ori_n80_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n134_), .B(ori_ori_n131_), .Y(ori04));
  NO2        o113(.A(ori_ori_n60_), .B(ori_ori_n39_), .Y(ori_ori_n136_));
  XO2        o114(.A(ori_ori_n136_), .B(ori_ori_n102_), .Y(ori05));
  NA2        o115(.A(ori_ori_n71_), .B(x07), .Y(ori_ori_n138_));
  BUFFER     o116(.A(ori_ori_n102_), .Y(ori_ori_n139_));
  NA3        o117(.A(ori_ori_n139_), .B(ori_ori_n35_), .C(x08), .Y(ori_ori_n140_));
  NO3        o118(.A(x03), .B(ori_ori_n140_), .C(ori_ori_n138_), .Y(ori06));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NO3        m026(.A(x02), .B(x11), .C(x09), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  INV        m029(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(x07), .Y(mai_mai_n53_));
  OAI210     m031(.A0(mai_mai_n53_), .A1(mai_mai_n49_), .B0(mai_mai_n47_), .Y(mai_mai_n54_));
  NOi21      m032(.An(x01), .B(x09), .Y(mai_mai_n55_));
  INV        m033(.A(x00), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n56_), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n57_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(x09), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  INV        m037(.A(x07), .Y(mai_mai_n60_));
  AOI220     m038(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n60_), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n58_), .Y(mai_mai_n62_));
  OAI220     m040(.A0(x02), .A1(mai_mai_n62_), .B0(mai_mai_n61_), .B1(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n60_), .B(mai_mai_n48_), .Y(mai_mai_n64_));
  OAI210     m042(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n64_), .Y(mai_mai_n65_));
  AOI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n58_), .B0(mai_mai_n63_), .B1(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n66_), .B(mai_mai_n54_), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n60_), .B(mai_mai_n23_), .Y(mai_mai_n68_));
  NA2        m046(.A(x09), .B(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x10), .B(x06), .Y(mai_mai_n70_));
  NA2        m048(.A(mai_mai_n70_), .B(mai_mai_n69_), .Y(mai_mai_n71_));
  OAI210     m049(.A0(mai_mai_n71_), .A1(mai_mai_n68_), .B0(x03), .Y(mai_mai_n72_));
  NOi31      m050(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n270_), .B(mai_mai_n24_), .Y(mai_mai_n74_));
  NA2        m052(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n48_), .B(mai_mai_n75_), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n77_));
  NO2        m055(.A(x08), .B(x01), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n78_), .A1(mai_mai_n77_), .B0(mai_mai_n35_), .Y(mai_mai_n79_));
  NO3        m057(.A(mai_mai_n79_), .B(mai_mai_n76_), .C(mai_mai_n74_), .Y(mai_mai_n80_));
  AN2        m058(.A(mai_mai_n80_), .B(mai_mai_n72_), .Y(mai_mai_n81_));
  INV        m059(.A(mai_mai_n79_), .Y(mai_mai_n82_));
  NO2        m060(.A(x06), .B(x05), .Y(mai_mai_n83_));
  NA2        m061(.A(x11), .B(x00), .Y(mai_mai_n84_));
  NO2        m062(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n85_));
  NOi21      m063(.An(mai_mai_n84_), .B(mai_mai_n85_), .Y(mai_mai_n86_));
  INV        m064(.A(mai_mai_n86_), .Y(mai_mai_n87_));
  NO2        m065(.A(mai_mai_n29_), .B(mai_mai_n56_), .Y(mai_mai_n88_));
  NO2        m066(.A(mai_mai_n87_), .B(x07), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n81_), .C(mai_mai_n67_), .Y(mai01));
  INV        m068(.A(x12), .Y(mai_mai_n91_));
  INV        m069(.A(x13), .Y(mai_mai_n92_));
  NA2        m070(.A(x08), .B(x04), .Y(mai_mai_n93_));
  NO2        m071(.A(x10), .B(x01), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n95_));
  NA2        m073(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n55_), .B(x05), .Y(mai_mai_n98_));
  NO2        m076(.A(x04), .B(x05), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n35_), .B(mai_mai_n56_), .Y(mai_mai_n100_));
  INV        m078(.A(mai_mai_n70_), .Y(mai_mai_n101_));
  NA2        m079(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n59_), .B(x05), .Y(mai_mai_n103_));
  NO2        m081(.A(x06), .B(x03), .Y(mai_mai_n104_));
  NO3        m082(.A(mai_mai_n104_), .B(mai_mai_n101_), .C(mai_mai_n97_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n106_));
  NO2        m084(.A(x09), .B(x05), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n107_), .B(mai_mai_n47_), .Y(mai_mai_n108_));
  NA2        m086(.A(x09), .B(x00), .Y(mai_mai_n109_));
  NA2        m087(.A(mai_mai_n98_), .B(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(x03), .B(x02), .Y(mai_mai_n111_));
  INV        m089(.A(mai_mai_n111_), .Y(mai_mai_n112_));
  OA210      m090(.A0(x02), .A1(x11), .B0(mai_mai_n112_), .Y(mai_mai_n113_));
  OAI210     m091(.A0(mai_mai_n105_), .A1(mai_mai_n23_), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  NOi21      m092(.An(x01), .B(x13), .Y(mai_mai_n115_));
  INV        m093(.A(mai_mai_n115_), .Y(mai_mai_n116_));
  NO2        m094(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n92_), .B(x01), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n119_), .B(x08), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n117_), .B(x02), .Y(mai_mai_n121_));
  NA2        m099(.A(x10), .B(x05), .Y(mai_mai_n122_));
  NO2        m100(.A(x09), .B(x01), .Y(mai_mai_n123_));
  NAi21      m101(.An(x13), .B(x00), .Y(mai_mai_n124_));
  AOI210     m102(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  AOI220     m103(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n126_));
  OAI210     m104(.A0(mai_mai_n122_), .A1(mai_mai_n35_), .B0(mai_mai_n126_), .Y(mai_mai_n127_));
  AN2        m105(.A(mai_mai_n127_), .B(mai_mai_n125_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n124_), .B(mai_mai_n36_), .Y(mai_mai_n129_));
  INV        m107(.A(mai_mai_n129_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n128_), .B(x03), .Y(mai_mai_n131_));
  NOi21      m109(.An(x09), .B(x00), .Y(mai_mai_n132_));
  NO3        m110(.A(mai_mai_n77_), .B(mai_mai_n132_), .C(mai_mai_n47_), .Y(mai_mai_n133_));
  INV        m111(.A(mai_mai_n133_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n272_), .B(mai_mai_n134_), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n92_), .B(x12), .Y(mai_mai_n136_));
  AOI210     m114(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n136_), .Y(mai_mai_n137_));
  NO2        m115(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n138_));
  NA2        m116(.A(mai_mai_n137_), .B(mai_mai_n135_), .Y(mai_mai_n139_));
  NA3        m117(.A(mai_mai_n139_), .B(mai_mai_n131_), .C(mai_mai_n121_), .Y(mai_mai_n140_));
  AOI210     m118(.A0(mai_mai_n114_), .A1(mai_mai_n91_), .B0(mai_mai_n140_), .Y(mai_mai_n141_));
  INV        m119(.A(mai_mai_n73_), .Y(mai_mai_n142_));
  NO2        m120(.A(x05), .B(mai_mai_n50_), .Y(mai_mai_n143_));
  OAI210     m121(.A0(mai_mai_n143_), .A1(mai_mai_n116_), .B0(mai_mai_n56_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n144_), .B(mai_mai_n142_), .Y(mai_mai_n145_));
  AOI210     m123(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n50_), .Y(mai_mai_n146_));
  NO2        m124(.A(mai_mai_n146_), .B(mai_mai_n41_), .Y(mai_mai_n147_));
  NA3        m125(.A(mai_mai_n55_), .B(mai_mai_n36_), .C(x04), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n106_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n149_), .A1(mai_mai_n147_), .B0(x02), .Y(mai_mai_n150_));
  AOI210     m128(.A0(mai_mai_n150_), .A1(mai_mai_n145_), .B0(mai_mai_n23_), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n273_), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  INV        m130(.A(mai_mai_n85_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n153_), .B(x12), .Y(mai_mai_n154_));
  NO2        m132(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n155_));
  OAI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n127_), .B0(mai_mai_n125_), .Y(mai_mai_n156_));
  AOI210     m134(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n157_), .B(mai_mai_n41_), .Y(mai_mai_n158_));
  OAI210     m136(.A0(mai_mai_n93_), .A1(mai_mai_n109_), .B0(mai_mai_n70_), .Y(mai_mai_n159_));
  NO2        m137(.A(mai_mai_n159_), .B(mai_mai_n158_), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n161_));
  NA2        m139(.A(mai_mai_n161_), .B(x03), .Y(mai_mai_n162_));
  OA210      m140(.A0(mai_mai_n162_), .A1(mai_mai_n160_), .B0(mai_mai_n156_), .Y(mai_mai_n163_));
  NA2        m141(.A(x13), .B(mai_mai_n91_), .Y(mai_mai_n164_));
  NA2        m142(.A(x12), .B(mai_mai_n86_), .Y(mai_mai_n165_));
  OAI210     m143(.A0(mai_mai_n163_), .A1(x01), .B0(mai_mai_n165_), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n154_), .B(mai_mai_n166_), .Y(mai_mai_n167_));
  AOI210     m145(.A0(mai_mai_n167_), .A1(mai_mai_n152_), .B0(x07), .Y(mai_mai_n168_));
  NO2        m146(.A(x08), .B(x05), .Y(mai_mai_n169_));
  NO2        m147(.A(x12), .B(x02), .Y(mai_mai_n170_));
  NO2        m148(.A(x05), .B(x01), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n92_), .B(x04), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n57_), .B(x05), .Y(mai_mai_n173_));
  INV        m151(.A(mai_mai_n168_), .Y(mai_mai_n174_));
  OAI210     m152(.A0(mai_mai_n141_), .A1(mai_mai_n60_), .B0(mai_mai_n174_), .Y(mai02));
  NA2        m153(.A(x04), .B(mai_mai_n55_), .Y(mai_mai_n176_));
  NA2        m154(.A(mai_mai_n32_), .B(mai_mai_n176_), .Y(mai_mai_n177_));
  INV        m155(.A(mai_mai_n177_), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n122_), .Y(mai_mai_n179_));
  NA2        m157(.A(x13), .B(mai_mai_n179_), .Y(mai_mai_n180_));
  AOI210     m158(.A0(mai_mai_n180_), .A1(mai_mai_n178_), .B0(mai_mai_n48_), .Y(mai_mai_n181_));
  AOI210     m159(.A0(mai_mai_n169_), .A1(mai_mai_n57_), .B0(mai_mai_n55_), .Y(mai_mai_n182_));
  NOi21      m160(.An(x04), .B(mai_mai_n182_), .Y(mai_mai_n183_));
  INV        m161(.A(mai_mai_n183_), .Y(mai_mai_n184_));
  AOI210     m162(.A0(mai_mai_n184_), .A1(x02), .B0(mai_mai_n106_), .Y(mai_mai_n185_));
  NO2        m163(.A(mai_mai_n161_), .B(mai_mai_n47_), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n186_), .Y(mai_mai_n187_));
  OAI210     m165(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n48_), .B(mai_mai_n88_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n187_), .Y(mai_mai_n190_));
  NO3        m168(.A(mai_mai_n190_), .B(mai_mai_n185_), .C(mai_mai_n181_), .Y(mai_mai_n191_));
  NA2        m169(.A(x09), .B(x03), .Y(mai_mai_n192_));
  INV        m170(.A(mai_mai_n124_), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n35_), .B(mai_mai_n36_), .Y(mai_mai_n194_));
  AOI220     m172(.A0(mai_mai_n194_), .A1(mai_mai_n193_), .B0(mai_mai_n138_), .B1(x08), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n195_), .B(mai_mai_n192_), .Y(mai_mai_n196_));
  NA2        m174(.A(mai_mai_n196_), .B(mai_mai_n94_), .Y(mai_mai_n197_));
  OAI210     m175(.A0(mai_mai_n55_), .A1(x05), .B0(mai_mai_n95_), .Y(mai_mai_n198_));
  NA3        m176(.A(mai_mai_n198_), .B(mai_mai_n197_), .C(mai_mai_n48_), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n138_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n136_), .B(x04), .Y(mai_mai_n201_));
  INV        m179(.A(mai_mai_n201_), .Y(mai_mai_n202_));
  NO3        m180(.A(mai_mai_n126_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n203_));
  OAI210     m181(.A0(mai_mai_n203_), .A1(mai_mai_n202_), .B0(mai_mai_n88_), .Y(mai_mai_n204_));
  NO3        m182(.A(mai_mai_n136_), .B(mai_mai_n118_), .C(mai_mai_n51_), .Y(mai_mai_n205_));
  OAI210     m183(.A0(x12), .A1(mai_mai_n133_), .B0(mai_mai_n205_), .Y(mai_mai_n206_));
  NA3        m184(.A(mai_mai_n206_), .B(mai_mai_n204_), .C(x06), .Y(mai_mai_n207_));
  NO3        m185(.A(mai_mai_n173_), .B(x01), .C(x08), .Y(mai_mai_n208_));
  INV        m186(.A(mai_mai_n208_), .Y(mai_mai_n209_));
  NA2        m187(.A(mai_mai_n205_), .B(x05), .Y(mai_mai_n210_));
  OAI210     m188(.A0(mai_mai_n209_), .A1(mai_mai_n28_), .B0(mai_mai_n210_), .Y(mai_mai_n211_));
  AN2        m189(.A(mai_mai_n211_), .B(x04), .Y(mai_mai_n212_));
  AOI210     m190(.A0(mai_mai_n207_), .A1(mai_mai_n199_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  OAI210     m191(.A0(mai_mai_n191_), .A1(x12), .B0(mai_mai_n213_), .Y(mai03));
  NA2        m192(.A(mai_mai_n274_), .B(x05), .Y(mai_mai_n215_));
  NO2        m193(.A(x08), .B(mai_mai_n99_), .Y(mai_mai_n216_));
  OAI220     m194(.A0(mai_mai_n216_), .A1(mai_mai_n58_), .B0(x02), .B1(mai_mai_n182_), .Y(mai_mai_n217_));
  OAI210     m195(.A0(mai_mai_n217_), .A1(x05), .B0(mai_mai_n91_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n123_), .B(mai_mai_n103_), .Y(mai_mai_n219_));
  OAI220     m197(.A0(mai_mai_n219_), .A1(mai_mai_n37_), .B0(mai_mai_n110_), .B1(x13), .Y(mai_mai_n220_));
  OAI210     m198(.A0(mai_mai_n220_), .A1(mai_mai_n275_), .B0(x04), .Y(mai_mai_n221_));
  AOI210     m199(.A0(mai_mai_n130_), .A1(mai_mai_n91_), .B0(mai_mai_n108_), .Y(mai_mai_n222_));
  OA210      m200(.A0(mai_mai_n120_), .A1(x12), .B0(mai_mai_n103_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n223_), .B(mai_mai_n222_), .Y(mai_mai_n224_));
  NA4        m202(.A(mai_mai_n224_), .B(mai_mai_n221_), .C(mai_mai_n218_), .D(mai_mai_n215_), .Y(mai04));
  NO2        m203(.A(mai_mai_n82_), .B(mai_mai_n39_), .Y(mai_mai_n226_));
  XO2        m204(.A(mai_mai_n226_), .B(mai_mai_n164_), .Y(mai05));
  NA2        m205(.A(mai_mai_n69_), .B(mai_mai_n51_), .Y(mai_mai_n228_));
  AOI210     m206(.A0(mai_mai_n228_), .A1(mai_mai_n188_), .B0(mai_mai_n25_), .Y(mai_mai_n229_));
  NA3        m207(.A(mai_mai_n106_), .B(mai_mai_n102_), .C(mai_mai_n31_), .Y(mai_mai_n230_));
  AOI210     m208(.A0(mai_mai_n271_), .A1(mai_mai_n230_), .B0(mai_mai_n24_), .Y(mai_mai_n231_));
  OAI210     m209(.A0(mai_mai_n231_), .A1(mai_mai_n229_), .B0(mai_mai_n91_), .Y(mai_mai_n232_));
  NA2        m210(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n234_));
  NA2        m212(.A(x10), .B(x03), .Y(mai_mai_n235_));
  OAI220     m213(.A0(mai_mai_n235_), .A1(mai_mai_n234_), .B0(mai_mai_n233_), .B1(mai_mai_n75_), .Y(mai_mai_n236_));
  OAI210     m214(.A0(mai_mai_n26_), .A1(mai_mai_n91_), .B0(x07), .Y(mai_mai_n237_));
  AOI210     m215(.A0(mai_mai_n236_), .A1(x06), .B0(mai_mai_n237_), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n33_), .B(mai_mai_n91_), .Y(mai_mai_n239_));
  AOI210     m217(.A0(mai_mai_n239_), .A1(mai_mai_n85_), .B0(x07), .Y(mai_mai_n240_));
  AOI210     m218(.A0(mai_mai_n238_), .A1(mai_mai_n232_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  AOI210     m219(.A0(mai_mai_n201_), .A1(mai_mai_n96_), .B0(mai_mai_n170_), .Y(mai_mai_n242_));
  NOi21      m220(.An(mai_mai_n192_), .B(mai_mai_n103_), .Y(mai_mai_n243_));
  OAI210     m221(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n244_));
  AOI210     m222(.A0(mai_mai_n164_), .A1(mai_mai_n47_), .B0(mai_mai_n244_), .Y(mai_mai_n245_));
  NO3        m223(.A(mai_mai_n245_), .B(mai_mai_n242_), .C(x08), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n102_), .B(mai_mai_n28_), .Y(mai_mai_n247_));
  NO2        m225(.A(mai_mai_n247_), .B(mai_mai_n171_), .Y(mai_mai_n248_));
  NA3        m226(.A(mai_mai_n200_), .B(mai_mai_n100_), .C(x12), .Y(mai_mai_n249_));
  AO210      m227(.A0(mai_mai_n200_), .A1(mai_mai_n100_), .B0(mai_mai_n164_), .Y(mai_mai_n250_));
  NA3        m228(.A(mai_mai_n250_), .B(mai_mai_n249_), .C(x08), .Y(mai_mai_n251_));
  INV        m229(.A(mai_mai_n251_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n246_), .B(mai_mai_n252_), .Y(mai_mai_n253_));
  INV        m231(.A(x03), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n107_), .B(mai_mai_n43_), .Y(mai_mai_n255_));
  OAI210     m233(.A0(mai_mai_n255_), .A1(mai_mai_n254_), .B0(mai_mai_n129_), .Y(mai_mai_n256_));
  NA3        m234(.A(mai_mai_n248_), .B(mai_mai_n243_), .C(x12), .Y(mai_mai_n257_));
  INV        m235(.A(x14), .Y(mai_mai_n258_));
  NO3        m236(.A(mai_mai_n119_), .B(x05), .C(mai_mai_n56_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n259_), .B(mai_mai_n258_), .Y(mai_mai_n260_));
  NA3        m238(.A(mai_mai_n260_), .B(mai_mai_n257_), .C(mai_mai_n256_), .Y(mai_mai_n261_));
  NA2        m239(.A(mai_mai_n239_), .B(mai_mai_n60_), .Y(mai_mai_n262_));
  NOi21      m240(.An(mai_mai_n172_), .B(mai_mai_n110_), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n264_));
  OAI210     m242(.A0(mai_mai_n264_), .A1(mai_mai_n263_), .B0(mai_mai_n91_), .Y(mai_mai_n265_));
  OAI210     m243(.A0(mai_mai_n262_), .A1(mai_mai_n84_), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  NO4        m244(.A(mai_mai_n266_), .B(mai_mai_n261_), .C(mai_mai_n253_), .D(mai_mai_n241_), .Y(mai06));
  INV        m245(.A(x07), .Y(mai_mai_n270_));
  INV        m246(.A(mai_mai_n83_), .Y(mai_mai_n271_));
  INV        m247(.A(x12), .Y(mai_mai_n272_));
  INV        m248(.A(x12), .Y(mai_mai_n273_));
  INV        m249(.A(mai_mai_n42_), .Y(mai_mai_n274_));
  INV        m250(.A(mai_mai_n38_), .Y(mai_mai_n275_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  INV        u003(.A(x02), .Y(men_men_n26_));
  INV        u004(.A(x10), .Y(men_men_n27_));
  NA2        u005(.A(men_men_n27_), .B(men_men_n26_), .Y(men_men_n28_));
  INV        u006(.A(x03), .Y(men_men_n29_));
  NA2        u007(.A(x10), .B(men_men_n29_), .Y(men_men_n30_));
  INV        u008(.A(x04), .Y(men_men_n31_));
  INV        u009(.A(x08), .Y(men_men_n32_));
  NA2        u010(.A(x08), .B(x03), .Y(men_men_n33_));
  NO2        u011(.A(men_men_n33_), .B(men_men_n31_), .Y(men_men_n34_));
  NA2        u012(.A(x09), .B(men_men_n29_), .Y(men_men_n35_));
  INV        u013(.A(x05), .Y(men_men_n36_));
  NO2        u014(.A(x09), .B(x02), .Y(men_men_n37_));
  NO2        u015(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NA2        u016(.A(men_men_n38_), .B(men_men_n35_), .Y(men_men_n39_));
  INV        u017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u018(.A(men_men_n40_), .B(men_men_n34_), .Y(men00));
  INV        u019(.A(x01), .Y(men_men_n42_));
  INV        u020(.A(x06), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n26_), .Y(men_men_n44_));
  INV        u022(.A(x09), .Y(men_men_n45_));
  NO2        u023(.A(x10), .B(x02), .Y(men_men_n46_));
  NO2        u024(.A(x09), .B(x07), .Y(men_men_n47_));
  OAI210     u025(.A0(men_men_n47_), .A1(men_men_n43_), .B0(men_men_n42_), .Y(men_men_n48_));
  NOi21      u026(.An(x01), .B(x09), .Y(men_men_n49_));
  INV        u027(.A(x00), .Y(men_men_n50_));
  NO2        u028(.A(men_men_n45_), .B(men_men_n50_), .Y(men_men_n51_));
  NO2        u029(.A(men_men_n51_), .B(men_men_n49_), .Y(men_men_n52_));
  NA2        u030(.A(x09), .B(men_men_n50_), .Y(men_men_n53_));
  INV        u031(.A(x07), .Y(men_men_n54_));
  NA2        u032(.A(men_men_n27_), .B(x02), .Y(men_men_n55_));
  NA2        u033(.A(men_men_n52_), .B(men_men_n29_), .Y(men_men_n56_));
  AOI210     u034(.A0(men_men_n56_), .A1(men_men_n48_), .B0(x05), .Y(men_men_n57_));
  NA2        u035(.A(x10), .B(x09), .Y(men_men_n58_));
  NA2        u036(.A(x09), .B(x05), .Y(men_men_n59_));
  NA2        u037(.A(x10), .B(x06), .Y(men_men_n60_));
  NA3        u038(.A(men_men_n60_), .B(men_men_n59_), .C(men_men_n26_), .Y(men_men_n61_));
  NO2        u039(.A(men_men_n54_), .B(men_men_n36_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n61_), .B(x03), .Y(men_men_n63_));
  NOi31      u041(.An(x08), .B(x04), .C(x00), .Y(men_men_n64_));
  NO2        u042(.A(x10), .B(x09), .Y(men_men_n65_));
  NO2        u043(.A(x09), .B(men_men_n36_), .Y(men_men_n66_));
  NO2        u044(.A(men_men_n66_), .B(men_men_n32_), .Y(men_men_n67_));
  OAI210     u045(.A0(men_men_n66_), .A1(men_men_n27_), .B0(x02), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n67_), .A1(men_men_n43_), .B0(men_men_n68_), .Y(men_men_n69_));
  NO2        u047(.A(men_men_n32_), .B(x00), .Y(men_men_n70_));
  NO2        u048(.A(x08), .B(x01), .Y(men_men_n71_));
  OAI210     u049(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n31_), .Y(men_men_n72_));
  NA2        u050(.A(men_men_n45_), .B(men_men_n32_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n72_), .B(men_men_n69_), .Y(men_men_n74_));
  AN2        u052(.A(men_men_n74_), .B(men_men_n63_), .Y(men_men_n75_));
  INV        u053(.A(men_men_n72_), .Y(men_men_n76_));
  NO2        u054(.A(x06), .B(x05), .Y(men_men_n77_));
  NA2        u055(.A(x11), .B(x00), .Y(men_men_n78_));
  NO2        u056(.A(x11), .B(men_men_n42_), .Y(men_men_n79_));
  NOi21      u057(.An(men_men_n78_), .B(men_men_n79_), .Y(men_men_n80_));
  AOI210     u058(.A0(men_men_n77_), .A1(men_men_n76_), .B0(men_men_n80_), .Y(men_men_n81_));
  NOi21      u059(.An(x01), .B(x10), .Y(men_men_n82_));
  NO2        u060(.A(men_men_n27_), .B(men_men_n50_), .Y(men_men_n83_));
  NO3        u061(.A(men_men_n83_), .B(men_men_n82_), .C(x06), .Y(men_men_n84_));
  INV        u062(.A(men_men_n84_), .Y(men_men_n85_));
  OAI210     u063(.A0(men_men_n81_), .A1(x07), .B0(men_men_n85_), .Y(men_men_n86_));
  NO3        u064(.A(men_men_n86_), .B(men_men_n75_), .C(men_men_n57_), .Y(men01));
  INV        u065(.A(x12), .Y(men_men_n88_));
  INV        u066(.A(x13), .Y(men_men_n89_));
  NA2        u067(.A(x08), .B(x04), .Y(men_men_n90_));
  NO2        u068(.A(men_men_n90_), .B(men_men_n50_), .Y(men_men_n91_));
  NA2        u069(.A(men_men_n91_), .B(men_men_n77_), .Y(men_men_n92_));
  NA2        u070(.A(men_men_n82_), .B(men_men_n26_), .Y(men_men_n93_));
  NO2        u071(.A(men_men_n93_), .B(men_men_n59_), .Y(men_men_n94_));
  NO2        u072(.A(x10), .B(x01), .Y(men_men_n95_));
  NO2        u073(.A(men_men_n27_), .B(x00), .Y(men_men_n96_));
  NO2        u074(.A(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  NA2        u075(.A(x04), .B(men_men_n26_), .Y(men_men_n98_));
  NO3        u076(.A(men_men_n98_), .B(men_men_n32_), .C(men_men_n36_), .Y(men_men_n99_));
  AOI210     u077(.A0(men_men_n99_), .A1(men_men_n97_), .B0(men_men_n94_), .Y(men_men_n100_));
  AOI210     u078(.A0(men_men_n100_), .A1(men_men_n92_), .B0(men_men_n89_), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n49_), .B(x05), .Y(men_men_n102_));
  NOi21      u080(.An(men_men_n102_), .B(men_men_n51_), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n31_), .B(x02), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n89_), .B(men_men_n32_), .Y(men_men_n105_));
  NA3        u083(.A(men_men_n105_), .B(men_men_n104_), .C(x06), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n103_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n71_), .B(x13), .Y(men_men_n108_));
  NA2        u086(.A(x09), .B(men_men_n31_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n108_), .Y(men_men_n110_));
  NA2        u088(.A(x13), .B(men_men_n31_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n111_), .B(x05), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n112_), .B(men_men_n110_), .Y(men_men_n113_));
  NA2        u091(.A(men_men_n31_), .B(men_men_n50_), .Y(men_men_n114_));
  NA2        u092(.A(men_men_n114_), .B(men_men_n89_), .Y(men_men_n115_));
  AOI210     u093(.A0(men_men_n115_), .A1(men_men_n67_), .B0(men_men_n103_), .Y(men_men_n116_));
  AOI210     u094(.A0(men_men_n116_), .A1(men_men_n113_), .B0(men_men_n60_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n27_), .B(men_men_n42_), .Y(men_men_n118_));
  NA2        u096(.A(x10), .B(men_men_n50_), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n45_), .B(x05), .Y(men_men_n121_));
  NA2        u099(.A(men_men_n32_), .B(x04), .Y(men_men_n122_));
  NA3        u100(.A(men_men_n122_), .B(men_men_n121_), .C(x13), .Y(men_men_n123_));
  NO3        u101(.A(men_men_n114_), .B(men_men_n66_), .C(men_men_n32_), .Y(men_men_n124_));
  NO2        u102(.A(men_men_n53_), .B(x05), .Y(men_men_n125_));
  NOi41      u103(.An(men_men_n123_), .B(men_men_n125_), .C(men_men_n124_), .D(men_men_n120_), .Y(men_men_n126_));
  NO3        u104(.A(men_men_n126_), .B(x06), .C(x03), .Y(men_men_n127_));
  NO4        u105(.A(men_men_n127_), .B(men_men_n117_), .C(men_men_n107_), .D(men_men_n101_), .Y(men_men_n128_));
  NA2        u106(.A(x13), .B(men_men_n32_), .Y(men_men_n129_));
  OAI210     u107(.A0(men_men_n71_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n130_), .B(men_men_n129_), .Y(men_men_n131_));
  NOi21      u109(.An(men_men_n77_), .B(men_men_n50_), .Y(men_men_n132_));
  NO2        u110(.A(men_men_n31_), .B(men_men_n42_), .Y(men_men_n133_));
  OA210      u111(.A0(men_men_n132_), .A1(men_men_n65_), .B0(men_men_n133_), .Y(men_men_n134_));
  NO2        u112(.A(men_men_n45_), .B(men_men_n36_), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n27_), .B(x06), .Y(men_men_n136_));
  AOI210     u114(.A0(men_men_n136_), .A1(men_men_n44_), .B0(men_men_n135_), .Y(men_men_n137_));
  OA210      u115(.A0(men_men_n137_), .A1(men_men_n134_), .B0(men_men_n131_), .Y(men_men_n138_));
  NO2        u116(.A(x09), .B(x05), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(men_men_n42_), .Y(men_men_n140_));
  AOI210     u118(.A0(men_men_n140_), .A1(men_men_n97_), .B0(men_men_n44_), .Y(men_men_n141_));
  NA2        u119(.A(x09), .B(x00), .Y(men_men_n142_));
  NA2        u120(.A(men_men_n102_), .B(men_men_n142_), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n64_), .B(men_men_n45_), .Y(men_men_n144_));
  AOI210     u122(.A0(men_men_n144_), .A1(men_men_n143_), .B0(men_men_n136_), .Y(men_men_n145_));
  NO3        u123(.A(men_men_n145_), .B(men_men_n141_), .C(men_men_n138_), .Y(men_men_n146_));
  NO2        u124(.A(x03), .B(x02), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n72_), .B(men_men_n89_), .Y(men_men_n148_));
  OAI210     u126(.A0(men_men_n148_), .A1(men_men_n103_), .B0(men_men_n147_), .Y(men_men_n149_));
  OA210      u127(.A0(men_men_n146_), .A1(x11), .B0(men_men_n149_), .Y(men_men_n150_));
  OAI210     u128(.A0(men_men_n128_), .A1(men_men_n23_), .B0(men_men_n150_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n97_), .B(men_men_n35_), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n23_), .B(men_men_n32_), .Y(men_men_n153_));
  NAi21      u131(.An(x06), .B(x10), .Y(men_men_n154_));
  NOi21      u132(.An(x01), .B(x13), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  OR2        u134(.A(men_men_n156_), .B(men_men_n153_), .Y(men_men_n157_));
  AOI210     u135(.A0(men_men_n157_), .A1(men_men_n152_), .B0(men_men_n36_), .Y(men_men_n158_));
  NO2        u136(.A(men_men_n27_), .B(x03), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n89_), .B(x01), .Y(men_men_n160_));
  NO2        u138(.A(men_men_n160_), .B(x08), .Y(men_men_n161_));
  OAI210     u139(.A0(x05), .A1(men_men_n161_), .B0(men_men_n45_), .Y(men_men_n162_));
  AOI210     u140(.A0(men_men_n162_), .A1(men_men_n159_), .B0(men_men_n43_), .Y(men_men_n163_));
  AOI210     u141(.A0(x11), .A1(men_men_n29_), .B0(men_men_n26_), .Y(men_men_n164_));
  OAI210     u142(.A0(men_men_n163_), .A1(men_men_n158_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u143(.A(x04), .B(x02), .Y(men_men_n166_));
  NA2        u144(.A(x10), .B(x05), .Y(men_men_n167_));
  NA2        u145(.A(x09), .B(x06), .Y(men_men_n168_));
  AOI210     u146(.A0(men_men_n168_), .A1(men_men_n167_), .B0(men_men_n153_), .Y(men_men_n169_));
  NO2        u147(.A(x09), .B(x01), .Y(men_men_n170_));
  NO2        u148(.A(men_men_n170_), .B(men_men_n29_), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n171_), .A1(men_men_n169_), .B0(x00), .Y(men_men_n172_));
  NO2        u150(.A(men_men_n102_), .B(x08), .Y(men_men_n173_));
  NA3        u151(.A(men_men_n155_), .B(men_men_n154_), .C(men_men_n45_), .Y(men_men_n174_));
  NA2        u152(.A(men_men_n82_), .B(x05), .Y(men_men_n175_));
  OAI210     u153(.A0(men_men_n175_), .A1(men_men_n105_), .B0(men_men_n174_), .Y(men_men_n176_));
  AOI210     u154(.A0(men_men_n173_), .A1(x06), .B0(men_men_n176_), .Y(men_men_n177_));
  OAI210     u155(.A0(men_men_n177_), .A1(x11), .B0(men_men_n172_), .Y(men_men_n178_));
  NAi21      u156(.An(men_men_n166_), .B(men_men_n178_), .Y(men_men_n179_));
  INV        u157(.A(men_men_n25_), .Y(men_men_n180_));
  NAi21      u158(.An(x13), .B(x00), .Y(men_men_n181_));
  AOI210     u159(.A0(men_men_n27_), .A1(men_men_n43_), .B0(men_men_n181_), .Y(men_men_n182_));
  AOI220     u160(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n167_), .A1(men_men_n31_), .B0(men_men_n183_), .Y(men_men_n184_));
  AN2        u162(.A(men_men_n184_), .B(men_men_n182_), .Y(men_men_n185_));
  NO2        u163(.A(men_men_n83_), .B(x06), .Y(men_men_n186_));
  NO2        u164(.A(men_men_n181_), .B(men_men_n32_), .Y(men_men_n187_));
  INV        u165(.A(men_men_n187_), .Y(men_men_n188_));
  OAI220     u166(.A0(men_men_n188_), .A1(men_men_n168_), .B0(men_men_n186_), .B1(men_men_n59_), .Y(men_men_n189_));
  OAI210     u167(.A0(men_men_n189_), .A1(men_men_n185_), .B0(men_men_n180_), .Y(men_men_n190_));
  NOi21      u168(.An(x09), .B(x00), .Y(men_men_n191_));
  NA2        u169(.A(x10), .B(x08), .Y(men_men_n192_));
  INV        u170(.A(men_men_n192_), .Y(men_men_n193_));
  NA2        u171(.A(x06), .B(x05), .Y(men_men_n194_));
  OAI210     u172(.A0(men_men_n194_), .A1(men_men_n31_), .B0(men_men_n88_), .Y(men_men_n195_));
  AOI210     u173(.A0(men_men_n193_), .A1(men_men_n51_), .B0(men_men_n195_), .Y(men_men_n196_));
  INV        u174(.A(men_men_n196_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n89_), .B(x12), .Y(men_men_n198_));
  AOI210     u176(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n198_), .Y(men_men_n199_));
  NA2        u177(.A(men_men_n82_), .B(men_men_n45_), .Y(men_men_n200_));
  NO2        u178(.A(men_men_n31_), .B(men_men_n29_), .Y(men_men_n201_));
  NA2        u179(.A(men_men_n201_), .B(x02), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n202_), .B(men_men_n200_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n199_), .A1(men_men_n197_), .B0(men_men_n203_), .Y(men_men_n204_));
  NA4        u182(.A(men_men_n204_), .B(men_men_n190_), .C(men_men_n179_), .D(men_men_n165_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n151_), .A1(men_men_n88_), .B0(men_men_n205_), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n129_), .A1(x09), .B0(men_men_n61_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(men_men_n131_), .Y(men_men_n208_));
  NA2        u186(.A(men_men_n45_), .B(men_men_n42_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n209_), .B(men_men_n130_), .Y(men_men_n210_));
  AOI210     u188(.A0(men_men_n28_), .A1(x06), .B0(x05), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n118_), .B(x06), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n211_), .A1(men_men_n210_), .B0(men_men_n212_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n213_), .A1(men_men_n208_), .B0(x12), .Y(men_men_n214_));
  INV        u192(.A(men_men_n64_), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n192_), .A1(x05), .B0(men_men_n45_), .Y(men_men_n216_));
  OAI210     u194(.A0(men_men_n216_), .A1(men_men_n156_), .B0(men_men_n50_), .Y(men_men_n217_));
  NA2        u195(.A(men_men_n217_), .B(men_men_n215_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n82_), .B(x06), .Y(men_men_n219_));
  AOI210     u197(.A0(men_men_n32_), .A1(x04), .B0(men_men_n45_), .Y(men_men_n220_));
  NO3        u198(.A(men_men_n220_), .B(men_men_n219_), .C(men_men_n36_), .Y(men_men_n221_));
  NA4        u199(.A(men_men_n154_), .B(men_men_n49_), .C(men_men_n32_), .D(x04), .Y(men_men_n222_));
  NA2        u200(.A(men_men_n222_), .B(men_men_n136_), .Y(men_men_n223_));
  OAI210     u201(.A0(men_men_n223_), .A1(men_men_n221_), .B0(x02), .Y(men_men_n224_));
  AOI210     u202(.A0(men_men_n224_), .A1(men_men_n218_), .B0(men_men_n23_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n214_), .A1(men_men_n50_), .B0(men_men_n225_), .Y(men_men_n226_));
  INV        u204(.A(men_men_n136_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n45_), .B(x03), .Y(men_men_n228_));
  OAI210     u206(.A0(men_men_n66_), .A1(men_men_n32_), .B0(men_men_n109_), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n89_), .B(x03), .Y(men_men_n230_));
  AOI220     u208(.A0(men_men_n230_), .A1(men_men_n229_), .B0(men_men_n64_), .B1(men_men_n228_), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n30_), .B(x06), .Y(men_men_n232_));
  INV        u210(.A(men_men_n154_), .Y(men_men_n233_));
  NOi21      u211(.An(x13), .B(x04), .Y(men_men_n234_));
  NO3        u212(.A(men_men_n234_), .B(men_men_n64_), .C(men_men_n191_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n235_), .B(x05), .Y(men_men_n236_));
  AOI220     u214(.A0(men_men_n236_), .A1(men_men_n232_), .B0(men_men_n233_), .B1(men_men_n50_), .Y(men_men_n237_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n227_), .B0(men_men_n237_), .Y(men_men_n238_));
  INV        u216(.A(men_men_n79_), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n23_), .B(men_men_n42_), .Y(men_men_n240_));
  NO2        u218(.A(men_men_n45_), .B(men_men_n32_), .Y(men_men_n241_));
  OAI210     u219(.A0(men_men_n241_), .A1(men_men_n184_), .B0(men_men_n182_), .Y(men_men_n242_));
  AOI210     u220(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n243_));
  NO2        u221(.A(x06), .B(x00), .Y(men_men_n244_));
  NO3        u222(.A(men_men_n244_), .B(men_men_n243_), .C(men_men_n36_), .Y(men_men_n245_));
  OAI210     u223(.A0(men_men_n90_), .A1(men_men_n142_), .B0(men_men_n60_), .Y(men_men_n246_));
  NO2        u224(.A(men_men_n246_), .B(men_men_n245_), .Y(men_men_n247_));
  NA2        u225(.A(men_men_n27_), .B(men_men_n43_), .Y(men_men_n248_));
  INV        u226(.A(x03), .Y(men_men_n249_));
  OA210      u227(.A0(men_men_n249_), .A1(men_men_n247_), .B0(men_men_n242_), .Y(men_men_n250_));
  NA2        u228(.A(x13), .B(men_men_n88_), .Y(men_men_n251_));
  NA3        u229(.A(men_men_n251_), .B(men_men_n195_), .C(men_men_n80_), .Y(men_men_n252_));
  OAI210     u230(.A0(men_men_n250_), .A1(men_men_n240_), .B0(men_men_n252_), .Y(men_men_n253_));
  AOI210     u231(.A0(men_men_n79_), .A1(men_men_n238_), .B0(men_men_n253_), .Y(men_men_n254_));
  AOI210     u232(.A0(men_men_n254_), .A1(men_men_n226_), .B0(x07), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n59_), .B(men_men_n27_), .Y(men_men_n256_));
  NOi31      u234(.An(men_men_n129_), .B(men_men_n234_), .C(men_men_n191_), .Y(men_men_n257_));
  AOI210     u235(.A0(men_men_n257_), .A1(men_men_n144_), .B0(men_men_n256_), .Y(men_men_n258_));
  NO2        u236(.A(men_men_n89_), .B(x06), .Y(men_men_n259_));
  INV        u237(.A(men_men_n259_), .Y(men_men_n260_));
  NO2        u238(.A(x08), .B(x05), .Y(men_men_n261_));
  NO2        u239(.A(men_men_n261_), .B(men_men_n243_), .Y(men_men_n262_));
  OAI210     u240(.A0(men_men_n64_), .A1(x13), .B0(men_men_n29_), .Y(men_men_n263_));
  OAI210     u241(.A0(men_men_n262_), .A1(men_men_n260_), .B0(men_men_n263_), .Y(men_men_n264_));
  NO2        u242(.A(x12), .B(x02), .Y(men_men_n265_));
  INV        u243(.A(men_men_n265_), .Y(men_men_n266_));
  NO2        u244(.A(men_men_n266_), .B(men_men_n239_), .Y(men_men_n267_));
  OA210      u245(.A0(men_men_n264_), .A1(men_men_n258_), .B0(men_men_n267_), .Y(men_men_n268_));
  NA2        u246(.A(men_men_n45_), .B(men_men_n36_), .Y(men_men_n269_));
  NO2        u247(.A(men_men_n269_), .B(x01), .Y(men_men_n270_));
  NOi21      u248(.An(men_men_n71_), .B(men_men_n109_), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n271_), .B(men_men_n270_), .Y(men_men_n272_));
  AOI210     u250(.A0(men_men_n272_), .A1(men_men_n123_), .B0(men_men_n27_), .Y(men_men_n273_));
  NA2        u251(.A(men_men_n259_), .B(men_men_n229_), .Y(men_men_n274_));
  NA2        u252(.A(men_men_n89_), .B(x04), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n275_), .B(men_men_n26_), .Y(men_men_n276_));
  OAI210     u254(.A0(men_men_n276_), .A1(men_men_n108_), .B0(men_men_n274_), .Y(men_men_n277_));
  NO3        u255(.A(men_men_n78_), .B(x12), .C(x03), .Y(men_men_n278_));
  OAI210     u256(.A0(men_men_n277_), .A1(men_men_n273_), .B0(men_men_n278_), .Y(men_men_n279_));
  AOI210     u257(.A0(men_men_n200_), .A1(men_men_n194_), .B0(men_men_n90_), .Y(men_men_n280_));
  NOi21      u258(.An(men_men_n256_), .B(men_men_n219_), .Y(men_men_n281_));
  NO2        u259(.A(men_men_n25_), .B(x00), .Y(men_men_n282_));
  OAI210     u260(.A0(men_men_n281_), .A1(men_men_n280_), .B0(men_men_n282_), .Y(men_men_n283_));
  NO2        u261(.A(men_men_n51_), .B(x05), .Y(men_men_n284_));
  NO3        u262(.A(men_men_n284_), .B(men_men_n220_), .C(men_men_n186_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n240_), .B(men_men_n26_), .Y(men_men_n286_));
  OAI210     u264(.A0(men_men_n285_), .A1(men_men_n227_), .B0(men_men_n286_), .Y(men_men_n287_));
  NA3        u265(.A(men_men_n287_), .B(men_men_n283_), .C(men_men_n279_), .Y(men_men_n288_));
  NO3        u266(.A(men_men_n288_), .B(men_men_n268_), .C(men_men_n255_), .Y(men_men_n289_));
  OAI210     u267(.A0(men_men_n206_), .A1(men_men_n54_), .B0(men_men_n289_), .Y(men02));
  AOI210     u268(.A0(men_men_n129_), .A1(men_men_n72_), .B0(men_men_n121_), .Y(men_men_n291_));
  NOi21      u269(.An(men_men_n235_), .B(men_men_n170_), .Y(men_men_n292_));
  NA3        u270(.A(x13), .B(men_men_n193_), .C(men_men_n49_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n292_), .A1(men_men_n30_), .B0(men_men_n293_), .Y(men_men_n294_));
  OAI210     u272(.A0(men_men_n294_), .A1(men_men_n291_), .B0(men_men_n167_), .Y(men_men_n295_));
  INV        u273(.A(men_men_n167_), .Y(men_men_n296_));
  AOI210     u274(.A0(men_men_n104_), .A1(men_men_n73_), .B0(men_men_n220_), .Y(men_men_n297_));
  OAI220     u275(.A0(men_men_n297_), .A1(men_men_n89_), .B0(men_men_n72_), .B1(men_men_n45_), .Y(men_men_n298_));
  AOI220     u276(.A0(men_men_n298_), .A1(men_men_n296_), .B0(men_men_n148_), .B1(men_men_n147_), .Y(men_men_n299_));
  AOI210     u277(.A0(men_men_n299_), .A1(men_men_n295_), .B0(men_men_n43_), .Y(men_men_n300_));
  NO2        u278(.A(x05), .B(x02), .Y(men_men_n301_));
  OAI210     u279(.A0(men_men_n210_), .A1(men_men_n191_), .B0(men_men_n301_), .Y(men_men_n302_));
  NOi21      u280(.An(x13), .B(men_men_n445_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n234_), .A1(men_men_n66_), .B0(men_men_n303_), .Y(men_men_n304_));
  AOI210     u282(.A0(men_men_n304_), .A1(men_men_n302_), .B0(men_men_n136_), .Y(men_men_n305_));
  NAi21      u283(.An(men_men_n236_), .B(men_men_n231_), .Y(men_men_n306_));
  NO2        u284(.A(men_men_n248_), .B(men_men_n42_), .Y(men_men_n307_));
  NA2        u285(.A(men_men_n307_), .B(men_men_n306_), .Y(men_men_n308_));
  AN2        u286(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n309_));
  OAI210     u287(.A0(men_men_n37_), .A1(men_men_n36_), .B0(men_men_n43_), .Y(men_men_n310_));
  NA2        u288(.A(x13), .B(men_men_n26_), .Y(men_men_n311_));
  OA210      u289(.A0(men_men_n311_), .A1(x08), .B0(men_men_n140_), .Y(men_men_n312_));
  AOI210     u290(.A0(men_men_n312_), .A1(men_men_n130_), .B0(men_men_n310_), .Y(men_men_n313_));
  OAI210     u291(.A0(men_men_n313_), .A1(men_men_n309_), .B0(men_men_n83_), .Y(men_men_n314_));
  NA3        u292(.A(men_men_n83_), .B(men_men_n71_), .C(men_men_n228_), .Y(men_men_n315_));
  NA3        u293(.A(men_men_n82_), .B(men_men_n70_), .C(men_men_n37_), .Y(men_men_n316_));
  AOI210     u294(.A0(men_men_n316_), .A1(men_men_n315_), .B0(x04), .Y(men_men_n317_));
  NO2        u295(.A(men_men_n262_), .B(men_men_n93_), .Y(men_men_n318_));
  AOI210     u296(.A0(men_men_n318_), .A1(x13), .B0(men_men_n317_), .Y(men_men_n319_));
  NA3        u297(.A(men_men_n319_), .B(men_men_n314_), .C(men_men_n308_), .Y(men_men_n320_));
  NO3        u298(.A(men_men_n320_), .B(men_men_n305_), .C(men_men_n300_), .Y(men_men_n321_));
  NA2        u299(.A(men_men_n135_), .B(x03), .Y(men_men_n322_));
  INV        u300(.A(men_men_n181_), .Y(men_men_n323_));
  OAI210     u301(.A0(men_men_n45_), .A1(men_men_n31_), .B0(men_men_n32_), .Y(men_men_n324_));
  AOI220     u302(.A0(men_men_n324_), .A1(men_men_n323_), .B0(men_men_n201_), .B1(x08), .Y(men_men_n325_));
  NO2        u303(.A(men_men_n325_), .B(men_men_n284_), .Y(men_men_n326_));
  NA2        u304(.A(men_men_n326_), .B(men_men_n95_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n166_), .B(men_men_n160_), .Y(men_men_n328_));
  AN2        u306(.A(men_men_n328_), .B(men_men_n173_), .Y(men_men_n329_));
  NO2        u307(.A(men_men_n275_), .B(x09), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n330_), .A1(men_men_n329_), .B0(men_men_n96_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n275_), .B(men_men_n88_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n88_), .B(men_men_n36_), .Y(men_men_n333_));
  NA3        u311(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n120_), .Y(men_men_n334_));
  NA4        u312(.A(men_men_n334_), .B(men_men_n331_), .C(men_men_n327_), .D(men_men_n43_), .Y(men_men_n335_));
  INV        u313(.A(men_men_n201_), .Y(men_men_n336_));
  NO2        u314(.A(men_men_n161_), .B(men_men_n35_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n30_), .B(x05), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n337_), .B0(men_men_n336_), .B1(men_men_n52_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n339_), .B(x02), .Y(men_men_n340_));
  INV        u318(.A(men_men_n241_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n198_), .B(x04), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  NO3        u321(.A(men_men_n183_), .B(x13), .C(men_men_n29_), .Y(men_men_n344_));
  OAI210     u322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n83_), .Y(men_men_n345_));
  NO3        u323(.A(men_men_n198_), .B(men_men_n159_), .C(men_men_n46_), .Y(men_men_n346_));
  OAI210     u324(.A0(men_men_n142_), .A1(men_men_n32_), .B0(men_men_n88_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NA4        u326(.A(men_men_n348_), .B(men_men_n345_), .C(men_men_n340_), .D(x06), .Y(men_men_n349_));
  NA2        u327(.A(x09), .B(x03), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n350_), .A1(men_men_n119_), .B0(men_men_n209_), .B1(men_men_n55_), .Y(men_men_n351_));
  OAI220     u329(.A0(men_men_n160_), .A1(x09), .B0(x08), .B1(men_men_n36_), .Y(men_men_n352_));
  NO3        u330(.A(men_men_n284_), .B(men_men_n118_), .C(x08), .Y(men_men_n353_));
  AOI210     u331(.A0(men_men_n352_), .A1(men_men_n227_), .B0(men_men_n353_), .Y(men_men_n354_));
  NO2        u332(.A(men_men_n43_), .B(men_men_n36_), .Y(men_men_n355_));
  NO3        u333(.A(men_men_n102_), .B(men_men_n119_), .C(men_men_n33_), .Y(men_men_n356_));
  AOI210     u334(.A0(men_men_n346_), .A1(men_men_n355_), .B0(men_men_n356_), .Y(men_men_n357_));
  OAI210     u335(.A0(men_men_n354_), .A1(men_men_n26_), .B0(men_men_n357_), .Y(men_men_n358_));
  AO220      u336(.A0(men_men_n358_), .A1(x04), .B0(men_men_n351_), .B1(x05), .Y(men_men_n359_));
  AOI210     u337(.A0(men_men_n349_), .A1(men_men_n335_), .B0(men_men_n359_), .Y(men_men_n360_));
  OAI210     u338(.A0(men_men_n321_), .A1(x12), .B0(men_men_n360_), .Y(men03));
  OR2        u339(.A(men_men_n37_), .B(men_men_n228_), .Y(men_men_n362_));
  AOI210     u340(.A0(men_men_n148_), .A1(men_men_n88_), .B0(men_men_n362_), .Y(men_men_n363_));
  AO210      u341(.A0(men_men_n341_), .A1(men_men_n73_), .B0(men_men_n342_), .Y(men_men_n364_));
  INV        u342(.A(men_men_n364_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n363_), .B0(x05), .Y(men_men_n366_));
  NA2        u344(.A(men_men_n362_), .B(x05), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n130_), .A1(men_men_n215_), .B0(men_men_n367_), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n230_), .A1(men_men_n67_), .B0(men_men_n112_), .Y(men_men_n369_));
  OAI220     u347(.A0(men_men_n369_), .A1(men_men_n52_), .B0(men_men_n311_), .B1(men_men_n445_), .Y(men_men_n370_));
  OAI210     u348(.A0(men_men_n370_), .A1(men_men_n368_), .B0(men_men_n88_), .Y(men_men_n371_));
  NO2        u349(.A(men_men_n333_), .B(men_men_n72_), .Y(men_men_n372_));
  INV        u350(.A(men_men_n372_), .Y(men_men_n373_));
  NA4        u351(.A(men_men_n373_), .B(men_men_n143_), .C(men_men_n371_), .D(men_men_n366_), .Y(men04));
  NO2        u352(.A(men_men_n76_), .B(men_men_n34_), .Y(men_men_n375_));
  XO2        u353(.A(men_men_n375_), .B(men_men_n251_), .Y(men05));
  AOI210     u354(.A0(men_men_n59_), .A1(men_men_n46_), .B0(men_men_n212_), .Y(men_men_n377_));
  AOI210     u355(.A0(men_men_n377_), .A1(men_men_n310_), .B0(men_men_n25_), .Y(men_men_n378_));
  NAi41      u356(.An(men_men_n65_), .B(men_men_n136_), .C(men_men_n121_), .D(men_men_n29_), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n233_), .A1(men_men_n50_), .B0(men_men_n77_), .Y(men_men_n380_));
  AOI210     u358(.A0(men_men_n380_), .A1(men_men_n379_), .B0(men_men_n24_), .Y(men_men_n381_));
  OAI210     u359(.A0(men_men_n381_), .A1(men_men_n378_), .B0(men_men_n88_), .Y(men_men_n382_));
  NA2        u360(.A(x11), .B(men_men_n29_), .Y(men_men_n383_));
  NA2        u361(.A(men_men_n23_), .B(men_men_n26_), .Y(men_men_n384_));
  NA2        u362(.A(men_men_n256_), .B(x03), .Y(men_men_n385_));
  OAI220     u363(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n383_), .B1(men_men_n68_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n386_), .A1(x06), .B0(men_men_n446_), .Y(men_men_n387_));
  AOI220     u365(.A0(men_men_n68_), .A1(men_men_n29_), .B0(men_men_n46_), .B1(men_men_n45_), .Y(men_men_n388_));
  NO3        u366(.A(men_men_n388_), .B(men_men_n23_), .C(x00), .Y(men_men_n389_));
  NA2        u367(.A(men_men_n58_), .B(x02), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n390_), .A1(men_men_n385_), .B0(men_men_n259_), .Y(men_men_n391_));
  OR2        u369(.A(men_men_n391_), .B(men_men_n240_), .Y(men_men_n392_));
  NA2        u370(.A(men_men_n155_), .B(x05), .Y(men_men_n393_));
  NA3        u371(.A(men_men_n393_), .B(men_men_n244_), .C(men_men_n239_), .Y(men_men_n394_));
  NO2        u372(.A(men_men_n23_), .B(x10), .Y(men_men_n395_));
  OAI210     u373(.A0(x11), .A1(men_men_n27_), .B0(men_men_n43_), .Y(men_men_n396_));
  OR3        u374(.A(men_men_n396_), .B(men_men_n395_), .C(men_men_n39_), .Y(men_men_n397_));
  NA3        u375(.A(men_men_n397_), .B(men_men_n394_), .C(men_men_n392_), .Y(men_men_n398_));
  OAI210     u376(.A0(men_men_n398_), .A1(men_men_n389_), .B0(men_men_n88_), .Y(men_men_n399_));
  INV        u377(.A(x07), .Y(men_men_n400_));
  AOI220     u378(.A0(men_men_n400_), .A1(men_men_n399_), .B0(men_men_n387_), .B1(men_men_n382_), .Y(men_men_n401_));
  NA3        u379(.A(men_men_n23_), .B(men_men_n54_), .C(men_men_n43_), .Y(men_men_n402_));
  AO210      u380(.A0(men_men_n402_), .A1(men_men_n269_), .B0(men_men_n266_), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n395_), .A1(men_men_n62_), .B0(men_men_n135_), .Y(men_men_n404_));
  OR2        u382(.A(men_men_n404_), .B(x03), .Y(men_men_n405_));
  NA2        u383(.A(men_men_n355_), .B(men_men_n54_), .Y(men_men_n406_));
  NO2        u384(.A(men_men_n406_), .B(x11), .Y(men_men_n407_));
  NO3        u385(.A(men_men_n407_), .B(men_men_n139_), .C(men_men_n26_), .Y(men_men_n408_));
  AOI220     u386(.A0(men_men_n408_), .A1(men_men_n405_), .B0(men_men_n403_), .B1(men_men_n42_), .Y(men_men_n409_));
  NO4        u387(.A(men_men_n333_), .B(men_men_n30_), .C(x11), .D(x09), .Y(men_men_n410_));
  OAI210     u388(.A0(men_men_n410_), .A1(men_men_n409_), .B0(men_men_n89_), .Y(men_men_n411_));
  NOi21      u389(.An(men_men_n322_), .B(men_men_n125_), .Y(men_men_n412_));
  NO2        u390(.A(men_men_n412_), .B(men_men_n266_), .Y(men_men_n413_));
  NO2        u391(.A(men_men_n413_), .B(x08), .Y(men_men_n414_));
  AOI210     u392(.A0(men_men_n395_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n415_));
  NA2        u393(.A(x09), .B(men_men_n36_), .Y(men_men_n416_));
  OAI220     u394(.A0(men_men_n416_), .A1(men_men_n415_), .B0(men_men_n383_), .B1(x06), .Y(men_men_n417_));
  NO2        u395(.A(x13), .B(x12), .Y(men_men_n418_));
  NO2        u396(.A(men_men_n121_), .B(men_men_n26_), .Y(men_men_n419_));
  NO2        u397(.A(men_men_n419_), .B(men_men_n270_), .Y(men_men_n420_));
  OR3        u398(.A(men_men_n420_), .B(x12), .C(x03), .Y(men_men_n421_));
  NA2        u399(.A(men_men_n421_), .B(x08), .Y(men_men_n422_));
  AOI210     u400(.A0(men_men_n418_), .A1(men_men_n417_), .B0(men_men_n422_), .Y(men_men_n423_));
  AOI210     u401(.A0(men_men_n414_), .A1(men_men_n411_), .B0(men_men_n423_), .Y(men_men_n424_));
  OAI210     u402(.A0(men_men_n406_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n425_));
  NA2        u403(.A(men_men_n296_), .B(x07), .Y(men_men_n426_));
  OAI220     u404(.A0(men_men_n426_), .A1(men_men_n384_), .B0(men_men_n139_), .B1(men_men_n38_), .Y(men_men_n427_));
  OAI210     u405(.A0(men_men_n427_), .A1(men_men_n425_), .B0(men_men_n187_), .Y(men_men_n428_));
  NA3        u406(.A(men_men_n420_), .B(men_men_n412_), .C(men_men_n332_), .Y(men_men_n429_));
  INV        u407(.A(x14), .Y(men_men_n430_));
  NO3        u408(.A(men_men_n322_), .B(men_men_n93_), .C(x11), .Y(men_men_n431_));
  NO3        u409(.A(men_men_n160_), .B(men_men_n62_), .C(men_men_n50_), .Y(men_men_n432_));
  NO3        u410(.A(men_men_n402_), .B(men_men_n333_), .C(men_men_n181_), .Y(men_men_n433_));
  NO4        u411(.A(men_men_n433_), .B(men_men_n432_), .C(men_men_n431_), .D(men_men_n430_), .Y(men_men_n434_));
  NA3        u412(.A(men_men_n434_), .B(men_men_n429_), .C(men_men_n428_), .Y(men_men_n435_));
  NA2        u413(.A(men_men_n419_), .B(men_men_n159_), .Y(men_men_n436_));
  NO3        u414(.A(men_men_n118_), .B(men_men_n24_), .C(x06), .Y(men_men_n437_));
  AOI210     u415(.A0(men_men_n282_), .A1(men_men_n233_), .B0(men_men_n437_), .Y(men_men_n438_));
  INV        u416(.A(men_men_n438_), .Y(men_men_n439_));
  NA2        u417(.A(men_men_n439_), .B(men_men_n88_), .Y(men_men_n440_));
  OAI210     u418(.A0(men_men_n436_), .A1(men_men_n78_), .B0(men_men_n440_), .Y(men_men_n441_));
  NO4        u419(.A(men_men_n441_), .B(men_men_n435_), .C(men_men_n424_), .D(men_men_n401_), .Y(men06));
  INV        u420(.A(men_men_n261_), .Y(men_men_n445_));
  INV        u421(.A(x07), .Y(men_men_n446_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule