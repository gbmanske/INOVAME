//Benchmark atmr_max1024_476_0.5

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n474_, men_men_n475_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  INV        o003(.A(ori_ori_n19_), .Y(ori_ori_n20_));
  NA2        o004(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n21_));
  INV        o005(.A(x5), .Y(ori_ori_n22_));
  INV        o006(.A(ori_ori_n21_), .Y(ori_ori_n23_));
  NO2        o007(.A(x4), .B(x3), .Y(ori_ori_n24_));
  INV        o008(.A(ori_ori_n24_), .Y(ori_ori_n25_));
  NOi21      o009(.An(ori_ori_n20_), .B(ori_ori_n23_), .Y(ori00));
  NO2        o010(.A(x1), .B(x0), .Y(ori_ori_n27_));
  INV        o011(.A(x6), .Y(ori_ori_n28_));
  NA2        o012(.A(x4), .B(x3), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n20_), .B(ori_ori_n29_), .Y(ori_ori_n30_));
  NO2        o014(.A(x2), .B(x0), .Y(ori_ori_n31_));
  INV        o015(.A(x3), .Y(ori_ori_n32_));
  NO2        o016(.A(ori_ori_n32_), .B(ori_ori_n18_), .Y(ori_ori_n33_));
  INV        o017(.A(ori_ori_n33_), .Y(ori_ori_n34_));
  INV        o018(.A(x4), .Y(ori_ori_n35_));
  OAI210     o019(.A0(ori_ori_n35_), .A1(ori_ori_n34_), .B0(ori_ori_n31_), .Y(ori_ori_n36_));
  INV        o020(.A(x4), .Y(ori_ori_n37_));
  INV        o021(.A(ori_ori_n36_), .Y(ori_ori_n38_));
  INV        o022(.A(ori_ori_n27_), .Y(ori_ori_n39_));
  INV        o023(.A(x2), .Y(ori_ori_n40_));
  NO2        o024(.A(ori_ori_n40_), .B(ori_ori_n17_), .Y(ori_ori_n41_));
  NA2        o025(.A(ori_ori_n32_), .B(ori_ori_n18_), .Y(ori_ori_n42_));
  NA2        o026(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  OAI210     o027(.A0(ori_ori_n39_), .A1(ori_ori_n25_), .B0(ori_ori_n43_), .Y(ori_ori_n44_));
  NO3        o028(.A(ori_ori_n44_), .B(ori_ori_n38_), .C(ori_ori_n30_), .Y(ori01));
  NA2        o029(.A(ori_ori_n32_), .B(x1), .Y(ori_ori_n46_));
  NO2        o030(.A(ori_ori_n46_), .B(x5), .Y(ori_ori_n47_));
  OAI210     o031(.A0(ori_ori_n33_), .A1(ori_ori_n22_), .B0(ori_ori_n40_), .Y(ori_ori_n48_));
  NA2        o032(.A(ori_ori_n42_), .B(ori_ori_n48_), .Y(ori_ori_n49_));
  INV        o033(.A(ori_ori_n49_), .Y(ori_ori_n50_));
  NA2        o034(.A(ori_ori_n50_), .B(x4), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n37_), .B(x2), .Y(ori_ori_n52_));
  OAI210     o036(.A0(ori_ori_n52_), .A1(ori_ori_n42_), .B0(x0), .Y(ori_ori_n53_));
  NAi21      o037(.An(x4), .B(x3), .Y(ori_ori_n54_));
  NO2        o038(.A(x4), .B(x2), .Y(ori_ori_n55_));
  NO2        o039(.A(ori_ori_n54_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NO2        o040(.A(ori_ori_n56_), .B(ori_ori_n53_), .Y(ori_ori_n57_));
  NA2        o041(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n58_));
  NO2        o042(.A(ori_ori_n58_), .B(ori_ori_n22_), .Y(ori_ori_n59_));
  AOI210     o043(.A0(ori_ori_n42_), .A1(ori_ori_n22_), .B0(ori_ori_n40_), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n34_), .B(ori_ori_n37_), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n62_));
  NA2        o046(.A(x4), .B(ori_ori_n32_), .Y(ori_ori_n63_));
  NO2        o047(.A(ori_ori_n37_), .B(ori_ori_n40_), .Y(ori_ori_n64_));
  NO2        o048(.A(ori_ori_n63_), .B(x1), .Y(ori_ori_n65_));
  NA2        o049(.A(ori_ori_n40_), .B(x1), .Y(ori_ori_n66_));
  OAI210     o050(.A0(ori_ori_n66_), .A1(ori_ori_n29_), .B0(ori_ori_n17_), .Y(ori_ori_n67_));
  NO3        o051(.A(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n62_), .Y(ori_ori_n68_));
  AO210      o052(.A0(ori_ori_n57_), .A1(ori_ori_n51_), .B0(ori_ori_n68_), .Y(ori02));
  NO2        o053(.A(x4), .B(x1), .Y(ori_ori_n70_));
  NO2        o054(.A(x5), .B(ori_ori_n37_), .Y(ori_ori_n71_));
  NO2        o055(.A(ori_ori_n55_), .B(ori_ori_n64_), .Y(ori_ori_n72_));
  NA2        o056(.A(x5), .B(x0), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n37_), .B(x2), .Y(ori_ori_n74_));
  NO2        o058(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n75_));
  NA2        o059(.A(ori_ori_n22_), .B(ori_ori_n18_), .Y(ori_ori_n76_));
  NA2        o060(.A(ori_ori_n22_), .B(ori_ori_n17_), .Y(ori_ori_n77_));
  NA3        o061(.A(ori_ori_n77_), .B(ori_ori_n76_), .C(ori_ori_n21_), .Y(ori_ori_n78_));
  AN2        o062(.A(ori_ori_n78_), .B(ori_ori_n74_), .Y(ori_ori_n79_));
  NA2        o063(.A(x2), .B(x0), .Y(ori_ori_n80_));
  NA2        o064(.A(x4), .B(x1), .Y(ori_ori_n81_));
  NAi21      o065(.An(ori_ori_n70_), .B(ori_ori_n81_), .Y(ori_ori_n82_));
  NOi21      o066(.An(ori_ori_n82_), .B(ori_ori_n80_), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n79_), .C(ori_ori_n75_), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n84_), .B(ori_ori_n32_), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n78_), .B(ori_ori_n52_), .Y(ori_ori_n86_));
  INV        o070(.A(ori_ori_n71_), .Y(ori_ori_n87_));
  NO2        o071(.A(ori_ori_n66_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  NA2        o072(.A(ori_ori_n82_), .B(ori_ori_n31_), .Y(ori_ori_n89_));
  OAI210     o073(.A0(ori_ori_n77_), .A1(ori_ori_n72_), .B0(ori_ori_n89_), .Y(ori_ori_n90_));
  NO3        o074(.A(ori_ori_n90_), .B(ori_ori_n88_), .C(ori_ori_n86_), .Y(ori_ori_n91_));
  NO2        o075(.A(ori_ori_n91_), .B(x3), .Y(ori_ori_n92_));
  NO2        o076(.A(ori_ori_n92_), .B(ori_ori_n85_), .Y(ori03));
  NO2        o077(.A(x0), .B(x6), .Y(ori_ori_n94_));
  NOi21      o078(.An(ori_ori_n55_), .B(ori_ori_n94_), .Y(ori_ori_n95_));
  INV        o079(.A(ori_ori_n95_), .Y(ori_ori_n96_));
  OR2        o080(.A(ori_ori_n96_), .B(x5), .Y(ori_ori_n97_));
  NA2        o081(.A(ori_ori_n74_), .B(ori_ori_n59_), .Y(ori_ori_n98_));
  NA2        o082(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n99_));
  NA3        o083(.A(ori_ori_n99_), .B(ori_ori_n98_), .C(ori_ori_n97_), .Y(ori_ori_n100_));
  INV        o084(.A(ori_ori_n100_), .Y(ori_ori_n101_));
  NA2        o085(.A(x3), .B(x2), .Y(ori_ori_n102_));
  INV        o086(.A(ori_ori_n33_), .Y(ori_ori_n103_));
  NO2        o087(.A(ori_ori_n103_), .B(ori_ori_n87_), .Y(ori_ori_n104_));
  NA2        o088(.A(x3), .B(x2), .Y(ori_ori_n105_));
  NAi21      o089(.An(x4), .B(x0), .Y(ori_ori_n106_));
  NO3        o090(.A(ori_ori_n106_), .B(ori_ori_n33_), .C(x2), .Y(ori_ori_n107_));
  INV        o091(.A(ori_ori_n107_), .Y(ori_ori_n108_));
  AOI220     o092(.A0(ori_ori_n17_), .A1(x3), .B0(ori_ori_n18_), .B1(ori_ori_n24_), .Y(ori_ori_n109_));
  AOI210     o093(.A0(ori_ori_n109_), .A1(ori_ori_n108_), .B0(ori_ori_n22_), .Y(ori_ori_n110_));
  NO2        o094(.A(ori_ori_n110_), .B(ori_ori_n104_), .Y(ori_ori_n111_));
  NA2        o095(.A(ori_ori_n101_), .B(ori_ori_n111_), .Y(ori04));
  INV        o096(.A(ori_ori_n106_), .Y(ori_ori_n113_));
  NO2        o097(.A(ori_ori_n40_), .B(ori_ori_n113_), .Y(ori_ori_n114_));
  NO2        o098(.A(ori_ori_n105_), .B(ori_ori_n135_), .Y(ori_ori_n115_));
  INV        o099(.A(ori_ori_n115_), .Y(ori_ori_n116_));
  NA2        o100(.A(ori_ori_n116_), .B(ori_ori_n114_), .Y(ori_ori_n117_));
  NA2        o101(.A(ori_ori_n117_), .B(x6), .Y(ori_ori_n118_));
  NA3        o102(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n119_), .B(x2), .Y(ori_ori_n120_));
  NA2        o104(.A(ori_ori_n120_), .B(x6), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n132_), .B(ori_ori_n40_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n122_), .B(ori_ori_n134_), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n123_), .B(ori_ori_n22_), .Y(ori_ori_n124_));
  NA2        o108(.A(ori_ori_n136_), .B(ori_ori_n102_), .Y(ori_ori_n125_));
  INV        o109(.A(ori_ori_n125_), .Y(ori_ori_n126_));
  OAI210     o110(.A0(ori_ori_n126_), .A1(ori_ori_n124_), .B0(ori_ori_n28_), .Y(ori_ori_n127_));
  NA2        o111(.A(ori_ori_n127_), .B(ori_ori_n121_), .Y(ori_ori_n128_));
  AOI210     o112(.A0(ori_ori_n133_), .A1(ori_ori_n22_), .B0(ori_ori_n128_), .Y(ori05));
  INV        o113(.A(x3), .Y(ori_ori_n132_));
  INV        o114(.A(ori_ori_n118_), .Y(ori_ori_n133_));
  INV        o115(.A(x0), .Y(ori_ori_n134_));
  INV        o116(.A(x0), .Y(ori_ori_n135_));
  INV        o117(.A(x0), .Y(ori_ori_n136_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  NAi21      m004(.An(mai_mai_n20_), .B(mai_mai_n19_), .Y(mai_mai_n21_));
  NA2        m005(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n22_));
  INV        m006(.A(x5), .Y(mai_mai_n23_));
  NA2        m007(.A(x7), .B(x6), .Y(mai_mai_n24_));
  NA2        m008(.A(x8), .B(x3), .Y(mai_mai_n25_));
  NA2        m009(.A(x4), .B(x2), .Y(mai_mai_n26_));
  NO4        m010(.A(mai_mai_n26_), .B(mai_mai_n25_), .C(mai_mai_n24_), .D(mai_mai_n23_), .Y(mai_mai_n27_));
  NO2        m011(.A(mai_mai_n27_), .B(mai_mai_n22_), .Y(mai_mai_n28_));
  NO2        m012(.A(x4), .B(x3), .Y(mai_mai_n29_));
  INV        m013(.A(mai_mai_n29_), .Y(mai_mai_n30_));
  OA210      m014(.A0(mai_mai_n30_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n31_));
  NOi31      m015(.An(mai_mai_n21_), .B(mai_mai_n31_), .C(mai_mai_n28_), .Y(mai00));
  NO2        m016(.A(x1), .B(x0), .Y(mai_mai_n33_));
  INV        m017(.A(x6), .Y(mai_mai_n34_));
  NA2        m018(.A(x4), .B(x3), .Y(mai_mai_n35_));
  AOI210     m019(.A0(mai_mai_n369_), .A1(mai_mai_n21_), .B0(mai_mai_n35_), .Y(mai_mai_n36_));
  NO2        m020(.A(x2), .B(x0), .Y(mai_mai_n37_));
  INV        m021(.A(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n39_));
  INV        m023(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(x5), .B(x4), .Y(mai_mai_n41_));
  OAI210     m025(.A0(mai_mai_n41_), .A1(mai_mai_n40_), .B0(mai_mai_n37_), .Y(mai_mai_n42_));
  INV        m026(.A(x4), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n44_));
  NA2        m028(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n45_));
  OAI210     m029(.A0(mai_mai_n45_), .A1(mai_mai_n20_), .B0(mai_mai_n42_), .Y(mai_mai_n46_));
  AOI220     m030(.A0(mai_mai_n23_), .A1(mai_mai_n33_), .B0(mai_mai_n20_), .B1(mai_mai_n19_), .Y(mai_mai_n47_));
  INV        m031(.A(x2), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n51_));
  OAI210     m035(.A0(mai_mai_n47_), .A1(mai_mai_n30_), .B0(mai_mai_n51_), .Y(mai_mai_n52_));
  NO3        m036(.A(mai_mai_n52_), .B(mai_mai_n46_), .C(mai_mai_n36_), .Y(mai01));
  NA2        m037(.A(x8), .B(x7), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n38_), .B(x1), .Y(mai_mai_n55_));
  INV        m039(.A(x9), .Y(mai_mai_n56_));
  NO2        m040(.A(mai_mai_n56_), .B(mai_mai_n34_), .Y(mai_mai_n57_));
  NO3        m041(.A(mai_mai_n34_), .B(mai_mai_n55_), .C(mai_mai_n54_), .Y(mai_mai_n58_));
  NO2        m042(.A(x7), .B(x6), .Y(mai_mai_n59_));
  NO2        m043(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n60_));
  NO2        m044(.A(x8), .B(x2), .Y(mai_mai_n61_));
  OA210      m045(.A0(mai_mai_n61_), .A1(mai_mai_n60_), .B0(mai_mai_n59_), .Y(mai_mai_n62_));
  OAI210     m046(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n48_), .Y(mai_mai_n63_));
  OAI210     m047(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n63_), .Y(mai_mai_n64_));
  NO2        m048(.A(mai_mai_n64_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n65_), .A1(mai_mai_n58_), .B0(x4), .Y(mai_mai_n66_));
  NA2        m050(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n67_));
  OAI210     m051(.A0(mai_mai_n67_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n68_));
  NA2        m052(.A(x5), .B(x3), .Y(mai_mai_n69_));
  NO2        m053(.A(x8), .B(x6), .Y(mai_mai_n70_));
  NO4        m054(.A(mai_mai_n70_), .B(mai_mai_n69_), .C(mai_mai_n59_), .D(mai_mai_n48_), .Y(mai_mai_n71_));
  NAi21      m055(.An(x4), .B(x3), .Y(mai_mai_n72_));
  INV        m056(.A(mai_mai_n72_), .Y(mai_mai_n73_));
  NO2        m057(.A(mai_mai_n73_), .B(mai_mai_n20_), .Y(mai_mai_n74_));
  NO2        m058(.A(x4), .B(x2), .Y(mai_mai_n75_));
  NO2        m059(.A(mai_mai_n75_), .B(x3), .Y(mai_mai_n76_));
  NO3        m060(.A(mai_mai_n76_), .B(mai_mai_n74_), .C(mai_mai_n18_), .Y(mai_mai_n77_));
  NO3        m061(.A(mai_mai_n77_), .B(mai_mai_n71_), .C(mai_mai_n68_), .Y(mai_mai_n78_));
  NO4        m062(.A(x7), .B(x6), .C(mai_mai_n38_), .D(x1), .Y(mai_mai_n79_));
  NA2        m063(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n80_), .B(mai_mai_n23_), .Y(mai_mai_n81_));
  INV        m065(.A(x8), .Y(mai_mai_n82_));
  NA2        m066(.A(x2), .B(x1), .Y(mai_mai_n83_));
  NO2        m067(.A(x2), .B(mai_mai_n81_), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(mai_mai_n24_), .Y(mai_mai_n85_));
  AOI210     m069(.A0(mai_mai_n50_), .A1(mai_mai_n23_), .B0(mai_mai_n48_), .Y(mai_mai_n86_));
  OAI210     m070(.A0(mai_mai_n40_), .A1(x5), .B0(mai_mai_n43_), .Y(mai_mai_n87_));
  NO3        m071(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(mai_mai_n85_), .Y(mai_mai_n88_));
  NA2        m072(.A(x4), .B(mai_mai_n38_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n43_), .B(mai_mai_n48_), .Y(mai_mai_n90_));
  OAI210     m074(.A0(mai_mai_n90_), .A1(mai_mai_n38_), .B0(mai_mai_n18_), .Y(mai_mai_n91_));
  AOI210     m075(.A0(mai_mai_n89_), .A1(mai_mai_n23_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NO2        m076(.A(x3), .B(x2), .Y(mai_mai_n93_));
  NA2        m077(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n94_));
  OAI210     m078(.A0(mai_mai_n94_), .A1(mai_mai_n35_), .B0(mai_mai_n17_), .Y(mai_mai_n95_));
  NO4        m079(.A(mai_mai_n95_), .B(mai_mai_n93_), .C(mai_mai_n92_), .D(mai_mai_n88_), .Y(mai_mai_n96_));
  AO220      m080(.A0(mai_mai_n96_), .A1(mai_mai_n368_), .B0(mai_mai_n78_), .B1(mai_mai_n66_), .Y(mai02));
  NO2        m081(.A(x3), .B(mai_mai_n48_), .Y(mai_mai_n98_));
  NA2        m082(.A(mai_mai_n38_), .B(x0), .Y(mai_mai_n99_));
  AOI220     m083(.A0(mai_mai_n43_), .A1(x1), .B0(mai_mai_n98_), .B1(x4), .Y(mai_mai_n100_));
  NO3        m084(.A(mai_mai_n100_), .B(x7), .C(x5), .Y(mai_mai_n101_));
  NA2        m085(.A(x9), .B(x2), .Y(mai_mai_n102_));
  OR2        m086(.A(x8), .B(x0), .Y(mai_mai_n103_));
  NAi21      m087(.An(x2), .B(x8), .Y(mai_mai_n104_));
  INV        m088(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m089(.A(x4), .B(x1), .Y(mai_mai_n106_));
  NA3        m090(.A(mai_mai_n106_), .B(x2), .C(mai_mai_n54_), .Y(mai_mai_n107_));
  NOi21      m091(.An(x0), .B(x1), .Y(mai_mai_n108_));
  NO3        m092(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n109_));
  NOi21      m093(.An(x0), .B(x4), .Y(mai_mai_n110_));
  NO2        m094(.A(x8), .B(mai_mai_n56_), .Y(mai_mai_n111_));
  AOI220     m095(.A0(mai_mai_n111_), .A1(mai_mai_n110_), .B0(mai_mai_n109_), .B1(mai_mai_n108_), .Y(mai_mai_n112_));
  AOI210     m096(.A0(mai_mai_n112_), .A1(mai_mai_n107_), .B0(mai_mai_n69_), .Y(mai_mai_n113_));
  NO2        m097(.A(x5), .B(mai_mai_n43_), .Y(mai_mai_n114_));
  NA2        m098(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n115_));
  AOI210     m099(.A0(mai_mai_n115_), .A1(mai_mai_n94_), .B0(mai_mai_n99_), .Y(mai_mai_n116_));
  OAI210     m100(.A0(mai_mai_n116_), .A1(mai_mai_n33_), .B0(mai_mai_n114_), .Y(mai_mai_n117_));
  NAi21      m101(.An(x0), .B(x4), .Y(mai_mai_n118_));
  NO2        m102(.A(mai_mai_n118_), .B(x1), .Y(mai_mai_n119_));
  NO2        m103(.A(x7), .B(x0), .Y(mai_mai_n120_));
  NO2        m104(.A(mai_mai_n75_), .B(mai_mai_n90_), .Y(mai_mai_n121_));
  NO2        m105(.A(mai_mai_n121_), .B(x3), .Y(mai_mai_n122_));
  OAI210     m106(.A0(mai_mai_n120_), .A1(mai_mai_n119_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NA2        m107(.A(x5), .B(x0), .Y(mai_mai_n124_));
  NO2        m108(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n125_));
  NA3        m109(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(x3), .Y(mai_mai_n126_));
  NA4        m110(.A(mai_mai_n126_), .B(mai_mai_n123_), .C(mai_mai_n117_), .D(mai_mai_n34_), .Y(mai_mai_n127_));
  NO3        m111(.A(mai_mai_n127_), .B(mai_mai_n113_), .C(mai_mai_n101_), .Y(mai_mai_n128_));
  NO3        m112(.A(mai_mai_n69_), .B(mai_mai_n67_), .C(mai_mai_n22_), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n26_), .B(mai_mai_n23_), .Y(mai_mai_n130_));
  AOI220     m114(.A0(mai_mai_n108_), .A1(mai_mai_n130_), .B0(mai_mai_n60_), .B1(mai_mai_n17_), .Y(mai_mai_n131_));
  NO3        m115(.A(mai_mai_n131_), .B(mai_mai_n54_), .C(mai_mai_n56_), .Y(mai_mai_n132_));
  NA2        m116(.A(x7), .B(x3), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n89_), .B(x5), .Y(mai_mai_n134_));
  NO2        m118(.A(x9), .B(x7), .Y(mai_mai_n135_));
  NOi21      m119(.An(x8), .B(x0), .Y(mai_mai_n136_));
  NO2        m120(.A(mai_mai_n38_), .B(x2), .Y(mai_mai_n137_));
  INV        m121(.A(x7), .Y(mai_mai_n138_));
  NA2        m122(.A(mai_mai_n138_), .B(mai_mai_n18_), .Y(mai_mai_n139_));
  AOI220     m123(.A0(mai_mai_n139_), .A1(mai_mai_n137_), .B0(mai_mai_n98_), .B1(x7), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n23_), .B(x4), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n141_), .B(mai_mai_n110_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n142_), .B(mai_mai_n140_), .Y(mai_mai_n143_));
  AOI210     m127(.A0(mai_mai_n136_), .A1(mai_mai_n134_), .B0(mai_mai_n143_), .Y(mai_mai_n144_));
  OAI210     m128(.A0(mai_mai_n133_), .A1(mai_mai_n45_), .B0(mai_mai_n144_), .Y(mai_mai_n145_));
  NA2        m129(.A(x5), .B(x1), .Y(mai_mai_n146_));
  INV        m130(.A(mai_mai_n146_), .Y(mai_mai_n147_));
  AOI210     m131(.A0(mai_mai_n147_), .A1(mai_mai_n110_), .B0(mai_mai_n34_), .Y(mai_mai_n148_));
  NAi31      m132(.An(mai_mai_n69_), .B(x7), .C(mai_mai_n33_), .Y(mai_mai_n149_));
  NA2        m133(.A(mai_mai_n149_), .B(mai_mai_n148_), .Y(mai_mai_n150_));
  NO4        m134(.A(mai_mai_n150_), .B(mai_mai_n145_), .C(mai_mai_n132_), .D(mai_mai_n129_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n151_), .B(mai_mai_n128_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n124_), .B(mai_mai_n121_), .Y(mai_mai_n153_));
  NA2        m137(.A(mai_mai_n23_), .B(mai_mai_n18_), .Y(mai_mai_n154_));
  NA2        m138(.A(mai_mai_n23_), .B(mai_mai_n17_), .Y(mai_mai_n155_));
  NA3        m139(.A(mai_mai_n155_), .B(mai_mai_n154_), .C(mai_mai_n22_), .Y(mai_mai_n156_));
  AN2        m140(.A(mai_mai_n156_), .B(mai_mai_n125_), .Y(mai_mai_n157_));
  NA2        m141(.A(x8), .B(x0), .Y(mai_mai_n158_));
  NO2        m142(.A(mai_mai_n138_), .B(mai_mai_n23_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n108_), .B(x4), .Y(mai_mai_n160_));
  NA2        m144(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  AOI210     m145(.A0(mai_mai_n158_), .A1(mai_mai_n115_), .B0(mai_mai_n161_), .Y(mai_mai_n162_));
  NA2        m146(.A(x2), .B(x0), .Y(mai_mai_n163_));
  NA2        m147(.A(x4), .B(x1), .Y(mai_mai_n164_));
  BUFFER     m148(.A(mai_mai_n106_), .Y(mai_mai_n165_));
  NOi31      m149(.An(mai_mai_n165_), .B(mai_mai_n141_), .C(mai_mai_n163_), .Y(mai_mai_n166_));
  NO4        m150(.A(mai_mai_n166_), .B(mai_mai_n162_), .C(mai_mai_n157_), .D(mai_mai_n153_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n167_), .B(mai_mai_n38_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n156_), .B(mai_mai_n67_), .Y(mai_mai_n169_));
  INV        m153(.A(mai_mai_n114_), .Y(mai_mai_n170_));
  NO3        m154(.A(mai_mai_n360_), .B(mai_mai_n170_), .C(x7), .Y(mai_mai_n171_));
  NO2        m155(.A(mai_mai_n155_), .B(mai_mai_n121_), .Y(mai_mai_n172_));
  NO3        m156(.A(mai_mai_n172_), .B(mai_mai_n171_), .C(mai_mai_n169_), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n173_), .B(x3), .Y(mai_mai_n174_));
  NO3        m158(.A(mai_mai_n174_), .B(mai_mai_n168_), .C(mai_mai_n152_), .Y(mai03));
  NO2        m159(.A(mai_mai_n43_), .B(x3), .Y(mai_mai_n176_));
  NO2        m160(.A(x6), .B(mai_mai_n23_), .Y(mai_mai_n177_));
  INV        m161(.A(mai_mai_n176_), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n69_), .B(x6), .Y(mai_mai_n179_));
  NA2        m163(.A(x6), .B(mai_mai_n23_), .Y(mai_mai_n180_));
  NO2        m164(.A(mai_mai_n180_), .B(x4), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n182_));
  AO220      m166(.A0(mai_mai_n182_), .A1(mai_mai_n181_), .B0(mai_mai_n179_), .B1(mai_mai_n49_), .Y(mai_mai_n183_));
  NA2        m167(.A(mai_mai_n183_), .B(mai_mai_n56_), .Y(mai_mai_n184_));
  NA2        m168(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n185_), .B(mai_mai_n180_), .Y(mai_mai_n186_));
  NA2        m170(.A(mai_mai_n180_), .B(mai_mai_n72_), .Y(mai_mai_n187_));
  AOI210     m171(.A0(mai_mai_n23_), .A1(x3), .B0(mai_mai_n163_), .Y(mai_mai_n188_));
  AOI220     m172(.A0(mai_mai_n188_), .A1(mai_mai_n187_), .B0(x9), .B1(mai_mai_n186_), .Y(mai_mai_n189_));
  NO2        m173(.A(x5), .B(x1), .Y(mai_mai_n190_));
  AOI220     m174(.A0(mai_mai_n190_), .A1(mai_mai_n17_), .B0(mai_mai_n93_), .B1(x5), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n185_), .B(mai_mai_n154_), .Y(mai_mai_n192_));
  NO3        m176(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n193_), .B(mai_mai_n192_), .Y(mai_mai_n194_));
  OAI210     m178(.A0(mai_mai_n191_), .A1(mai_mai_n34_), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  NA2        m179(.A(mai_mai_n195_), .B(mai_mai_n43_), .Y(mai_mai_n196_));
  NA4        m180(.A(mai_mai_n196_), .B(mai_mai_n189_), .C(mai_mai_n184_), .D(mai_mai_n178_), .Y(mai_mai_n197_));
  NO2        m181(.A(mai_mai_n43_), .B(mai_mai_n38_), .Y(mai_mai_n198_));
  NO2        m182(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n199_));
  NO2        m183(.A(mai_mai_n199_), .B(x6), .Y(mai_mai_n200_));
  NA2        m184(.A(mai_mai_n56_), .B(mai_mai_n82_), .Y(mai_mai_n201_));
  NA2        m185(.A(mai_mai_n38_), .B(mai_mai_n48_), .Y(mai_mai_n202_));
  NO2        m186(.A(mai_mai_n202_), .B(mai_mai_n23_), .Y(mai_mai_n203_));
  NO3        m187(.A(mai_mai_n164_), .B(mai_mai_n56_), .C(x6), .Y(mai_mai_n204_));
  AOI220     m188(.A0(mai_mai_n204_), .A1(mai_mai_n203_), .B0(mai_mai_n125_), .B1(mai_mai_n81_), .Y(mai_mai_n205_));
  NA2        m189(.A(x6), .B(mai_mai_n43_), .Y(mai_mai_n206_));
  AOI210     m190(.A0(mai_mai_n365_), .A1(mai_mai_n206_), .B0(mai_mai_n69_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n146_), .B(mai_mai_n38_), .Y(mai_mai_n208_));
  NO2        m192(.A(mai_mai_n208_), .B(mai_mai_n192_), .Y(mai_mai_n209_));
  NA2        m193(.A(mai_mai_n177_), .B(mai_mai_n119_), .Y(mai_mai_n210_));
  NA3        m194(.A(mai_mai_n185_), .B(mai_mai_n114_), .C(x6), .Y(mai_mai_n211_));
  NA3        m195(.A(mai_mai_n211_), .B(mai_mai_n210_), .C(mai_mai_n209_), .Y(mai_mai_n212_));
  OAI210     m196(.A0(mai_mai_n212_), .A1(mai_mai_n207_), .B0(x2), .Y(mai_mai_n213_));
  NA3        m197(.A(mai_mai_n213_), .B(mai_mai_n205_), .C(x7), .Y(mai_mai_n214_));
  AOI210     m198(.A0(mai_mai_n197_), .A1(x8), .B0(mai_mai_n214_), .Y(mai_mai_n215_));
  NA2        m199(.A(mai_mai_n200_), .B(mai_mai_n141_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n216_), .B(x2), .Y(mai_mai_n217_));
  NO2        m201(.A(x4), .B(mai_mai_n48_), .Y(mai_mai_n218_));
  NA2        m202(.A(mai_mai_n218_), .B(mai_mai_n60_), .Y(mai_mai_n219_));
  NA2        m203(.A(mai_mai_n56_), .B(x6), .Y(mai_mai_n220_));
  NA3        m204(.A(mai_mai_n23_), .B(x3), .C(x2), .Y(mai_mai_n221_));
  AOI210     m205(.A0(mai_mai_n221_), .A1(mai_mai_n124_), .B0(mai_mai_n220_), .Y(mai_mai_n222_));
  NA2        m206(.A(mai_mai_n38_), .B(mai_mai_n17_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n222_), .B(mai_mai_n106_), .Y(mai_mai_n224_));
  NO2        m208(.A(mai_mai_n185_), .B(x6), .Y(mai_mai_n225_));
  NA3        m209(.A(mai_mai_n185_), .B(mai_mai_n361_), .C(mai_mai_n130_), .Y(mai_mai_n226_));
  NA4        m210(.A(mai_mai_n226_), .B(mai_mai_n224_), .C(mai_mai_n219_), .D(mai_mai_n138_), .Y(mai_mai_n227_));
  NA2        m211(.A(mai_mai_n177_), .B(mai_mai_n199_), .Y(mai_mai_n228_));
  NO2        m212(.A(mai_mai_n124_), .B(mai_mai_n18_), .Y(mai_mai_n229_));
  NAi21      m213(.An(mai_mai_n229_), .B(mai_mai_n221_), .Y(mai_mai_n230_));
  NAi21      m214(.An(x1), .B(x4), .Y(mai_mai_n231_));
  AOI210     m215(.A0(x3), .A1(x2), .B0(mai_mai_n43_), .Y(mai_mai_n232_));
  OAI210     m216(.A0(mai_mai_n124_), .A1(x3), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  AOI210     m217(.A0(mai_mai_n233_), .A1(mai_mai_n231_), .B0(mai_mai_n230_), .Y(mai_mai_n234_));
  NA2        m218(.A(mai_mai_n234_), .B(mai_mai_n228_), .Y(mai_mai_n235_));
  NA2        m219(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n236_));
  NO2        m220(.A(mai_mai_n236_), .B(mai_mai_n228_), .Y(mai_mai_n237_));
  NO3        m221(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n238_));
  NA2        m222(.A(x6), .B(x2), .Y(mai_mai_n239_));
  NO2        m223(.A(mai_mai_n239_), .B(mai_mai_n154_), .Y(mai_mai_n240_));
  AOI210     m224(.A0(mai_mai_n48_), .A1(mai_mai_n238_), .B0(mai_mai_n240_), .Y(mai_mai_n241_));
  OAI220     m225(.A0(mai_mai_n241_), .A1(mai_mai_n38_), .B0(mai_mai_n160_), .B1(mai_mai_n41_), .Y(mai_mai_n242_));
  OAI210     m226(.A0(mai_mai_n242_), .A1(mai_mai_n237_), .B0(mai_mai_n235_), .Y(mai_mai_n243_));
  NA2        m227(.A(x4), .B(x0), .Y(mai_mai_n244_));
  NA2        m228(.A(mai_mai_n134_), .B(mai_mai_n37_), .Y(mai_mai_n245_));
  AOI210     m229(.A0(mai_mai_n245_), .A1(mai_mai_n243_), .B0(x8), .Y(mai_mai_n246_));
  OAI210     m230(.A0(mai_mai_n229_), .A1(mai_mai_n190_), .B0(x6), .Y(mai_mai_n247_));
  AOI210     m231(.A0(mai_mai_n370_), .A1(mai_mai_n247_), .B0(mai_mai_n202_), .Y(mai_mai_n248_));
  NO4        m232(.A(mai_mai_n248_), .B(mai_mai_n246_), .C(mai_mai_n227_), .D(mai_mai_n217_), .Y(mai_mai_n249_));
  OAI210     m233(.A0(x6), .A1(mai_mai_n225_), .B0(x2), .Y(mai_mai_n250_));
  NA2        m234(.A(x6), .B(mai_mai_n39_), .Y(mai_mai_n251_));
  AOI210     m235(.A0(mai_mai_n251_), .A1(mai_mai_n250_), .B0(mai_mai_n170_), .Y(mai_mai_n252_));
  NOi21      m236(.An(mai_mai_n239_), .B(mai_mai_n17_), .Y(mai_mai_n253_));
  NA3        m237(.A(mai_mai_n253_), .B(mai_mai_n190_), .C(mai_mai_n35_), .Y(mai_mai_n254_));
  AOI210     m238(.A0(mai_mai_n34_), .A1(mai_mai_n48_), .B0(x0), .Y(mai_mai_n255_));
  NA3        m239(.A(mai_mai_n255_), .B(mai_mai_n147_), .C(mai_mai_n30_), .Y(mai_mai_n256_));
  NA2        m240(.A(x3), .B(x2), .Y(mai_mai_n257_));
  AOI220     m241(.A0(mai_mai_n257_), .A1(mai_mai_n202_), .B0(mai_mai_n256_), .B1(mai_mai_n254_), .Y(mai_mai_n258_));
  NAi21      m242(.An(x4), .B(x0), .Y(mai_mai_n259_));
  NO3        m243(.A(mai_mai_n259_), .B(mai_mai_n39_), .C(x2), .Y(mai_mai_n260_));
  NO2        m244(.A(x9), .B(x8), .Y(mai_mai_n261_));
  NA2        m245(.A(x0), .B(mai_mai_n73_), .Y(mai_mai_n262_));
  NO2        m246(.A(mai_mai_n262_), .B(mai_mai_n23_), .Y(mai_mai_n263_));
  NA3        m247(.A(mai_mai_n34_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n264_));
  OAI210     m248(.A0(mai_mai_n255_), .A1(mai_mai_n253_), .B0(mai_mai_n264_), .Y(mai_mai_n265_));
  INV        m249(.A(mai_mai_n192_), .Y(mai_mai_n266_));
  NA2        m250(.A(mai_mai_n34_), .B(mai_mai_n38_), .Y(mai_mai_n267_));
  OR2        m251(.A(mai_mai_n267_), .B(mai_mai_n244_), .Y(mai_mai_n268_));
  OAI220     m252(.A0(mai_mai_n268_), .A1(mai_mai_n146_), .B0(mai_mai_n206_), .B1(mai_mai_n266_), .Y(mai_mai_n269_));
  AO210      m253(.A0(mai_mai_n265_), .A1(mai_mai_n134_), .B0(mai_mai_n269_), .Y(mai_mai_n270_));
  NO4        m254(.A(mai_mai_n270_), .B(mai_mai_n263_), .C(mai_mai_n258_), .D(mai_mai_n252_), .Y(mai_mai_n271_));
  OAI210     m255(.A0(mai_mai_n249_), .A1(mai_mai_n215_), .B0(mai_mai_n271_), .Y(mai04));
  NO2        m256(.A(mai_mai_n236_), .B(mai_mai_n80_), .Y(mai_mai_n273_));
  NO2        m257(.A(mai_mai_n273_), .B(mai_mai_n34_), .Y(mai_mai_n274_));
  NO2        m258(.A(mai_mai_n257_), .B(mai_mai_n182_), .Y(mai_mai_n275_));
  NA2        m259(.A(mai_mai_n275_), .B(mai_mai_n82_), .Y(mai_mai_n276_));
  NA2        m260(.A(mai_mai_n276_), .B(mai_mai_n274_), .Y(mai_mai_n277_));
  NA2        m261(.A(mai_mai_n277_), .B(x6), .Y(mai_mai_n278_));
  NOi21      m262(.An(mai_mai_n136_), .B(mai_mai_n115_), .Y(mai_mai_n279_));
  AOI210     m263(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n280_));
  OAI220     m264(.A0(mai_mai_n280_), .A1(mai_mai_n267_), .B0(mai_mai_n236_), .B1(mai_mai_n264_), .Y(mai_mai_n281_));
  AOI210     m265(.A0(mai_mai_n279_), .A1(mai_mai_n57_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n94_), .A1(mai_mai_n17_), .B0(mai_mai_n366_), .Y(mai_mai_n283_));
  AOI220     m267(.A0(mai_mai_n283_), .A1(mai_mai_n70_), .B0(mai_mai_n273_), .B1(mai_mai_n82_), .Y(mai_mai_n284_));
  NA2        m268(.A(mai_mai_n284_), .B(mai_mai_n282_), .Y(mai_mai_n285_));
  OAI210     m269(.A0(x1), .A1(x3), .B0(mai_mai_n260_), .Y(mai_mai_n286_));
  NA2        m270(.A(mai_mai_n286_), .B(mai_mai_n138_), .Y(mai_mai_n287_));
  AOI210     m271(.A0(mai_mai_n285_), .A1(x4), .B0(mai_mai_n287_), .Y(mai_mai_n288_));
  NOi21      m272(.An(x4), .B(x0), .Y(mai_mai_n289_));
  XO2        m273(.A(x4), .B(x0), .Y(mai_mai_n290_));
  OAI210     m274(.A0(mai_mai_n290_), .A1(mai_mai_n102_), .B0(mai_mai_n231_), .Y(mai_mai_n291_));
  AOI220     m275(.A0(mai_mai_n291_), .A1(x8), .B0(mai_mai_n289_), .B1(mai_mai_n83_), .Y(mai_mai_n292_));
  NO2        m276(.A(mai_mai_n292_), .B(x3), .Y(mai_mai_n293_));
  NO2        m277(.A(mai_mai_n82_), .B(x4), .Y(mai_mai_n294_));
  NA2        m278(.A(mai_mai_n294_), .B(mai_mai_n39_), .Y(mai_mai_n295_));
  NO3        m279(.A(mai_mai_n201_), .B(mai_mai_n26_), .C(mai_mai_n22_), .Y(mai_mai_n296_));
  INV        m280(.A(mai_mai_n296_), .Y(mai_mai_n297_));
  NA3        m281(.A(mai_mai_n297_), .B(mai_mai_n295_), .C(x6), .Y(mai_mai_n298_));
  NO2        m282(.A(mai_mai_n136_), .B(mai_mai_n72_), .Y(mai_mai_n299_));
  NO2        m283(.A(mai_mai_n33_), .B(x2), .Y(mai_mai_n300_));
  NOi21      m284(.An(mai_mai_n106_), .B(mai_mai_n25_), .Y(mai_mai_n301_));
  AOI210     m285(.A0(mai_mai_n300_), .A1(mai_mai_n299_), .B0(mai_mai_n301_), .Y(mai_mai_n302_));
  OAI210     m286(.A0(mai_mai_n363_), .A1(mai_mai_n56_), .B0(mai_mai_n302_), .Y(mai_mai_n303_));
  OAI220     m287(.A0(mai_mai_n303_), .A1(x6), .B0(mai_mai_n298_), .B1(mai_mai_n293_), .Y(mai_mai_n304_));
  INV        m288(.A(mai_mai_n268_), .Y(mai_mai_n305_));
  AOI210     m289(.A0(mai_mai_n305_), .A1(mai_mai_n18_), .B0(mai_mai_n138_), .Y(mai_mai_n306_));
  AO220      m290(.A0(mai_mai_n306_), .A1(mai_mai_n304_), .B0(mai_mai_n288_), .B1(mai_mai_n278_), .Y(mai_mai_n307_));
  NA2        m291(.A(mai_mai_n300_), .B(x6), .Y(mai_mai_n308_));
  NA2        m292(.A(mai_mai_n294_), .B(x0), .Y(mai_mai_n309_));
  NA2        m293(.A(mai_mai_n75_), .B(x6), .Y(mai_mai_n310_));
  OAI210     m294(.A0(mai_mai_n309_), .A1(mai_mai_n367_), .B0(mai_mai_n310_), .Y(mai_mai_n311_));
  AOI220     m295(.A0(mai_mai_n311_), .A1(mai_mai_n308_), .B0(mai_mai_n193_), .B1(mai_mai_n44_), .Y(mai_mai_n312_));
  NA2        m296(.A(mai_mai_n312_), .B(mai_mai_n307_), .Y(mai_mai_n313_));
  NA3        m297(.A(mai_mai_n105_), .B(mai_mai_n198_), .C(x0), .Y(mai_mai_n314_));
  AOI210     m298(.A0(mai_mai_n104_), .A1(mai_mai_n103_), .B0(mai_mai_n37_), .Y(mai_mai_n315_));
  NOi31      m299(.An(mai_mai_n315_), .B(x3), .C(mai_mai_n164_), .Y(mai_mai_n316_));
  OAI210     m300(.A0(mai_mai_n316_), .A1(x5), .B0(mai_mai_n135_), .Y(mai_mai_n317_));
  NA3        m301(.A(mai_mai_n23_), .B(mai_mai_n317_), .C(mai_mai_n314_), .Y(mai_mai_n318_));
  OAI210     m302(.A0(mai_mai_n318_), .A1(x5), .B0(x6), .Y(mai_mai_n319_));
  NA3        m303(.A(mai_mai_n49_), .B(x7), .C(mai_mai_n29_), .Y(mai_mai_n320_));
  NO2        m304(.A(mai_mai_n320_), .B(mai_mai_n30_), .Y(mai_mai_n321_));
  NA2        m305(.A(mai_mai_n176_), .B(mai_mai_n138_), .Y(mai_mai_n322_));
  AOI210     m306(.A0(mai_mai_n111_), .A1(mai_mai_n218_), .B0(x1), .Y(mai_mai_n323_));
  OAI210     m307(.A0(mai_mai_n322_), .A1(x8), .B0(mai_mai_n323_), .Y(mai_mai_n324_));
  NA3        m308(.A(x0), .B(mai_mai_n133_), .C(x9), .Y(mai_mai_n325_));
  NO4        m309(.A(x8), .B(mai_mai_n259_), .C(x9), .D(x2), .Y(mai_mai_n326_));
  NOi21      m310(.An(mai_mai_n109_), .B(mai_mai_n163_), .Y(mai_mai_n327_));
  NO3        m311(.A(mai_mai_n327_), .B(mai_mai_n326_), .C(mai_mai_n18_), .Y(mai_mai_n328_));
  NA2        m312(.A(mai_mai_n299_), .B(mai_mai_n138_), .Y(mai_mai_n329_));
  NA4        m313(.A(mai_mai_n329_), .B(mai_mai_n328_), .C(mai_mai_n325_), .D(mai_mai_n45_), .Y(mai_mai_n330_));
  OAI210     m314(.A0(mai_mai_n324_), .A1(mai_mai_n321_), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  NO2        m315(.A(mai_mai_n109_), .B(mai_mai_n38_), .Y(mai_mai_n332_));
  NO3        m316(.A(mai_mai_n364_), .B(mai_mai_n332_), .C(x2), .Y(mai_mai_n333_));
  OAI220     m317(.A0(mai_mai_n290_), .A1(mai_mai_n261_), .B0(mai_mai_n259_), .B1(mai_mai_n38_), .Y(mai_mai_n334_));
  NA2        m318(.A(mai_mai_n334_), .B(mai_mai_n138_), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n335_), .B(mai_mai_n48_), .Y(mai_mai_n336_));
  NO2        m320(.A(mai_mai_n336_), .B(mai_mai_n333_), .Y(mai_mai_n337_));
  AOI210     m321(.A0(mai_mai_n337_), .A1(mai_mai_n331_), .B0(mai_mai_n23_), .Y(mai_mai_n338_));
  NA2        m322(.A(mai_mai_n359_), .B(mai_mai_n315_), .Y(mai_mai_n339_));
  NO2        m323(.A(mai_mai_n339_), .B(mai_mai_n93_), .Y(mai_mai_n340_));
  NO3        m324(.A(mai_mai_n236_), .B(mai_mai_n158_), .C(mai_mai_n35_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n341_), .A1(mai_mai_n340_), .B0(x7), .Y(mai_mai_n342_));
  INV        m326(.A(mai_mai_n342_), .Y(mai_mai_n343_));
  OAI210     m327(.A0(mai_mai_n343_), .A1(mai_mai_n338_), .B0(mai_mai_n34_), .Y(mai_mai_n344_));
  INV        m328(.A(mai_mai_n182_), .Y(mai_mai_n345_));
  NO4        m329(.A(mai_mai_n345_), .B(mai_mai_n69_), .C(x4), .D(mai_mai_n48_), .Y(mai_mai_n346_));
  NA2        m330(.A(mai_mai_n223_), .B(x7), .Y(mai_mai_n347_));
  NO2        m331(.A(mai_mai_n146_), .B(mai_mai_n120_), .Y(mai_mai_n348_));
  NA2        m332(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  AOI210     m333(.A0(mai_mai_n349_), .A1(mai_mai_n149_), .B0(mai_mai_n26_), .Y(mai_mai_n350_));
  AOI210     m334(.A0(mai_mai_n362_), .A1(mai_mai_n23_), .B0(mai_mai_n206_), .Y(mai_mai_n351_));
  NA2        m335(.A(x9), .B(x5), .Y(mai_mai_n352_));
  NO4        m336(.A(mai_mai_n94_), .B(mai_mai_n352_), .C(mai_mai_n54_), .D(mai_mai_n30_), .Y(mai_mai_n353_));
  NO4        m337(.A(mai_mai_n353_), .B(mai_mai_n351_), .C(mai_mai_n350_), .D(mai_mai_n346_), .Y(mai_mai_n354_));
  NA3        m338(.A(mai_mai_n354_), .B(mai_mai_n344_), .C(mai_mai_n319_), .Y(mai_mai_n355_));
  AOI210     m339(.A0(mai_mai_n313_), .A1(mai_mai_n23_), .B0(mai_mai_n355_), .Y(mai05));
  INV        m340(.A(x4), .Y(mai_mai_n359_));
  INV        m341(.A(mai_mai_n33_), .Y(mai_mai_n360_));
  INV        m342(.A(x6), .Y(mai_mai_n361_));
  INV        m343(.A(x5), .Y(mai_mai_n362_));
  INV        m344(.A(x0), .Y(mai_mai_n363_));
  INV        m345(.A(x0), .Y(mai_mai_n364_));
  INV        m346(.A(x0), .Y(mai_mai_n365_));
  INV        m347(.A(x2), .Y(mai_mai_n366_));
  INV        m348(.A(x1), .Y(mai_mai_n367_));
  INV        m349(.A(mai_mai_n79_), .Y(mai_mai_n368_));
  INV        m350(.A(mai_mai_n33_), .Y(mai_mai_n369_));
  INV        m351(.A(x4), .Y(mai_mai_n370_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO2        u012(.A(x4), .B(men_men_n24_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n23_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n25_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA3        u020(.A(men_men_n36_), .B(men_men_n35_), .C(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n23_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n35_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n50_));
  AOI220     u034(.A0(men_men_n50_), .A1(men_men_n33_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  INV        u037(.A(men_men_n53_), .Y(men_men_n54_));
  OAI210     u038(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n54_), .Y(men_men_n55_));
  NO3        u039(.A(men_men_n55_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u040(.A(x8), .B(x7), .Y(men_men_n57_));
  NA2        u041(.A(men_men_n41_), .B(x1), .Y(men_men_n58_));
  INV        u042(.A(x9), .Y(men_men_n59_));
  NO2        u043(.A(men_men_n59_), .B(men_men_n34_), .Y(men_men_n60_));
  INV        u044(.A(men_men_n60_), .Y(men_men_n61_));
  NO2        u045(.A(x7), .B(x6), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n58_), .B(x5), .Y(men_men_n63_));
  NO2        u047(.A(x8), .B(x2), .Y(men_men_n64_));
  INV        u048(.A(men_men_n64_), .Y(men_men_n65_));
  NO2        u049(.A(men_men_n65_), .B(x1), .Y(men_men_n66_));
  OA210      u050(.A0(men_men_n66_), .A1(men_men_n63_), .B0(men_men_n62_), .Y(men_men_n67_));
  OAI210     u051(.A0(men_men_n42_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n68_));
  INV        u052(.A(men_men_n68_), .Y(men_men_n69_));
  NAi31      u053(.An(x1), .B(x9), .C(x5), .Y(men_men_n70_));
  OAI220     u054(.A0(men_men_n70_), .A1(men_men_n41_), .B0(men_men_n69_), .B1(men_men_n67_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n71_), .A1(men_men_n60_), .B0(x4), .Y(men_men_n72_));
  NA2        u056(.A(men_men_n46_), .B(x2), .Y(men_men_n73_));
  INV        u057(.A(x0), .Y(men_men_n74_));
  NA2        u058(.A(x5), .B(x3), .Y(men_men_n75_));
  NO2        u059(.A(x8), .B(x6), .Y(men_men_n76_));
  NO4        u060(.A(men_men_n76_), .B(men_men_n75_), .C(men_men_n62_), .D(men_men_n52_), .Y(men_men_n77_));
  NAi21      u061(.An(x4), .B(x3), .Y(men_men_n78_));
  INV        u062(.A(men_men_n78_), .Y(men_men_n79_));
  NO2        u063(.A(x4), .B(x2), .Y(men_men_n80_));
  NO2        u064(.A(men_men_n80_), .B(x3), .Y(men_men_n81_));
  NO3        u065(.A(men_men_n81_), .B(men_men_n21_), .C(men_men_n18_), .Y(men_men_n82_));
  NO3        u066(.A(men_men_n82_), .B(men_men_n77_), .C(men_men_n74_), .Y(men_men_n83_));
  NO4        u067(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n84_));
  NA2        u068(.A(men_men_n59_), .B(men_men_n46_), .Y(men_men_n85_));
  INV        u069(.A(men_men_n85_), .Y(men_men_n86_));
  OAI210     u070(.A0(men_men_n84_), .A1(men_men_n63_), .B0(men_men_n86_), .Y(men_men_n87_));
  NA2        u071(.A(x3), .B(men_men_n18_), .Y(men_men_n88_));
  NO2        u072(.A(men_men_n88_), .B(men_men_n25_), .Y(men_men_n89_));
  INV        u073(.A(x8), .Y(men_men_n90_));
  NA2        u074(.A(x2), .B(x1), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n89_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n26_), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n25_), .B(men_men_n52_), .Y(men_men_n95_));
  OAI210     u079(.A0(men_men_n43_), .A1(men_men_n35_), .B0(men_men_n46_), .Y(men_men_n96_));
  NO3        u080(.A(men_men_n96_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n97_));
  NA2        u081(.A(x4), .B(men_men_n41_), .Y(men_men_n98_));
  NO2        u082(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n99_));
  NO2        u083(.A(men_men_n50_), .B(men_men_n52_), .Y(men_men_n100_));
  NO2        u084(.A(x3), .B(x2), .Y(men_men_n101_));
  NA3        u085(.A(men_men_n101_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n102_));
  AOI210     u086(.A0(x8), .A1(x6), .B0(men_men_n102_), .Y(men_men_n103_));
  NA2        u087(.A(men_men_n52_), .B(x1), .Y(men_men_n104_));
  NO4        u088(.A(x0), .B(men_men_n103_), .C(men_men_n100_), .D(men_men_n97_), .Y(men_men_n105_));
  AO220      u089(.A0(men_men_n105_), .A1(men_men_n87_), .B0(men_men_n83_), .B1(men_men_n72_), .Y(men02));
  NO2        u090(.A(x3), .B(men_men_n52_), .Y(men_men_n107_));
  NO2        u091(.A(x8), .B(men_men_n18_), .Y(men_men_n108_));
  NA2        u092(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n109_));
  NA2        u093(.A(men_men_n41_), .B(x0), .Y(men_men_n110_));
  OAI210     u094(.A0(men_men_n85_), .A1(men_men_n109_), .B0(men_men_n110_), .Y(men_men_n111_));
  AOI220     u095(.A0(men_men_n111_), .A1(men_men_n108_), .B0(men_men_n107_), .B1(x4), .Y(men_men_n112_));
  NO3        u096(.A(men_men_n112_), .B(x7), .C(x5), .Y(men_men_n113_));
  NA2        u097(.A(x9), .B(x2), .Y(men_men_n114_));
  OR2        u098(.A(x8), .B(x0), .Y(men_men_n115_));
  INV        u099(.A(men_men_n115_), .Y(men_men_n116_));
  NAi21      u100(.An(x2), .B(x8), .Y(men_men_n117_));
  INV        u101(.A(men_men_n117_), .Y(men_men_n118_));
  OAI220     u102(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n114_), .B1(x7), .Y(men_men_n119_));
  NO2        u103(.A(x4), .B(x1), .Y(men_men_n120_));
  NA3        u104(.A(men_men_n120_), .B(men_men_n119_), .C(men_men_n57_), .Y(men_men_n121_));
  NOi21      u105(.An(x0), .B(x1), .Y(men_men_n122_));
  NO3        u106(.A(x9), .B(x8), .C(x7), .Y(men_men_n123_));
  NOi21      u107(.An(x0), .B(x4), .Y(men_men_n124_));
  NAi21      u108(.An(x8), .B(x7), .Y(men_men_n125_));
  NO2        u109(.A(men_men_n125_), .B(men_men_n59_), .Y(men_men_n126_));
  AOI220     u110(.A0(men_men_n126_), .A1(men_men_n124_), .B0(men_men_n123_), .B1(men_men_n122_), .Y(men_men_n127_));
  AOI210     u111(.A0(men_men_n127_), .A1(men_men_n121_), .B0(men_men_n75_), .Y(men_men_n128_));
  NO2        u112(.A(x5), .B(men_men_n46_), .Y(men_men_n129_));
  OAI210     u113(.A0(men_men_n18_), .A1(men_men_n33_), .B0(men_men_n129_), .Y(men_men_n130_));
  NAi21      u114(.An(x0), .B(x4), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n131_), .B(x1), .Y(men_men_n132_));
  NO2        u116(.A(x7), .B(x0), .Y(men_men_n133_));
  NO2        u117(.A(men_men_n80_), .B(men_men_n99_), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x3), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n133_), .A1(men_men_n132_), .B0(men_men_n135_), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n137_));
  NA2        u121(.A(x5), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n46_), .B(x2), .Y(men_men_n139_));
  NA3        u123(.A(men_men_n139_), .B(men_men_n138_), .C(men_men_n137_), .Y(men_men_n140_));
  NA4        u124(.A(men_men_n140_), .B(men_men_n136_), .C(men_men_n130_), .D(men_men_n34_), .Y(men_men_n141_));
  NO3        u125(.A(men_men_n141_), .B(men_men_n128_), .C(men_men_n113_), .Y(men_men_n142_));
  NO3        u126(.A(men_men_n75_), .B(men_men_n73_), .C(men_men_n24_), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n144_));
  AOI220     u128(.A0(men_men_n122_), .A1(men_men_n144_), .B0(men_men_n63_), .B1(men_men_n17_), .Y(men_men_n145_));
  NO3        u129(.A(men_men_n145_), .B(men_men_n57_), .C(men_men_n59_), .Y(men_men_n146_));
  NA2        u130(.A(x7), .B(x3), .Y(men_men_n147_));
  NO2        u131(.A(men_men_n98_), .B(x5), .Y(men_men_n148_));
  NO2        u132(.A(x9), .B(x7), .Y(men_men_n149_));
  NOi21      u133(.An(x8), .B(x0), .Y(men_men_n150_));
  OA210      u134(.A0(men_men_n149_), .A1(x1), .B0(men_men_n150_), .Y(men_men_n151_));
  NO2        u135(.A(men_men_n41_), .B(x2), .Y(men_men_n152_));
  INV        u136(.A(x7), .Y(men_men_n153_));
  NA2        u137(.A(men_men_n153_), .B(men_men_n18_), .Y(men_men_n154_));
  AOI220     u138(.A0(men_men_n154_), .A1(men_men_n152_), .B0(men_men_n107_), .B1(men_men_n36_), .Y(men_men_n155_));
  NO2        u139(.A(men_men_n25_), .B(x4), .Y(men_men_n156_));
  NO2        u140(.A(x4), .B(men_men_n155_), .Y(men_men_n157_));
  AOI210     u141(.A0(men_men_n151_), .A1(men_men_n148_), .B0(men_men_n157_), .Y(men_men_n158_));
  OAI210     u142(.A0(men_men_n147_), .A1(men_men_n48_), .B0(men_men_n158_), .Y(men_men_n159_));
  NA2        u143(.A(x5), .B(x1), .Y(men_men_n160_));
  INV        u144(.A(men_men_n160_), .Y(men_men_n161_));
  AOI210     u145(.A0(men_men_n161_), .A1(men_men_n124_), .B0(men_men_n34_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n59_), .B(men_men_n90_), .Y(men_men_n163_));
  NAi21      u147(.An(x2), .B(x7), .Y(men_men_n164_));
  NO3        u148(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n46_), .Y(men_men_n165_));
  NA2        u149(.A(men_men_n165_), .B(men_men_n63_), .Y(men_men_n166_));
  NAi31      u150(.An(men_men_n75_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n167_));
  NA3        u151(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n162_), .Y(men_men_n168_));
  NO4        u152(.A(men_men_n168_), .B(men_men_n159_), .C(men_men_n146_), .D(men_men_n143_), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n169_), .B(men_men_n142_), .Y(men_men_n170_));
  NA2        u154(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n172_));
  NA2        u156(.A(x8), .B(x0), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n153_), .B(men_men_n25_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n122_), .B(x4), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  INV        u160(.A(men_men_n176_), .Y(men_men_n177_));
  NA2        u161(.A(x2), .B(x0), .Y(men_men_n178_));
  NA2        u162(.A(x4), .B(x1), .Y(men_men_n179_));
  NAi21      u163(.An(men_men_n120_), .B(men_men_n179_), .Y(men_men_n180_));
  NOi31      u164(.An(men_men_n180_), .B(men_men_n156_), .C(men_men_n178_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n181_), .B(men_men_n177_), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n182_), .B(men_men_n41_), .Y(men_men_n183_));
  INV        u167(.A(men_men_n129_), .Y(men_men_n184_));
  NO2        u168(.A(men_men_n104_), .B(men_men_n17_), .Y(men_men_n185_));
  AOI210     u169(.A0(men_men_n33_), .A1(men_men_n90_), .B0(men_men_n185_), .Y(men_men_n186_));
  NO3        u170(.A(men_men_n186_), .B(men_men_n184_), .C(x7), .Y(men_men_n187_));
  NA3        u171(.A(men_men_n180_), .B(men_men_n184_), .C(men_men_n40_), .Y(men_men_n188_));
  OAI210     u172(.A0(men_men_n172_), .A1(men_men_n134_), .B0(men_men_n188_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n189_), .B(men_men_n187_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(x3), .Y(men_men_n191_));
  NO3        u175(.A(men_men_n191_), .B(men_men_n183_), .C(men_men_n170_), .Y(men03));
  NO2        u176(.A(men_men_n46_), .B(x3), .Y(men_men_n193_));
  NO2        u177(.A(x6), .B(men_men_n25_), .Y(men_men_n194_));
  INV        u178(.A(men_men_n194_), .Y(men_men_n195_));
  NO2        u179(.A(men_men_n52_), .B(x1), .Y(men_men_n196_));
  OAI210     u180(.A0(men_men_n196_), .A1(men_men_n25_), .B0(men_men_n60_), .Y(men_men_n197_));
  OAI220     u181(.A0(men_men_n197_), .A1(men_men_n17_), .B0(men_men_n195_), .B1(men_men_n104_), .Y(men_men_n198_));
  NA2        u182(.A(men_men_n198_), .B(men_men_n193_), .Y(men_men_n199_));
  NO2        u183(.A(men_men_n75_), .B(x6), .Y(men_men_n200_));
  NA2        u184(.A(x6), .B(men_men_n25_), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n201_), .B(x4), .Y(men_men_n202_));
  NO2        u186(.A(men_men_n18_), .B(x0), .Y(men_men_n203_));
  AO220      u187(.A0(men_men_n203_), .A1(men_men_n202_), .B0(men_men_n200_), .B1(men_men_n53_), .Y(men_men_n204_));
  NA2        u188(.A(men_men_n204_), .B(men_men_n59_), .Y(men_men_n205_));
  NA2        u189(.A(x3), .B(men_men_n17_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n206_), .B(men_men_n201_), .Y(men_men_n207_));
  NA2        u191(.A(x9), .B(men_men_n52_), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n208_), .B(x4), .Y(men_men_n209_));
  NA2        u193(.A(men_men_n201_), .B(men_men_n78_), .Y(men_men_n210_));
  AOI210     u194(.A0(men_men_n25_), .A1(x3), .B0(men_men_n178_), .Y(men_men_n211_));
  AOI220     u195(.A0(men_men_n211_), .A1(men_men_n210_), .B0(men_men_n209_), .B1(men_men_n207_), .Y(men_men_n212_));
  NO3        u196(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n213_));
  NO2        u197(.A(x5), .B(x1), .Y(men_men_n214_));
  AOI220     u198(.A0(men_men_n214_), .A1(men_men_n17_), .B0(men_men_n101_), .B1(x5), .Y(men_men_n215_));
  NO2        u199(.A(men_men_n206_), .B(men_men_n171_), .Y(men_men_n216_));
  NO3        u200(.A(x3), .B(x2), .C(x1), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  OAI210     u202(.A0(men_men_n215_), .A1(men_men_n61_), .B0(men_men_n218_), .Y(men_men_n219_));
  AOI220     u203(.A0(men_men_n219_), .A1(men_men_n46_), .B0(men_men_n213_), .B1(men_men_n129_), .Y(men_men_n220_));
  NA4        u204(.A(men_men_n220_), .B(men_men_n212_), .C(men_men_n205_), .D(men_men_n199_), .Y(men_men_n221_));
  NO2        u205(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n222_), .B(men_men_n19_), .Y(men_men_n223_));
  NO2        u207(.A(x3), .B(men_men_n17_), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n224_), .B(x6), .Y(men_men_n225_));
  NOi21      u209(.An(men_men_n80_), .B(men_men_n225_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n59_), .B(men_men_n90_), .Y(men_men_n227_));
  NA3        u211(.A(men_men_n227_), .B(men_men_n224_), .C(x6), .Y(men_men_n228_));
  AOI210     u212(.A0(men_men_n228_), .A1(men_men_n226_), .B0(men_men_n153_), .Y(men_men_n229_));
  AO210      u213(.A0(men_men_n229_), .A1(men_men_n223_), .B0(men_men_n174_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n25_), .B0(men_men_n172_), .Y(men_men_n232_));
  NO3        u216(.A(men_men_n179_), .B(men_men_n59_), .C(x6), .Y(men_men_n233_));
  NA2        u217(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  NA2        u218(.A(x6), .B(men_men_n46_), .Y(men_men_n235_));
  OAI210     u219(.A0(men_men_n116_), .A1(men_men_n76_), .B0(x4), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n75_), .Y(men_men_n237_));
  NO2        u221(.A(men_men_n59_), .B(x6), .Y(men_men_n238_));
  NO2        u222(.A(men_men_n160_), .B(men_men_n41_), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n239_), .A1(men_men_n216_), .B0(men_men_n238_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n194_), .B(men_men_n132_), .Y(men_men_n241_));
  NA3        u225(.A(men_men_n206_), .B(men_men_n129_), .C(x6), .Y(men_men_n242_));
  OAI210     u226(.A0(men_men_n90_), .A1(men_men_n34_), .B0(men_men_n63_), .Y(men_men_n243_));
  NA4        u227(.A(men_men_n243_), .B(men_men_n242_), .C(men_men_n241_), .D(men_men_n240_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n237_), .B0(x2), .Y(men_men_n245_));
  NA3        u229(.A(men_men_n245_), .B(men_men_n234_), .C(men_men_n230_), .Y(men_men_n246_));
  AOI210     u230(.A0(men_men_n221_), .A1(x8), .B0(men_men_n246_), .Y(men_men_n247_));
  NO2        u231(.A(men_men_n90_), .B(x3), .Y(men_men_n248_));
  NA2        u232(.A(men_men_n248_), .B(men_men_n202_), .Y(men_men_n249_));
  NO3        u233(.A(men_men_n88_), .B(men_men_n76_), .C(men_men_n25_), .Y(men_men_n250_));
  AOI210     u234(.A0(men_men_n225_), .A1(men_men_n156_), .B0(men_men_n250_), .Y(men_men_n251_));
  AOI210     u235(.A0(men_men_n251_), .A1(men_men_n249_), .B0(x2), .Y(men_men_n252_));
  NO2        u236(.A(x4), .B(men_men_n52_), .Y(men_men_n253_));
  AOI220     u237(.A0(men_men_n202_), .A1(men_men_n185_), .B0(men_men_n253_), .B1(men_men_n63_), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n59_), .B(x6), .Y(men_men_n255_));
  NA3        u239(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n256_));
  AOI210     u240(.A0(men_men_n256_), .A1(men_men_n138_), .B0(men_men_n255_), .Y(men_men_n257_));
  NA2        u241(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n258_), .B(men_men_n25_), .Y(men_men_n259_));
  OAI210     u243(.A0(men_men_n259_), .A1(men_men_n257_), .B0(men_men_n120_), .Y(men_men_n260_));
  NO2        u244(.A(men_men_n206_), .B(x6), .Y(men_men_n261_));
  NAi21      u245(.An(men_men_n163_), .B(men_men_n261_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n262_), .B(men_men_n144_), .Y(men_men_n263_));
  NA4        u247(.A(men_men_n263_), .B(men_men_n260_), .C(men_men_n254_), .D(men_men_n153_), .Y(men_men_n264_));
  NA2        u248(.A(men_men_n194_), .B(men_men_n224_), .Y(men_men_n265_));
  NO2        u249(.A(x9), .B(x6), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n138_), .B(men_men_n18_), .Y(men_men_n267_));
  NAi21      u251(.An(men_men_n267_), .B(men_men_n256_), .Y(men_men_n268_));
  NAi21      u252(.An(x1), .B(x4), .Y(men_men_n269_));
  AOI210     u253(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n270_));
  OAI210     u254(.A0(men_men_n138_), .A1(x3), .B0(men_men_n270_), .Y(men_men_n271_));
  AOI220     u255(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n268_), .B1(men_men_n266_), .Y(men_men_n272_));
  NA2        u256(.A(men_men_n272_), .B(men_men_n265_), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n59_), .B(x2), .Y(men_men_n274_));
  NO2        u258(.A(men_men_n274_), .B(men_men_n265_), .Y(men_men_n275_));
  NO3        u259(.A(x9), .B(x6), .C(x0), .Y(men_men_n276_));
  NA2        u260(.A(men_men_n104_), .B(men_men_n25_), .Y(men_men_n277_));
  NA2        u261(.A(x6), .B(x2), .Y(men_men_n278_));
  NO2        u262(.A(men_men_n278_), .B(men_men_n171_), .Y(men_men_n279_));
  AOI210     u263(.A0(men_men_n277_), .A1(men_men_n276_), .B0(men_men_n279_), .Y(men_men_n280_));
  OAI220     u264(.A0(men_men_n280_), .A1(men_men_n41_), .B0(men_men_n175_), .B1(men_men_n44_), .Y(men_men_n281_));
  OAI210     u265(.A0(men_men_n281_), .A1(men_men_n275_), .B0(men_men_n273_), .Y(men_men_n282_));
  NA2        u266(.A(x9), .B(men_men_n41_), .Y(men_men_n283_));
  NO2        u267(.A(men_men_n283_), .B(men_men_n201_), .Y(men_men_n284_));
  OR3        u268(.A(men_men_n284_), .B(men_men_n200_), .C(men_men_n148_), .Y(men_men_n285_));
  NA2        u269(.A(x4), .B(x0), .Y(men_men_n286_));
  NO3        u270(.A(men_men_n70_), .B(men_men_n286_), .C(x6), .Y(men_men_n287_));
  AOI210     u271(.A0(men_men_n285_), .A1(men_men_n40_), .B0(men_men_n287_), .Y(men_men_n288_));
  AOI210     u272(.A0(men_men_n288_), .A1(men_men_n282_), .B0(x8), .Y(men_men_n289_));
  INV        u273(.A(men_men_n255_), .Y(men_men_n290_));
  OAI210     u274(.A0(men_men_n267_), .A1(men_men_n214_), .B0(men_men_n290_), .Y(men_men_n291_));
  INV        u275(.A(men_men_n173_), .Y(men_men_n292_));
  OAI210     u276(.A0(men_men_n292_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n293_));
  AOI210     u277(.A0(men_men_n293_), .A1(men_men_n291_), .B0(men_men_n231_), .Y(men_men_n294_));
  NO4        u278(.A(men_men_n294_), .B(men_men_n289_), .C(men_men_n264_), .D(men_men_n252_), .Y(men_men_n295_));
  NO2        u279(.A(men_men_n163_), .B(x1), .Y(men_men_n296_));
  NO3        u280(.A(men_men_n296_), .B(x3), .C(men_men_n34_), .Y(men_men_n297_));
  OAI210     u281(.A0(men_men_n297_), .A1(men_men_n261_), .B0(x2), .Y(men_men_n298_));
  OAI210     u282(.A0(men_men_n292_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n299_));
  AOI210     u283(.A0(men_men_n299_), .A1(men_men_n298_), .B0(men_men_n184_), .Y(men_men_n300_));
  NOi21      u284(.An(men_men_n278_), .B(men_men_n17_), .Y(men_men_n301_));
  NA3        u285(.A(men_men_n301_), .B(men_men_n214_), .C(men_men_n38_), .Y(men_men_n302_));
  AOI210     u286(.A0(men_men_n34_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n303_));
  NA3        u287(.A(men_men_n303_), .B(men_men_n161_), .C(men_men_n31_), .Y(men_men_n304_));
  NA2        u288(.A(x3), .B(x2), .Y(men_men_n305_));
  AOI220     u289(.A0(men_men_n305_), .A1(men_men_n231_), .B0(men_men_n304_), .B1(men_men_n302_), .Y(men_men_n306_));
  NAi21      u290(.An(x4), .B(x0), .Y(men_men_n307_));
  NO3        u291(.A(men_men_n307_), .B(men_men_n42_), .C(x2), .Y(men_men_n308_));
  OAI210     u292(.A0(x6), .A1(men_men_n18_), .B0(men_men_n308_), .Y(men_men_n309_));
  OAI220     u293(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n310_));
  NO2        u294(.A(x9), .B(x8), .Y(men_men_n311_));
  NA3        u295(.A(men_men_n311_), .B(men_men_n34_), .C(men_men_n52_), .Y(men_men_n312_));
  OAI210     u296(.A0(men_men_n303_), .A1(men_men_n301_), .B0(men_men_n312_), .Y(men_men_n313_));
  AOI220     u297(.A0(men_men_n313_), .A1(men_men_n79_), .B0(men_men_n310_), .B1(men_men_n30_), .Y(men_men_n314_));
  AOI210     u298(.A0(men_men_n314_), .A1(men_men_n309_), .B0(men_men_n25_), .Y(men_men_n315_));
  NA3        u299(.A(men_men_n34_), .B(x1), .C(men_men_n17_), .Y(men_men_n316_));
  OAI210     u300(.A0(men_men_n303_), .A1(men_men_n301_), .B0(men_men_n316_), .Y(men_men_n317_));
  INV        u301(.A(men_men_n216_), .Y(men_men_n318_));
  NA2        u302(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n319_));
  OR2        u303(.A(men_men_n319_), .B(men_men_n286_), .Y(men_men_n320_));
  OAI220     u304(.A0(men_men_n320_), .A1(men_men_n160_), .B0(men_men_n235_), .B1(men_men_n318_), .Y(men_men_n321_));
  AO210      u305(.A0(men_men_n317_), .A1(men_men_n148_), .B0(men_men_n321_), .Y(men_men_n322_));
  NO4        u306(.A(men_men_n322_), .B(men_men_n315_), .C(men_men_n306_), .D(men_men_n300_), .Y(men_men_n323_));
  OAI210     u307(.A0(men_men_n295_), .A1(men_men_n247_), .B0(men_men_n323_), .Y(men04));
  OAI210     u308(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n325_));
  NA3        u309(.A(men_men_n325_), .B(men_men_n276_), .C(men_men_n81_), .Y(men_men_n326_));
  NO2        u310(.A(x2), .B(x1), .Y(men_men_n327_));
  OAI210     u311(.A0(men_men_n258_), .A1(men_men_n327_), .B0(men_men_n34_), .Y(men_men_n328_));
  NO2        u312(.A(men_men_n327_), .B(men_men_n307_), .Y(men_men_n329_));
  AOI210     u313(.A0(men_men_n59_), .A1(x4), .B0(men_men_n109_), .Y(men_men_n330_));
  OAI210     u314(.A0(men_men_n330_), .A1(men_men_n329_), .B0(men_men_n248_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n274_), .B(men_men_n88_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n332_), .B(men_men_n34_), .Y(men_men_n333_));
  NA2        u317(.A(x9), .B(x0), .Y(men_men_n334_));
  AOI210     u318(.A0(men_men_n88_), .A1(men_men_n73_), .B0(men_men_n334_), .Y(men_men_n335_));
  OAI210     u319(.A0(men_men_n335_), .A1(men_men_n475_), .B0(men_men_n90_), .Y(men_men_n336_));
  NA3        u320(.A(men_men_n336_), .B(men_men_n333_), .C(men_men_n331_), .Y(men_men_n337_));
  NA2        u321(.A(men_men_n337_), .B(men_men_n328_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n208_), .B(men_men_n110_), .Y(men_men_n339_));
  NO3        u323(.A(men_men_n255_), .B(men_men_n117_), .C(men_men_n18_), .Y(men_men_n340_));
  NO2        u324(.A(men_men_n340_), .B(men_men_n339_), .Y(men_men_n341_));
  OAI210     u325(.A0(men_men_n115_), .A1(men_men_n104_), .B0(men_men_n173_), .Y(men_men_n342_));
  NA3        u326(.A(men_men_n342_), .B(x6), .C(x3), .Y(men_men_n343_));
  AOI210     u327(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n344_));
  OAI220     u328(.A0(men_men_n344_), .A1(men_men_n319_), .B0(men_men_n274_), .B1(men_men_n316_), .Y(men_men_n345_));
  AOI210     u329(.A0(x2), .A1(men_men_n60_), .B0(men_men_n345_), .Y(men_men_n346_));
  NA2        u330(.A(x2), .B(men_men_n17_), .Y(men_men_n347_));
  OAI210     u331(.A0(men_men_n104_), .A1(men_men_n17_), .B0(men_men_n347_), .Y(men_men_n348_));
  AOI220     u332(.A0(men_men_n348_), .A1(men_men_n76_), .B0(men_men_n332_), .B1(men_men_n90_), .Y(men_men_n349_));
  NA4        u333(.A(men_men_n349_), .B(men_men_n346_), .C(men_men_n343_), .D(men_men_n341_), .Y(men_men_n350_));
  OAI210     u334(.A0(men_men_n108_), .A1(x3), .B0(men_men_n308_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n227_), .B(men_men_n213_), .C(men_men_n80_), .Y(men_men_n352_));
  NA3        u336(.A(men_men_n352_), .B(men_men_n351_), .C(men_men_n153_), .Y(men_men_n353_));
  AOI210     u337(.A0(men_men_n350_), .A1(x4), .B0(men_men_n353_), .Y(men_men_n354_));
  NA3        u338(.A(men_men_n329_), .B(men_men_n208_), .C(men_men_n90_), .Y(men_men_n355_));
  NOi21      u339(.An(x4), .B(x0), .Y(men_men_n356_));
  XO2        u340(.A(x4), .B(x0), .Y(men_men_n357_));
  OAI210     u341(.A0(men_men_n357_), .A1(men_men_n114_), .B0(men_men_n269_), .Y(men_men_n358_));
  AOI210     u342(.A0(men_men_n358_), .A1(x8), .B0(men_men_n356_), .Y(men_men_n359_));
  AOI210     u343(.A0(men_men_n359_), .A1(men_men_n355_), .B0(x3), .Y(men_men_n360_));
  INV        u344(.A(men_men_n91_), .Y(men_men_n361_));
  NO2        u345(.A(men_men_n90_), .B(x4), .Y(men_men_n362_));
  NO3        u346(.A(men_men_n357_), .B(men_men_n163_), .C(x2), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n28_), .B(men_men_n24_), .Y(men_men_n364_));
  NO2        u348(.A(men_men_n364_), .B(men_men_n363_), .Y(men_men_n365_));
  NA4        u349(.A(men_men_n365_), .B(men_men_n91_), .C(men_men_n223_), .D(x6), .Y(men_men_n366_));
  OAI220     u350(.A0(men_men_n307_), .A1(men_men_n88_), .B0(men_men_n178_), .B1(men_men_n90_), .Y(men_men_n367_));
  NO2        u351(.A(men_men_n41_), .B(x0), .Y(men_men_n368_));
  OR2        u352(.A(men_men_n362_), .B(men_men_n368_), .Y(men_men_n369_));
  NO2        u353(.A(men_men_n150_), .B(men_men_n104_), .Y(men_men_n370_));
  AOI220     u354(.A0(men_men_n370_), .A1(men_men_n369_), .B0(men_men_n367_), .B1(men_men_n58_), .Y(men_men_n371_));
  NO2        u355(.A(men_men_n150_), .B(men_men_n78_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n33_), .B(x2), .Y(men_men_n373_));
  NOi21      u357(.An(men_men_n120_), .B(men_men_n27_), .Y(men_men_n374_));
  AOI210     u358(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n374_), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n371_), .A1(men_men_n59_), .B0(men_men_n375_), .Y(men_men_n376_));
  OAI220     u360(.A0(men_men_n376_), .A1(x6), .B0(men_men_n366_), .B1(men_men_n360_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n60_), .A1(men_men_n46_), .B0(men_men_n40_), .Y(men_men_n378_));
  OAI210     u362(.A0(men_men_n378_), .A1(men_men_n90_), .B0(men_men_n320_), .Y(men_men_n379_));
  AOI210     u363(.A0(men_men_n379_), .A1(men_men_n18_), .B0(men_men_n153_), .Y(men_men_n380_));
  AO220      u364(.A0(men_men_n380_), .A1(men_men_n377_), .B0(men_men_n354_), .B1(men_men_n338_), .Y(men_men_n381_));
  AOI210     u365(.A0(x6), .A1(x1), .B0(men_men_n152_), .Y(men_men_n382_));
  NA2        u366(.A(men_men_n362_), .B(x0), .Y(men_men_n383_));
  NO2        u367(.A(men_men_n383_), .B(men_men_n382_), .Y(men_men_n384_));
  AOI220     u368(.A0(men_men_n384_), .A1(men_men_n474_), .B0(men_men_n217_), .B1(men_men_n47_), .Y(men_men_n385_));
  NA3        u369(.A(men_men_n385_), .B(men_men_n381_), .C(men_men_n326_), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n196_), .A1(x8), .B0(men_men_n108_), .Y(men_men_n387_));
  NA2        u371(.A(men_men_n387_), .B(men_men_n347_), .Y(men_men_n388_));
  NA3        u372(.A(men_men_n388_), .B(men_men_n193_), .C(men_men_n153_), .Y(men_men_n389_));
  OAI210     u373(.A0(men_men_n28_), .A1(x1), .B0(men_men_n231_), .Y(men_men_n390_));
  AO220      u374(.A0(men_men_n390_), .A1(men_men_n149_), .B0(men_men_n107_), .B1(x4), .Y(men_men_n391_));
  NA3        u375(.A(x7), .B(x3), .C(x0), .Y(men_men_n392_));
  NA2        u376(.A(men_men_n222_), .B(x0), .Y(men_men_n393_));
  OAI220     u377(.A0(men_men_n393_), .A1(men_men_n208_), .B0(men_men_n392_), .B1(men_men_n361_), .Y(men_men_n394_));
  AOI210     u378(.A0(men_men_n391_), .A1(men_men_n116_), .B0(men_men_n394_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n395_), .A1(men_men_n389_), .B0(men_men_n25_), .Y(men_men_n396_));
  NA3        u380(.A(men_men_n118_), .B(men_men_n222_), .C(x0), .Y(men_men_n397_));
  OAI210     u381(.A0(men_men_n193_), .A1(men_men_n64_), .B0(men_men_n203_), .Y(men_men_n398_));
  NA3        u382(.A(men_men_n196_), .B(men_men_n224_), .C(x8), .Y(men_men_n399_));
  AOI210     u383(.A0(men_men_n399_), .A1(men_men_n398_), .B0(men_men_n25_), .Y(men_men_n400_));
  AOI210     u384(.A0(men_men_n117_), .A1(men_men_n115_), .B0(men_men_n40_), .Y(men_men_n401_));
  NOi31      u385(.An(men_men_n401_), .B(men_men_n368_), .C(men_men_n179_), .Y(men_men_n402_));
  OAI210     u386(.A0(men_men_n402_), .A1(men_men_n400_), .B0(men_men_n149_), .Y(men_men_n403_));
  NAi31      u387(.An(men_men_n48_), .B(men_men_n296_), .C(men_men_n174_), .Y(men_men_n404_));
  NA3        u388(.A(men_men_n404_), .B(men_men_n403_), .C(men_men_n397_), .Y(men_men_n405_));
  OAI210     u389(.A0(men_men_n405_), .A1(men_men_n396_), .B0(x6), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n163_), .A1(men_men_n46_), .B0(men_men_n133_), .Y(men_men_n407_));
  NA3        u391(.A(men_men_n53_), .B(men_men_n36_), .C(men_men_n30_), .Y(men_men_n408_));
  AOI220     u392(.A0(men_men_n408_), .A1(men_men_n407_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n409_));
  NO2        u393(.A(men_men_n153_), .B(x0), .Y(men_men_n410_));
  NA2        u394(.A(men_men_n193_), .B(men_men_n153_), .Y(men_men_n411_));
  AOI210     u395(.A0(men_men_n126_), .A1(men_men_n253_), .B0(x1), .Y(men_men_n412_));
  OAI210     u396(.A0(men_men_n411_), .A1(x8), .B0(men_men_n412_), .Y(men_men_n413_));
  NAi31      u397(.An(x2), .B(x8), .C(x0), .Y(men_men_n414_));
  OAI210     u398(.A0(men_men_n414_), .A1(x4), .B0(men_men_n164_), .Y(men_men_n415_));
  NA3        u399(.A(men_men_n415_), .B(men_men_n147_), .C(x9), .Y(men_men_n416_));
  NO4        u400(.A(men_men_n125_), .B(men_men_n307_), .C(x9), .D(x2), .Y(men_men_n417_));
  NOi21      u401(.An(men_men_n123_), .B(men_men_n178_), .Y(men_men_n418_));
  NO3        u402(.A(men_men_n418_), .B(men_men_n417_), .C(men_men_n18_), .Y(men_men_n419_));
  NO3        u403(.A(x9), .B(men_men_n153_), .C(x0), .Y(men_men_n420_));
  AOI220     u404(.A0(men_men_n420_), .A1(men_men_n248_), .B0(men_men_n372_), .B1(men_men_n153_), .Y(men_men_n421_));
  NA4        u405(.A(men_men_n421_), .B(men_men_n419_), .C(men_men_n416_), .D(men_men_n48_), .Y(men_men_n422_));
  OAI210     u406(.A0(men_men_n413_), .A1(men_men_n409_), .B0(men_men_n422_), .Y(men_men_n423_));
  NOi31      u407(.An(men_men_n410_), .B(men_men_n31_), .C(x8), .Y(men_men_n424_));
  AOI210     u408(.A0(men_men_n36_), .A1(x9), .B0(men_men_n131_), .Y(men_men_n425_));
  NO3        u409(.A(men_men_n425_), .B(men_men_n123_), .C(men_men_n41_), .Y(men_men_n426_));
  NOi31      u410(.An(x1), .B(x8), .C(x7), .Y(men_men_n427_));
  AOI220     u411(.A0(men_men_n427_), .A1(men_men_n356_), .B0(men_men_n124_), .B1(x3), .Y(men_men_n428_));
  AOI210     u412(.A0(men_men_n269_), .A1(men_men_n57_), .B0(men_men_n122_), .Y(men_men_n429_));
  OAI210     u413(.A0(men_men_n429_), .A1(x3), .B0(men_men_n428_), .Y(men_men_n430_));
  NO3        u414(.A(men_men_n430_), .B(men_men_n426_), .C(x2), .Y(men_men_n431_));
  OAI220     u415(.A0(men_men_n357_), .A1(men_men_n311_), .B0(men_men_n307_), .B1(men_men_n41_), .Y(men_men_n432_));
  AOI210     u416(.A0(x9), .A1(men_men_n46_), .B0(men_men_n392_), .Y(men_men_n433_));
  AOI220     u417(.A0(men_men_n433_), .A1(men_men_n90_), .B0(men_men_n432_), .B1(men_men_n153_), .Y(men_men_n434_));
  NO2        u418(.A(men_men_n434_), .B(men_men_n52_), .Y(men_men_n435_));
  NO3        u419(.A(men_men_n435_), .B(men_men_n431_), .C(men_men_n424_), .Y(men_men_n436_));
  AOI210     u420(.A0(men_men_n436_), .A1(men_men_n423_), .B0(men_men_n25_), .Y(men_men_n437_));
  NA4        u421(.A(men_men_n30_), .B(men_men_n90_), .C(x2), .D(men_men_n17_), .Y(men_men_n438_));
  NO3        u422(.A(men_men_n59_), .B(x4), .C(x1), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n64_), .B(men_men_n18_), .C(x0), .Y(men_men_n440_));
  AOI220     u424(.A0(men_men_n440_), .A1(men_men_n270_), .B0(men_men_n439_), .B1(men_men_n401_), .Y(men_men_n441_));
  NO2        u425(.A(men_men_n441_), .B(men_men_n101_), .Y(men_men_n442_));
  NO3        u426(.A(men_men_n274_), .B(men_men_n173_), .C(men_men_n38_), .Y(men_men_n443_));
  OAI210     u427(.A0(men_men_n443_), .A1(men_men_n442_), .B0(x7), .Y(men_men_n444_));
  NA2        u428(.A(men_men_n227_), .B(x7), .Y(men_men_n445_));
  NA3        u429(.A(men_men_n445_), .B(men_men_n152_), .C(men_men_n132_), .Y(men_men_n446_));
  NA3        u430(.A(men_men_n446_), .B(men_men_n444_), .C(men_men_n438_), .Y(men_men_n447_));
  OAI210     u431(.A0(men_men_n447_), .A1(men_men_n437_), .B0(men_men_n34_), .Y(men_men_n448_));
  NO2        u432(.A(men_men_n420_), .B(men_men_n203_), .Y(men_men_n449_));
  NO4        u433(.A(men_men_n449_), .B(men_men_n75_), .C(x4), .D(men_men_n52_), .Y(men_men_n450_));
  NA2        u434(.A(men_men_n258_), .B(men_men_n21_), .Y(men_men_n451_));
  NO2        u435(.A(men_men_n160_), .B(men_men_n133_), .Y(men_men_n452_));
  NA2        u436(.A(men_men_n452_), .B(men_men_n451_), .Y(men_men_n453_));
  AOI210     u437(.A0(men_men_n453_), .A1(men_men_n167_), .B0(men_men_n28_), .Y(men_men_n454_));
  AOI220     u438(.A0(men_men_n368_), .A1(men_men_n90_), .B0(men_men_n150_), .B1(men_men_n196_), .Y(men_men_n455_));
  NA3        u439(.A(men_men_n455_), .B(men_men_n414_), .C(men_men_n88_), .Y(men_men_n456_));
  NA2        u440(.A(men_men_n456_), .B(men_men_n174_), .Y(men_men_n457_));
  OAI220     u441(.A0(men_men_n283_), .A1(men_men_n65_), .B0(men_men_n160_), .B1(men_men_n41_), .Y(men_men_n458_));
  NA2        u442(.A(x3), .B(men_men_n52_), .Y(men_men_n459_));
  AOI210     u443(.A0(men_men_n164_), .A1(men_men_n27_), .B0(men_men_n70_), .Y(men_men_n460_));
  OAI210     u444(.A0(men_men_n149_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n461_));
  NO3        u445(.A(men_men_n427_), .B(x3), .C(men_men_n52_), .Y(men_men_n462_));
  AOI210     u446(.A0(men_men_n462_), .A1(men_men_n461_), .B0(men_men_n460_), .Y(men_men_n463_));
  OAI210     u447(.A0(men_men_n154_), .A1(men_men_n459_), .B0(men_men_n463_), .Y(men_men_n464_));
  AOI220     u448(.A0(men_men_n464_), .A1(x0), .B0(men_men_n458_), .B1(men_men_n133_), .Y(men_men_n465_));
  AOI210     u449(.A0(men_men_n465_), .A1(men_men_n457_), .B0(men_men_n235_), .Y(men_men_n466_));
  NA2        u450(.A(x9), .B(x5), .Y(men_men_n467_));
  NO4        u451(.A(men_men_n104_), .B(men_men_n467_), .C(men_men_n57_), .D(men_men_n31_), .Y(men_men_n468_));
  NO4        u452(.A(men_men_n468_), .B(men_men_n466_), .C(men_men_n454_), .D(men_men_n450_), .Y(men_men_n469_));
  NA3        u453(.A(men_men_n469_), .B(men_men_n448_), .C(men_men_n406_), .Y(men_men_n470_));
  AOI210     u454(.A0(men_men_n386_), .A1(men_men_n25_), .B0(men_men_n470_), .Y(men05));
  INV        u455(.A(x6), .Y(men_men_n474_));
  INV        u456(.A(men_men_n305_), .Y(men_men_n475_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule