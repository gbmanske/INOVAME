// Benchmark "top" written by ABC on Thu Jun 20 14:00:08 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n143_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1077_, new_new_n1078_, new_new_n1079_,
    new_new_n1080_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  OAI210     g0067(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n89_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_10_), .Y(new_new_n91_));
  NA2        g0069(.A(i_6_), .B(i_9_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n91_), .B0(new_new_n64_), .Y(new_new_n93_));
  NA2        g0071(.A(i_2_), .B(i_6_), .Y(new_new_n94_));
  NO3        g0072(.A(new_new_n94_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n95_));
  NO2        g0073(.A(new_new_n95_), .B(new_new_n93_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n90_), .B0(new_new_n81_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n63_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n87_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  NO3        g0088(.A(new_new_n110_), .B(new_new_n91_), .C(new_new_n54_), .Y(new_new_n111_));
  AN2        g0089(.A(i_2_), .B(i_10_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n112_), .B(i_7_), .Y(new_new_n113_));
  OR2        g0091(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n114_));
  NO2        g0092(.A(i_8_), .B(new_new_n103_), .Y(new_new_n115_));
  NO3        g0093(.A(new_new_n115_), .B(new_new_n114_), .C(new_new_n113_), .Y(new_new_n116_));
  NA2        g0094(.A(i_12_), .B(i_7_), .Y(new_new_n117_));
  NO2        g0095(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n118_));
  NA2        g0096(.A(new_new_n118_), .B(i_0_), .Y(new_new_n119_));
  NA2        g0097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  OAI210     g0098(.A0(new_new_n119_), .A1(new_new_n117_), .B0(new_new_n120_), .Y(new_new_n121_));
  NO2        g0099(.A(new_new_n121_), .B(new_new_n116_), .Y(new_new_n122_));
  NAi41      g0100(.An(new_new_n111_), .B(new_new_n122_), .C(new_new_n109_), .D(new_new_n102_), .Y(new_new_n123_));
  NOi21      g0101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g0104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g0106(.A(new_new_n128_), .B(new_new_n47_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n92_), .B(new_new_n91_), .Y(new_new_n130_));
  NAi21      g0108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n131_), .B(new_new_n63_), .Y(new_new_n132_));
  NOi31      g0110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g0111(.A(i_1_), .B(new_new_n87_), .Y(new_new_n134_));
  NO2        g0112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g0113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g0114(.A0(new_new_n136_), .A1(new_new_n48_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g0115(.A0(new_new_n137_), .A1(new_new_n110_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g0116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n97_), .Y(new_new_n139_));
  NA3        g0117(.A(new_new_n139_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g0118(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g0119(.A(i_6_), .B(new_new_n25_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(new_new_n141_), .Y(new_new_n143_));
  NA4        g0121(.A(new_new_n143_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g0122(.A(i_8_), .B(i_7_), .Y(new_new_n145_));
  NA2        g0123(.A(new_new_n145_), .B(i_6_), .Y(new_new_n146_));
  NO2        g0124(.A(i_12_), .B(i_13_), .Y(new_new_n147_));
  NAi21      g0125(.An(i_5_), .B(i_11_), .Y(new_new_n148_));
  NOi21      g0126(.An(new_new_n147_), .B(new_new_n148_), .Y(new_new_n149_));
  NO2        g0127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NA2        g0128(.A(i_2_), .B(i_3_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(i_4_), .Y(new_new_n152_));
  NA3        g0130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  AN2        g0131(.A(new_new_n147_), .B(new_new_n84_), .Y(new_new_n154_));
  NO2        g0132(.A(new_new_n154_), .B(new_new_n27_), .Y(new_new_n155_));
  NA2        g0133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  NO2        g0134(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n157_));
  NA2        g0135(.A(new_new_n157_), .B(new_new_n36_), .Y(new_new_n158_));
  NO3        g0136(.A(new_new_n158_), .B(new_new_n156_), .C(new_new_n155_), .Y(new_new_n159_));
  OR2        g0137(.A(i_0_), .B(i_1_), .Y(new_new_n160_));
  NO3        g0138(.A(new_new_n160_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n161_));
  NAi32      g0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n162_));
  NAi21      g0140(.An(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NOi21      g0141(.An(i_4_), .B(i_10_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n40_), .Y(new_new_n165_));
  NO2        g0143(.A(i_3_), .B(i_5_), .Y(new_new_n166_));
  NO3        g0144(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n167_));
  NA2        g0145(.A(new_new_n167_), .B(new_new_n166_), .Y(new_new_n168_));
  OAI210     g0146(.A0(new_new_n168_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n169_));
  NO2        g0147(.A(new_new_n169_), .B(new_new_n159_), .Y(new_new_n170_));
  AOI210     g0148(.A0(new_new_n170_), .A1(new_new_n153_), .B0(new_new_n146_), .Y(new_new_n171_));
  NA3        g0149(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n172_));
  NA2        g0150(.A(i_3_), .B(new_new_n49_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_4_), .B(i_9_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_11_), .B(i_13_), .Y(new_new_n175_));
  NA2        g0153(.A(new_new_n175_), .B(new_new_n174_), .Y(new_new_n176_));
  OR2        g0154(.A(new_new_n176_), .B(new_new_n173_), .Y(new_new_n177_));
  NO2        g0155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g0156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n84_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n172_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n183_), .B(new_new_n47_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n36_), .B(i_5_), .Y(new_new_n185_));
  NAi31      g0163(.An(new_new_n185_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n186_));
  NA2        g0164(.A(i_3_), .B(i_5_), .Y(new_new_n187_));
  OR2        g0165(.A(new_new_n187_), .B(new_new_n176_), .Y(new_new_n188_));
  AOI210     g0166(.A0(new_new_n188_), .A1(new_new_n186_), .B0(new_new_n184_), .Y(new_new_n189_));
  NO2        g0167(.A(new_new_n74_), .B(i_5_), .Y(new_new_n190_));
  NO2        g0168(.A(i_13_), .B(i_10_), .Y(new_new_n191_));
  NA3        g0169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n45_), .Y(new_new_n192_));
  NO2        g0170(.A(i_2_), .B(i_1_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_3_), .Y(new_new_n194_));
  NAi21      g0172(.An(i_4_), .B(i_12_), .Y(new_new_n195_));
  NO4        g0173(.A(new_new_n195_), .B(new_new_n194_), .C(new_new_n192_), .D(new_new_n25_), .Y(new_new_n196_));
  NO3        g0174(.A(new_new_n196_), .B(new_new_n189_), .C(new_new_n182_), .Y(new_new_n197_));
  INV        g0175(.A(i_8_), .Y(new_new_n198_));
  NO2        g0176(.A(new_new_n198_), .B(i_7_), .Y(new_new_n199_));
  NA2        g0177(.A(new_new_n199_), .B(i_6_), .Y(new_new_n200_));
  NO3        g0178(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n201_));
  NA2        g0179(.A(new_new_n201_), .B(new_new_n115_), .Y(new_new_n202_));
  NO3        g0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n204_));
  NO3        g0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n205_));
  OAI210     g0183(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n205_), .Y(new_new_n206_));
  AOI210     g0184(.A0(new_new_n206_), .A1(new_new_n204_), .B0(new_new_n202_), .Y(new_new_n207_));
  NO2        g0185(.A(i_3_), .B(i_8_), .Y(new_new_n208_));
  NO3        g0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n105_), .B(new_new_n59_), .Y(new_new_n210_));
  NO2        g0188(.A(i_13_), .B(i_9_), .Y(new_new_n211_));
  NA3        g0189(.A(new_new_n211_), .B(i_6_), .C(new_new_n198_), .Y(new_new_n212_));
  NAi21      g0190(.An(i_12_), .B(i_3_), .Y(new_new_n213_));
  NO2        g0191(.A(new_new_n45_), .B(i_5_), .Y(new_new_n214_));
  NO3        g0192(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n215_));
  NA3        g0193(.A(new_new_n215_), .B(new_new_n214_), .C(i_10_), .Y(new_new_n216_));
  NO2        g0194(.A(new_new_n216_), .B(new_new_n212_), .Y(new_new_n217_));
  AOI210     g0195(.A0(new_new_n217_), .A1(i_7_), .B0(new_new_n207_), .Y(new_new_n218_));
  OAI220     g0196(.A0(new_new_n218_), .A1(i_4_), .B0(new_new_n200_), .B1(new_new_n197_), .Y(new_new_n219_));
  NAi21      g0197(.An(i_12_), .B(i_7_), .Y(new_new_n220_));
  NA3        g0198(.A(i_13_), .B(new_new_n198_), .C(i_10_), .Y(new_new_n221_));
  NA2        g0199(.A(i_0_), .B(i_5_), .Y(new_new_n222_));
  NAi31      g0200(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n36_), .B(i_13_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n225_));
  NO2        g0203(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n226_));
  NA3        g0204(.A(new_new_n226_), .B(new_new_n225_), .C(new_new_n224_), .Y(new_new_n227_));
  INV        g0205(.A(i_13_), .Y(new_new_n228_));
  NO2        g0206(.A(i_12_), .B(new_new_n228_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n227_), .B(new_new_n223_), .Y(new_new_n230_));
  NA2        g0208(.A(new_new_n230_), .B(new_new_n145_), .Y(new_new_n231_));
  NO2        g0209(.A(i_12_), .B(new_new_n37_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n187_), .B(i_4_), .Y(new_new_n233_));
  NA2        g0211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  OR2        g0212(.A(i_8_), .B(i_7_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n235_), .B(new_new_n87_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n54_), .B(i_1_), .Y(new_new_n237_));
  NA2        g0215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  INV        g0216(.A(i_12_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n45_), .B(new_new_n239_), .Y(new_new_n240_));
  NO3        g0218(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n241_));
  NA2        g0219(.A(i_2_), .B(i_1_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n238_), .B(new_new_n234_), .Y(new_new_n243_));
  NO3        g0221(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n244_));
  NAi21      g0222(.An(i_4_), .B(i_3_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n245_), .B(new_new_n76_), .Y(new_new_n246_));
  NO2        g0224(.A(i_0_), .B(i_6_), .Y(new_new_n247_));
  NOi41      g0225(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n248_));
  NA2        g0226(.A(new_new_n248_), .B(new_new_n247_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n242_), .B(new_new_n187_), .Y(new_new_n250_));
  NAi21      g0228(.An(new_new_n249_), .B(new_new_n250_), .Y(new_new_n251_));
  INV        g0229(.A(new_new_n251_), .Y(new_new_n252_));
  AOI220     g0230(.A0(new_new_n252_), .A1(new_new_n40_), .B0(new_new_n243_), .B1(new_new_n211_), .Y(new_new_n253_));
  NO2        g0231(.A(i_11_), .B(new_new_n228_), .Y(new_new_n254_));
  NOi21      g0232(.An(i_1_), .B(i_6_), .Y(new_new_n255_));
  NAi21      g0233(.An(i_3_), .B(i_7_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n239_), .B(i_9_), .Y(new_new_n257_));
  OR4        g0235(.A(new_new_n257_), .B(new_new_n256_), .C(new_new_n255_), .D(new_new_n190_), .Y(new_new_n258_));
  NO2        g0236(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n259_));
  NO2        g0237(.A(i_12_), .B(i_3_), .Y(new_new_n260_));
  NA2        g0238(.A(new_new_n74_), .B(i_5_), .Y(new_new_n261_));
  NA2        g0239(.A(i_3_), .B(i_9_), .Y(new_new_n262_));
  NAi21      g0240(.An(i_7_), .B(i_10_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n263_), .B(new_new_n262_), .Y(new_new_n264_));
  NA3        g0242(.A(new_new_n264_), .B(new_new_n261_), .C(new_new_n65_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n265_), .B(new_new_n258_), .Y(new_new_n266_));
  NA3        g0244(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n267_));
  INV        g0245(.A(new_new_n146_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n239_), .B(i_13_), .Y(new_new_n269_));
  NO2        g0247(.A(new_new_n269_), .B(new_new_n76_), .Y(new_new_n270_));
  AOI220     g0248(.A0(new_new_n270_), .A1(new_new_n268_), .B0(new_new_n266_), .B1(new_new_n254_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n235_), .B(new_new_n37_), .Y(new_new_n272_));
  NA2        g0250(.A(i_12_), .B(i_6_), .Y(new_new_n273_));
  OR2        g0251(.A(i_13_), .B(i_9_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n245_), .B(i_2_), .Y(new_new_n275_));
  NA2        g0253(.A(new_new_n254_), .B(i_9_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n157_), .B(new_new_n64_), .Y(new_new_n277_));
  NO3        g0255(.A(i_11_), .B(new_new_n228_), .C(new_new_n25_), .Y(new_new_n278_));
  NO2        g0256(.A(new_new_n256_), .B(i_8_), .Y(new_new_n279_));
  NO2        g0257(.A(i_6_), .B(new_new_n49_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n278_), .Y(new_new_n281_));
  NO3        g0259(.A(new_new_n26_), .B(new_new_n87_), .C(i_5_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n272_), .C(new_new_n229_), .Y(new_new_n283_));
  AOI210     g0261(.A0(new_new_n283_), .A1(new_new_n281_), .B0(new_new_n277_), .Y(new_new_n284_));
  INV        g0262(.A(new_new_n284_), .Y(new_new_n285_));
  NA4        g0263(.A(new_new_n285_), .B(new_new_n271_), .C(new_new_n253_), .D(new_new_n231_), .Y(new_new_n286_));
  NO3        g0264(.A(i_12_), .B(new_new_n228_), .C(new_new_n37_), .Y(new_new_n287_));
  INV        g0265(.A(new_new_n287_), .Y(new_new_n288_));
  NA2        g0266(.A(i_8_), .B(new_new_n103_), .Y(new_new_n289_));
  NOi21      g0267(.An(new_new_n166_), .B(new_new_n87_), .Y(new_new_n290_));
  NO3        g0268(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n291_));
  AOI220     g0269(.A0(new_new_n291_), .A1(new_new_n201_), .B0(new_new_n290_), .B1(new_new_n237_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n292_), .B(new_new_n289_), .Y(new_new_n293_));
  NO3        g0271(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n242_), .B(i_0_), .Y(new_new_n295_));
  AOI220     g0273(.A0(new_new_n295_), .A1(new_new_n199_), .B0(new_new_n294_), .B1(new_new_n145_), .Y(new_new_n296_));
  NA2        g0274(.A(new_new_n280_), .B(new_new_n26_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(new_new_n296_), .Y(new_new_n298_));
  NA2        g0276(.A(i_0_), .B(i_1_), .Y(new_new_n299_));
  NO2        g0277(.A(new_new_n299_), .B(i_2_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n60_), .B(i_6_), .Y(new_new_n301_));
  NA3        g0279(.A(new_new_n301_), .B(new_new_n300_), .C(new_new_n166_), .Y(new_new_n302_));
  OAI210     g0280(.A0(new_new_n168_), .A1(new_new_n146_), .B0(new_new_n302_), .Y(new_new_n303_));
  NO3        g0281(.A(new_new_n303_), .B(new_new_n298_), .C(new_new_n293_), .Y(new_new_n304_));
  NO2        g0282(.A(i_3_), .B(i_10_), .Y(new_new_n305_));
  NA3        g0283(.A(new_new_n305_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n306_));
  NO2        g0284(.A(i_2_), .B(new_new_n103_), .Y(new_new_n307_));
  NA2        g0285(.A(i_1_), .B(new_new_n36_), .Y(new_new_n308_));
  NO2        g0286(.A(new_new_n308_), .B(i_8_), .Y(new_new_n309_));
  NA2        g0287(.A(new_new_n309_), .B(new_new_n307_), .Y(new_new_n310_));
  AN2        g0288(.A(i_3_), .B(i_10_), .Y(new_new_n311_));
  NA4        g0289(.A(new_new_n311_), .B(new_new_n203_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n312_));
  NO2        g0290(.A(i_5_), .B(new_new_n37_), .Y(new_new_n313_));
  NO2        g0291(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n314_));
  OR2        g0292(.A(new_new_n310_), .B(new_new_n306_), .Y(new_new_n315_));
  OAI220     g0293(.A0(new_new_n315_), .A1(i_6_), .B0(new_new_n304_), .B1(new_new_n288_), .Y(new_new_n316_));
  NO4        g0294(.A(new_new_n316_), .B(new_new_n286_), .C(new_new_n219_), .D(new_new_n171_), .Y(new_new_n317_));
  NO3        g0295(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n318_));
  NO2        g0296(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n319_));
  NA2        g0297(.A(new_new_n295_), .B(new_new_n319_), .Y(new_new_n320_));
  NO3        g0298(.A(i_6_), .B(new_new_n198_), .C(i_7_), .Y(new_new_n321_));
  NA2        g0299(.A(new_new_n321_), .B(new_new_n203_), .Y(new_new_n322_));
  AOI210     g0300(.A0(new_new_n322_), .A1(new_new_n320_), .B0(new_new_n173_), .Y(new_new_n323_));
  NO2        g0301(.A(i_2_), .B(i_3_), .Y(new_new_n324_));
  OR2        g0302(.A(i_0_), .B(i_5_), .Y(new_new_n325_));
  NA2        g0303(.A(new_new_n222_), .B(new_new_n325_), .Y(new_new_n326_));
  NA4        g0304(.A(new_new_n326_), .B(new_new_n236_), .C(new_new_n324_), .D(i_1_), .Y(new_new_n327_));
  NA3        g0305(.A(new_new_n295_), .B(new_new_n290_), .C(new_new_n115_), .Y(new_new_n328_));
  NAi21      g0306(.An(i_8_), .B(i_7_), .Y(new_new_n329_));
  NO2        g0307(.A(new_new_n329_), .B(i_6_), .Y(new_new_n330_));
  NO2        g0308(.A(new_new_n160_), .B(new_new_n47_), .Y(new_new_n331_));
  NA3        g0309(.A(new_new_n331_), .B(new_new_n330_), .C(new_new_n166_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n332_), .B(new_new_n328_), .C(new_new_n327_), .Y(new_new_n333_));
  OAI210     g0311(.A0(new_new_n333_), .A1(new_new_n323_), .B0(i_4_), .Y(new_new_n334_));
  NO2        g0312(.A(i_12_), .B(i_10_), .Y(new_new_n335_));
  NOi21      g0313(.An(i_5_), .B(i_0_), .Y(new_new_n336_));
  AOI210     g0314(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n103_), .Y(new_new_n337_));
  NO4        g0315(.A(new_new_n337_), .B(new_new_n308_), .C(new_new_n336_), .D(new_new_n131_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n338_), .B(new_new_n335_), .Y(new_new_n339_));
  NO2        g0317(.A(i_6_), .B(i_8_), .Y(new_new_n340_));
  NOi21      g0318(.An(i_0_), .B(i_2_), .Y(new_new_n341_));
  AN2        g0319(.A(new_new_n341_), .B(new_new_n340_), .Y(new_new_n342_));
  NO2        g0320(.A(i_1_), .B(i_7_), .Y(new_new_n343_));
  AO220      g0321(.A0(new_new_n343_), .A1(new_new_n342_), .B0(new_new_n330_), .B1(new_new_n237_), .Y(new_new_n344_));
  NA3        g0322(.A(new_new_n344_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n345_));
  NA3        g0323(.A(new_new_n345_), .B(new_new_n339_), .C(new_new_n334_), .Y(new_new_n346_));
  NO3        g0324(.A(new_new_n235_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n347_));
  NO3        g0325(.A(new_new_n329_), .B(i_2_), .C(i_1_), .Y(new_new_n348_));
  OAI210     g0326(.A0(new_new_n348_), .A1(new_new_n347_), .B0(i_6_), .Y(new_new_n349_));
  NA3        g0327(.A(new_new_n255_), .B(new_new_n307_), .C(new_new_n198_), .Y(new_new_n350_));
  AOI210     g0328(.A0(new_new_n350_), .A1(new_new_n349_), .B0(new_new_n326_), .Y(new_new_n351_));
  NOi21      g0329(.An(new_new_n156_), .B(new_new_n106_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n352_), .B(new_new_n127_), .Y(new_new_n353_));
  OAI210     g0331(.A0(new_new_n353_), .A1(new_new_n351_), .B0(i_3_), .Y(new_new_n354_));
  INV        g0332(.A(new_new_n85_), .Y(new_new_n355_));
  NO2        g0333(.A(new_new_n299_), .B(new_new_n82_), .Y(new_new_n356_));
  NA2        g0334(.A(new_new_n356_), .B(new_new_n135_), .Y(new_new_n357_));
  NO2        g0335(.A(new_new_n94_), .B(new_new_n198_), .Y(new_new_n358_));
  NA2        g0336(.A(new_new_n358_), .B(new_new_n64_), .Y(new_new_n359_));
  AOI210     g0337(.A0(new_new_n359_), .A1(new_new_n357_), .B0(new_new_n355_), .Y(new_new_n360_));
  NO2        g0338(.A(new_new_n198_), .B(i_9_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n210_), .Y(new_new_n362_));
  NO2        g0340(.A(new_new_n362_), .B(new_new_n47_), .Y(new_new_n363_));
  NO3        g0341(.A(new_new_n363_), .B(new_new_n360_), .C(new_new_n298_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n364_), .A1(new_new_n354_), .B0(new_new_n165_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n346_), .A1(new_new_n318_), .B0(new_new_n365_), .Y(new_new_n366_));
  NOi32      g0344(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n367_));
  INV        g0345(.A(new_new_n367_), .Y(new_new_n368_));
  NAi21      g0346(.An(i_0_), .B(i_6_), .Y(new_new_n369_));
  NAi21      g0347(.An(i_1_), .B(i_5_), .Y(new_new_n370_));
  NA2        g0348(.A(new_new_n370_), .B(new_new_n369_), .Y(new_new_n371_));
  NAi41      g0349(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n372_));
  OAI220     g0350(.A0(new_new_n372_), .A1(new_new_n370_), .B0(new_new_n223_), .B1(new_new_n162_), .Y(new_new_n373_));
  AOI210     g0351(.A0(new_new_n372_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n374_));
  NOi32      g0352(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n375_));
  NAi21      g0353(.An(i_6_), .B(i_1_), .Y(new_new_n376_));
  NA3        g0354(.A(new_new_n376_), .B(new_new_n375_), .C(new_new_n47_), .Y(new_new_n377_));
  NO2        g0355(.A(new_new_n377_), .B(i_0_), .Y(new_new_n378_));
  OR3        g0356(.A(new_new_n378_), .B(new_new_n374_), .C(new_new_n373_), .Y(new_new_n379_));
  NO2        g0357(.A(i_1_), .B(new_new_n103_), .Y(new_new_n380_));
  NAi21      g0358(.An(i_3_), .B(i_4_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n381_), .B(i_9_), .Y(new_new_n382_));
  AN2        g0360(.A(i_6_), .B(i_7_), .Y(new_new_n383_));
  OAI210     g0361(.A0(new_new_n383_), .A1(new_new_n380_), .B0(new_new_n382_), .Y(new_new_n384_));
  NA2        g0362(.A(i_2_), .B(i_7_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n381_), .B(i_10_), .Y(new_new_n386_));
  NA3        g0364(.A(new_new_n386_), .B(new_new_n385_), .C(new_new_n247_), .Y(new_new_n387_));
  AOI210     g0365(.A0(new_new_n387_), .A1(new_new_n384_), .B0(new_new_n190_), .Y(new_new_n388_));
  AOI210     g0366(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n389_));
  OAI210     g0367(.A0(new_new_n389_), .A1(new_new_n193_), .B0(new_new_n386_), .Y(new_new_n390_));
  AOI220     g0368(.A0(new_new_n386_), .A1(new_new_n343_), .B0(new_new_n241_), .B1(new_new_n193_), .Y(new_new_n391_));
  AOI210     g0369(.A0(new_new_n391_), .A1(new_new_n390_), .B0(i_5_), .Y(new_new_n392_));
  NO4        g0370(.A(new_new_n392_), .B(new_new_n388_), .C(new_new_n379_), .D(new_new_n1079_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n393_), .B(new_new_n368_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n395_));
  AN2        g0373(.A(i_12_), .B(i_5_), .Y(new_new_n396_));
  NO2        g0374(.A(i_4_), .B(new_new_n26_), .Y(new_new_n397_));
  NA2        g0375(.A(new_new_n397_), .B(new_new_n396_), .Y(new_new_n398_));
  NO2        g0376(.A(i_11_), .B(i_6_), .Y(new_new_n399_));
  NA3        g0377(.A(new_new_n399_), .B(new_new_n331_), .C(new_new_n228_), .Y(new_new_n400_));
  NO2        g0378(.A(new_new_n400_), .B(new_new_n398_), .Y(new_new_n401_));
  NO2        g0379(.A(new_new_n245_), .B(i_5_), .Y(new_new_n402_));
  NO2        g0380(.A(i_5_), .B(i_10_), .Y(new_new_n403_));
  AOI220     g0381(.A0(new_new_n403_), .A1(new_new_n275_), .B0(new_new_n402_), .B1(new_new_n203_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n147_), .B(new_new_n46_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n405_), .B(new_new_n404_), .Y(new_new_n406_));
  OAI210     g0384(.A0(new_new_n406_), .A1(new_new_n401_), .B0(new_new_n395_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n408_));
  NO3        g0386(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n409_));
  NO2        g0387(.A(i_3_), .B(new_new_n103_), .Y(new_new_n410_));
  NA4        g0388(.A(new_new_n305_), .B(new_new_n92_), .C(new_new_n76_), .D(new_new_n55_), .Y(new_new_n411_));
  NO2        g0389(.A(i_11_), .B(i_12_), .Y(new_new_n412_));
  NA2        g0390(.A(new_new_n412_), .B(new_new_n36_), .Y(new_new_n413_));
  NO2        g0391(.A(new_new_n411_), .B(new_new_n413_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n403_), .B(new_new_n239_), .Y(new_new_n415_));
  NA3        g0393(.A(new_new_n115_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n416_));
  NO2        g0394(.A(new_new_n416_), .B(new_new_n223_), .Y(new_new_n417_));
  NAi21      g0395(.An(i_13_), .B(i_0_), .Y(new_new_n418_));
  NO2        g0396(.A(new_new_n418_), .B(new_new_n242_), .Y(new_new_n419_));
  OAI210     g0397(.A0(new_new_n417_), .A1(new_new_n414_), .B0(new_new_n419_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n420_), .B(new_new_n407_), .Y(new_new_n421_));
  NO3        g0399(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n422_));
  NO2        g0400(.A(i_0_), .B(i_11_), .Y(new_new_n423_));
  INV        g0401(.A(i_5_), .Y(new_new_n424_));
  AN2        g0402(.A(i_1_), .B(i_6_), .Y(new_new_n425_));
  NOi21      g0403(.An(i_2_), .B(i_12_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n426_), .B(new_new_n425_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(new_new_n424_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n145_), .B(i_9_), .Y(new_new_n429_));
  NO2        g0407(.A(new_new_n429_), .B(i_4_), .Y(new_new_n430_));
  NA2        g0408(.A(new_new_n428_), .B(new_new_n430_), .Y(new_new_n431_));
  NAi21      g0409(.An(i_9_), .B(i_4_), .Y(new_new_n432_));
  OR2        g0410(.A(i_13_), .B(i_10_), .Y(new_new_n433_));
  NO3        g0411(.A(new_new_n433_), .B(new_new_n120_), .C(new_new_n432_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n176_), .B(new_new_n126_), .Y(new_new_n435_));
  OR2        g0413(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n287_), .B(new_new_n437_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n280_), .B(new_new_n215_), .Y(new_new_n439_));
  OAI220     g0417(.A0(new_new_n439_), .A1(new_new_n436_), .B0(new_new_n438_), .B1(new_new_n352_), .Y(new_new_n440_));
  INV        g0418(.A(new_new_n440_), .Y(new_new_n441_));
  AOI210     g0419(.A0(new_new_n441_), .A1(new_new_n431_), .B0(new_new_n26_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n328_), .B(new_new_n327_), .Y(new_new_n443_));
  AOI220     g0421(.A0(new_new_n301_), .A1(new_new_n291_), .B0(new_new_n295_), .B1(new_new_n319_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(new_new_n173_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n187_), .B(new_new_n87_), .Y(new_new_n446_));
  AOI220     g0424(.A0(new_new_n446_), .A1(new_new_n300_), .B0(new_new_n282_), .B1(new_new_n215_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(new_new_n289_), .Y(new_new_n448_));
  NO3        g0426(.A(new_new_n448_), .B(new_new_n445_), .C(new_new_n443_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n201_), .B(new_new_n98_), .Y(new_new_n450_));
  NA3        g0428(.A(new_new_n331_), .B(new_new_n166_), .C(new_new_n87_), .Y(new_new_n451_));
  AOI210     g0429(.A0(new_new_n451_), .A1(new_new_n450_), .B0(new_new_n329_), .Y(new_new_n452_));
  NA2        g0430(.A(new_new_n198_), .B(i_10_), .Y(new_new_n453_));
  NA3        g0431(.A(new_new_n261_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n301_), .B(new_new_n237_), .Y(new_new_n455_));
  OAI220     g0433(.A0(new_new_n455_), .A1(new_new_n187_), .B0(new_new_n454_), .B1(new_new_n453_), .Y(new_new_n456_));
  NO2        g0434(.A(i_3_), .B(new_new_n49_), .Y(new_new_n457_));
  NA3        g0435(.A(new_new_n343_), .B(new_new_n342_), .C(new_new_n457_), .Y(new_new_n458_));
  NA2        g0436(.A(new_new_n321_), .B(new_new_n326_), .Y(new_new_n459_));
  OAI210     g0437(.A0(new_new_n459_), .A1(new_new_n194_), .B0(new_new_n458_), .Y(new_new_n460_));
  NO3        g0438(.A(new_new_n460_), .B(new_new_n456_), .C(new_new_n452_), .Y(new_new_n461_));
  AOI210     g0439(.A0(new_new_n461_), .A1(new_new_n449_), .B0(new_new_n276_), .Y(new_new_n462_));
  NO4        g0440(.A(new_new_n462_), .B(new_new_n442_), .C(new_new_n421_), .D(new_new_n394_), .Y(new_new_n463_));
  NO2        g0441(.A(new_new_n64_), .B(i_4_), .Y(new_new_n464_));
  NO2        g0442(.A(new_new_n74_), .B(i_13_), .Y(new_new_n465_));
  NO2        g0443(.A(i_10_), .B(i_9_), .Y(new_new_n466_));
  NAi21      g0444(.An(i_12_), .B(i_8_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n467_), .B(i_3_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n314_), .B(i_0_), .Y(new_new_n469_));
  NO3        g0447(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n273_), .B(new_new_n99_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n471_), .B(new_new_n470_), .Y(new_new_n472_));
  NA2        g0450(.A(i_8_), .B(i_9_), .Y(new_new_n473_));
  AOI210     g0451(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n474_));
  OR2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n287_), .B(new_new_n210_), .Y(new_new_n476_));
  NO2        g0454(.A(new_new_n476_), .B(new_new_n475_), .Y(new_new_n477_));
  NA2        g0455(.A(new_new_n254_), .B(new_new_n313_), .Y(new_new_n478_));
  NO3        g0456(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n479_));
  INV        g0457(.A(new_new_n479_), .Y(new_new_n480_));
  NA3        g0458(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n481_));
  NA4        g0459(.A(new_new_n148_), .B(new_new_n118_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n482_));
  OAI220     g0460(.A0(new_new_n482_), .A1(new_new_n481_), .B0(new_new_n480_), .B1(new_new_n478_), .Y(new_new_n483_));
  NO2        g0461(.A(new_new_n483_), .B(new_new_n477_), .Y(new_new_n484_));
  NA2        g0462(.A(new_new_n300_), .B(new_new_n110_), .Y(new_new_n485_));
  OR2        g0463(.A(new_new_n485_), .B(new_new_n212_), .Y(new_new_n486_));
  BUFFER     g0464(.A(new_new_n302_), .Y(new_new_n487_));
  OA220      g0465(.A0(new_new_n487_), .A1(new_new_n165_), .B0(new_new_n486_), .B1(new_new_n234_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n98_), .B(i_13_), .Y(new_new_n489_));
  NO2        g0467(.A(i_2_), .B(i_13_), .Y(new_new_n490_));
  NO3        g0468(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n491_));
  NO2        g0469(.A(i_6_), .B(i_7_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n492_), .B(new_new_n491_), .Y(new_new_n493_));
  NO2        g0471(.A(i_11_), .B(i_1_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n74_), .B(i_3_), .Y(new_new_n495_));
  OR2        g0473(.A(i_11_), .B(i_8_), .Y(new_new_n496_));
  NOi21      g0474(.An(i_2_), .B(i_7_), .Y(new_new_n497_));
  NAi31      g0475(.An(new_new_n496_), .B(new_new_n497_), .C(new_new_n495_), .Y(new_new_n498_));
  NO2        g0476(.A(new_new_n433_), .B(i_6_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n464_), .C(new_new_n76_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n500_), .B(new_new_n498_), .Y(new_new_n501_));
  NO2        g0479(.A(i_3_), .B(new_new_n198_), .Y(new_new_n502_));
  NO2        g0480(.A(i_6_), .B(i_10_), .Y(new_new_n503_));
  NA4        g0481(.A(new_new_n503_), .B(new_new_n318_), .C(new_new_n502_), .D(new_new_n239_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n504_), .B(new_new_n158_), .Y(new_new_n505_));
  NA3        g0483(.A(new_new_n248_), .B(new_new_n175_), .C(new_new_n135_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n507_));
  NO2        g0485(.A(new_new_n160_), .B(i_3_), .Y(new_new_n508_));
  NAi31      g0486(.An(new_new_n507_), .B(new_new_n508_), .C(new_new_n229_), .Y(new_new_n509_));
  NA3        g0487(.A(new_new_n408_), .B(new_new_n183_), .C(new_new_n152_), .Y(new_new_n510_));
  NA3        g0488(.A(new_new_n510_), .B(new_new_n509_), .C(new_new_n506_), .Y(new_new_n511_));
  NO3        g0489(.A(new_new_n511_), .B(new_new_n505_), .C(new_new_n501_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n470_), .B(new_new_n396_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n479_), .B(new_new_n403_), .Y(new_new_n514_));
  NO2        g0492(.A(new_new_n514_), .B(new_new_n227_), .Y(new_new_n515_));
  NAi21      g0493(.An(new_new_n221_), .B(new_new_n412_), .Y(new_new_n516_));
  NO2        g0494(.A(new_new_n26_), .B(i_5_), .Y(new_new_n517_));
  NO2        g0495(.A(i_0_), .B(new_new_n87_), .Y(new_new_n518_));
  NA3        g0496(.A(new_new_n518_), .B(new_new_n517_), .C(new_new_n145_), .Y(new_new_n519_));
  OR3        g0497(.A(new_new_n308_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n520_));
  NO2        g0498(.A(new_new_n520_), .B(new_new_n519_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n27_), .B(i_10_), .Y(new_new_n522_));
  NA2        g0500(.A(new_new_n318_), .B(new_new_n241_), .Y(new_new_n523_));
  OAI220     g0501(.A0(new_new_n523_), .A1(new_new_n454_), .B0(new_new_n522_), .B1(new_new_n489_), .Y(new_new_n524_));
  NA4        g0502(.A(new_new_n311_), .B(new_new_n226_), .C(new_new_n74_), .D(new_new_n239_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n493_), .Y(new_new_n526_));
  NO4        g0504(.A(new_new_n526_), .B(new_new_n524_), .C(new_new_n521_), .D(new_new_n515_), .Y(new_new_n527_));
  NA4        g0505(.A(new_new_n527_), .B(new_new_n512_), .C(new_new_n488_), .D(new_new_n484_), .Y(new_new_n528_));
  NA3        g0506(.A(new_new_n311_), .B(new_new_n180_), .C(new_new_n178_), .Y(new_new_n529_));
  OAI210     g0507(.A0(new_new_n306_), .A1(new_new_n185_), .B0(new_new_n529_), .Y(new_new_n530_));
  AN2        g0508(.A(new_new_n291_), .B(new_new_n236_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n531_), .B(new_new_n530_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n318_), .B(new_new_n167_), .Y(new_new_n533_));
  OAI210     g0511(.A0(new_new_n533_), .A1(new_new_n234_), .B0(new_new_n312_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n534_), .B(new_new_n330_), .Y(new_new_n535_));
  NA2        g0513(.A(new_new_n396_), .B(new_new_n228_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n367_), .B(new_new_n74_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n383_), .B(new_new_n375_), .Y(new_new_n538_));
  OR2        g0516(.A(new_new_n536_), .B(new_new_n538_), .Y(new_new_n539_));
  NO2        g0517(.A(new_new_n36_), .B(i_8_), .Y(new_new_n540_));
  NAi41      g0518(.An(new_new_n537_), .B(new_new_n503_), .C(new_new_n540_), .D(new_new_n47_), .Y(new_new_n541_));
  AOI210     g0519(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n434_), .Y(new_new_n542_));
  NA3        g0520(.A(new_new_n542_), .B(new_new_n541_), .C(new_new_n539_), .Y(new_new_n543_));
  INV        g0521(.A(new_new_n543_), .Y(new_new_n544_));
  INV        g0522(.A(new_new_n137_), .Y(new_new_n545_));
  AOI210     g0523(.A0(new_new_n199_), .A1(i_9_), .B0(new_new_n272_), .Y(new_new_n546_));
  NO2        g0524(.A(new_new_n546_), .B(new_new_n204_), .Y(new_new_n547_));
  OR2        g0525(.A(new_new_n187_), .B(i_4_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n548_), .B(new_new_n87_), .Y(new_new_n549_));
  AOI220     g0527(.A0(new_new_n549_), .A1(new_new_n547_), .B0(new_new_n545_), .B1(new_new_n435_), .Y(new_new_n550_));
  NA4        g0528(.A(new_new_n550_), .B(new_new_n544_), .C(new_new_n535_), .D(new_new_n532_), .Y(new_new_n551_));
  NA2        g0529(.A(new_new_n402_), .B(new_new_n300_), .Y(new_new_n552_));
  OAI210     g0530(.A0(new_new_n398_), .A1(new_new_n172_), .B0(new_new_n552_), .Y(new_new_n553_));
  NO2        g0531(.A(i_12_), .B(new_new_n198_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n228_), .Y(new_new_n555_));
  NA3        g0533(.A(new_new_n503_), .B(new_new_n178_), .C(new_new_n27_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n556_), .B(new_new_n555_), .Y(new_new_n557_));
  NOi31      g0535(.An(new_new_n321_), .B(new_new_n433_), .C(new_new_n38_), .Y(new_new_n558_));
  OAI210     g0536(.A0(new_new_n558_), .A1(new_new_n557_), .B0(new_new_n553_), .Y(new_new_n559_));
  NO2        g0537(.A(i_8_), .B(i_7_), .Y(new_new_n560_));
  OAI210     g0538(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n561_));
  NA2        g0539(.A(new_new_n561_), .B(new_new_n226_), .Y(new_new_n562_));
  AOI220     g0540(.A0(new_new_n331_), .A1(new_new_n40_), .B0(new_new_n237_), .B1(new_new_n211_), .Y(new_new_n563_));
  OAI220     g0541(.A0(new_new_n563_), .A1(new_new_n548_), .B0(new_new_n562_), .B1(new_new_n245_), .Y(new_new_n564_));
  NA2        g0542(.A(new_new_n45_), .B(i_10_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n565_), .B(i_6_), .Y(new_new_n566_));
  NA3        g0544(.A(new_new_n566_), .B(new_new_n564_), .C(new_new_n560_), .Y(new_new_n567_));
  NOi31      g0545(.An(new_new_n295_), .B(new_new_n306_), .C(new_new_n185_), .Y(new_new_n568_));
  NO2        g0546(.A(new_new_n160_), .B(i_5_), .Y(new_new_n569_));
  NA2        g0547(.A(new_new_n568_), .B(new_new_n479_), .Y(new_new_n570_));
  NA3        g0548(.A(new_new_n570_), .B(new_new_n567_), .C(new_new_n559_), .Y(new_new_n571_));
  NA3        g0549(.A(new_new_n222_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n572_));
  NA2        g0550(.A(new_new_n287_), .B(new_new_n85_), .Y(new_new_n573_));
  AOI210     g0551(.A0(new_new_n572_), .A1(new_new_n357_), .B0(new_new_n573_), .Y(new_new_n574_));
  NA2        g0552(.A(new_new_n301_), .B(new_new_n291_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n575_), .B(new_new_n177_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n226_), .B(new_new_n225_), .Y(new_new_n577_));
  NA2        g0555(.A(new_new_n466_), .B(new_new_n224_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n577_), .B(new_new_n578_), .Y(new_new_n579_));
  AOI210     g0557(.A0(new_new_n376_), .A1(new_new_n47_), .B0(new_new_n380_), .Y(new_new_n580_));
  NA2        g0558(.A(i_0_), .B(new_new_n49_), .Y(new_new_n581_));
  NA3        g0559(.A(new_new_n554_), .B(new_new_n278_), .C(new_new_n581_), .Y(new_new_n582_));
  NO2        g0560(.A(new_new_n580_), .B(new_new_n582_), .Y(new_new_n583_));
  NO4        g0561(.A(new_new_n583_), .B(new_new_n579_), .C(new_new_n576_), .D(new_new_n574_), .Y(new_new_n584_));
  NO4        g0562(.A(new_new_n255_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n585_));
  NO3        g0563(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n235_), .B(new_new_n36_), .Y(new_new_n587_));
  AN2        g0565(.A(new_new_n587_), .B(new_new_n586_), .Y(new_new_n588_));
  OA210      g0566(.A0(new_new_n588_), .A1(new_new_n585_), .B0(new_new_n367_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n433_), .B(i_1_), .Y(new_new_n590_));
  NOi31      g0568(.An(new_new_n590_), .B(new_new_n471_), .C(new_new_n74_), .Y(new_new_n591_));
  AN4        g0569(.A(new_new_n591_), .B(new_new_n430_), .C(new_new_n517_), .D(i_2_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n444_), .B(new_new_n181_), .Y(new_new_n593_));
  NO3        g0571(.A(new_new_n593_), .B(new_new_n592_), .C(new_new_n589_), .Y(new_new_n594_));
  NOi21      g0572(.An(i_10_), .B(i_6_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n597_));
  NA2        g0575(.A(new_new_n321_), .B(new_new_n167_), .Y(new_new_n598_));
  AOI220     g0576(.A0(new_new_n598_), .A1(new_new_n455_), .B0(new_new_n188_), .B1(new_new_n186_), .Y(new_new_n599_));
  INV        g0577(.A(new_new_n599_), .Y(new_new_n600_));
  NO2        g0578(.A(i_12_), .B(new_new_n87_), .Y(new_new_n601_));
  NA2        g0579(.A(new_new_n178_), .B(i_0_), .Y(new_new_n602_));
  NO3        g0580(.A(new_new_n602_), .B(new_new_n349_), .C(new_new_n306_), .Y(new_new_n603_));
  OR2        g0581(.A(i_2_), .B(i_5_), .Y(new_new_n604_));
  OR2        g0582(.A(new_new_n604_), .B(new_new_n425_), .Y(new_new_n605_));
  AOI210     g0583(.A0(new_new_n385_), .A1(new_new_n247_), .B0(new_new_n203_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n606_), .A1(new_new_n605_), .B0(new_new_n516_), .Y(new_new_n607_));
  NO2        g0585(.A(new_new_n607_), .B(new_new_n603_), .Y(new_new_n608_));
  NA4        g0586(.A(new_new_n608_), .B(new_new_n600_), .C(new_new_n594_), .D(new_new_n584_), .Y(new_new_n609_));
  NO4        g0587(.A(new_new_n609_), .B(new_new_n571_), .C(new_new_n551_), .D(new_new_n528_), .Y(new_new_n610_));
  NA4        g0588(.A(new_new_n610_), .B(new_new_n463_), .C(new_new_n366_), .D(new_new_n317_), .Y(mai7));
  NO2        g0589(.A(new_new_n94_), .B(new_new_n55_), .Y(new_new_n612_));
  NA2        g0590(.A(new_new_n503_), .B(new_new_n85_), .Y(new_new_n613_));
  NA2        g0591(.A(i_11_), .B(new_new_n198_), .Y(new_new_n614_));
  NA2        g0592(.A(new_new_n147_), .B(new_new_n614_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n615_), .B(new_new_n613_), .Y(new_new_n616_));
  NA3        g0594(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n617_));
  NO2        g0595(.A(new_new_n239_), .B(i_4_), .Y(new_new_n618_));
  NA2        g0596(.A(new_new_n618_), .B(i_8_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n107_), .B(new_new_n617_), .Y(new_new_n620_));
  NA2        g0598(.A(i_2_), .B(new_new_n87_), .Y(new_new_n621_));
  OAI210     g0599(.A0(new_new_n88_), .A1(new_new_n208_), .B0(new_new_n209_), .Y(new_new_n622_));
  NO2        g0600(.A(i_7_), .B(new_new_n37_), .Y(new_new_n623_));
  NA2        g0601(.A(i_4_), .B(i_8_), .Y(new_new_n624_));
  AOI210     g0602(.A0(new_new_n624_), .A1(new_new_n311_), .B0(new_new_n623_), .Y(new_new_n625_));
  OAI220     g0603(.A0(new_new_n625_), .A1(new_new_n621_), .B0(new_new_n622_), .B1(i_13_), .Y(new_new_n626_));
  NO4        g0604(.A(new_new_n626_), .B(new_new_n620_), .C(new_new_n616_), .D(new_new_n612_), .Y(new_new_n627_));
  AOI210     g0605(.A0(new_new_n131_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n628_));
  AOI210     g0606(.A0(new_new_n628_), .A1(new_new_n239_), .B0(new_new_n164_), .Y(new_new_n629_));
  OR2        g0607(.A(i_6_), .B(i_10_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n630_), .B(new_new_n23_), .Y(new_new_n631_));
  OR3        g0609(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n632_));
  NO3        g0610(.A(new_new_n632_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n633_));
  INV        g0611(.A(new_new_n205_), .Y(new_new_n634_));
  OR2        g0612(.A(new_new_n629_), .B(new_new_n274_), .Y(new_new_n635_));
  AOI210     g0613(.A0(new_new_n635_), .A1(new_new_n627_), .B0(new_new_n64_), .Y(new_new_n636_));
  NOi21      g0614(.An(i_11_), .B(i_7_), .Y(new_new_n637_));
  AO210      g0615(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n638_));
  NO2        g0616(.A(new_new_n638_), .B(new_new_n637_), .Y(new_new_n639_));
  NA2        g0617(.A(new_new_n639_), .B(new_new_n211_), .Y(new_new_n640_));
  NA3        g0618(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n641_));
  NO2        g0619(.A(new_new_n640_), .B(new_new_n64_), .Y(new_new_n642_));
  OR2        g0620(.A(new_new_n391_), .B(new_new_n41_), .Y(new_new_n643_));
  NO3        g0621(.A(new_new_n263_), .B(new_new_n213_), .C(new_new_n614_), .Y(new_new_n644_));
  OAI210     g0622(.A0(new_new_n644_), .A1(new_new_n229_), .B0(new_new_n64_), .Y(new_new_n645_));
  NA2        g0623(.A(new_new_n426_), .B(new_new_n31_), .Y(new_new_n646_));
  OR2        g0624(.A(new_new_n213_), .B(new_new_n110_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n647_), .B(new_new_n646_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n64_), .B(i_9_), .Y(new_new_n649_));
  NO2        g0627(.A(new_new_n649_), .B(i_4_), .Y(new_new_n650_));
  NA2        g0628(.A(new_new_n650_), .B(new_new_n648_), .Y(new_new_n651_));
  NO2        g0629(.A(i_1_), .B(i_12_), .Y(new_new_n652_));
  NA3        g0630(.A(new_new_n651_), .B(new_new_n645_), .C(new_new_n643_), .Y(new_new_n653_));
  OAI210     g0631(.A0(new_new_n653_), .A1(new_new_n642_), .B0(i_6_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n641_), .B(new_new_n110_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n655_), .B(new_new_n601_), .Y(new_new_n656_));
  NO2        g0634(.A(i_6_), .B(i_11_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n656_), .B(new_new_n472_), .Y(new_new_n658_));
  NO4        g0636(.A(new_new_n220_), .B(new_new_n131_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n659_), .B(new_new_n649_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n239_), .B(i_6_), .Y(new_new_n661_));
  NO3        g0639(.A(new_new_n630_), .B(new_new_n235_), .C(new_new_n23_), .Y(new_new_n662_));
  AOI210     g0640(.A0(i_1_), .A1(new_new_n264_), .B0(new_new_n662_), .Y(new_new_n663_));
  OAI210     g0641(.A0(new_new_n663_), .A1(new_new_n45_), .B0(new_new_n660_), .Y(new_new_n664_));
  NA3        g0642(.A(new_new_n560_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n141_), .B(i_9_), .Y(new_new_n666_));
  NA3        g0644(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n47_), .B(i_1_), .Y(new_new_n668_));
  NA3        g0646(.A(new_new_n668_), .B(new_new_n273_), .C(new_new_n45_), .Y(new_new_n669_));
  OAI220     g0647(.A0(new_new_n669_), .A1(new_new_n667_), .B0(new_new_n666_), .B1(new_new_n1078_), .Y(new_new_n670_));
  NA3        g0648(.A(new_new_n649_), .B(new_new_n324_), .C(i_6_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n671_), .B(new_new_n23_), .Y(new_new_n672_));
  AOI210     g0650(.A0(new_new_n494_), .A1(new_new_n437_), .B0(new_new_n244_), .Y(new_new_n673_));
  NO2        g0651(.A(new_new_n673_), .B(new_new_n621_), .Y(new_new_n674_));
  NAi21      g0652(.An(new_new_n665_), .B(new_new_n93_), .Y(new_new_n675_));
  NA2        g0653(.A(new_new_n668_), .B(new_new_n273_), .Y(new_new_n676_));
  NO2        g0654(.A(i_11_), .B(new_new_n37_), .Y(new_new_n677_));
  NA2        g0655(.A(new_new_n677_), .B(new_new_n24_), .Y(new_new_n678_));
  OAI210     g0656(.A0(new_new_n678_), .A1(new_new_n676_), .B0(new_new_n675_), .Y(new_new_n679_));
  OR4        g0657(.A(new_new_n679_), .B(new_new_n674_), .C(new_new_n672_), .D(new_new_n670_), .Y(new_new_n680_));
  NO3        g0658(.A(new_new_n680_), .B(new_new_n664_), .C(new_new_n658_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n239_), .B(new_new_n103_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n682_), .B(new_new_n637_), .Y(new_new_n683_));
  NA2        g0661(.A(new_new_n683_), .B(i_1_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n684_), .B(new_new_n632_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n432_), .B(new_new_n87_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n685_), .B(new_new_n47_), .Y(new_new_n687_));
  NA2        g0665(.A(i_3_), .B(new_new_n198_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(new_new_n117_), .Y(new_new_n689_));
  AN2        g0667(.A(new_new_n689_), .B(new_new_n566_), .Y(new_new_n690_));
  NO2        g0668(.A(new_new_n235_), .B(new_new_n45_), .Y(new_new_n691_));
  NO3        g0669(.A(new_new_n691_), .B(new_new_n314_), .C(new_new_n240_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n693_), .B(i_6_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n87_), .B(i_9_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n64_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n652_), .Y(new_new_n697_));
  NO4        g0675(.A(new_new_n697_), .B(new_new_n694_), .C(new_new_n692_), .D(i_4_), .Y(new_new_n698_));
  NA2        g0676(.A(i_1_), .B(i_3_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n473_), .B(new_new_n94_), .Y(new_new_n700_));
  AOI210     g0678(.A0(new_new_n691_), .A1(new_new_n595_), .B0(new_new_n700_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n701_), .B(new_new_n699_), .Y(new_new_n702_));
  NO3        g0680(.A(new_new_n702_), .B(new_new_n698_), .C(new_new_n690_), .Y(new_new_n703_));
  NA4        g0681(.A(new_new_n703_), .B(new_new_n687_), .C(new_new_n681_), .D(new_new_n654_), .Y(new_new_n704_));
  NO3        g0682(.A(new_new_n496_), .B(i_3_), .C(i_7_), .Y(new_new_n705_));
  NOi21      g0683(.An(new_new_n705_), .B(i_10_), .Y(new_new_n706_));
  OA210      g0684(.A0(new_new_n706_), .A1(new_new_n248_), .B0(new_new_n87_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n383_), .B(new_new_n382_), .Y(new_new_n708_));
  NA3        g0686(.A(new_new_n503_), .B(new_new_n540_), .C(new_new_n47_), .Y(new_new_n709_));
  NO3        g0687(.A(new_new_n497_), .B(new_new_n624_), .C(new_new_n87_), .Y(new_new_n710_));
  NA2        g0688(.A(new_new_n710_), .B(new_new_n25_), .Y(new_new_n711_));
  NA3        g0689(.A(new_new_n711_), .B(new_new_n709_), .C(new_new_n708_), .Y(new_new_n712_));
  OAI210     g0690(.A0(new_new_n712_), .A1(new_new_n707_), .B0(i_1_), .Y(new_new_n713_));
  AOI210     g0691(.A0(new_new_n273_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n714_));
  NO2        g0692(.A(new_new_n381_), .B(i_2_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n715_), .B(new_new_n714_), .Y(new_new_n716_));
  OAI210     g0694(.A0(new_new_n671_), .A1(new_new_n467_), .B0(new_new_n716_), .Y(new_new_n717_));
  INV        g0695(.A(new_new_n717_), .Y(new_new_n718_));
  AOI210     g0696(.A0(new_new_n718_), .A1(new_new_n713_), .B0(i_13_), .Y(new_new_n719_));
  OR2        g0697(.A(i_11_), .B(i_7_), .Y(new_new_n720_));
  AOI210     g0698(.A0(new_new_n667_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n721_));
  NO2        g0699(.A(new_new_n497_), .B(new_new_n24_), .Y(new_new_n722_));
  AOI220     g0700(.A0(new_new_n722_), .A1(new_new_n686_), .B0(new_new_n248_), .B1(new_new_n134_), .Y(new_new_n723_));
  OAI220     g0701(.A0(new_new_n723_), .A1(new_new_n41_), .B0(new_new_n1077_), .B1(new_new_n94_), .Y(new_new_n724_));
  INV        g0702(.A(new_new_n724_), .Y(new_new_n725_));
  INV        g0703(.A(new_new_n117_), .Y(new_new_n726_));
  AOI220     g0704(.A0(new_new_n726_), .A1(new_new_n73_), .B0(new_new_n399_), .B1(new_new_n668_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n727_), .B(new_new_n245_), .Y(new_new_n728_));
  AOI210     g0706(.A0(new_new_n467_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n729_));
  NOi31      g0707(.An(new_new_n729_), .B(new_new_n613_), .C(new_new_n45_), .Y(new_new_n730_));
  NA2        g0708(.A(new_new_n130_), .B(i_13_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n667_), .B(new_new_n117_), .Y(new_new_n732_));
  INV        g0710(.A(new_new_n732_), .Y(new_new_n733_));
  OAI220     g0711(.A0(new_new_n733_), .A1(new_new_n72_), .B0(new_new_n731_), .B1(new_new_n714_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n26_), .B(new_new_n198_), .Y(new_new_n735_));
  NA2        g0713(.A(new_new_n735_), .B(i_7_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n497_), .B(new_new_n239_), .C(new_new_n87_), .Y(new_new_n737_));
  NA2        g0715(.A(new_new_n737_), .B(new_new_n736_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n399_), .A1(new_new_n668_), .B0(new_new_n93_), .B1(new_new_n104_), .Y(new_new_n739_));
  OAI220     g0717(.A0(new_new_n739_), .A1(new_new_n619_), .B0(new_new_n738_), .B1(new_new_n634_), .Y(new_new_n740_));
  NO4        g0718(.A(new_new_n740_), .B(new_new_n734_), .C(new_new_n730_), .D(new_new_n728_), .Y(new_new_n741_));
  OR2        g0719(.A(i_11_), .B(i_6_), .Y(new_new_n742_));
  NA3        g0720(.A(new_new_n618_), .B(new_new_n735_), .C(i_7_), .Y(new_new_n743_));
  AOI210     g0721(.A0(new_new_n743_), .A1(new_new_n733_), .B0(new_new_n742_), .Y(new_new_n744_));
  NA3        g0722(.A(new_new_n426_), .B(new_new_n623_), .C(new_new_n99_), .Y(new_new_n745_));
  NA2        g0723(.A(new_new_n657_), .B(i_13_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n104_), .B(new_new_n735_), .Y(new_new_n747_));
  NAi21      g0725(.An(i_11_), .B(i_12_), .Y(new_new_n748_));
  NOi41      g0726(.An(new_new_n113_), .B(new_new_n748_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n749_));
  NO3        g0727(.A(new_new_n497_), .B(new_new_n601_), .C(new_new_n624_), .Y(new_new_n750_));
  AOI220     g0728(.A0(new_new_n750_), .A1(new_new_n318_), .B0(new_new_n749_), .B1(new_new_n747_), .Y(new_new_n751_));
  NA3        g0729(.A(new_new_n751_), .B(new_new_n746_), .C(new_new_n745_), .Y(new_new_n752_));
  OAI210     g0730(.A0(new_new_n752_), .A1(new_new_n744_), .B0(new_new_n64_), .Y(new_new_n753_));
  NO2        g0731(.A(i_2_), .B(i_12_), .Y(new_new_n754_));
  NA2        g0732(.A(new_new_n380_), .B(new_new_n754_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n382_), .B(new_new_n380_), .Y(new_new_n756_));
  NO2        g0734(.A(new_new_n131_), .B(i_2_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n757_), .B(new_new_n652_), .Y(new_new_n758_));
  NA3        g0736(.A(new_new_n758_), .B(new_new_n756_), .C(new_new_n755_), .Y(new_new_n759_));
  NA3        g0737(.A(new_new_n759_), .B(new_new_n46_), .C(new_new_n228_), .Y(new_new_n760_));
  NA4        g0738(.A(new_new_n760_), .B(new_new_n753_), .C(new_new_n741_), .D(new_new_n725_), .Y(new_new_n761_));
  OR4        g0739(.A(new_new_n761_), .B(new_new_n719_), .C(new_new_n704_), .D(new_new_n636_), .Y(mai5));
  NA2        g0740(.A(new_new_n683_), .B(new_new_n275_), .Y(new_new_n763_));
  AN2        g0741(.A(new_new_n24_), .B(i_10_), .Y(new_new_n764_));
  NA3        g0742(.A(new_new_n764_), .B(new_new_n754_), .C(new_new_n110_), .Y(new_new_n765_));
  NO2        g0743(.A(new_new_n619_), .B(i_11_), .Y(new_new_n766_));
  NA2        g0744(.A(new_new_n88_), .B(new_new_n766_), .Y(new_new_n767_));
  NA3        g0745(.A(new_new_n767_), .B(new_new_n765_), .C(new_new_n763_), .Y(new_new_n768_));
  NO3        g0746(.A(i_11_), .B(new_new_n239_), .C(i_13_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n770_));
  NA2        g0748(.A(i_12_), .B(i_8_), .Y(new_new_n771_));
  OAI210     g0749(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n771_), .Y(new_new_n772_));
  INV        g0750(.A(new_new_n466_), .Y(new_new_n773_));
  AOI220     g0751(.A0(new_new_n324_), .A1(new_new_n597_), .B0(new_new_n772_), .B1(new_new_n770_), .Y(new_new_n774_));
  INV        g0752(.A(new_new_n774_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n775_), .B(new_new_n768_), .Y(new_new_n776_));
  INV        g0754(.A(new_new_n175_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n248_), .Y(new_new_n778_));
  OAI210     g0756(.A0(new_new_n715_), .A1(new_new_n468_), .B0(new_new_n113_), .Y(new_new_n779_));
  AOI210     g0757(.A0(new_new_n779_), .A1(new_new_n778_), .B0(new_new_n777_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n473_), .B(new_new_n26_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n781_), .B(new_new_n437_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n782_), .B(i_2_), .Y(new_new_n783_));
  INV        g0761(.A(new_new_n783_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n433_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n785_), .A1(new_new_n784_), .B0(new_new_n780_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n195_), .B(new_new_n128_), .Y(new_new_n787_));
  OAI210     g0765(.A0(new_new_n787_), .A1(new_new_n770_), .B0(i_2_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n176_), .Y(new_new_n789_));
  NO3        g0767(.A(new_new_n638_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n789_), .A1(new_new_n88_), .B0(new_new_n790_), .Y(new_new_n791_));
  AOI210     g0769(.A0(new_new_n791_), .A1(new_new_n788_), .B0(new_new_n198_), .Y(new_new_n792_));
  OA210      g0770(.A0(new_new_n639_), .A1(new_new_n129_), .B0(i_13_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n205_), .B(new_new_n208_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n154_), .B(new_new_n614_), .Y(new_new_n795_));
  AOI210     g0773(.A0(new_new_n795_), .A1(new_new_n794_), .B0(new_new_n385_), .Y(new_new_n796_));
  AOI210     g0774(.A0(new_new_n213_), .A1(new_new_n151_), .B0(new_new_n540_), .Y(new_new_n797_));
  NA2        g0775(.A(new_new_n797_), .B(new_new_n437_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n307_), .Y(new_new_n800_));
  NA4        g0778(.A(new_new_n800_), .B(new_new_n311_), .C(new_new_n127_), .D(new_new_n43_), .Y(new_new_n801_));
  OAI210     g0779(.A0(new_new_n801_), .A1(new_new_n799_), .B0(new_new_n798_), .Y(new_new_n802_));
  NO4        g0780(.A(new_new_n802_), .B(new_new_n796_), .C(new_new_n793_), .D(new_new_n792_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n597_), .B(new_new_n28_), .Y(new_new_n804_));
  NA2        g0782(.A(new_new_n769_), .B(new_new_n279_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n805_), .B(new_new_n804_), .Y(new_new_n806_));
  NO2        g0784(.A(new_new_n63_), .B(i_12_), .Y(new_new_n807_));
  NO2        g0785(.A(new_new_n807_), .B(new_new_n129_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n808_), .B(new_new_n614_), .Y(new_new_n809_));
  AOI220     g0787(.A0(new_new_n809_), .A1(new_new_n36_), .B0(new_new_n806_), .B1(new_new_n47_), .Y(new_new_n810_));
  NA4        g0788(.A(new_new_n810_), .B(new_new_n803_), .C(new_new_n786_), .D(new_new_n776_), .Y(mai6));
  NO3        g0789(.A(new_new_n259_), .B(new_new_n313_), .C(i_1_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n190_), .B(new_new_n142_), .Y(new_new_n813_));
  OAI210     g0791(.A0(new_new_n813_), .A1(new_new_n812_), .B0(new_new_n757_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n223_), .B(new_new_n507_), .Y(new_new_n815_));
  NO2        g0793(.A(i_11_), .B(i_9_), .Y(new_new_n816_));
  INV        g0794(.A(new_new_n336_), .Y(new_new_n817_));
  AO210      g0795(.A0(new_new_n817_), .A1(new_new_n814_), .B0(i_12_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n386_), .B(new_new_n343_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n601_), .B(new_new_n64_), .Y(new_new_n820_));
  NA2        g0798(.A(new_new_n706_), .B(new_new_n72_), .Y(new_new_n821_));
  NA3        g0799(.A(new_new_n821_), .B(new_new_n820_), .C(new_new_n819_), .Y(new_new_n822_));
  INV        g0800(.A(new_new_n202_), .Y(new_new_n823_));
  AOI220     g0801(.A0(new_new_n823_), .A1(new_new_n816_), .B0(new_new_n822_), .B1(new_new_n74_), .Y(new_new_n824_));
  INV        g0802(.A(new_new_n335_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n76_), .B(new_new_n134_), .Y(new_new_n826_));
  INV        g0804(.A(new_new_n127_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n827_), .B(new_new_n47_), .Y(new_new_n828_));
  AOI210     g0806(.A0(new_new_n828_), .A1(new_new_n826_), .B0(new_new_n825_), .Y(new_new_n829_));
  NO2        g0807(.A(new_new_n255_), .B(i_9_), .Y(new_new_n830_));
  NA2        g0808(.A(new_new_n830_), .B(new_new_n807_), .Y(new_new_n831_));
  AOI210     g0809(.A0(new_new_n831_), .A1(new_new_n538_), .B0(new_new_n190_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n32_), .B(i_11_), .Y(new_new_n833_));
  NA3        g0811(.A(new_new_n833_), .B(new_new_n492_), .C(new_new_n403_), .Y(new_new_n834_));
  NAi32      g0812(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n835_));
  NO2        g0813(.A(new_new_n742_), .B(new_new_n835_), .Y(new_new_n836_));
  OAI210     g0814(.A0(new_new_n705_), .A1(new_new_n587_), .B0(new_new_n586_), .Y(new_new_n837_));
  NAi31      g0815(.An(new_new_n836_), .B(new_new_n837_), .C(new_new_n834_), .Y(new_new_n838_));
  OR3        g0816(.A(new_new_n838_), .B(new_new_n832_), .C(new_new_n829_), .Y(new_new_n839_));
  NO2        g0817(.A(new_new_n720_), .B(i_2_), .Y(new_new_n840_));
  NA2        g0818(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n841_), .B(new_new_n425_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n842_), .B(new_new_n840_), .Y(new_new_n843_));
  AO220      g0821(.A0(new_new_n371_), .A1(new_new_n361_), .B0(new_new_n409_), .B1(new_new_n614_), .Y(new_new_n844_));
  NA3        g0822(.A(new_new_n844_), .B(new_new_n260_), .C(i_7_), .Y(new_new_n845_));
  OR2        g0823(.A(new_new_n639_), .B(new_new_n468_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n846_), .B(new_new_n150_), .C(new_new_n70_), .Y(new_new_n847_));
  AO210      g0825(.A0(new_new_n514_), .A1(new_new_n773_), .B0(new_new_n36_), .Y(new_new_n848_));
  NA4        g0826(.A(new_new_n848_), .B(new_new_n847_), .C(new_new_n845_), .D(new_new_n843_), .Y(new_new_n849_));
  NO2        g0827(.A(i_6_), .B(i_11_), .Y(new_new_n850_));
  AOI220     g0828(.A0(new_new_n850_), .A1(new_new_n586_), .B0(new_new_n815_), .B1(new_new_n736_), .Y(new_new_n851_));
  NA3        g0829(.A(new_new_n385_), .B(new_new_n241_), .C(new_new_n150_), .Y(new_new_n852_));
  NA2        g0830(.A(new_new_n409_), .B(new_new_n71_), .Y(new_new_n853_));
  NA4        g0831(.A(new_new_n853_), .B(new_new_n852_), .C(new_new_n851_), .D(new_new_n622_), .Y(new_new_n854_));
  AN2        g0832(.A(new_new_n540_), .B(new_new_n47_), .Y(new_new_n855_));
  NA3        g0833(.A(new_new_n855_), .B(new_new_n503_), .C(new_new_n222_), .Y(new_new_n856_));
  AOI210     g0834(.A0(new_new_n468_), .A1(new_new_n466_), .B0(new_new_n585_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n630_), .B(new_new_n104_), .Y(new_new_n858_));
  OAI210     g0836(.A0(new_new_n858_), .A1(new_new_n114_), .B0(new_new_n423_), .Y(new_new_n859_));
  INV        g0837(.A(new_new_n605_), .Y(new_new_n860_));
  NA3        g0838(.A(new_new_n860_), .B(new_new_n335_), .C(i_7_), .Y(new_new_n861_));
  NA4        g0839(.A(new_new_n861_), .B(new_new_n859_), .C(new_new_n857_), .D(new_new_n856_), .Y(new_new_n862_));
  NO4        g0840(.A(new_new_n862_), .B(new_new_n854_), .C(new_new_n849_), .D(new_new_n839_), .Y(new_new_n863_));
  NA4        g0841(.A(new_new_n863_), .B(new_new_n824_), .C(new_new_n818_), .D(new_new_n393_), .Y(mai3));
  NA2        g0842(.A(i_12_), .B(i_10_), .Y(new_new_n865_));
  NA2        g0843(.A(i_6_), .B(i_7_), .Y(new_new_n866_));
  NO2        g0844(.A(new_new_n866_), .B(i_0_), .Y(new_new_n867_));
  NO2        g0845(.A(i_11_), .B(new_new_n239_), .Y(new_new_n868_));
  OAI210     g0846(.A0(new_new_n867_), .A1(new_new_n295_), .B0(new_new_n868_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n869_), .B(new_new_n198_), .Y(new_new_n870_));
  NO3        g0848(.A(new_new_n469_), .B(new_new_n91_), .C(new_new_n45_), .Y(new_new_n871_));
  OA210      g0849(.A0(new_new_n871_), .A1(new_new_n870_), .B0(new_new_n178_), .Y(new_new_n872_));
  NA3        g0850(.A(new_new_n852_), .B(new_new_n622_), .C(new_new_n384_), .Y(new_new_n873_));
  NA2        g0851(.A(new_new_n873_), .B(new_new_n40_), .Y(new_new_n874_));
  NOi21      g0852(.An(new_new_n98_), .B(new_new_n782_), .Y(new_new_n875_));
  NO3        g0853(.A(new_new_n647_), .B(new_new_n473_), .C(new_new_n134_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n426_), .B(new_new_n46_), .Y(new_new_n877_));
  AN2        g0855(.A(new_new_n471_), .B(new_new_n56_), .Y(new_new_n878_));
  NO3        g0856(.A(new_new_n878_), .B(new_new_n876_), .C(new_new_n875_), .Y(new_new_n879_));
  AOI210     g0857(.A0(new_new_n879_), .A1(new_new_n874_), .B0(new_new_n49_), .Y(new_new_n880_));
  NO4        g0858(.A(new_new_n389_), .B(new_new_n396_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n190_), .B(new_new_n595_), .Y(new_new_n882_));
  NOi21      g0860(.An(new_new_n882_), .B(new_new_n881_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n729_), .B(new_new_n695_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n341_), .B(new_new_n457_), .Y(new_new_n885_));
  OAI220     g0863(.A0(new_new_n885_), .A1(new_new_n884_), .B0(new_new_n883_), .B1(new_new_n64_), .Y(new_new_n886_));
  NOi21      g0864(.An(i_5_), .B(i_9_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n887_), .B(new_new_n465_), .Y(new_new_n888_));
  BUFFER     g0866(.A(new_new_n273_), .Y(new_new_n889_));
  AOI210     g0867(.A0(new_new_n889_), .A1(new_new_n494_), .B0(new_new_n710_), .Y(new_new_n890_));
  NO3        g0868(.A(new_new_n429_), .B(new_new_n273_), .C(new_new_n74_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n179_), .B(new_new_n151_), .Y(new_new_n892_));
  AOI210     g0870(.A0(new_new_n892_), .A1(new_new_n247_), .B0(new_new_n891_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n185_), .B0(new_new_n890_), .B1(new_new_n888_), .Y(new_new_n894_));
  NO4        g0872(.A(new_new_n894_), .B(new_new_n886_), .C(new_new_n880_), .D(new_new_n872_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n190_), .B(new_new_n24_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n318_), .B(new_new_n132_), .Y(new_new_n897_));
  NO2        g0875(.A(new_new_n897_), .B(new_new_n415_), .Y(new_new_n898_));
  INV        g0876(.A(new_new_n898_), .Y(new_new_n899_));
  NO2        g0877(.A(new_new_n403_), .B(new_new_n299_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n900_), .B(new_new_n732_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n596_), .B(i_0_), .Y(new_new_n902_));
  NO4        g0880(.A(new_new_n604_), .B(new_new_n220_), .C(new_new_n433_), .D(new_new_n425_), .Y(new_new_n903_));
  NA2        g0881(.A(new_new_n903_), .B(i_11_), .Y(new_new_n904_));
  AN2        g0882(.A(new_new_n98_), .B(new_new_n246_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n769_), .B(new_new_n336_), .Y(new_new_n906_));
  AOI210     g0884(.A0(new_new_n503_), .A1(new_new_n88_), .B0(new_new_n59_), .Y(new_new_n907_));
  OAI220     g0885(.A0(new_new_n907_), .A1(new_new_n906_), .B0(new_new_n678_), .B1(new_new_n562_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n257_), .B(new_new_n156_), .Y(new_new_n909_));
  NA2        g0887(.A(i_0_), .B(i_10_), .Y(new_new_n910_));
  OAI210     g0888(.A0(new_new_n910_), .A1(new_new_n87_), .B0(new_new_n565_), .Y(new_new_n911_));
  NO4        g0889(.A(new_new_n117_), .B(new_new_n59_), .C(new_new_n688_), .D(i_5_), .Y(new_new_n912_));
  AO220      g0890(.A0(new_new_n912_), .A1(new_new_n911_), .B0(new_new_n909_), .B1(i_6_), .Y(new_new_n913_));
  AOI220     g0891(.A0(new_new_n341_), .A1(new_new_n100_), .B0(new_new_n190_), .B1(new_new_n85_), .Y(new_new_n914_));
  NA2        g0892(.A(new_new_n590_), .B(i_4_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n193_), .B(new_new_n208_), .Y(new_new_n916_));
  OAI220     g0894(.A0(new_new_n916_), .A1(new_new_n906_), .B0(new_new_n915_), .B1(new_new_n914_), .Y(new_new_n917_));
  NO4        g0895(.A(new_new_n917_), .B(new_new_n913_), .C(new_new_n908_), .D(new_new_n905_), .Y(new_new_n918_));
  NA4        g0896(.A(new_new_n918_), .B(new_new_n904_), .C(new_new_n901_), .D(new_new_n899_), .Y(new_new_n919_));
  NA2        g0897(.A(i_11_), .B(i_9_), .Y(new_new_n920_));
  NO2        g0898(.A(new_new_n49_), .B(i_7_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n408_), .B(new_new_n183_), .Y(new_new_n922_));
  NA2        g0900(.A(new_new_n922_), .B(new_new_n163_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n920_), .B(new_new_n74_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n179_), .B(i_0_), .Y(new_new_n925_));
  INV        g0903(.A(new_new_n925_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n492_), .B(new_new_n233_), .Y(new_new_n927_));
  AOI210     g0905(.A0(new_new_n383_), .A1(new_new_n42_), .B0(new_new_n422_), .Y(new_new_n928_));
  OAI220     g0906(.A0(new_new_n928_), .A1(new_new_n888_), .B0(new_new_n927_), .B1(new_new_n926_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n929_), .B(new_new_n923_), .Y(new_new_n930_));
  NA2        g0908(.A(new_new_n677_), .B(new_new_n124_), .Y(new_new_n931_));
  NO2        g0909(.A(i_6_), .B(new_new_n931_), .Y(new_new_n932_));
  AOI210     g0910(.A0(new_new_n467_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n933_));
  NA2        g0911(.A(new_new_n175_), .B(new_new_n105_), .Y(new_new_n934_));
  NOi32      g0912(.An(new_new_n933_), .Bn(new_new_n193_), .C(new_new_n934_), .Y(new_new_n935_));
  NA2        g0913(.A(new_new_n623_), .B(new_new_n336_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n936_), .B(new_new_n877_), .Y(new_new_n937_));
  NO3        g0915(.A(new_new_n937_), .B(new_new_n935_), .C(new_new_n932_), .Y(new_new_n938_));
  NOi21      g0916(.An(i_7_), .B(i_5_), .Y(new_new_n939_));
  OR2        g0917(.A(new_new_n934_), .B(new_new_n538_), .Y(new_new_n940_));
  NO3        g0918(.A(new_new_n418_), .B(new_new_n372_), .C(new_new_n370_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n267_), .B(new_new_n325_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n748_), .B(new_new_n262_), .Y(new_new_n943_));
  AOI210     g0921(.A0(new_new_n943_), .A1(new_new_n942_), .B0(new_new_n941_), .Y(new_new_n944_));
  NA4        g0922(.A(new_new_n944_), .B(new_new_n940_), .C(new_new_n938_), .D(new_new_n930_), .Y(new_new_n945_));
  NO2        g0923(.A(new_new_n896_), .B(new_new_n242_), .Y(new_new_n946_));
  AN2        g0924(.A(new_new_n340_), .B(new_new_n336_), .Y(new_new_n947_));
  AN2        g0925(.A(new_new_n947_), .B(new_new_n892_), .Y(new_new_n948_));
  OAI210     g0926(.A0(new_new_n948_), .A1(new_new_n946_), .B0(i_10_), .Y(new_new_n949_));
  NO2        g0927(.A(new_new_n865_), .B(new_new_n324_), .Y(new_new_n950_));
  OA210      g0928(.A0(new_new_n492_), .A1(new_new_n226_), .B0(new_new_n491_), .Y(new_new_n951_));
  NA2        g0929(.A(new_new_n950_), .B(new_new_n924_), .Y(new_new_n952_));
  NO2        g0930(.A(new_new_n260_), .B(new_new_n47_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n924_), .B(new_new_n311_), .Y(new_new_n954_));
  OAI210     g0932(.A0(new_new_n953_), .A1(new_new_n192_), .B0(new_new_n954_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n955_), .B(new_new_n492_), .Y(new_new_n956_));
  NA2        g0934(.A(new_new_n94_), .B(new_new_n45_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n76_), .B(new_new_n771_), .Y(new_new_n958_));
  NA2        g0936(.A(new_new_n958_), .B(new_new_n957_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n959_), .B(new_new_n48_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n722_), .B(new_new_n569_), .Y(new_new_n961_));
  NAi21      g0939(.An(i_9_), .B(i_5_), .Y(new_new_n962_));
  NO2        g0940(.A(new_new_n962_), .B(new_new_n418_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n617_), .B(new_new_n107_), .Y(new_new_n964_));
  AOI220     g0942(.A0(new_new_n964_), .A1(i_0_), .B0(new_new_n963_), .B1(new_new_n639_), .Y(new_new_n965_));
  OAI220     g0943(.A0(new_new_n965_), .A1(new_new_n87_), .B0(new_new_n961_), .B1(new_new_n176_), .Y(new_new_n966_));
  NO3        g0944(.A(new_new_n966_), .B(new_new_n960_), .C(new_new_n543_), .Y(new_new_n967_));
  NA4        g0945(.A(new_new_n967_), .B(new_new_n956_), .C(new_new_n952_), .D(new_new_n949_), .Y(new_new_n968_));
  NO3        g0946(.A(new_new_n968_), .B(new_new_n945_), .C(new_new_n919_), .Y(new_new_n969_));
  NO2        g0947(.A(i_0_), .B(new_new_n748_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n910_), .B(new_new_n971_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n973_));
  AO220      g0951(.A0(new_new_n973_), .A1(new_new_n972_), .B0(new_new_n970_), .B1(new_new_n178_), .Y(new_new_n974_));
  AOI210     g0952(.A0(new_new_n820_), .A1(new_new_n708_), .B0(new_new_n934_), .Y(new_new_n975_));
  AOI210     g0953(.A0(new_new_n974_), .A1(new_new_n358_), .B0(new_new_n975_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n757_), .B(new_new_n149_), .Y(new_new_n977_));
  INV        g0955(.A(new_new_n977_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n978_), .B(new_new_n695_), .C(new_new_n74_), .Y(new_new_n979_));
  NO2        g0957(.A(new_new_n837_), .B(new_new_n418_), .Y(new_new_n980_));
  NA3        g0958(.A(new_new_n867_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n868_), .B(i_9_), .Y(new_new_n982_));
  AOI210     g0960(.A0(new_new_n981_), .A1(new_new_n519_), .B0(new_new_n982_), .Y(new_new_n983_));
  OAI210     g0961(.A0(new_new_n247_), .A1(i_9_), .B0(new_new_n232_), .Y(new_new_n984_));
  AOI210     g0962(.A0(new_new_n984_), .A1(new_new_n902_), .B0(new_new_n156_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n985_), .B(new_new_n983_), .C(new_new_n980_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n986_), .B(new_new_n979_), .C(new_new_n976_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n947_), .B(new_new_n385_), .Y(new_new_n988_));
  AOI210     g0966(.A0(new_new_n306_), .A1(new_new_n165_), .B0(new_new_n988_), .Y(new_new_n989_));
  NA3        g0967(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n990_));
  NA2        g0968(.A(new_new_n921_), .B(new_new_n508_), .Y(new_new_n991_));
  AOI210     g0969(.A0(new_new_n990_), .A1(new_new_n165_), .B0(new_new_n991_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n992_), .B(new_new_n989_), .Y(new_new_n993_));
  NO3        g0971(.A(new_new_n910_), .B(new_new_n887_), .C(new_new_n195_), .Y(new_new_n994_));
  AOI220     g0972(.A0(new_new_n994_), .A1(i_11_), .B0(new_new_n591_), .B1(new_new_n76_), .Y(new_new_n995_));
  NO3        g0973(.A(new_new_n214_), .B(new_new_n396_), .C(i_0_), .Y(new_new_n996_));
  OAI210     g0974(.A0(new_new_n996_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n997_));
  INV        g0975(.A(new_new_n222_), .Y(new_new_n998_));
  OAI220     g0976(.A0(new_new_n555_), .A1(new_new_n142_), .B0(new_new_n661_), .B1(new_new_n634_), .Y(new_new_n999_));
  NA3        g0977(.A(new_new_n999_), .B(new_new_n410_), .C(new_new_n998_), .Y(new_new_n1000_));
  NA4        g0978(.A(new_new_n1000_), .B(new_new_n997_), .C(new_new_n995_), .D(new_new_n993_), .Y(new_new_n1001_));
  INV        g0979(.A(new_new_n111_), .Y(new_new_n1002_));
  AOI220     g0980(.A0(new_new_n939_), .A1(new_new_n508_), .B0(new_new_n867_), .B1(new_new_n166_), .Y(new_new_n1003_));
  NA2        g0981(.A(new_new_n361_), .B(new_new_n180_), .Y(new_new_n1004_));
  OA220      g0982(.A0(new_new_n1004_), .A1(new_new_n1003_), .B0(new_new_n1002_), .B1(i_5_), .Y(new_new_n1005_));
  AOI210     g0983(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n1006_));
  NA2        g0984(.A(new_new_n1006_), .B(new_new_n951_), .Y(new_new_n1007_));
  NA3        g0985(.A(new_new_n631_), .B(new_new_n190_), .C(new_new_n85_), .Y(new_new_n1008_));
  INV        g0986(.A(new_new_n1008_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n877_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1010_));
  NA2        g0988(.A(new_new_n513_), .B(new_new_n506_), .Y(new_new_n1011_));
  NO3        g0989(.A(new_new_n1011_), .B(new_new_n1010_), .C(new_new_n1009_), .Y(new_new_n1012_));
  NA3        g0990(.A(new_new_n403_), .B(new_new_n175_), .C(new_new_n174_), .Y(new_new_n1013_));
  NA3        g0991(.A(new_new_n403_), .B(new_new_n342_), .C(new_new_n224_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n1014_), .Y(new_new_n1015_));
  NOi31      g0993(.An(new_new_n402_), .B(new_new_n971_), .C(new_new_n242_), .Y(new_new_n1016_));
  NO3        g0994(.A(new_new_n920_), .B(new_new_n222_), .C(new_new_n195_), .Y(new_new_n1017_));
  NO4        g0995(.A(new_new_n1017_), .B(new_new_n1016_), .C(new_new_n1015_), .D(new_new_n1080_), .Y(new_new_n1018_));
  NA4        g0996(.A(new_new_n1018_), .B(new_new_n1012_), .C(new_new_n1007_), .D(new_new_n1005_), .Y(new_new_n1019_));
  INV        g0997(.A(new_new_n633_), .Y(new_new_n1020_));
  NO3        g0998(.A(new_new_n1020_), .B(new_new_n581_), .C(new_new_n355_), .Y(new_new_n1021_));
  NO2        g0999(.A(new_new_n87_), .B(i_5_), .Y(new_new_n1022_));
  NA3        g1000(.A(new_new_n868_), .B(new_new_n112_), .C(new_new_n127_), .Y(new_new_n1023_));
  INV        g1001(.A(new_new_n1023_), .Y(new_new_n1024_));
  AOI210     g1002(.A0(new_new_n1024_), .A1(new_new_n1022_), .B0(new_new_n1021_), .Y(new_new_n1025_));
  NAi21      g1003(.An(new_new_n244_), .B(new_new_n245_), .Y(new_new_n1026_));
  NO4        g1004(.A(new_new_n242_), .B(new_new_n214_), .C(i_0_), .D(i_12_), .Y(new_new_n1027_));
  NA2        g1005(.A(new_new_n1027_), .B(new_new_n1026_), .Y(new_new_n1028_));
  AN2        g1006(.A(new_new_n910_), .B(new_new_n156_), .Y(new_new_n1029_));
  NO4        g1007(.A(new_new_n1029_), .B(i_12_), .C(new_new_n665_), .D(new_new_n134_), .Y(new_new_n1030_));
  NA2        g1008(.A(new_new_n1030_), .B(new_new_n222_), .Y(new_new_n1031_));
  NA3        g1009(.A(new_new_n100_), .B(new_new_n595_), .C(i_11_), .Y(new_new_n1032_));
  NO2        g1010(.A(new_new_n1032_), .B(new_new_n158_), .Y(new_new_n1033_));
  NA2        g1011(.A(new_new_n939_), .B(new_new_n490_), .Y(new_new_n1034_));
  NO2        g1012(.A(new_new_n1034_), .B(new_new_n696_), .Y(new_new_n1035_));
  AOI210     g1013(.A0(new_new_n1035_), .A1(new_new_n925_), .B0(new_new_n1033_), .Y(new_new_n1036_));
  NA4        g1014(.A(new_new_n1036_), .B(new_new_n1031_), .C(new_new_n1028_), .D(new_new_n1025_), .Y(new_new_n1037_));
  NO4        g1015(.A(new_new_n1037_), .B(new_new_n1019_), .C(new_new_n1001_), .D(new_new_n987_), .Y(new_new_n1038_));
  OAI210     g1016(.A0(new_new_n840_), .A1(new_new_n833_), .B0(new_new_n37_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n933_), .B(new_new_n380_), .C(i_5_), .Y(new_new_n1040_));
  NA3        g1018(.A(new_new_n1040_), .B(new_new_n1039_), .C(new_new_n629_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n1041_), .B(new_new_n211_), .Y(new_new_n1042_));
  BUFFER     g1020(.A(new_new_n381_), .Y(new_new_n1043_));
  NA2        g1021(.A(new_new_n191_), .B(new_new_n193_), .Y(new_new_n1044_));
  AO210      g1022(.A0(new_new_n1043_), .A1(new_new_n33_), .B0(new_new_n1044_), .Y(new_new_n1045_));
  OAI210     g1023(.A0(new_new_n633_), .A1(new_new_n631_), .B0(new_new_n324_), .Y(new_new_n1046_));
  NAi31      g1024(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1047_));
  AOI210     g1025(.A0(new_new_n120_), .A1(new_new_n71_), .B0(new_new_n1047_), .Y(new_new_n1048_));
  NO2        g1026(.A(new_new_n1048_), .B(new_new_n662_), .Y(new_new_n1049_));
  NA3        g1027(.A(new_new_n1049_), .B(new_new_n1046_), .C(new_new_n1045_), .Y(new_new_n1050_));
  NO2        g1028(.A(new_new_n481_), .B(new_new_n273_), .Y(new_new_n1051_));
  NO4        g1029(.A(new_new_n235_), .B(new_new_n148_), .C(new_new_n699_), .D(new_new_n37_), .Y(new_new_n1052_));
  NO3        g1030(.A(new_new_n1052_), .B(new_new_n1051_), .C(new_new_n903_), .Y(new_new_n1053_));
  OAI210     g1031(.A0(new_new_n1032_), .A1(new_new_n151_), .B0(new_new_n1053_), .Y(new_new_n1054_));
  AOI210     g1032(.A0(new_new_n1050_), .A1(new_new_n49_), .B0(new_new_n1054_), .Y(new_new_n1055_));
  AOI210     g1033(.A0(new_new_n1055_), .A1(new_new_n1042_), .B0(new_new_n74_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n588_), .B(new_new_n392_), .Y(new_new_n1057_));
  NO2        g1035(.A(new_new_n1057_), .B(new_new_n777_), .Y(new_new_n1058_));
  NA2        g1036(.A(new_new_n267_), .B(new_new_n58_), .Y(new_new_n1059_));
  AOI220     g1037(.A0(new_new_n1059_), .A1(new_new_n77_), .B0(new_new_n356_), .B1(new_new_n259_), .Y(new_new_n1060_));
  NO2        g1038(.A(new_new_n1060_), .B(new_new_n239_), .Y(new_new_n1061_));
  NA3        g1039(.A(new_new_n98_), .B(new_new_n313_), .C(new_new_n31_), .Y(new_new_n1062_));
  INV        g1040(.A(new_new_n1062_), .Y(new_new_n1063_));
  NO2        g1041(.A(new_new_n1063_), .B(new_new_n1061_), .Y(new_new_n1064_));
  NA2        g1042(.A(new_new_n161_), .B(new_new_n88_), .Y(new_new_n1065_));
  NO2        g1043(.A(new_new_n1065_), .B(i_11_), .Y(new_new_n1066_));
  NO4        g1044(.A(new_new_n962_), .B(new_new_n496_), .C(new_new_n256_), .D(new_new_n255_), .Y(new_new_n1067_));
  NO2        g1045(.A(new_new_n1067_), .B(new_new_n585_), .Y(new_new_n1068_));
  INV        g1046(.A(new_new_n373_), .Y(new_new_n1069_));
  AOI210     g1047(.A0(new_new_n1069_), .A1(new_new_n1068_), .B0(new_new_n41_), .Y(new_new_n1070_));
  NO2        g1048(.A(new_new_n1070_), .B(new_new_n1066_), .Y(new_new_n1071_));
  OAI210     g1049(.A0(new_new_n1064_), .A1(i_4_), .B0(new_new_n1071_), .Y(new_new_n1072_));
  NO3        g1050(.A(new_new_n1072_), .B(new_new_n1058_), .C(new_new_n1056_), .Y(new_new_n1073_));
  NA4        g1051(.A(new_new_n1073_), .B(new_new_n1038_), .C(new_new_n969_), .D(new_new_n895_), .Y(mai4));
  INV        g1052(.A(new_new_n721_), .Y(new_new_n1077_));
  INV        g1053(.A(i_2_), .Y(new_new_n1078_));
  INV        g1054(.A(new_new_n249_), .Y(new_new_n1079_));
  INV        g1055(.A(new_new_n1013_), .Y(new_new_n1080_));
endmodule


