library verilog;
use verilog.vl_types.all;
entity decodificador2x4_vlg_vec_tst is
end decodificador2x4_vlg_vec_tst;
