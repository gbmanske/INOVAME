library verilog;
use verilog.vl_types.all;
entity divisordefreq2_vlg_vec_tst is
end divisordefreq2_vlg_vec_tst;
