// Benchmark "top" written by ABC on Thu Jun 20 14:59:19 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n132_, new_new_n133_, new_new_n134_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n697_, new_new_n698_, new_new_n699_,
    new_new_n700_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n712_, new_new_n713_, new_new_n714_, new_new_n715_,
    new_new_n716_, new_new_n717_, new_new_n718_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n925_, new_new_n926_, new_new_n927_,
    new_new_n928_, new_new_n929_, new_new_n930_, new_new_n931_,
    new_new_n932_, new_new_n933_, new_new_n934_, new_new_n935_,
    new_new_n936_, new_new_n937_, new_new_n938_, new_new_n939_,
    new_new_n940_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NO2        g028(.A(new_new_n47_), .B(new_new_n46_), .Y(new_new_n51_));
  NA2        g029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n51_), .B(new_new_n45_), .Y(new_new_n54_));
  NA3        g032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  OAI210     g035(.A0(new_new_n57_), .A1(new_new_n56_), .B0(new_new_n55_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi31      g043(.An(new_new_n65_), .B(new_new_n63_), .C(new_new_n59_), .Y(new_new_n66_));
  NA2        g044(.A(new_new_n50_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  INV        g053(.A(new_new_n75_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  INV        g059(.A(i_6_), .Y(new_new_n82_));
  OR4        g060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n83_));
  INV        g061(.A(new_new_n83_), .Y(new_new_n84_));
  NO2        g062(.A(i_2_), .B(i_7_), .Y(new_new_n85_));
  NO2        g063(.A(new_new_n84_), .B(new_new_n85_), .Y(new_new_n86_));
  NA2        g064(.A(i_1_), .B(new_new_n86_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_10_), .Y(new_new_n88_));
  NA2        g066(.A(i_6_), .B(i_9_), .Y(new_new_n89_));
  AOI210     g067(.A0(new_new_n89_), .A1(new_new_n88_), .B0(new_new_n61_), .Y(new_new_n90_));
  NA2        g068(.A(i_2_), .B(i_6_), .Y(new_new_n91_));
  INV        g069(.A(new_new_n90_), .Y(new_new_n92_));
  AOI210     g070(.A0(new_new_n92_), .A1(new_new_n87_), .B0(new_new_n78_), .Y(new_new_n93_));
  AN3        g071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NO2        g073(.A(i_5_), .B(i_8_), .Y(new_new_n96_));
  NOi21      g074(.An(new_new_n96_), .B(new_new_n95_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n97_), .B(new_new_n60_), .Y(new_new_n98_));
  INV        g076(.A(i_7_), .Y(new_new_n99_));
  NA2        g077(.A(new_new_n46_), .B(new_new_n99_), .Y(new_new_n100_));
  NO2        g078(.A(i_0_), .B(i_5_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(new_new_n82_), .Y(new_new_n102_));
  NA2        g080(.A(i_12_), .B(i_3_), .Y(new_new_n103_));
  INV        g081(.A(new_new_n103_), .Y(new_new_n104_));
  NA3        g082(.A(new_new_n104_), .B(new_new_n102_), .C(new_new_n100_), .Y(new_new_n105_));
  NAi21      g083(.An(i_7_), .B(i_11_), .Y(new_new_n106_));
  AN2        g084(.A(i_2_), .B(i_10_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n107_), .B(i_7_), .Y(new_new_n108_));
  OR2        g086(.A(new_new_n78_), .B(new_new_n56_), .Y(new_new_n109_));
  NO2        g087(.A(i_8_), .B(new_new_n99_), .Y(new_new_n110_));
  NO3        g088(.A(new_new_n110_), .B(new_new_n109_), .C(new_new_n108_), .Y(new_new_n111_));
  NA2        g089(.A(i_12_), .B(i_7_), .Y(new_new_n112_));
  NA2        g090(.A(i_11_), .B(i_12_), .Y(new_new_n113_));
  INV        g091(.A(new_new_n113_), .Y(new_new_n114_));
  NO2        g092(.A(new_new_n114_), .B(new_new_n111_), .Y(new_new_n115_));
  NA3        g093(.A(new_new_n115_), .B(new_new_n105_), .C(new_new_n98_), .Y(new_new_n116_));
  NOi21      g094(.An(i_1_), .B(i_5_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(i_11_), .Y(new_new_n118_));
  NA2        g096(.A(i_7_), .B(new_new_n25_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_10_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(new_new_n46_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n89_), .B(new_new_n88_), .Y(new_new_n122_));
  NAi21      g100(.An(i_3_), .B(i_8_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n60_), .Y(new_new_n124_));
  NOi31      g102(.An(new_new_n124_), .B(new_new_n122_), .C(new_new_n121_), .Y(new_new_n125_));
  NO2        g103(.A(i_1_), .B(new_new_n82_), .Y(new_new_n126_));
  NO2        g104(.A(i_6_), .B(i_5_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(i_3_), .Y(new_new_n128_));
  NO2        g106(.A(new_new_n125_), .B(new_new_n118_), .Y(new_new_n129_));
  NO3        g107(.A(new_new_n129_), .B(new_new_n116_), .C(new_new_n93_), .Y(new_new_n130_));
  NA3        g108(.A(new_new_n130_), .B(new_new_n77_), .C(new_new_n54_), .Y(mai2));
  NO2        g109(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n132_));
  NA2        g110(.A(i_6_), .B(new_new_n25_), .Y(new_new_n133_));
  NA2        g111(.A(new_new_n133_), .B(new_new_n132_), .Y(new_new_n134_));
  NA4        g112(.A(new_new_n134_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(mai0));
  AN2        g113(.A(i_8_), .B(i_7_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_6_), .Y(new_new_n137_));
  NO2        g115(.A(i_12_), .B(i_13_), .Y(new_new_n138_));
  NAi21      g116(.An(i_5_), .B(i_11_), .Y(new_new_n139_));
  NOi21      g117(.An(new_new_n138_), .B(new_new_n139_), .Y(new_new_n140_));
  NO2        g118(.A(i_0_), .B(i_1_), .Y(new_new_n141_));
  NA2        g119(.A(i_2_), .B(i_3_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n142_), .B(i_4_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n140_), .Y(new_new_n144_));
  AN2        g122(.A(new_new_n138_), .B(new_new_n80_), .Y(new_new_n145_));
  NO2        g123(.A(new_new_n145_), .B(new_new_n27_), .Y(new_new_n146_));
  NA2        g124(.A(i_1_), .B(i_5_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n71_), .B(new_new_n46_), .Y(new_new_n148_));
  NA2        g126(.A(new_new_n148_), .B(new_new_n36_), .Y(new_new_n149_));
  NO3        g127(.A(new_new_n149_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n150_));
  OR2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NO3        g129(.A(new_new_n151_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n152_));
  NAi32      g130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n153_));
  NAi21      g131(.An(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  NOi21      g132(.An(i_4_), .B(i_10_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n40_), .Y(new_new_n156_));
  NO2        g134(.A(i_3_), .B(i_5_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n157_), .Y(new_new_n159_));
  OAI210     g137(.A0(new_new_n159_), .A1(new_new_n156_), .B0(new_new_n154_), .Y(new_new_n160_));
  NO2        g138(.A(new_new_n160_), .B(new_new_n150_), .Y(new_new_n161_));
  AOI210     g139(.A0(new_new_n161_), .A1(new_new_n144_), .B0(new_new_n137_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n46_), .B(i_1_), .Y(new_new_n163_));
  NOi21      g141(.An(i_4_), .B(i_9_), .Y(new_new_n164_));
  NOi21      g142(.An(i_11_), .B(i_13_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  BUFFER     g144(.A(new_new_n166_), .Y(new_new_n167_));
  NO2        g145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NA3        g148(.A(new_new_n170_), .B(new_new_n168_), .C(new_new_n80_), .Y(new_new_n171_));
  AOI210     g149(.A0(new_new_n171_), .A1(new_new_n167_), .B0(new_new_n163_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n71_), .B(new_new_n61_), .Y(new_new_n173_));
  INV        g151(.A(new_new_n173_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n36_), .B(i_5_), .Y(new_new_n175_));
  NAi31      g153(.An(new_new_n175_), .B(new_new_n145_), .C(i_11_), .Y(new_new_n176_));
  NA2        g154(.A(i_3_), .B(i_5_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n176_), .B(new_new_n174_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n71_), .B(i_5_), .Y(new_new_n179_));
  NO2        g157(.A(i_13_), .B(i_10_), .Y(new_new_n180_));
  NA3        g158(.A(new_new_n180_), .B(new_new_n179_), .C(new_new_n44_), .Y(new_new_n181_));
  NO2        g159(.A(i_2_), .B(i_1_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(i_3_), .Y(new_new_n183_));
  NAi21      g161(.An(i_4_), .B(i_12_), .Y(new_new_n184_));
  NO3        g162(.A(new_new_n184_), .B(new_new_n183_), .C(new_new_n181_), .Y(new_new_n185_));
  NO3        g163(.A(new_new_n185_), .B(new_new_n178_), .C(new_new_n172_), .Y(new_new_n186_));
  INV        g164(.A(i_8_), .Y(new_new_n187_));
  NA2        g165(.A(i_8_), .B(i_6_), .Y(new_new_n188_));
  NO3        g166(.A(i_3_), .B(new_new_n82_), .C(new_new_n48_), .Y(new_new_n189_));
  NA2        g167(.A(new_new_n189_), .B(new_new_n110_), .Y(new_new_n190_));
  NO3        g168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n191_));
  NA3        g169(.A(new_new_n191_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n193_));
  INV        g171(.A(new_new_n193_), .Y(new_new_n194_));
  AOI210     g172(.A0(new_new_n194_), .A1(new_new_n192_), .B0(new_new_n190_), .Y(new_new_n195_));
  NO2        g173(.A(i_3_), .B(i_8_), .Y(new_new_n196_));
  NO3        g174(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n197_));
  NO2        g175(.A(i_13_), .B(i_9_), .Y(new_new_n198_));
  NA2        g176(.A(new_new_n198_), .B(i_6_), .Y(new_new_n199_));
  NAi21      g177(.An(i_12_), .B(i_3_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n44_), .B(i_5_), .Y(new_new_n201_));
  NO3        g179(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n202_));
  INV        g180(.A(new_new_n195_), .Y(new_new_n203_));
  OAI220     g181(.A0(new_new_n203_), .A1(i_4_), .B0(new_new_n188_), .B1(new_new_n186_), .Y(new_new_n204_));
  NA3        g182(.A(i_13_), .B(new_new_n187_), .C(i_10_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n205_), .B(i_12_), .Y(new_new_n206_));
  NA2        g184(.A(i_0_), .B(i_5_), .Y(new_new_n207_));
  NA2        g185(.A(new_new_n207_), .B(new_new_n102_), .Y(new_new_n208_));
  OAI220     g186(.A0(new_new_n208_), .A1(new_new_n183_), .B0(new_new_n174_), .B1(new_new_n128_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n36_), .B(i_13_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n46_), .B(new_new_n61_), .Y(new_new_n212_));
  NA3        g190(.A(new_new_n212_), .B(new_new_n211_), .C(new_new_n210_), .Y(new_new_n213_));
  INV        g191(.A(i_13_), .Y(new_new_n214_));
  NO2        g192(.A(i_12_), .B(new_new_n214_), .Y(new_new_n215_));
  NA3        g193(.A(new_new_n215_), .B(new_new_n191_), .C(new_new_n189_), .Y(new_new_n216_));
  OAI210     g194(.A0(new_new_n213_), .A1(i_9_), .B0(new_new_n216_), .Y(new_new_n217_));
  AOI220     g195(.A0(new_new_n217_), .A1(new_new_n136_), .B0(new_new_n209_), .B1(new_new_n206_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n177_), .B(i_4_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n219_), .B(new_new_n934_), .Y(new_new_n220_));
  OR2        g198(.A(i_8_), .B(i_7_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n52_), .B(i_1_), .Y(new_new_n222_));
  NA2        g200(.A(new_new_n222_), .B(i_6_), .Y(new_new_n223_));
  INV        g201(.A(i_12_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n44_), .B(new_new_n224_), .Y(new_new_n225_));
  NO3        g203(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n226_));
  NA2        g204(.A(i_2_), .B(i_1_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n223_), .B(new_new_n220_), .Y(new_new_n228_));
  NAi21      g206(.An(i_4_), .B(i_3_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n229_), .B(new_new_n73_), .Y(new_new_n230_));
  NO2        g208(.A(i_0_), .B(i_6_), .Y(new_new_n231_));
  NOi41      g209(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  AOI210     g211(.A0(new_new_n932_), .A1(new_new_n40_), .B0(new_new_n228_), .Y(new_new_n234_));
  NO2        g212(.A(i_11_), .B(new_new_n214_), .Y(new_new_n235_));
  NOi21      g213(.An(i_1_), .B(i_6_), .Y(new_new_n236_));
  NAi21      g214(.An(i_3_), .B(i_7_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n224_), .B(i_9_), .Y(new_new_n238_));
  OR4        g216(.A(new_new_n238_), .B(new_new_n237_), .C(new_new_n236_), .D(new_new_n179_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n240_));
  NO2        g218(.A(i_12_), .B(i_3_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n71_), .B(i_5_), .Y(new_new_n242_));
  NA2        g220(.A(i_3_), .B(i_9_), .Y(new_new_n243_));
  NAi21      g221(.An(i_7_), .B(i_10_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n244_), .B(new_new_n243_), .Y(new_new_n245_));
  NA3        g223(.A(new_new_n245_), .B(new_new_n242_), .C(new_new_n62_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n246_), .B(new_new_n239_), .Y(new_new_n247_));
  NA3        g225(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n248_));
  INV        g226(.A(new_new_n137_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n224_), .B(i_13_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n250_), .B(new_new_n73_), .Y(new_new_n251_));
  AOI220     g229(.A0(new_new_n251_), .A1(new_new_n249_), .B0(new_new_n247_), .B1(new_new_n235_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n221_), .B(new_new_n37_), .Y(new_new_n253_));
  NA2        g231(.A(i_12_), .B(i_6_), .Y(new_new_n254_));
  NO3        g232(.A(i_9_), .B(new_new_n254_), .C(new_new_n48_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n229_), .B(i_2_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n235_), .B(i_9_), .Y(new_new_n257_));
  NA2        g235(.A(new_new_n148_), .B(new_new_n61_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n237_), .B(i_8_), .Y(new_new_n259_));
  NO2        g237(.A(i_6_), .B(new_new_n48_), .Y(new_new_n260_));
  NA3        g238(.A(new_new_n260_), .B(new_new_n259_), .C(i_9_), .Y(new_new_n261_));
  NA3        g239(.A(i_6_), .B(new_new_n253_), .C(new_new_n215_), .Y(new_new_n262_));
  AOI210     g240(.A0(new_new_n262_), .A1(new_new_n261_), .B0(new_new_n258_), .Y(new_new_n263_));
  INV        g241(.A(new_new_n263_), .Y(new_new_n264_));
  NA4        g242(.A(new_new_n264_), .B(new_new_n252_), .C(new_new_n234_), .D(new_new_n218_), .Y(new_new_n265_));
  NO3        g243(.A(i_12_), .B(new_new_n214_), .C(new_new_n37_), .Y(new_new_n266_));
  INV        g244(.A(new_new_n266_), .Y(new_new_n267_));
  NA2        g245(.A(i_8_), .B(new_new_n99_), .Y(new_new_n268_));
  NO3        g246(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n269_));
  AOI220     g247(.A0(new_new_n269_), .A1(new_new_n189_), .B0(i_6_), .B1(new_new_n222_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n270_), .B(new_new_n268_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n227_), .B(i_0_), .Y(new_new_n272_));
  AOI220     g250(.A0(new_new_n272_), .A1(i_8_), .B0(i_1_), .B1(new_new_n136_), .Y(new_new_n273_));
  NA2        g251(.A(new_new_n260_), .B(new_new_n26_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n274_), .B(new_new_n273_), .Y(new_new_n275_));
  NA2        g253(.A(i_0_), .B(i_1_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(i_2_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n57_), .B(i_6_), .Y(new_new_n278_));
  NA3        g256(.A(new_new_n278_), .B(new_new_n277_), .C(new_new_n157_), .Y(new_new_n279_));
  OAI210     g257(.A0(new_new_n159_), .A1(new_new_n137_), .B0(new_new_n279_), .Y(new_new_n280_));
  NO3        g258(.A(new_new_n280_), .B(new_new_n275_), .C(new_new_n271_), .Y(new_new_n281_));
  NO2        g259(.A(i_3_), .B(i_10_), .Y(new_new_n282_));
  NA3        g260(.A(new_new_n282_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n283_));
  NA2        g261(.A(i_1_), .B(new_new_n36_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(i_8_), .Y(new_new_n285_));
  NA2        g263(.A(new_new_n285_), .B(i_7_), .Y(new_new_n286_));
  AN2        g264(.A(i_3_), .B(i_10_), .Y(new_new_n287_));
  NA3        g265(.A(new_new_n287_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n288_));
  NO2        g266(.A(i_5_), .B(new_new_n37_), .Y(new_new_n289_));
  NO2        g267(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n290_));
  OR2        g268(.A(new_new_n286_), .B(new_new_n283_), .Y(new_new_n291_));
  OAI220     g269(.A0(new_new_n291_), .A1(i_6_), .B0(new_new_n281_), .B1(new_new_n267_), .Y(new_new_n292_));
  NO4        g270(.A(new_new_n292_), .B(new_new_n265_), .C(new_new_n204_), .D(new_new_n162_), .Y(new_new_n293_));
  NO3        g271(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n57_), .B(new_new_n82_), .Y(new_new_n295_));
  NA2        g273(.A(new_new_n272_), .B(new_new_n295_), .Y(new_new_n296_));
  NO3        g274(.A(i_6_), .B(new_new_n187_), .C(i_7_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n297_), .B(new_new_n191_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n298_), .B(new_new_n296_), .Y(new_new_n299_));
  NO2        g277(.A(i_2_), .B(i_3_), .Y(new_new_n300_));
  OR2        g278(.A(i_0_), .B(i_5_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n207_), .B(new_new_n301_), .Y(new_new_n302_));
  NA4        g280(.A(new_new_n302_), .B(i_6_), .C(new_new_n300_), .D(i_1_), .Y(new_new_n303_));
  NA3        g281(.A(new_new_n272_), .B(i_6_), .C(new_new_n110_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n151_), .B(new_new_n46_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n305_), .B(i_7_), .C(new_new_n157_), .Y(new_new_n306_));
  NA3        g284(.A(new_new_n306_), .B(new_new_n304_), .C(new_new_n303_), .Y(new_new_n307_));
  OAI210     g285(.A0(new_new_n307_), .A1(new_new_n299_), .B0(i_4_), .Y(new_new_n308_));
  NO2        g286(.A(i_12_), .B(i_10_), .Y(new_new_n309_));
  NOi21      g287(.An(i_5_), .B(i_0_), .Y(new_new_n310_));
  NO3        g288(.A(new_new_n284_), .B(new_new_n310_), .C(new_new_n123_), .Y(new_new_n311_));
  NA4        g289(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n82_), .D(i_8_), .Y(new_new_n312_));
  NA2        g290(.A(new_new_n311_), .B(new_new_n309_), .Y(new_new_n313_));
  NO2        g291(.A(i_6_), .B(i_8_), .Y(new_new_n314_));
  NOi21      g292(.An(i_0_), .B(i_2_), .Y(new_new_n315_));
  AN2        g293(.A(new_new_n315_), .B(new_new_n314_), .Y(new_new_n316_));
  NO2        g294(.A(i_1_), .B(i_7_), .Y(new_new_n317_));
  AO220      g295(.A0(new_new_n317_), .A1(new_new_n316_), .B0(i_7_), .B1(new_new_n222_), .Y(new_new_n318_));
  NA3        g296(.A(new_new_n318_), .B(i_4_), .C(i_5_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n319_), .B(new_new_n313_), .C(new_new_n308_), .Y(new_new_n320_));
  NO3        g298(.A(new_new_n221_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n321_));
  OAI210     g299(.A0(i_7_), .A1(new_new_n321_), .B0(i_6_), .Y(new_new_n322_));
  AOI210     g300(.A0(new_new_n99_), .A1(new_new_n322_), .B0(new_new_n302_), .Y(new_new_n323_));
  NOi21      g301(.An(new_new_n147_), .B(new_new_n102_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n324_), .B(new_new_n119_), .Y(new_new_n325_));
  OAI210     g303(.A0(new_new_n325_), .A1(new_new_n323_), .B0(i_3_), .Y(new_new_n326_));
  INV        g304(.A(new_new_n81_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n276_), .B(new_new_n79_), .Y(new_new_n328_));
  INV        g306(.A(new_new_n328_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n91_), .B(new_new_n187_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n330_), .B(new_new_n61_), .Y(new_new_n331_));
  AOI210     g309(.A0(new_new_n331_), .A1(new_new_n329_), .B0(new_new_n327_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n187_), .B(i_9_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n332_), .B(new_new_n275_), .Y(new_new_n334_));
  AOI210     g312(.A0(new_new_n334_), .A1(new_new_n326_), .B0(new_new_n156_), .Y(new_new_n335_));
  AOI210     g313(.A0(new_new_n320_), .A1(new_new_n294_), .B0(new_new_n335_), .Y(new_new_n336_));
  NOi32      g314(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n337_));
  INV        g315(.A(new_new_n337_), .Y(new_new_n338_));
  NAi21      g316(.An(i_0_), .B(i_6_), .Y(new_new_n339_));
  NAi21      g317(.An(i_1_), .B(i_5_), .Y(new_new_n340_));
  NA2        g318(.A(new_new_n340_), .B(new_new_n339_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n25_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n342_), .B(new_new_n153_), .Y(new_new_n343_));
  NAi41      g321(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n344_), .A1(new_new_n153_), .B0(new_new_n151_), .Y(new_new_n345_));
  NOi32      g323(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n346_));
  NO2        g324(.A(i_1_), .B(new_new_n99_), .Y(new_new_n347_));
  NAi21      g325(.An(i_3_), .B(i_4_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(i_9_), .Y(new_new_n349_));
  AN2        g327(.A(i_6_), .B(i_7_), .Y(new_new_n350_));
  OAI210     g328(.A0(new_new_n350_), .A1(new_new_n347_), .B0(new_new_n349_), .Y(new_new_n351_));
  NA2        g329(.A(i_2_), .B(i_7_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n348_), .B(i_10_), .Y(new_new_n353_));
  NA3        g331(.A(new_new_n353_), .B(new_new_n352_), .C(new_new_n231_), .Y(new_new_n354_));
  AOI210     g332(.A0(new_new_n354_), .A1(new_new_n351_), .B0(new_new_n179_), .Y(new_new_n355_));
  AOI210     g333(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n356_));
  OAI210     g334(.A0(new_new_n356_), .A1(new_new_n182_), .B0(new_new_n353_), .Y(new_new_n357_));
  AOI220     g335(.A0(new_new_n353_), .A1(new_new_n317_), .B0(new_new_n226_), .B1(new_new_n182_), .Y(new_new_n358_));
  AOI210     g336(.A0(new_new_n358_), .A1(new_new_n357_), .B0(i_5_), .Y(new_new_n359_));
  NO4        g337(.A(new_new_n359_), .B(new_new_n355_), .C(new_new_n345_), .D(new_new_n343_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n360_), .B(new_new_n338_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n362_));
  AN2        g340(.A(i_12_), .B(i_5_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n937_), .B(new_new_n363_), .Y(new_new_n364_));
  NO2        g342(.A(i_11_), .B(i_6_), .Y(new_new_n365_));
  NA3        g343(.A(new_new_n365_), .B(new_new_n305_), .C(new_new_n214_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n366_), .B(new_new_n364_), .Y(new_new_n367_));
  NO2        g345(.A(i_5_), .B(i_10_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n138_), .B(new_new_n45_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(new_new_n229_), .Y(new_new_n370_));
  OAI210     g348(.A0(new_new_n370_), .A1(new_new_n367_), .B0(new_new_n362_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n367_), .B(new_new_n372_), .Y(new_new_n373_));
  NO3        g351(.A(new_new_n82_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n374_));
  NO2        g352(.A(i_11_), .B(i_12_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n368_), .B(new_new_n224_), .Y(new_new_n376_));
  NA3        g354(.A(new_new_n110_), .B(i_4_), .C(i_11_), .Y(new_new_n377_));
  INV        g355(.A(new_new_n377_), .Y(new_new_n378_));
  NAi21      g356(.An(i_13_), .B(i_0_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n227_), .Y(new_new_n380_));
  NA2        g358(.A(new_new_n378_), .B(new_new_n380_), .Y(new_new_n381_));
  NA3        g359(.A(new_new_n381_), .B(new_new_n373_), .C(new_new_n371_), .Y(new_new_n382_));
  NO3        g360(.A(i_1_), .B(i_12_), .C(new_new_n82_), .Y(new_new_n383_));
  NO2        g361(.A(i_0_), .B(i_11_), .Y(new_new_n384_));
  AN2        g362(.A(i_1_), .B(i_6_), .Y(new_new_n385_));
  NOi21      g363(.An(i_2_), .B(i_12_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  INV        g365(.A(new_new_n387_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n136_), .B(i_9_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(i_4_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n388_), .B(new_new_n390_), .Y(new_new_n391_));
  NAi21      g369(.An(i_9_), .B(i_4_), .Y(new_new_n392_));
  OR2        g370(.A(i_13_), .B(i_10_), .Y(new_new_n393_));
  NO3        g371(.A(new_new_n393_), .B(new_new_n113_), .C(new_new_n392_), .Y(new_new_n394_));
  BUFFER     g372(.A(new_new_n205_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n99_), .B(new_new_n25_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n266_), .B(new_new_n396_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n260_), .B(new_new_n202_), .Y(new_new_n398_));
  OAI220     g376(.A0(new_new_n398_), .A1(new_new_n395_), .B0(new_new_n397_), .B1(new_new_n324_), .Y(new_new_n399_));
  INV        g377(.A(new_new_n399_), .Y(new_new_n400_));
  AOI210     g378(.A0(new_new_n400_), .A1(new_new_n391_), .B0(new_new_n26_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n304_), .B(new_new_n303_), .Y(new_new_n402_));
  AOI220     g380(.A0(new_new_n278_), .A1(new_new_n269_), .B0(new_new_n272_), .B1(new_new_n295_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n403_), .B(i_5_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n177_), .B(new_new_n82_), .Y(new_new_n405_));
  AOI220     g383(.A0(new_new_n405_), .A1(new_new_n277_), .B0(i_6_), .B1(new_new_n202_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n406_), .B(new_new_n268_), .Y(new_new_n407_));
  NO3        g385(.A(new_new_n407_), .B(new_new_n404_), .C(new_new_n402_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n189_), .B(new_new_n94_), .Y(new_new_n409_));
  NA3        g387(.A(new_new_n305_), .B(new_new_n157_), .C(new_new_n82_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n410_), .A1(new_new_n409_), .B0(i_8_), .Y(new_new_n411_));
  INV        g389(.A(i_10_), .Y(new_new_n412_));
  NA3        g390(.A(new_new_n242_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n278_), .B(new_new_n222_), .Y(new_new_n414_));
  OAI220     g392(.A0(new_new_n414_), .A1(new_new_n177_), .B0(new_new_n413_), .B1(new_new_n412_), .Y(new_new_n415_));
  NA3        g393(.A(new_new_n317_), .B(new_new_n316_), .C(i_5_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n297_), .B(new_new_n302_), .Y(new_new_n417_));
  OAI210     g395(.A0(new_new_n417_), .A1(new_new_n183_), .B0(new_new_n416_), .Y(new_new_n418_));
  NO3        g396(.A(new_new_n418_), .B(new_new_n415_), .C(new_new_n411_), .Y(new_new_n419_));
  AOI210     g397(.A0(new_new_n419_), .A1(new_new_n408_), .B0(new_new_n257_), .Y(new_new_n420_));
  NO4        g398(.A(new_new_n420_), .B(new_new_n401_), .C(new_new_n382_), .D(new_new_n361_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n71_), .B(i_13_), .Y(new_new_n422_));
  NO2        g400(.A(i_10_), .B(i_9_), .Y(new_new_n423_));
  NAi21      g401(.An(i_12_), .B(i_8_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n424_), .B(i_3_), .Y(new_new_n425_));
  NO3        g403(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n254_), .B(new_new_n95_), .Y(new_new_n427_));
  NA2        g405(.A(i_8_), .B(i_9_), .Y(new_new_n428_));
  NO3        g406(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n429_));
  NA3        g407(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n430_));
  OR2        g408(.A(new_new_n276_), .B(new_new_n199_), .Y(new_new_n431_));
  BUFFER     g409(.A(new_new_n279_), .Y(new_new_n432_));
  OA220      g410(.A0(new_new_n432_), .A1(new_new_n156_), .B0(new_new_n431_), .B1(new_new_n220_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n94_), .B(i_13_), .Y(new_new_n434_));
  INV        g412(.A(new_new_n362_), .Y(new_new_n435_));
  NO2        g413(.A(i_2_), .B(i_13_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n435_), .B(new_new_n434_), .Y(new_new_n437_));
  NO3        g415(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n438_));
  NO2        g416(.A(i_6_), .B(i_7_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n439_), .B(new_new_n438_), .Y(new_new_n440_));
  NO2        g418(.A(i_11_), .B(i_1_), .Y(new_new_n441_));
  NOi21      g419(.An(i_2_), .B(i_7_), .Y(new_new_n442_));
  NAi31      g420(.An(i_11_), .B(new_new_n442_), .C(new_new_n930_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n393_), .B(i_6_), .Y(new_new_n444_));
  NA3        g422(.A(new_new_n444_), .B(new_new_n935_), .C(new_new_n73_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n445_), .B(new_new_n443_), .Y(new_new_n446_));
  NO2        g424(.A(i_6_), .B(i_10_), .Y(new_new_n447_));
  NA3        g425(.A(new_new_n447_), .B(new_new_n294_), .C(i_8_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n448_), .B(new_new_n149_), .Y(new_new_n449_));
  NA3        g427(.A(new_new_n232_), .B(new_new_n165_), .C(new_new_n127_), .Y(new_new_n450_));
  NA2        g428(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n151_), .B(i_3_), .Y(new_new_n452_));
  NAi31      g430(.An(new_new_n451_), .B(new_new_n452_), .C(new_new_n215_), .Y(new_new_n453_));
  NA3        g431(.A(new_new_n372_), .B(new_new_n173_), .C(new_new_n143_), .Y(new_new_n454_));
  NA3        g432(.A(new_new_n454_), .B(new_new_n453_), .C(new_new_n450_), .Y(new_new_n455_));
  NO4        g433(.A(new_new_n455_), .B(new_new_n449_), .C(new_new_n446_), .D(new_new_n437_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n426_), .B(new_new_n363_), .Y(new_new_n457_));
  NO2        g435(.A(i_8_), .B(new_new_n213_), .Y(new_new_n458_));
  NAi21      g436(.An(new_new_n205_), .B(new_new_n375_), .Y(new_new_n459_));
  NO2        g437(.A(i_0_), .B(new_new_n82_), .Y(new_new_n460_));
  NA3        g438(.A(new_new_n460_), .B(new_new_n931_), .C(new_new_n136_), .Y(new_new_n461_));
  OR3        g439(.A(new_new_n284_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n461_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n27_), .B(i_10_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n294_), .B(new_new_n226_), .Y(new_new_n465_));
  OAI220     g443(.A0(new_new_n465_), .A1(new_new_n413_), .B0(new_new_n464_), .B1(new_new_n434_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n287_), .B(new_new_n212_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n467_), .B(new_new_n440_), .Y(new_new_n468_));
  NO4        g446(.A(new_new_n468_), .B(new_new_n466_), .C(new_new_n463_), .D(new_new_n458_), .Y(new_new_n469_));
  NA3        g447(.A(new_new_n469_), .B(new_new_n456_), .C(new_new_n433_), .Y(new_new_n470_));
  NA3        g448(.A(new_new_n287_), .B(new_new_n170_), .C(new_new_n168_), .Y(new_new_n471_));
  OAI210     g449(.A0(new_new_n283_), .A1(new_new_n175_), .B0(new_new_n471_), .Y(new_new_n472_));
  BUFFER     g450(.A(new_new_n269_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n118_), .B(new_new_n109_), .Y(new_new_n475_));
  AN2        g453(.A(new_new_n475_), .B(new_new_n426_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n294_), .B(new_new_n158_), .Y(new_new_n477_));
  OAI210     g455(.A0(new_new_n477_), .A1(new_new_n220_), .B0(new_new_n288_), .Y(new_new_n478_));
  AOI220     g456(.A0(new_new_n478_), .A1(i_7_), .B0(new_new_n476_), .B1(new_new_n290_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n363_), .B(new_new_n214_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n337_), .B(new_new_n71_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n350_), .B(new_new_n346_), .Y(new_new_n482_));
  OR2        g460(.A(new_new_n480_), .B(new_new_n482_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n36_), .B(i_8_), .Y(new_new_n484_));
  NAi41      g462(.An(new_new_n481_), .B(new_new_n447_), .C(new_new_n484_), .D(new_new_n46_), .Y(new_new_n485_));
  AOI210     g463(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n394_), .Y(new_new_n486_));
  NA3        g464(.A(new_new_n486_), .B(new_new_n485_), .C(new_new_n483_), .Y(new_new_n487_));
  INV        g465(.A(new_new_n487_), .Y(new_new_n488_));
  INV        g466(.A(new_new_n192_), .Y(new_new_n489_));
  OR2        g467(.A(new_new_n177_), .B(i_4_), .Y(new_new_n490_));
  NO2        g468(.A(new_new_n490_), .B(new_new_n82_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n491_), .B(new_new_n489_), .Y(new_new_n492_));
  NA4        g470(.A(new_new_n492_), .B(new_new_n488_), .C(new_new_n479_), .D(new_new_n474_), .Y(new_new_n493_));
  INV        g471(.A(new_new_n277_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n364_), .A1(new_new_n163_), .B0(new_new_n494_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n926_), .B(new_new_n214_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n447_), .B(new_new_n27_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n497_), .B(new_new_n496_), .Y(new_new_n498_));
  NOi31      g476(.An(new_new_n297_), .B(new_new_n393_), .C(new_new_n38_), .Y(new_new_n499_));
  OAI210     g477(.A0(new_new_n499_), .A1(new_new_n498_), .B0(new_new_n495_), .Y(new_new_n500_));
  NO2        g478(.A(i_8_), .B(i_7_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n46_), .B(new_new_n229_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n44_), .B(i_10_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(i_6_), .Y(new_new_n504_));
  NA3        g482(.A(new_new_n504_), .B(new_new_n502_), .C(new_new_n501_), .Y(new_new_n505_));
  OAI210     g483(.A0(new_new_n177_), .A1(new_new_n250_), .B0(new_new_n434_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n506_), .B(new_new_n253_), .Y(new_new_n507_));
  NOi31      g485(.An(new_new_n272_), .B(new_new_n283_), .C(new_new_n175_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n210_), .B(new_new_n44_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n151_), .B(i_5_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n510_), .B(new_new_n300_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n511_), .B(new_new_n509_), .Y(new_new_n512_));
  OAI210     g490(.A0(new_new_n512_), .A1(new_new_n508_), .B0(new_new_n429_), .Y(new_new_n513_));
  NA4        g491(.A(new_new_n513_), .B(new_new_n507_), .C(new_new_n505_), .D(new_new_n500_), .Y(new_new_n514_));
  NA2        g492(.A(new_new_n69_), .B(new_new_n44_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n266_), .B(new_new_n81_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n515_), .A1(new_new_n329_), .B0(new_new_n516_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n278_), .B(new_new_n269_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(new_new_n167_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n423_), .B(new_new_n210_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n520_), .B(new_new_n521_), .Y(new_new_n522_));
  NO3        g500(.A(new_new_n522_), .B(new_new_n519_), .C(new_new_n517_), .Y(new_new_n523_));
  NO4        g501(.A(new_new_n236_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n524_));
  NO3        g502(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n221_), .B(new_new_n36_), .Y(new_new_n526_));
  AN2        g504(.A(new_new_n526_), .B(new_new_n525_), .Y(new_new_n527_));
  OA210      g505(.A0(new_new_n527_), .A1(new_new_n524_), .B0(new_new_n337_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n393_), .B(i_1_), .Y(new_new_n529_));
  NOi31      g507(.An(new_new_n529_), .B(new_new_n427_), .C(new_new_n71_), .Y(new_new_n530_));
  AN3        g508(.A(new_new_n530_), .B(new_new_n390_), .C(i_2_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n403_), .B(new_new_n171_), .Y(new_new_n532_));
  NO3        g510(.A(new_new_n532_), .B(new_new_n531_), .C(new_new_n528_), .Y(new_new_n533_));
  NOi21      g511(.An(i_10_), .B(i_6_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n535_));
  NA2        g513(.A(new_new_n297_), .B(new_new_n158_), .Y(new_new_n536_));
  AOI220     g514(.A0(new_new_n536_), .A1(new_new_n414_), .B0(new_new_n166_), .B1(new_new_n176_), .Y(new_new_n537_));
  NOi31      g515(.An(new_new_n140_), .B(i_1_), .C(new_new_n312_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n538_), .B(new_new_n537_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n481_), .B(new_new_n358_), .Y(new_new_n540_));
  NO2        g518(.A(i_12_), .B(new_new_n82_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n168_), .B(i_0_), .Y(new_new_n542_));
  NO3        g520(.A(new_new_n542_), .B(new_new_n322_), .C(new_new_n283_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n352_), .B(new_new_n231_), .Y(new_new_n544_));
  AOI210     g522(.A0(new_new_n544_), .A1(i_5_), .B0(new_new_n459_), .Y(new_new_n545_));
  NO3        g523(.A(new_new_n545_), .B(new_new_n543_), .C(new_new_n540_), .Y(new_new_n546_));
  NA4        g524(.A(new_new_n546_), .B(new_new_n539_), .C(new_new_n533_), .D(new_new_n523_), .Y(new_new_n547_));
  NO4        g525(.A(new_new_n547_), .B(new_new_n514_), .C(new_new_n493_), .D(new_new_n470_), .Y(new_new_n548_));
  NA4        g526(.A(new_new_n548_), .B(new_new_n421_), .C(new_new_n336_), .D(new_new_n293_), .Y(mai7));
  NO2        g527(.A(new_new_n91_), .B(new_new_n53_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n447_), .B(new_new_n81_), .Y(new_new_n551_));
  NA3        g529(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n224_), .B(i_4_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n553_), .B(i_8_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n103_), .B(new_new_n552_), .Y(new_new_n555_));
  NA2        g533(.A(i_2_), .B(new_new_n82_), .Y(new_new_n556_));
  OAI210     g534(.A0(new_new_n85_), .A1(new_new_n196_), .B0(new_new_n197_), .Y(new_new_n557_));
  NO2        g535(.A(i_7_), .B(new_new_n37_), .Y(new_new_n558_));
  NA2        g536(.A(i_4_), .B(i_8_), .Y(new_new_n559_));
  AOI210     g537(.A0(new_new_n559_), .A1(new_new_n287_), .B0(new_new_n558_), .Y(new_new_n560_));
  OAI220     g538(.A0(new_new_n560_), .A1(new_new_n556_), .B0(new_new_n557_), .B1(i_13_), .Y(new_new_n561_));
  NO3        g539(.A(new_new_n561_), .B(new_new_n555_), .C(new_new_n550_), .Y(new_new_n562_));
  OR2        g540(.A(i_6_), .B(i_10_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n563_), .B(new_new_n23_), .Y(new_new_n564_));
  OR3        g542(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n565_));
  NO3        g543(.A(new_new_n565_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n566_));
  INV        g544(.A(new_new_n193_), .Y(new_new_n567_));
  NO2        g545(.A(new_new_n566_), .B(new_new_n564_), .Y(new_new_n568_));
  OR2        g546(.A(new_new_n568_), .B(i_3_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n569_), .A1(new_new_n562_), .B0(new_new_n61_), .Y(new_new_n570_));
  NOi21      g548(.An(i_11_), .B(i_7_), .Y(new_new_n571_));
  AO210      g549(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n572_));
  NO2        g550(.A(new_new_n572_), .B(new_new_n571_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n573_), .B(new_new_n198_), .Y(new_new_n574_));
  NA3        g552(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n575_));
  NO2        g553(.A(new_new_n574_), .B(new_new_n61_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n84_), .B(new_new_n61_), .Y(new_new_n577_));
  AO210      g555(.A0(new_new_n577_), .A1(new_new_n358_), .B0(new_new_n41_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n215_), .B(new_new_n61_), .Y(new_new_n579_));
  OR2        g557(.A(new_new_n200_), .B(new_new_n106_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n61_), .B(i_9_), .Y(new_new_n581_));
  NO2        g559(.A(i_1_), .B(i_12_), .Y(new_new_n582_));
  NA2        g560(.A(new_new_n579_), .B(new_new_n578_), .Y(new_new_n583_));
  OAI210     g561(.A0(new_new_n583_), .A1(new_new_n576_), .B0(i_6_), .Y(new_new_n584_));
  NO2        g562(.A(new_new_n575_), .B(new_new_n106_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n585_), .B(new_new_n541_), .Y(new_new_n586_));
  NO2        g564(.A(i_6_), .B(i_11_), .Y(new_new_n587_));
  INV        g565(.A(new_new_n586_), .Y(new_new_n588_));
  NO4        g566(.A(i_12_), .B(new_new_n123_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n589_), .B(new_new_n581_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n224_), .B(i_6_), .Y(new_new_n591_));
  NO3        g569(.A(new_new_n563_), .B(new_new_n221_), .C(new_new_n23_), .Y(new_new_n592_));
  AOI210     g570(.A0(i_1_), .A1(new_new_n245_), .B0(new_new_n592_), .Y(new_new_n593_));
  OAI210     g571(.A0(new_new_n593_), .A1(new_new_n44_), .B0(new_new_n590_), .Y(new_new_n594_));
  NA3        g572(.A(new_new_n501_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n132_), .B(i_9_), .Y(new_new_n596_));
  NA3        g574(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n597_));
  NA3        g575(.A(i_2_), .B(new_new_n254_), .C(new_new_n44_), .Y(new_new_n598_));
  OAI220     g576(.A0(new_new_n598_), .A1(new_new_n597_), .B0(new_new_n596_), .B1(new_new_n925_), .Y(new_new_n599_));
  NA3        g577(.A(new_new_n581_), .B(new_new_n300_), .C(i_6_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n600_), .B(new_new_n23_), .Y(new_new_n601_));
  NA2        g579(.A(i_2_), .B(new_new_n254_), .Y(new_new_n602_));
  NO2        g580(.A(i_11_), .B(new_new_n37_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n603_), .B(new_new_n24_), .Y(new_new_n604_));
  NO2        g582(.A(new_new_n604_), .B(new_new_n602_), .Y(new_new_n605_));
  OR3        g583(.A(new_new_n605_), .B(new_new_n601_), .C(new_new_n599_), .Y(new_new_n606_));
  NO3        g584(.A(new_new_n606_), .B(new_new_n594_), .C(new_new_n588_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n224_), .B(new_new_n99_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n608_), .B(new_new_n571_), .Y(new_new_n609_));
  NA2        g587(.A(new_new_n609_), .B(i_1_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n610_), .B(new_new_n565_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n392_), .B(new_new_n82_), .Y(new_new_n612_));
  INV        g590(.A(new_new_n611_), .Y(new_new_n613_));
  NO2        g591(.A(new_new_n221_), .B(new_new_n44_), .Y(new_new_n614_));
  NO3        g592(.A(new_new_n614_), .B(new_new_n290_), .C(new_new_n225_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n113_), .B(new_new_n37_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n616_), .B(i_6_), .Y(new_new_n617_));
  NO2        g595(.A(new_new_n82_), .B(i_9_), .Y(new_new_n618_));
  NO2        g596(.A(new_new_n618_), .B(new_new_n61_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n619_), .B(new_new_n582_), .Y(new_new_n620_));
  NO4        g598(.A(new_new_n620_), .B(new_new_n617_), .C(new_new_n615_), .D(i_4_), .Y(new_new_n621_));
  NA2        g599(.A(i_1_), .B(i_3_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n428_), .B(new_new_n91_), .Y(new_new_n623_));
  AOI210     g601(.A0(new_new_n614_), .A1(new_new_n534_), .B0(new_new_n623_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n624_), .B(new_new_n622_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n621_), .Y(new_new_n626_));
  NA4        g604(.A(new_new_n626_), .B(new_new_n613_), .C(new_new_n607_), .D(new_new_n584_), .Y(new_new_n627_));
  NO3        g605(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n628_));
  NOi21      g606(.An(new_new_n628_), .B(i_10_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n350_), .B(new_new_n349_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n447_), .B(new_new_n484_), .Y(new_new_n631_));
  NA2        g609(.A(new_new_n631_), .B(new_new_n630_), .Y(new_new_n632_));
  NA2        g610(.A(new_new_n632_), .B(i_1_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n254_), .A1(new_new_n95_), .B0(i_1_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n348_), .B(i_2_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n635_), .B(new_new_n634_), .Y(new_new_n636_));
  AOI210     g614(.A0(new_new_n636_), .A1(new_new_n633_), .B0(i_13_), .Y(new_new_n637_));
  OR2        g615(.A(i_11_), .B(i_7_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n53_), .B(i_12_), .Y(new_new_n639_));
  INV        g617(.A(new_new_n639_), .Y(new_new_n640_));
  AOI220     g618(.A0(i_7_), .A1(new_new_n612_), .B0(new_new_n232_), .B1(new_new_n126_), .Y(new_new_n641_));
  OAI220     g619(.A0(new_new_n641_), .A1(new_new_n41_), .B0(new_new_n640_), .B1(new_new_n91_), .Y(new_new_n642_));
  INV        g620(.A(new_new_n642_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n424_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n644_));
  NOi31      g622(.An(new_new_n644_), .B(new_new_n551_), .C(new_new_n44_), .Y(new_new_n645_));
  NA2        g623(.A(new_new_n122_), .B(i_13_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n597_), .B(new_new_n112_), .Y(new_new_n647_));
  INV        g625(.A(new_new_n647_), .Y(new_new_n648_));
  OAI220     g626(.A0(new_new_n648_), .A1(new_new_n69_), .B0(new_new_n646_), .B1(new_new_n634_), .Y(new_new_n649_));
  AOI220     g627(.A0(new_new_n365_), .A1(i_2_), .B0(new_new_n90_), .B1(new_new_n100_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n650_), .B(new_new_n554_), .Y(new_new_n651_));
  NO3        g629(.A(new_new_n651_), .B(new_new_n649_), .C(new_new_n645_), .Y(new_new_n652_));
  OR2        g630(.A(i_11_), .B(i_6_), .Y(new_new_n653_));
  NA2        g631(.A(new_new_n553_), .B(i_7_), .Y(new_new_n654_));
  AOI210     g632(.A0(new_new_n654_), .A1(new_new_n648_), .B0(new_new_n653_), .Y(new_new_n655_));
  NA3        g633(.A(new_new_n386_), .B(new_new_n558_), .C(new_new_n95_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n587_), .B(i_13_), .Y(new_new_n657_));
  NAi21      g635(.An(i_11_), .B(i_12_), .Y(new_new_n658_));
  NOi41      g636(.An(new_new_n108_), .B(new_new_n658_), .C(i_13_), .D(new_new_n82_), .Y(new_new_n659_));
  INV        g637(.A(new_new_n659_), .Y(new_new_n660_));
  NA3        g638(.A(new_new_n660_), .B(new_new_n657_), .C(new_new_n656_), .Y(new_new_n661_));
  OAI210     g639(.A0(new_new_n661_), .A1(new_new_n655_), .B0(new_new_n61_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n936_), .B(new_new_n347_), .Y(new_new_n663_));
  NO2        g641(.A(new_new_n123_), .B(i_2_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n664_), .B(new_new_n582_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n665_), .B(new_new_n663_), .Y(new_new_n666_));
  NA3        g644(.A(new_new_n666_), .B(new_new_n45_), .C(new_new_n214_), .Y(new_new_n667_));
  NA4        g645(.A(new_new_n667_), .B(new_new_n662_), .C(new_new_n652_), .D(new_new_n643_), .Y(new_new_n668_));
  OR4        g646(.A(new_new_n668_), .B(new_new_n637_), .C(new_new_n627_), .D(new_new_n570_), .Y(mai5));
  NA2        g647(.A(new_new_n609_), .B(new_new_n256_), .Y(new_new_n670_));
  NO2        g648(.A(new_new_n554_), .B(i_11_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n85_), .B(new_new_n671_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n672_), .B(new_new_n670_), .Y(new_new_n673_));
  NO3        g651(.A(i_11_), .B(new_new_n224_), .C(i_13_), .Y(new_new_n674_));
  NA2        g652(.A(i_12_), .B(i_8_), .Y(new_new_n675_));
  INV        g653(.A(new_new_n423_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n535_), .B(new_new_n673_), .Y(new_new_n677_));
  INV        g655(.A(new_new_n165_), .Y(new_new_n678_));
  INV        g656(.A(new_new_n232_), .Y(new_new_n679_));
  OAI210     g657(.A0(new_new_n635_), .A1(new_new_n425_), .B0(new_new_n108_), .Y(new_new_n680_));
  AOI210     g658(.A0(new_new_n680_), .A1(new_new_n679_), .B0(new_new_n678_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n428_), .B(new_new_n26_), .Y(new_new_n682_));
  NO2        g660(.A(new_new_n682_), .B(new_new_n396_), .Y(new_new_n683_));
  AOI210     g661(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n393_), .Y(new_new_n684_));
  AOI210     g662(.A0(new_new_n684_), .A1(i_2_), .B0(new_new_n681_), .Y(new_new_n685_));
  NO3        g663(.A(new_new_n572_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n686_));
  OA210      g664(.A0(new_new_n573_), .A1(new_new_n121_), .B0(i_13_), .Y(new_new_n687_));
  INV        g665(.A(new_new_n145_), .Y(new_new_n688_));
  NO2        g666(.A(new_new_n688_), .B(new_new_n352_), .Y(new_new_n689_));
  NA2        g667(.A(i_2_), .B(new_new_n396_), .Y(new_new_n690_));
  NA3        g668(.A(new_new_n287_), .B(new_new_n119_), .C(new_new_n42_), .Y(new_new_n691_));
  OAI210     g669(.A0(new_new_n691_), .A1(new_new_n46_), .B0(new_new_n690_), .Y(new_new_n692_));
  NO4        g670(.A(new_new_n692_), .B(new_new_n689_), .C(new_new_n687_), .D(new_new_n686_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n674_), .B(new_new_n259_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n60_), .B(i_12_), .Y(new_new_n695_));
  NA4        g673(.A(new_new_n694_), .B(new_new_n693_), .C(new_new_n685_), .D(new_new_n677_), .Y(mai6));
  NO3        g674(.A(new_new_n240_), .B(new_new_n289_), .C(i_1_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n179_), .B(new_new_n133_), .Y(new_new_n698_));
  OAI210     g676(.A0(new_new_n698_), .A1(new_new_n697_), .B0(new_new_n664_), .Y(new_new_n699_));
  INV        g677(.A(new_new_n310_), .Y(new_new_n700_));
  AO210      g678(.A0(new_new_n700_), .A1(new_new_n699_), .B0(i_12_), .Y(new_new_n701_));
  NA2        g679(.A(new_new_n353_), .B(new_new_n317_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n541_), .B(new_new_n61_), .Y(new_new_n703_));
  NA2        g681(.A(new_new_n629_), .B(new_new_n69_), .Y(new_new_n704_));
  BUFFER     g682(.A(new_new_n577_), .Y(new_new_n705_));
  NA4        g683(.A(new_new_n705_), .B(new_new_n704_), .C(new_new_n703_), .D(new_new_n702_), .Y(new_new_n706_));
  NA2        g684(.A(new_new_n706_), .B(new_new_n71_), .Y(new_new_n707_));
  INV        g685(.A(new_new_n309_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n73_), .B(new_new_n126_), .Y(new_new_n709_));
  AOI210     g687(.A0(new_new_n119_), .A1(new_new_n709_), .B0(new_new_n708_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n236_), .B(i_9_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n711_), .B(new_new_n695_), .Y(new_new_n712_));
  AOI210     g690(.A0(new_new_n712_), .A1(new_new_n482_), .B0(new_new_n179_), .Y(new_new_n713_));
  NO2        g691(.A(new_new_n32_), .B(i_11_), .Y(new_new_n714_));
  NA3        g692(.A(new_new_n714_), .B(new_new_n439_), .C(new_new_n368_), .Y(new_new_n715_));
  NAi32      g693(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n653_), .B(new_new_n716_), .Y(new_new_n717_));
  OAI210     g695(.A0(new_new_n628_), .A1(new_new_n526_), .B0(new_new_n525_), .Y(new_new_n718_));
  NAi31      g696(.An(new_new_n717_), .B(new_new_n718_), .C(new_new_n715_), .Y(new_new_n719_));
  OR3        g697(.A(new_new_n719_), .B(new_new_n713_), .C(new_new_n710_), .Y(new_new_n720_));
  NO2        g698(.A(new_new_n638_), .B(i_2_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n722_), .B(new_new_n385_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n723_), .B(new_new_n721_), .Y(new_new_n724_));
  AO210      g702(.A0(new_new_n341_), .A1(new_new_n333_), .B0(new_new_n374_), .Y(new_new_n725_));
  NA3        g703(.A(new_new_n725_), .B(new_new_n241_), .C(i_7_), .Y(new_new_n726_));
  OR2        g704(.A(new_new_n573_), .B(new_new_n425_), .Y(new_new_n727_));
  NA2        g705(.A(new_new_n727_), .B(new_new_n141_), .Y(new_new_n728_));
  OR2        g706(.A(new_new_n676_), .B(new_new_n36_), .Y(new_new_n729_));
  NA4        g707(.A(new_new_n729_), .B(new_new_n728_), .C(new_new_n726_), .D(new_new_n724_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n933_), .B(new_new_n525_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n374_), .B(new_new_n68_), .Y(new_new_n732_));
  NA3        g710(.A(new_new_n732_), .B(new_new_n731_), .C(new_new_n557_), .Y(new_new_n733_));
  OR2        g711(.A(new_new_n484_), .B(new_new_n84_), .Y(new_new_n734_));
  NA3        g712(.A(new_new_n734_), .B(new_new_n447_), .C(new_new_n207_), .Y(new_new_n735_));
  AOI210     g713(.A0(new_new_n425_), .A1(new_new_n423_), .B0(new_new_n524_), .Y(new_new_n736_));
  OAI210     g714(.A0(new_new_n939_), .A1(new_new_n109_), .B0(new_new_n384_), .Y(new_new_n737_));
  NA3        g715(.A(new_new_n737_), .B(new_new_n736_), .C(new_new_n735_), .Y(new_new_n738_));
  NO4        g716(.A(new_new_n738_), .B(new_new_n733_), .C(new_new_n730_), .D(new_new_n720_), .Y(new_new_n739_));
  NA4        g717(.A(new_new_n739_), .B(new_new_n707_), .C(new_new_n701_), .D(new_new_n360_), .Y(mai3));
  NA2        g718(.A(i_12_), .B(i_10_), .Y(new_new_n741_));
  INV        g719(.A(i_0_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n272_), .B(new_new_n940_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n743_), .Y(new_new_n744_));
  NO3        g722(.A(new_new_n928_), .B(new_new_n88_), .C(new_new_n44_), .Y(new_new_n745_));
  OA210      g723(.A0(new_new_n745_), .A1(new_new_n744_), .B0(new_new_n168_), .Y(new_new_n746_));
  NOi21      g724(.An(new_new_n94_), .B(new_new_n683_), .Y(new_new_n747_));
  NO3        g725(.A(new_new_n580_), .B(new_new_n428_), .C(new_new_n126_), .Y(new_new_n748_));
  NO2        g726(.A(new_new_n748_), .B(new_new_n747_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n749_), .B(new_new_n48_), .Y(new_new_n750_));
  NO4        g728(.A(new_new_n356_), .B(new_new_n363_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n751_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n644_), .B(new_new_n618_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n315_), .B(i_5_), .Y(new_new_n754_));
  OAI220     g732(.A0(new_new_n754_), .A1(new_new_n753_), .B0(new_new_n752_), .B1(new_new_n61_), .Y(new_new_n755_));
  NOi21      g733(.An(i_5_), .B(i_9_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n756_), .B(new_new_n422_), .Y(new_new_n757_));
  BUFFER     g735(.A(new_new_n254_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n758_), .B(new_new_n441_), .Y(new_new_n759_));
  NO2        g737(.A(new_new_n169_), .B(new_new_n142_), .Y(new_new_n760_));
  INV        g738(.A(new_new_n760_), .Y(new_new_n761_));
  OAI220     g739(.A0(new_new_n761_), .A1(new_new_n175_), .B0(new_new_n759_), .B1(new_new_n757_), .Y(new_new_n762_));
  NO4        g740(.A(new_new_n762_), .B(new_new_n755_), .C(new_new_n750_), .D(new_new_n746_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n179_), .B(new_new_n24_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n294_), .B(new_new_n124_), .Y(new_new_n765_));
  NAi21      g743(.An(new_new_n156_), .B(i_5_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n765_), .B(new_new_n376_), .Y(new_new_n767_));
  INV        g745(.A(new_new_n767_), .Y(new_new_n768_));
  NO2        g746(.A(new_new_n368_), .B(new_new_n276_), .Y(new_new_n769_));
  NA2        g747(.A(new_new_n769_), .B(new_new_n647_), .Y(new_new_n770_));
  AN2        g748(.A(new_new_n94_), .B(new_new_n230_), .Y(new_new_n771_));
  NA2        g749(.A(new_new_n674_), .B(new_new_n310_), .Y(new_new_n772_));
  AOI210     g750(.A0(new_new_n447_), .A1(new_new_n85_), .B0(new_new_n56_), .Y(new_new_n773_));
  NO2        g751(.A(new_new_n773_), .B(new_new_n772_), .Y(new_new_n774_));
  NO2        g752(.A(new_new_n238_), .B(new_new_n147_), .Y(new_new_n775_));
  NA2        g753(.A(i_0_), .B(i_10_), .Y(new_new_n776_));
  AN2        g754(.A(new_new_n775_), .B(i_6_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n315_), .B(new_new_n96_), .Y(new_new_n778_));
  NA2        g756(.A(new_new_n529_), .B(i_4_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n182_), .B(new_new_n196_), .Y(new_new_n780_));
  OAI220     g758(.A0(new_new_n780_), .A1(new_new_n772_), .B0(new_new_n779_), .B1(new_new_n778_), .Y(new_new_n781_));
  NO4        g759(.A(new_new_n781_), .B(new_new_n777_), .C(new_new_n774_), .D(new_new_n771_), .Y(new_new_n782_));
  NA3        g760(.A(new_new_n782_), .B(new_new_n770_), .C(new_new_n768_), .Y(new_new_n783_));
  NA2        g761(.A(i_11_), .B(i_9_), .Y(new_new_n784_));
  NO2        g762(.A(new_new_n48_), .B(i_7_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n372_), .B(new_new_n173_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n786_), .B(new_new_n154_), .Y(new_new_n787_));
  NO2        g765(.A(new_new_n784_), .B(new_new_n71_), .Y(new_new_n788_));
  NO2        g766(.A(new_new_n169_), .B(i_0_), .Y(new_new_n789_));
  NA2        g767(.A(new_new_n439_), .B(new_new_n219_), .Y(new_new_n790_));
  INV        g768(.A(new_new_n383_), .Y(new_new_n791_));
  OAI220     g769(.A0(new_new_n791_), .A1(new_new_n757_), .B0(new_new_n790_), .B1(new_new_n169_), .Y(new_new_n792_));
  NO2        g770(.A(new_new_n792_), .B(new_new_n787_), .Y(new_new_n793_));
  NA2        g771(.A(new_new_n603_), .B(new_new_n117_), .Y(new_new_n794_));
  NO2        g772(.A(i_6_), .B(new_new_n794_), .Y(new_new_n795_));
  AOI210     g773(.A0(new_new_n424_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n796_));
  NA2        g774(.A(new_new_n165_), .B(new_new_n101_), .Y(new_new_n797_));
  NOi32      g775(.An(new_new_n796_), .Bn(new_new_n182_), .C(new_new_n797_), .Y(new_new_n798_));
  NO2        g776(.A(new_new_n798_), .B(new_new_n795_), .Y(new_new_n799_));
  NOi21      g777(.An(i_7_), .B(i_5_), .Y(new_new_n800_));
  NOi31      g778(.An(new_new_n800_), .B(i_0_), .C(new_new_n658_), .Y(new_new_n801_));
  NA3        g779(.A(new_new_n801_), .B(new_new_n937_), .C(i_6_), .Y(new_new_n802_));
  OA210      g780(.A0(new_new_n797_), .A1(new_new_n482_), .B0(new_new_n802_), .Y(new_new_n803_));
  NO3        g781(.A(new_new_n379_), .B(new_new_n344_), .C(new_new_n340_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n248_), .B(new_new_n301_), .Y(new_new_n805_));
  NO2        g783(.A(new_new_n658_), .B(new_new_n243_), .Y(new_new_n806_));
  AOI210     g784(.A0(new_new_n806_), .A1(new_new_n805_), .B0(new_new_n804_), .Y(new_new_n807_));
  NA4        g785(.A(new_new_n807_), .B(new_new_n803_), .C(new_new_n799_), .D(new_new_n793_), .Y(new_new_n808_));
  NO2        g786(.A(new_new_n764_), .B(new_new_n227_), .Y(new_new_n809_));
  AN2        g787(.A(new_new_n314_), .B(new_new_n310_), .Y(new_new_n810_));
  AN2        g788(.A(new_new_n810_), .B(new_new_n760_), .Y(new_new_n811_));
  OAI210     g789(.A0(new_new_n811_), .A1(new_new_n809_), .B0(i_10_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n741_), .B(new_new_n300_), .Y(new_new_n813_));
  OA210      g791(.A0(new_new_n439_), .A1(new_new_n212_), .B0(new_new_n438_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n813_), .B(new_new_n788_), .Y(new_new_n815_));
  NA3        g793(.A(new_new_n438_), .B(new_new_n386_), .C(new_new_n45_), .Y(new_new_n816_));
  OAI210     g794(.A0(new_new_n766_), .A1(i_6_), .B0(new_new_n816_), .Y(new_new_n817_));
  NO2        g795(.A(new_new_n241_), .B(new_new_n46_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n818_), .B(new_new_n181_), .Y(new_new_n819_));
  AOI220     g797(.A0(new_new_n819_), .A1(new_new_n439_), .B0(new_new_n817_), .B1(new_new_n71_), .Y(new_new_n820_));
  NA3        g798(.A(new_new_n722_), .B(new_new_n362_), .C(i_6_), .Y(new_new_n821_));
  NA2        g799(.A(new_new_n91_), .B(new_new_n44_), .Y(new_new_n822_));
  NO2        g800(.A(new_new_n73_), .B(new_new_n675_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n823_), .B(new_new_n822_), .Y(new_new_n824_));
  AOI210     g802(.A0(new_new_n824_), .A1(new_new_n821_), .B0(new_new_n47_), .Y(new_new_n825_));
  NO2        g803(.A(new_new_n552_), .B(new_new_n103_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n826_), .B(i_0_), .Y(new_new_n827_));
  NO2        g805(.A(new_new_n827_), .B(new_new_n82_), .Y(new_new_n828_));
  NO3        g806(.A(new_new_n828_), .B(new_new_n825_), .C(new_new_n487_), .Y(new_new_n829_));
  NA4        g807(.A(new_new_n829_), .B(new_new_n820_), .C(new_new_n815_), .D(new_new_n812_), .Y(new_new_n830_));
  NO3        g808(.A(new_new_n830_), .B(new_new_n808_), .C(new_new_n783_), .Y(new_new_n831_));
  AOI210     g809(.A0(new_new_n703_), .A1(new_new_n630_), .B0(new_new_n797_), .Y(new_new_n832_));
  AOI210     g810(.A0(new_new_n168_), .A1(new_new_n330_), .B0(new_new_n832_), .Y(new_new_n833_));
  NO2        g811(.A(new_new_n718_), .B(new_new_n379_), .Y(new_new_n834_));
  NA3        g812(.A(new_new_n742_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n835_));
  NA2        g813(.A(new_new_n940_), .B(i_9_), .Y(new_new_n836_));
  AOI210     g814(.A0(new_new_n835_), .A1(new_new_n461_), .B0(new_new_n836_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n834_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n833_), .Y(new_new_n839_));
  NA2        g817(.A(new_new_n810_), .B(new_new_n352_), .Y(new_new_n840_));
  AOI210     g818(.A0(new_new_n283_), .A1(new_new_n156_), .B0(new_new_n840_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n785_), .B(new_new_n452_), .Y(new_new_n842_));
  AOI210     g820(.A0(i_11_), .A1(new_new_n156_), .B0(new_new_n842_), .Y(new_new_n843_));
  NO2        g821(.A(new_new_n843_), .B(new_new_n841_), .Y(new_new_n844_));
  NO3        g822(.A(new_new_n776_), .B(new_new_n756_), .C(new_new_n184_), .Y(new_new_n845_));
  AOI220     g823(.A0(new_new_n845_), .A1(i_11_), .B0(new_new_n530_), .B1(new_new_n73_), .Y(new_new_n846_));
  NO3        g824(.A(new_new_n201_), .B(new_new_n363_), .C(i_0_), .Y(new_new_n847_));
  OAI210     g825(.A0(new_new_n847_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n848_));
  OAI220     g826(.A0(new_new_n496_), .A1(new_new_n133_), .B0(new_new_n591_), .B1(new_new_n567_), .Y(new_new_n849_));
  NA3        g827(.A(new_new_n849_), .B(i_7_), .C(i_0_), .Y(new_new_n850_));
  NA4        g828(.A(new_new_n850_), .B(new_new_n848_), .C(new_new_n846_), .D(new_new_n844_), .Y(new_new_n851_));
  NA2        g829(.A(new_new_n333_), .B(new_new_n170_), .Y(new_new_n852_));
  OR2        g830(.A(new_new_n852_), .B(new_new_n929_), .Y(new_new_n853_));
  AOI210     g831(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n854_), .B(new_new_n814_), .Y(new_new_n855_));
  NA3        g833(.A(new_new_n564_), .B(new_new_n179_), .C(new_new_n81_), .Y(new_new_n856_));
  INV        g834(.A(new_new_n856_), .Y(new_new_n857_));
  NO3        g835(.A(new_new_n938_), .B(new_new_n53_), .C(new_new_n48_), .Y(new_new_n858_));
  NA2        g836(.A(new_new_n457_), .B(new_new_n450_), .Y(new_new_n859_));
  NO3        g837(.A(new_new_n859_), .B(new_new_n858_), .C(new_new_n857_), .Y(new_new_n860_));
  NA3        g838(.A(new_new_n368_), .B(new_new_n165_), .C(new_new_n164_), .Y(new_new_n861_));
  INV        g839(.A(new_new_n861_), .Y(new_new_n862_));
  NA3        g840(.A(new_new_n368_), .B(new_new_n316_), .C(new_new_n210_), .Y(new_new_n863_));
  INV        g841(.A(new_new_n863_), .Y(new_new_n864_));
  NO3        g842(.A(new_new_n784_), .B(new_new_n207_), .C(new_new_n184_), .Y(new_new_n865_));
  NO3        g843(.A(new_new_n865_), .B(new_new_n864_), .C(new_new_n862_), .Y(new_new_n866_));
  NA4        g844(.A(new_new_n866_), .B(new_new_n860_), .C(new_new_n855_), .D(new_new_n853_), .Y(new_new_n867_));
  INV        g845(.A(new_new_n566_), .Y(new_new_n868_));
  NO3        g846(.A(new_new_n868_), .B(i_5_), .C(new_new_n327_), .Y(new_new_n869_));
  INV        g847(.A(new_new_n869_), .Y(new_new_n870_));
  NA2        g848(.A(new_new_n287_), .B(i_5_), .Y(new_new_n871_));
  NO4        g849(.A(new_new_n227_), .B(new_new_n201_), .C(i_0_), .D(i_12_), .Y(new_new_n872_));
  NA2        g850(.A(new_new_n872_), .B(i_10_), .Y(new_new_n873_));
  AN2        g851(.A(new_new_n776_), .B(new_new_n147_), .Y(new_new_n874_));
  NO4        g852(.A(new_new_n874_), .B(i_12_), .C(new_new_n595_), .D(new_new_n126_), .Y(new_new_n875_));
  INV        g853(.A(new_new_n875_), .Y(new_new_n876_));
  NA3        g854(.A(new_new_n96_), .B(new_new_n534_), .C(i_11_), .Y(new_new_n877_));
  NA2        g855(.A(new_new_n800_), .B(new_new_n436_), .Y(new_new_n878_));
  OAI220     g856(.A0(i_7_), .A1(new_new_n871_), .B0(new_new_n878_), .B1(new_new_n619_), .Y(new_new_n879_));
  NA2        g857(.A(new_new_n879_), .B(new_new_n789_), .Y(new_new_n880_));
  NA4        g858(.A(new_new_n880_), .B(new_new_n876_), .C(new_new_n873_), .D(new_new_n870_), .Y(new_new_n881_));
  NO4        g859(.A(new_new_n881_), .B(new_new_n867_), .C(new_new_n851_), .D(new_new_n839_), .Y(new_new_n882_));
  OAI210     g860(.A0(new_new_n721_), .A1(new_new_n714_), .B0(new_new_n37_), .Y(new_new_n883_));
  NA3        g861(.A(new_new_n796_), .B(new_new_n347_), .C(i_5_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n884_), .B(new_new_n883_), .Y(new_new_n885_));
  NA2        g863(.A(new_new_n885_), .B(new_new_n198_), .Y(new_new_n886_));
  BUFFER     g864(.A(new_new_n348_), .Y(new_new_n887_));
  NA2        g865(.A(new_new_n180_), .B(new_new_n182_), .Y(new_new_n888_));
  AO210      g866(.A0(new_new_n887_), .A1(new_new_n33_), .B0(new_new_n888_), .Y(new_new_n889_));
  OAI210     g867(.A0(new_new_n566_), .A1(new_new_n564_), .B0(new_new_n300_), .Y(new_new_n890_));
  NAi31      g868(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n891_));
  NO2        g869(.A(new_new_n68_), .B(new_new_n891_), .Y(new_new_n892_));
  NO2        g870(.A(new_new_n892_), .B(new_new_n592_), .Y(new_new_n893_));
  NA3        g871(.A(new_new_n893_), .B(new_new_n890_), .C(new_new_n889_), .Y(new_new_n894_));
  NO2        g872(.A(new_new_n430_), .B(new_new_n254_), .Y(new_new_n895_));
  NO4        g873(.A(new_new_n221_), .B(new_new_n139_), .C(new_new_n622_), .D(new_new_n37_), .Y(new_new_n896_));
  NO2        g874(.A(new_new_n896_), .B(new_new_n895_), .Y(new_new_n897_));
  OAI210     g875(.A0(new_new_n877_), .A1(new_new_n142_), .B0(new_new_n897_), .Y(new_new_n898_));
  AOI210     g876(.A0(new_new_n894_), .A1(new_new_n48_), .B0(new_new_n898_), .Y(new_new_n899_));
  AOI210     g877(.A0(new_new_n899_), .A1(new_new_n886_), .B0(new_new_n71_), .Y(new_new_n900_));
  NO2        g878(.A(new_new_n527_), .B(new_new_n359_), .Y(new_new_n901_));
  NO2        g879(.A(new_new_n901_), .B(new_new_n678_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n53_), .B(new_new_n106_), .Y(new_new_n903_));
  NA2        g881(.A(new_new_n903_), .B(new_new_n74_), .Y(new_new_n904_));
  AOI210     g882(.A0(new_new_n854_), .A1(new_new_n785_), .B0(new_new_n801_), .Y(new_new_n905_));
  AOI210     g883(.A0(new_new_n905_), .A1(new_new_n904_), .B0(new_new_n622_), .Y(new_new_n906_));
  NA2        g884(.A(new_new_n248_), .B(new_new_n55_), .Y(new_new_n907_));
  AOI220     g885(.A0(new_new_n907_), .A1(new_new_n74_), .B0(new_new_n328_), .B1(new_new_n240_), .Y(new_new_n908_));
  NO2        g886(.A(new_new_n908_), .B(new_new_n224_), .Y(new_new_n909_));
  NA3        g887(.A(new_new_n94_), .B(new_new_n289_), .C(new_new_n31_), .Y(new_new_n910_));
  INV        g888(.A(new_new_n910_), .Y(new_new_n911_));
  NO3        g889(.A(new_new_n911_), .B(new_new_n909_), .C(new_new_n906_), .Y(new_new_n912_));
  OAI210     g890(.A0(new_new_n255_), .A1(new_new_n152_), .B0(new_new_n85_), .Y(new_new_n913_));
  NA3        g891(.A(new_new_n682_), .B(new_new_n272_), .C(new_new_n78_), .Y(new_new_n914_));
  AOI210     g892(.A0(new_new_n914_), .A1(new_new_n913_), .B0(i_11_), .Y(new_new_n915_));
  OAI210     g893(.A0(new_new_n927_), .A1(new_new_n796_), .B0(new_new_n198_), .Y(new_new_n916_));
  NA2        g894(.A(new_new_n158_), .B(i_5_), .Y(new_new_n917_));
  NO2        g895(.A(new_new_n916_), .B(new_new_n917_), .Y(new_new_n918_));
  NO2        g896(.A(new_new_n918_), .B(new_new_n915_), .Y(new_new_n919_));
  OAI210     g897(.A0(new_new_n912_), .A1(i_4_), .B0(new_new_n919_), .Y(new_new_n920_));
  NO3        g898(.A(new_new_n920_), .B(new_new_n902_), .C(new_new_n900_), .Y(new_new_n921_));
  NA4        g899(.A(new_new_n921_), .B(new_new_n882_), .C(new_new_n831_), .D(new_new_n763_), .Y(mai4));
  INV        g900(.A(i_2_), .Y(new_new_n925_));
  INV        g901(.A(i_12_), .Y(new_new_n926_));
  INV        g902(.A(i_12_), .Y(new_new_n927_));
  INV        g903(.A(i_0_), .Y(new_new_n928_));
  INV        g904(.A(new_new_n157_), .Y(new_new_n929_));
  INV        g905(.A(i_3_), .Y(new_new_n930_));
  INV        g906(.A(i_5_), .Y(new_new_n931_));
  INV        g907(.A(new_new_n233_), .Y(new_new_n932_));
  INV        g908(.A(i_11_), .Y(new_new_n933_));
  INV        g909(.A(i_12_), .Y(new_new_n934_));
  INV        g910(.A(i_4_), .Y(new_new_n935_));
  INV        g911(.A(i_9_), .Y(new_new_n936_));
  INV        g912(.A(i_4_), .Y(new_new_n937_));
  INV        g913(.A(new_new_n386_), .Y(new_new_n938_));
  INV        g914(.A(new_new_n563_), .Y(new_new_n939_));
  INV        g915(.A(i_11_), .Y(new_new_n940_));
endmodule


