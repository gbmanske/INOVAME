module ex4(
	input[3:0] A,B,
	input[2:0] C,D,
	output [5:0] S6,
	output [4:0] S5,
	output [3:0] S4,
	output [2:0] S3
);

	assign S6 = A+B;
	
	assign S5 = A+B;
	
	assign S4 = A+B;
	
	assign S3 = C+D;
	
	
	
endmodule



