//Benchmark atmr_intb_466_0.25

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n230_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n295_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n350_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  INV        o026(.A(x09), .Y(ori_ori_n49_));
  NO2        o027(.A(x10), .B(x02), .Y(ori_ori_n50_));
  NOi21      o028(.An(x01), .B(x09), .Y(ori_ori_n51_));
  INV        o029(.A(x00), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n49_), .B(ori_ori_n52_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(ori_ori_n51_), .Y(ori_ori_n54_));
  NA2        o032(.A(x09), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  INV        o033(.A(x07), .Y(ori_ori_n56_));
  INV        o034(.A(ori_ori_n54_), .Y(ori_ori_n57_));
  NA2        o035(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(ori_ori_n24_), .Y(ori_ori_n59_));
  NO2        o037(.A(ori_ori_n59_), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n56_), .B(ori_ori_n48_), .Y(ori_ori_n61_));
  OAI210     o039(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n61_), .Y(ori_ori_n62_));
  AOI220     o040(.A0(ori_ori_n62_), .A1(ori_ori_n54_), .B0(ori_ori_n60_), .B1(ori_ori_n31_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(x05), .Y(ori_ori_n64_));
  NA2        o042(.A(x09), .B(x05), .Y(ori_ori_n65_));
  NA2        o043(.A(x10), .B(x06), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n67_), .B(x03), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n69_));
  NO2        o047(.A(x08), .B(x01), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n35_), .Y(ori_ori_n71_));
  NA2        o049(.A(ori_ori_n49_), .B(ori_ori_n36_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n71_), .B(x02), .Y(ori_ori_n73_));
  AN2        o051(.A(ori_ori_n73_), .B(ori_ori_n68_), .Y(ori_ori_n74_));
  INV        o052(.A(ori_ori_n71_), .Y(ori_ori_n75_));
  NA2        o053(.A(x11), .B(x00), .Y(ori_ori_n76_));
  NO2        o054(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n77_));
  NOi21      o055(.An(ori_ori_n76_), .B(ori_ori_n77_), .Y(ori_ori_n78_));
  INV        o056(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NOi21      o057(.An(x01), .B(x10), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n29_), .B(ori_ori_n52_), .Y(ori_ori_n81_));
  NO3        o059(.A(ori_ori_n81_), .B(ori_ori_n80_), .C(x06), .Y(ori_ori_n82_));
  NA2        o060(.A(ori_ori_n82_), .B(ori_ori_n27_), .Y(ori_ori_n83_));
  OAI210     o061(.A0(ori_ori_n79_), .A1(x07), .B0(ori_ori_n83_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n74_), .C(ori_ori_n64_), .Y(ori01));
  INV        o063(.A(x12), .Y(ori_ori_n86_));
  INV        o064(.A(x13), .Y(ori_ori_n87_));
  NO2        o065(.A(x10), .B(x01), .Y(ori_ori_n88_));
  NO2        o066(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n89_));
  NOi21      o067(.An(ori_ori_n89_), .B(ori_ori_n53_), .Y(ori_ori_n90_));
  INV        o068(.A(x13), .Y(ori_ori_n91_));
  NA2        o069(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(x05), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n94_));
  NA2        o072(.A(x10), .B(ori_ori_n52_), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n95_), .B(ori_ori_n94_), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n55_), .B(x05), .Y(ori_ori_n97_));
  NO3        o075(.A(ori_ori_n94_), .B(x06), .C(x03), .Y(ori_ori_n98_));
  INV        o076(.A(ori_ori_n98_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n49_), .B(ori_ori_n41_), .Y(ori_ori_n100_));
  NA2        o078(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n101_));
  NO2        o079(.A(x09), .B(x05), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n102_), .B(ori_ori_n47_), .Y(ori_ori_n103_));
  NA2        o081(.A(x09), .B(x00), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n89_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o083(.A(x03), .B(x02), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n71_), .B(ori_ori_n87_), .Y(ori_ori_n107_));
  OAI210     o085(.A0(ori_ori_n107_), .A1(ori_ori_n90_), .B0(ori_ori_n106_), .Y(ori_ori_n108_));
  OAI210     o086(.A0(ori_ori_n99_), .A1(ori_ori_n23_), .B0(ori_ori_n108_), .Y(ori_ori_n109_));
  NAi21      o087(.An(x06), .B(x10), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n111_));
  INV        o089(.A(x05), .Y(ori_ori_n112_));
  NO2        o090(.A(x09), .B(x01), .Y(ori_ori_n113_));
  NAi21      o091(.An(x13), .B(x00), .Y(ori_ori_n114_));
  INV        o092(.A(ori_ori_n81_), .Y(ori_ori_n115_));
  NOi21      o093(.An(x09), .B(x00), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n47_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n117_), .B(ori_ori_n95_), .Y(ori_ori_n118_));
  NA2        o096(.A(x06), .B(x05), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(ori_ori_n86_), .Y(ori_ori_n120_));
  AOI210     o098(.A0(x10), .A1(ori_ori_n53_), .B0(ori_ori_n120_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n121_), .B(ori_ori_n118_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n87_), .B(x12), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n124_), .B(ori_ori_n122_), .Y(ori_ori_n126_));
  INV        o104(.A(ori_ori_n126_), .Y(ori_ori_n127_));
  AOI210     o105(.A0(ori_ori_n109_), .A1(ori_ori_n86_), .B0(ori_ori_n127_), .Y(ori_ori_n128_));
  NO2        o106(.A(ori_ori_n80_), .B(x06), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n129_), .B(ori_ori_n41_), .Y(ori_ori_n130_));
  INV        o108(.A(ori_ori_n101_), .Y(ori_ori_n131_));
  OAI210     o109(.A0(ori_ori_n131_), .A1(ori_ori_n130_), .B0(x02), .Y(ori_ori_n132_));
  AOI210     o110(.A0(ori_ori_n132_), .A1(ori_ori_n52_), .B0(ori_ori_n23_), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n52_), .B(ori_ori_n133_), .Y(ori_ori_n134_));
  INV        o112(.A(ori_ori_n101_), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n49_), .B(x03), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n137_));
  INV        o115(.A(ori_ori_n110_), .Y(ori_ori_n138_));
  NOi21      o116(.An(x13), .B(x04), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n139_), .B(ori_ori_n116_), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n140_), .B(x05), .Y(ori_ori_n141_));
  AOI220     o119(.A0(ori_ori_n141_), .A1(ori_ori_n137_), .B0(ori_ori_n138_), .B1(ori_ori_n52_), .Y(ori_ori_n142_));
  INV        o120(.A(ori_ori_n142_), .Y(ori_ori_n143_));
  INV        o121(.A(ori_ori_n77_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n144_), .B(x12), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n49_), .B(ori_ori_n36_), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n148_));
  NA2        o126(.A(x13), .B(ori_ori_n86_), .Y(ori_ori_n149_));
  NA3        o127(.A(ori_ori_n149_), .B(ori_ori_n120_), .C(ori_ori_n78_), .Y(ori_ori_n150_));
  INV        o128(.A(ori_ori_n150_), .Y(ori_ori_n151_));
  AOI210     o129(.A0(ori_ori_n145_), .A1(ori_ori_n143_), .B0(ori_ori_n151_), .Y(ori_ori_n152_));
  AOI210     o130(.A0(ori_ori_n152_), .A1(ori_ori_n134_), .B0(x07), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n65_), .B(ori_ori_n29_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n139_), .B(ori_ori_n116_), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NO2        o134(.A(x12), .B(x02), .Y(ori_ori_n157_));
  INV        o135(.A(ori_ori_n157_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n158_), .B(ori_ori_n144_), .Y(ori_ori_n159_));
  AN2        o137(.A(ori_ori_n156_), .B(ori_ori_n159_), .Y(ori_ori_n160_));
  NO2        o138(.A(x02), .B(ori_ori_n91_), .Y(ori_ori_n161_));
  NO3        o139(.A(ori_ori_n76_), .B(x12), .C(x03), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n161_), .B(ori_ori_n162_), .Y(ori_ori_n163_));
  NOi21      o141(.An(ori_ori_n154_), .B(ori_ori_n129_), .Y(ori_ori_n164_));
  NO2        o142(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n164_), .B(ori_ori_n165_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n53_), .B(x05), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n167_), .B(ori_ori_n115_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n146_), .B(ori_ori_n28_), .Y(ori_ori_n169_));
  OAI210     o147(.A0(ori_ori_n168_), .A1(ori_ori_n135_), .B0(ori_ori_n169_), .Y(ori_ori_n170_));
  NA3        o148(.A(ori_ori_n170_), .B(ori_ori_n166_), .C(ori_ori_n163_), .Y(ori_ori_n171_));
  NO3        o149(.A(ori_ori_n171_), .B(ori_ori_n160_), .C(ori_ori_n153_), .Y(ori_ori_n172_));
  OAI210     o150(.A0(ori_ori_n128_), .A1(ori_ori_n56_), .B0(ori_ori_n172_), .Y(ori02));
  INV        o151(.A(ori_ori_n113_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n174_), .B(ori_ori_n32_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n112_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n107_), .B(ori_ori_n106_), .Y(ori_ori_n177_));
  AOI210     o155(.A0(ori_ori_n177_), .A1(ori_ori_n176_), .B0(ori_ori_n48_), .Y(ori_ori_n178_));
  NO2        o156(.A(x05), .B(x02), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n116_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n180_), .B(ori_ori_n101_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n148_), .B(ori_ori_n47_), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n182_), .B(ori_ori_n141_), .Y(ori_ori_n183_));
  BUFFER     o161(.A(ori_ori_n103_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n184_), .B(x06), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n185_), .B(ori_ori_n81_), .Y(ori_ori_n186_));
  INV        o164(.A(ori_ori_n106_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n187_), .B(ori_ori_n96_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n188_), .B(x13), .Y(ori_ori_n189_));
  NA3        o167(.A(ori_ori_n189_), .B(ori_ori_n186_), .C(ori_ori_n183_), .Y(ori_ori_n190_));
  NO3        o168(.A(ori_ori_n190_), .B(ori_ori_n181_), .C(ori_ori_n178_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n100_), .B(x03), .Y(ori_ori_n192_));
  OAI210     o170(.A0(ori_ori_n114_), .A1(ori_ori_n167_), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n193_), .B(ori_ori_n88_), .Y(ori_ori_n194_));
  NA2        o172(.A(x12), .B(ori_ori_n96_), .Y(ori_ori_n195_));
  NA3        o173(.A(ori_ori_n195_), .B(ori_ori_n194_), .C(ori_ori_n48_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n125_), .Y(ori_ori_n197_));
  NA2        o175(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n198_));
  OAI210     o176(.A0(ori_ori_n197_), .A1(ori_ori_n54_), .B0(ori_ori_n198_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n199_), .B(x02), .Y(ori_ori_n200_));
  INV        o178(.A(ori_ori_n147_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n123_), .B(x04), .Y(ori_ori_n202_));
  NO3        o180(.A(ori_ori_n123_), .B(ori_ori_n111_), .C(ori_ori_n50_), .Y(ori_ori_n203_));
  OAI210     o181(.A0(ori_ori_n104_), .A1(ori_ori_n36_), .B0(ori_ori_n86_), .Y(ori_ori_n204_));
  OAI210     o182(.A0(ori_ori_n204_), .A1(ori_ori_n117_), .B0(ori_ori_n203_), .Y(ori_ori_n205_));
  NA3        o183(.A(ori_ori_n205_), .B(ori_ori_n200_), .C(x06), .Y(ori_ori_n206_));
  NA2        o184(.A(x09), .B(x03), .Y(ori_ori_n207_));
  OAI220     o185(.A0(ori_ori_n207_), .A1(ori_ori_n95_), .B0(x01), .B1(ori_ori_n58_), .Y(ori_ori_n208_));
  NO3        o186(.A(ori_ori_n89_), .B(ori_ori_n95_), .C(ori_ori_n38_), .Y(ori_ori_n209_));
  AO220      o187(.A0(ori_ori_n209_), .A1(x04), .B0(ori_ori_n208_), .B1(x05), .Y(ori_ori_n210_));
  AOI210     o188(.A0(ori_ori_n206_), .A1(ori_ori_n196_), .B0(ori_ori_n210_), .Y(ori_ori_n211_));
  OAI210     o189(.A0(ori_ori_n191_), .A1(x12), .B0(ori_ori_n211_), .Y(ori03));
  OR2        o190(.A(ori_ori_n42_), .B(ori_ori_n136_), .Y(ori_ori_n213_));
  AOI210     o191(.A0(ori_ori_n107_), .A1(ori_ori_n86_), .B0(ori_ori_n213_), .Y(ori_ori_n214_));
  AO210      o192(.A0(ori_ori_n201_), .A1(ori_ori_n72_), .B0(ori_ori_n202_), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n123_), .B(ori_ori_n106_), .Y(ori_ori_n216_));
  NA2        o194(.A(ori_ori_n216_), .B(ori_ori_n215_), .Y(ori_ori_n217_));
  OAI210     o195(.A0(ori_ori_n217_), .A1(ori_ori_n214_), .B0(x05), .Y(ori_ori_n218_));
  INV        o196(.A(ori_ori_n93_), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n219_), .B(ori_ori_n54_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n220_), .B(ori_ori_n86_), .Y(ori_ori_n221_));
  AOI210     o199(.A0(ori_ori_n103_), .A1(ori_ori_n55_), .B0(ori_ori_n38_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n113_), .B(ori_ori_n97_), .Y(ori_ori_n223_));
  OAI220     o201(.A0(ori_ori_n223_), .A1(ori_ori_n37_), .B0(ori_ori_n105_), .B1(x13), .Y(ori_ori_n224_));
  OAI210     o202(.A0(ori_ori_n224_), .A1(ori_ori_n222_), .B0(x04), .Y(ori_ori_n225_));
  AOI210     o203(.A0(ori_ori_n114_), .A1(ori_ori_n86_), .B0(ori_ori_n103_), .Y(ori_ori_n226_));
  AN2        o204(.A(x12), .B(ori_ori_n97_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  NA4        o206(.A(ori_ori_n228_), .B(ori_ori_n225_), .C(ori_ori_n221_), .D(ori_ori_n218_), .Y(ori04));
  NO2        o207(.A(ori_ori_n75_), .B(ori_ori_n39_), .Y(ori_ori_n230_));
  XO2        o208(.A(ori_ori_n230_), .B(ori_ori_n149_), .Y(ori05));
  NA2        o209(.A(ori_ori_n86_), .B(x07), .Y(ori_ori_n232_));
  INV        o210(.A(x08), .Y(ori_ori_n233_));
  NA2        o211(.A(x14), .B(ori_ori_n114_), .Y(ori_ori_n234_));
  INV        o212(.A(ori_ori_n44_), .Y(ori_ori_n235_));
  OAI210     o213(.A0(ori_ori_n235_), .A1(ori_ori_n89_), .B0(ori_ori_n86_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NO4        o215(.A(ori_ori_n237_), .B(ori_ori_n234_), .C(ori_ori_n233_), .D(ori_ori_n232_), .Y(ori06));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  INV        m030(.A(mai_mai_n52_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA3        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n28_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(x11), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n338_), .B(mai_mai_n24_), .Y(mai_mai_n76_));
  NO2        m054(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n77_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n48_), .B(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n80_));
  NO2        m058(.A(x08), .B(x01), .Y(mai_mai_n81_));
  OAI210     m059(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n35_), .Y(mai_mai_n82_));
  NO3        m060(.A(mai_mai_n82_), .B(mai_mai_n79_), .C(mai_mai_n76_), .Y(mai_mai_n83_));
  AN2        m061(.A(mai_mai_n83_), .B(mai_mai_n74_), .Y(mai_mai_n84_));
  INV        m062(.A(mai_mai_n82_), .Y(mai_mai_n85_));
  NO2        m063(.A(x06), .B(x05), .Y(mai_mai_n86_));
  NA2        m064(.A(x11), .B(x00), .Y(mai_mai_n87_));
  NO2        m065(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n88_));
  NOi21      m066(.An(mai_mai_n87_), .B(mai_mai_n88_), .Y(mai_mai_n89_));
  AOI210     m067(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NOi21      m068(.An(x01), .B(x10), .Y(mai_mai_n91_));
  NO2        m069(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n92_));
  NO3        m070(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(x06), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n93_), .B(mai_mai_n27_), .Y(mai_mai_n94_));
  OAI210     m072(.A0(mai_mai_n90_), .A1(x07), .B0(mai_mai_n94_), .Y(mai_mai_n95_));
  NO3        m073(.A(mai_mai_n95_), .B(mai_mai_n84_), .C(mai_mai_n70_), .Y(mai01));
  INV        m074(.A(x12), .Y(mai_mai_n97_));
  INV        m075(.A(x13), .Y(mai_mai_n98_));
  NA2        m076(.A(x08), .B(x04), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n91_), .B(mai_mai_n28_), .Y(mai_mai_n100_));
  NO2        m078(.A(x10), .B(x01), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n343_), .B(mai_mai_n36_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n106_));
  INV        m084(.A(mai_mai_n72_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n108_));
  NA2        m086(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n109_));
  NA2        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NA2        m088(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n112_));
  NO2        m090(.A(x06), .B(x03), .Y(mai_mai_n113_));
  NO3        m091(.A(mai_mai_n113_), .B(mai_mai_n107_), .C(mai_mai_n104_), .Y(mai_mai_n114_));
  NA2        m092(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n115_));
  OAI210     m093(.A0(mai_mai_n81_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n119_));
  AOI210     m097(.A0(mai_mai_n119_), .A1(mai_mai_n49_), .B0(mai_mai_n118_), .Y(mai_mai_n120_));
  AN2        m098(.A(mai_mai_n120_), .B(mai_mai_n117_), .Y(mai_mai_n121_));
  NO2        m099(.A(x09), .B(x05), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n122_), .B(mai_mai_n47_), .Y(mai_mai_n123_));
  AOI210     m101(.A0(mai_mai_n123_), .A1(mai_mai_n103_), .B0(mai_mai_n49_), .Y(mai_mai_n124_));
  NA2        m102(.A(x09), .B(x00), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n105_), .B(mai_mai_n125_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n75_), .B(mai_mai_n51_), .Y(mai_mai_n127_));
  AOI210     m105(.A0(mai_mai_n127_), .A1(mai_mai_n126_), .B0(mai_mai_n119_), .Y(mai_mai_n128_));
  NO3        m106(.A(mai_mai_n128_), .B(mai_mai_n124_), .C(mai_mai_n121_), .Y(mai_mai_n129_));
  OR2        m107(.A(mai_mai_n129_), .B(x11), .Y(mai_mai_n130_));
  OAI210     m108(.A0(mai_mai_n114_), .A1(mai_mai_n23_), .B0(mai_mai_n130_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n103_), .B(mai_mai_n40_), .Y(mai_mai_n132_));
  NOi21      m110(.An(x01), .B(x13), .Y(mai_mai_n133_));
  INV        m111(.A(mai_mai_n133_), .Y(mai_mai_n134_));
  NO2        m112(.A(mai_mai_n132_), .B(mai_mai_n41_), .Y(mai_mai_n135_));
  NO2        m113(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n98_), .B(x01), .Y(mai_mai_n137_));
  OAI210     m115(.A0(x05), .A1(mai_mai_n98_), .B0(mai_mai_n51_), .Y(mai_mai_n138_));
  AOI210     m116(.A0(mai_mai_n138_), .A1(mai_mai_n136_), .B0(mai_mai_n48_), .Y(mai_mai_n139_));
  AOI210     m117(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n140_));
  OAI210     m118(.A0(mai_mai_n139_), .A1(mai_mai_n135_), .B0(mai_mai_n140_), .Y(mai_mai_n141_));
  NA2        m119(.A(x04), .B(x02), .Y(mai_mai_n142_));
  NA2        m120(.A(x10), .B(x05), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n105_), .B(x08), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n91_), .B(x05), .Y(mai_mai_n145_));
  OAI210     m123(.A0(mai_mai_n145_), .A1(x08), .B0(x13), .Y(mai_mai_n146_));
  AOI210     m124(.A0(mai_mai_n144_), .A1(x06), .B0(mai_mai_n146_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n147_), .B(x11), .Y(mai_mai_n148_));
  NAi21      m126(.An(mai_mai_n142_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  INV        m127(.A(mai_mai_n25_), .Y(mai_mai_n150_));
  NAi21      m128(.An(x13), .B(x00), .Y(mai_mai_n151_));
  AOI210     m129(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  AN2        m130(.A(x04), .B(mai_mai_n152_), .Y(mai_mai_n153_));
  INV        m131(.A(x06), .Y(mai_mai_n154_));
  NO2        m132(.A(mai_mai_n151_), .B(mai_mai_n36_), .Y(mai_mai_n155_));
  OAI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n153_), .B0(mai_mai_n150_), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n80_), .B(mai_mai_n47_), .Y(mai_mai_n157_));
  NA2        m135(.A(mai_mai_n157_), .B(mai_mai_n109_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n97_), .B(mai_mai_n158_), .Y(mai_mai_n159_));
  NO2        m137(.A(mai_mai_n98_), .B(x12), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n161_), .B(mai_mai_n159_), .Y(mai_mai_n163_));
  NA4        m141(.A(mai_mai_n163_), .B(mai_mai_n156_), .C(mai_mai_n149_), .D(mai_mai_n141_), .Y(mai_mai_n164_));
  AOI210     m142(.A0(mai_mai_n131_), .A1(mai_mai_n97_), .B0(mai_mai_n164_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n166_), .B(mai_mai_n116_), .Y(mai_mai_n167_));
  AOI210     m145(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n168_));
  NO2        m146(.A(mai_mai_n108_), .B(x06), .Y(mai_mai_n169_));
  AOI210     m147(.A0(mai_mai_n168_), .A1(mai_mai_n167_), .B0(mai_mai_n169_), .Y(mai_mai_n170_));
  AOI210     m148(.A0(mai_mai_n170_), .A1(mai_mai_n73_), .B0(x12), .Y(mai_mai_n171_));
  INV        m149(.A(mai_mai_n75_), .Y(mai_mai_n172_));
  NA2        m150(.A(mai_mai_n134_), .B(mai_mai_n57_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  AOI210     m152(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n175_));
  NA2        m153(.A(mai_mai_n56_), .B(x02), .Y(mai_mai_n176_));
  AOI210     m154(.A0(mai_mai_n176_), .A1(mai_mai_n174_), .B0(mai_mai_n23_), .Y(mai_mai_n177_));
  OAI210     m155(.A0(mai_mai_n171_), .A1(mai_mai_n57_), .B0(mai_mai_n177_), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n119_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n98_), .B(x03), .Y(mai_mai_n181_));
  NO2        m159(.A(mai_mai_n75_), .B(mai_mai_n181_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n182_), .B(mai_mai_n179_), .Y(mai_mai_n183_));
  INV        m161(.A(mai_mai_n88_), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n184_), .B(x12), .Y(mai_mai_n185_));
  NA2        m163(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n186_));
  OAI210     m164(.A0(x08), .A1(x04), .B0(mai_mai_n152_), .Y(mai_mai_n187_));
  AOI210     m165(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n188_), .B(mai_mai_n41_), .Y(mai_mai_n189_));
  OAI210     m167(.A0(mai_mai_n99_), .A1(mai_mai_n125_), .B0(mai_mai_n72_), .Y(mai_mai_n190_));
  NO2        m168(.A(mai_mai_n190_), .B(mai_mai_n189_), .Y(mai_mai_n191_));
  NA2        m169(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n192_));
  INV        m170(.A(x03), .Y(mai_mai_n193_));
  OA210      m171(.A0(mai_mai_n193_), .A1(mai_mai_n191_), .B0(mai_mai_n187_), .Y(mai_mai_n194_));
  NA2        m172(.A(x13), .B(mai_mai_n97_), .Y(mai_mai_n195_));
  NA3        m173(.A(mai_mai_n195_), .B(x12), .C(mai_mai_n89_), .Y(mai_mai_n196_));
  OAI210     m174(.A0(mai_mai_n194_), .A1(mai_mai_n186_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  AOI210     m175(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(mai_mai_n197_), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n198_), .A1(mai_mai_n178_), .B0(x07), .Y(mai_mai_n199_));
  NA2        m177(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n200_));
  AOI210     m178(.A0(mai_mai_n115_), .A1(mai_mai_n127_), .B0(mai_mai_n200_), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n98_), .B(x06), .Y(mai_mai_n202_));
  INV        m180(.A(mai_mai_n202_), .Y(mai_mai_n203_));
  NO2        m181(.A(x08), .B(x05), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(mai_mai_n188_), .Y(mai_mai_n205_));
  OAI210     m183(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n206_));
  OAI210     m184(.A0(mai_mai_n205_), .A1(mai_mai_n203_), .B0(mai_mai_n206_), .Y(mai_mai_n207_));
  NO2        m185(.A(x12), .B(x02), .Y(mai_mai_n208_));
  INV        m186(.A(mai_mai_n208_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n209_), .B(mai_mai_n184_), .Y(mai_mai_n210_));
  OA210      m188(.A0(mai_mai_n207_), .A1(mai_mai_n201_), .B0(mai_mai_n210_), .Y(mai_mai_n211_));
  NO2        m189(.A(x05), .B(x01), .Y(mai_mai_n212_));
  NA2        m190(.A(mai_mai_n98_), .B(x04), .Y(mai_mai_n213_));
  NA2        m191(.A(x02), .B(x06), .Y(mai_mai_n214_));
  NO3        m192(.A(mai_mai_n87_), .B(x12), .C(x03), .Y(mai_mai_n215_));
  OAI210     m193(.A0(mai_mai_n214_), .A1(x10), .B0(mai_mai_n215_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n340_), .B(mai_mai_n217_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n219_));
  NO3        m197(.A(mai_mai_n219_), .B(mai_mai_n175_), .C(mai_mai_n154_), .Y(mai_mai_n220_));
  NO2        m198(.A(mai_mai_n186_), .B(mai_mai_n28_), .Y(mai_mai_n221_));
  NA2        m199(.A(mai_mai_n220_), .B(mai_mai_n221_), .Y(mai_mai_n222_));
  NA3        m200(.A(mai_mai_n222_), .B(mai_mai_n218_), .C(mai_mai_n216_), .Y(mai_mai_n223_));
  NO3        m201(.A(mai_mai_n223_), .B(mai_mai_n211_), .C(mai_mai_n199_), .Y(mai_mai_n224_));
  OAI210     m202(.A0(mai_mai_n165_), .A1(mai_mai_n61_), .B0(mai_mai_n224_), .Y(mai02));
  AOI210     m203(.A0(mai_mai_n115_), .A1(mai_mai_n82_), .B0(mai_mai_n111_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n98_), .B(mai_mai_n35_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n32_), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n143_), .Y(mai_mai_n229_));
  INV        m207(.A(mai_mai_n143_), .Y(mai_mai_n230_));
  NA2        m208(.A(x09), .B(mai_mai_n230_), .Y(mai_mai_n231_));
  AOI210     m209(.A0(mai_mai_n231_), .A1(mai_mai_n229_), .B0(mai_mai_n48_), .Y(mai_mai_n232_));
  NO2        m210(.A(x05), .B(x02), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n167_), .B(mai_mai_n233_), .Y(mai_mai_n234_));
  AOI220     m212(.A0(mai_mai_n204_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n235_));
  NOi21      m213(.An(mai_mai_n227_), .B(mai_mai_n235_), .Y(mai_mai_n236_));
  AOI210     m214(.A0(x13), .A1(mai_mai_n77_), .B0(mai_mai_n236_), .Y(mai_mai_n237_));
  AOI210     m215(.A0(mai_mai_n237_), .A1(mai_mai_n234_), .B0(mai_mai_n119_), .Y(mai_mai_n238_));
  INV        m216(.A(mai_mai_n182_), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n192_), .B(mai_mai_n47_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n240_), .B(mai_mai_n239_), .Y(mai_mai_n241_));
  OAI210     m219(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n242_));
  OA210      m220(.A0(mai_mai_n344_), .A1(x08), .B0(mai_mai_n123_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n243_), .A1(mai_mai_n116_), .B0(mai_mai_n242_), .Y(mai_mai_n244_));
  OAI210     m222(.A0(mai_mai_n244_), .A1(mai_mai_n181_), .B0(mai_mai_n92_), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n92_), .B(mai_mai_n180_), .Y(mai_mai_n246_));
  NA3        m224(.A(mai_mai_n91_), .B(mai_mai_n80_), .C(mai_mai_n42_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n247_), .A1(mai_mai_n246_), .B0(x04), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n205_), .B(mai_mai_n100_), .Y(mai_mai_n249_));
  AOI210     m227(.A0(mai_mai_n249_), .A1(x13), .B0(mai_mai_n248_), .Y(mai_mai_n250_));
  NA3        m228(.A(mai_mai_n250_), .B(mai_mai_n245_), .C(mai_mai_n241_), .Y(mai_mai_n251_));
  NO3        m229(.A(mai_mai_n251_), .B(mai_mai_n238_), .C(mai_mai_n232_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n118_), .B(x03), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n162_), .B(mai_mai_n101_), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n142_), .B(mai_mai_n137_), .Y(mai_mai_n255_));
  AN2        m233(.A(mai_mai_n255_), .B(mai_mai_n144_), .Y(mai_mai_n256_));
  OAI220     m234(.A0(mai_mai_n213_), .A1(x09), .B0(mai_mai_n111_), .B1(mai_mai_n28_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n257_), .A1(mai_mai_n256_), .B0(mai_mai_n102_), .Y(mai_mai_n258_));
  NA2        m236(.A(mai_mai_n213_), .B(mai_mai_n97_), .Y(mai_mai_n259_));
  NA2        m237(.A(mai_mai_n259_), .B(mai_mai_n110_), .Y(mai_mai_n260_));
  NA4        m238(.A(mai_mai_n260_), .B(mai_mai_n258_), .C(mai_mai_n254_), .D(mai_mai_n48_), .Y(mai_mai_n261_));
  INV        m239(.A(mai_mai_n162_), .Y(mai_mai_n262_));
  OAI220     m240(.A0(mai_mai_n339_), .A1(mai_mai_n31_), .B0(mai_mai_n262_), .B1(mai_mai_n59_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n263_), .B(x02), .Y(mai_mai_n264_));
  INV        m242(.A(x08), .Y(mai_mai_n265_));
  NA2        m243(.A(mai_mai_n160_), .B(x04), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n266_), .B(mai_mai_n265_), .Y(mai_mai_n267_));
  NO2        m245(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n268_));
  OAI210     m246(.A0(mai_mai_n268_), .A1(mai_mai_n267_), .B0(mai_mai_n92_), .Y(mai_mai_n269_));
  NO3        m247(.A(mai_mai_n160_), .B(mai_mai_n136_), .C(mai_mai_n52_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(x12), .A1(mai_mai_n157_), .B0(mai_mai_n270_), .Y(mai_mai_n271_));
  NA4        m249(.A(mai_mai_n271_), .B(mai_mai_n269_), .C(mai_mai_n264_), .D(x06), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n166_), .B(mai_mai_n64_), .Y(mai_mai_n273_));
  NO3        m251(.A(mai_mai_n219_), .B(mai_mai_n108_), .C(x08), .Y(mai_mai_n274_));
  INV        m252(.A(mai_mai_n274_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n270_), .B(x06), .Y(mai_mai_n276_));
  OAI210     m254(.A0(mai_mai_n275_), .A1(mai_mai_n28_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  AO220      m255(.A0(mai_mai_n277_), .A1(x04), .B0(mai_mai_n273_), .B1(x05), .Y(mai_mai_n278_));
  AOI210     m256(.A0(mai_mai_n272_), .A1(mai_mai_n261_), .B0(mai_mai_n278_), .Y(mai_mai_n279_));
  OAI210     m257(.A0(mai_mai_n252_), .A1(x12), .B0(mai_mai_n279_), .Y(mai03));
  OR2        m258(.A(mai_mai_n42_), .B(mai_mai_n180_), .Y(mai_mai_n281_));
  AOI210     m259(.A0(x13), .A1(mai_mai_n97_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n341_), .A1(mai_mai_n282_), .B0(x05), .Y(mai_mai_n283_));
  NA2        m261(.A(mai_mai_n281_), .B(x05), .Y(mai_mai_n284_));
  AOI210     m262(.A0(mai_mai_n116_), .A1(mai_mai_n172_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  OAI220     m263(.A0(mai_mai_n342_), .A1(mai_mai_n59_), .B0(mai_mai_n344_), .B1(mai_mai_n235_), .Y(mai_mai_n286_));
  OAI210     m264(.A0(mai_mai_n286_), .A1(mai_mai_n285_), .B0(mai_mai_n97_), .Y(mai_mai_n287_));
  INV        m265(.A(mai_mai_n126_), .Y(mai_mai_n288_));
  NA2        m266(.A(mai_mai_n288_), .B(x04), .Y(mai_mai_n289_));
  NO3        m267(.A(x12), .B(mai_mai_n82_), .C(mai_mai_n59_), .Y(mai_mai_n290_));
  NO2        m268(.A(mai_mai_n97_), .B(mai_mai_n123_), .Y(mai_mai_n291_));
  OA210      m269(.A0(mai_mai_n98_), .A1(x12), .B0(mai_mai_n112_), .Y(mai_mai_n292_));
  NO3        m270(.A(mai_mai_n292_), .B(mai_mai_n291_), .C(mai_mai_n290_), .Y(mai_mai_n293_));
  NA4        m271(.A(mai_mai_n293_), .B(mai_mai_n289_), .C(mai_mai_n287_), .D(mai_mai_n283_), .Y(mai04));
  NO2        m272(.A(mai_mai_n85_), .B(mai_mai_n39_), .Y(mai_mai_n295_));
  XO2        m273(.A(mai_mai_n295_), .B(mai_mai_n195_), .Y(mai05));
  NA2        m274(.A(mai_mai_n71_), .B(mai_mai_n52_), .Y(mai_mai_n297_));
  AOI210     m275(.A0(mai_mai_n297_), .A1(mai_mai_n242_), .B0(mai_mai_n25_), .Y(mai_mai_n298_));
  NA3        m276(.A(mai_mai_n119_), .B(mai_mai_n111_), .C(mai_mai_n31_), .Y(mai_mai_n299_));
  INV        m277(.A(mai_mai_n86_), .Y(mai_mai_n300_));
  AOI210     m278(.A0(mai_mai_n300_), .A1(mai_mai_n299_), .B0(mai_mai_n24_), .Y(mai_mai_n301_));
  OAI210     m279(.A0(mai_mai_n301_), .A1(mai_mai_n298_), .B0(mai_mai_n97_), .Y(mai_mai_n302_));
  NA2        m280(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n303_));
  NA2        m281(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n304_));
  NA2        m282(.A(mai_mai_n200_), .B(x03), .Y(mai_mai_n305_));
  OAI220     m283(.A0(mai_mai_n305_), .A1(mai_mai_n304_), .B0(mai_mai_n303_), .B1(mai_mai_n78_), .Y(mai_mai_n306_));
  OAI210     m284(.A0(mai_mai_n26_), .A1(mai_mai_n97_), .B0(x07), .Y(mai_mai_n307_));
  AOI210     m285(.A0(mai_mai_n306_), .A1(x06), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  NA2        m286(.A(mai_mai_n33_), .B(mai_mai_n97_), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n309_), .A1(mai_mai_n88_), .B0(x07), .Y(mai_mai_n310_));
  AOI210     m288(.A0(mai_mai_n308_), .A1(mai_mai_n302_), .B0(mai_mai_n310_), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n118_), .Y(mai_mai_n312_));
  OR2        m290(.A(mai_mai_n312_), .B(x03), .Y(mai_mai_n313_));
  NO2        m291(.A(mai_mai_n122_), .B(mai_mai_n28_), .Y(mai_mai_n314_));
  AOI210     m292(.A0(mai_mai_n314_), .A1(mai_mai_n313_), .B0(mai_mai_n47_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n315_), .B(mai_mai_n98_), .Y(mai_mai_n316_));
  NOi21      m294(.An(mai_mai_n253_), .B(mai_mai_n112_), .Y(mai_mai_n317_));
  NO2        m295(.A(mai_mai_n317_), .B(mai_mai_n209_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n319_));
  AOI210     m297(.A0(mai_mai_n195_), .A1(mai_mai_n47_), .B0(mai_mai_n319_), .Y(mai_mai_n320_));
  NO3        m298(.A(mai_mai_n320_), .B(mai_mai_n318_), .C(x08), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n111_), .B(mai_mai_n28_), .Y(mai_mai_n322_));
  NO2        m300(.A(mai_mai_n322_), .B(mai_mai_n212_), .Y(mai_mai_n323_));
  NA3        m301(.A(mai_mai_n262_), .B(mai_mai_n106_), .C(x12), .Y(mai_mai_n324_));
  AO210      m302(.A0(mai_mai_n262_), .A1(mai_mai_n106_), .B0(mai_mai_n195_), .Y(mai_mai_n325_));
  NA3        m303(.A(mai_mai_n325_), .B(mai_mai_n324_), .C(x08), .Y(mai_mai_n326_));
  INV        m304(.A(mai_mai_n326_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n316_), .B0(mai_mai_n327_), .Y(mai_mai_n328_));
  NA3        m306(.A(mai_mai_n323_), .B(mai_mai_n317_), .C(mai_mai_n259_), .Y(mai_mai_n329_));
  NA2        m307(.A(x14), .B(mai_mai_n329_), .Y(mai_mai_n330_));
  NA2        m308(.A(mai_mai_n309_), .B(mai_mai_n61_), .Y(mai_mai_n331_));
  NOi21      m309(.An(mai_mai_n213_), .B(mai_mai_n126_), .Y(mai_mai_n332_));
  NA2        m310(.A(mai_mai_n332_), .B(mai_mai_n97_), .Y(mai_mai_n333_));
  OAI210     m311(.A0(mai_mai_n331_), .A1(mai_mai_n87_), .B0(mai_mai_n333_), .Y(mai_mai_n334_));
  NO4        m312(.A(mai_mai_n334_), .B(mai_mai_n330_), .C(mai_mai_n328_), .D(mai_mai_n311_), .Y(mai06));
  INV        m313(.A(x07), .Y(mai_mai_n338_));
  INV        m314(.A(x05), .Y(mai_mai_n339_));
  INV        m315(.A(mai_mai_n99_), .Y(mai_mai_n340_));
  INV        m316(.A(mai_mai_n266_), .Y(mai_mai_n341_));
  INV        m317(.A(mai_mai_n181_), .Y(mai_mai_n342_));
  INV        m318(.A(x04), .Y(mai_mai_n343_));
  INV        m319(.A(x13), .Y(mai_mai_n344_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  INV        u007(.A(x03), .Y(men_men_n30_));
  NA2        u008(.A(x10), .B(men_men_n30_), .Y(men_men_n31_));
  NA3        u009(.A(men_men_n31_), .B(x02), .C(x06), .Y(men_men_n32_));
  NA2        u010(.A(men_men_n32_), .B(men_men_n27_), .Y(men_men_n33_));
  INV        u011(.A(x04), .Y(men_men_n34_));
  INV        u012(.A(x08), .Y(men_men_n35_));
  NA2        u013(.A(men_men_n35_), .B(x02), .Y(men_men_n36_));
  NA2        u014(.A(x08), .B(x03), .Y(men_men_n37_));
  AOI210     u015(.A0(men_men_n37_), .A1(men_men_n36_), .B0(men_men_n34_), .Y(men_men_n38_));
  NA2        u016(.A(x09), .B(men_men_n30_), .Y(men_men_n39_));
  INV        u017(.A(x05), .Y(men_men_n40_));
  NO2        u018(.A(x09), .B(x02), .Y(men_men_n41_));
  NO2        u019(.A(men_men_n41_), .B(men_men_n40_), .Y(men_men_n42_));
  NA2        u020(.A(men_men_n42_), .B(men_men_n39_), .Y(men_men_n43_));
  INV        u021(.A(men_men_n43_), .Y(men_men_n44_));
  NO3        u022(.A(men_men_n44_), .B(men_men_n38_), .C(men_men_n33_), .Y(men00));
  INV        u023(.A(x01), .Y(men_men_n46_));
  INV        u024(.A(x06), .Y(men_men_n47_));
  NO2        u025(.A(x02), .B(x11), .Y(men_men_n48_));
  INV        u026(.A(x09), .Y(men_men_n49_));
  NO2        u027(.A(x10), .B(x02), .Y(men_men_n50_));
  NO2        u028(.A(x09), .B(x07), .Y(men_men_n51_));
  OAI210     u029(.A0(men_men_n51_), .A1(men_men_n48_), .B0(men_men_n46_), .Y(men_men_n52_));
  NOi21      u030(.An(x01), .B(x09), .Y(men_men_n53_));
  INV        u031(.A(x00), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n49_), .B(men_men_n54_), .Y(men_men_n55_));
  NO2        u033(.A(men_men_n55_), .B(men_men_n53_), .Y(men_men_n56_));
  NA2        u034(.A(x09), .B(men_men_n54_), .Y(men_men_n57_));
  INV        u035(.A(x07), .Y(men_men_n58_));
  NA2        u036(.A(men_men_n56_), .B(men_men_n30_), .Y(men_men_n59_));
  AOI210     u037(.A0(men_men_n59_), .A1(men_men_n52_), .B0(x05), .Y(men_men_n60_));
  NA2        u038(.A(x10), .B(x09), .Y(men_men_n61_));
  NA2        u039(.A(x09), .B(x05), .Y(men_men_n62_));
  NA2        u040(.A(x10), .B(x06), .Y(men_men_n63_));
  NO2        u041(.A(men_men_n58_), .B(men_men_n40_), .Y(men_men_n64_));
  NA2        u042(.A(x07), .B(x03), .Y(men_men_n65_));
  NOi31      u043(.An(x08), .B(x04), .C(x00), .Y(men_men_n66_));
  NO2        u044(.A(x09), .B(men_men_n40_), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n67_), .B(men_men_n35_), .Y(men_men_n68_));
  OAI210     u046(.A0(men_men_n67_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n69_));
  AOI210     u047(.A0(men_men_n68_), .A1(men_men_n47_), .B0(men_men_n69_), .Y(men_men_n70_));
  NO2        u048(.A(men_men_n35_), .B(x00), .Y(men_men_n71_));
  NO2        u049(.A(x08), .B(x01), .Y(men_men_n72_));
  OAI210     u050(.A0(men_men_n72_), .A1(men_men_n71_), .B0(men_men_n34_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n73_), .B(men_men_n70_), .Y(men_men_n74_));
  AN2        u052(.A(men_men_n74_), .B(men_men_n65_), .Y(men_men_n75_));
  INV        u053(.A(men_men_n73_), .Y(men_men_n76_));
  NO2        u054(.A(x06), .B(x05), .Y(men_men_n77_));
  NA2        u055(.A(x11), .B(x00), .Y(men_men_n78_));
  NO2        u056(.A(x11), .B(men_men_n46_), .Y(men_men_n79_));
  NOi21      u057(.An(men_men_n78_), .B(men_men_n79_), .Y(men_men_n80_));
  NOi21      u058(.An(x01), .B(x10), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n29_), .B(men_men_n54_), .Y(men_men_n82_));
  NO3        u060(.A(men_men_n82_), .B(men_men_n81_), .C(x06), .Y(men_men_n83_));
  NA2        u061(.A(men_men_n83_), .B(men_men_n27_), .Y(men_men_n84_));
  OAI210     u062(.A0(men_men_n422_), .A1(x07), .B0(men_men_n84_), .Y(men_men_n85_));
  NO3        u063(.A(men_men_n85_), .B(men_men_n75_), .C(men_men_n60_), .Y(men01));
  INV        u064(.A(x12), .Y(men_men_n87_));
  INV        u065(.A(x13), .Y(men_men_n88_));
  NA2        u066(.A(x08), .B(x04), .Y(men_men_n89_));
  NA2        u067(.A(men_men_n81_), .B(men_men_n28_), .Y(men_men_n90_));
  NO2        u068(.A(men_men_n90_), .B(men_men_n62_), .Y(men_men_n91_));
  NO2        u069(.A(x10), .B(x01), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n29_), .B(x00), .Y(men_men_n93_));
  NO2        u071(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NA2        u072(.A(x04), .B(men_men_n28_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n35_), .C(men_men_n40_), .Y(men_men_n96_));
  AOI210     u074(.A0(men_men_n96_), .A1(men_men_n94_), .B0(men_men_n91_), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n97_), .B(men_men_n88_), .Y(men_men_n98_));
  NO2        u076(.A(men_men_n53_), .B(x05), .Y(men_men_n99_));
  NOi21      u077(.An(men_men_n99_), .B(men_men_n55_), .Y(men_men_n100_));
  NO2        u078(.A(men_men_n34_), .B(x02), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n88_), .B(men_men_n35_), .Y(men_men_n102_));
  NA3        u080(.A(men_men_n102_), .B(men_men_n101_), .C(x06), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n103_), .B(men_men_n100_), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n72_), .B(x13), .Y(men_men_n105_));
  NA2        u083(.A(x09), .B(men_men_n34_), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NA2        u085(.A(x13), .B(men_men_n34_), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n108_), .B(x05), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n107_), .Y(men_men_n110_));
  NA2        u088(.A(men_men_n34_), .B(men_men_n54_), .Y(men_men_n111_));
  NA2        u089(.A(men_men_n111_), .B(men_men_n88_), .Y(men_men_n112_));
  AOI210     u090(.A0(men_men_n112_), .A1(men_men_n68_), .B0(men_men_n100_), .Y(men_men_n113_));
  AOI210     u091(.A0(men_men_n113_), .A1(men_men_n110_), .B0(men_men_n63_), .Y(men_men_n114_));
  NA2        u092(.A(men_men_n29_), .B(men_men_n46_), .Y(men_men_n115_));
  NA2        u093(.A(x10), .B(men_men_n54_), .Y(men_men_n116_));
  NA2        u094(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n49_), .B(x05), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n35_), .B(x04), .Y(men_men_n119_));
  NA3        u097(.A(men_men_n119_), .B(men_men_n118_), .C(x13), .Y(men_men_n120_));
  NO3        u098(.A(men_men_n111_), .B(men_men_n67_), .C(men_men_n35_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n57_), .B(x05), .Y(men_men_n122_));
  NOi41      u100(.An(men_men_n120_), .B(men_men_n122_), .C(men_men_n121_), .D(men_men_n117_), .Y(men_men_n123_));
  NO3        u101(.A(men_men_n123_), .B(x06), .C(x03), .Y(men_men_n124_));
  NO4        u102(.A(men_men_n124_), .B(men_men_n114_), .C(men_men_n104_), .D(men_men_n98_), .Y(men_men_n125_));
  NA2        u103(.A(x13), .B(men_men_n35_), .Y(men_men_n126_));
  OAI210     u104(.A0(men_men_n72_), .A1(x13), .B0(men_men_n34_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n127_), .B(men_men_n126_), .Y(men_men_n128_));
  NO2        u106(.A(men_men_n49_), .B(men_men_n40_), .Y(men_men_n129_));
  NA2        u107(.A(men_men_n29_), .B(x06), .Y(men_men_n130_));
  OA210      u108(.A0(men_men_n28_), .A1(x04), .B0(men_men_n128_), .Y(men_men_n131_));
  NO2        u109(.A(x09), .B(x05), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n132_), .B(men_men_n46_), .Y(men_men_n133_));
  NA2        u111(.A(x09), .B(x00), .Y(men_men_n134_));
  INV        u112(.A(men_men_n130_), .Y(men_men_n135_));
  NO3        u113(.A(men_men_n135_), .B(men_men_n424_), .C(men_men_n131_), .Y(men_men_n136_));
  NO2        u114(.A(x03), .B(x02), .Y(men_men_n137_));
  NA2        u115(.A(men_men_n73_), .B(men_men_n88_), .Y(men_men_n138_));
  OAI210     u116(.A0(men_men_n138_), .A1(men_men_n100_), .B0(men_men_n137_), .Y(men_men_n139_));
  OA210      u117(.A0(men_men_n136_), .A1(x11), .B0(men_men_n139_), .Y(men_men_n140_));
  OAI210     u118(.A0(men_men_n125_), .A1(men_men_n23_), .B0(men_men_n140_), .Y(men_men_n141_));
  NA2        u119(.A(men_men_n94_), .B(men_men_n39_), .Y(men_men_n142_));
  NAi21      u120(.An(x06), .B(x10), .Y(men_men_n143_));
  NOi21      u121(.An(x01), .B(x13), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n145_));
  OR2        u123(.A(men_men_n145_), .B(x08), .Y(men_men_n146_));
  AOI210     u124(.A0(men_men_n146_), .A1(men_men_n142_), .B0(men_men_n40_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n29_), .B(x03), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n88_), .B(x01), .Y(men_men_n149_));
  NO2        u127(.A(men_men_n149_), .B(x08), .Y(men_men_n150_));
  OAI210     u128(.A0(x05), .A1(men_men_n150_), .B0(men_men_n49_), .Y(men_men_n151_));
  AOI210     u129(.A0(men_men_n151_), .A1(men_men_n148_), .B0(men_men_n47_), .Y(men_men_n152_));
  AOI210     u130(.A0(x11), .A1(men_men_n30_), .B0(men_men_n28_), .Y(men_men_n153_));
  OAI210     u131(.A0(men_men_n152_), .A1(men_men_n147_), .B0(men_men_n153_), .Y(men_men_n154_));
  NA2        u132(.A(x04), .B(x02), .Y(men_men_n155_));
  NA2        u133(.A(x10), .B(x05), .Y(men_men_n156_));
  NA2        u134(.A(x09), .B(x06), .Y(men_men_n157_));
  NO2        u135(.A(x09), .B(x01), .Y(men_men_n158_));
  NO3        u136(.A(men_men_n158_), .B(men_men_n92_), .C(men_men_n30_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n159_), .B(x00), .Y(men_men_n160_));
  NA3        u138(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n49_), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n81_), .B(x05), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n162_), .A1(men_men_n102_), .B0(men_men_n161_), .Y(men_men_n163_));
  INV        u141(.A(men_men_n163_), .Y(men_men_n164_));
  OAI210     u142(.A0(men_men_n164_), .A1(x11), .B0(men_men_n160_), .Y(men_men_n165_));
  NAi21      u143(.An(men_men_n155_), .B(men_men_n165_), .Y(men_men_n166_));
  NAi21      u144(.An(x13), .B(x00), .Y(men_men_n167_));
  AOI210     u145(.A0(men_men_n29_), .A1(men_men_n47_), .B0(men_men_n167_), .Y(men_men_n168_));
  AOI220     u146(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n169_));
  OAI210     u147(.A0(men_men_n156_), .A1(men_men_n34_), .B0(men_men_n169_), .Y(men_men_n170_));
  AN2        u148(.A(men_men_n170_), .B(men_men_n168_), .Y(men_men_n171_));
  NO2        u149(.A(men_men_n82_), .B(x06), .Y(men_men_n172_));
  NO2        u150(.A(men_men_n167_), .B(men_men_n35_), .Y(men_men_n173_));
  INV        u151(.A(men_men_n173_), .Y(men_men_n174_));
  OAI220     u152(.A0(men_men_n174_), .A1(men_men_n157_), .B0(men_men_n172_), .B1(men_men_n62_), .Y(men_men_n175_));
  OAI210     u153(.A0(men_men_n175_), .A1(men_men_n171_), .B0(x03), .Y(men_men_n176_));
  NOi21      u154(.An(x09), .B(x00), .Y(men_men_n177_));
  NA2        u155(.A(x10), .B(x08), .Y(men_men_n178_));
  INV        u156(.A(men_men_n178_), .Y(men_men_n179_));
  NA2        u157(.A(x06), .B(x05), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(men_men_n34_), .B0(men_men_n87_), .Y(men_men_n181_));
  AOI210     u159(.A0(men_men_n179_), .A1(men_men_n55_), .B0(men_men_n181_), .Y(men_men_n182_));
  INV        u160(.A(men_men_n182_), .Y(men_men_n183_));
  NO2        u161(.A(men_men_n88_), .B(x12), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n184_), .Y(men_men_n185_));
  NA2        u163(.A(men_men_n81_), .B(men_men_n49_), .Y(men_men_n186_));
  NO2        u164(.A(men_men_n34_), .B(men_men_n30_), .Y(men_men_n187_));
  NA2        u165(.A(men_men_n187_), .B(x02), .Y(men_men_n188_));
  NO2        u166(.A(men_men_n188_), .B(men_men_n186_), .Y(men_men_n189_));
  AOI210     u167(.A0(men_men_n185_), .A1(men_men_n183_), .B0(men_men_n189_), .Y(men_men_n190_));
  NA4        u168(.A(men_men_n190_), .B(men_men_n176_), .C(men_men_n166_), .D(men_men_n154_), .Y(men_men_n191_));
  AOI210     u169(.A0(men_men_n141_), .A1(men_men_n87_), .B0(men_men_n191_), .Y(men_men_n192_));
  NA2        u170(.A(men_men_n28_), .B(men_men_n128_), .Y(men_men_n193_));
  NA2        u171(.A(men_men_n49_), .B(men_men_n46_), .Y(men_men_n194_));
  NA2        u172(.A(men_men_n194_), .B(men_men_n127_), .Y(men_men_n195_));
  NO2        u173(.A(men_men_n115_), .B(x06), .Y(men_men_n196_));
  AOI210     u174(.A0(men_men_n423_), .A1(men_men_n195_), .B0(men_men_n196_), .Y(men_men_n197_));
  AOI210     u175(.A0(men_men_n197_), .A1(men_men_n193_), .B0(x12), .Y(men_men_n198_));
  INV        u176(.A(men_men_n66_), .Y(men_men_n199_));
  AOI210     u177(.A0(men_men_n178_), .A1(x05), .B0(men_men_n49_), .Y(men_men_n200_));
  OAI210     u178(.A0(men_men_n200_), .A1(men_men_n145_), .B0(men_men_n54_), .Y(men_men_n201_));
  NA2        u179(.A(men_men_n201_), .B(men_men_n199_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n81_), .B(x06), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n35_), .A1(x04), .B0(men_men_n49_), .Y(men_men_n204_));
  NO3        u182(.A(men_men_n204_), .B(men_men_n203_), .C(men_men_n40_), .Y(men_men_n205_));
  NA4        u183(.A(men_men_n143_), .B(men_men_n53_), .C(men_men_n35_), .D(x04), .Y(men_men_n206_));
  NA2        u184(.A(men_men_n206_), .B(men_men_n130_), .Y(men_men_n207_));
  OAI210     u185(.A0(men_men_n207_), .A1(men_men_n205_), .B0(x02), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n208_), .A1(men_men_n202_), .B0(men_men_n23_), .Y(men_men_n209_));
  OAI210     u187(.A0(men_men_n198_), .A1(men_men_n54_), .B0(men_men_n209_), .Y(men_men_n210_));
  INV        u188(.A(men_men_n130_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n49_), .B(x03), .Y(men_men_n212_));
  OAI210     u190(.A0(men_men_n67_), .A1(men_men_n35_), .B0(men_men_n106_), .Y(men_men_n213_));
  NO2        u191(.A(men_men_n88_), .B(x03), .Y(men_men_n214_));
  AOI220     u192(.A0(men_men_n214_), .A1(men_men_n213_), .B0(men_men_n66_), .B1(men_men_n212_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n31_), .B(x06), .Y(men_men_n216_));
  INV        u194(.A(men_men_n143_), .Y(men_men_n217_));
  NOi21      u195(.An(x13), .B(x04), .Y(men_men_n218_));
  NO3        u196(.A(men_men_n218_), .B(men_men_n66_), .C(men_men_n177_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n219_), .B(x05), .Y(men_men_n220_));
  AOI220     u198(.A0(men_men_n220_), .A1(men_men_n216_), .B0(men_men_n217_), .B1(men_men_n54_), .Y(men_men_n221_));
  NA2        u199(.A(men_men_n215_), .B(men_men_n221_), .Y(men_men_n222_));
  INV        u200(.A(men_men_n79_), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n23_), .B(men_men_n46_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n49_), .B(men_men_n35_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n225_), .A1(men_men_n170_), .B0(men_men_n168_), .Y(men_men_n226_));
  AOI210     u204(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n227_));
  NO2        u205(.A(x06), .B(x00), .Y(men_men_n228_));
  NO3        u206(.A(men_men_n228_), .B(men_men_n227_), .C(men_men_n40_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n89_), .A1(men_men_n134_), .B0(men_men_n63_), .Y(men_men_n230_));
  NO2        u208(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n232_), .B(x03), .Y(men_men_n233_));
  OA210      u211(.A0(men_men_n233_), .A1(men_men_n231_), .B0(men_men_n226_), .Y(men_men_n234_));
  NA2        u212(.A(x13), .B(men_men_n87_), .Y(men_men_n235_));
  NA3        u213(.A(men_men_n235_), .B(men_men_n181_), .C(men_men_n80_), .Y(men_men_n236_));
  OAI210     u214(.A0(men_men_n234_), .A1(men_men_n224_), .B0(men_men_n236_), .Y(men_men_n237_));
  AOI210     u215(.A0(men_men_n79_), .A1(men_men_n222_), .B0(men_men_n237_), .Y(men_men_n238_));
  AOI210     u216(.A0(men_men_n238_), .A1(men_men_n210_), .B0(x07), .Y(men_men_n239_));
  NA2        u217(.A(men_men_n62_), .B(men_men_n29_), .Y(men_men_n240_));
  INV        u218(.A(men_men_n240_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n88_), .B(x06), .Y(men_men_n242_));
  NO2        u220(.A(x08), .B(x05), .Y(men_men_n243_));
  NO2        u221(.A(men_men_n243_), .B(men_men_n227_), .Y(men_men_n244_));
  OAI210     u222(.A0(men_men_n244_), .A1(x06), .B0(x03), .Y(men_men_n245_));
  NO2        u223(.A(x12), .B(x02), .Y(men_men_n246_));
  INV        u224(.A(men_men_n246_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n247_), .B(men_men_n223_), .Y(men_men_n248_));
  OA210      u226(.A0(men_men_n245_), .A1(men_men_n241_), .B0(men_men_n248_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n49_), .B(men_men_n40_), .Y(men_men_n250_));
  NO2        u228(.A(men_men_n250_), .B(x01), .Y(men_men_n251_));
  NOi21      u229(.An(men_men_n72_), .B(men_men_n106_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(men_men_n251_), .Y(men_men_n253_));
  AOI210     u231(.A0(men_men_n253_), .A1(men_men_n120_), .B0(men_men_n29_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n242_), .B(men_men_n213_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n88_), .B(x04), .Y(men_men_n256_));
  INV        u234(.A(men_men_n255_), .Y(men_men_n257_));
  NO3        u235(.A(men_men_n78_), .B(x12), .C(x03), .Y(men_men_n258_));
  OAI210     u236(.A0(men_men_n257_), .A1(men_men_n254_), .B0(men_men_n258_), .Y(men_men_n259_));
  AOI210     u237(.A0(men_men_n186_), .A1(men_men_n180_), .B0(men_men_n89_), .Y(men_men_n260_));
  NOi21      u238(.An(men_men_n240_), .B(men_men_n203_), .Y(men_men_n261_));
  NO2        u239(.A(men_men_n25_), .B(x00), .Y(men_men_n262_));
  OAI210     u240(.A0(men_men_n261_), .A1(men_men_n260_), .B0(men_men_n262_), .Y(men_men_n263_));
  NO2        u241(.A(men_men_n55_), .B(x05), .Y(men_men_n264_));
  NO3        u242(.A(men_men_n264_), .B(men_men_n204_), .C(men_men_n172_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n224_), .B(men_men_n28_), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n265_), .A1(men_men_n211_), .B0(men_men_n266_), .Y(men_men_n267_));
  NA3        u245(.A(men_men_n267_), .B(men_men_n263_), .C(men_men_n259_), .Y(men_men_n268_));
  NO3        u246(.A(men_men_n268_), .B(men_men_n249_), .C(men_men_n239_), .Y(men_men_n269_));
  OAI210     u247(.A0(men_men_n192_), .A1(men_men_n58_), .B0(men_men_n269_), .Y(men02));
  AOI210     u248(.A0(men_men_n126_), .A1(men_men_n73_), .B0(men_men_n118_), .Y(men_men_n271_));
  NOi21      u249(.An(men_men_n219_), .B(men_men_n158_), .Y(men_men_n272_));
  NA3        u250(.A(x13), .B(men_men_n179_), .C(men_men_n53_), .Y(men_men_n273_));
  OAI210     u251(.A0(men_men_n272_), .A1(men_men_n31_), .B0(men_men_n273_), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n274_), .A1(men_men_n271_), .B0(men_men_n156_), .Y(men_men_n275_));
  INV        u253(.A(men_men_n156_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n101_), .B(men_men_n204_), .Y(men_men_n277_));
  OAI220     u255(.A0(men_men_n277_), .A1(men_men_n88_), .B0(men_men_n73_), .B1(men_men_n49_), .Y(men_men_n278_));
  AOI220     u256(.A0(men_men_n278_), .A1(men_men_n276_), .B0(men_men_n138_), .B1(men_men_n137_), .Y(men_men_n279_));
  AOI210     u257(.A0(men_men_n279_), .A1(men_men_n275_), .B0(men_men_n47_), .Y(men_men_n280_));
  NO2        u258(.A(x05), .B(x02), .Y(men_men_n281_));
  OAI210     u259(.A0(men_men_n195_), .A1(men_men_n177_), .B0(men_men_n281_), .Y(men_men_n282_));
  AOI220     u260(.A0(men_men_n243_), .A1(men_men_n55_), .B0(men_men_n53_), .B1(men_men_n35_), .Y(men_men_n283_));
  NOi21      u261(.An(x13), .B(men_men_n283_), .Y(men_men_n284_));
  AOI210     u262(.A0(men_men_n218_), .A1(men_men_n67_), .B0(men_men_n284_), .Y(men_men_n285_));
  AOI210     u263(.A0(men_men_n285_), .A1(men_men_n282_), .B0(men_men_n130_), .Y(men_men_n286_));
  NAi21      u264(.An(men_men_n220_), .B(men_men_n215_), .Y(men_men_n287_));
  NO2        u265(.A(men_men_n232_), .B(men_men_n46_), .Y(men_men_n288_));
  NA2        u266(.A(men_men_n288_), .B(men_men_n287_), .Y(men_men_n289_));
  AN2        u267(.A(men_men_n214_), .B(men_men_n213_), .Y(men_men_n290_));
  OAI210     u268(.A0(men_men_n41_), .A1(men_men_n40_), .B0(men_men_n47_), .Y(men_men_n291_));
  NA2        u269(.A(x13), .B(men_men_n28_), .Y(men_men_n292_));
  AOI210     u270(.A0(men_men_n292_), .A1(men_men_n127_), .B0(men_men_n291_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n293_), .A1(men_men_n290_), .B0(men_men_n82_), .Y(men_men_n294_));
  NA3        u272(.A(men_men_n82_), .B(men_men_n72_), .C(men_men_n212_), .Y(men_men_n295_));
  NO2        u273(.A(men_men_n295_), .B(x04), .Y(men_men_n296_));
  NO2        u274(.A(men_men_n244_), .B(men_men_n90_), .Y(men_men_n297_));
  NO2        u275(.A(men_men_n297_), .B(men_men_n296_), .Y(men_men_n298_));
  NA3        u276(.A(men_men_n298_), .B(men_men_n294_), .C(men_men_n289_), .Y(men_men_n299_));
  NO3        u277(.A(men_men_n299_), .B(men_men_n286_), .C(men_men_n280_), .Y(men_men_n300_));
  NA2        u278(.A(men_men_n129_), .B(x03), .Y(men_men_n301_));
  INV        u279(.A(men_men_n167_), .Y(men_men_n302_));
  OAI210     u280(.A0(men_men_n49_), .A1(men_men_n34_), .B0(men_men_n35_), .Y(men_men_n303_));
  AOI220     u281(.A0(men_men_n303_), .A1(men_men_n302_), .B0(men_men_n187_), .B1(x08), .Y(men_men_n304_));
  OAI210     u282(.A0(men_men_n304_), .A1(men_men_n264_), .B0(men_men_n301_), .Y(men_men_n305_));
  NA2        u283(.A(men_men_n305_), .B(men_men_n92_), .Y(men_men_n306_));
  OAI210     u284(.A0(men_men_n53_), .A1(x05), .B0(men_men_n93_), .Y(men_men_n307_));
  NA2        u285(.A(men_men_n256_), .B(men_men_n87_), .Y(men_men_n308_));
  NA2        u286(.A(men_men_n87_), .B(men_men_n40_), .Y(men_men_n309_));
  NA3        u287(.A(men_men_n309_), .B(men_men_n308_), .C(men_men_n117_), .Y(men_men_n310_));
  NA4        u288(.A(men_men_n310_), .B(men_men_n307_), .C(men_men_n306_), .D(men_men_n47_), .Y(men_men_n311_));
  INV        u289(.A(men_men_n187_), .Y(men_men_n312_));
  INV        u290(.A(men_men_n225_), .Y(men_men_n313_));
  NA2        u291(.A(men_men_n184_), .B(x04), .Y(men_men_n314_));
  NO2        u292(.A(men_men_n314_), .B(men_men_n313_), .Y(men_men_n315_));
  NO3        u293(.A(men_men_n169_), .B(x13), .C(men_men_n30_), .Y(men_men_n316_));
  OAI210     u294(.A0(men_men_n316_), .A1(men_men_n315_), .B0(men_men_n82_), .Y(men_men_n317_));
  NO3        u295(.A(men_men_n184_), .B(men_men_n148_), .C(men_men_n50_), .Y(men_men_n318_));
  OAI210     u296(.A0(men_men_n134_), .A1(men_men_n35_), .B0(men_men_n87_), .Y(men_men_n319_));
  NA2        u297(.A(men_men_n319_), .B(men_men_n318_), .Y(men_men_n320_));
  NA3        u298(.A(men_men_n320_), .B(men_men_n317_), .C(x06), .Y(men_men_n321_));
  OAI220     u299(.A0(men_men_n149_), .A1(x09), .B0(x08), .B1(men_men_n40_), .Y(men_men_n322_));
  NO3        u300(.A(men_men_n264_), .B(men_men_n115_), .C(x08), .Y(men_men_n323_));
  AOI210     u301(.A0(men_men_n322_), .A1(men_men_n211_), .B0(men_men_n323_), .Y(men_men_n324_));
  NO2        u302(.A(men_men_n47_), .B(men_men_n40_), .Y(men_men_n325_));
  NO3        u303(.A(men_men_n99_), .B(men_men_n116_), .C(men_men_n37_), .Y(men_men_n326_));
  AOI210     u304(.A0(men_men_n318_), .A1(men_men_n325_), .B0(men_men_n326_), .Y(men_men_n327_));
  OAI210     u305(.A0(men_men_n324_), .A1(men_men_n28_), .B0(men_men_n327_), .Y(men_men_n328_));
  AN2        u306(.A(men_men_n328_), .B(x04), .Y(men_men_n329_));
  AOI210     u307(.A0(men_men_n321_), .A1(men_men_n311_), .B0(men_men_n329_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n300_), .A1(x12), .B0(men_men_n330_), .Y(men03));
  OR2        u309(.A(men_men_n41_), .B(men_men_n212_), .Y(men_men_n332_));
  AOI210     u310(.A0(men_men_n138_), .A1(men_men_n87_), .B0(men_men_n332_), .Y(men_men_n333_));
  INV        u311(.A(men_men_n188_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n334_), .A1(men_men_n333_), .B0(x05), .Y(men_men_n335_));
  NA2        u313(.A(men_men_n332_), .B(x05), .Y(men_men_n336_));
  AOI210     u314(.A0(men_men_n127_), .A1(men_men_n199_), .B0(men_men_n336_), .Y(men_men_n337_));
  AOI210     u315(.A0(men_men_n214_), .A1(men_men_n68_), .B0(men_men_n109_), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n56_), .B0(men_men_n292_), .B1(men_men_n283_), .Y(men_men_n339_));
  OAI210     u317(.A0(men_men_n339_), .A1(men_men_n337_), .B0(men_men_n87_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n133_), .A1(men_men_n57_), .B0(men_men_n37_), .Y(men_men_n341_));
  NO2        u319(.A(men_men_n158_), .B(men_men_n122_), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n36_), .Y(men_men_n343_));
  OAI210     u321(.A0(men_men_n343_), .A1(men_men_n341_), .B0(x04), .Y(men_men_n344_));
  NO3        u322(.A(men_men_n309_), .B(men_men_n73_), .C(men_men_n56_), .Y(men_men_n345_));
  AOI210     u323(.A0(men_men_n174_), .A1(men_men_n87_), .B0(men_men_n133_), .Y(men_men_n346_));
  OA210      u324(.A0(men_men_n150_), .A1(x12), .B0(men_men_n122_), .Y(men_men_n347_));
  NO3        u325(.A(men_men_n347_), .B(men_men_n346_), .C(men_men_n345_), .Y(men_men_n348_));
  NA4        u326(.A(men_men_n348_), .B(men_men_n344_), .C(men_men_n340_), .D(men_men_n335_), .Y(men04));
  NO2        u327(.A(men_men_n76_), .B(men_men_n38_), .Y(men_men_n350_));
  XO2        u328(.A(men_men_n350_), .B(men_men_n235_), .Y(men05));
  AOI210     u329(.A0(men_men_n62_), .A1(men_men_n50_), .B0(men_men_n196_), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n352_), .A1(men_men_n291_), .B0(men_men_n25_), .Y(men_men_n353_));
  NA3        u331(.A(men_men_n130_), .B(men_men_n118_), .C(men_men_n30_), .Y(men_men_n354_));
  AOI210     u332(.A0(men_men_n217_), .A1(men_men_n54_), .B0(men_men_n77_), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n24_), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n356_), .A1(men_men_n353_), .B0(men_men_n87_), .Y(men_men_n357_));
  NA2        u335(.A(x11), .B(men_men_n30_), .Y(men_men_n358_));
  NA2        u336(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n359_));
  NA2        u337(.A(men_men_n240_), .B(x03), .Y(men_men_n360_));
  OAI220     u338(.A0(men_men_n360_), .A1(men_men_n359_), .B0(men_men_n358_), .B1(men_men_n69_), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n361_), .A1(x06), .B0(men_men_n425_), .Y(men_men_n362_));
  AOI220     u340(.A0(men_men_n69_), .A1(men_men_n30_), .B0(men_men_n50_), .B1(men_men_n49_), .Y(men_men_n363_));
  NO3        u341(.A(men_men_n363_), .B(men_men_n23_), .C(x00), .Y(men_men_n364_));
  NA2        u342(.A(men_men_n61_), .B(x02), .Y(men_men_n365_));
  AOI210     u343(.A0(men_men_n365_), .A1(men_men_n360_), .B0(men_men_n242_), .Y(men_men_n366_));
  OR2        u344(.A(men_men_n366_), .B(men_men_n224_), .Y(men_men_n367_));
  NA2        u345(.A(men_men_n144_), .B(x05), .Y(men_men_n368_));
  NA3        u346(.A(men_men_n368_), .B(men_men_n228_), .C(men_men_n223_), .Y(men_men_n369_));
  NO2        u347(.A(men_men_n23_), .B(x10), .Y(men_men_n370_));
  OAI210     u348(.A0(x11), .A1(men_men_n29_), .B0(men_men_n47_), .Y(men_men_n371_));
  OR3        u349(.A(men_men_n371_), .B(men_men_n370_), .C(men_men_n43_), .Y(men_men_n372_));
  NA3        u350(.A(men_men_n372_), .B(men_men_n369_), .C(men_men_n367_), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n364_), .B0(men_men_n87_), .Y(men_men_n374_));
  INV        u352(.A(x07), .Y(men_men_n375_));
  AOI220     u353(.A0(men_men_n375_), .A1(men_men_n374_), .B0(men_men_n362_), .B1(men_men_n357_), .Y(men_men_n376_));
  NA3        u354(.A(men_men_n23_), .B(men_men_n58_), .C(men_men_n47_), .Y(men_men_n377_));
  AO210      u355(.A0(men_men_n377_), .A1(men_men_n250_), .B0(men_men_n247_), .Y(men_men_n378_));
  AOI210     u356(.A0(men_men_n370_), .A1(men_men_n64_), .B0(men_men_n129_), .Y(men_men_n379_));
  OR2        u357(.A(men_men_n379_), .B(x03), .Y(men_men_n380_));
  NA2        u358(.A(men_men_n325_), .B(men_men_n58_), .Y(men_men_n381_));
  NO2        u359(.A(men_men_n381_), .B(x11), .Y(men_men_n382_));
  NO3        u360(.A(men_men_n382_), .B(men_men_n132_), .C(men_men_n28_), .Y(men_men_n383_));
  AOI220     u361(.A0(men_men_n383_), .A1(men_men_n380_), .B0(men_men_n378_), .B1(men_men_n46_), .Y(men_men_n384_));
  NO4        u362(.A(men_men_n309_), .B(men_men_n31_), .C(x11), .D(x09), .Y(men_men_n385_));
  OAI210     u363(.A0(men_men_n385_), .A1(men_men_n384_), .B0(men_men_n88_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n314_), .A1(men_men_n95_), .B0(men_men_n246_), .Y(men_men_n387_));
  NOi21      u365(.An(men_men_n301_), .B(men_men_n122_), .Y(men_men_n388_));
  NO2        u366(.A(men_men_n387_), .B(x08), .Y(men_men_n389_));
  AOI210     u367(.A0(men_men_n370_), .A1(men_men_n28_), .B0(men_men_n30_), .Y(men_men_n390_));
  NA2        u368(.A(x09), .B(men_men_n40_), .Y(men_men_n391_));
  OAI220     u369(.A0(men_men_n391_), .A1(men_men_n390_), .B0(men_men_n358_), .B1(x06), .Y(men_men_n392_));
  NO2        u370(.A(x13), .B(x12), .Y(men_men_n393_));
  NO2        u371(.A(men_men_n118_), .B(men_men_n28_), .Y(men_men_n394_));
  NO2        u372(.A(men_men_n394_), .B(men_men_n251_), .Y(men_men_n395_));
  OR3        u373(.A(men_men_n395_), .B(x12), .C(x03), .Y(men_men_n396_));
  NA3        u374(.A(men_men_n312_), .B(men_men_n111_), .C(x12), .Y(men_men_n397_));
  AO210      u375(.A0(men_men_n312_), .A1(men_men_n111_), .B0(men_men_n235_), .Y(men_men_n398_));
  NA4        u376(.A(men_men_n398_), .B(men_men_n397_), .C(men_men_n396_), .D(x08), .Y(men_men_n399_));
  AOI210     u377(.A0(men_men_n393_), .A1(men_men_n392_), .B0(men_men_n399_), .Y(men_men_n400_));
  AOI210     u378(.A0(men_men_n389_), .A1(men_men_n386_), .B0(men_men_n400_), .Y(men_men_n401_));
  OAI210     u379(.A0(men_men_n381_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n402_));
  NA2        u380(.A(men_men_n276_), .B(x07), .Y(men_men_n403_));
  OAI220     u381(.A0(men_men_n403_), .A1(men_men_n359_), .B0(men_men_n132_), .B1(men_men_n42_), .Y(men_men_n404_));
  OAI210     u382(.A0(men_men_n404_), .A1(men_men_n402_), .B0(men_men_n173_), .Y(men_men_n405_));
  NA3        u383(.A(men_men_n395_), .B(men_men_n388_), .C(men_men_n308_), .Y(men_men_n406_));
  INV        u384(.A(x14), .Y(men_men_n407_));
  NO3        u385(.A(men_men_n301_), .B(men_men_n90_), .C(x11), .Y(men_men_n408_));
  NO3        u386(.A(men_men_n149_), .B(men_men_n64_), .C(men_men_n54_), .Y(men_men_n409_));
  NO3        u387(.A(men_men_n377_), .B(men_men_n309_), .C(men_men_n167_), .Y(men_men_n410_));
  NO4        u388(.A(men_men_n410_), .B(men_men_n409_), .C(men_men_n408_), .D(men_men_n407_), .Y(men_men_n411_));
  NA3        u389(.A(men_men_n411_), .B(men_men_n406_), .C(men_men_n405_), .Y(men_men_n412_));
  NA2        u390(.A(men_men_n394_), .B(men_men_n148_), .Y(men_men_n413_));
  NO3        u391(.A(men_men_n115_), .B(men_men_n24_), .C(x06), .Y(men_men_n414_));
  AOI210     u392(.A0(men_men_n262_), .A1(men_men_n217_), .B0(men_men_n414_), .Y(men_men_n415_));
  OAI210     u393(.A0(men_men_n43_), .A1(x04), .B0(men_men_n415_), .Y(men_men_n416_));
  NA2        u394(.A(men_men_n416_), .B(men_men_n87_), .Y(men_men_n417_));
  OAI210     u395(.A0(men_men_n413_), .A1(men_men_n78_), .B0(men_men_n417_), .Y(men_men_n418_));
  NO4        u396(.A(men_men_n418_), .B(men_men_n412_), .C(men_men_n401_), .D(men_men_n376_), .Y(men06));
  INV        u397(.A(men_men_n80_), .Y(men_men_n422_));
  INV        u398(.A(x05), .Y(men_men_n423_));
  INV        u399(.A(x02), .Y(men_men_n424_));
  INV        u400(.A(x07), .Y(men_men_n425_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule