//Benchmark atmr_alu4_1266_0.5

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n122_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n97_, mai_mai_n98_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n140_, men_men_n141_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1146_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o00(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o01(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o02(.A(i_9_), .Y(ori_ori_n25_));
  INV        o03(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o04(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o05(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o06(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o07(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o08(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o09(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o10(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o11(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o12(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o13(.A(i_4_), .Y(ori_ori_n36_));
  INV        o14(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o15(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o16(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  INV        o17(.A(ori_ori_n35_), .Y(ori1));
  INV        o18(.A(i_11_), .Y(ori_ori_n41_));
  INV        o19(.A(i_2_), .Y(ori_ori_n42_));
  INV        o20(.A(i_5_), .Y(ori_ori_n43_));
  NO2        o21(.A(i_7_), .B(i_10_), .Y(ori_ori_n44_));
  AOI210     o22(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n44_), .Y(ori_ori_n45_));
  INV        o23(.A(i_5_), .Y(ori_ori_n46_));
  NA2        o24(.A(ori_ori_n46_), .B(i_11_), .Y(ori_ori_n47_));
  INV        o25(.A(i_1_), .Y(ori_ori_n48_));
  NA2        o26(.A(ori_ori_n45_), .B(i_2_), .Y(ori_ori_n49_));
  NA2        o27(.A(i_1_), .B(i_6_), .Y(ori_ori_n50_));
  NO2        o28(.A(ori_ori_n50_), .B(ori_ori_n25_), .Y(ori_ori_n51_));
  INV        o29(.A(i_0_), .Y(ori_ori_n52_));
  NAi21      o30(.An(i_5_), .B(i_10_), .Y(ori_ori_n53_));
  NA2        o31(.A(i_5_), .B(i_9_), .Y(ori_ori_n54_));
  AOI210     o32(.A0(ori_ori_n54_), .A1(ori_ori_n53_), .B0(ori_ori_n52_), .Y(ori_ori_n55_));
  NO2        o33(.A(ori_ori_n55_), .B(ori_ori_n51_), .Y(ori_ori_n56_));
  NA2        o34(.A(i_12_), .B(i_5_), .Y(ori_ori_n57_));
  NA2        o35(.A(i_6_), .B(i_9_), .Y(ori_ori_n58_));
  INV        o36(.A(i_7_), .Y(ori_ori_n59_));
  NA2        o37(.A(ori_ori_n59_), .B(ori_ori_n37_), .Y(ori_ori_n60_));
  NA2        o38(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n61_));
  NA2        o39(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n62_));
  NO2        o40(.A(ori_ori_n62_), .B(ori_ori_n42_), .Y(ori_ori_n63_));
  NA3        o41(.A(ori_ori_n57_), .B(ori_ori_n52_), .C(ori_ori_n47_), .Y(ori2));
  NO2        o42(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n65_));
  INV        o43(.A(i_6_), .Y(ori_ori_n66_));
  NA2        o44(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NA4        o45(.A(ori_ori_n67_), .B(ori_ori_n56_), .C(ori_ori_n49_), .D(ori_ori_n30_), .Y(ori0));
  NA2        o46(.A(i_1_), .B(i_5_), .Y(ori_ori_n69_));
  NO2        o47(.A(ori_ori_n41_), .B(i_5_), .Y(ori_ori_n70_));
  INV        o48(.A(i_12_), .Y(ori_ori_n71_));
  AN2        o49(.A(i_3_), .B(i_10_), .Y(ori_ori_n72_));
  NOi21      o50(.An(i_5_), .B(i_0_), .Y(ori_ori_n73_));
  AN2        o51(.A(i_12_), .B(i_5_), .Y(ori_ori_n74_));
  NO2        o52(.A(i_0_), .B(i_11_), .Y(ori_ori_n75_));
  NO2        o53(.A(i_10_), .B(i_9_), .Y(ori_ori_n76_));
  NA2        o54(.A(ori_ori_n39_), .B(i_13_), .Y(ori_ori_n77_));
  NO2        o55(.A(ori_ori_n37_), .B(i_6_), .Y(ori_ori_n78_));
  INV        o56(.A(ori_ori_n78_), .Y(ori_ori_n79_));
  NO2        o57(.A(ori_ori_n79_), .B(ori_ori_n48_), .Y(ori_ori_n80_));
  NOi21      o58(.An(i_11_), .B(i_7_), .Y(ori_ori_n81_));
  AO210      o59(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n82_));
  NO2        o60(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n83_));
  NA2        o61(.A(ori_ori_n71_), .B(ori_ori_n48_), .Y(ori_ori_n84_));
  INV        o62(.A(ori_ori_n84_), .Y(ori_ori_n85_));
  NA2        o63(.A(ori_ori_n85_), .B(i_6_), .Y(ori_ori_n86_));
  NO2        o64(.A(i_6_), .B(i_11_), .Y(ori_ori_n87_));
  INV        o65(.A(ori_ori_n86_), .Y(ori_ori_n88_));
  INV        o66(.A(i_1_), .Y(ori_ori_n89_));
  NO2        o67(.A(ori_ori_n58_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  INV        o68(.A(ori_ori_n90_), .Y(ori_ori_n91_));
  NA2        o69(.A(ori_ori_n87_), .B(ori_ori_n48_), .Y(ori_ori_n92_));
  NA2        o70(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  OR3        o71(.A(ori_ori_n93_), .B(ori_ori_n88_), .C(ori_ori_n80_), .Y(ori5));
  INV        o72(.A(ori_ori_n76_), .Y(ori_ori_n95_));
  OA210      o73(.A0(ori_ori_n83_), .A1(ori_ori_n63_), .B0(i_13_), .Y(ori_ori_n96_));
  NA2        o74(.A(ori_ori_n72_), .B(ori_ori_n61_), .Y(ori_ori_n97_));
  NO2        o75(.A(ori_ori_n97_), .B(ori_ori_n122_), .Y(ori_ori_n98_));
  NO2        o76(.A(ori_ori_n98_), .B(ori_ori_n96_), .Y(ori_ori_n99_));
  INV        o77(.A(ori_ori_n73_), .Y(ori_ori_n100_));
  OR2        o78(.A(ori_ori_n100_), .B(i_12_), .Y(ori_ori_n101_));
  OR2        o79(.A(ori_ori_n95_), .B(ori_ori_n36_), .Y(ori_ori_n102_));
  INV        o80(.A(ori_ori_n102_), .Y(ori_ori_n103_));
  NA2        o81(.A(ori_ori_n57_), .B(ori_ori_n75_), .Y(ori_ori_n104_));
  INV        o82(.A(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o83(.A(ori_ori_n105_), .B(ori_ori_n103_), .Y(ori_ori_n106_));
  NA2        o84(.A(ori_ori_n106_), .B(ori_ori_n101_), .Y(ori3));
  NA2        o85(.A(i_9_), .B(i_0_), .Y(ori_ori_n108_));
  NO2        o86(.A(ori_ori_n108_), .B(ori_ori_n69_), .Y(ori_ori_n109_));
  NO3        o87(.A(ori_ori_n70_), .B(ori_ori_n74_), .C(i_0_), .Y(ori_ori_n110_));
  OAI210     o88(.A0(ori_ori_n110_), .A1(ori_ori_n55_), .B0(i_13_), .Y(ori_ori_n111_));
  INV        o89(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  NO2        o90(.A(ori_ori_n112_), .B(ori_ori_n109_), .Y(ori_ori_n113_));
  NA2        o91(.A(i_10_), .B(ori_ori_n43_), .Y(ori_ori_n114_));
  NO2        o92(.A(ori_ori_n114_), .B(ori_ori_n52_), .Y(ori_ori_n115_));
  INV        o93(.A(ori_ori_n115_), .Y(ori_ori_n116_));
  NA2        o94(.A(ori_ori_n116_), .B(ori_ori_n113_), .Y(ori4));
  INV        o95(.A(ori_ori_n77_), .Y(ori7));
  INV        o96(.A(ori_ori_n99_), .Y(ori6));
  INV        o97(.A(i_2_), .Y(ori_ori_n122_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NOi21      m016(.An(i_12_), .B(i_13_), .Y(mai_mai_n39_));
  INV        m017(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NAi31      m018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n41_));
  INV        m019(.A(mai_mai_n35_), .Y(mai1));
  INV        m020(.A(i_11_), .Y(mai_mai_n43_));
  NO2        m021(.A(mai_mai_n43_), .B(i_6_), .Y(mai_mai_n44_));
  INV        m022(.A(i_2_), .Y(mai_mai_n45_));
  NA2        m023(.A(i_0_), .B(i_3_), .Y(mai_mai_n46_));
  INV        m024(.A(i_5_), .Y(mai_mai_n47_));
  NO2        m025(.A(i_7_), .B(i_10_), .Y(mai_mai_n48_));
  AOI210     m026(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n48_), .Y(mai_mai_n49_));
  NA2        m027(.A(i_0_), .B(i_2_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_7_), .B(i_9_), .Y(mai_mai_n51_));
  NO2        m029(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NA3        m030(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n53_));
  NO2        m031(.A(i_1_), .B(i_6_), .Y(mai_mai_n54_));
  NA2        m032(.A(i_8_), .B(i_7_), .Y(mai_mai_n55_));
  INV        m033(.A(i_1_), .Y(mai_mai_n56_));
  NA2        m034(.A(mai_mai_n49_), .B(i_2_), .Y(mai_mai_n57_));
  AOI210     m035(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n58_));
  NA2        m036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NO2        m037(.A(mai_mai_n59_), .B(mai_mai_n25_), .Y(mai_mai_n60_));
  INV        m038(.A(i_0_), .Y(mai_mai_n61_));
  NAi21      m039(.An(i_5_), .B(i_10_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_5_), .B(i_9_), .Y(mai_mai_n63_));
  AOI210     m041(.A0(mai_mai_n63_), .A1(mai_mai_n62_), .B0(mai_mai_n61_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(mai_mai_n60_), .Y(mai_mai_n65_));
  NA2        m043(.A(i_12_), .B(i_5_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_2_), .B(i_8_), .Y(mai_mai_n67_));
  NO2        m045(.A(i_3_), .B(i_9_), .Y(mai_mai_n68_));
  NO2        m046(.A(i_3_), .B(i_7_), .Y(mai_mai_n69_));
  INV        m047(.A(i_6_), .Y(mai_mai_n70_));
  INV        m048(.A(i_11_), .Y(mai_mai_n71_));
  NO2        m049(.A(i_2_), .B(i_7_), .Y(mai_mai_n72_));
  NAi21      m050(.An(i_6_), .B(i_10_), .Y(mai_mai_n73_));
  NA2        m051(.A(i_6_), .B(i_9_), .Y(mai_mai_n74_));
  NA2        m052(.A(i_2_), .B(i_6_), .Y(mai_mai_n75_));
  AN3        m053(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n76_));
  NAi21      m054(.An(i_6_), .B(i_11_), .Y(mai_mai_n77_));
  NA2        m055(.A(mai_mai_n76_), .B(mai_mai_n32_), .Y(mai_mai_n78_));
  INV        m056(.A(i_7_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_0_), .B(i_5_), .Y(mai_mai_n80_));
  NA2        m058(.A(i_12_), .B(i_3_), .Y(mai_mai_n81_));
  NAi21      m059(.An(i_7_), .B(i_11_), .Y(mai_mai_n82_));
  AN2        m060(.A(i_2_), .B(i_10_), .Y(mai_mai_n83_));
  NO2        m061(.A(mai_mai_n83_), .B(i_7_), .Y(mai_mai_n84_));
  NA2        m062(.A(i_12_), .B(i_7_), .Y(mai_mai_n85_));
  NO2        m063(.A(mai_mai_n56_), .B(mai_mai_n26_), .Y(mai_mai_n86_));
  NA2        m064(.A(i_11_), .B(i_12_), .Y(mai_mai_n87_));
  NA2        m065(.A(mai_mai_n87_), .B(mai_mai_n78_), .Y(mai_mai_n88_));
  NA2        m066(.A(mai_mai_n79_), .B(mai_mai_n37_), .Y(mai_mai_n89_));
  NA2        m067(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n90_));
  NA2        m068(.A(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  NO2        m069(.A(mai_mai_n91_), .B(mai_mai_n45_), .Y(mai_mai_n92_));
  NA2        m070(.A(mai_mai_n74_), .B(mai_mai_n73_), .Y(mai_mai_n93_));
  NO2        m071(.A(i_1_), .B(mai_mai_n70_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_6_), .B(i_5_), .Y(mai_mai_n95_));
  NA2        m073(.A(mai_mai_n750_), .B(mai_mai_n745_), .Y(mai2));
  NO2        m074(.A(mai_mai_n56_), .B(mai_mai_n37_), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n752_), .B(mai_mai_n97_), .Y(mai_mai_n98_));
  NA4        m076(.A(mai_mai_n98_), .B(mai_mai_n65_), .C(mai_mai_n57_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m077(.A(i_8_), .B(i_7_), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n100_), .B(i_6_), .Y(mai_mai_n101_));
  NO2        m079(.A(i_12_), .B(i_13_), .Y(mai_mai_n102_));
  NAi21      m080(.An(i_5_), .B(i_11_), .Y(mai_mai_n103_));
  NOi21      m081(.An(mai_mai_n102_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m082(.A(i_0_), .B(i_1_), .Y(mai_mai_n105_));
  NA2        m083(.A(i_2_), .B(i_3_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(i_4_), .Y(mai_mai_n107_));
  NA3        m085(.A(mai_mai_n107_), .B(mai_mai_n105_), .C(mai_mai_n104_), .Y(mai_mai_n108_));
  AN2        m086(.A(mai_mai_n102_), .B(mai_mai_n68_), .Y(mai_mai_n109_));
  NA2        m087(.A(i_1_), .B(i_5_), .Y(mai_mai_n110_));
  NA2        m088(.A(i_2_), .B(mai_mai_n36_), .Y(mai_mai_n111_));
  NO3        m089(.A(mai_mai_n111_), .B(mai_mai_n110_), .C(i_13_), .Y(mai_mai_n112_));
  OR2        m090(.A(i_0_), .B(i_1_), .Y(mai_mai_n113_));
  NO3        m091(.A(mai_mai_n113_), .B(mai_mai_n66_), .C(i_13_), .Y(mai_mai_n114_));
  NAi32      m092(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n115_));
  NAi21      m093(.An(mai_mai_n115_), .B(mai_mai_n114_), .Y(mai_mai_n116_));
  NOi21      m094(.An(i_4_), .B(i_10_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(mai_mai_n39_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n118_), .B(mai_mai_n116_), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n119_), .B(mai_mai_n112_), .Y(mai_mai_n120_));
  AOI210     m098(.A0(mai_mai_n120_), .A1(mai_mai_n108_), .B0(mai_mai_n101_), .Y(mai_mai_n121_));
  NOi21      m099(.An(i_4_), .B(i_9_), .Y(mai_mai_n122_));
  NOi21      m100(.An(i_11_), .B(i_13_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(mai_mai_n122_), .Y(mai_mai_n124_));
  BUFFER     m102(.A(mai_mai_n124_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_4_), .B(i_5_), .Y(mai_mai_n126_));
  NAi21      m104(.An(i_12_), .B(i_11_), .Y(mai_mai_n127_));
  NO2        m105(.A(mai_mai_n127_), .B(i_13_), .Y(mai_mai_n128_));
  NA3        m106(.A(mai_mai_n128_), .B(mai_mai_n126_), .C(mai_mai_n68_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n129_), .B(mai_mai_n125_), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n61_), .B(mai_mai_n56_), .Y(mai_mai_n131_));
  NAi31      m109(.An(mai_mai_n741_), .B(mai_mai_n109_), .C(i_11_), .Y(mai_mai_n132_));
  NA2        m110(.A(i_3_), .B(i_5_), .Y(mai_mai_n133_));
  AOI210     m111(.A0(mai_mai_n124_), .A1(mai_mai_n132_), .B0(mai_mai_n56_), .Y(mai_mai_n134_));
  NO2        m112(.A(mai_mai_n61_), .B(i_5_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_13_), .B(i_10_), .Y(mai_mai_n136_));
  NA3        m114(.A(mai_mai_n136_), .B(mai_mai_n135_), .C(mai_mai_n43_), .Y(mai_mai_n137_));
  NO2        m115(.A(i_2_), .B(i_1_), .Y(mai_mai_n138_));
  NAi21      m116(.An(i_4_), .B(i_12_), .Y(mai_mai_n139_));
  NO4        m117(.A(mai_mai_n139_), .B(i_2_), .C(mai_mai_n137_), .D(mai_mai_n25_), .Y(mai_mai_n140_));
  NO3        m118(.A(mai_mai_n140_), .B(mai_mai_n134_), .C(mai_mai_n130_), .Y(mai_mai_n141_));
  INV        m119(.A(i_8_), .Y(mai_mai_n142_));
  NO3        m120(.A(i_3_), .B(mai_mai_n70_), .C(mai_mai_n47_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(i_7_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n39_), .B(mai_mai_n43_), .Y(mai_mai_n145_));
  NO3        m123(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n146_));
  OAI210     m124(.A0(mai_mai_n76_), .A1(i_12_), .B0(mai_mai_n146_), .Y(mai_mai_n147_));
  AOI210     m125(.A0(mai_mai_n147_), .A1(mai_mai_n145_), .B0(mai_mai_n144_), .Y(mai_mai_n148_));
  NO3        m126(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n149_), .B(mai_mai_n39_), .Y(mai_mai_n150_));
  NO2        m128(.A(i_13_), .B(i_9_), .Y(mai_mai_n151_));
  NAi21      m129(.An(i_12_), .B(i_3_), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n43_), .B(i_5_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n54_), .B(mai_mai_n150_), .Y(mai_mai_n154_));
  AOI210     m132(.A0(mai_mai_n154_), .A1(i_7_), .B0(mai_mai_n148_), .Y(mai_mai_n155_));
  OAI210     m133(.A0(mai_mai_n155_), .A1(i_4_), .B0(mai_mai_n141_), .Y(mai_mai_n156_));
  NA3        m134(.A(i_13_), .B(mai_mai_n142_), .C(i_10_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n157_), .B(i_12_), .Y(mai_mai_n158_));
  NA2        m136(.A(i_0_), .B(i_5_), .Y(mai_mai_n159_));
  NAi31      m137(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n45_), .B(mai_mai_n56_), .Y(mai_mai_n161_));
  INV        m139(.A(i_13_), .Y(mai_mai_n162_));
  NO2        m140(.A(i_12_), .B(mai_mai_n162_), .Y(mai_mai_n163_));
  NA2        m141(.A(mai_mai_n163_), .B(mai_mai_n143_), .Y(mai_mai_n164_));
  INV        m142(.A(mai_mai_n164_), .Y(mai_mai_n165_));
  AOI210     m143(.A0(mai_mai_n165_), .A1(mai_mai_n100_), .B0(mai_mai_n158_), .Y(mai_mai_n166_));
  NO2        m144(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n133_), .B(i_4_), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  OR2        m147(.A(i_8_), .B(i_7_), .Y(mai_mai_n170_));
  INV        m148(.A(i_12_), .Y(mai_mai_n171_));
  NO3        m149(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n172_));
  NA2        m150(.A(i_2_), .B(i_1_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n174_));
  NO3        m152(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n175_));
  NAi21      m153(.An(i_4_), .B(i_3_), .Y(mai_mai_n176_));
  NO2        m154(.A(i_0_), .B(i_6_), .Y(mai_mai_n177_));
  NOi41      m155(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n178_));
  NA2        m156(.A(mai_mai_n178_), .B(mai_mai_n177_), .Y(mai_mai_n179_));
  AOI220     m157(.A0(mai_mai_n178_), .A1(mai_mai_n39_), .B0(mai_mai_n174_), .B1(mai_mai_n151_), .Y(mai_mai_n180_));
  NO2        m158(.A(i_11_), .B(mai_mai_n162_), .Y(mai_mai_n181_));
  NOi21      m159(.An(i_1_), .B(i_6_), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n171_), .B(i_9_), .Y(mai_mai_n183_));
  NO2        m161(.A(i_12_), .B(i_3_), .Y(mai_mai_n184_));
  NA2        m162(.A(i_3_), .B(i_9_), .Y(mai_mai_n185_));
  NAi21      m163(.An(i_7_), .B(i_10_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NA3        m165(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n188_));
  INV        m166(.A(mai_mai_n101_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n171_), .B(i_13_), .Y(mai_mai_n190_));
  NO2        m168(.A(mai_mai_n190_), .B(mai_mai_n63_), .Y(mai_mai_n191_));
  AOI220     m169(.A0(mai_mai_n191_), .A1(mai_mai_n189_), .B0(i_9_), .B1(mai_mai_n181_), .Y(mai_mai_n192_));
  NO2        m170(.A(mai_mai_n170_), .B(mai_mai_n37_), .Y(mai_mai_n193_));
  NA2        m171(.A(i_12_), .B(i_6_), .Y(mai_mai_n194_));
  OR2        m172(.A(i_13_), .B(i_9_), .Y(mai_mai_n195_));
  NO3        m173(.A(mai_mai_n195_), .B(mai_mai_n194_), .C(mai_mai_n47_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n176_), .B(i_2_), .Y(mai_mai_n197_));
  NA3        m175(.A(mai_mai_n197_), .B(mai_mai_n196_), .C(mai_mai_n43_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n181_), .B(i_9_), .Y(mai_mai_n199_));
  OAI210     m177(.A0(mai_mai_n56_), .A1(mai_mai_n199_), .B0(mai_mai_n198_), .Y(mai_mai_n200_));
  NO3        m178(.A(i_11_), .B(mai_mai_n162_), .C(mai_mai_n25_), .Y(mai_mai_n201_));
  INV        m179(.A(mai_mai_n201_), .Y(mai_mai_n202_));
  NA3        m180(.A(i_6_), .B(mai_mai_n193_), .C(mai_mai_n163_), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n203_), .A1(mai_mai_n202_), .B0(mai_mai_n45_), .Y(mai_mai_n204_));
  AOI210     m182(.A0(mai_mai_n200_), .A1(mai_mai_n193_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  NA4        m183(.A(mai_mai_n205_), .B(mai_mai_n192_), .C(mai_mai_n180_), .D(mai_mai_n166_), .Y(mai_mai_n206_));
  NO3        m184(.A(i_12_), .B(mai_mai_n162_), .C(mai_mai_n37_), .Y(mai_mai_n207_));
  INV        m185(.A(mai_mai_n207_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n173_), .B(i_0_), .Y(mai_mai_n209_));
  NO2        m187(.A(i_3_), .B(i_10_), .Y(mai_mai_n210_));
  NA3        m188(.A(mai_mai_n210_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n211_));
  AN2        m189(.A(i_3_), .B(i_10_), .Y(mai_mai_n212_));
  NO2        m190(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n45_), .B(mai_mai_n26_), .Y(mai_mai_n214_));
  OAI220     m192(.A0(mai_mai_n211_), .A1(i_6_), .B0(i_3_), .B1(mai_mai_n208_), .Y(mai_mai_n215_));
  NO4        m193(.A(mai_mai_n215_), .B(mai_mai_n206_), .C(mai_mai_n156_), .D(mai_mai_n121_), .Y(mai_mai_n216_));
  NO3        m194(.A(mai_mai_n43_), .B(i_13_), .C(i_9_), .Y(mai_mai_n217_));
  NO2        m195(.A(i_2_), .B(i_3_), .Y(mai_mai_n218_));
  NO2        m196(.A(i_12_), .B(i_10_), .Y(mai_mai_n219_));
  NOi21      m197(.An(i_5_), .B(i_0_), .Y(mai_mai_n220_));
  NA3        m198(.A(mai_mai_n36_), .B(mai_mai_n70_), .C(i_8_), .Y(mai_mai_n221_));
  NO2        m199(.A(i_6_), .B(i_8_), .Y(mai_mai_n222_));
  NO2        m200(.A(i_1_), .B(i_7_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n75_), .B(mai_mai_n142_), .Y(mai_mai_n224_));
  AOI210     m202(.A0(mai_mai_n54_), .A1(i_3_), .B0(mai_mai_n118_), .Y(mai_mai_n225_));
  AOI210     m203(.A0(i_12_), .A1(mai_mai_n217_), .B0(mai_mai_n225_), .Y(mai_mai_n226_));
  NOi32      m204(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n227_), .Y(mai_mai_n228_));
  NAi21      m206(.An(i_1_), .B(i_5_), .Y(mai_mai_n229_));
  OAI210     m207(.A0(i_9_), .A1(mai_mai_n115_), .B0(mai_mai_n179_), .Y(mai_mai_n230_));
  NAi41      m208(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n231_));
  OAI220     m209(.A0(mai_mai_n231_), .A1(mai_mai_n229_), .B0(mai_mai_n160_), .B1(mai_mai_n115_), .Y(mai_mai_n232_));
  AOI210     m210(.A0(mai_mai_n231_), .A1(mai_mai_n115_), .B0(mai_mai_n113_), .Y(mai_mai_n233_));
  NOi32      m211(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n234_));
  NA2        m212(.A(mai_mai_n234_), .B(mai_mai_n45_), .Y(mai_mai_n235_));
  NO2        m213(.A(mai_mai_n235_), .B(i_0_), .Y(mai_mai_n236_));
  OR3        m214(.A(mai_mai_n236_), .B(mai_mai_n233_), .C(mai_mai_n232_), .Y(mai_mai_n237_));
  NAi21      m215(.An(i_3_), .B(i_4_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n238_), .B(i_9_), .Y(mai_mai_n239_));
  INV        m217(.A(mai_mai_n239_), .Y(mai_mai_n240_));
  NA2        m218(.A(i_2_), .B(i_7_), .Y(mai_mai_n241_));
  NO2        m219(.A(mai_mai_n238_), .B(i_10_), .Y(mai_mai_n242_));
  NA3        m220(.A(mai_mai_n242_), .B(mai_mai_n241_), .C(mai_mai_n177_), .Y(mai_mai_n243_));
  AOI210     m221(.A0(mai_mai_n243_), .A1(mai_mai_n240_), .B0(mai_mai_n135_), .Y(mai_mai_n244_));
  AOI210     m222(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n245_));
  INV        m223(.A(mai_mai_n242_), .Y(mai_mai_n246_));
  AOI220     m224(.A0(mai_mai_n242_), .A1(mai_mai_n223_), .B0(mai_mai_n172_), .B1(mai_mai_n138_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n247_), .A1(mai_mai_n246_), .B0(i_5_), .Y(mai_mai_n248_));
  NO4        m226(.A(mai_mai_n248_), .B(mai_mai_n244_), .C(mai_mai_n237_), .D(mai_mai_n230_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n249_), .B(mai_mai_n228_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n55_), .B(mai_mai_n25_), .Y(mai_mai_n251_));
  AN2        m229(.A(i_12_), .B(i_5_), .Y(mai_mai_n252_));
  NO2        m230(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n253_), .B(mai_mai_n252_), .Y(mai_mai_n254_));
  NO2        m232(.A(i_11_), .B(mai_mai_n254_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n176_), .B(i_5_), .Y(mai_mai_n256_));
  NO2        m234(.A(i_5_), .B(i_10_), .Y(mai_mai_n257_));
  NO2        m235(.A(i_11_), .B(mai_mai_n176_), .Y(mai_mai_n258_));
  OAI210     m236(.A0(mai_mai_n258_), .A1(mai_mai_n255_), .B0(mai_mai_n251_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n108_), .B(mai_mai_n70_), .Y(mai_mai_n261_));
  OAI210     m239(.A0(mai_mai_n261_), .A1(mai_mai_n255_), .B0(mai_mai_n260_), .Y(mai_mai_n262_));
  NO3        m240(.A(mai_mai_n70_), .B(mai_mai_n47_), .C(i_9_), .Y(mai_mai_n263_));
  NO2        m241(.A(i_11_), .B(i_12_), .Y(mai_mai_n264_));
  NO2        m242(.A(i_10_), .B(i_11_), .Y(mai_mai_n265_));
  NAi21      m243(.An(i_13_), .B(i_0_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n266_), .B(mai_mai_n173_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n740_), .A1(mai_mai_n265_), .B0(mai_mai_n267_), .Y(mai_mai_n268_));
  NA3        m246(.A(mai_mai_n268_), .B(mai_mai_n262_), .C(mai_mai_n259_), .Y(mai_mai_n269_));
  NO2        m247(.A(i_0_), .B(i_11_), .Y(mai_mai_n270_));
  AN2        m248(.A(i_1_), .B(i_6_), .Y(mai_mai_n271_));
  NOi21      m249(.An(i_2_), .B(i_12_), .Y(mai_mai_n272_));
  NA2        m250(.A(mai_mai_n100_), .B(i_9_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n273_), .B(i_4_), .Y(mai_mai_n274_));
  NA2        m252(.A(mai_mai_n272_), .B(mai_mai_n274_), .Y(mai_mai_n275_));
  OR2        m253(.A(i_13_), .B(i_10_), .Y(mai_mai_n276_));
  NO3        m254(.A(mai_mai_n276_), .B(mai_mai_n87_), .C(i_9_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n124_), .B(mai_mai_n89_), .Y(mai_mai_n278_));
  BUFFER     m256(.A(mai_mai_n157_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n79_), .B(mai_mai_n25_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n207_), .B(mai_mai_n280_), .Y(mai_mai_n281_));
  NA2        m259(.A(i_5_), .B(i_1_), .Y(mai_mai_n282_));
  OAI220     m260(.A0(mai_mai_n282_), .A1(mai_mai_n279_), .B0(mai_mai_n281_), .B1(mai_mai_n80_), .Y(mai_mai_n283_));
  INV        m261(.A(mai_mai_n283_), .Y(mai_mai_n284_));
  AOI210     m262(.A0(mai_mai_n284_), .A1(mai_mai_n275_), .B0(mai_mai_n26_), .Y(mai_mai_n285_));
  NO4        m263(.A(mai_mai_n748_), .B(mai_mai_n285_), .C(mai_mai_n269_), .D(mai_mai_n250_), .Y(mai_mai_n286_));
  NO2        m264(.A(mai_mai_n61_), .B(i_13_), .Y(mai_mai_n287_));
  NO2        m265(.A(i_10_), .B(i_9_), .Y(mai_mai_n288_));
  NO2        m266(.A(i_12_), .B(i_3_), .Y(mai_mai_n289_));
  NO2        m267(.A(i_4_), .B(mai_mai_n150_), .Y(mai_mai_n290_));
  NO3        m268(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n291_));
  NA2        m269(.A(mai_mai_n194_), .B(mai_mai_n77_), .Y(mai_mai_n292_));
  NA2        m270(.A(mai_mai_n292_), .B(mai_mai_n291_), .Y(mai_mai_n293_));
  NA2        m271(.A(i_8_), .B(i_9_), .Y(mai_mai_n294_));
  INV        m272(.A(mai_mai_n207_), .Y(mai_mai_n295_));
  OAI220     m273(.A0(mai_mai_n295_), .A1(mai_mai_n294_), .B0(mai_mai_n293_), .B1(mai_mai_n214_), .Y(mai_mai_n296_));
  NA2        m274(.A(mai_mai_n181_), .B(mai_mai_n213_), .Y(mai_mai_n297_));
  NO3        m275(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n298_));
  AOI210     m276(.A0(mai_mai_n184_), .A1(mai_mai_n138_), .B0(mai_mai_n298_), .Y(mai_mai_n299_));
  NA3        m277(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n300_));
  NA4        m278(.A(mai_mai_n103_), .B(mai_mai_n86_), .C(mai_mai_n66_), .D(mai_mai_n23_), .Y(mai_mai_n301_));
  OAI220     m279(.A0(mai_mai_n301_), .A1(mai_mai_n300_), .B0(mai_mai_n299_), .B1(mai_mai_n297_), .Y(mai_mai_n302_));
  NO3        m280(.A(mai_mai_n302_), .B(mai_mai_n296_), .C(mai_mai_n290_), .Y(mai_mai_n303_));
  OR2        m281(.A(i_8_), .B(mai_mai_n169_), .Y(mai_mai_n304_));
  NA2        m282(.A(mai_mai_n76_), .B(i_13_), .Y(mai_mai_n305_));
  NA2        m283(.A(i_3_), .B(mai_mai_n251_), .Y(mai_mai_n306_));
  NO2        m284(.A(i_2_), .B(i_13_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n306_), .B(mai_mai_n305_), .Y(mai_mai_n308_));
  NO3        m286(.A(i_4_), .B(mai_mai_n47_), .C(i_8_), .Y(mai_mai_n309_));
  NO2        m287(.A(i_6_), .B(i_7_), .Y(mai_mai_n310_));
  NO2        m288(.A(i_11_), .B(i_1_), .Y(mai_mai_n311_));
  OR2        m289(.A(i_11_), .B(i_8_), .Y(mai_mai_n312_));
  NOi21      m290(.An(i_2_), .B(i_7_), .Y(mai_mai_n313_));
  NAi31      m291(.An(mai_mai_n312_), .B(mai_mai_n313_), .C(i_0_), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n276_), .B(mai_mai_n314_), .Y(mai_mai_n315_));
  NO2        m293(.A(i_6_), .B(i_10_), .Y(mai_mai_n316_));
  NA3        m294(.A(mai_mai_n178_), .B(mai_mai_n123_), .C(mai_mai_n95_), .Y(mai_mai_n317_));
  NO2        m295(.A(mai_mai_n113_), .B(i_3_), .Y(mai_mai_n318_));
  NAi31      m296(.An(i_11_), .B(mai_mai_n318_), .C(mai_mai_n163_), .Y(mai_mai_n319_));
  NA3        m297(.A(mai_mai_n260_), .B(mai_mai_n131_), .C(mai_mai_n107_), .Y(mai_mai_n320_));
  NA3        m298(.A(mai_mai_n320_), .B(mai_mai_n319_), .C(mai_mai_n317_), .Y(mai_mai_n321_));
  NO4        m299(.A(mai_mai_n321_), .B(mai_mai_n217_), .C(mai_mai_n315_), .D(mai_mai_n308_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n291_), .B(mai_mai_n252_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n298_), .B(mai_mai_n257_), .Y(mai_mai_n324_));
  INV        m302(.A(mai_mai_n323_), .Y(mai_mai_n325_));
  NAi21      m303(.An(mai_mai_n157_), .B(mai_mai_n264_), .Y(mai_mai_n326_));
  NA3        m304(.A(i_6_), .B(i_3_), .C(mai_mai_n100_), .Y(mai_mai_n327_));
  OAI220     m305(.A0(mai_mai_n38_), .A1(mai_mai_n327_), .B0(i_1_), .B1(mai_mai_n326_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n217_), .B(mai_mai_n172_), .Y(mai_mai_n330_));
  OAI210     m308(.A0(mai_mai_n329_), .A1(mai_mai_n305_), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  NO3        m309(.A(mai_mai_n331_), .B(mai_mai_n328_), .C(mai_mai_n325_), .Y(mai_mai_n332_));
  NA4        m310(.A(mai_mai_n332_), .B(mai_mai_n322_), .C(mai_mai_n304_), .D(mai_mai_n303_), .Y(mai_mai_n333_));
  NA3        m311(.A(mai_mai_n212_), .B(mai_mai_n128_), .C(mai_mai_n126_), .Y(mai_mai_n334_));
  OAI210     m312(.A0(mai_mai_n211_), .A1(mai_mai_n741_), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  INV        m313(.A(mai_mai_n335_), .Y(mai_mai_n336_));
  NA2        m314(.A(mai_mai_n252_), .B(mai_mai_n162_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n227_), .B(mai_mai_n61_), .Y(mai_mai_n338_));
  NA2        m316(.A(i_6_), .B(mai_mai_n234_), .Y(mai_mai_n339_));
  AO210      m317(.A0(mai_mai_n338_), .A1(mai_mai_n337_), .B0(mai_mai_n339_), .Y(mai_mai_n340_));
  NO2        m318(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n341_));
  NAi31      m319(.An(mai_mai_n338_), .B(mai_mai_n316_), .C(mai_mai_n45_), .Y(mai_mai_n342_));
  INV        m320(.A(mai_mai_n277_), .Y(mai_mai_n343_));
  NA3        m321(.A(mai_mai_n343_), .B(mai_mai_n342_), .C(mai_mai_n340_), .Y(mai_mai_n344_));
  INV        m322(.A(mai_mai_n344_), .Y(mai_mai_n345_));
  NO2        m323(.A(i_7_), .B(mai_mai_n145_), .Y(mai_mai_n346_));
  NO2        m324(.A(mai_mai_n133_), .B(mai_mai_n70_), .Y(mai_mai_n347_));
  AOI210     m325(.A0(mai_mai_n347_), .A1(mai_mai_n346_), .B0(mai_mai_n278_), .Y(mai_mai_n348_));
  NA3        m326(.A(mai_mai_n348_), .B(mai_mai_n345_), .C(mai_mai_n336_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n276_), .B(mai_mai_n38_), .Y(mai_mai_n350_));
  NA2        m328(.A(mai_mai_n350_), .B(mai_mai_n253_), .Y(mai_mai_n351_));
  NO2        m329(.A(i_8_), .B(i_7_), .Y(mai_mai_n352_));
  INV        m330(.A(mai_mai_n161_), .Y(mai_mai_n353_));
  NA2        m331(.A(mai_mai_n43_), .B(i_10_), .Y(mai_mai_n354_));
  NO2        m332(.A(mai_mai_n354_), .B(i_6_), .Y(mai_mai_n355_));
  NA3        m333(.A(mai_mai_n355_), .B(mai_mai_n739_), .C(mai_mai_n352_), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n133_), .A1(mai_mai_n190_), .B0(mai_mai_n305_), .Y(mai_mai_n357_));
  NA2        m335(.A(mai_mai_n357_), .B(mai_mai_n193_), .Y(mai_mai_n358_));
  NOi31      m336(.An(mai_mai_n209_), .B(mai_mai_n211_), .C(mai_mai_n741_), .Y(mai_mai_n359_));
  NA3        m337(.A(mai_mai_n212_), .B(mai_mai_n126_), .C(mai_mai_n76_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n113_), .B(i_5_), .Y(mai_mai_n361_));
  NA2        m339(.A(mai_mai_n361_), .B(mai_mai_n218_), .Y(mai_mai_n362_));
  NA2        m340(.A(mai_mai_n362_), .B(mai_mai_n360_), .Y(mai_mai_n363_));
  OAI210     m341(.A0(mai_mai_n363_), .A1(mai_mai_n359_), .B0(mai_mai_n298_), .Y(mai_mai_n364_));
  NA4        m342(.A(mai_mai_n364_), .B(mai_mai_n358_), .C(mai_mai_n356_), .D(mai_mai_n351_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n207_), .B(mai_mai_n69_), .Y(mai_mai_n366_));
  AOI210     m344(.A0(i_11_), .A1(mai_mai_n67_), .B0(mai_mai_n366_), .Y(mai_mai_n367_));
  NA2        m345(.A(i_0_), .B(mai_mai_n47_), .Y(mai_mai_n368_));
  NO2        m346(.A(mai_mai_n201_), .B(mai_mai_n367_), .Y(mai_mai_n369_));
  NO4        m347(.A(mai_mai_n182_), .B(mai_mai_n41_), .C(i_2_), .D(mai_mai_n47_), .Y(mai_mai_n370_));
  NO3        m348(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n371_));
  OA210      m349(.A0(mai_mai_n371_), .A1(mai_mai_n370_), .B0(mai_mai_n227_), .Y(mai_mai_n372_));
  NO2        m350(.A(mai_mai_n276_), .B(i_1_), .Y(mai_mai_n373_));
  NOi31      m351(.An(mai_mai_n373_), .B(mai_mai_n292_), .C(mai_mai_n61_), .Y(mai_mai_n374_));
  AN4        m352(.A(mai_mai_n374_), .B(mai_mai_n274_), .C(i_3_), .D(i_2_), .Y(mai_mai_n375_));
  INV        m353(.A(mai_mai_n129_), .Y(mai_mai_n376_));
  NO3        m354(.A(mai_mai_n376_), .B(mai_mai_n375_), .C(mai_mai_n372_), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n70_), .B(mai_mai_n25_), .Y(mai_mai_n378_));
  AOI220     m356(.A0(mai_mai_n207_), .A1(mai_mai_n378_), .B0(mai_mai_n201_), .B1(i_6_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(mai_mai_n214_), .Y(mai_mai_n380_));
  NO2        m358(.A(mai_mai_n85_), .B(mai_mai_n23_), .Y(mai_mai_n381_));
  NA2        m359(.A(mai_mai_n124_), .B(mai_mai_n132_), .Y(mai_mai_n382_));
  NOi21      m360(.An(mai_mai_n104_), .B(mai_mai_n221_), .Y(mai_mai_n383_));
  NO3        m361(.A(mai_mai_n383_), .B(mai_mai_n382_), .C(mai_mai_n380_), .Y(mai_mai_n384_));
  NO2        m362(.A(mai_mai_n338_), .B(mai_mai_n247_), .Y(mai_mai_n385_));
  NA2        m363(.A(i_6_), .B(mai_mai_n201_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n207_), .B(mai_mai_n159_), .Y(mai_mai_n387_));
  AOI210     m365(.A0(mai_mai_n387_), .A1(mai_mai_n386_), .B0(i_3_), .Y(mai_mai_n388_));
  NO3        m366(.A(i_4_), .B(i_8_), .C(mai_mai_n211_), .Y(mai_mai_n389_));
  INV        m367(.A(mai_mai_n326_), .Y(mai_mai_n390_));
  NO4        m368(.A(mai_mai_n390_), .B(mai_mai_n389_), .C(mai_mai_n388_), .D(mai_mai_n385_), .Y(mai_mai_n391_));
  NA4        m369(.A(mai_mai_n391_), .B(mai_mai_n384_), .C(mai_mai_n377_), .D(mai_mai_n369_), .Y(mai_mai_n392_));
  NO4        m370(.A(mai_mai_n392_), .B(mai_mai_n365_), .C(mai_mai_n349_), .D(mai_mai_n333_), .Y(mai_mai_n393_));
  NA4        m371(.A(mai_mai_n393_), .B(mai_mai_n286_), .C(mai_mai_n226_), .D(mai_mai_n216_), .Y(mai7));
  NA2        m372(.A(mai_mai_n316_), .B(mai_mai_n69_), .Y(mai_mai_n395_));
  NA2        m373(.A(i_11_), .B(mai_mai_n142_), .Y(mai_mai_n396_));
  NO2        m374(.A(i_13_), .B(mai_mai_n395_), .Y(mai_mai_n397_));
  NA3        m375(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n398_));
  NO2        m376(.A(mai_mai_n171_), .B(i_4_), .Y(mai_mai_n399_));
  NA2        m377(.A(mai_mai_n399_), .B(i_8_), .Y(mai_mai_n400_));
  NA2        m378(.A(i_2_), .B(mai_mai_n70_), .Y(mai_mai_n401_));
  INV        m379(.A(mai_mai_n149_), .Y(mai_mai_n402_));
  NO2        m380(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n402_), .B(i_13_), .Y(mai_mai_n404_));
  NO2        m382(.A(mai_mai_n404_), .B(mai_mai_n397_), .Y(mai_mai_n405_));
  OR2        m383(.A(i_6_), .B(i_10_), .Y(mai_mai_n406_));
  NO2        m384(.A(mai_mai_n406_), .B(mai_mai_n23_), .Y(mai_mai_n407_));
  OR3        m385(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n408_));
  INV        m386(.A(mai_mai_n146_), .Y(mai_mai_n409_));
  OA220      m387(.A0(mai_mai_n408_), .A1(i_3_), .B0(i_10_), .B1(mai_mai_n195_), .Y(mai_mai_n410_));
  AOI210     m388(.A0(mai_mai_n410_), .A1(mai_mai_n405_), .B0(mai_mai_n56_), .Y(mai_mai_n411_));
  NOi21      m389(.An(i_11_), .B(i_7_), .Y(mai_mai_n412_));
  AO210      m390(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n413_));
  NO2        m391(.A(mai_mai_n413_), .B(mai_mai_n412_), .Y(mai_mai_n414_));
  NA2        m392(.A(mai_mai_n71_), .B(mai_mai_n56_), .Y(mai_mai_n415_));
  AO210      m393(.A0(mai_mai_n415_), .A1(mai_mai_n247_), .B0(mai_mai_n40_), .Y(mai_mai_n416_));
  NA2        m394(.A(mai_mai_n163_), .B(mai_mai_n56_), .Y(mai_mai_n417_));
  OR2        m395(.A(mai_mai_n152_), .B(mai_mai_n82_), .Y(mai_mai_n418_));
  NO2        m396(.A(mai_mai_n56_), .B(i_9_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n417_), .B(mai_mai_n416_), .Y(mai_mai_n420_));
  NA2        m398(.A(mai_mai_n420_), .B(i_6_), .Y(mai_mai_n421_));
  NO2        m399(.A(mai_mai_n171_), .B(mai_mai_n70_), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n422_), .B(i_11_), .Y(mai_mai_n423_));
  NA2        m401(.A(mai_mai_n343_), .B(mai_mai_n293_), .Y(mai_mai_n424_));
  NO3        m402(.A(i_12_), .B(i_13_), .C(mai_mai_n70_), .Y(mai_mai_n425_));
  NA2        m403(.A(mai_mai_n425_), .B(mai_mai_n419_), .Y(mai_mai_n426_));
  NO3        m404(.A(mai_mai_n406_), .B(mai_mai_n170_), .C(mai_mai_n23_), .Y(mai_mai_n427_));
  AOI210     m405(.A0(i_1_), .A1(mai_mai_n187_), .B0(mai_mai_n427_), .Y(mai_mai_n428_));
  OAI210     m406(.A0(mai_mai_n428_), .A1(mai_mai_n43_), .B0(mai_mai_n426_), .Y(mai_mai_n429_));
  NA3        m407(.A(mai_mai_n352_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n430_));
  INV        m408(.A(i_2_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n97_), .B(i_9_), .Y(mai_mai_n432_));
  NO2        m410(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  NA3        m411(.A(mai_mai_n419_), .B(mai_mai_n218_), .C(i_6_), .Y(mai_mai_n434_));
  NO2        m412(.A(mai_mai_n434_), .B(mai_mai_n23_), .Y(mai_mai_n435_));
  AOI210     m413(.A0(mai_mai_n311_), .A1(mai_mai_n280_), .B0(mai_mai_n175_), .Y(mai_mai_n436_));
  NO2        m414(.A(mai_mai_n436_), .B(mai_mai_n401_), .Y(mai_mai_n437_));
  NO2        m415(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n438_));
  NA2        m416(.A(mai_mai_n438_), .B(mai_mai_n24_), .Y(mai_mai_n439_));
  OR3        m417(.A(mai_mai_n437_), .B(mai_mai_n435_), .C(mai_mai_n433_), .Y(mai_mai_n440_));
  NO3        m418(.A(mai_mai_n440_), .B(mai_mai_n429_), .C(mai_mai_n424_), .Y(mai_mai_n441_));
  NO2        m419(.A(mai_mai_n171_), .B(mai_mai_n79_), .Y(mai_mai_n442_));
  NO2        m420(.A(mai_mai_n442_), .B(mai_mai_n412_), .Y(mai_mai_n443_));
  NO2        m421(.A(mai_mai_n757_), .B(mai_mai_n408_), .Y(mai_mai_n444_));
  NO2        m422(.A(i_9_), .B(mai_mai_n70_), .Y(mai_mai_n445_));
  NA2        m423(.A(mai_mai_n444_), .B(mai_mai_n45_), .Y(mai_mai_n446_));
  NA2        m424(.A(i_3_), .B(mai_mai_n142_), .Y(mai_mai_n447_));
  NA2        m425(.A(i_1_), .B(i_3_), .Y(mai_mai_n448_));
  NA3        m426(.A(mai_mai_n446_), .B(mai_mai_n441_), .C(mai_mai_n421_), .Y(mai_mai_n449_));
  AN2        m427(.A(mai_mai_n178_), .B(mai_mai_n70_), .Y(mai_mai_n450_));
  NA2        m428(.A(i_6_), .B(mai_mai_n239_), .Y(mai_mai_n451_));
  NA2        m429(.A(mai_mai_n316_), .B(mai_mai_n45_), .Y(mai_mai_n452_));
  NA2        m430(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n453_));
  NA3        m431(.A(mai_mai_n117_), .B(mai_mai_n69_), .C(mai_mai_n70_), .Y(mai_mai_n454_));
  NA4        m432(.A(mai_mai_n454_), .B(mai_mai_n453_), .C(mai_mai_n452_), .D(mai_mai_n451_), .Y(mai_mai_n455_));
  OAI210     m433(.A0(mai_mai_n455_), .A1(mai_mai_n450_), .B0(i_1_), .Y(mai_mai_n456_));
  AOI210     m434(.A0(mai_mai_n194_), .A1(mai_mai_n77_), .B0(i_1_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n238_), .B(i_2_), .Y(mai_mai_n458_));
  NA2        m436(.A(mai_mai_n458_), .B(mai_mai_n457_), .Y(mai_mai_n459_));
  OAI210     m437(.A0(mai_mai_n434_), .A1(i_12_), .B0(mai_mai_n459_), .Y(mai_mai_n460_));
  INV        m438(.A(mai_mai_n460_), .Y(mai_mai_n461_));
  AOI210     m439(.A0(mai_mai_n461_), .A1(mai_mai_n456_), .B0(i_13_), .Y(mai_mai_n462_));
  NA2        m440(.A(mai_mai_n307_), .B(mai_mai_n117_), .Y(mai_mai_n463_));
  NO2        m441(.A(mai_mai_n463_), .B(mai_mai_n43_), .Y(mai_mai_n464_));
  NO2        m442(.A(mai_mai_n51_), .B(i_12_), .Y(mai_mai_n465_));
  AOI210     m443(.A0(mai_mai_n178_), .A1(mai_mai_n94_), .B0(mai_mai_n445_), .Y(mai_mai_n466_));
  OAI220     m444(.A0(mai_mai_n466_), .A1(mai_mai_n40_), .B0(mai_mai_n736_), .B1(mai_mai_n75_), .Y(mai_mai_n467_));
  AOI210     m445(.A0(mai_mai_n464_), .A1(mai_mai_n222_), .B0(mai_mai_n467_), .Y(mai_mai_n468_));
  NOi31      m446(.An(mai_mai_n753_), .B(mai_mai_n395_), .C(mai_mai_n43_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n93_), .B(i_13_), .Y(mai_mai_n470_));
  NO2        m448(.A(mai_mai_n470_), .B(mai_mai_n457_), .Y(mai_mai_n471_));
  NO2        m449(.A(mai_mai_n59_), .B(mai_mai_n79_), .Y(mai_mai_n472_));
  NO3        m450(.A(mai_mai_n313_), .B(mai_mai_n171_), .C(mai_mai_n70_), .Y(mai_mai_n473_));
  NO2        m451(.A(mai_mai_n473_), .B(mai_mai_n472_), .Y(mai_mai_n474_));
  NO2        m452(.A(mai_mai_n474_), .B(mai_mai_n409_), .Y(mai_mai_n475_));
  NO3        m453(.A(mai_mai_n475_), .B(mai_mai_n471_), .C(mai_mai_n469_), .Y(mai_mai_n476_));
  NA3        m454(.A(mai_mai_n272_), .B(mai_mai_n403_), .C(mai_mai_n77_), .Y(mai_mai_n477_));
  NA2        m455(.A(mai_mai_n423_), .B(i_13_), .Y(mai_mai_n478_));
  NAi21      m456(.An(i_11_), .B(i_12_), .Y(mai_mai_n479_));
  NOi41      m457(.An(mai_mai_n84_), .B(mai_mai_n479_), .C(i_13_), .D(mai_mai_n70_), .Y(mai_mai_n480_));
  AOI210     m458(.A0(mai_mai_n755_), .A1(mai_mai_n217_), .B0(mai_mai_n480_), .Y(mai_mai_n481_));
  NA3        m459(.A(mai_mai_n481_), .B(mai_mai_n478_), .C(mai_mai_n477_), .Y(mai_mai_n482_));
  NA2        m460(.A(mai_mai_n482_), .B(mai_mai_n56_), .Y(mai_mai_n483_));
  NO2        m461(.A(i_2_), .B(i_12_), .Y(mai_mai_n484_));
  NO2        m462(.A(i_3_), .B(i_2_), .Y(mai_mai_n485_));
  NA3        m463(.A(mai_mai_n756_), .B(mai_mai_n44_), .C(mai_mai_n162_), .Y(mai_mai_n486_));
  NA4        m464(.A(mai_mai_n486_), .B(mai_mai_n483_), .C(mai_mai_n476_), .D(mai_mai_n468_), .Y(mai_mai_n487_));
  OR4        m465(.A(mai_mai_n487_), .B(mai_mai_n462_), .C(mai_mai_n449_), .D(mai_mai_n411_), .Y(mai5));
  AOI210     m466(.A0(mai_mai_n443_), .A1(mai_mai_n197_), .B0(mai_mai_n278_), .Y(mai_mai_n489_));
  AO210      m467(.A0(mai_mai_n24_), .A1(i_10_), .B0(mai_mai_n181_), .Y(mai_mai_n490_));
  NA2        m468(.A(mai_mai_n490_), .B(mai_mai_n484_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n400_), .B(i_11_), .Y(mai_mai_n492_));
  OAI210     m470(.A0(mai_mai_n403_), .A1(mai_mai_n72_), .B0(mai_mai_n492_), .Y(mai_mai_n493_));
  NA4        m471(.A(mai_mai_n493_), .B(mai_mai_n491_), .C(mai_mai_n489_), .D(mai_mai_n343_), .Y(mai_mai_n494_));
  NO3        m472(.A(i_11_), .B(mai_mai_n171_), .C(i_13_), .Y(mai_mai_n495_));
  NO2        m473(.A(mai_mai_n90_), .B(mai_mai_n23_), .Y(mai_mai_n496_));
  NA2        m474(.A(i_12_), .B(i_8_), .Y(mai_mai_n497_));
  OAI210     m475(.A0(mai_mai_n45_), .A1(i_3_), .B0(mai_mai_n497_), .Y(mai_mai_n498_));
  INV        m476(.A(mai_mai_n288_), .Y(mai_mai_n499_));
  AOI220     m477(.A0(mai_mai_n218_), .A1(mai_mai_n381_), .B0(mai_mai_n498_), .B1(mai_mai_n496_), .Y(mai_mai_n500_));
  INV        m478(.A(mai_mai_n500_), .Y(mai_mai_n501_));
  NO2        m479(.A(mai_mai_n501_), .B(mai_mai_n494_), .Y(mai_mai_n502_));
  INV        m480(.A(mai_mai_n123_), .Y(mai_mai_n503_));
  INV        m481(.A(mai_mai_n178_), .Y(mai_mai_n504_));
  OAI210     m482(.A0(mai_mai_n458_), .A1(mai_mai_n289_), .B0(mai_mai_n84_), .Y(mai_mai_n505_));
  AOI210     m483(.A0(mai_mai_n505_), .A1(mai_mai_n504_), .B0(mai_mai_n503_), .Y(mai_mai_n506_));
  NO2        m484(.A(mai_mai_n294_), .B(mai_mai_n26_), .Y(mai_mai_n507_));
  NO2        m485(.A(mai_mai_n507_), .B(mai_mai_n280_), .Y(mai_mai_n508_));
  NA2        m486(.A(mai_mai_n508_), .B(i_2_), .Y(mai_mai_n509_));
  INV        m487(.A(mai_mai_n509_), .Y(mai_mai_n510_));
  AOI210     m488(.A0(mai_mai_n754_), .A1(mai_mai_n510_), .B0(mai_mai_n506_), .Y(mai_mai_n511_));
  NO2        m489(.A(mai_mai_n139_), .B(mai_mai_n91_), .Y(mai_mai_n512_));
  OAI210     m490(.A0(mai_mai_n512_), .A1(mai_mai_n496_), .B0(i_2_), .Y(mai_mai_n513_));
  INV        m491(.A(mai_mai_n124_), .Y(mai_mai_n514_));
  NO3        m492(.A(mai_mai_n413_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n515_));
  AOI210     m493(.A0(mai_mai_n514_), .A1(mai_mai_n72_), .B0(mai_mai_n515_), .Y(mai_mai_n516_));
  AOI210     m494(.A0(mai_mai_n516_), .A1(mai_mai_n513_), .B0(mai_mai_n142_), .Y(mai_mai_n517_));
  OA210      m495(.A0(mai_mai_n414_), .A1(mai_mai_n92_), .B0(i_13_), .Y(mai_mai_n518_));
  INV        m496(.A(mai_mai_n146_), .Y(mai_mai_n519_));
  NA2        m497(.A(mai_mai_n109_), .B(mai_mai_n396_), .Y(mai_mai_n520_));
  AOI210     m498(.A0(mai_mai_n520_), .A1(mai_mai_n519_), .B0(mai_mai_n241_), .Y(mai_mai_n521_));
  AOI210     m499(.A0(mai_mai_n152_), .A1(mai_mai_n106_), .B0(mai_mai_n341_), .Y(mai_mai_n522_));
  OAI210     m500(.A0(mai_mai_n522_), .A1(mai_mai_n163_), .B0(mai_mai_n280_), .Y(mai_mai_n523_));
  NO2        m501(.A(i_2_), .B(mai_mai_n43_), .Y(mai_mai_n524_));
  NA3        m502(.A(mai_mai_n212_), .B(mai_mai_n90_), .C(mai_mai_n41_), .Y(mai_mai_n525_));
  OAI210     m503(.A0(mai_mai_n525_), .A1(mai_mai_n524_), .B0(mai_mai_n523_), .Y(mai_mai_n526_));
  NO4        m504(.A(mai_mai_n526_), .B(mai_mai_n521_), .C(mai_mai_n518_), .D(mai_mai_n517_), .Y(mai_mai_n527_));
  INV        m505(.A(mai_mai_n381_), .Y(mai_mai_n528_));
  NA2        m506(.A(mai_mai_n495_), .B(i_7_), .Y(mai_mai_n529_));
  NA2        m507(.A(mai_mai_n529_), .B(mai_mai_n528_), .Y(mai_mai_n530_));
  NO2        m508(.A(i_2_), .B(i_12_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n531_), .B(mai_mai_n92_), .Y(mai_mai_n532_));
  NO2        m510(.A(mai_mai_n532_), .B(mai_mai_n396_), .Y(mai_mai_n533_));
  AOI220     m511(.A0(mai_mai_n533_), .A1(mai_mai_n36_), .B0(mai_mai_n530_), .B1(mai_mai_n45_), .Y(mai_mai_n534_));
  NA4        m512(.A(mai_mai_n534_), .B(mai_mai_n527_), .C(mai_mai_n511_), .D(mai_mai_n502_), .Y(mai6));
  OAI210     m513(.A0(mai_mai_n25_), .A1(mai_mai_n742_), .B0(mai_mai_n485_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n160_), .B(i_11_), .Y(mai_mai_n537_));
  NO2        m515(.A(i_11_), .B(i_9_), .Y(mai_mai_n538_));
  OR2        m516(.A(mai_mai_n536_), .B(i_12_), .Y(mai_mai_n539_));
  NA2        m517(.A(mai_mai_n242_), .B(mai_mai_n223_), .Y(mai_mai_n540_));
  NA4        m518(.A(mai_mai_n415_), .B(mai_mai_n312_), .C(i_12_), .D(mai_mai_n540_), .Y(mai_mai_n541_));
  AOI220     m519(.A0(mai_mai_n143_), .A1(mai_mai_n538_), .B0(mai_mai_n541_), .B1(mai_mai_n61_), .Y(mai_mai_n542_));
  INV        m520(.A(mai_mai_n219_), .Y(mai_mai_n543_));
  AOI210     m521(.A0(mai_mai_n90_), .A1(i_5_), .B0(mai_mai_n543_), .Y(mai_mai_n544_));
  NA2        m522(.A(mai_mai_n737_), .B(mai_mai_n531_), .Y(mai_mai_n545_));
  AOI210     m523(.A0(mai_mai_n545_), .A1(mai_mai_n339_), .B0(mai_mai_n135_), .Y(mai_mai_n546_));
  INV        m524(.A(i_11_), .Y(mai_mai_n547_));
  NA3        m525(.A(mai_mai_n547_), .B(mai_mai_n310_), .C(mai_mai_n257_), .Y(mai_mai_n548_));
  NAi32      m526(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n549_));
  AOI210     m527(.A0(i_11_), .A1(i_11_), .B0(mai_mai_n549_), .Y(mai_mai_n550_));
  NA2        m528(.A(i_4_), .B(mai_mai_n371_), .Y(mai_mai_n551_));
  NAi31      m529(.An(mai_mai_n550_), .B(mai_mai_n551_), .C(mai_mai_n548_), .Y(mai_mai_n552_));
  OR3        m530(.A(mai_mai_n552_), .B(mai_mai_n546_), .C(mai_mai_n544_), .Y(mai_mai_n553_));
  NA3        m531(.A(mai_mai_n749_), .B(mai_mai_n184_), .C(i_7_), .Y(mai_mai_n554_));
  OR2        m532(.A(mai_mai_n414_), .B(mai_mai_n289_), .Y(mai_mai_n555_));
  NA2        m533(.A(mai_mai_n555_), .B(mai_mai_n105_), .Y(mai_mai_n556_));
  AO210      m534(.A0(mai_mai_n324_), .A1(mai_mai_n499_), .B0(mai_mai_n36_), .Y(mai_mai_n557_));
  NA3        m535(.A(mai_mai_n557_), .B(mai_mai_n556_), .C(mai_mai_n554_), .Y(mai_mai_n558_));
  AOI210     m536(.A0(mai_mai_n738_), .A1(mai_mai_n371_), .B0(mai_mai_n537_), .Y(mai_mai_n559_));
  NA3        m537(.A(mai_mai_n241_), .B(mai_mai_n172_), .C(mai_mai_n105_), .Y(mai_mai_n560_));
  OAI210     m538(.A0(mai_mai_n263_), .A1(mai_mai_n149_), .B0(mai_mai_n58_), .Y(mai_mai_n561_));
  NA4        m539(.A(mai_mai_n561_), .B(mai_mai_n560_), .C(mai_mai_n559_), .D(mai_mai_n402_), .Y(mai_mai_n562_));
  AO210      m540(.A0(mai_mai_n341_), .A1(mai_mai_n45_), .B0(mai_mai_n71_), .Y(mai_mai_n563_));
  NA3        m541(.A(mai_mai_n563_), .B(mai_mai_n316_), .C(mai_mai_n159_), .Y(mai_mai_n564_));
  AOI210     m542(.A0(mai_mai_n289_), .A1(mai_mai_n288_), .B0(mai_mai_n370_), .Y(mai_mai_n565_));
  NA3        m543(.A(mai_mai_n744_), .B(mai_mai_n219_), .C(i_7_), .Y(mai_mai_n566_));
  NA4        m544(.A(mai_mai_n566_), .B(mai_mai_n743_), .C(mai_mai_n565_), .D(mai_mai_n564_), .Y(mai_mai_n567_));
  NO4        m545(.A(mai_mai_n567_), .B(mai_mai_n562_), .C(mai_mai_n558_), .D(mai_mai_n553_), .Y(mai_mai_n568_));
  NA4        m546(.A(mai_mai_n568_), .B(mai_mai_n542_), .C(mai_mai_n539_), .D(mai_mai_n249_), .Y(mai3));
  NA2        m547(.A(i_12_), .B(i_10_), .Y(mai_mai_n570_));
  NA2        m548(.A(i_6_), .B(i_7_), .Y(mai_mai_n571_));
  NO2        m549(.A(mai_mai_n571_), .B(i_0_), .Y(mai_mai_n572_));
  NO2        m550(.A(i_11_), .B(mai_mai_n171_), .Y(mai_mai_n573_));
  OAI210     m551(.A0(mai_mai_n572_), .A1(mai_mai_n209_), .B0(mai_mai_n573_), .Y(mai_mai_n574_));
  NA3        m552(.A(mai_mai_n560_), .B(mai_mai_n402_), .C(mai_mai_n240_), .Y(mai_mai_n575_));
  NA2        m553(.A(mai_mai_n575_), .B(mai_mai_n39_), .Y(mai_mai_n576_));
  NO3        m554(.A(mai_mai_n418_), .B(mai_mai_n294_), .C(mai_mai_n94_), .Y(mai_mai_n577_));
  NA2        m555(.A(mai_mai_n272_), .B(mai_mai_n44_), .Y(mai_mai_n578_));
  NO2        m556(.A(mai_mai_n52_), .B(mai_mai_n577_), .Y(mai_mai_n579_));
  AOI210     m557(.A0(mai_mai_n579_), .A1(mai_mai_n576_), .B0(mai_mai_n47_), .Y(mai_mai_n580_));
  NO3        m558(.A(mai_mai_n245_), .B(mai_mai_n38_), .C(i_0_), .Y(mai_mai_n581_));
  INV        m559(.A(mai_mai_n581_), .Y(mai_mai_n582_));
  NA2        m560(.A(mai_mai_n753_), .B(mai_mai_n746_), .Y(mai_mai_n583_));
  NA2        m561(.A(i_0_), .B(i_5_), .Y(mai_mai_n584_));
  OAI220     m562(.A0(mai_mai_n584_), .A1(mai_mai_n583_), .B0(mai_mai_n582_), .B1(mai_mai_n56_), .Y(mai_mai_n585_));
  NOi21      m563(.An(i_5_), .B(i_9_), .Y(mai_mai_n586_));
  NA2        m564(.A(mai_mai_n586_), .B(mai_mai_n287_), .Y(mai_mai_n587_));
  NO3        m565(.A(mai_mai_n273_), .B(mai_mai_n194_), .C(mai_mai_n61_), .Y(mai_mai_n588_));
  NO2        m566(.A(mai_mai_n127_), .B(mai_mai_n106_), .Y(mai_mai_n589_));
  AOI210     m567(.A0(mai_mai_n589_), .A1(mai_mai_n177_), .B0(mai_mai_n588_), .Y(mai_mai_n590_));
  OAI220     m568(.A0(mai_mai_n590_), .A1(mai_mai_n741_), .B0(i_12_), .B1(mai_mai_n587_), .Y(mai_mai_n591_));
  NO4        m569(.A(mai_mai_n591_), .B(mai_mai_n585_), .C(mai_mai_n580_), .D(mai_mai_n751_), .Y(mai_mai_n592_));
  INV        m570(.A(mai_mai_n217_), .Y(mai_mai_n593_));
  OAI220     m571(.A0(mai_mai_n118_), .A1(i_0_), .B0(mai_mai_n593_), .B1(i_10_), .Y(mai_mai_n594_));
  INV        m572(.A(mai_mai_n594_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n378_), .B(i_0_), .Y(mai_mai_n596_));
  NO3        m574(.A(mai_mai_n596_), .B(mai_mai_n254_), .C(mai_mai_n72_), .Y(mai_mai_n597_));
  NO4        m575(.A(i_5_), .B(i_12_), .C(mai_mai_n276_), .D(mai_mai_n271_), .Y(mai_mai_n598_));
  AOI210     m576(.A0(mai_mai_n598_), .A1(i_11_), .B0(mai_mai_n597_), .Y(mai_mai_n599_));
  NA2        m577(.A(mai_mai_n495_), .B(mai_mai_n220_), .Y(mai_mai_n600_));
  OAI220     m578(.A0(i_6_), .A1(mai_mai_n600_), .B0(mai_mai_n439_), .B1(mai_mai_n353_), .Y(mai_mai_n601_));
  NO2        m579(.A(mai_mai_n183_), .B(mai_mai_n110_), .Y(mai_mai_n602_));
  NO4        m580(.A(mai_mai_n85_), .B(mai_mai_n54_), .C(mai_mai_n447_), .D(i_5_), .Y(mai_mai_n603_));
  AO220      m581(.A0(mai_mai_n603_), .A1(mai_mai_n43_), .B0(mai_mai_n602_), .B1(i_6_), .Y(mai_mai_n604_));
  NO2        m582(.A(i_3_), .B(mai_mai_n600_), .Y(mai_mai_n605_));
  NO3        m583(.A(mai_mai_n605_), .B(mai_mai_n604_), .C(mai_mai_n601_), .Y(mai_mai_n606_));
  NA3        m584(.A(mai_mai_n606_), .B(mai_mai_n599_), .C(mai_mai_n595_), .Y(mai_mai_n607_));
  NA2        m585(.A(i_11_), .B(i_9_), .Y(mai_mai_n608_));
  NO3        m586(.A(i_12_), .B(mai_mai_n608_), .C(mai_mai_n401_), .Y(mai_mai_n609_));
  AO220      m587(.A0(mai_mai_n609_), .A1(i_10_), .B0(mai_mai_n196_), .B1(mai_mai_n71_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n608_), .B(mai_mai_n61_), .Y(mai_mai_n611_));
  NO2        m589(.A(mai_mai_n127_), .B(i_0_), .Y(mai_mai_n612_));
  NA2        m590(.A(mai_mai_n310_), .B(mai_mai_n168_), .Y(mai_mai_n613_));
  OAI220     m591(.A0(i_12_), .A1(mai_mai_n587_), .B0(mai_mai_n613_), .B1(mai_mai_n127_), .Y(mai_mai_n614_));
  NO3        m592(.A(mai_mai_n614_), .B(mai_mai_n114_), .C(mai_mai_n610_), .Y(mai_mai_n615_));
  NA2        m593(.A(mai_mai_n438_), .B(i_1_), .Y(mai_mai_n616_));
  NO2        m594(.A(i_6_), .B(mai_mai_n616_), .Y(mai_mai_n617_));
  NA2        m595(.A(mai_mai_n123_), .B(mai_mai_n80_), .Y(mai_mai_n618_));
  NOi21      m596(.An(mai_mai_n138_), .B(mai_mai_n618_), .Y(mai_mai_n619_));
  NO2        m597(.A(i_0_), .B(mai_mai_n578_), .Y(mai_mai_n620_));
  NO3        m598(.A(mai_mai_n620_), .B(mai_mai_n619_), .C(mai_mai_n617_), .Y(mai_mai_n621_));
  NOi21      m599(.An(i_7_), .B(mai_mai_n479_), .Y(mai_mai_n622_));
  NA3        m600(.A(mai_mai_n622_), .B(mai_mai_n253_), .C(i_6_), .Y(mai_mai_n623_));
  OA210      m601(.A0(mai_mai_n618_), .A1(mai_mai_n339_), .B0(mai_mai_n623_), .Y(mai_mai_n624_));
  NO3        m602(.A(mai_mai_n266_), .B(mai_mai_n231_), .C(mai_mai_n229_), .Y(mai_mai_n625_));
  INV        m603(.A(mai_mai_n188_), .Y(mai_mai_n626_));
  NO2        m604(.A(mai_mai_n479_), .B(mai_mai_n185_), .Y(mai_mai_n627_));
  AOI210     m605(.A0(mai_mai_n627_), .A1(mai_mai_n626_), .B0(mai_mai_n625_), .Y(mai_mai_n628_));
  NA4        m606(.A(mai_mai_n628_), .B(mai_mai_n624_), .C(mai_mai_n621_), .D(mai_mai_n615_), .Y(mai_mai_n629_));
  AN2        m607(.A(mai_mai_n220_), .B(mai_mai_n589_), .Y(mai_mai_n630_));
  NA2        m608(.A(mai_mai_n630_), .B(i_10_), .Y(mai_mai_n631_));
  NO2        m609(.A(mai_mai_n570_), .B(mai_mai_n218_), .Y(mai_mai_n632_));
  OA210      m610(.A0(mai_mai_n310_), .A1(mai_mai_n161_), .B0(mai_mai_n309_), .Y(mai_mai_n633_));
  OAI210     m611(.A0(mai_mai_n633_), .A1(mai_mai_n632_), .B0(mai_mai_n611_), .Y(mai_mai_n634_));
  NA3        m612(.A(mai_mai_n309_), .B(mai_mai_n272_), .C(mai_mai_n44_), .Y(mai_mai_n635_));
  OAI210     m613(.A0(mai_mai_n118_), .A1(i_7_), .B0(mai_mai_n635_), .Y(mai_mai_n636_));
  NA2        m614(.A(mai_mai_n611_), .B(mai_mai_n212_), .Y(mai_mai_n637_));
  NA2        m615(.A(mai_mai_n137_), .B(mai_mai_n637_), .Y(mai_mai_n638_));
  AOI220     m616(.A0(mai_mai_n638_), .A1(mai_mai_n310_), .B0(mai_mai_n636_), .B1(mai_mai_n61_), .Y(mai_mai_n639_));
  NA3        m617(.A(i_5_), .B(mai_mai_n251_), .C(mai_mai_n422_), .Y(mai_mai_n640_));
  NA2        m618(.A(mai_mai_n75_), .B(mai_mai_n43_), .Y(mai_mai_n641_));
  NO2        m619(.A(mai_mai_n63_), .B(mai_mai_n497_), .Y(mai_mai_n642_));
  NA2        m620(.A(mai_mai_n642_), .B(mai_mai_n641_), .Y(mai_mai_n643_));
  AOI210     m621(.A0(mai_mai_n643_), .A1(mai_mai_n640_), .B0(mai_mai_n46_), .Y(mai_mai_n644_));
  NAi21      m622(.An(i_9_), .B(i_5_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n645_), .B(mai_mai_n266_), .Y(mai_mai_n646_));
  NO2        m624(.A(mai_mai_n398_), .B(mai_mai_n81_), .Y(mai_mai_n647_));
  AOI220     m625(.A0(mai_mai_n647_), .A1(i_0_), .B0(mai_mai_n646_), .B1(mai_mai_n414_), .Y(mai_mai_n648_));
  OAI220     m626(.A0(mai_mai_n648_), .A1(mai_mai_n70_), .B0(i_0_), .B1(mai_mai_n124_), .Y(mai_mai_n649_));
  NO3        m627(.A(mai_mai_n649_), .B(mai_mai_n644_), .C(mai_mai_n344_), .Y(mai_mai_n650_));
  NA4        m628(.A(mai_mai_n650_), .B(mai_mai_n639_), .C(mai_mai_n634_), .D(mai_mai_n631_), .Y(mai_mai_n651_));
  NO3        m629(.A(mai_mai_n651_), .B(mai_mai_n629_), .C(mai_mai_n607_), .Y(mai_mai_n652_));
  INV        m630(.A(mai_mai_n479_), .Y(mai_mai_n653_));
  NO3        m631(.A(mai_mai_n81_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n654_));
  AO220      m632(.A0(mai_mai_n654_), .A1(mai_mai_n43_), .B0(mai_mai_n653_), .B1(mai_mai_n126_), .Y(mai_mai_n655_));
  AOI210     m633(.A0(i_12_), .A1(mai_mai_n451_), .B0(mai_mai_n618_), .Y(mai_mai_n656_));
  AOI210     m634(.A0(mai_mai_n655_), .A1(mai_mai_n224_), .B0(mai_mai_n656_), .Y(mai_mai_n657_));
  NA3        m635(.A(mai_mai_n104_), .B(mai_mai_n746_), .C(mai_mai_n61_), .Y(mai_mai_n658_));
  NO2        m636(.A(mai_mai_n551_), .B(mai_mai_n266_), .Y(mai_mai_n659_));
  NA2        m637(.A(mai_mai_n573_), .B(i_9_), .Y(mai_mai_n660_));
  AOI210     m638(.A0(i_0_), .A1(mai_mai_n327_), .B0(mai_mai_n660_), .Y(mai_mai_n661_));
  OAI210     m639(.A0(mai_mai_n177_), .A1(i_9_), .B0(mai_mai_n167_), .Y(mai_mai_n662_));
  NO2        m640(.A(mai_mai_n662_), .B(mai_mai_n110_), .Y(mai_mai_n663_));
  NO3        m641(.A(mai_mai_n663_), .B(mai_mai_n661_), .C(mai_mai_n659_), .Y(mai_mai_n664_));
  NA3        m642(.A(mai_mai_n664_), .B(mai_mai_n658_), .C(mai_mai_n657_), .Y(mai_mai_n665_));
  NA2        m643(.A(mai_mai_n220_), .B(mai_mai_n241_), .Y(mai_mai_n666_));
  AOI210     m644(.A0(mai_mai_n211_), .A1(mai_mai_n118_), .B0(mai_mai_n666_), .Y(mai_mai_n667_));
  INV        m645(.A(mai_mai_n667_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n374_), .B(mai_mai_n63_), .Y(mai_mai_n669_));
  NO3        m647(.A(mai_mai_n153_), .B(mai_mai_n252_), .C(i_0_), .Y(mai_mai_n670_));
  OAI210     m648(.A0(mai_mai_n670_), .A1(mai_mai_n64_), .B0(i_13_), .Y(mai_mai_n671_));
  INV        m649(.A(mai_mai_n159_), .Y(mai_mai_n672_));
  NO2        m650(.A(i_12_), .B(mai_mai_n409_), .Y(mai_mai_n673_));
  NA3        m651(.A(mai_mai_n673_), .B(i_7_), .C(mai_mai_n672_), .Y(mai_mai_n674_));
  NA4        m652(.A(mai_mai_n674_), .B(mai_mai_n671_), .C(mai_mai_n669_), .D(mai_mai_n668_), .Y(mai_mai_n675_));
  NO2        m653(.A(mai_mai_n176_), .B(mai_mai_n75_), .Y(mai_mai_n676_));
  NA2        m654(.A(mai_mai_n676_), .B(mai_mai_n653_), .Y(mai_mai_n677_));
  NA2        m655(.A(mai_mai_n749_), .B(mai_mai_n128_), .Y(mai_mai_n678_));
  OA220      m656(.A0(mai_mai_n678_), .A1(i_0_), .B0(mai_mai_n677_), .B1(i_5_), .Y(mai_mai_n679_));
  AOI210     m657(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n127_), .Y(mai_mai_n680_));
  NA2        m658(.A(mai_mai_n680_), .B(mai_mai_n633_), .Y(mai_mai_n681_));
  NA2        m659(.A(mai_mai_n407_), .B(mai_mai_n135_), .Y(mai_mai_n682_));
  NA2        m660(.A(mai_mai_n682_), .B(mai_mai_n360_), .Y(mai_mai_n683_));
  NO3        m661(.A(mai_mai_n578_), .B(mai_mai_n51_), .C(mai_mai_n47_), .Y(mai_mai_n684_));
  NA2        m662(.A(mai_mai_n323_), .B(mai_mai_n317_), .Y(mai_mai_n685_));
  NO3        m663(.A(mai_mai_n685_), .B(mai_mai_n684_), .C(mai_mai_n683_), .Y(mai_mai_n686_));
  NA3        m664(.A(mai_mai_n257_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n687_));
  INV        m665(.A(mai_mai_n687_), .Y(mai_mai_n688_));
  NOi31      m666(.An(mai_mai_n256_), .B(i_11_), .C(mai_mai_n173_), .Y(mai_mai_n689_));
  NO3        m667(.A(mai_mai_n608_), .B(mai_mai_n159_), .C(mai_mai_n139_), .Y(mai_mai_n690_));
  NO3        m668(.A(mai_mai_n690_), .B(mai_mai_n689_), .C(mai_mai_n688_), .Y(mai_mai_n691_));
  NA4        m669(.A(mai_mai_n691_), .B(mai_mai_n686_), .C(mai_mai_n681_), .D(mai_mai_n679_), .Y(mai_mai_n692_));
  NO3        m670(.A(mai_mai_n408_), .B(mai_mai_n368_), .C(i_7_), .Y(mai_mai_n693_));
  NA3        m671(.A(mai_mai_n573_), .B(mai_mai_n83_), .C(mai_mai_n90_), .Y(mai_mai_n694_));
  INV        m672(.A(mai_mai_n694_), .Y(mai_mai_n695_));
  AOI210     m673(.A0(mai_mai_n695_), .A1(i_6_), .B0(mai_mai_n693_), .Y(mai_mai_n696_));
  NAi21      m674(.An(mai_mai_n175_), .B(mai_mai_n176_), .Y(mai_mai_n697_));
  NO3        m675(.A(mai_mai_n173_), .B(i_0_), .C(i_12_), .Y(mai_mai_n698_));
  AOI220     m676(.A0(mai_mai_n698_), .A1(mai_mai_n697_), .B0(mai_mai_n257_), .B1(mai_mai_n128_), .Y(mai_mai_n699_));
  NO3        m677(.A(i_12_), .B(mai_mai_n430_), .C(mai_mai_n94_), .Y(mai_mai_n700_));
  NA2        m678(.A(mai_mai_n700_), .B(mai_mai_n159_), .Y(mai_mai_n701_));
  NA2        m679(.A(mai_mai_n307_), .B(mai_mai_n612_), .Y(mai_mai_n702_));
  NA4        m680(.A(mai_mai_n702_), .B(mai_mai_n701_), .C(mai_mai_n699_), .D(mai_mai_n696_), .Y(mai_mai_n703_));
  NO4        m681(.A(mai_mai_n703_), .B(mai_mai_n692_), .C(mai_mai_n675_), .D(mai_mai_n665_), .Y(mai_mai_n704_));
  NA2        m682(.A(mai_mai_n747_), .B(mai_mai_n151_), .Y(mai_mai_n705_));
  NO2        m683(.A(mai_mai_n300_), .B(mai_mai_n194_), .Y(mai_mai_n706_));
  NO2        m684(.A(mai_mai_n706_), .B(mai_mai_n598_), .Y(mai_mai_n707_));
  INV        m685(.A(mai_mai_n707_), .Y(mai_mai_n708_));
  AOI210     m686(.A0(mai_mai_n136_), .A1(mai_mai_n47_), .B0(mai_mai_n708_), .Y(mai_mai_n709_));
  AOI210     m687(.A0(mai_mai_n709_), .A1(mai_mai_n705_), .B0(mai_mai_n61_), .Y(mai_mai_n710_));
  NO2        m688(.A(mai_mai_n371_), .B(mai_mai_n248_), .Y(mai_mai_n711_));
  NO2        m689(.A(mai_mai_n711_), .B(mai_mai_n503_), .Y(mai_mai_n712_));
  INV        m690(.A(mai_mai_n622_), .Y(mai_mai_n713_));
  NO2        m691(.A(mai_mai_n713_), .B(mai_mai_n448_), .Y(mai_mai_n714_));
  INV        m692(.A(mai_mai_n53_), .Y(mai_mai_n715_));
  NA2        m693(.A(mai_mai_n715_), .B(mai_mai_n64_), .Y(mai_mai_n716_));
  NO2        m694(.A(mai_mai_n716_), .B(mai_mai_n171_), .Y(mai_mai_n717_));
  NO2        m695(.A(mai_mai_n717_), .B(mai_mai_n714_), .Y(mai_mai_n718_));
  OAI210     m696(.A0(mai_mai_n196_), .A1(mai_mai_n114_), .B0(mai_mai_n72_), .Y(mai_mai_n719_));
  NA3        m697(.A(mai_mai_n507_), .B(mai_mai_n209_), .C(mai_mai_n66_), .Y(mai_mai_n720_));
  AOI210     m698(.A0(mai_mai_n720_), .A1(mai_mai_n719_), .B0(i_11_), .Y(mai_mai_n721_));
  INV        m699(.A(mai_mai_n151_), .Y(mai_mai_n722_));
  NA2        m700(.A(i_0_), .B(i_5_), .Y(mai_mai_n723_));
  AOI210     m701(.A0(mai_mai_n722_), .A1(mai_mai_n519_), .B0(mai_mai_n723_), .Y(mai_mai_n724_));
  NO3        m702(.A(mai_mai_n55_), .B(mai_mai_n54_), .C(i_4_), .Y(mai_mai_n725_));
  OAI210     m703(.A0(mai_mai_n626_), .A1(mai_mai_n213_), .B0(mai_mai_n725_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n726_), .B(mai_mai_n479_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n550_), .B(mai_mai_n232_), .Y(mai_mai_n728_));
  NO2        m706(.A(mai_mai_n728_), .B(mai_mai_n40_), .Y(mai_mai_n729_));
  NO4        m707(.A(mai_mai_n729_), .B(mai_mai_n727_), .C(mai_mai_n724_), .D(mai_mai_n721_), .Y(mai_mai_n730_));
  OAI210     m708(.A0(mai_mai_n718_), .A1(i_4_), .B0(mai_mai_n730_), .Y(mai_mai_n731_));
  NO3        m709(.A(mai_mai_n731_), .B(mai_mai_n712_), .C(mai_mai_n710_), .Y(mai_mai_n732_));
  NA4        m710(.A(mai_mai_n732_), .B(mai_mai_n704_), .C(mai_mai_n652_), .D(mai_mai_n592_), .Y(mai4));
  INV        m711(.A(mai_mai_n465_), .Y(mai_mai_n736_));
  INV        m712(.A(i_9_), .Y(mai_mai_n737_));
  INV        m713(.A(i_11_), .Y(mai_mai_n738_));
  INV        m714(.A(mai_mai_n176_), .Y(mai_mai_n739_));
  INV        m715(.A(mai_mai_n160_), .Y(mai_mai_n740_));
  INV        m716(.A(i_5_), .Y(mai_mai_n741_));
  INV        m717(.A(i_9_), .Y(mai_mai_n742_));
  INV        m718(.A(mai_mai_n270_), .Y(mai_mai_n743_));
  INV        m719(.A(i_5_), .Y(mai_mai_n744_));
  INV        m720(.A(mai_mai_n64_), .Y(mai_mai_n745_));
  INV        m721(.A(i_9_), .Y(mai_mai_n746_));
  INV        m722(.A(i_10_), .Y(mai_mai_n747_));
  INV        m723(.A(mai_mai_n199_), .Y(mai_mai_n748_));
  INV        m724(.A(i_9_), .Y(mai_mai_n749_));
  INV        m725(.A(mai_mai_n88_), .Y(mai_mai_n750_));
  INV        m726(.A(mai_mai_n574_), .Y(mai_mai_n751_));
  INV        m727(.A(i_6_), .Y(mai_mai_n752_));
  INV        m728(.A(i_13_), .Y(mai_mai_n753_));
  INV        m729(.A(mai_mai_n276_), .Y(mai_mai_n754_));
  INV        m730(.A(i_6_), .Y(mai_mai_n755_));
  INV        m731(.A(i_1_), .Y(mai_mai_n756_));
  INV        m732(.A(i_1_), .Y(mai_mai_n757_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  NOi21      u0006(.An(i_11_), .B(i_8_), .Y(men_men_n29_));
  AO210      u0007(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n30_));
  OR2        u0008(.A(men_men_n30_), .B(men_men_n29_), .Y(men_men_n31_));
  NA2        u0009(.A(men_men_n31_), .B(men_men_n26_), .Y(men_men_n32_));
  XO2        u0010(.A(men_men_n32_), .B(men_men_n23_), .Y(men_men_n33_));
  INV        u0011(.A(i_4_), .Y(men_men_n34_));
  INV        u0012(.A(i_10_), .Y(men_men_n35_));
  NAi21      u0013(.An(i_11_), .B(i_9_), .Y(men_men_n36_));
  NOi21      u0014(.An(i_12_), .B(i_13_), .Y(men_men_n37_));
  INV        u0015(.A(men_men_n37_), .Y(men_men_n38_));
  NO2        u0016(.A(men_men_n34_), .B(i_3_), .Y(men_men_n39_));
  NAi31      u0017(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n33_), .Y(men1));
  INV        u0019(.A(i_11_), .Y(men_men_n42_));
  NO2        u0020(.A(men_men_n42_), .B(i_6_), .Y(men_men_n43_));
  INV        u0021(.A(i_2_), .Y(men_men_n44_));
  NA2        u0022(.A(i_0_), .B(i_3_), .Y(men_men_n45_));
  INV        u0023(.A(i_5_), .Y(men_men_n46_));
  NO2        u0024(.A(i_7_), .B(i_10_), .Y(men_men_n47_));
  AOI210     u0025(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n47_), .Y(men_men_n48_));
  OAI210     u0026(.A0(men_men_n48_), .A1(i_3_), .B0(men_men_n46_), .Y(men_men_n49_));
  AOI210     u0027(.A0(men_men_n49_), .A1(men_men_n45_), .B0(men_men_n44_), .Y(men_men_n50_));
  NA2        u0028(.A(i_0_), .B(i_2_), .Y(men_men_n51_));
  NA2        u0029(.A(i_7_), .B(i_9_), .Y(men_men_n52_));
  NO2        u0030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  OAI210     u0031(.A0(men_men_n53_), .A1(men_men_n50_), .B0(men_men_n43_), .Y(men_men_n54_));
  NA3        u0032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n55_));
  NO2        u0033(.A(i_1_), .B(i_6_), .Y(men_men_n56_));
  NA2        u0034(.A(i_8_), .B(i_7_), .Y(men_men_n57_));
  OAI210     u0035(.A0(men_men_n57_), .A1(men_men_n56_), .B0(men_men_n55_), .Y(men_men_n58_));
  NA2        u0036(.A(men_men_n58_), .B(i_12_), .Y(men_men_n59_));
  NAi21      u0037(.An(i_2_), .B(i_7_), .Y(men_men_n60_));
  INV        u0038(.A(i_1_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_6_), .Y(men_men_n62_));
  NA3        u0040(.A(men_men_n62_), .B(men_men_n60_), .C(men_men_n29_), .Y(men_men_n63_));
  NA2        u0041(.A(i_1_), .B(i_10_), .Y(men_men_n64_));
  NO2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NAi31      u0043(.An(men_men_n65_), .B(men_men_n63_), .C(men_men_n59_), .Y(men_men_n66_));
  NA2        u0044(.A(men_men_n48_), .B(i_2_), .Y(men_men_n67_));
  AOI210     u0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n68_));
  NA2        u0046(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO2        u0047(.A(men_men_n69_), .B(men_men_n25_), .Y(men_men_n70_));
  INV        u0048(.A(i_0_), .Y(men_men_n71_));
  NAi21      u0049(.An(i_5_), .B(i_10_), .Y(men_men_n72_));
  NA2        u0050(.A(i_5_), .B(i_9_), .Y(men_men_n73_));
  AOI210     u0051(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n71_), .Y(men_men_n74_));
  NO2        u0052(.A(men_men_n74_), .B(men_men_n70_), .Y(men_men_n75_));
  OAI210     u0053(.A0(men_men_n68_), .A1(men_men_n67_), .B0(men_men_n75_), .Y(men_men_n76_));
  OAI210     u0054(.A0(men_men_n76_), .A1(men_men_n66_), .B0(i_0_), .Y(men_men_n77_));
  NA2        u0055(.A(i_12_), .B(i_5_), .Y(men_men_n78_));
  NA2        u0056(.A(i_2_), .B(i_8_), .Y(men_men_n79_));
  NO2        u0057(.A(men_men_n79_), .B(men_men_n56_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_9_), .Y(men_men_n81_));
  NO2        u0059(.A(i_3_), .B(i_7_), .Y(men_men_n82_));
  NO3        u0060(.A(men_men_n82_), .B(men_men_n81_), .C(men_men_n61_), .Y(men_men_n83_));
  INV        u0061(.A(i_6_), .Y(men_men_n84_));
  OR4        u0062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n85_));
  INV        u0063(.A(men_men_n85_), .Y(men_men_n86_));
  NO2        u0064(.A(i_2_), .B(i_7_), .Y(men_men_n87_));
  AOI210     u0065(.A0(men_men_n86_), .A1(men_men_n84_), .B0(men_men_n87_), .Y(men_men_n88_));
  OAI210     u0066(.A0(men_men_n83_), .A1(men_men_n80_), .B0(men_men_n88_), .Y(men_men_n89_));
  NAi21      u0067(.An(i_6_), .B(i_10_), .Y(men_men_n90_));
  NA2        u0068(.A(i_6_), .B(i_9_), .Y(men_men_n91_));
  AOI210     u0069(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n61_), .Y(men_men_n92_));
  NA2        u0070(.A(i_2_), .B(i_6_), .Y(men_men_n93_));
  NO3        u0071(.A(men_men_n93_), .B(men_men_n47_), .C(men_men_n25_), .Y(men_men_n94_));
  NO2        u0072(.A(men_men_n94_), .B(men_men_n92_), .Y(men_men_n95_));
  AOI210     u0073(.A0(men_men_n95_), .A1(men_men_n89_), .B0(men_men_n78_), .Y(men_men_n96_));
  AN3        u0074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n97_));
  NAi21      u0075(.An(i_6_), .B(i_11_), .Y(men_men_n98_));
  NO2        u0076(.A(i_5_), .B(i_8_), .Y(men_men_n99_));
  NOi21      u0077(.An(men_men_n99_), .B(men_men_n98_), .Y(men_men_n100_));
  AOI220     u0078(.A0(men_men_n100_), .A1(men_men_n60_), .B0(men_men_n97_), .B1(men_men_n30_), .Y(men_men_n101_));
  INV        u0079(.A(i_7_), .Y(men_men_n102_));
  NA2        u0080(.A(men_men_n44_), .B(men_men_n102_), .Y(men_men_n103_));
  NO2        u0081(.A(i_0_), .B(i_5_), .Y(men_men_n104_));
  NO2        u0082(.A(men_men_n104_), .B(men_men_n84_), .Y(men_men_n105_));
  NA2        u0083(.A(i_12_), .B(i_3_), .Y(men_men_n106_));
  INV        u0084(.A(men_men_n106_), .Y(men_men_n107_));
  NA3        u0085(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n103_), .Y(men_men_n108_));
  NAi21      u0086(.An(i_7_), .B(i_11_), .Y(men_men_n109_));
  NO3        u0087(.A(men_men_n109_), .B(men_men_n90_), .C(men_men_n51_), .Y(men_men_n110_));
  AN2        u0088(.A(i_2_), .B(i_10_), .Y(men_men_n111_));
  NO2        u0089(.A(men_men_n111_), .B(i_7_), .Y(men_men_n112_));
  OR2        u0090(.A(men_men_n78_), .B(men_men_n56_), .Y(men_men_n113_));
  NO2        u0091(.A(i_8_), .B(men_men_n102_), .Y(men_men_n114_));
  NO3        u0092(.A(men_men_n114_), .B(men_men_n113_), .C(men_men_n112_), .Y(men_men_n115_));
  NA2        u0093(.A(i_12_), .B(i_7_), .Y(men_men_n116_));
  NO2        u0094(.A(men_men_n61_), .B(men_men_n26_), .Y(men_men_n117_));
  NA2        u0095(.A(men_men_n117_), .B(i_0_), .Y(men_men_n118_));
  NA2        u0096(.A(i_11_), .B(i_12_), .Y(men_men_n119_));
  OAI210     u0097(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n119_), .Y(men_men_n120_));
  NO2        u0098(.A(men_men_n120_), .B(men_men_n115_), .Y(men_men_n121_));
  NAi41      u0099(.An(men_men_n110_), .B(men_men_n121_), .C(men_men_n108_), .D(men_men_n101_), .Y(men_men_n122_));
  NOi21      u0100(.An(i_1_), .B(i_5_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n123_), .B(i_11_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n102_), .B(men_men_n35_), .Y(men_men_n125_));
  NA2        u0103(.A(i_7_), .B(men_men_n25_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n126_), .B(men_men_n125_), .Y(men_men_n127_));
  NO2        u0105(.A(men_men_n127_), .B(men_men_n44_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n129_));
  NAi21      u0107(.An(i_3_), .B(i_8_), .Y(men_men_n130_));
  NA2        u0108(.A(men_men_n130_), .B(men_men_n60_), .Y(men_men_n131_));
  NOi31      u0109(.An(men_men_n131_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n132_));
  NO2        u0110(.A(i_1_), .B(men_men_n84_), .Y(men_men_n133_));
  NO2        u0111(.A(i_6_), .B(i_5_), .Y(men_men_n134_));
  NA2        u0112(.A(men_men_n134_), .B(i_3_), .Y(men_men_n135_));
  AO210      u0113(.A0(men_men_n135_), .A1(men_men_n45_), .B0(men_men_n133_), .Y(men_men_n136_));
  OAI220     u0114(.A0(men_men_n136_), .A1(men_men_n109_), .B0(men_men_n132_), .B1(men_men_n124_), .Y(men_men_n137_));
  NO3        u0115(.A(men_men_n137_), .B(men_men_n122_), .C(men_men_n96_), .Y(men_men_n138_));
  NA3        u0116(.A(men_men_n138_), .B(men_men_n77_), .C(men_men_n54_), .Y(men2));
  NO2        u0117(.A(men_men_n61_), .B(men_men_n35_), .Y(men_men_n140_));
  NA2        u0118(.A(i_6_), .B(men_men_n25_), .Y(men_men_n141_));
  NA3        u0119(.A(men_men_n75_), .B(men_men_n67_), .C(men_men_n26_), .Y(men0));
  AN2        u0120(.A(i_8_), .B(i_7_), .Y(men_men_n143_));
  NA2        u0121(.A(men_men_n143_), .B(i_6_), .Y(men_men_n144_));
  NO2        u0122(.A(i_12_), .B(i_13_), .Y(men_men_n145_));
  NAi21      u0123(.An(i_5_), .B(i_11_), .Y(men_men_n146_));
  NOi21      u0124(.An(men_men_n145_), .B(men_men_n146_), .Y(men_men_n147_));
  NO2        u0125(.A(i_0_), .B(i_1_), .Y(men_men_n148_));
  NA2        u0126(.A(i_2_), .B(i_3_), .Y(men_men_n149_));
  NO2        u0127(.A(men_men_n149_), .B(i_4_), .Y(men_men_n150_));
  NA3        u0128(.A(men_men_n150_), .B(men_men_n148_), .C(men_men_n147_), .Y(men_men_n151_));
  OR2        u0129(.A(men_men_n151_), .B(men_men_n25_), .Y(men_men_n152_));
  AN2        u0130(.A(men_men_n145_), .B(men_men_n81_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n153_), .B(men_men_n27_), .Y(men_men_n154_));
  NA2        u0132(.A(i_1_), .B(i_5_), .Y(men_men_n155_));
  NO2        u0133(.A(men_men_n71_), .B(men_men_n44_), .Y(men_men_n156_));
  NA2        u0134(.A(men_men_n156_), .B(men_men_n34_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n155_), .C(men_men_n154_), .Y(men_men_n158_));
  OR2        u0136(.A(i_0_), .B(i_1_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n159_), .B(men_men_n78_), .C(i_13_), .Y(men_men_n160_));
  NAi32      u0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n161_));
  NAi21      u0139(.An(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NOi21      u0140(.An(i_4_), .B(i_10_), .Y(men_men_n163_));
  NA2        u0141(.A(men_men_n163_), .B(men_men_n37_), .Y(men_men_n164_));
  NO2        u0142(.A(i_3_), .B(i_5_), .Y(men_men_n165_));
  NO3        u0143(.A(men_men_n71_), .B(i_2_), .C(i_1_), .Y(men_men_n166_));
  NA2        u0144(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  OAI210     u0145(.A0(men_men_n167_), .A1(men_men_n164_), .B0(men_men_n162_), .Y(men_men_n168_));
  NO2        u0146(.A(men_men_n168_), .B(men_men_n158_), .Y(men_men_n169_));
  AOI210     u0147(.A0(men_men_n169_), .A1(men_men_n152_), .B0(men_men_n144_), .Y(men_men_n170_));
  NA3        u0148(.A(men_men_n71_), .B(men_men_n44_), .C(i_1_), .Y(men_men_n171_));
  NA2        u0149(.A(i_3_), .B(men_men_n46_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_4_), .B(i_9_), .Y(men_men_n173_));
  NOi21      u0151(.An(i_11_), .B(i_13_), .Y(men_men_n174_));
  NA2        u0152(.A(men_men_n174_), .B(men_men_n173_), .Y(men_men_n175_));
  OR2        u0153(.A(men_men_n175_), .B(men_men_n172_), .Y(men_men_n176_));
  NO2        u0154(.A(i_4_), .B(i_5_), .Y(men_men_n177_));
  NAi21      u0155(.An(i_12_), .B(i_11_), .Y(men_men_n178_));
  NO2        u0156(.A(men_men_n178_), .B(i_13_), .Y(men_men_n179_));
  NA3        u0157(.A(men_men_n179_), .B(men_men_n177_), .C(men_men_n81_), .Y(men_men_n180_));
  AOI210     u0158(.A0(men_men_n180_), .A1(men_men_n176_), .B0(men_men_n171_), .Y(men_men_n181_));
  NO2        u0159(.A(men_men_n71_), .B(men_men_n61_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n182_), .B(men_men_n44_), .Y(men_men_n183_));
  NA2        u0161(.A(men_men_n34_), .B(i_5_), .Y(men_men_n184_));
  NAi31      u0162(.An(men_men_n184_), .B(men_men_n153_), .C(i_11_), .Y(men_men_n185_));
  NA2        u0163(.A(i_3_), .B(i_5_), .Y(men_men_n186_));
  OR2        u0164(.A(men_men_n186_), .B(men_men_n175_), .Y(men_men_n187_));
  AOI210     u0165(.A0(men_men_n187_), .A1(men_men_n185_), .B0(men_men_n183_), .Y(men_men_n188_));
  NO2        u0166(.A(men_men_n71_), .B(i_5_), .Y(men_men_n189_));
  NO2        u0167(.A(i_13_), .B(i_10_), .Y(men_men_n190_));
  NA3        u0168(.A(men_men_n190_), .B(men_men_n189_), .C(men_men_n42_), .Y(men_men_n191_));
  NO2        u0169(.A(i_2_), .B(i_1_), .Y(men_men_n192_));
  NA2        u0170(.A(men_men_n192_), .B(i_3_), .Y(men_men_n193_));
  NAi21      u0171(.An(i_4_), .B(i_12_), .Y(men_men_n194_));
  NO4        u0172(.A(men_men_n194_), .B(men_men_n193_), .C(men_men_n191_), .D(men_men_n25_), .Y(men_men_n195_));
  NO3        u0173(.A(men_men_n195_), .B(men_men_n188_), .C(men_men_n181_), .Y(men_men_n196_));
  INV        u0174(.A(i_8_), .Y(men_men_n197_));
  NO2        u0175(.A(men_men_n197_), .B(i_7_), .Y(men_men_n198_));
  NA2        u0176(.A(men_men_n198_), .B(i_6_), .Y(men_men_n199_));
  NO3        u0177(.A(i_3_), .B(men_men_n84_), .C(men_men_n46_), .Y(men_men_n200_));
  NA2        u0178(.A(men_men_n200_), .B(men_men_n114_), .Y(men_men_n201_));
  NO3        u0179(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n202_));
  NA3        u0180(.A(men_men_n202_), .B(men_men_n37_), .C(men_men_n42_), .Y(men_men_n203_));
  NO3        u0181(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n204_));
  OAI210     u0182(.A0(men_men_n97_), .A1(i_12_), .B0(men_men_n204_), .Y(men_men_n205_));
  AOI210     u0183(.A0(men_men_n205_), .A1(men_men_n203_), .B0(men_men_n201_), .Y(men_men_n206_));
  NO2        u0184(.A(i_3_), .B(i_8_), .Y(men_men_n207_));
  NO3        u0185(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n208_));
  NA3        u0186(.A(men_men_n208_), .B(men_men_n207_), .C(men_men_n37_), .Y(men_men_n209_));
  NO2        u0187(.A(men_men_n104_), .B(men_men_n56_), .Y(men_men_n210_));
  NA2        u0188(.A(men_men_n210_), .B(men_men_n159_), .Y(men_men_n211_));
  NO2        u0189(.A(i_13_), .B(i_9_), .Y(men_men_n212_));
  NA3        u0190(.A(men_men_n212_), .B(i_6_), .C(men_men_n197_), .Y(men_men_n213_));
  NAi21      u0191(.An(i_12_), .B(i_3_), .Y(men_men_n214_));
  OR2        u0192(.A(men_men_n214_), .B(men_men_n213_), .Y(men_men_n215_));
  NO2        u0193(.A(men_men_n42_), .B(i_5_), .Y(men_men_n216_));
  NO3        u0194(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n217_));
  NA3        u0195(.A(men_men_n217_), .B(men_men_n216_), .C(i_10_), .Y(men_men_n218_));
  OAI220     u0196(.A0(men_men_n218_), .A1(men_men_n215_), .B0(men_men_n211_), .B1(men_men_n209_), .Y(men_men_n219_));
  AOI210     u0197(.A0(men_men_n219_), .A1(i_7_), .B0(men_men_n206_), .Y(men_men_n220_));
  OAI220     u0198(.A0(men_men_n220_), .A1(i_4_), .B0(men_men_n199_), .B1(men_men_n196_), .Y(men_men_n221_));
  NAi21      u0199(.An(i_12_), .B(i_7_), .Y(men_men_n222_));
  NA3        u0200(.A(i_13_), .B(men_men_n197_), .C(i_10_), .Y(men_men_n223_));
  NO2        u0201(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  NA2        u0202(.A(i_0_), .B(i_5_), .Y(men_men_n225_));
  NA2        u0203(.A(men_men_n225_), .B(men_men_n105_), .Y(men_men_n226_));
  OAI220     u0204(.A0(men_men_n226_), .A1(men_men_n193_), .B0(men_men_n183_), .B1(men_men_n135_), .Y(men_men_n227_));
  NAi31      u0205(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n228_));
  NO2        u0206(.A(men_men_n34_), .B(i_13_), .Y(men_men_n229_));
  NO2        u0207(.A(men_men_n71_), .B(men_men_n26_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n44_), .B(men_men_n61_), .Y(men_men_n231_));
  NA3        u0209(.A(men_men_n231_), .B(men_men_n230_), .C(men_men_n229_), .Y(men_men_n232_));
  INV        u0210(.A(i_13_), .Y(men_men_n233_));
  NO2        u0211(.A(i_12_), .B(men_men_n233_), .Y(men_men_n234_));
  NA3        u0212(.A(men_men_n234_), .B(men_men_n202_), .C(men_men_n200_), .Y(men_men_n235_));
  OAI210     u0213(.A0(men_men_n232_), .A1(men_men_n228_), .B0(men_men_n235_), .Y(men_men_n236_));
  AOI220     u0214(.A0(men_men_n236_), .A1(men_men_n143_), .B0(men_men_n227_), .B1(men_men_n224_), .Y(men_men_n237_));
  NO2        u0215(.A(i_12_), .B(men_men_n35_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n186_), .B(i_4_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  OR2        u0218(.A(i_8_), .B(i_7_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n241_), .B(men_men_n84_), .Y(men_men_n242_));
  NO2        u0220(.A(men_men_n51_), .B(i_1_), .Y(men_men_n243_));
  NA2        u0221(.A(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  INV        u0222(.A(i_12_), .Y(men_men_n245_));
  NO2        u0223(.A(men_men_n42_), .B(men_men_n245_), .Y(men_men_n246_));
  NO3        u0224(.A(men_men_n34_), .B(i_8_), .C(i_10_), .Y(men_men_n247_));
  NA2        u0225(.A(i_2_), .B(i_1_), .Y(men_men_n248_));
  NO2        u0226(.A(men_men_n244_), .B(men_men_n240_), .Y(men_men_n249_));
  NO3        u0227(.A(i_11_), .B(i_7_), .C(men_men_n35_), .Y(men_men_n250_));
  NAi21      u0228(.An(i_4_), .B(i_3_), .Y(men_men_n251_));
  NO2        u0229(.A(men_men_n251_), .B(men_men_n73_), .Y(men_men_n252_));
  NO2        u0230(.A(i_0_), .B(i_6_), .Y(men_men_n253_));
  NOi41      u0231(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n254_));
  NA2        u0232(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NO2        u0233(.A(men_men_n248_), .B(men_men_n186_), .Y(men_men_n256_));
  NAi21      u0234(.An(men_men_n255_), .B(men_men_n256_), .Y(men_men_n257_));
  INV        u0235(.A(men_men_n257_), .Y(men_men_n258_));
  AOI220     u0236(.A0(men_men_n258_), .A1(men_men_n37_), .B0(men_men_n249_), .B1(men_men_n212_), .Y(men_men_n259_));
  NO2        u0237(.A(i_11_), .B(men_men_n233_), .Y(men_men_n260_));
  NOi21      u0238(.An(i_1_), .B(i_6_), .Y(men_men_n261_));
  NAi21      u0239(.An(i_3_), .B(i_7_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n245_), .B(i_9_), .Y(men_men_n263_));
  OR4        u0241(.A(men_men_n263_), .B(men_men_n262_), .C(men_men_n261_), .D(men_men_n189_), .Y(men_men_n264_));
  NO2        u0242(.A(men_men_n46_), .B(men_men_n25_), .Y(men_men_n265_));
  NO2        u0243(.A(i_12_), .B(i_3_), .Y(men_men_n266_));
  NA2        u0244(.A(men_men_n71_), .B(i_5_), .Y(men_men_n267_));
  NA2        u0245(.A(i_3_), .B(i_9_), .Y(men_men_n268_));
  NAi21      u0246(.An(i_7_), .B(i_10_), .Y(men_men_n269_));
  NO2        u0247(.A(men_men_n269_), .B(men_men_n268_), .Y(men_men_n270_));
  NA3        u0248(.A(men_men_n270_), .B(men_men_n267_), .C(men_men_n62_), .Y(men_men_n271_));
  NA2        u0249(.A(men_men_n271_), .B(men_men_n264_), .Y(men_men_n272_));
  NA3        u0250(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n273_));
  INV        u0251(.A(men_men_n144_), .Y(men_men_n274_));
  NA2        u0252(.A(men_men_n245_), .B(i_13_), .Y(men_men_n275_));
  NO2        u0253(.A(men_men_n275_), .B(men_men_n73_), .Y(men_men_n276_));
  AOI220     u0254(.A0(men_men_n276_), .A1(men_men_n274_), .B0(men_men_n272_), .B1(men_men_n260_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n241_), .B(men_men_n35_), .Y(men_men_n278_));
  NA2        u0256(.A(i_12_), .B(i_6_), .Y(men_men_n279_));
  OR2        u0257(.A(i_13_), .B(i_9_), .Y(men_men_n280_));
  NO3        u0258(.A(men_men_n280_), .B(men_men_n279_), .C(men_men_n46_), .Y(men_men_n281_));
  NO2        u0259(.A(men_men_n251_), .B(i_2_), .Y(men_men_n282_));
  NA3        u0260(.A(men_men_n282_), .B(men_men_n281_), .C(men_men_n42_), .Y(men_men_n283_));
  NA2        u0261(.A(men_men_n260_), .B(i_9_), .Y(men_men_n284_));
  NA3        u0262(.A(men_men_n267_), .B(men_men_n159_), .C(men_men_n62_), .Y(men_men_n285_));
  OAI210     u0263(.A0(men_men_n285_), .A1(men_men_n284_), .B0(men_men_n283_), .Y(men_men_n286_));
  NA2        u0264(.A(men_men_n156_), .B(men_men_n61_), .Y(men_men_n287_));
  NO3        u0265(.A(i_11_), .B(men_men_n233_), .C(men_men_n25_), .Y(men_men_n288_));
  NO2        u0266(.A(men_men_n262_), .B(i_8_), .Y(men_men_n289_));
  NO2        u0267(.A(i_6_), .B(men_men_n46_), .Y(men_men_n290_));
  NA3        u0268(.A(men_men_n290_), .B(men_men_n289_), .C(men_men_n288_), .Y(men_men_n291_));
  NO3        u0269(.A(men_men_n26_), .B(men_men_n84_), .C(i_5_), .Y(men_men_n292_));
  NA3        u0270(.A(men_men_n292_), .B(men_men_n278_), .C(men_men_n234_), .Y(men_men_n293_));
  AOI210     u0271(.A0(men_men_n293_), .A1(men_men_n291_), .B0(men_men_n287_), .Y(men_men_n294_));
  AOI210     u0272(.A0(men_men_n286_), .A1(men_men_n278_), .B0(men_men_n294_), .Y(men_men_n295_));
  NA4        u0273(.A(men_men_n295_), .B(men_men_n277_), .C(men_men_n259_), .D(men_men_n237_), .Y(men_men_n296_));
  NO3        u0274(.A(i_12_), .B(men_men_n233_), .C(men_men_n35_), .Y(men_men_n297_));
  INV        u0275(.A(men_men_n297_), .Y(men_men_n298_));
  NA2        u0276(.A(i_8_), .B(men_men_n102_), .Y(men_men_n299_));
  NOi21      u0277(.An(men_men_n165_), .B(men_men_n84_), .Y(men_men_n300_));
  NO3        u0278(.A(i_0_), .B(men_men_n44_), .C(i_1_), .Y(men_men_n301_));
  AOI220     u0279(.A0(men_men_n301_), .A1(men_men_n200_), .B0(men_men_n300_), .B1(men_men_n243_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n302_), .B(men_men_n299_), .Y(men_men_n303_));
  NO3        u0281(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n248_), .B(i_0_), .Y(men_men_n305_));
  AOI220     u0283(.A0(men_men_n305_), .A1(men_men_n198_), .B0(men_men_n304_), .B1(men_men_n143_), .Y(men_men_n306_));
  NA2        u0284(.A(men_men_n290_), .B(men_men_n26_), .Y(men_men_n307_));
  NO2        u0285(.A(men_men_n307_), .B(men_men_n306_), .Y(men_men_n308_));
  NA2        u0286(.A(i_0_), .B(i_1_), .Y(men_men_n309_));
  NO2        u0287(.A(men_men_n309_), .B(i_2_), .Y(men_men_n310_));
  NO2        u0288(.A(men_men_n57_), .B(i_6_), .Y(men_men_n311_));
  NA3        u0289(.A(men_men_n311_), .B(men_men_n310_), .C(men_men_n165_), .Y(men_men_n312_));
  OAI210     u0290(.A0(men_men_n167_), .A1(men_men_n144_), .B0(men_men_n312_), .Y(men_men_n313_));
  NO3        u0291(.A(men_men_n313_), .B(men_men_n308_), .C(men_men_n303_), .Y(men_men_n314_));
  NO2        u0292(.A(i_3_), .B(i_10_), .Y(men_men_n315_));
  NA3        u0293(.A(men_men_n315_), .B(men_men_n37_), .C(men_men_n42_), .Y(men_men_n316_));
  NO2        u0294(.A(i_2_), .B(men_men_n102_), .Y(men_men_n317_));
  NA2        u0295(.A(i_1_), .B(men_men_n34_), .Y(men_men_n318_));
  NO2        u0296(.A(men_men_n318_), .B(i_8_), .Y(men_men_n319_));
  NOi21      u0297(.An(men_men_n225_), .B(men_men_n104_), .Y(men_men_n320_));
  NA3        u0298(.A(men_men_n320_), .B(men_men_n319_), .C(men_men_n317_), .Y(men_men_n321_));
  AN2        u0299(.A(i_3_), .B(i_10_), .Y(men_men_n322_));
  NA4        u0300(.A(men_men_n322_), .B(men_men_n202_), .C(men_men_n179_), .D(men_men_n177_), .Y(men_men_n323_));
  NO2        u0301(.A(i_5_), .B(men_men_n35_), .Y(men_men_n324_));
  NO2        u0302(.A(men_men_n44_), .B(men_men_n26_), .Y(men_men_n325_));
  OR2        u0303(.A(men_men_n321_), .B(men_men_n316_), .Y(men_men_n326_));
  OAI220     u0304(.A0(men_men_n326_), .A1(i_6_), .B0(men_men_n314_), .B1(men_men_n298_), .Y(men_men_n327_));
  NO4        u0305(.A(men_men_n327_), .B(men_men_n296_), .C(men_men_n221_), .D(men_men_n170_), .Y(men_men_n328_));
  NO3        u0306(.A(men_men_n42_), .B(i_13_), .C(i_9_), .Y(men_men_n329_));
  NO2        u0307(.A(men_men_n57_), .B(men_men_n84_), .Y(men_men_n330_));
  NA2        u0308(.A(men_men_n305_), .B(men_men_n330_), .Y(men_men_n331_));
  NO3        u0309(.A(i_6_), .B(men_men_n197_), .C(i_7_), .Y(men_men_n332_));
  NA2        u0310(.A(men_men_n332_), .B(men_men_n202_), .Y(men_men_n333_));
  AOI210     u0311(.A0(men_men_n333_), .A1(men_men_n331_), .B0(men_men_n172_), .Y(men_men_n334_));
  NO2        u0312(.A(i_2_), .B(i_3_), .Y(men_men_n335_));
  OR2        u0313(.A(i_0_), .B(i_5_), .Y(men_men_n336_));
  NA2        u0314(.A(men_men_n225_), .B(men_men_n336_), .Y(men_men_n337_));
  NA4        u0315(.A(men_men_n337_), .B(men_men_n242_), .C(men_men_n335_), .D(i_1_), .Y(men_men_n338_));
  NA3        u0316(.A(men_men_n305_), .B(men_men_n300_), .C(men_men_n114_), .Y(men_men_n339_));
  NAi21      u0317(.An(i_8_), .B(i_7_), .Y(men_men_n340_));
  NO2        u0318(.A(men_men_n340_), .B(i_6_), .Y(men_men_n341_));
  NO2        u0319(.A(men_men_n159_), .B(men_men_n44_), .Y(men_men_n342_));
  NA3        u0320(.A(men_men_n342_), .B(men_men_n341_), .C(men_men_n165_), .Y(men_men_n343_));
  NA3        u0321(.A(men_men_n343_), .B(men_men_n339_), .C(men_men_n338_), .Y(men_men_n344_));
  OAI210     u0322(.A0(men_men_n344_), .A1(men_men_n334_), .B0(i_4_), .Y(men_men_n345_));
  NO2        u0323(.A(i_12_), .B(i_10_), .Y(men_men_n346_));
  NOi21      u0324(.An(i_5_), .B(i_0_), .Y(men_men_n347_));
  AOI210     u0325(.A0(i_2_), .A1(men_men_n46_), .B0(men_men_n102_), .Y(men_men_n348_));
  NO4        u0326(.A(men_men_n348_), .B(men_men_n318_), .C(men_men_n347_), .D(men_men_n130_), .Y(men_men_n349_));
  NA4        u0327(.A(men_men_n82_), .B(men_men_n34_), .C(men_men_n84_), .D(i_8_), .Y(men_men_n350_));
  NA2        u0328(.A(men_men_n349_), .B(men_men_n346_), .Y(men_men_n351_));
  NO2        u0329(.A(i_6_), .B(i_8_), .Y(men_men_n352_));
  NOi21      u0330(.An(i_0_), .B(i_2_), .Y(men_men_n353_));
  AN2        u0331(.A(men_men_n353_), .B(men_men_n352_), .Y(men_men_n354_));
  NO2        u0332(.A(i_1_), .B(i_7_), .Y(men_men_n355_));
  AO220      u0333(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n341_), .B1(men_men_n243_), .Y(men_men_n356_));
  NA3        u0334(.A(men_men_n356_), .B(men_men_n39_), .C(i_5_), .Y(men_men_n357_));
  NA3        u0335(.A(men_men_n357_), .B(men_men_n351_), .C(men_men_n345_), .Y(men_men_n358_));
  NO3        u0336(.A(men_men_n241_), .B(men_men_n44_), .C(i_1_), .Y(men_men_n359_));
  NO3        u0337(.A(men_men_n340_), .B(i_2_), .C(i_1_), .Y(men_men_n360_));
  OAI210     u0338(.A0(men_men_n360_), .A1(men_men_n359_), .B0(i_6_), .Y(men_men_n361_));
  NA3        u0339(.A(men_men_n261_), .B(men_men_n317_), .C(men_men_n197_), .Y(men_men_n362_));
  AOI210     u0340(.A0(men_men_n362_), .A1(men_men_n361_), .B0(men_men_n337_), .Y(men_men_n363_));
  NOi21      u0341(.An(men_men_n155_), .B(men_men_n105_), .Y(men_men_n364_));
  NO2        u0342(.A(men_men_n364_), .B(men_men_n126_), .Y(men_men_n365_));
  OAI210     u0343(.A0(men_men_n365_), .A1(men_men_n363_), .B0(i_3_), .Y(men_men_n366_));
  INV        u0344(.A(men_men_n82_), .Y(men_men_n367_));
  NO2        u0345(.A(men_men_n309_), .B(men_men_n79_), .Y(men_men_n368_));
  NA2        u0346(.A(men_men_n368_), .B(men_men_n134_), .Y(men_men_n369_));
  NO2        u0347(.A(men_men_n93_), .B(men_men_n197_), .Y(men_men_n370_));
  NA3        u0348(.A(men_men_n320_), .B(men_men_n370_), .C(men_men_n61_), .Y(men_men_n371_));
  AOI210     u0349(.A0(men_men_n371_), .A1(men_men_n369_), .B0(men_men_n367_), .Y(men_men_n372_));
  NO2        u0350(.A(men_men_n197_), .B(i_9_), .Y(men_men_n373_));
  NA3        u0351(.A(men_men_n373_), .B(men_men_n210_), .C(men_men_n159_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n374_), .B(men_men_n44_), .Y(men_men_n375_));
  NO3        u0353(.A(men_men_n375_), .B(men_men_n372_), .C(men_men_n308_), .Y(men_men_n376_));
  AOI210     u0354(.A0(men_men_n376_), .A1(men_men_n366_), .B0(men_men_n164_), .Y(men_men_n377_));
  AOI210     u0355(.A0(men_men_n358_), .A1(men_men_n329_), .B0(men_men_n377_), .Y(men_men_n378_));
  NOi32      u0356(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n379_));
  INV        u0357(.A(men_men_n379_), .Y(men_men_n380_));
  NAi21      u0358(.An(i_0_), .B(i_6_), .Y(men_men_n381_));
  NAi21      u0359(.An(i_1_), .B(i_5_), .Y(men_men_n382_));
  NA2        u0360(.A(men_men_n382_), .B(men_men_n381_), .Y(men_men_n383_));
  NA2        u0361(.A(men_men_n383_), .B(men_men_n25_), .Y(men_men_n384_));
  OAI210     u0362(.A0(men_men_n384_), .A1(men_men_n161_), .B0(men_men_n255_), .Y(men_men_n385_));
  NAi41      u0363(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n386_));
  OAI220     u0364(.A0(men_men_n386_), .A1(men_men_n382_), .B0(men_men_n228_), .B1(men_men_n161_), .Y(men_men_n387_));
  AOI210     u0365(.A0(men_men_n386_), .A1(men_men_n161_), .B0(men_men_n159_), .Y(men_men_n388_));
  NOi32      u0366(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n389_));
  NAi21      u0367(.An(i_6_), .B(i_1_), .Y(men_men_n390_));
  NA3        u0368(.A(men_men_n390_), .B(men_men_n389_), .C(men_men_n44_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n391_), .B(i_0_), .Y(men_men_n392_));
  OR3        u0370(.A(men_men_n392_), .B(men_men_n388_), .C(men_men_n387_), .Y(men_men_n393_));
  NO2        u0371(.A(i_1_), .B(men_men_n102_), .Y(men_men_n394_));
  NAi21      u0372(.An(i_3_), .B(i_4_), .Y(men_men_n395_));
  NO2        u0373(.A(men_men_n395_), .B(i_9_), .Y(men_men_n396_));
  AN2        u0374(.A(i_6_), .B(i_7_), .Y(men_men_n397_));
  OAI210     u0375(.A0(men_men_n397_), .A1(men_men_n394_), .B0(men_men_n396_), .Y(men_men_n398_));
  NA2        u0376(.A(i_2_), .B(i_7_), .Y(men_men_n399_));
  NO2        u0377(.A(men_men_n395_), .B(i_10_), .Y(men_men_n400_));
  NA3        u0378(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n253_), .Y(men_men_n401_));
  AOI210     u0379(.A0(men_men_n401_), .A1(men_men_n398_), .B0(men_men_n189_), .Y(men_men_n402_));
  AOI210     u0380(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n403_));
  OAI210     u0381(.A0(men_men_n403_), .A1(men_men_n192_), .B0(men_men_n400_), .Y(men_men_n404_));
  AOI220     u0382(.A0(men_men_n400_), .A1(men_men_n355_), .B0(men_men_n247_), .B1(men_men_n192_), .Y(men_men_n405_));
  AOI210     u0383(.A0(men_men_n405_), .A1(men_men_n404_), .B0(i_5_), .Y(men_men_n406_));
  NO4        u0384(.A(men_men_n406_), .B(men_men_n402_), .C(men_men_n393_), .D(men_men_n385_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n407_), .B(men_men_n380_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n57_), .B(men_men_n25_), .Y(men_men_n409_));
  AN2        u0387(.A(i_12_), .B(i_5_), .Y(men_men_n410_));
  NO2        u0388(.A(i_4_), .B(men_men_n26_), .Y(men_men_n411_));
  NA2        u0389(.A(men_men_n411_), .B(men_men_n410_), .Y(men_men_n412_));
  NO2        u0390(.A(i_11_), .B(i_6_), .Y(men_men_n413_));
  NA3        u0391(.A(men_men_n413_), .B(men_men_n342_), .C(men_men_n233_), .Y(men_men_n414_));
  NO2        u0392(.A(men_men_n414_), .B(men_men_n412_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n251_), .B(i_5_), .Y(men_men_n416_));
  NO2        u0394(.A(i_5_), .B(i_10_), .Y(men_men_n417_));
  AOI220     u0395(.A0(men_men_n417_), .A1(men_men_n282_), .B0(men_men_n416_), .B1(men_men_n202_), .Y(men_men_n418_));
  NA2        u0396(.A(men_men_n145_), .B(men_men_n43_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n419_), .B(men_men_n418_), .Y(men_men_n420_));
  OAI210     u0398(.A0(men_men_n420_), .A1(men_men_n415_), .B0(men_men_n409_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n35_), .B(men_men_n25_), .Y(men_men_n422_));
  NO2        u0400(.A(men_men_n151_), .B(men_men_n84_), .Y(men_men_n423_));
  OAI210     u0401(.A0(men_men_n423_), .A1(men_men_n415_), .B0(men_men_n422_), .Y(men_men_n424_));
  NO3        u0402(.A(men_men_n84_), .B(men_men_n46_), .C(i_9_), .Y(men_men_n425_));
  NO2        u0403(.A(i_3_), .B(men_men_n102_), .Y(men_men_n426_));
  NO2        u0404(.A(i_11_), .B(i_12_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n417_), .B(men_men_n245_), .Y(men_men_n428_));
  NA3        u0406(.A(men_men_n114_), .B(men_men_n39_), .C(i_11_), .Y(men_men_n429_));
  OAI220     u0407(.A0(men_men_n429_), .A1(men_men_n228_), .B0(men_men_n428_), .B1(men_men_n350_), .Y(men_men_n430_));
  NAi21      u0408(.An(i_13_), .B(i_0_), .Y(men_men_n431_));
  NO2        u0409(.A(men_men_n431_), .B(men_men_n248_), .Y(men_men_n432_));
  NA2        u0410(.A(men_men_n430_), .B(men_men_n432_), .Y(men_men_n433_));
  NA3        u0411(.A(men_men_n433_), .B(men_men_n424_), .C(men_men_n421_), .Y(men_men_n434_));
  NA2        u0412(.A(men_men_n42_), .B(men_men_n233_), .Y(men_men_n435_));
  NO3        u0413(.A(i_1_), .B(i_12_), .C(men_men_n84_), .Y(men_men_n436_));
  NO2        u0414(.A(i_0_), .B(i_11_), .Y(men_men_n437_));
  AN2        u0415(.A(i_1_), .B(i_6_), .Y(men_men_n438_));
  NOi21      u0416(.An(i_2_), .B(i_12_), .Y(men_men_n439_));
  NA2        u0417(.A(men_men_n439_), .B(men_men_n438_), .Y(men_men_n440_));
  NO2        u0418(.A(men_men_n440_), .B(men_men_n1146_), .Y(men_men_n441_));
  NA2        u0419(.A(men_men_n143_), .B(i_9_), .Y(men_men_n442_));
  NO2        u0420(.A(men_men_n442_), .B(i_4_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n441_), .B(men_men_n443_), .Y(men_men_n444_));
  NAi21      u0422(.An(i_9_), .B(i_4_), .Y(men_men_n445_));
  OR2        u0423(.A(i_13_), .B(i_10_), .Y(men_men_n446_));
  NO3        u0424(.A(men_men_n446_), .B(men_men_n119_), .C(men_men_n445_), .Y(men_men_n447_));
  NO2        u0425(.A(men_men_n175_), .B(men_men_n125_), .Y(men_men_n448_));
  OR2        u0426(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n449_));
  NO2        u0427(.A(men_men_n102_), .B(men_men_n25_), .Y(men_men_n450_));
  NA2        u0428(.A(men_men_n297_), .B(men_men_n450_), .Y(men_men_n451_));
  NA2        u0429(.A(men_men_n290_), .B(men_men_n217_), .Y(men_men_n452_));
  OAI220     u0430(.A0(men_men_n452_), .A1(men_men_n449_), .B0(men_men_n451_), .B1(men_men_n364_), .Y(men_men_n453_));
  INV        u0431(.A(men_men_n453_), .Y(men_men_n454_));
  AOI210     u0432(.A0(men_men_n454_), .A1(men_men_n444_), .B0(men_men_n26_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n339_), .B(men_men_n338_), .Y(men_men_n456_));
  AOI220     u0434(.A0(men_men_n311_), .A1(men_men_n301_), .B0(men_men_n305_), .B1(men_men_n330_), .Y(men_men_n457_));
  NO2        u0435(.A(men_men_n457_), .B(men_men_n172_), .Y(men_men_n458_));
  NO2        u0436(.A(men_men_n186_), .B(men_men_n84_), .Y(men_men_n459_));
  AOI220     u0437(.A0(men_men_n459_), .A1(men_men_n310_), .B0(men_men_n292_), .B1(men_men_n217_), .Y(men_men_n460_));
  NO2        u0438(.A(men_men_n460_), .B(men_men_n299_), .Y(men_men_n461_));
  NO3        u0439(.A(men_men_n461_), .B(men_men_n458_), .C(men_men_n456_), .Y(men_men_n462_));
  NA2        u0440(.A(men_men_n200_), .B(men_men_n97_), .Y(men_men_n463_));
  NA3        u0441(.A(men_men_n342_), .B(men_men_n165_), .C(men_men_n84_), .Y(men_men_n464_));
  AOI210     u0442(.A0(men_men_n464_), .A1(men_men_n463_), .B0(men_men_n340_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n197_), .B(i_10_), .Y(men_men_n466_));
  NA3        u0444(.A(men_men_n267_), .B(men_men_n62_), .C(i_2_), .Y(men_men_n467_));
  NA2        u0445(.A(men_men_n311_), .B(men_men_n243_), .Y(men_men_n468_));
  OAI220     u0446(.A0(men_men_n468_), .A1(men_men_n186_), .B0(men_men_n467_), .B1(men_men_n466_), .Y(men_men_n469_));
  NO2        u0447(.A(i_3_), .B(men_men_n46_), .Y(men_men_n470_));
  NA3        u0448(.A(men_men_n355_), .B(men_men_n354_), .C(men_men_n470_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n332_), .B(men_men_n337_), .Y(men_men_n472_));
  OAI210     u0450(.A0(men_men_n472_), .A1(men_men_n193_), .B0(men_men_n471_), .Y(men_men_n473_));
  NO3        u0451(.A(men_men_n473_), .B(men_men_n469_), .C(men_men_n465_), .Y(men_men_n474_));
  AOI210     u0452(.A0(men_men_n474_), .A1(men_men_n462_), .B0(men_men_n284_), .Y(men_men_n475_));
  NO4        u0453(.A(men_men_n475_), .B(men_men_n455_), .C(men_men_n434_), .D(men_men_n408_), .Y(men_men_n476_));
  NO2        u0454(.A(men_men_n61_), .B(i_4_), .Y(men_men_n477_));
  NO2        u0455(.A(men_men_n71_), .B(i_13_), .Y(men_men_n478_));
  NA3        u0456(.A(men_men_n478_), .B(men_men_n477_), .C(i_2_), .Y(men_men_n479_));
  NO2        u0457(.A(i_10_), .B(i_9_), .Y(men_men_n480_));
  NAi21      u0458(.An(i_12_), .B(i_8_), .Y(men_men_n481_));
  NO2        u0459(.A(men_men_n481_), .B(i_3_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n482_), .B(men_men_n480_), .Y(men_men_n483_));
  NO2        u0461(.A(men_men_n44_), .B(i_4_), .Y(men_men_n484_));
  NA2        u0462(.A(men_men_n484_), .B(men_men_n105_), .Y(men_men_n485_));
  OAI220     u0463(.A0(men_men_n485_), .A1(men_men_n209_), .B0(men_men_n483_), .B1(men_men_n479_), .Y(men_men_n486_));
  NA2        u0464(.A(men_men_n325_), .B(i_0_), .Y(men_men_n487_));
  NO3        u0465(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n279_), .B(men_men_n98_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n490_));
  NA2        u0468(.A(i_8_), .B(i_9_), .Y(men_men_n491_));
  AOI210     u0469(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n492_));
  OR2        u0470(.A(men_men_n492_), .B(men_men_n491_), .Y(men_men_n493_));
  NA2        u0471(.A(men_men_n297_), .B(men_men_n210_), .Y(men_men_n494_));
  OAI220     u0472(.A0(men_men_n494_), .A1(men_men_n493_), .B0(men_men_n490_), .B1(men_men_n487_), .Y(men_men_n495_));
  NA2        u0473(.A(men_men_n260_), .B(men_men_n324_), .Y(men_men_n496_));
  NO3        u0474(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n497_));
  AOI210     u0475(.A0(men_men_n266_), .A1(men_men_n192_), .B0(men_men_n497_), .Y(men_men_n498_));
  NA3        u0476(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n499_));
  NA4        u0477(.A(men_men_n146_), .B(men_men_n117_), .C(men_men_n78_), .D(men_men_n23_), .Y(men_men_n500_));
  OAI220     u0478(.A0(men_men_n500_), .A1(men_men_n499_), .B0(men_men_n498_), .B1(men_men_n496_), .Y(men_men_n501_));
  NO3        u0479(.A(men_men_n501_), .B(men_men_n495_), .C(men_men_n486_), .Y(men_men_n502_));
  NA2        u0480(.A(men_men_n310_), .B(men_men_n109_), .Y(men_men_n503_));
  OR2        u0481(.A(men_men_n503_), .B(men_men_n213_), .Y(men_men_n504_));
  OA210      u0482(.A0(men_men_n374_), .A1(men_men_n102_), .B0(men_men_n312_), .Y(men_men_n505_));
  OA220      u0483(.A0(men_men_n505_), .A1(men_men_n164_), .B0(men_men_n504_), .B1(men_men_n240_), .Y(men_men_n506_));
  NA2        u0484(.A(men_men_n97_), .B(i_13_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n459_), .B(men_men_n409_), .Y(men_men_n508_));
  NO2        u0486(.A(i_2_), .B(i_13_), .Y(men_men_n509_));
  NA3        u0487(.A(men_men_n509_), .B(men_men_n163_), .C(men_men_n100_), .Y(men_men_n510_));
  OAI220     u0488(.A0(men_men_n510_), .A1(men_men_n245_), .B0(men_men_n508_), .B1(men_men_n507_), .Y(men_men_n511_));
  NO3        u0489(.A(i_4_), .B(men_men_n46_), .C(i_8_), .Y(men_men_n512_));
  NO2        u0490(.A(i_6_), .B(i_7_), .Y(men_men_n513_));
  NA2        u0491(.A(men_men_n513_), .B(men_men_n512_), .Y(men_men_n514_));
  NO2        u0492(.A(i_11_), .B(i_1_), .Y(men_men_n515_));
  NO2        u0493(.A(men_men_n71_), .B(i_3_), .Y(men_men_n516_));
  OR2        u0494(.A(i_11_), .B(i_8_), .Y(men_men_n517_));
  NOi21      u0495(.An(i_2_), .B(i_7_), .Y(men_men_n518_));
  NAi31      u0496(.An(men_men_n517_), .B(men_men_n518_), .C(men_men_n516_), .Y(men_men_n519_));
  NO2        u0497(.A(men_men_n446_), .B(i_6_), .Y(men_men_n520_));
  NA3        u0498(.A(men_men_n520_), .B(men_men_n477_), .C(men_men_n73_), .Y(men_men_n521_));
  NO2        u0499(.A(men_men_n521_), .B(men_men_n519_), .Y(men_men_n522_));
  NO2        u0500(.A(i_3_), .B(men_men_n197_), .Y(men_men_n523_));
  NO2        u0501(.A(i_6_), .B(i_10_), .Y(men_men_n524_));
  NA4        u0502(.A(men_men_n524_), .B(men_men_n329_), .C(men_men_n523_), .D(men_men_n245_), .Y(men_men_n525_));
  NO2        u0503(.A(men_men_n525_), .B(men_men_n157_), .Y(men_men_n526_));
  NA3        u0504(.A(men_men_n254_), .B(men_men_n174_), .C(men_men_n134_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n44_), .B(men_men_n42_), .Y(men_men_n528_));
  NO2        u0506(.A(men_men_n159_), .B(i_3_), .Y(men_men_n529_));
  NAi31      u0507(.An(men_men_n528_), .B(men_men_n529_), .C(men_men_n234_), .Y(men_men_n530_));
  NA3        u0508(.A(men_men_n422_), .B(men_men_n182_), .C(men_men_n150_), .Y(men_men_n531_));
  NA3        u0509(.A(men_men_n531_), .B(men_men_n530_), .C(men_men_n527_), .Y(men_men_n532_));
  NO4        u0510(.A(men_men_n532_), .B(men_men_n526_), .C(men_men_n522_), .D(men_men_n511_), .Y(men_men_n533_));
  NA2        u0511(.A(men_men_n488_), .B(men_men_n410_), .Y(men_men_n534_));
  NA2        u0512(.A(men_men_n497_), .B(men_men_n417_), .Y(men_men_n535_));
  OAI220     u0513(.A0(men_men_n535_), .A1(men_men_n232_), .B0(men_men_n534_), .B1(men_men_n55_), .Y(men_men_n536_));
  NAi21      u0514(.An(men_men_n223_), .B(men_men_n427_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n355_), .B(men_men_n225_), .Y(men_men_n538_));
  NO2        u0516(.A(men_men_n26_), .B(i_5_), .Y(men_men_n539_));
  NO2        u0517(.A(i_0_), .B(men_men_n84_), .Y(men_men_n540_));
  NA3        u0518(.A(men_men_n540_), .B(men_men_n539_), .C(men_men_n143_), .Y(men_men_n541_));
  OR3        u0519(.A(men_men_n318_), .B(men_men_n36_), .C(men_men_n44_), .Y(men_men_n542_));
  OAI220     u0520(.A0(men_men_n542_), .A1(men_men_n541_), .B0(men_men_n538_), .B1(men_men_n537_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n27_), .B(i_10_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n329_), .B(men_men_n247_), .Y(men_men_n545_));
  OAI220     u0523(.A0(men_men_n545_), .A1(men_men_n467_), .B0(men_men_n544_), .B1(men_men_n507_), .Y(men_men_n546_));
  NA4        u0524(.A(men_men_n322_), .B(men_men_n231_), .C(men_men_n71_), .D(men_men_n245_), .Y(men_men_n547_));
  NO2        u0525(.A(men_men_n547_), .B(men_men_n514_), .Y(men_men_n548_));
  NO4        u0526(.A(men_men_n548_), .B(men_men_n546_), .C(men_men_n543_), .D(men_men_n536_), .Y(men_men_n549_));
  NA4        u0527(.A(men_men_n549_), .B(men_men_n533_), .C(men_men_n506_), .D(men_men_n502_), .Y(men_men_n550_));
  NA3        u0528(.A(men_men_n322_), .B(men_men_n179_), .C(men_men_n177_), .Y(men_men_n551_));
  OAI210     u0529(.A0(men_men_n316_), .A1(men_men_n184_), .B0(men_men_n551_), .Y(men_men_n552_));
  AN2        u0530(.A(men_men_n301_), .B(men_men_n242_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n553_), .B(men_men_n552_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n124_), .B(men_men_n113_), .Y(men_men_n555_));
  AO220      u0533(.A0(men_men_n555_), .A1(men_men_n488_), .B0(men_men_n447_), .B1(i_6_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n329_), .B(men_men_n166_), .Y(men_men_n557_));
  OAI210     u0535(.A0(men_men_n557_), .A1(men_men_n240_), .B0(men_men_n323_), .Y(men_men_n558_));
  AOI220     u0536(.A0(men_men_n558_), .A1(men_men_n341_), .B0(men_men_n556_), .B1(men_men_n325_), .Y(men_men_n559_));
  NA4        u0537(.A(men_men_n478_), .B(men_men_n477_), .C(men_men_n207_), .D(i_2_), .Y(men_men_n560_));
  INV        u0538(.A(men_men_n560_), .Y(men_men_n561_));
  NA2        u0539(.A(men_men_n410_), .B(men_men_n233_), .Y(men_men_n562_));
  NA2        u0540(.A(men_men_n379_), .B(men_men_n71_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n397_), .B(men_men_n389_), .Y(men_men_n564_));
  AO210      u0542(.A0(men_men_n563_), .A1(men_men_n562_), .B0(men_men_n564_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n34_), .B(i_8_), .Y(men_men_n566_));
  INV        u0544(.A(men_men_n447_), .Y(men_men_n567_));
  NA2        u0545(.A(men_men_n567_), .B(men_men_n565_), .Y(men_men_n568_));
  AOI210     u0546(.A0(men_men_n561_), .A1(men_men_n208_), .B0(men_men_n568_), .Y(men_men_n569_));
  NA2        u0547(.A(men_men_n267_), .B(men_men_n62_), .Y(men_men_n570_));
  OAI210     u0548(.A0(i_8_), .A1(men_men_n570_), .B0(men_men_n136_), .Y(men_men_n571_));
  AOI210     u0549(.A0(men_men_n198_), .A1(i_9_), .B0(men_men_n278_), .Y(men_men_n572_));
  NO2        u0550(.A(men_men_n572_), .B(men_men_n203_), .Y(men_men_n573_));
  OR2        u0551(.A(men_men_n186_), .B(i_4_), .Y(men_men_n574_));
  NO2        u0552(.A(men_men_n574_), .B(men_men_n84_), .Y(men_men_n575_));
  AOI220     u0553(.A0(men_men_n575_), .A1(men_men_n573_), .B0(men_men_n571_), .B1(men_men_n448_), .Y(men_men_n576_));
  NA4        u0554(.A(men_men_n576_), .B(men_men_n569_), .C(men_men_n559_), .D(men_men_n554_), .Y(men_men_n577_));
  NA2        u0555(.A(men_men_n416_), .B(men_men_n310_), .Y(men_men_n578_));
  OAI210     u0556(.A0(men_men_n412_), .A1(men_men_n171_), .B0(men_men_n578_), .Y(men_men_n579_));
  NO2        u0557(.A(i_12_), .B(men_men_n197_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n580_), .B(men_men_n233_), .Y(men_men_n581_));
  NA3        u0559(.A(men_men_n524_), .B(men_men_n177_), .C(men_men_n27_), .Y(men_men_n582_));
  NO3        u0560(.A(men_men_n582_), .B(men_men_n581_), .C(men_men_n503_), .Y(men_men_n583_));
  NOi31      u0561(.An(men_men_n332_), .B(men_men_n446_), .C(men_men_n36_), .Y(men_men_n584_));
  OAI210     u0562(.A0(men_men_n584_), .A1(men_men_n583_), .B0(men_men_n579_), .Y(men_men_n585_));
  NO2        u0563(.A(i_8_), .B(i_7_), .Y(men_men_n586_));
  OAI210     u0564(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n587_));
  NA2        u0565(.A(men_men_n587_), .B(men_men_n231_), .Y(men_men_n588_));
  AOI220     u0566(.A0(men_men_n342_), .A1(men_men_n37_), .B0(men_men_n243_), .B1(men_men_n212_), .Y(men_men_n589_));
  OAI220     u0567(.A0(men_men_n589_), .A1(men_men_n574_), .B0(men_men_n588_), .B1(men_men_n251_), .Y(men_men_n590_));
  NA2        u0568(.A(men_men_n42_), .B(i_10_), .Y(men_men_n591_));
  NO2        u0569(.A(men_men_n591_), .B(i_6_), .Y(men_men_n592_));
  NA3        u0570(.A(men_men_n592_), .B(men_men_n590_), .C(men_men_n586_), .Y(men_men_n593_));
  AOI220     u0571(.A0(men_men_n459_), .A1(men_men_n342_), .B0(men_men_n256_), .B1(men_men_n253_), .Y(men_men_n594_));
  OAI220     u0572(.A0(men_men_n594_), .A1(men_men_n275_), .B0(men_men_n507_), .B1(men_men_n135_), .Y(men_men_n595_));
  NA2        u0573(.A(men_men_n595_), .B(men_men_n278_), .Y(men_men_n596_));
  NOi31      u0574(.An(men_men_n305_), .B(men_men_n316_), .C(men_men_n184_), .Y(men_men_n597_));
  NA3        u0575(.A(men_men_n322_), .B(men_men_n177_), .C(men_men_n97_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n229_), .B(men_men_n42_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n159_), .B(i_5_), .Y(men_men_n600_));
  NA3        u0578(.A(men_men_n600_), .B(men_men_n435_), .C(men_men_n335_), .Y(men_men_n601_));
  OAI210     u0579(.A0(men_men_n601_), .A1(men_men_n599_), .B0(men_men_n598_), .Y(men_men_n602_));
  OAI210     u0580(.A0(men_men_n602_), .A1(men_men_n597_), .B0(men_men_n497_), .Y(men_men_n603_));
  NA4        u0581(.A(men_men_n603_), .B(men_men_n596_), .C(men_men_n593_), .D(men_men_n585_), .Y(men_men_n604_));
  NA3        u0582(.A(men_men_n225_), .B(men_men_n69_), .C(men_men_n42_), .Y(men_men_n605_));
  NA2        u0583(.A(men_men_n297_), .B(men_men_n82_), .Y(men_men_n606_));
  AOI210     u0584(.A0(men_men_n605_), .A1(men_men_n369_), .B0(men_men_n606_), .Y(men_men_n607_));
  NA2        u0585(.A(men_men_n311_), .B(men_men_n301_), .Y(men_men_n608_));
  NO2        u0586(.A(men_men_n608_), .B(men_men_n176_), .Y(men_men_n609_));
  NA2        u0587(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n610_));
  NA2        u0588(.A(men_men_n480_), .B(men_men_n229_), .Y(men_men_n611_));
  NO2        u0589(.A(men_men_n610_), .B(men_men_n611_), .Y(men_men_n612_));
  AOI210     u0590(.A0(men_men_n390_), .A1(men_men_n44_), .B0(men_men_n394_), .Y(men_men_n613_));
  NA2        u0591(.A(i_0_), .B(men_men_n46_), .Y(men_men_n614_));
  NA3        u0592(.A(men_men_n580_), .B(men_men_n288_), .C(men_men_n614_), .Y(men_men_n615_));
  NO2        u0593(.A(men_men_n613_), .B(men_men_n615_), .Y(men_men_n616_));
  NO4        u0594(.A(men_men_n616_), .B(men_men_n612_), .C(men_men_n609_), .D(men_men_n607_), .Y(men_men_n617_));
  NO4        u0595(.A(men_men_n261_), .B(men_men_n40_), .C(i_2_), .D(men_men_n46_), .Y(men_men_n618_));
  NO3        u0596(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n619_));
  NO2        u0597(.A(men_men_n241_), .B(men_men_n34_), .Y(men_men_n620_));
  AN2        u0598(.A(men_men_n620_), .B(men_men_n619_), .Y(men_men_n621_));
  OA210      u0599(.A0(men_men_n621_), .A1(men_men_n618_), .B0(men_men_n379_), .Y(men_men_n622_));
  NO2        u0600(.A(men_men_n446_), .B(i_1_), .Y(men_men_n623_));
  NOi31      u0601(.An(men_men_n623_), .B(men_men_n489_), .C(men_men_n71_), .Y(men_men_n624_));
  AN4        u0602(.A(men_men_n624_), .B(men_men_n443_), .C(men_men_n539_), .D(i_2_), .Y(men_men_n625_));
  NO2        u0603(.A(men_men_n457_), .B(men_men_n180_), .Y(men_men_n626_));
  NO3        u0604(.A(men_men_n626_), .B(men_men_n625_), .C(men_men_n622_), .Y(men_men_n627_));
  NOi21      u0605(.An(i_10_), .B(i_6_), .Y(men_men_n628_));
  NO2        u0606(.A(men_men_n84_), .B(men_men_n25_), .Y(men_men_n629_));
  AOI220     u0607(.A0(men_men_n297_), .A1(men_men_n629_), .B0(men_men_n288_), .B1(men_men_n628_), .Y(men_men_n630_));
  NO2        u0608(.A(men_men_n630_), .B(men_men_n487_), .Y(men_men_n631_));
  NO2        u0609(.A(men_men_n116_), .B(men_men_n23_), .Y(men_men_n632_));
  NA2        u0610(.A(men_men_n332_), .B(men_men_n166_), .Y(men_men_n633_));
  AOI220     u0611(.A0(men_men_n633_), .A1(men_men_n468_), .B0(men_men_n187_), .B1(men_men_n185_), .Y(men_men_n634_));
  NO2        u0612(.A(men_men_n202_), .B(men_men_n35_), .Y(men_men_n635_));
  NOi31      u0613(.An(men_men_n147_), .B(men_men_n635_), .C(men_men_n350_), .Y(men_men_n636_));
  NO3        u0614(.A(men_men_n636_), .B(men_men_n634_), .C(men_men_n631_), .Y(men_men_n637_));
  NO2        u0615(.A(men_men_n563_), .B(men_men_n405_), .Y(men_men_n638_));
  INV        u0616(.A(men_men_n335_), .Y(men_men_n639_));
  NO2        u0617(.A(i_12_), .B(men_men_n84_), .Y(men_men_n640_));
  NA3        u0618(.A(men_men_n640_), .B(men_men_n288_), .C(men_men_n614_), .Y(men_men_n641_));
  NA3        u0619(.A(men_men_n413_), .B(men_men_n297_), .C(men_men_n225_), .Y(men_men_n642_));
  AOI210     u0620(.A0(men_men_n642_), .A1(men_men_n641_), .B0(men_men_n639_), .Y(men_men_n643_));
  NA2        u0621(.A(men_men_n177_), .B(i_0_), .Y(men_men_n644_));
  NO3        u0622(.A(men_men_n644_), .B(men_men_n361_), .C(men_men_n316_), .Y(men_men_n645_));
  OR2        u0623(.A(i_2_), .B(i_5_), .Y(men_men_n646_));
  OR2        u0624(.A(men_men_n646_), .B(men_men_n438_), .Y(men_men_n647_));
  AOI210     u0625(.A0(men_men_n399_), .A1(men_men_n253_), .B0(men_men_n202_), .Y(men_men_n648_));
  AOI210     u0626(.A0(men_men_n648_), .A1(men_men_n647_), .B0(men_men_n537_), .Y(men_men_n649_));
  NO4        u0627(.A(men_men_n649_), .B(men_men_n645_), .C(men_men_n643_), .D(men_men_n638_), .Y(men_men_n650_));
  NA4        u0628(.A(men_men_n650_), .B(men_men_n637_), .C(men_men_n627_), .D(men_men_n617_), .Y(men_men_n651_));
  NO4        u0629(.A(men_men_n651_), .B(men_men_n604_), .C(men_men_n577_), .D(men_men_n550_), .Y(men_men_n652_));
  NA4        u0630(.A(men_men_n652_), .B(men_men_n476_), .C(men_men_n378_), .D(men_men_n328_), .Y(men7));
  OAI220     u0631(.A0(men_men_n544_), .A1(men_men_n119_), .B0(men_men_n93_), .B1(men_men_n52_), .Y(men_men_n654_));
  NO2        u0632(.A(men_men_n109_), .B(men_men_n90_), .Y(men_men_n655_));
  NA2        u0633(.A(men_men_n411_), .B(men_men_n655_), .Y(men_men_n656_));
  NA2        u0634(.A(men_men_n524_), .B(men_men_n82_), .Y(men_men_n657_));
  NA2        u0635(.A(i_11_), .B(men_men_n197_), .Y(men_men_n658_));
  NA2        u0636(.A(men_men_n145_), .B(men_men_n658_), .Y(men_men_n659_));
  OAI210     u0637(.A0(men_men_n659_), .A1(men_men_n657_), .B0(men_men_n656_), .Y(men_men_n660_));
  NA3        u0638(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n661_));
  NO2        u0639(.A(men_men_n245_), .B(i_4_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(i_8_), .Y(men_men_n663_));
  AOI210     u0641(.A0(men_men_n663_), .A1(men_men_n106_), .B0(men_men_n661_), .Y(men_men_n664_));
  NA2        u0642(.A(i_2_), .B(men_men_n84_), .Y(men_men_n665_));
  OAI210     u0643(.A0(men_men_n87_), .A1(men_men_n207_), .B0(men_men_n208_), .Y(men_men_n666_));
  NO2        u0644(.A(i_7_), .B(men_men_n35_), .Y(men_men_n667_));
  NA2        u0645(.A(i_4_), .B(i_8_), .Y(men_men_n668_));
  AOI210     u0646(.A0(men_men_n668_), .A1(men_men_n322_), .B0(men_men_n667_), .Y(men_men_n669_));
  OAI220     u0647(.A0(men_men_n669_), .A1(men_men_n665_), .B0(men_men_n666_), .B1(i_13_), .Y(men_men_n670_));
  NO4        u0648(.A(men_men_n670_), .B(men_men_n664_), .C(men_men_n660_), .D(men_men_n654_), .Y(men_men_n671_));
  AOI210     u0649(.A0(men_men_n130_), .A1(men_men_n60_), .B0(i_10_), .Y(men_men_n672_));
  AOI210     u0650(.A0(men_men_n672_), .A1(men_men_n245_), .B0(men_men_n163_), .Y(men_men_n673_));
  OR2        u0651(.A(i_6_), .B(i_10_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(men_men_n23_), .Y(men_men_n675_));
  OR3        u0653(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n676_));
  NO3        u0654(.A(men_men_n676_), .B(i_8_), .C(men_men_n29_), .Y(men_men_n677_));
  INV        u0655(.A(men_men_n204_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n677_), .B(men_men_n675_), .Y(men_men_n679_));
  OA220      u0657(.A0(men_men_n679_), .A1(men_men_n639_), .B0(men_men_n673_), .B1(men_men_n280_), .Y(men_men_n680_));
  AOI210     u0658(.A0(men_men_n680_), .A1(men_men_n671_), .B0(men_men_n61_), .Y(men_men_n681_));
  NOi21      u0659(.An(i_11_), .B(i_7_), .Y(men_men_n682_));
  AO210      u0660(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n683_));
  NO2        u0661(.A(men_men_n683_), .B(men_men_n682_), .Y(men_men_n684_));
  NA2        u0662(.A(men_men_n684_), .B(men_men_n212_), .Y(men_men_n685_));
  NA3        u0663(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n686_));
  NAi31      u0664(.An(men_men_n686_), .B(men_men_n222_), .C(i_11_), .Y(men_men_n687_));
  AOI210     u0665(.A0(men_men_n687_), .A1(men_men_n685_), .B0(men_men_n61_), .Y(men_men_n688_));
  NA2        u0666(.A(men_men_n86_), .B(men_men_n61_), .Y(men_men_n689_));
  AO210      u0667(.A0(men_men_n689_), .A1(men_men_n405_), .B0(men_men_n38_), .Y(men_men_n690_));
  NO3        u0668(.A(men_men_n269_), .B(men_men_n214_), .C(men_men_n658_), .Y(men_men_n691_));
  OAI210     u0669(.A0(men_men_n691_), .A1(men_men_n234_), .B0(men_men_n61_), .Y(men_men_n692_));
  NA2        u0670(.A(men_men_n439_), .B(men_men_n29_), .Y(men_men_n693_));
  OR2        u0671(.A(men_men_n214_), .B(men_men_n109_), .Y(men_men_n694_));
  NA2        u0672(.A(men_men_n694_), .B(men_men_n693_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n61_), .B(i_9_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n696_), .B(i_4_), .Y(men_men_n697_));
  NA2        u0675(.A(men_men_n697_), .B(men_men_n695_), .Y(men_men_n698_));
  NO2        u0676(.A(i_1_), .B(i_12_), .Y(men_men_n699_));
  NA3        u0677(.A(men_men_n699_), .B(men_men_n111_), .C(men_men_n24_), .Y(men_men_n700_));
  NA4        u0678(.A(men_men_n700_), .B(men_men_n698_), .C(men_men_n692_), .D(men_men_n690_), .Y(men_men_n701_));
  OAI210     u0679(.A0(men_men_n701_), .A1(men_men_n688_), .B0(i_6_), .Y(men_men_n702_));
  OAI210     u0680(.A0(men_men_n686_), .A1(men_men_n109_), .B0(men_men_n499_), .Y(men_men_n703_));
  NA2        u0681(.A(men_men_n703_), .B(men_men_n640_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n245_), .B(men_men_n84_), .Y(men_men_n705_));
  NA3        u0683(.A(men_men_n704_), .B(men_men_n567_), .C(men_men_n490_), .Y(men_men_n706_));
  NO4        u0684(.A(men_men_n222_), .B(men_men_n130_), .C(i_13_), .D(men_men_n84_), .Y(men_men_n707_));
  NA2        u0685(.A(men_men_n707_), .B(men_men_n696_), .Y(men_men_n708_));
  NA2        u0686(.A(men_men_n245_), .B(i_6_), .Y(men_men_n709_));
  NO3        u0687(.A(men_men_n674_), .B(men_men_n241_), .C(men_men_n23_), .Y(men_men_n710_));
  AOI210     u0688(.A0(i_1_), .A1(men_men_n270_), .B0(men_men_n710_), .Y(men_men_n711_));
  OAI210     u0689(.A0(men_men_n711_), .A1(men_men_n42_), .B0(men_men_n708_), .Y(men_men_n712_));
  NA3        u0690(.A(men_men_n586_), .B(i_11_), .C(men_men_n34_), .Y(men_men_n713_));
  NA3        u0691(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n714_));
  NO2        u0692(.A(men_men_n44_), .B(i_1_), .Y(men_men_n715_));
  NA3        u0693(.A(men_men_n715_), .B(men_men_n279_), .C(men_men_n42_), .Y(men_men_n716_));
  NO2        u0694(.A(men_men_n716_), .B(men_men_n714_), .Y(men_men_n717_));
  NA3        u0695(.A(men_men_n696_), .B(men_men_n335_), .C(i_6_), .Y(men_men_n718_));
  NO2        u0696(.A(men_men_n718_), .B(men_men_n23_), .Y(men_men_n719_));
  NAi21      u0697(.An(men_men_n713_), .B(men_men_n92_), .Y(men_men_n720_));
  NA2        u0698(.A(men_men_n715_), .B(men_men_n279_), .Y(men_men_n721_));
  NO2        u0699(.A(i_11_), .B(men_men_n35_), .Y(men_men_n722_));
  NA2        u0700(.A(men_men_n722_), .B(men_men_n24_), .Y(men_men_n723_));
  OAI210     u0701(.A0(men_men_n723_), .A1(men_men_n721_), .B0(men_men_n720_), .Y(men_men_n724_));
  OR3        u0702(.A(men_men_n724_), .B(men_men_n719_), .C(men_men_n717_), .Y(men_men_n725_));
  NO3        u0703(.A(men_men_n725_), .B(men_men_n712_), .C(men_men_n706_), .Y(men_men_n726_));
  NO2        u0704(.A(men_men_n245_), .B(men_men_n102_), .Y(men_men_n727_));
  NO2        u0705(.A(men_men_n727_), .B(men_men_n682_), .Y(men_men_n728_));
  NA2        u0706(.A(men_men_n728_), .B(i_1_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n729_), .B(men_men_n676_), .Y(men_men_n730_));
  NO2        u0708(.A(men_men_n445_), .B(men_men_n84_), .Y(men_men_n731_));
  NA2        u0709(.A(men_men_n730_), .B(men_men_n44_), .Y(men_men_n732_));
  NA2        u0710(.A(i_3_), .B(men_men_n197_), .Y(men_men_n733_));
  AOI210     u0711(.A0(men_men_n268_), .A1(men_men_n733_), .B0(men_men_n116_), .Y(men_men_n734_));
  AN2        u0712(.A(men_men_n734_), .B(men_men_n592_), .Y(men_men_n735_));
  NO2        u0713(.A(men_men_n241_), .B(men_men_n42_), .Y(men_men_n736_));
  NO3        u0714(.A(men_men_n736_), .B(men_men_n325_), .C(men_men_n246_), .Y(men_men_n737_));
  NO2        u0715(.A(men_men_n119_), .B(men_men_n35_), .Y(men_men_n738_));
  NO2        u0716(.A(men_men_n738_), .B(i_6_), .Y(men_men_n739_));
  NO2        u0717(.A(men_men_n84_), .B(i_9_), .Y(men_men_n740_));
  NO2        u0718(.A(men_men_n740_), .B(men_men_n61_), .Y(men_men_n741_));
  NO2        u0719(.A(men_men_n741_), .B(men_men_n699_), .Y(men_men_n742_));
  NO4        u0720(.A(men_men_n742_), .B(men_men_n739_), .C(men_men_n737_), .D(i_4_), .Y(men_men_n743_));
  NA2        u0721(.A(i_1_), .B(i_3_), .Y(men_men_n744_));
  NO2        u0722(.A(men_men_n491_), .B(men_men_n93_), .Y(men_men_n745_));
  AOI210     u0723(.A0(men_men_n736_), .A1(men_men_n628_), .B0(men_men_n745_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n746_), .B(men_men_n744_), .Y(men_men_n747_));
  NO3        u0725(.A(men_men_n747_), .B(men_men_n743_), .C(men_men_n735_), .Y(men_men_n748_));
  NA4        u0726(.A(men_men_n748_), .B(men_men_n732_), .C(men_men_n726_), .D(men_men_n702_), .Y(men_men_n749_));
  NO3        u0727(.A(men_men_n517_), .B(i_3_), .C(i_7_), .Y(men_men_n750_));
  NOi21      u0728(.An(men_men_n750_), .B(i_10_), .Y(men_men_n751_));
  OA210      u0729(.A0(men_men_n751_), .A1(men_men_n254_), .B0(men_men_n84_), .Y(men_men_n752_));
  NA2        u0730(.A(men_men_n397_), .B(men_men_n396_), .Y(men_men_n753_));
  NA3        u0731(.A(men_men_n524_), .B(men_men_n566_), .C(men_men_n44_), .Y(men_men_n754_));
  NO3        u0732(.A(men_men_n518_), .B(men_men_n668_), .C(men_men_n84_), .Y(men_men_n755_));
  NA2        u0733(.A(men_men_n755_), .B(men_men_n25_), .Y(men_men_n756_));
  NA3        u0734(.A(men_men_n163_), .B(men_men_n82_), .C(men_men_n84_), .Y(men_men_n757_));
  NA4        u0735(.A(men_men_n757_), .B(men_men_n756_), .C(men_men_n754_), .D(men_men_n753_), .Y(men_men_n758_));
  OAI210     u0736(.A0(men_men_n758_), .A1(men_men_n752_), .B0(i_1_), .Y(men_men_n759_));
  AOI210     u0737(.A0(men_men_n279_), .A1(men_men_n98_), .B0(i_1_), .Y(men_men_n760_));
  NO2        u0738(.A(men_men_n395_), .B(i_2_), .Y(men_men_n761_));
  NA2        u0739(.A(men_men_n761_), .B(men_men_n760_), .Y(men_men_n762_));
  OAI210     u0740(.A0(men_men_n718_), .A1(men_men_n481_), .B0(men_men_n762_), .Y(men_men_n763_));
  INV        u0741(.A(men_men_n763_), .Y(men_men_n764_));
  AOI210     u0742(.A0(men_men_n764_), .A1(men_men_n759_), .B0(i_13_), .Y(men_men_n765_));
  OR2        u0743(.A(i_11_), .B(i_7_), .Y(men_men_n766_));
  NA3        u0744(.A(men_men_n766_), .B(men_men_n107_), .C(men_men_n140_), .Y(men_men_n767_));
  AOI220     u0745(.A0(men_men_n509_), .A1(men_men_n163_), .B0(men_men_n484_), .B1(men_men_n140_), .Y(men_men_n768_));
  OAI210     u0746(.A0(men_men_n768_), .A1(men_men_n42_), .B0(men_men_n767_), .Y(men_men_n769_));
  NO3        u0747(.A(men_men_n518_), .B(men_men_n586_), .C(men_men_n24_), .Y(men_men_n770_));
  AOI220     u0748(.A0(men_men_n770_), .A1(men_men_n731_), .B0(men_men_n254_), .B1(men_men_n133_), .Y(men_men_n771_));
  NO2        u0749(.A(men_men_n771_), .B(men_men_n38_), .Y(men_men_n772_));
  AOI210     u0750(.A0(men_men_n769_), .A1(men_men_n352_), .B0(men_men_n772_), .Y(men_men_n773_));
  NA2        u0751(.A(men_men_n116_), .B(men_men_n109_), .Y(men_men_n774_));
  AOI220     u0752(.A0(men_men_n774_), .A1(men_men_n70_), .B0(men_men_n413_), .B1(men_men_n715_), .Y(men_men_n775_));
  NO2        u0753(.A(men_men_n775_), .B(men_men_n251_), .Y(men_men_n776_));
  AOI210     u0754(.A0(men_men_n481_), .A1(men_men_n34_), .B0(i_13_), .Y(men_men_n777_));
  NOi31      u0755(.An(men_men_n777_), .B(men_men_n657_), .C(men_men_n42_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n714_), .B(men_men_n116_), .Y(men_men_n779_));
  INV        u0757(.A(men_men_n779_), .Y(men_men_n780_));
  NO2        u0758(.A(men_men_n780_), .B(men_men_n69_), .Y(men_men_n781_));
  NO3        u0759(.A(men_men_n69_), .B(men_men_n30_), .C(men_men_n102_), .Y(men_men_n782_));
  NA2        u0760(.A(men_men_n26_), .B(men_men_n197_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(i_7_), .Y(men_men_n784_));
  NO3        u0762(.A(men_men_n518_), .B(men_men_n245_), .C(men_men_n84_), .Y(men_men_n785_));
  AOI210     u0763(.A0(men_men_n785_), .A1(men_men_n784_), .B0(men_men_n782_), .Y(men_men_n786_));
  AOI220     u0764(.A0(men_men_n413_), .A1(men_men_n715_), .B0(men_men_n92_), .B1(men_men_n103_), .Y(men_men_n787_));
  OAI220     u0765(.A0(men_men_n787_), .A1(men_men_n663_), .B0(men_men_n786_), .B1(men_men_n678_), .Y(men_men_n788_));
  NO4        u0766(.A(men_men_n788_), .B(men_men_n781_), .C(men_men_n778_), .D(men_men_n776_), .Y(men_men_n789_));
  OR2        u0767(.A(i_11_), .B(i_6_), .Y(men_men_n790_));
  NA3        u0768(.A(men_men_n662_), .B(men_men_n783_), .C(i_7_), .Y(men_men_n791_));
  AOI210     u0769(.A0(men_men_n791_), .A1(men_men_n780_), .B0(men_men_n790_), .Y(men_men_n792_));
  NA2        u0770(.A(men_men_n103_), .B(men_men_n783_), .Y(men_men_n793_));
  NAi21      u0771(.An(i_11_), .B(i_12_), .Y(men_men_n794_));
  NOi41      u0772(.An(men_men_n112_), .B(men_men_n794_), .C(i_13_), .D(men_men_n84_), .Y(men_men_n795_));
  NO3        u0773(.A(men_men_n518_), .B(men_men_n640_), .C(men_men_n668_), .Y(men_men_n796_));
  AOI220     u0774(.A0(men_men_n796_), .A1(men_men_n329_), .B0(men_men_n795_), .B1(men_men_n793_), .Y(men_men_n797_));
  INV        u0775(.A(men_men_n797_), .Y(men_men_n798_));
  OAI210     u0776(.A0(men_men_n798_), .A1(men_men_n792_), .B0(men_men_n61_), .Y(men_men_n799_));
  NO2        u0777(.A(i_2_), .B(i_12_), .Y(men_men_n800_));
  OAI210     u0778(.A0(men_men_n672_), .A1(men_men_n394_), .B0(men_men_n800_), .Y(men_men_n801_));
  NA2        u0779(.A(i_8_), .B(men_men_n25_), .Y(men_men_n802_));
  NO3        u0780(.A(men_men_n802_), .B(men_men_n411_), .C(men_men_n662_), .Y(men_men_n803_));
  OAI210     u0781(.A0(men_men_n803_), .A1(men_men_n396_), .B0(men_men_n394_), .Y(men_men_n804_));
  NO2        u0782(.A(men_men_n130_), .B(i_2_), .Y(men_men_n805_));
  NA2        u0783(.A(men_men_n805_), .B(men_men_n699_), .Y(men_men_n806_));
  NA3        u0784(.A(men_men_n806_), .B(men_men_n804_), .C(men_men_n801_), .Y(men_men_n807_));
  NA3        u0785(.A(men_men_n807_), .B(men_men_n43_), .C(men_men_n233_), .Y(men_men_n808_));
  NA4        u0786(.A(men_men_n808_), .B(men_men_n799_), .C(men_men_n789_), .D(men_men_n773_), .Y(men_men_n809_));
  OR4        u0787(.A(men_men_n809_), .B(men_men_n765_), .C(men_men_n749_), .D(men_men_n681_), .Y(men5));
  AOI210     u0788(.A0(men_men_n728_), .A1(men_men_n282_), .B0(men_men_n448_), .Y(men_men_n811_));
  NA3        u0789(.A(men_men_n24_), .B(men_men_n800_), .C(men_men_n109_), .Y(men_men_n812_));
  NO2        u0790(.A(men_men_n663_), .B(i_11_), .Y(men_men_n813_));
  OAI210     u0791(.A0(men_men_n667_), .A1(men_men_n87_), .B0(men_men_n813_), .Y(men_men_n814_));
  NA4        u0792(.A(men_men_n814_), .B(men_men_n812_), .C(men_men_n811_), .D(men_men_n567_), .Y(men_men_n815_));
  NO3        u0793(.A(i_11_), .B(men_men_n245_), .C(i_13_), .Y(men_men_n816_));
  NO2        u0794(.A(men_men_n126_), .B(men_men_n23_), .Y(men_men_n817_));
  NA2        u0795(.A(i_12_), .B(i_8_), .Y(men_men_n818_));
  OAI210     u0796(.A0(men_men_n44_), .A1(i_3_), .B0(men_men_n818_), .Y(men_men_n819_));
  AOI220     u0797(.A0(men_men_n335_), .A1(men_men_n632_), .B0(men_men_n819_), .B1(men_men_n817_), .Y(men_men_n820_));
  INV        u0798(.A(men_men_n820_), .Y(men_men_n821_));
  NO2        u0799(.A(men_men_n821_), .B(men_men_n815_), .Y(men_men_n822_));
  INV        u0800(.A(men_men_n174_), .Y(men_men_n823_));
  INV        u0801(.A(men_men_n254_), .Y(men_men_n824_));
  OAI210     u0802(.A0(men_men_n761_), .A1(men_men_n482_), .B0(men_men_n112_), .Y(men_men_n825_));
  AOI210     u0803(.A0(men_men_n825_), .A1(men_men_n824_), .B0(men_men_n823_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n491_), .B(men_men_n26_), .Y(men_men_n827_));
  NO2        u0805(.A(men_men_n827_), .B(men_men_n450_), .Y(men_men_n828_));
  AOI210     u0806(.A0(men_men_n31_), .A1(men_men_n34_), .B0(men_men_n446_), .Y(men_men_n829_));
  AOI210     u0807(.A0(men_men_n829_), .A1(i_2_), .B0(men_men_n826_), .Y(men_men_n830_));
  NO2        u0808(.A(men_men_n194_), .B(men_men_n127_), .Y(men_men_n831_));
  OAI210     u0809(.A0(men_men_n831_), .A1(men_men_n817_), .B0(i_2_), .Y(men_men_n832_));
  NO3        u0810(.A(men_men_n683_), .B(men_men_n36_), .C(men_men_n26_), .Y(men_men_n833_));
  AOI210     u0811(.A0(men_men_n173_), .A1(men_men_n87_), .B0(men_men_n833_), .Y(men_men_n834_));
  AOI210     u0812(.A0(men_men_n834_), .A1(men_men_n832_), .B0(men_men_n197_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n204_), .B(men_men_n207_), .Y(men_men_n836_));
  NA2        u0814(.A(men_men_n153_), .B(men_men_n658_), .Y(men_men_n837_));
  AOI210     u0815(.A0(men_men_n837_), .A1(men_men_n836_), .B0(men_men_n399_), .Y(men_men_n838_));
  AOI210     u0816(.A0(men_men_n214_), .A1(men_men_n149_), .B0(men_men_n566_), .Y(men_men_n839_));
  OAI210     u0817(.A0(men_men_n839_), .A1(men_men_n234_), .B0(men_men_n450_), .Y(men_men_n840_));
  NA4        u0818(.A(men_men_n102_), .B(men_men_n322_), .C(men_men_n126_), .D(men_men_n40_), .Y(men_men_n841_));
  OAI210     u0819(.A0(men_men_n841_), .A1(i_11_), .B0(men_men_n840_), .Y(men_men_n842_));
  NO3        u0820(.A(men_men_n842_), .B(men_men_n838_), .C(men_men_n835_), .Y(men_men_n843_));
  NA2        u0821(.A(men_men_n632_), .B(men_men_n28_), .Y(men_men_n844_));
  NA2        u0822(.A(men_men_n816_), .B(men_men_n289_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n845_), .B(men_men_n844_), .Y(men_men_n846_));
  NO2        u0824(.A(men_men_n60_), .B(i_12_), .Y(men_men_n847_));
  NO2        u0825(.A(men_men_n847_), .B(men_men_n128_), .Y(men_men_n848_));
  NO2        u0826(.A(men_men_n848_), .B(men_men_n658_), .Y(men_men_n849_));
  AOI220     u0827(.A0(men_men_n849_), .A1(men_men_n34_), .B0(men_men_n846_), .B1(men_men_n44_), .Y(men_men_n850_));
  NA4        u0828(.A(men_men_n850_), .B(men_men_n843_), .C(men_men_n830_), .D(men_men_n822_), .Y(men6));
  NO3        u0829(.A(men_men_n265_), .B(men_men_n324_), .C(i_1_), .Y(men_men_n852_));
  NO2        u0830(.A(men_men_n189_), .B(men_men_n141_), .Y(men_men_n853_));
  OAI210     u0831(.A0(men_men_n853_), .A1(men_men_n852_), .B0(men_men_n805_), .Y(men_men_n854_));
  NA4        u0832(.A(men_men_n417_), .B(men_men_n523_), .C(men_men_n69_), .D(men_men_n102_), .Y(men_men_n855_));
  INV        u0833(.A(men_men_n855_), .Y(men_men_n856_));
  NO2        u0834(.A(men_men_n228_), .B(men_men_n528_), .Y(men_men_n857_));
  NO2        u0835(.A(i_11_), .B(i_9_), .Y(men_men_n858_));
  AO210      u0836(.A0(men_men_n855_), .A1(men_men_n854_), .B0(i_12_), .Y(men_men_n859_));
  NA2        u0837(.A(men_men_n400_), .B(men_men_n355_), .Y(men_men_n860_));
  NA2        u0838(.A(men_men_n640_), .B(men_men_n61_), .Y(men_men_n861_));
  NA2        u0839(.A(men_men_n751_), .B(men_men_n69_), .Y(men_men_n862_));
  NA4        u0840(.A(men_men_n689_), .B(men_men_n862_), .C(men_men_n861_), .D(men_men_n860_), .Y(men_men_n863_));
  INV        u0841(.A(men_men_n201_), .Y(men_men_n864_));
  AOI220     u0842(.A0(men_men_n864_), .A1(men_men_n858_), .B0(men_men_n863_), .B1(men_men_n71_), .Y(men_men_n865_));
  INV        u0843(.A(men_men_n346_), .Y(men_men_n866_));
  NA2        u0844(.A(men_men_n73_), .B(men_men_n133_), .Y(men_men_n867_));
  OAI210     u0845(.A0(men_men_n790_), .A1(i_5_), .B0(men_men_n126_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n868_), .B(men_men_n44_), .Y(men_men_n869_));
  AOI210     u0847(.A0(men_men_n869_), .A1(men_men_n867_), .B0(men_men_n866_), .Y(men_men_n870_));
  NO3        u0848(.A(men_men_n261_), .B(men_men_n134_), .C(i_9_), .Y(men_men_n871_));
  NA2        u0849(.A(men_men_n871_), .B(men_men_n847_), .Y(men_men_n872_));
  AOI210     u0850(.A0(men_men_n872_), .A1(men_men_n564_), .B0(men_men_n189_), .Y(men_men_n873_));
  NO2        u0851(.A(men_men_n30_), .B(i_11_), .Y(men_men_n874_));
  NA3        u0852(.A(men_men_n874_), .B(men_men_n513_), .C(men_men_n417_), .Y(men_men_n875_));
  NAi32      u0853(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n876_));
  AOI210     u0854(.A0(men_men_n790_), .A1(men_men_n85_), .B0(men_men_n876_), .Y(men_men_n877_));
  OAI210     u0855(.A0(men_men_n750_), .A1(men_men_n620_), .B0(men_men_n619_), .Y(men_men_n878_));
  NAi31      u0856(.An(men_men_n877_), .B(men_men_n878_), .C(men_men_n875_), .Y(men_men_n879_));
  OR3        u0857(.A(men_men_n879_), .B(men_men_n873_), .C(men_men_n870_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n766_), .B(i_2_), .Y(men_men_n881_));
  NA2        u0859(.A(men_men_n46_), .B(men_men_n35_), .Y(men_men_n882_));
  OAI210     u0860(.A0(men_men_n882_), .A1(men_men_n438_), .B0(men_men_n384_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n883_), .B(men_men_n881_), .Y(men_men_n884_));
  AO220      u0862(.A0(men_men_n383_), .A1(men_men_n373_), .B0(men_men_n425_), .B1(men_men_n658_), .Y(men_men_n885_));
  NA3        u0863(.A(men_men_n885_), .B(men_men_n266_), .C(i_7_), .Y(men_men_n886_));
  OR2        u0864(.A(men_men_n684_), .B(men_men_n482_), .Y(men_men_n887_));
  NA3        u0865(.A(men_men_n887_), .B(men_men_n148_), .C(men_men_n67_), .Y(men_men_n888_));
  OR2        u0866(.A(men_men_n535_), .B(men_men_n34_), .Y(men_men_n889_));
  NA4        u0867(.A(men_men_n889_), .B(men_men_n888_), .C(men_men_n886_), .D(men_men_n884_), .Y(men_men_n890_));
  OAI210     u0868(.A0(men_men_n705_), .A1(i_11_), .B0(men_men_n85_), .Y(men_men_n891_));
  AOI220     u0869(.A0(men_men_n891_), .A1(men_men_n619_), .B0(men_men_n857_), .B1(men_men_n784_), .Y(men_men_n892_));
  NA3        u0870(.A(men_men_n399_), .B(men_men_n247_), .C(men_men_n148_), .Y(men_men_n893_));
  OAI210     u0871(.A0(men_men_n425_), .A1(men_men_n208_), .B0(men_men_n68_), .Y(men_men_n894_));
  NA4        u0872(.A(men_men_n894_), .B(men_men_n893_), .C(men_men_n892_), .D(men_men_n666_), .Y(men_men_n895_));
  AO210      u0873(.A0(men_men_n566_), .A1(men_men_n44_), .B0(men_men_n86_), .Y(men_men_n896_));
  NA3        u0874(.A(men_men_n896_), .B(men_men_n524_), .C(men_men_n225_), .Y(men_men_n897_));
  AOI210     u0875(.A0(men_men_n482_), .A1(men_men_n480_), .B0(men_men_n618_), .Y(men_men_n898_));
  NO2        u0876(.A(men_men_n674_), .B(men_men_n103_), .Y(men_men_n899_));
  OAI210     u0877(.A0(men_men_n899_), .A1(men_men_n113_), .B0(men_men_n437_), .Y(men_men_n900_));
  NA2        u0878(.A(men_men_n253_), .B(men_men_n44_), .Y(men_men_n901_));
  NA2        u0879(.A(men_men_n901_), .B(men_men_n647_), .Y(men_men_n902_));
  NA3        u0880(.A(men_men_n902_), .B(men_men_n346_), .C(i_7_), .Y(men_men_n903_));
  NA4        u0881(.A(men_men_n903_), .B(men_men_n900_), .C(men_men_n898_), .D(men_men_n897_), .Y(men_men_n904_));
  NO4        u0882(.A(men_men_n904_), .B(men_men_n895_), .C(men_men_n890_), .D(men_men_n880_), .Y(men_men_n905_));
  NA4        u0883(.A(men_men_n905_), .B(men_men_n865_), .C(men_men_n859_), .D(men_men_n407_), .Y(men3));
  NA2        u0884(.A(i_12_), .B(i_10_), .Y(men_men_n907_));
  NA2        u0885(.A(i_6_), .B(i_7_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n908_), .B(i_0_), .Y(men_men_n909_));
  NO2        u0887(.A(i_11_), .B(men_men_n245_), .Y(men_men_n910_));
  OAI210     u0888(.A0(men_men_n909_), .A1(men_men_n305_), .B0(men_men_n910_), .Y(men_men_n911_));
  NO2        u0889(.A(men_men_n911_), .B(men_men_n197_), .Y(men_men_n912_));
  NO3        u0890(.A(men_men_n487_), .B(men_men_n90_), .C(men_men_n42_), .Y(men_men_n913_));
  OA210      u0891(.A0(men_men_n913_), .A1(men_men_n912_), .B0(men_men_n177_), .Y(men_men_n914_));
  NA3        u0892(.A(men_men_n893_), .B(men_men_n666_), .C(men_men_n398_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n915_), .B(men_men_n37_), .Y(men_men_n916_));
  NOi21      u0894(.An(men_men_n97_), .B(men_men_n828_), .Y(men_men_n917_));
  NO3        u0895(.A(men_men_n694_), .B(men_men_n491_), .C(men_men_n133_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n439_), .B(men_men_n43_), .Y(men_men_n919_));
  AN2        u0897(.A(men_men_n489_), .B(men_men_n53_), .Y(men_men_n920_));
  NO3        u0898(.A(men_men_n920_), .B(men_men_n918_), .C(men_men_n917_), .Y(men_men_n921_));
  AOI210     u0899(.A0(men_men_n921_), .A1(men_men_n916_), .B0(men_men_n46_), .Y(men_men_n922_));
  NO4        u0900(.A(men_men_n403_), .B(men_men_n410_), .C(men_men_n36_), .D(i_0_), .Y(men_men_n923_));
  NA2        u0901(.A(men_men_n189_), .B(men_men_n628_), .Y(men_men_n924_));
  NOi21      u0902(.An(men_men_n924_), .B(men_men_n923_), .Y(men_men_n925_));
  NA2        u0903(.A(men_men_n777_), .B(men_men_n740_), .Y(men_men_n926_));
  NA2        u0904(.A(men_men_n353_), .B(men_men_n470_), .Y(men_men_n927_));
  OAI220     u0905(.A0(men_men_n927_), .A1(men_men_n926_), .B0(men_men_n925_), .B1(men_men_n61_), .Y(men_men_n928_));
  NOi21      u0906(.An(i_5_), .B(i_9_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n929_), .B(men_men_n478_), .Y(men_men_n930_));
  AOI210     u0908(.A0(men_men_n279_), .A1(men_men_n515_), .B0(men_men_n755_), .Y(men_men_n931_));
  NO3        u0909(.A(men_men_n442_), .B(men_men_n279_), .C(men_men_n71_), .Y(men_men_n932_));
  NO2        u0910(.A(men_men_n178_), .B(men_men_n149_), .Y(men_men_n933_));
  AOI210     u0911(.A0(men_men_n933_), .A1(men_men_n253_), .B0(men_men_n932_), .Y(men_men_n934_));
  OAI220     u0912(.A0(men_men_n934_), .A1(men_men_n184_), .B0(men_men_n931_), .B1(men_men_n930_), .Y(men_men_n935_));
  NO4        u0913(.A(men_men_n935_), .B(men_men_n928_), .C(men_men_n922_), .D(men_men_n914_), .Y(men_men_n936_));
  NOi21      u0914(.An(i_0_), .B(i_10_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n189_), .B(men_men_n24_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n738_), .B(men_men_n655_), .Y(men_men_n939_));
  NO2        u0917(.A(men_men_n939_), .B(men_men_n938_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n329_), .B(men_men_n131_), .Y(men_men_n941_));
  NAi21      u0919(.An(men_men_n164_), .B(men_men_n470_), .Y(men_men_n942_));
  OAI220     u0920(.A0(men_men_n942_), .A1(men_men_n901_), .B0(men_men_n941_), .B1(men_men_n428_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n943_), .B(men_men_n940_), .Y(men_men_n944_));
  NA2        u0922(.A(men_men_n629_), .B(i_0_), .Y(men_men_n945_));
  NO3        u0923(.A(men_men_n945_), .B(men_men_n412_), .C(men_men_n87_), .Y(men_men_n946_));
  NO4        u0924(.A(men_men_n646_), .B(men_men_n222_), .C(men_men_n446_), .D(men_men_n438_), .Y(men_men_n947_));
  AOI210     u0925(.A0(men_men_n947_), .A1(i_11_), .B0(men_men_n946_), .Y(men_men_n948_));
  INV        u0926(.A(men_men_n513_), .Y(men_men_n949_));
  AN2        u0927(.A(men_men_n97_), .B(men_men_n252_), .Y(men_men_n950_));
  NA2        u0928(.A(men_men_n816_), .B(men_men_n347_), .Y(men_men_n951_));
  AOI210     u0929(.A0(men_men_n524_), .A1(men_men_n87_), .B0(men_men_n56_), .Y(men_men_n952_));
  OAI220     u0930(.A0(men_men_n952_), .A1(men_men_n951_), .B0(men_men_n723_), .B1(men_men_n588_), .Y(men_men_n953_));
  NO2        u0931(.A(men_men_n263_), .B(men_men_n155_), .Y(men_men_n954_));
  NA2        u0932(.A(i_0_), .B(i_10_), .Y(men_men_n955_));
  INV        u0933(.A(men_men_n591_), .Y(men_men_n956_));
  NO4        u0934(.A(men_men_n116_), .B(men_men_n56_), .C(men_men_n733_), .D(i_5_), .Y(men_men_n957_));
  AO220      u0935(.A0(men_men_n957_), .A1(men_men_n956_), .B0(men_men_n954_), .B1(i_6_), .Y(men_men_n958_));
  AOI220     u0936(.A0(men_men_n353_), .A1(men_men_n99_), .B0(men_men_n189_), .B1(men_men_n82_), .Y(men_men_n959_));
  NA2        u0937(.A(men_men_n623_), .B(i_4_), .Y(men_men_n960_));
  NA2        u0938(.A(men_men_n192_), .B(men_men_n207_), .Y(men_men_n961_));
  OAI220     u0939(.A0(men_men_n961_), .A1(men_men_n951_), .B0(men_men_n960_), .B1(men_men_n959_), .Y(men_men_n962_));
  NO4        u0940(.A(men_men_n962_), .B(men_men_n958_), .C(men_men_n953_), .D(men_men_n950_), .Y(men_men_n963_));
  NA3        u0941(.A(men_men_n963_), .B(men_men_n948_), .C(men_men_n944_), .Y(men_men_n964_));
  NO2        u0942(.A(men_men_n104_), .B(men_men_n35_), .Y(men_men_n965_));
  NA2        u0943(.A(i_11_), .B(i_9_), .Y(men_men_n966_));
  NO3        u0944(.A(i_12_), .B(men_men_n966_), .C(men_men_n665_), .Y(men_men_n967_));
  AO220      u0945(.A0(men_men_n967_), .A1(men_men_n965_), .B0(men_men_n281_), .B1(men_men_n86_), .Y(men_men_n968_));
  NO2        u0946(.A(men_men_n46_), .B(i_7_), .Y(men_men_n969_));
  NA2        u0947(.A(men_men_n422_), .B(men_men_n182_), .Y(men_men_n970_));
  NAi41      u0948(.An(men_men_n276_), .B(men_men_n970_), .C(men_men_n496_), .D(men_men_n162_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n966_), .B(men_men_n71_), .Y(men_men_n972_));
  NO2        u0950(.A(men_men_n178_), .B(i_0_), .Y(men_men_n973_));
  INV        u0951(.A(men_men_n973_), .Y(men_men_n974_));
  NA2        u0952(.A(men_men_n513_), .B(men_men_n239_), .Y(men_men_n975_));
  AOI210     u0953(.A0(men_men_n397_), .A1(men_men_n39_), .B0(men_men_n436_), .Y(men_men_n976_));
  OAI220     u0954(.A0(men_men_n976_), .A1(men_men_n930_), .B0(men_men_n975_), .B1(men_men_n974_), .Y(men_men_n977_));
  NO3        u0955(.A(men_men_n977_), .B(men_men_n971_), .C(men_men_n968_), .Y(men_men_n978_));
  NA2        u0956(.A(men_men_n722_), .B(men_men_n123_), .Y(men_men_n979_));
  NO2        u0957(.A(i_6_), .B(men_men_n979_), .Y(men_men_n980_));
  AOI210     u0958(.A0(men_men_n481_), .A1(men_men_n34_), .B0(i_3_), .Y(men_men_n981_));
  NA2        u0959(.A(men_men_n174_), .B(men_men_n104_), .Y(men_men_n982_));
  NOi32      u0960(.An(men_men_n981_), .Bn(men_men_n192_), .C(men_men_n982_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n667_), .A1(men_men_n347_), .B0(men_men_n252_), .Y(men_men_n984_));
  NO2        u0962(.A(men_men_n984_), .B(men_men_n919_), .Y(men_men_n985_));
  NO3        u0963(.A(men_men_n985_), .B(men_men_n983_), .C(men_men_n980_), .Y(men_men_n986_));
  NOi21      u0964(.An(i_7_), .B(i_5_), .Y(men_men_n987_));
  NOi31      u0965(.An(men_men_n987_), .B(men_men_n937_), .C(men_men_n794_), .Y(men_men_n988_));
  NA3        u0966(.A(men_men_n988_), .B(men_men_n411_), .C(i_6_), .Y(men_men_n989_));
  OA210      u0967(.A0(men_men_n982_), .A1(men_men_n564_), .B0(men_men_n989_), .Y(men_men_n990_));
  NO3        u0968(.A(men_men_n431_), .B(men_men_n386_), .C(men_men_n382_), .Y(men_men_n991_));
  NO2        u0969(.A(men_men_n273_), .B(men_men_n336_), .Y(men_men_n992_));
  NO2        u0970(.A(men_men_n794_), .B(men_men_n268_), .Y(men_men_n993_));
  AOI210     u0971(.A0(men_men_n993_), .A1(men_men_n992_), .B0(men_men_n991_), .Y(men_men_n994_));
  NA4        u0972(.A(men_men_n994_), .B(men_men_n990_), .C(men_men_n986_), .D(men_men_n978_), .Y(men_men_n995_));
  NO2        u0973(.A(men_men_n938_), .B(men_men_n248_), .Y(men_men_n996_));
  AN2        u0974(.A(men_men_n352_), .B(men_men_n347_), .Y(men_men_n997_));
  AO220      u0975(.A0(men_men_n997_), .A1(men_men_n933_), .B0(men_men_n368_), .B1(men_men_n27_), .Y(men_men_n998_));
  OAI210     u0976(.A0(men_men_n998_), .A1(men_men_n996_), .B0(i_10_), .Y(men_men_n999_));
  NO2        u0977(.A(men_men_n907_), .B(men_men_n335_), .Y(men_men_n1000_));
  OA210      u0978(.A0(men_men_n513_), .A1(men_men_n231_), .B0(men_men_n512_), .Y(men_men_n1001_));
  OAI210     u0979(.A0(men_men_n1001_), .A1(men_men_n1000_), .B0(men_men_n972_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n512_), .B(men_men_n439_), .C(men_men_n43_), .Y(men_men_n1003_));
  OAI210     u0981(.A0(men_men_n942_), .A1(men_men_n949_), .B0(men_men_n1003_), .Y(men_men_n1004_));
  NO2        u0982(.A(men_men_n266_), .B(men_men_n44_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n972_), .B(men_men_n322_), .Y(men_men_n1006_));
  OAI210     u0984(.A0(men_men_n1005_), .A1(men_men_n191_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  AOI220     u0985(.A0(men_men_n1007_), .A1(men_men_n513_), .B0(men_men_n1004_), .B1(men_men_n71_), .Y(men_men_n1008_));
  NA3        u0986(.A(men_men_n882_), .B(men_men_n409_), .C(men_men_n705_), .Y(men_men_n1009_));
  NA2        u0987(.A(men_men_n93_), .B(men_men_n42_), .Y(men_men_n1010_));
  NO2        u0988(.A(men_men_n73_), .B(men_men_n818_), .Y(men_men_n1011_));
  AOI220     u0989(.A0(men_men_n1011_), .A1(men_men_n1010_), .B0(men_men_n177_), .B1(men_men_n655_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n1012_), .A1(men_men_n1009_), .B0(men_men_n45_), .Y(men_men_n1013_));
  NO3        u0991(.A(men_men_n646_), .B(men_men_n381_), .C(men_men_n24_), .Y(men_men_n1014_));
  AOI210     u0992(.A0(men_men_n770_), .A1(men_men_n600_), .B0(men_men_n1014_), .Y(men_men_n1015_));
  NAi21      u0993(.An(i_9_), .B(i_5_), .Y(men_men_n1016_));
  NO2        u0994(.A(men_men_n1016_), .B(men_men_n431_), .Y(men_men_n1017_));
  NO2        u0995(.A(men_men_n661_), .B(men_men_n106_), .Y(men_men_n1018_));
  AOI220     u0996(.A0(men_men_n1018_), .A1(i_0_), .B0(men_men_n1017_), .B1(men_men_n684_), .Y(men_men_n1019_));
  OAI220     u0997(.A0(men_men_n1019_), .A1(men_men_n84_), .B0(men_men_n1015_), .B1(men_men_n175_), .Y(men_men_n1020_));
  NO3        u0998(.A(men_men_n1020_), .B(men_men_n1013_), .C(men_men_n568_), .Y(men_men_n1021_));
  NA4        u0999(.A(men_men_n1021_), .B(men_men_n1008_), .C(men_men_n1002_), .D(men_men_n999_), .Y(men_men_n1022_));
  NO3        u1000(.A(men_men_n1022_), .B(men_men_n995_), .C(men_men_n964_), .Y(men_men_n1023_));
  NO2        u1001(.A(men_men_n937_), .B(men_men_n794_), .Y(men_men_n1024_));
  NA2        u1002(.A(men_men_n71_), .B(men_men_n42_), .Y(men_men_n1025_));
  INV        u1003(.A(men_men_n1025_), .Y(men_men_n1026_));
  NO3        u1004(.A(men_men_n106_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n1027_));
  AO220      u1005(.A0(men_men_n1027_), .A1(men_men_n1026_), .B0(men_men_n1024_), .B1(men_men_n177_), .Y(men_men_n1028_));
  AOI210     u1006(.A0(men_men_n861_), .A1(men_men_n753_), .B0(men_men_n982_), .Y(men_men_n1029_));
  AOI210     u1007(.A0(men_men_n1028_), .A1(men_men_n370_), .B0(men_men_n1029_), .Y(men_men_n1030_));
  NA2        u1008(.A(men_men_n805_), .B(men_men_n147_), .Y(men_men_n1031_));
  INV        u1009(.A(men_men_n1031_), .Y(men_men_n1032_));
  NA3        u1010(.A(men_men_n1032_), .B(men_men_n740_), .C(men_men_n71_), .Y(men_men_n1033_));
  NO2        u1011(.A(men_men_n878_), .B(men_men_n431_), .Y(men_men_n1034_));
  NA3        u1012(.A(men_men_n909_), .B(i_2_), .C(men_men_n46_), .Y(men_men_n1035_));
  NA2        u1013(.A(men_men_n910_), .B(i_9_), .Y(men_men_n1036_));
  AOI210     u1014(.A0(men_men_n1035_), .A1(men_men_n541_), .B0(men_men_n1036_), .Y(men_men_n1037_));
  OAI210     u1015(.A0(men_men_n253_), .A1(i_9_), .B0(men_men_n238_), .Y(men_men_n1038_));
  AOI210     u1016(.A0(men_men_n1038_), .A1(men_men_n945_), .B0(men_men_n155_), .Y(men_men_n1039_));
  NO3        u1017(.A(men_men_n1039_), .B(men_men_n1037_), .C(men_men_n1034_), .Y(men_men_n1040_));
  NA3        u1018(.A(men_men_n1040_), .B(men_men_n1033_), .C(men_men_n1030_), .Y(men_men_n1041_));
  NA2        u1019(.A(men_men_n997_), .B(men_men_n399_), .Y(men_men_n1042_));
  AOI210     u1020(.A0(men_men_n316_), .A1(men_men_n164_), .B0(men_men_n1042_), .Y(men_men_n1043_));
  NA3        u1021(.A(men_men_n37_), .B(men_men_n28_), .C(men_men_n42_), .Y(men_men_n1044_));
  NA2        u1022(.A(men_men_n969_), .B(men_men_n529_), .Y(men_men_n1045_));
  AOI210     u1023(.A0(men_men_n1044_), .A1(men_men_n164_), .B0(men_men_n1045_), .Y(men_men_n1046_));
  NO2        u1024(.A(men_men_n1046_), .B(men_men_n1043_), .Y(men_men_n1047_));
  NO3        u1025(.A(men_men_n955_), .B(men_men_n929_), .C(men_men_n194_), .Y(men_men_n1048_));
  AOI220     u1026(.A0(men_men_n1048_), .A1(i_11_), .B0(men_men_n624_), .B1(men_men_n73_), .Y(men_men_n1049_));
  INV        u1027(.A(men_men_n225_), .Y(men_men_n1050_));
  OAI220     u1028(.A0(men_men_n581_), .A1(men_men_n141_), .B0(men_men_n709_), .B1(men_men_n678_), .Y(men_men_n1051_));
  NA3        u1029(.A(men_men_n1051_), .B(men_men_n426_), .C(men_men_n1050_), .Y(men_men_n1052_));
  NA3        u1030(.A(men_men_n1052_), .B(men_men_n1049_), .C(men_men_n1047_), .Y(men_men_n1053_));
  NO2        u1031(.A(men_men_n251_), .B(men_men_n93_), .Y(men_men_n1054_));
  AOI210     u1032(.A0(men_men_n1054_), .A1(men_men_n1024_), .B0(men_men_n110_), .Y(men_men_n1055_));
  AOI220     u1033(.A0(men_men_n987_), .A1(men_men_n529_), .B0(men_men_n909_), .B1(men_men_n165_), .Y(men_men_n1056_));
  NA2        u1034(.A(men_men_n373_), .B(men_men_n179_), .Y(men_men_n1057_));
  OA220      u1035(.A0(men_men_n1057_), .A1(men_men_n1056_), .B0(men_men_n1055_), .B1(i_5_), .Y(men_men_n1058_));
  AOI210     u1036(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n178_), .Y(men_men_n1059_));
  NA2        u1037(.A(men_men_n1059_), .B(men_men_n1001_), .Y(men_men_n1060_));
  NA3        u1038(.A(men_men_n675_), .B(men_men_n189_), .C(men_men_n82_), .Y(men_men_n1061_));
  NA2        u1039(.A(men_men_n1061_), .B(men_men_n598_), .Y(men_men_n1062_));
  NO3        u1040(.A(men_men_n919_), .B(men_men_n52_), .C(men_men_n46_), .Y(men_men_n1063_));
  NA3        u1041(.A(men_men_n534_), .B(men_men_n527_), .C(men_men_n510_), .Y(men_men_n1064_));
  NO3        u1042(.A(men_men_n1064_), .B(men_men_n1063_), .C(men_men_n1062_), .Y(men_men_n1065_));
  NA3        u1043(.A(men_men_n417_), .B(men_men_n174_), .C(men_men_n173_), .Y(men_men_n1066_));
  NA3        u1044(.A(men_men_n969_), .B(men_men_n305_), .C(men_men_n238_), .Y(men_men_n1067_));
  NA2        u1045(.A(men_men_n1067_), .B(men_men_n1066_), .Y(men_men_n1068_));
  NA3        u1046(.A(men_men_n417_), .B(men_men_n354_), .C(men_men_n229_), .Y(men_men_n1069_));
  INV        u1047(.A(men_men_n1069_), .Y(men_men_n1070_));
  NOi31      u1048(.An(men_men_n416_), .B(men_men_n1025_), .C(men_men_n248_), .Y(men_men_n1071_));
  NO3        u1049(.A(men_men_n966_), .B(men_men_n225_), .C(men_men_n194_), .Y(men_men_n1072_));
  NO4        u1050(.A(men_men_n1072_), .B(men_men_n1071_), .C(men_men_n1070_), .D(men_men_n1068_), .Y(men_men_n1073_));
  NA4        u1051(.A(men_men_n1073_), .B(men_men_n1065_), .C(men_men_n1060_), .D(men_men_n1058_), .Y(men_men_n1074_));
  AOI210     u1052(.A0(men_men_n623_), .A1(men_men_n580_), .B0(men_men_n677_), .Y(men_men_n1075_));
  NO3        u1053(.A(men_men_n1075_), .B(men_men_n614_), .C(men_men_n367_), .Y(men_men_n1076_));
  NO2        u1054(.A(men_men_n84_), .B(i_5_), .Y(men_men_n1077_));
  NA3        u1055(.A(men_men_n910_), .B(men_men_n111_), .C(men_men_n126_), .Y(men_men_n1078_));
  INV        u1056(.A(men_men_n1078_), .Y(men_men_n1079_));
  AOI210     u1057(.A0(men_men_n1079_), .A1(men_men_n1077_), .B0(men_men_n1076_), .Y(men_men_n1080_));
  NA3        u1058(.A(men_men_n322_), .B(i_5_), .C(men_men_n197_), .Y(men_men_n1081_));
  NAi31      u1059(.An(men_men_n250_), .B(men_men_n1081_), .C(men_men_n251_), .Y(men_men_n1082_));
  NO4        u1060(.A(men_men_n248_), .B(men_men_n216_), .C(i_0_), .D(i_12_), .Y(men_men_n1083_));
  AOI220     u1061(.A0(men_men_n1083_), .A1(men_men_n1082_), .B0(men_men_n856_), .B1(men_men_n179_), .Y(men_men_n1084_));
  BUFFER     u1062(.A(men_men_n155_), .Y(men_men_n1085_));
  NO4        u1063(.A(men_men_n1085_), .B(i_12_), .C(men_men_n713_), .D(men_men_n133_), .Y(men_men_n1086_));
  NA2        u1064(.A(men_men_n1086_), .B(men_men_n225_), .Y(men_men_n1087_));
  NA3        u1065(.A(men_men_n99_), .B(men_men_n628_), .C(i_11_), .Y(men_men_n1088_));
  NO2        u1066(.A(men_men_n1088_), .B(men_men_n157_), .Y(men_men_n1089_));
  NA2        u1067(.A(men_men_n987_), .B(men_men_n509_), .Y(men_men_n1090_));
  NA2        u1068(.A(men_men_n62_), .B(men_men_n102_), .Y(men_men_n1091_));
  OAI220     u1069(.A0(men_men_n1091_), .A1(men_men_n1081_), .B0(men_men_n1090_), .B1(men_men_n741_), .Y(men_men_n1092_));
  AOI210     u1070(.A0(men_men_n1092_), .A1(men_men_n973_), .B0(men_men_n1089_), .Y(men_men_n1093_));
  NA4        u1071(.A(men_men_n1093_), .B(men_men_n1087_), .C(men_men_n1084_), .D(men_men_n1080_), .Y(men_men_n1094_));
  NO4        u1072(.A(men_men_n1094_), .B(men_men_n1074_), .C(men_men_n1053_), .D(men_men_n1041_), .Y(men_men_n1095_));
  OAI210     u1073(.A0(men_men_n881_), .A1(men_men_n874_), .B0(men_men_n35_), .Y(men_men_n1096_));
  NA3        u1074(.A(men_men_n981_), .B(men_men_n394_), .C(i_5_), .Y(men_men_n1097_));
  NA3        u1075(.A(men_men_n1097_), .B(men_men_n1096_), .C(men_men_n673_), .Y(men_men_n1098_));
  NA2        u1076(.A(men_men_n1098_), .B(men_men_n212_), .Y(men_men_n1099_));
  AN2        u1077(.A(men_men_n766_), .B(men_men_n395_), .Y(men_men_n1100_));
  NA2        u1078(.A(men_men_n190_), .B(men_men_n192_), .Y(men_men_n1101_));
  AO210      u1079(.A0(men_men_n1100_), .A1(men_men_n31_), .B0(men_men_n1101_), .Y(men_men_n1102_));
  OAI210     u1080(.A0(men_men_n677_), .A1(men_men_n675_), .B0(men_men_n335_), .Y(men_men_n1103_));
  NAi31      u1081(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1104_));
  AOI210     u1082(.A0(men_men_n119_), .A1(men_men_n68_), .B0(men_men_n1104_), .Y(men_men_n1105_));
  NO2        u1083(.A(men_men_n1105_), .B(men_men_n710_), .Y(men_men_n1106_));
  NA3        u1084(.A(men_men_n1106_), .B(men_men_n1103_), .C(men_men_n1102_), .Y(men_men_n1107_));
  NO2        u1085(.A(men_men_n499_), .B(men_men_n279_), .Y(men_men_n1108_));
  NO4        u1086(.A(men_men_n241_), .B(men_men_n146_), .C(men_men_n744_), .D(men_men_n35_), .Y(men_men_n1109_));
  NO3        u1087(.A(men_men_n1109_), .B(men_men_n1108_), .C(men_men_n947_), .Y(men_men_n1110_));
  OAI210     u1088(.A0(men_men_n1088_), .A1(men_men_n149_), .B0(men_men_n1110_), .Y(men_men_n1111_));
  AOI210     u1089(.A0(men_men_n1107_), .A1(men_men_n46_), .B0(men_men_n1111_), .Y(men_men_n1112_));
  AOI210     u1090(.A0(men_men_n1112_), .A1(men_men_n1099_), .B0(men_men_n71_), .Y(men_men_n1113_));
  NO2        u1091(.A(men_men_n621_), .B(men_men_n406_), .Y(men_men_n1114_));
  NO2        u1092(.A(men_men_n1114_), .B(men_men_n823_), .Y(men_men_n1115_));
  OAI210     u1093(.A0(men_men_n78_), .A1(men_men_n52_), .B0(men_men_n109_), .Y(men_men_n1116_));
  NA2        u1094(.A(men_men_n1116_), .B(men_men_n74_), .Y(men_men_n1117_));
  AOI210     u1095(.A0(men_men_n1059_), .A1(men_men_n969_), .B0(men_men_n988_), .Y(men_men_n1118_));
  AOI210     u1096(.A0(men_men_n1118_), .A1(men_men_n1117_), .B0(men_men_n744_), .Y(men_men_n1119_));
  INV        u1097(.A(men_men_n55_), .Y(men_men_n1120_));
  AOI220     u1098(.A0(men_men_n1120_), .A1(men_men_n74_), .B0(men_men_n368_), .B1(men_men_n265_), .Y(men_men_n1121_));
  NO2        u1099(.A(men_men_n1121_), .B(men_men_n245_), .Y(men_men_n1122_));
  NA3        u1100(.A(men_men_n97_), .B(men_men_n324_), .C(men_men_n29_), .Y(men_men_n1123_));
  INV        u1101(.A(men_men_n1123_), .Y(men_men_n1124_));
  NO3        u1102(.A(men_men_n1124_), .B(men_men_n1122_), .C(men_men_n1119_), .Y(men_men_n1125_));
  OAI210     u1103(.A0(men_men_n281_), .A1(men_men_n160_), .B0(men_men_n87_), .Y(men_men_n1126_));
  NA3        u1104(.A(men_men_n827_), .B(men_men_n305_), .C(men_men_n78_), .Y(men_men_n1127_));
  AOI210     u1105(.A0(men_men_n1127_), .A1(men_men_n1126_), .B0(i_11_), .Y(men_men_n1128_));
  NA2        u1106(.A(men_men_n668_), .B(men_men_n222_), .Y(men_men_n1129_));
  OAI210     u1107(.A0(men_men_n1129_), .A1(men_men_n981_), .B0(men_men_n212_), .Y(men_men_n1130_));
  NA2        u1108(.A(men_men_n166_), .B(i_5_), .Y(men_men_n1131_));
  AOI210     u1109(.A0(men_men_n1130_), .A1(men_men_n836_), .B0(men_men_n1131_), .Y(men_men_n1132_));
  NO3        u1110(.A(men_men_n57_), .B(men_men_n56_), .C(i_4_), .Y(men_men_n1133_));
  OAI210     u1111(.A0(men_men_n992_), .A1(men_men_n324_), .B0(men_men_n1133_), .Y(men_men_n1134_));
  NO2        u1112(.A(men_men_n1134_), .B(men_men_n794_), .Y(men_men_n1135_));
  NO4        u1113(.A(men_men_n1016_), .B(men_men_n517_), .C(men_men_n262_), .D(men_men_n261_), .Y(men_men_n1136_));
  NO2        u1114(.A(men_men_n1136_), .B(men_men_n618_), .Y(men_men_n1137_));
  NO2        u1115(.A(men_men_n877_), .B(men_men_n387_), .Y(men_men_n1138_));
  AOI210     u1116(.A0(men_men_n1138_), .A1(men_men_n1137_), .B0(men_men_n38_), .Y(men_men_n1139_));
  NO4        u1117(.A(men_men_n1139_), .B(men_men_n1135_), .C(men_men_n1132_), .D(men_men_n1128_), .Y(men_men_n1140_));
  OAI210     u1118(.A0(men_men_n1125_), .A1(i_4_), .B0(men_men_n1140_), .Y(men_men_n1141_));
  NO3        u1119(.A(men_men_n1141_), .B(men_men_n1115_), .C(men_men_n1113_), .Y(men_men_n1142_));
  NA4        u1120(.A(men_men_n1142_), .B(men_men_n1095_), .C(men_men_n1023_), .D(men_men_n936_), .Y(men4));
  INV        u1121(.A(i_5_), .Y(men_men_n1146_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule