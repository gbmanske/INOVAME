//Benchmark atmr_alu4_1266_0.0156

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1045_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1057_, men_men_n1058_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NA3        o034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n57_));
  NO2        o035(.A(i_1_), .B(i_6_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  OAI210     o037(.A0(ori_ori_n59_), .A1(ori_ori_n58_), .B0(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n61_));
  NAi21      o039(.An(i_2_), .B(i_7_), .Y(ori_ori_n62_));
  INV        o040(.A(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NA3        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .C(ori_ori_n31_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_1_), .B(i_10_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(i_6_), .Y(ori_ori_n67_));
  NAi31      o045(.An(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n61_), .Y(ori_ori_n68_));
  NA2        o046(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_1_), .B(i_6_), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n71_), .B(ori_ori_n25_), .Y(ori_ori_n72_));
  INV        o050(.A(i_0_), .Y(ori_ori_n73_));
  NAi21      o051(.An(i_5_), .B(i_10_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_5_), .B(i_9_), .Y(ori_ori_n75_));
  AOI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n73_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  OAI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n68_), .B0(i_0_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_12_), .B(i_5_), .Y(ori_ori_n80_));
  NA2        o058(.A(i_2_), .B(i_8_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n81_), .B(ori_ori_n58_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_9_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_3_), .B(i_7_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(ori_ori_n63_), .Y(ori_ori_n85_));
  INV        o063(.A(i_6_), .Y(ori_ori_n86_));
  OR4        o064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NO2        o066(.A(i_2_), .B(i_7_), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n88_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  OAI210     o068(.A0(ori_ori_n85_), .A1(ori_ori_n82_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NAi21      o069(.An(i_6_), .B(i_10_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_6_), .B(i_9_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n93_), .A1(ori_ori_n92_), .B0(ori_ori_n63_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_2_), .B(i_6_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n96_), .B(ori_ori_n94_), .Y(ori_ori_n97_));
  AOI210     o075(.A0(ori_ori_n97_), .A1(ori_ori_n91_), .B0(ori_ori_n80_), .Y(ori_ori_n98_));
  AN3        o076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n99_));
  NAi21      o077(.An(i_6_), .B(i_11_), .Y(ori_ori_n100_));
  NO2        o078(.A(i_5_), .B(i_8_), .Y(ori_ori_n101_));
  NOi21      o079(.An(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  AOI220     o080(.A0(ori_ori_n102_), .A1(ori_ori_n62_), .B0(ori_ori_n99_), .B1(ori_ori_n32_), .Y(ori_ori_n103_));
  INV        o081(.A(i_7_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n46_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o083(.A(i_0_), .B(i_5_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n86_), .Y(ori_ori_n107_));
  NA2        o085(.A(i_12_), .B(i_3_), .Y(ori_ori_n108_));
  INV        o086(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NA3        o087(.A(ori_ori_n109_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n110_));
  NAi21      o088(.An(i_7_), .B(i_11_), .Y(ori_ori_n111_));
  NO3        o089(.A(ori_ori_n111_), .B(ori_ori_n92_), .C(ori_ori_n53_), .Y(ori_ori_n112_));
  AN2        o090(.A(i_2_), .B(i_10_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(i_7_), .Y(ori_ori_n114_));
  OR2        o092(.A(ori_ori_n80_), .B(ori_ori_n58_), .Y(ori_ori_n115_));
  NO2        o093(.A(i_8_), .B(ori_ori_n104_), .Y(ori_ori_n116_));
  NO3        o094(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(ori_ori_n114_), .Y(ori_ori_n117_));
  NA2        o095(.A(i_12_), .B(i_7_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n63_), .B(ori_ori_n26_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(i_0_), .Y(ori_ori_n120_));
  NA2        o098(.A(i_11_), .B(i_12_), .Y(ori_ori_n121_));
  OAI210     o099(.A0(ori_ori_n120_), .A1(ori_ori_n118_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n122_), .B(ori_ori_n117_), .Y(ori_ori_n123_));
  NAi41      o101(.An(ori_ori_n112_), .B(ori_ori_n123_), .C(ori_ori_n110_), .D(ori_ori_n103_), .Y(ori_ori_n124_));
  NOi21      o102(.An(i_1_), .B(i_5_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(i_11_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n127_));
  NA2        o105(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n127_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n129_), .B(ori_ori_n46_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n93_), .B(ori_ori_n92_), .Y(ori_ori_n131_));
  NAi21      o109(.An(i_3_), .B(i_8_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n62_), .Y(ori_ori_n133_));
  NOi31      o111(.An(ori_ori_n133_), .B(ori_ori_n131_), .C(ori_ori_n130_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_1_), .B(ori_ori_n86_), .Y(ori_ori_n135_));
  NO2        o113(.A(i_6_), .B(i_5_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(i_3_), .Y(ori_ori_n137_));
  AO210      o115(.A0(ori_ori_n137_), .A1(ori_ori_n47_), .B0(ori_ori_n135_), .Y(ori_ori_n138_));
  OAI220     o116(.A0(ori_ori_n138_), .A1(ori_ori_n111_), .B0(ori_ori_n134_), .B1(ori_ori_n126_), .Y(ori_ori_n139_));
  NO3        o117(.A(ori_ori_n139_), .B(ori_ori_n124_), .C(ori_ori_n98_), .Y(ori_ori_n140_));
  NA3        o118(.A(ori_ori_n140_), .B(ori_ori_n79_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o119(.A(ori_ori_n63_), .B(ori_ori_n37_), .Y(ori_ori_n142_));
  NA2        o120(.A(i_6_), .B(ori_ori_n25_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(ori_ori_n142_), .Y(ori_ori_n144_));
  NA4        o122(.A(ori_ori_n144_), .B(ori_ori_n77_), .C(ori_ori_n69_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o123(.A(i_8_), .B(i_7_), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n146_), .B(i_6_), .Y(ori_ori_n147_));
  NO2        o125(.A(i_12_), .B(i_13_), .Y(ori_ori_n148_));
  NAi21      o126(.An(i_5_), .B(i_11_), .Y(ori_ori_n149_));
  NOi21      o127(.An(ori_ori_n148_), .B(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o128(.A(i_0_), .B(i_1_), .Y(ori_ori_n151_));
  NA2        o129(.A(i_2_), .B(i_3_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n152_), .B(i_4_), .Y(ori_ori_n153_));
  NA3        o131(.A(ori_ori_n153_), .B(ori_ori_n151_), .C(ori_ori_n150_), .Y(ori_ori_n154_));
  OR2        o132(.A(ori_ori_n154_), .B(ori_ori_n25_), .Y(ori_ori_n155_));
  AN2        o133(.A(ori_ori_n148_), .B(ori_ori_n83_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n156_), .B(ori_ori_n27_), .Y(ori_ori_n157_));
  NA2        o135(.A(i_1_), .B(i_5_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n73_), .B(ori_ori_n46_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n159_), .B(ori_ori_n36_), .Y(ori_ori_n160_));
  NO3        o138(.A(ori_ori_n160_), .B(ori_ori_n158_), .C(ori_ori_n157_), .Y(ori_ori_n161_));
  OR2        o139(.A(i_0_), .B(i_1_), .Y(ori_ori_n162_));
  NO3        o140(.A(ori_ori_n162_), .B(ori_ori_n80_), .C(i_13_), .Y(ori_ori_n163_));
  NAi32      o141(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n164_));
  NAi21      o142(.An(ori_ori_n164_), .B(ori_ori_n163_), .Y(ori_ori_n165_));
  NOi21      o143(.An(i_4_), .B(i_10_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n166_), .B(ori_ori_n40_), .Y(ori_ori_n167_));
  NO2        o145(.A(i_3_), .B(i_5_), .Y(ori_ori_n168_));
  NO3        o146(.A(ori_ori_n73_), .B(i_2_), .C(i_1_), .Y(ori_ori_n169_));
  NA2        o147(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  OAI210     o148(.A0(ori_ori_n170_), .A1(ori_ori_n167_), .B0(ori_ori_n165_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n171_), .B(ori_ori_n161_), .Y(ori_ori_n172_));
  AOI210     o150(.A0(ori_ori_n172_), .A1(ori_ori_n155_), .B0(ori_ori_n147_), .Y(ori_ori_n173_));
  NA2        o151(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n174_));
  NOi21      o152(.An(i_4_), .B(i_9_), .Y(ori_ori_n175_));
  NOi21      o153(.An(i_11_), .B(i_13_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(ori_ori_n175_), .Y(ori_ori_n177_));
  NO2        o155(.A(i_4_), .B(i_5_), .Y(ori_ori_n178_));
  NAi21      o156(.An(i_12_), .B(i_11_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n179_), .B(i_13_), .Y(ori_ori_n180_));
  NA3        o158(.A(ori_ori_n180_), .B(ori_ori_n178_), .C(ori_ori_n83_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n73_), .B(ori_ori_n63_), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n182_), .B(ori_ori_n46_), .Y(ori_ori_n183_));
  NA2        o161(.A(ori_ori_n36_), .B(i_5_), .Y(ori_ori_n184_));
  NAi31      o162(.An(ori_ori_n184_), .B(ori_ori_n156_), .C(i_11_), .Y(ori_ori_n185_));
  NA2        o163(.A(i_3_), .B(i_5_), .Y(ori_ori_n186_));
  OR2        o164(.A(ori_ori_n186_), .B(ori_ori_n177_), .Y(ori_ori_n187_));
  AOI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n185_), .B0(ori_ori_n183_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n189_));
  NO2        o167(.A(i_13_), .B(i_10_), .Y(ori_ori_n190_));
  NO2        o168(.A(i_2_), .B(i_1_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n191_), .B(i_3_), .Y(ori_ori_n192_));
  NAi21      o170(.An(i_4_), .B(i_12_), .Y(ori_ori_n193_));
  INV        o171(.A(ori_ori_n188_), .Y(ori_ori_n194_));
  INV        o172(.A(i_8_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n195_), .B(i_7_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n196_), .B(i_6_), .Y(ori_ori_n197_));
  NO3        o175(.A(i_3_), .B(ori_ori_n86_), .C(ori_ori_n48_), .Y(ori_ori_n198_));
  NA2        o176(.A(ori_ori_n198_), .B(ori_ori_n116_), .Y(ori_ori_n199_));
  NO3        o177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n200_));
  NA3        o178(.A(ori_ori_n200_), .B(ori_ori_n40_), .C(ori_ori_n44_), .Y(ori_ori_n201_));
  NO3        o179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n202_));
  OAI210     o180(.A0(ori_ori_n99_), .A1(i_12_), .B0(ori_ori_n202_), .Y(ori_ori_n203_));
  AOI210     o181(.A0(ori_ori_n203_), .A1(ori_ori_n201_), .B0(ori_ori_n199_), .Y(ori_ori_n204_));
  NO2        o182(.A(i_3_), .B(i_8_), .Y(ori_ori_n205_));
  NO3        o183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n206_));
  NA3        o184(.A(ori_ori_n206_), .B(ori_ori_n205_), .C(ori_ori_n40_), .Y(ori_ori_n207_));
  NO2        o185(.A(ori_ori_n106_), .B(ori_ori_n58_), .Y(ori_ori_n208_));
  INV        o186(.A(ori_ori_n208_), .Y(ori_ori_n209_));
  NO2        o187(.A(i_13_), .B(i_9_), .Y(ori_ori_n210_));
  NAi21      o188(.An(i_12_), .B(i_3_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n212_));
  NO3        o190(.A(i_0_), .B(i_2_), .C(ori_ori_n63_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n209_), .B(ori_ori_n207_), .Y(ori_ori_n214_));
  AOI210     o192(.A0(ori_ori_n214_), .A1(i_7_), .B0(ori_ori_n204_), .Y(ori_ori_n215_));
  OAI220     o193(.A0(ori_ori_n215_), .A1(i_4_), .B0(ori_ori_n197_), .B1(ori_ori_n194_), .Y(ori_ori_n216_));
  NAi21      o194(.An(i_12_), .B(i_7_), .Y(ori_ori_n217_));
  NA3        o195(.A(i_13_), .B(ori_ori_n195_), .C(i_10_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  NA2        o197(.A(i_0_), .B(i_5_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n220_), .B(ori_ori_n107_), .Y(ori_ori_n221_));
  OAI220     o199(.A0(ori_ori_n221_), .A1(ori_ori_n192_), .B0(ori_ori_n183_), .B1(ori_ori_n137_), .Y(ori_ori_n222_));
  NAi31      o200(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n73_), .B(ori_ori_n26_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n46_), .B(ori_ori_n63_), .Y(ori_ori_n226_));
  NA3        o204(.A(ori_ori_n226_), .B(ori_ori_n225_), .C(ori_ori_n224_), .Y(ori_ori_n227_));
  INV        o205(.A(i_13_), .Y(ori_ori_n228_));
  NO2        o206(.A(i_12_), .B(ori_ori_n228_), .Y(ori_ori_n229_));
  NA3        o207(.A(ori_ori_n229_), .B(ori_ori_n200_), .C(ori_ori_n198_), .Y(ori_ori_n230_));
  OAI210     o208(.A0(ori_ori_n227_), .A1(ori_ori_n223_), .B0(ori_ori_n230_), .Y(ori_ori_n231_));
  AOI220     o209(.A0(ori_ori_n231_), .A1(ori_ori_n146_), .B0(ori_ori_n222_), .B1(ori_ori_n219_), .Y(ori_ori_n232_));
  NO2        o210(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n186_), .B(i_4_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n234_), .B(ori_ori_n233_), .Y(ori_ori_n235_));
  OR2        o213(.A(i_8_), .B(i_7_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n86_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n53_), .B(i_1_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n238_), .B(ori_ori_n237_), .Y(ori_ori_n239_));
  INV        o217(.A(i_12_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n44_), .B(ori_ori_n240_), .Y(ori_ori_n241_));
  NO3        o219(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n242_));
  NA2        o220(.A(i_2_), .B(i_1_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n239_), .B(ori_ori_n235_), .Y(ori_ori_n244_));
  NO3        o222(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n245_));
  NAi21      o223(.An(i_4_), .B(i_3_), .Y(ori_ori_n246_));
  NO2        o224(.A(ori_ori_n246_), .B(ori_ori_n75_), .Y(ori_ori_n247_));
  NO2        o225(.A(i_0_), .B(i_6_), .Y(ori_ori_n248_));
  NOi41      o226(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n249_), .B(ori_ori_n248_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n243_), .B(ori_ori_n186_), .Y(ori_ori_n251_));
  NA2        o229(.A(ori_ori_n244_), .B(ori_ori_n210_), .Y(ori_ori_n252_));
  NO2        o230(.A(i_11_), .B(ori_ori_n228_), .Y(ori_ori_n253_));
  NOi21      o231(.An(i_1_), .B(i_6_), .Y(ori_ori_n254_));
  NAi21      o232(.An(i_3_), .B(i_7_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n240_), .B(i_9_), .Y(ori_ori_n256_));
  OR4        o234(.A(ori_ori_n256_), .B(ori_ori_n255_), .C(ori_ori_n254_), .D(ori_ori_n189_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n48_), .B(ori_ori_n25_), .Y(ori_ori_n258_));
  NO2        o236(.A(i_12_), .B(i_3_), .Y(ori_ori_n259_));
  NA2        o237(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n260_));
  NA2        o238(.A(i_3_), .B(i_9_), .Y(ori_ori_n261_));
  NAi21      o239(.An(i_7_), .B(i_10_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n261_), .Y(ori_ori_n263_));
  NA3        o241(.A(ori_ori_n263_), .B(ori_ori_n260_), .C(ori_ori_n64_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n257_), .Y(ori_ori_n265_));
  NA3        o243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(ori_ori_n266_));
  INV        o244(.A(ori_ori_n147_), .Y(ori_ori_n267_));
  NA2        o245(.A(ori_ori_n240_), .B(i_13_), .Y(ori_ori_n268_));
  NO2        o246(.A(ori_ori_n268_), .B(ori_ori_n75_), .Y(ori_ori_n269_));
  AOI220     o247(.A0(ori_ori_n269_), .A1(ori_ori_n267_), .B0(ori_ori_n265_), .B1(ori_ori_n253_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n236_), .B(ori_ori_n37_), .Y(ori_ori_n271_));
  NA2        o249(.A(i_12_), .B(i_6_), .Y(ori_ori_n272_));
  OR2        o250(.A(i_13_), .B(i_9_), .Y(ori_ori_n273_));
  NO3        o251(.A(ori_ori_n273_), .B(ori_ori_n272_), .C(ori_ori_n48_), .Y(ori_ori_n274_));
  NO2        o252(.A(ori_ori_n246_), .B(i_2_), .Y(ori_ori_n275_));
  NA3        o253(.A(ori_ori_n275_), .B(ori_ori_n274_), .C(ori_ori_n44_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n253_), .B(i_9_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n260_), .B(ori_ori_n64_), .Y(ori_ori_n278_));
  OAI210     o256(.A0(ori_ori_n278_), .A1(ori_ori_n277_), .B0(ori_ori_n276_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n159_), .B(ori_ori_n63_), .Y(ori_ori_n280_));
  NO3        o258(.A(i_11_), .B(ori_ori_n228_), .C(ori_ori_n25_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n255_), .B(i_8_), .Y(ori_ori_n282_));
  NO2        o260(.A(i_6_), .B(ori_ori_n48_), .Y(ori_ori_n283_));
  NA3        o261(.A(ori_ori_n283_), .B(ori_ori_n282_), .C(ori_ori_n281_), .Y(ori_ori_n284_));
  NO3        o262(.A(ori_ori_n26_), .B(ori_ori_n86_), .C(i_5_), .Y(ori_ori_n285_));
  NA3        o263(.A(ori_ori_n285_), .B(ori_ori_n271_), .C(ori_ori_n229_), .Y(ori_ori_n286_));
  AOI210     o264(.A0(ori_ori_n286_), .A1(ori_ori_n284_), .B0(ori_ori_n280_), .Y(ori_ori_n287_));
  AOI210     o265(.A0(ori_ori_n279_), .A1(ori_ori_n271_), .B0(ori_ori_n287_), .Y(ori_ori_n288_));
  NA4        o266(.A(ori_ori_n288_), .B(ori_ori_n270_), .C(ori_ori_n252_), .D(ori_ori_n232_), .Y(ori_ori_n289_));
  NO3        o267(.A(i_12_), .B(ori_ori_n228_), .C(ori_ori_n37_), .Y(ori_ori_n290_));
  INV        o268(.A(ori_ori_n290_), .Y(ori_ori_n291_));
  NA2        o269(.A(i_8_), .B(ori_ori_n104_), .Y(ori_ori_n292_));
  NOi21      o270(.An(ori_ori_n168_), .B(ori_ori_n86_), .Y(ori_ori_n293_));
  NO3        o271(.A(i_0_), .B(ori_ori_n46_), .C(i_1_), .Y(ori_ori_n294_));
  AOI220     o272(.A0(ori_ori_n294_), .A1(ori_ori_n198_), .B0(ori_ori_n293_), .B1(ori_ori_n238_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n295_), .B(ori_ori_n292_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n243_), .B(i_0_), .Y(ori_ori_n297_));
  NA2        o275(.A(i_0_), .B(i_1_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(i_2_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n59_), .B(i_6_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n170_), .B(ori_ori_n147_), .Y(ori_ori_n301_));
  NO2        o279(.A(ori_ori_n301_), .B(ori_ori_n296_), .Y(ori_ori_n302_));
  NO2        o280(.A(i_3_), .B(i_10_), .Y(ori_ori_n303_));
  NA3        o281(.A(ori_ori_n303_), .B(ori_ori_n40_), .C(ori_ori_n44_), .Y(ori_ori_n304_));
  NO2        o282(.A(i_2_), .B(ori_ori_n104_), .Y(ori_ori_n305_));
  NA2        o283(.A(i_1_), .B(ori_ori_n36_), .Y(ori_ori_n306_));
  AN2        o284(.A(i_3_), .B(i_10_), .Y(ori_ori_n307_));
  NA4        o285(.A(ori_ori_n307_), .B(ori_ori_n200_), .C(ori_ori_n180_), .D(ori_ori_n178_), .Y(ori_ori_n308_));
  NO2        o286(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n302_), .B(ori_ori_n291_), .Y(ori_ori_n311_));
  NO4        o289(.A(ori_ori_n311_), .B(ori_ori_n289_), .C(ori_ori_n216_), .D(ori_ori_n173_), .Y(ori_ori_n312_));
  NO3        o290(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n59_), .B(ori_ori_n86_), .Y(ori_ori_n314_));
  NO3        o292(.A(i_6_), .B(ori_ori_n195_), .C(i_7_), .Y(ori_ori_n315_));
  NO2        o293(.A(i_2_), .B(i_3_), .Y(ori_ori_n316_));
  OR2        o294(.A(i_0_), .B(i_5_), .Y(ori_ori_n317_));
  NA2        o295(.A(ori_ori_n220_), .B(ori_ori_n317_), .Y(ori_ori_n318_));
  NA4        o296(.A(ori_ori_n318_), .B(ori_ori_n237_), .C(ori_ori_n316_), .D(i_1_), .Y(ori_ori_n319_));
  NA3        o297(.A(ori_ori_n297_), .B(ori_ori_n293_), .C(ori_ori_n116_), .Y(ori_ori_n320_));
  NAi21      o298(.An(i_8_), .B(i_7_), .Y(ori_ori_n321_));
  NO2        o299(.A(ori_ori_n321_), .B(i_6_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n162_), .B(ori_ori_n46_), .Y(ori_ori_n323_));
  NA3        o301(.A(ori_ori_n323_), .B(ori_ori_n322_), .C(ori_ori_n168_), .Y(ori_ori_n324_));
  NA3        o302(.A(ori_ori_n324_), .B(ori_ori_n320_), .C(ori_ori_n319_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n325_), .B(i_4_), .Y(ori_ori_n326_));
  NO2        o304(.A(i_12_), .B(i_10_), .Y(ori_ori_n327_));
  NOi21      o305(.An(i_5_), .B(i_0_), .Y(ori_ori_n328_));
  NA4        o306(.A(ori_ori_n84_), .B(ori_ori_n36_), .C(ori_ori_n86_), .D(i_8_), .Y(ori_ori_n329_));
  NO2        o307(.A(i_6_), .B(i_8_), .Y(ori_ori_n330_));
  NOi21      o308(.An(i_0_), .B(i_2_), .Y(ori_ori_n331_));
  AN2        o309(.A(ori_ori_n331_), .B(ori_ori_n330_), .Y(ori_ori_n332_));
  NO2        o310(.A(i_1_), .B(i_7_), .Y(ori_ori_n333_));
  INV        o311(.A(ori_ori_n326_), .Y(ori_ori_n334_));
  NO3        o312(.A(ori_ori_n236_), .B(ori_ori_n46_), .C(i_1_), .Y(ori_ori_n335_));
  NO3        o313(.A(ori_ori_n321_), .B(i_2_), .C(i_1_), .Y(ori_ori_n336_));
  OAI210     o314(.A0(ori_ori_n336_), .A1(ori_ori_n335_), .B0(i_6_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n254_), .B(ori_ori_n305_), .C(ori_ori_n195_), .Y(ori_ori_n338_));
  AOI210     o316(.A0(ori_ori_n338_), .A1(ori_ori_n337_), .B0(ori_ori_n318_), .Y(ori_ori_n339_));
  NOi21      o317(.An(ori_ori_n158_), .B(ori_ori_n107_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n340_), .B(ori_ori_n128_), .Y(ori_ori_n341_));
  OAI210     o319(.A0(ori_ori_n341_), .A1(ori_ori_n339_), .B0(i_3_), .Y(ori_ori_n342_));
  NO2        o320(.A(ori_ori_n298_), .B(ori_ori_n81_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n343_), .B(ori_ori_n136_), .Y(ori_ori_n344_));
  NO2        o322(.A(ori_ori_n344_), .B(i_3_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n195_), .B(i_9_), .Y(ori_ori_n346_));
  NA2        o324(.A(ori_ori_n346_), .B(ori_ori_n208_), .Y(ori_ori_n347_));
  NO2        o325(.A(ori_ori_n347_), .B(ori_ori_n46_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(ori_ori_n345_), .Y(ori_ori_n349_));
  AOI210     o327(.A0(ori_ori_n349_), .A1(ori_ori_n342_), .B0(ori_ori_n167_), .Y(ori_ori_n350_));
  AOI210     o328(.A0(ori_ori_n334_), .A1(ori_ori_n313_), .B0(ori_ori_n350_), .Y(ori_ori_n351_));
  NOi32      o329(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n352_));
  INV        o330(.A(ori_ori_n352_), .Y(ori_ori_n353_));
  NAi21      o331(.An(i_0_), .B(i_6_), .Y(ori_ori_n354_));
  NAi21      o332(.An(i_1_), .B(i_5_), .Y(ori_ori_n355_));
  NA2        o333(.A(ori_ori_n355_), .B(ori_ori_n354_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(ori_ori_n25_), .Y(ori_ori_n357_));
  OAI210     o335(.A0(ori_ori_n357_), .A1(ori_ori_n164_), .B0(ori_ori_n250_), .Y(ori_ori_n358_));
  NAi41      o336(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n359_));
  OAI220     o337(.A0(ori_ori_n359_), .A1(ori_ori_n355_), .B0(ori_ori_n223_), .B1(ori_ori_n164_), .Y(ori_ori_n360_));
  AOI210     o338(.A0(ori_ori_n359_), .A1(ori_ori_n164_), .B0(ori_ori_n162_), .Y(ori_ori_n361_));
  NOi32      o339(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n362_));
  NAi21      o340(.An(i_6_), .B(i_1_), .Y(ori_ori_n363_));
  OR2        o341(.A(ori_ori_n361_), .B(ori_ori_n360_), .Y(ori_ori_n364_));
  NO2        o342(.A(i_1_), .B(ori_ori_n104_), .Y(ori_ori_n365_));
  NAi21      o343(.An(i_3_), .B(i_4_), .Y(ori_ori_n366_));
  NO2        o344(.A(ori_ori_n366_), .B(i_9_), .Y(ori_ori_n367_));
  AN2        o345(.A(i_6_), .B(i_7_), .Y(ori_ori_n368_));
  OAI210     o346(.A0(ori_ori_n368_), .A1(ori_ori_n365_), .B0(ori_ori_n367_), .Y(ori_ori_n369_));
  NA2        o347(.A(i_2_), .B(i_7_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n366_), .B(i_10_), .Y(ori_ori_n371_));
  NA3        o349(.A(ori_ori_n371_), .B(ori_ori_n370_), .C(ori_ori_n248_), .Y(ori_ori_n372_));
  AOI210     o350(.A0(ori_ori_n372_), .A1(ori_ori_n369_), .B0(ori_ori_n189_), .Y(ori_ori_n373_));
  AOI210     o351(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n374_));
  OAI210     o352(.A0(ori_ori_n374_), .A1(ori_ori_n191_), .B0(ori_ori_n371_), .Y(ori_ori_n375_));
  AOI220     o353(.A0(ori_ori_n371_), .A1(ori_ori_n333_), .B0(ori_ori_n242_), .B1(ori_ori_n191_), .Y(ori_ori_n376_));
  AOI210     o354(.A0(ori_ori_n376_), .A1(ori_ori_n375_), .B0(i_5_), .Y(ori_ori_n377_));
  NO4        o355(.A(ori_ori_n377_), .B(ori_ori_n373_), .C(ori_ori_n364_), .D(ori_ori_n358_), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n378_), .B(ori_ori_n353_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n59_), .B(ori_ori_n25_), .Y(ori_ori_n380_));
  AN2        o358(.A(i_12_), .B(i_5_), .Y(ori_ori_n381_));
  NO2        o359(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n382_));
  NO2        o360(.A(i_11_), .B(i_6_), .Y(ori_ori_n383_));
  NO2        o361(.A(i_5_), .B(i_10_), .Y(ori_ori_n384_));
  NO2        o362(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n154_), .B(ori_ori_n86_), .Y(ori_ori_n386_));
  NA2        o364(.A(ori_ori_n386_), .B(ori_ori_n385_), .Y(ori_ori_n387_));
  NO3        o365(.A(ori_ori_n86_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n388_));
  NO2        o366(.A(i_3_), .B(ori_ori_n104_), .Y(ori_ori_n389_));
  NO2        o367(.A(i_11_), .B(i_12_), .Y(ori_ori_n390_));
  NAi21      o368(.An(i_13_), .B(i_0_), .Y(ori_ori_n391_));
  INV        o369(.A(ori_ori_n387_), .Y(ori_ori_n392_));
  NO3        o370(.A(i_1_), .B(i_12_), .C(ori_ori_n86_), .Y(ori_ori_n393_));
  NO2        o371(.A(i_0_), .B(i_11_), .Y(ori_ori_n394_));
  INV        o372(.A(i_5_), .Y(ori_ori_n395_));
  AN2        o373(.A(i_1_), .B(i_6_), .Y(ori_ori_n396_));
  NOi21      o374(.An(i_2_), .B(i_12_), .Y(ori_ori_n397_));
  NA2        o375(.A(ori_ori_n397_), .B(ori_ori_n396_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n395_), .Y(ori_ori_n399_));
  NA2        o377(.A(ori_ori_n146_), .B(i_9_), .Y(ori_ori_n400_));
  NO2        o378(.A(ori_ori_n400_), .B(i_4_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n399_), .B(ori_ori_n401_), .Y(ori_ori_n402_));
  NAi21      o380(.An(i_9_), .B(i_4_), .Y(ori_ori_n403_));
  OR2        o381(.A(i_13_), .B(i_10_), .Y(ori_ori_n404_));
  NO3        o382(.A(ori_ori_n404_), .B(ori_ori_n121_), .C(ori_ori_n403_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n177_), .B(ori_ori_n127_), .Y(ori_ori_n406_));
  OR2        o384(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n104_), .B(ori_ori_n25_), .Y(ori_ori_n408_));
  NA2        o386(.A(ori_ori_n290_), .B(ori_ori_n408_), .Y(ori_ori_n409_));
  NA2        o387(.A(ori_ori_n283_), .B(ori_ori_n213_), .Y(ori_ori_n410_));
  OAI220     o388(.A0(ori_ori_n410_), .A1(ori_ori_n407_), .B0(ori_ori_n409_), .B1(ori_ori_n340_), .Y(ori_ori_n411_));
  INV        o389(.A(ori_ori_n411_), .Y(ori_ori_n412_));
  AOI210     o390(.A0(ori_ori_n412_), .A1(ori_ori_n402_), .B0(ori_ori_n26_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n320_), .B(ori_ori_n319_), .Y(ori_ori_n414_));
  AOI220     o392(.A0(ori_ori_n300_), .A1(ori_ori_n294_), .B0(ori_ori_n297_), .B1(ori_ori_n314_), .Y(ori_ori_n415_));
  NO2        o393(.A(ori_ori_n415_), .B(ori_ori_n174_), .Y(ori_ori_n416_));
  NO2        o394(.A(ori_ori_n186_), .B(ori_ori_n86_), .Y(ori_ori_n417_));
  AOI220     o395(.A0(ori_ori_n417_), .A1(ori_ori_n299_), .B0(ori_ori_n285_), .B1(ori_ori_n213_), .Y(ori_ori_n418_));
  NO2        o396(.A(ori_ori_n418_), .B(ori_ori_n292_), .Y(ori_ori_n419_));
  NO3        o397(.A(ori_ori_n419_), .B(ori_ori_n416_), .C(ori_ori_n414_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n198_), .B(ori_ori_n99_), .Y(ori_ori_n421_));
  NA3        o399(.A(ori_ori_n323_), .B(ori_ori_n168_), .C(ori_ori_n86_), .Y(ori_ori_n422_));
  AOI210     o400(.A0(ori_ori_n422_), .A1(ori_ori_n421_), .B0(ori_ori_n321_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n195_), .B(i_10_), .Y(ori_ori_n424_));
  NA3        o402(.A(ori_ori_n260_), .B(ori_ori_n64_), .C(i_2_), .Y(ori_ori_n425_));
  NA2        o403(.A(ori_ori_n300_), .B(ori_ori_n238_), .Y(ori_ori_n426_));
  OAI220     o404(.A0(ori_ori_n426_), .A1(ori_ori_n186_), .B0(ori_ori_n425_), .B1(ori_ori_n424_), .Y(ori_ori_n427_));
  NO2        o405(.A(ori_ori_n427_), .B(ori_ori_n423_), .Y(ori_ori_n428_));
  AOI210     o406(.A0(ori_ori_n428_), .A1(ori_ori_n420_), .B0(ori_ori_n277_), .Y(ori_ori_n429_));
  NO4        o407(.A(ori_ori_n429_), .B(ori_ori_n413_), .C(ori_ori_n392_), .D(ori_ori_n379_), .Y(ori_ori_n430_));
  NO2        o408(.A(ori_ori_n63_), .B(i_4_), .Y(ori_ori_n431_));
  NO2        o409(.A(ori_ori_n73_), .B(i_13_), .Y(ori_ori_n432_));
  NA3        o410(.A(ori_ori_n432_), .B(ori_ori_n431_), .C(i_2_), .Y(ori_ori_n433_));
  NO2        o411(.A(i_10_), .B(i_9_), .Y(ori_ori_n434_));
  NAi21      o412(.An(i_12_), .B(i_8_), .Y(ori_ori_n435_));
  NO2        o413(.A(ori_ori_n435_), .B(i_3_), .Y(ori_ori_n436_));
  NA2        o414(.A(ori_ori_n436_), .B(ori_ori_n434_), .Y(ori_ori_n437_));
  NO2        o415(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n438_), .B(ori_ori_n107_), .Y(ori_ori_n439_));
  OAI220     o417(.A0(ori_ori_n439_), .A1(ori_ori_n207_), .B0(ori_ori_n437_), .B1(ori_ori_n433_), .Y(ori_ori_n440_));
  NA2        o418(.A(ori_ori_n310_), .B(i_0_), .Y(ori_ori_n441_));
  NO3        o419(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n272_), .B(ori_ori_n100_), .Y(ori_ori_n443_));
  NA2        o421(.A(ori_ori_n443_), .B(ori_ori_n442_), .Y(ori_ori_n444_));
  NA2        o422(.A(i_8_), .B(i_9_), .Y(ori_ori_n445_));
  AOI210     o423(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n446_));
  OR2        o424(.A(ori_ori_n446_), .B(ori_ori_n445_), .Y(ori_ori_n447_));
  NA2        o425(.A(ori_ori_n290_), .B(ori_ori_n208_), .Y(ori_ori_n448_));
  NO2        o426(.A(ori_ori_n448_), .B(ori_ori_n447_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n253_), .B(ori_ori_n309_), .Y(ori_ori_n450_));
  NO3        o428(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n451_));
  INV        o429(.A(ori_ori_n451_), .Y(ori_ori_n452_));
  NA3        o430(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n453_));
  NA4        o431(.A(ori_ori_n149_), .B(ori_ori_n119_), .C(ori_ori_n80_), .D(ori_ori_n23_), .Y(ori_ori_n454_));
  OAI220     o432(.A0(ori_ori_n454_), .A1(ori_ori_n453_), .B0(ori_ori_n452_), .B1(ori_ori_n450_), .Y(ori_ori_n455_));
  NO3        o433(.A(ori_ori_n455_), .B(ori_ori_n449_), .C(ori_ori_n440_), .Y(ori_ori_n456_));
  NA2        o434(.A(ori_ori_n99_), .B(i_13_), .Y(ori_ori_n457_));
  NA2        o435(.A(ori_ori_n417_), .B(ori_ori_n380_), .Y(ori_ori_n458_));
  NO2        o436(.A(i_2_), .B(i_13_), .Y(ori_ori_n459_));
  NO2        o437(.A(ori_ori_n458_), .B(ori_ori_n457_), .Y(ori_ori_n460_));
  NO3        o438(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n461_));
  NO2        o439(.A(i_6_), .B(i_7_), .Y(ori_ori_n462_));
  NO2        o440(.A(i_11_), .B(i_1_), .Y(ori_ori_n463_));
  NOi21      o441(.An(i_2_), .B(i_7_), .Y(ori_ori_n464_));
  NO2        o442(.A(i_3_), .B(ori_ori_n195_), .Y(ori_ori_n465_));
  NO2        o443(.A(i_6_), .B(i_10_), .Y(ori_ori_n466_));
  NA4        o444(.A(ori_ori_n466_), .B(ori_ori_n313_), .C(ori_ori_n465_), .D(ori_ori_n240_), .Y(ori_ori_n467_));
  NO2        o445(.A(ori_ori_n467_), .B(ori_ori_n160_), .Y(ori_ori_n468_));
  NA3        o446(.A(ori_ori_n249_), .B(ori_ori_n176_), .C(ori_ori_n136_), .Y(ori_ori_n469_));
  NA2        o447(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n470_));
  NO2        o448(.A(ori_ori_n162_), .B(i_3_), .Y(ori_ori_n471_));
  NAi31      o449(.An(ori_ori_n470_), .B(ori_ori_n471_), .C(ori_ori_n229_), .Y(ori_ori_n472_));
  NA3        o450(.A(ori_ori_n385_), .B(ori_ori_n182_), .C(ori_ori_n153_), .Y(ori_ori_n473_));
  NA3        o451(.A(ori_ori_n473_), .B(ori_ori_n472_), .C(ori_ori_n469_), .Y(ori_ori_n474_));
  NO3        o452(.A(ori_ori_n474_), .B(ori_ori_n468_), .C(ori_ori_n460_), .Y(ori_ori_n475_));
  NA2        o453(.A(ori_ori_n442_), .B(ori_ori_n381_), .Y(ori_ori_n476_));
  NA2        o454(.A(ori_ori_n451_), .B(ori_ori_n384_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n477_), .B(ori_ori_n227_), .Y(ori_ori_n478_));
  NAi21      o456(.An(ori_ori_n218_), .B(ori_ori_n390_), .Y(ori_ori_n479_));
  NA2        o457(.A(ori_ori_n333_), .B(ori_ori_n220_), .Y(ori_ori_n480_));
  NO2        o458(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n481_));
  NO2        o459(.A(i_0_), .B(ori_ori_n86_), .Y(ori_ori_n482_));
  NA3        o460(.A(ori_ori_n482_), .B(ori_ori_n481_), .C(ori_ori_n146_), .Y(ori_ori_n483_));
  OR3        o461(.A(ori_ori_n306_), .B(ori_ori_n38_), .C(ori_ori_n46_), .Y(ori_ori_n484_));
  OAI220     o462(.A0(ori_ori_n484_), .A1(ori_ori_n483_), .B0(ori_ori_n480_), .B1(ori_ori_n479_), .Y(ori_ori_n485_));
  NA2        o463(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n486_));
  NA2        o464(.A(ori_ori_n313_), .B(ori_ori_n242_), .Y(ori_ori_n487_));
  OAI220     o465(.A0(ori_ori_n487_), .A1(ori_ori_n425_), .B0(ori_ori_n486_), .B1(ori_ori_n457_), .Y(ori_ori_n488_));
  NO3        o466(.A(ori_ori_n488_), .B(ori_ori_n485_), .C(ori_ori_n478_), .Y(ori_ori_n489_));
  NA3        o467(.A(ori_ori_n489_), .B(ori_ori_n475_), .C(ori_ori_n456_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n126_), .B(ori_ori_n115_), .Y(ori_ori_n491_));
  AN2        o469(.A(ori_ori_n491_), .B(ori_ori_n442_), .Y(ori_ori_n492_));
  NA2        o470(.A(ori_ori_n313_), .B(ori_ori_n169_), .Y(ori_ori_n493_));
  OAI210     o471(.A0(ori_ori_n493_), .A1(ori_ori_n235_), .B0(ori_ori_n308_), .Y(ori_ori_n494_));
  AOI220     o472(.A0(ori_ori_n494_), .A1(ori_ori_n322_), .B0(ori_ori_n492_), .B1(ori_ori_n310_), .Y(ori_ori_n495_));
  NA4        o473(.A(ori_ori_n432_), .B(ori_ori_n431_), .C(ori_ori_n205_), .D(i_2_), .Y(ori_ori_n496_));
  INV        o474(.A(ori_ori_n496_), .Y(ori_ori_n497_));
  NA2        o475(.A(ori_ori_n381_), .B(ori_ori_n228_), .Y(ori_ori_n498_));
  NA2        o476(.A(ori_ori_n368_), .B(ori_ori_n362_), .Y(ori_ori_n499_));
  OR2        o477(.A(ori_ori_n498_), .B(ori_ori_n499_), .Y(ori_ori_n500_));
  NO2        o478(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n501_));
  AOI210     o479(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n405_), .Y(ori_ori_n502_));
  NA2        o480(.A(ori_ori_n502_), .B(ori_ori_n500_), .Y(ori_ori_n503_));
  AOI210     o481(.A0(ori_ori_n497_), .A1(ori_ori_n206_), .B0(ori_ori_n503_), .Y(ori_ori_n504_));
  NA2        o482(.A(ori_ori_n260_), .B(ori_ori_n64_), .Y(ori_ori_n505_));
  OAI210     o483(.A0(i_8_), .A1(ori_ori_n505_), .B0(ori_ori_n138_), .Y(ori_ori_n506_));
  AOI210     o484(.A0(ori_ori_n196_), .A1(i_9_), .B0(ori_ori_n271_), .Y(ori_ori_n507_));
  NO2        o485(.A(ori_ori_n507_), .B(ori_ori_n201_), .Y(ori_ori_n508_));
  OR2        o486(.A(ori_ori_n186_), .B(i_4_), .Y(ori_ori_n509_));
  NO2        o487(.A(ori_ori_n509_), .B(ori_ori_n86_), .Y(ori_ori_n510_));
  AOI220     o488(.A0(ori_ori_n510_), .A1(ori_ori_n508_), .B0(ori_ori_n506_), .B1(ori_ori_n406_), .Y(ori_ori_n511_));
  NA3        o489(.A(ori_ori_n511_), .B(ori_ori_n504_), .C(ori_ori_n495_), .Y(ori_ori_n512_));
  NO2        o490(.A(i_12_), .B(ori_ori_n195_), .Y(ori_ori_n513_));
  NA2        o491(.A(ori_ori_n513_), .B(ori_ori_n228_), .Y(ori_ori_n514_));
  NO2        o492(.A(i_8_), .B(i_7_), .Y(ori_ori_n515_));
  OAI210     o493(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(ori_ori_n516_));
  NA2        o494(.A(ori_ori_n516_), .B(ori_ori_n226_), .Y(ori_ori_n517_));
  AOI220     o495(.A0(ori_ori_n323_), .A1(ori_ori_n40_), .B0(ori_ori_n238_), .B1(ori_ori_n210_), .Y(ori_ori_n518_));
  OAI220     o496(.A0(ori_ori_n518_), .A1(ori_ori_n509_), .B0(ori_ori_n517_), .B1(ori_ori_n246_), .Y(ori_ori_n519_));
  NA2        o497(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n520_));
  NO2        o498(.A(ori_ori_n520_), .B(i_6_), .Y(ori_ori_n521_));
  NA3        o499(.A(ori_ori_n521_), .B(ori_ori_n519_), .C(ori_ori_n515_), .Y(ori_ori_n522_));
  AOI220     o500(.A0(ori_ori_n417_), .A1(ori_ori_n323_), .B0(ori_ori_n251_), .B1(ori_ori_n248_), .Y(ori_ori_n523_));
  OAI220     o501(.A0(ori_ori_n523_), .A1(ori_ori_n268_), .B0(ori_ori_n457_), .B1(ori_ori_n137_), .Y(ori_ori_n524_));
  NA2        o502(.A(ori_ori_n524_), .B(ori_ori_n271_), .Y(ori_ori_n525_));
  NOi31      o503(.An(ori_ori_n297_), .B(ori_ori_n304_), .C(ori_ori_n184_), .Y(ori_ori_n526_));
  NA3        o504(.A(ori_ori_n307_), .B(ori_ori_n178_), .C(ori_ori_n99_), .Y(ori_ori_n527_));
  OAI210     o505(.A0(ori_ori_n1013_), .A1(ori_ori_n526_), .B0(ori_ori_n451_), .Y(ori_ori_n528_));
  NA3        o506(.A(ori_ori_n528_), .B(ori_ori_n525_), .C(ori_ori_n522_), .Y(ori_ori_n529_));
  NA3        o507(.A(ori_ori_n220_), .B(ori_ori_n71_), .C(ori_ori_n44_), .Y(ori_ori_n530_));
  NA2        o508(.A(ori_ori_n290_), .B(ori_ori_n84_), .Y(ori_ori_n531_));
  AOI210     o509(.A0(ori_ori_n530_), .A1(ori_ori_n344_), .B0(ori_ori_n531_), .Y(ori_ori_n532_));
  NA2        o510(.A(ori_ori_n226_), .B(ori_ori_n225_), .Y(ori_ori_n533_));
  NA2        o511(.A(ori_ori_n434_), .B(ori_ori_n224_), .Y(ori_ori_n534_));
  NO2        o512(.A(ori_ori_n533_), .B(ori_ori_n534_), .Y(ori_ori_n535_));
  AOI210     o513(.A0(ori_ori_n363_), .A1(ori_ori_n46_), .B0(ori_ori_n365_), .Y(ori_ori_n536_));
  NA2        o514(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n537_));
  NA3        o515(.A(ori_ori_n513_), .B(ori_ori_n281_), .C(ori_ori_n537_), .Y(ori_ori_n538_));
  NO2        o516(.A(ori_ori_n536_), .B(ori_ori_n538_), .Y(ori_ori_n539_));
  NO3        o517(.A(ori_ori_n539_), .B(ori_ori_n535_), .C(ori_ori_n532_), .Y(ori_ori_n540_));
  NO4        o518(.A(ori_ori_n254_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n541_));
  NO3        o519(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n542_));
  NO2        o520(.A(ori_ori_n236_), .B(ori_ori_n36_), .Y(ori_ori_n543_));
  NO2        o521(.A(ori_ori_n404_), .B(i_1_), .Y(ori_ori_n544_));
  NOi31      o522(.An(ori_ori_n544_), .B(ori_ori_n443_), .C(ori_ori_n73_), .Y(ori_ori_n545_));
  AN4        o523(.A(ori_ori_n545_), .B(ori_ori_n401_), .C(ori_ori_n481_), .D(i_2_), .Y(ori_ori_n546_));
  NO2        o524(.A(ori_ori_n415_), .B(ori_ori_n181_), .Y(ori_ori_n547_));
  NO2        o525(.A(ori_ori_n547_), .B(ori_ori_n546_), .Y(ori_ori_n548_));
  NOi21      o526(.An(i_10_), .B(i_6_), .Y(ori_ori_n549_));
  NO2        o527(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n550_));
  NO2        o528(.A(ori_ori_n118_), .B(ori_ori_n23_), .Y(ori_ori_n551_));
  NA2        o529(.A(ori_ori_n315_), .B(ori_ori_n169_), .Y(ori_ori_n552_));
  AOI220     o530(.A0(ori_ori_n552_), .A1(ori_ori_n426_), .B0(ori_ori_n187_), .B1(ori_ori_n185_), .Y(ori_ori_n553_));
  NO2        o531(.A(ori_ori_n200_), .B(ori_ori_n37_), .Y(ori_ori_n554_));
  NOi31      o532(.An(ori_ori_n150_), .B(ori_ori_n554_), .C(ori_ori_n329_), .Y(ori_ori_n555_));
  NO2        o533(.A(ori_ori_n555_), .B(ori_ori_n553_), .Y(ori_ori_n556_));
  INV        o534(.A(ori_ori_n316_), .Y(ori_ori_n557_));
  NO2        o535(.A(i_12_), .B(ori_ori_n86_), .Y(ori_ori_n558_));
  NA3        o536(.A(ori_ori_n558_), .B(ori_ori_n281_), .C(ori_ori_n537_), .Y(ori_ori_n559_));
  NA3        o537(.A(ori_ori_n383_), .B(ori_ori_n290_), .C(ori_ori_n220_), .Y(ori_ori_n560_));
  AOI210     o538(.A0(ori_ori_n560_), .A1(ori_ori_n559_), .B0(ori_ori_n557_), .Y(ori_ori_n561_));
  NA2        o539(.A(ori_ori_n178_), .B(i_0_), .Y(ori_ori_n562_));
  NO3        o540(.A(ori_ori_n562_), .B(ori_ori_n337_), .C(ori_ori_n304_), .Y(ori_ori_n563_));
  OR2        o541(.A(i_2_), .B(i_5_), .Y(ori_ori_n564_));
  OR2        o542(.A(ori_ori_n564_), .B(ori_ori_n396_), .Y(ori_ori_n565_));
  NO2        o543(.A(ori_ori_n565_), .B(ori_ori_n479_), .Y(ori_ori_n566_));
  NO3        o544(.A(ori_ori_n566_), .B(ori_ori_n563_), .C(ori_ori_n561_), .Y(ori_ori_n567_));
  NA4        o545(.A(ori_ori_n567_), .B(ori_ori_n556_), .C(ori_ori_n548_), .D(ori_ori_n540_), .Y(ori_ori_n568_));
  NO4        o546(.A(ori_ori_n568_), .B(ori_ori_n529_), .C(ori_ori_n512_), .D(ori_ori_n490_), .Y(ori_ori_n569_));
  NA4        o547(.A(ori_ori_n569_), .B(ori_ori_n430_), .C(ori_ori_n351_), .D(ori_ori_n312_), .Y(ori7));
  NO2        o548(.A(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n571_));
  NO2        o549(.A(ori_ori_n111_), .B(ori_ori_n92_), .Y(ori_ori_n572_));
  NA2        o550(.A(ori_ori_n382_), .B(ori_ori_n572_), .Y(ori_ori_n573_));
  NA2        o551(.A(ori_ori_n466_), .B(ori_ori_n84_), .Y(ori_ori_n574_));
  NA2        o552(.A(i_11_), .B(ori_ori_n195_), .Y(ori_ori_n575_));
  NA2        o553(.A(ori_ori_n148_), .B(ori_ori_n575_), .Y(ori_ori_n576_));
  OAI210     o554(.A0(ori_ori_n576_), .A1(ori_ori_n574_), .B0(ori_ori_n573_), .Y(ori_ori_n577_));
  NA3        o555(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n578_));
  NO2        o556(.A(ori_ori_n240_), .B(i_4_), .Y(ori_ori_n579_));
  NA2        o557(.A(ori_ori_n579_), .B(i_8_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n108_), .B(ori_ori_n578_), .Y(ori_ori_n581_));
  NA2        o559(.A(i_2_), .B(ori_ori_n86_), .Y(ori_ori_n582_));
  OAI210     o560(.A0(ori_ori_n89_), .A1(ori_ori_n205_), .B0(ori_ori_n206_), .Y(ori_ori_n583_));
  NO2        o561(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n584_));
  NA2        o562(.A(i_4_), .B(i_8_), .Y(ori_ori_n585_));
  AOI210     o563(.A0(ori_ori_n585_), .A1(ori_ori_n307_), .B0(ori_ori_n584_), .Y(ori_ori_n586_));
  OAI220     o564(.A0(ori_ori_n586_), .A1(ori_ori_n582_), .B0(ori_ori_n583_), .B1(i_13_), .Y(ori_ori_n587_));
  NO4        o565(.A(ori_ori_n587_), .B(ori_ori_n581_), .C(ori_ori_n577_), .D(ori_ori_n571_), .Y(ori_ori_n588_));
  AOI210     o566(.A0(ori_ori_n132_), .A1(ori_ori_n62_), .B0(i_10_), .Y(ori_ori_n589_));
  AOI210     o567(.A0(ori_ori_n589_), .A1(ori_ori_n240_), .B0(ori_ori_n166_), .Y(ori_ori_n590_));
  OR2        o568(.A(i_6_), .B(i_10_), .Y(ori_ori_n591_));
  NO2        o569(.A(ori_ori_n591_), .B(ori_ori_n23_), .Y(ori_ori_n592_));
  OR3        o570(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n593_));
  INV        o571(.A(ori_ori_n202_), .Y(ori_ori_n594_));
  INV        o572(.A(ori_ori_n592_), .Y(ori_ori_n595_));
  OA220      o573(.A0(ori_ori_n595_), .A1(ori_ori_n557_), .B0(ori_ori_n590_), .B1(ori_ori_n273_), .Y(ori_ori_n596_));
  AOI210     o574(.A0(ori_ori_n596_), .A1(ori_ori_n588_), .B0(ori_ori_n63_), .Y(ori_ori_n597_));
  NOi21      o575(.An(i_11_), .B(i_7_), .Y(ori_ori_n598_));
  AO210      o576(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n599_));
  NO2        o577(.A(ori_ori_n599_), .B(ori_ori_n598_), .Y(ori_ori_n600_));
  NA2        o578(.A(ori_ori_n600_), .B(ori_ori_n210_), .Y(ori_ori_n601_));
  NO2        o579(.A(ori_ori_n601_), .B(ori_ori_n63_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n88_), .B(ori_ori_n63_), .Y(ori_ori_n603_));
  AO210      o581(.A0(ori_ori_n603_), .A1(ori_ori_n376_), .B0(ori_ori_n41_), .Y(ori_ori_n604_));
  NO3        o582(.A(ori_ori_n262_), .B(ori_ori_n211_), .C(ori_ori_n575_), .Y(ori_ori_n605_));
  OAI210     o583(.A0(ori_ori_n605_), .A1(ori_ori_n229_), .B0(ori_ori_n63_), .Y(ori_ori_n606_));
  NA2        o584(.A(ori_ori_n397_), .B(ori_ori_n31_), .Y(ori_ori_n607_));
  OR2        o585(.A(ori_ori_n211_), .B(ori_ori_n111_), .Y(ori_ori_n608_));
  NA2        o586(.A(ori_ori_n608_), .B(ori_ori_n607_), .Y(ori_ori_n609_));
  NO2        o587(.A(ori_ori_n63_), .B(i_9_), .Y(ori_ori_n610_));
  NO2        o588(.A(ori_ori_n610_), .B(i_4_), .Y(ori_ori_n611_));
  NA2        o589(.A(ori_ori_n611_), .B(ori_ori_n609_), .Y(ori_ori_n612_));
  NO2        o590(.A(i_1_), .B(i_12_), .Y(ori_ori_n613_));
  NA3        o591(.A(ori_ori_n612_), .B(ori_ori_n606_), .C(ori_ori_n604_), .Y(ori_ori_n614_));
  OAI210     o592(.A0(ori_ori_n614_), .A1(ori_ori_n602_), .B0(i_6_), .Y(ori_ori_n615_));
  NO2        o593(.A(ori_ori_n240_), .B(ori_ori_n86_), .Y(ori_ori_n616_));
  NO2        o594(.A(ori_ori_n616_), .B(i_11_), .Y(ori_ori_n617_));
  INV        o595(.A(ori_ori_n444_), .Y(ori_ori_n618_));
  NO4        o596(.A(ori_ori_n217_), .B(ori_ori_n132_), .C(i_13_), .D(ori_ori_n86_), .Y(ori_ori_n619_));
  NA2        o597(.A(ori_ori_n619_), .B(ori_ori_n610_), .Y(ori_ori_n620_));
  NA2        o598(.A(ori_ori_n240_), .B(i_6_), .Y(ori_ori_n621_));
  NO3        o599(.A(ori_ori_n591_), .B(ori_ori_n236_), .C(ori_ori_n23_), .Y(ori_ori_n622_));
  AOI210     o600(.A0(i_1_), .A1(ori_ori_n263_), .B0(ori_ori_n622_), .Y(ori_ori_n623_));
  OAI210     o601(.A0(ori_ori_n623_), .A1(ori_ori_n44_), .B0(ori_ori_n620_), .Y(ori_ori_n624_));
  NA3        o602(.A(ori_ori_n515_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n625_));
  INV        o603(.A(i_2_), .Y(ori_ori_n626_));
  NA2        o604(.A(ori_ori_n142_), .B(i_9_), .Y(ori_ori_n627_));
  NA3        o605(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n628_));
  NO2        o606(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n629_));
  NA3        o607(.A(ori_ori_n629_), .B(ori_ori_n272_), .C(ori_ori_n44_), .Y(ori_ori_n630_));
  OAI220     o608(.A0(ori_ori_n630_), .A1(ori_ori_n628_), .B0(ori_ori_n627_), .B1(ori_ori_n626_), .Y(ori_ori_n631_));
  NA3        o609(.A(ori_ori_n610_), .B(ori_ori_n316_), .C(i_6_), .Y(ori_ori_n632_));
  NO2        o610(.A(ori_ori_n632_), .B(ori_ori_n23_), .Y(ori_ori_n633_));
  AOI210     o611(.A0(ori_ori_n463_), .A1(ori_ori_n408_), .B0(ori_ori_n245_), .Y(ori_ori_n634_));
  NO2        o612(.A(ori_ori_n634_), .B(ori_ori_n582_), .Y(ori_ori_n635_));
  NAi21      o613(.An(ori_ori_n625_), .B(ori_ori_n94_), .Y(ori_ori_n636_));
  NA2        o614(.A(ori_ori_n629_), .B(ori_ori_n272_), .Y(ori_ori_n637_));
  NO2        o615(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n638_));
  NA2        o616(.A(ori_ori_n638_), .B(ori_ori_n24_), .Y(ori_ori_n639_));
  OAI210     o617(.A0(ori_ori_n639_), .A1(ori_ori_n637_), .B0(ori_ori_n636_), .Y(ori_ori_n640_));
  OR4        o618(.A(ori_ori_n640_), .B(ori_ori_n635_), .C(ori_ori_n633_), .D(ori_ori_n631_), .Y(ori_ori_n641_));
  NO3        o619(.A(ori_ori_n641_), .B(ori_ori_n624_), .C(ori_ori_n618_), .Y(ori_ori_n642_));
  NO2        o620(.A(ori_ori_n240_), .B(ori_ori_n104_), .Y(ori_ori_n643_));
  NO2        o621(.A(ori_ori_n643_), .B(ori_ori_n598_), .Y(ori_ori_n644_));
  NA2        o622(.A(ori_ori_n644_), .B(i_1_), .Y(ori_ori_n645_));
  NO2        o623(.A(ori_ori_n645_), .B(ori_ori_n593_), .Y(ori_ori_n646_));
  NO2        o624(.A(ori_ori_n403_), .B(ori_ori_n86_), .Y(ori_ori_n647_));
  NA2        o625(.A(ori_ori_n646_), .B(ori_ori_n46_), .Y(ori_ori_n648_));
  NA2        o626(.A(i_3_), .B(ori_ori_n195_), .Y(ori_ori_n649_));
  NO2        o627(.A(ori_ori_n649_), .B(ori_ori_n118_), .Y(ori_ori_n650_));
  AN2        o628(.A(ori_ori_n650_), .B(ori_ori_n521_), .Y(ori_ori_n651_));
  NO2        o629(.A(ori_ori_n236_), .B(ori_ori_n44_), .Y(ori_ori_n652_));
  NO3        o630(.A(ori_ori_n652_), .B(ori_ori_n310_), .C(ori_ori_n241_), .Y(ori_ori_n653_));
  NO2        o631(.A(ori_ori_n121_), .B(ori_ori_n37_), .Y(ori_ori_n654_));
  NO2        o632(.A(ori_ori_n654_), .B(i_6_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n86_), .B(i_9_), .Y(ori_ori_n656_));
  NO2        o634(.A(ori_ori_n656_), .B(ori_ori_n63_), .Y(ori_ori_n657_));
  NO2        o635(.A(ori_ori_n657_), .B(ori_ori_n613_), .Y(ori_ori_n658_));
  NO4        o636(.A(ori_ori_n658_), .B(ori_ori_n655_), .C(ori_ori_n653_), .D(i_4_), .Y(ori_ori_n659_));
  NA2        o637(.A(i_1_), .B(i_3_), .Y(ori_ori_n660_));
  NO2        o638(.A(ori_ori_n445_), .B(ori_ori_n95_), .Y(ori_ori_n661_));
  AOI210     o639(.A0(ori_ori_n652_), .A1(ori_ori_n549_), .B0(ori_ori_n661_), .Y(ori_ori_n662_));
  NO2        o640(.A(ori_ori_n662_), .B(ori_ori_n660_), .Y(ori_ori_n663_));
  NO3        o641(.A(ori_ori_n663_), .B(ori_ori_n659_), .C(ori_ori_n651_), .Y(ori_ori_n664_));
  NA4        o642(.A(ori_ori_n664_), .B(ori_ori_n648_), .C(ori_ori_n642_), .D(ori_ori_n615_), .Y(ori_ori_n665_));
  NO3        o643(.A(i_11_), .B(i_3_), .C(i_7_), .Y(ori_ori_n666_));
  AN2        o644(.A(ori_ori_n249_), .B(ori_ori_n86_), .Y(ori_ori_n667_));
  NA2        o645(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n668_));
  NA3        o646(.A(ori_ori_n466_), .B(ori_ori_n501_), .C(ori_ori_n46_), .Y(ori_ori_n669_));
  NO3        o647(.A(ori_ori_n464_), .B(ori_ori_n585_), .C(ori_ori_n86_), .Y(ori_ori_n670_));
  NA2        o648(.A(ori_ori_n670_), .B(ori_ori_n25_), .Y(ori_ori_n671_));
  NA3        o649(.A(ori_ori_n671_), .B(ori_ori_n669_), .C(ori_ori_n668_), .Y(ori_ori_n672_));
  OAI210     o650(.A0(ori_ori_n672_), .A1(ori_ori_n667_), .B0(i_1_), .Y(ori_ori_n673_));
  AOI210     o651(.A0(ori_ori_n272_), .A1(ori_ori_n100_), .B0(i_1_), .Y(ori_ori_n674_));
  NO2        o652(.A(ori_ori_n366_), .B(i_2_), .Y(ori_ori_n675_));
  NA2        o653(.A(ori_ori_n675_), .B(ori_ori_n674_), .Y(ori_ori_n676_));
  OAI210     o654(.A0(ori_ori_n632_), .A1(ori_ori_n435_), .B0(ori_ori_n676_), .Y(ori_ori_n677_));
  INV        o655(.A(ori_ori_n677_), .Y(ori_ori_n678_));
  AOI210     o656(.A0(ori_ori_n678_), .A1(ori_ori_n673_), .B0(i_13_), .Y(ori_ori_n679_));
  OR2        o657(.A(i_11_), .B(i_7_), .Y(ori_ori_n680_));
  AOI210     o658(.A0(ori_ori_n628_), .A1(ori_ori_n54_), .B0(i_12_), .Y(ori_ori_n681_));
  NO2        o659(.A(ori_ori_n464_), .B(ori_ori_n24_), .Y(ori_ori_n682_));
  AOI220     o660(.A0(ori_ori_n682_), .A1(ori_ori_n647_), .B0(ori_ori_n249_), .B1(ori_ori_n135_), .Y(ori_ori_n683_));
  OAI220     o661(.A0(ori_ori_n683_), .A1(ori_ori_n41_), .B0(ori_ori_n1012_), .B1(ori_ori_n95_), .Y(ori_ori_n684_));
  INV        o662(.A(ori_ori_n684_), .Y(ori_ori_n685_));
  INV        o663(.A(ori_ori_n118_), .Y(ori_ori_n686_));
  AOI220     o664(.A0(ori_ori_n686_), .A1(ori_ori_n72_), .B0(ori_ori_n383_), .B1(ori_ori_n629_), .Y(ori_ori_n687_));
  NO2        o665(.A(ori_ori_n687_), .B(ori_ori_n246_), .Y(ori_ori_n688_));
  AOI210     o666(.A0(ori_ori_n435_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n689_));
  NOi31      o667(.An(ori_ori_n689_), .B(ori_ori_n574_), .C(ori_ori_n44_), .Y(ori_ori_n690_));
  NA2        o668(.A(ori_ori_n131_), .B(i_13_), .Y(ori_ori_n691_));
  NO2        o669(.A(ori_ori_n628_), .B(ori_ori_n118_), .Y(ori_ori_n692_));
  INV        o670(.A(ori_ori_n692_), .Y(ori_ori_n693_));
  OAI220     o671(.A0(ori_ori_n693_), .A1(ori_ori_n71_), .B0(ori_ori_n691_), .B1(ori_ori_n674_), .Y(ori_ori_n694_));
  NO3        o672(.A(ori_ori_n71_), .B(ori_ori_n32_), .C(ori_ori_n104_), .Y(ori_ori_n695_));
  NA2        o673(.A(ori_ori_n26_), .B(ori_ori_n195_), .Y(ori_ori_n696_));
  NA2        o674(.A(ori_ori_n696_), .B(i_7_), .Y(ori_ori_n697_));
  AOI220     o675(.A0(ori_ori_n383_), .A1(ori_ori_n629_), .B0(ori_ori_n94_), .B1(ori_ori_n105_), .Y(ori_ori_n698_));
  OAI220     o676(.A0(ori_ori_n698_), .A1(ori_ori_n580_), .B0(ori_ori_n1014_), .B1(ori_ori_n594_), .Y(ori_ori_n699_));
  NO4        o677(.A(ori_ori_n699_), .B(ori_ori_n694_), .C(ori_ori_n690_), .D(ori_ori_n688_), .Y(ori_ori_n700_));
  OR2        o678(.A(i_11_), .B(i_6_), .Y(ori_ori_n701_));
  NA3        o679(.A(ori_ori_n579_), .B(ori_ori_n696_), .C(i_7_), .Y(ori_ori_n702_));
  AOI210     o680(.A0(ori_ori_n702_), .A1(ori_ori_n693_), .B0(ori_ori_n701_), .Y(ori_ori_n703_));
  NA3        o681(.A(ori_ori_n397_), .B(ori_ori_n584_), .C(ori_ori_n100_), .Y(ori_ori_n704_));
  NA2        o682(.A(ori_ori_n617_), .B(i_13_), .Y(ori_ori_n705_));
  NA2        o683(.A(ori_ori_n105_), .B(ori_ori_n696_), .Y(ori_ori_n706_));
  NAi21      o684(.An(i_11_), .B(i_12_), .Y(ori_ori_n707_));
  NOi41      o685(.An(ori_ori_n114_), .B(ori_ori_n707_), .C(i_13_), .D(ori_ori_n86_), .Y(ori_ori_n708_));
  NA2        o686(.A(ori_ori_n708_), .B(ori_ori_n706_), .Y(ori_ori_n709_));
  NA3        o687(.A(ori_ori_n709_), .B(ori_ori_n705_), .C(ori_ori_n704_), .Y(ori_ori_n710_));
  OAI210     o688(.A0(ori_ori_n710_), .A1(ori_ori_n703_), .B0(ori_ori_n63_), .Y(ori_ori_n711_));
  NO2        o689(.A(i_2_), .B(i_12_), .Y(ori_ori_n712_));
  NA2        o690(.A(ori_ori_n365_), .B(ori_ori_n712_), .Y(ori_ori_n713_));
  NA2        o691(.A(i_8_), .B(ori_ori_n25_), .Y(ori_ori_n714_));
  NO3        o692(.A(ori_ori_n714_), .B(ori_ori_n382_), .C(ori_ori_n579_), .Y(ori_ori_n715_));
  OAI210     o693(.A0(ori_ori_n715_), .A1(ori_ori_n367_), .B0(ori_ori_n365_), .Y(ori_ori_n716_));
  NO2        o694(.A(ori_ori_n132_), .B(i_2_), .Y(ori_ori_n717_));
  NA2        o695(.A(ori_ori_n717_), .B(ori_ori_n613_), .Y(ori_ori_n718_));
  NA3        o696(.A(ori_ori_n718_), .B(ori_ori_n716_), .C(ori_ori_n713_), .Y(ori_ori_n719_));
  NA3        o697(.A(ori_ori_n719_), .B(ori_ori_n45_), .C(ori_ori_n228_), .Y(ori_ori_n720_));
  NA4        o698(.A(ori_ori_n720_), .B(ori_ori_n711_), .C(ori_ori_n700_), .D(ori_ori_n685_), .Y(ori_ori_n721_));
  OR4        o699(.A(ori_ori_n721_), .B(ori_ori_n679_), .C(ori_ori_n665_), .D(ori_ori_n597_), .Y(ori5));
  NA2        o700(.A(ori_ori_n644_), .B(ori_ori_n275_), .Y(ori_ori_n723_));
  AN2        o701(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n724_));
  NA3        o702(.A(ori_ori_n724_), .B(ori_ori_n712_), .C(ori_ori_n111_), .Y(ori_ori_n725_));
  NO2        o703(.A(ori_ori_n580_), .B(i_11_), .Y(ori_ori_n726_));
  NA2        o704(.A(ori_ori_n89_), .B(ori_ori_n726_), .Y(ori_ori_n727_));
  NA3        o705(.A(ori_ori_n727_), .B(ori_ori_n725_), .C(ori_ori_n723_), .Y(ori_ori_n728_));
  NO3        o706(.A(i_11_), .B(ori_ori_n240_), .C(i_13_), .Y(ori_ori_n729_));
  NO2        o707(.A(ori_ori_n128_), .B(ori_ori_n23_), .Y(ori_ori_n730_));
  NA2        o708(.A(i_12_), .B(i_8_), .Y(ori_ori_n731_));
  OAI210     o709(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n731_), .Y(ori_ori_n732_));
  INV        o710(.A(ori_ori_n434_), .Y(ori_ori_n733_));
  AOI220     o711(.A0(ori_ori_n316_), .A1(ori_ori_n551_), .B0(ori_ori_n732_), .B1(ori_ori_n730_), .Y(ori_ori_n734_));
  INV        o712(.A(ori_ori_n734_), .Y(ori_ori_n735_));
  NO2        o713(.A(ori_ori_n735_), .B(ori_ori_n728_), .Y(ori_ori_n736_));
  INV        o714(.A(ori_ori_n176_), .Y(ori_ori_n737_));
  INV        o715(.A(ori_ori_n249_), .Y(ori_ori_n738_));
  OAI210     o716(.A0(ori_ori_n675_), .A1(ori_ori_n436_), .B0(ori_ori_n114_), .Y(ori_ori_n739_));
  AOI210     o717(.A0(ori_ori_n739_), .A1(ori_ori_n738_), .B0(ori_ori_n737_), .Y(ori_ori_n740_));
  NO2        o718(.A(ori_ori_n445_), .B(ori_ori_n26_), .Y(ori_ori_n741_));
  NO2        o719(.A(ori_ori_n741_), .B(ori_ori_n408_), .Y(ori_ori_n742_));
  NA2        o720(.A(ori_ori_n742_), .B(i_2_), .Y(ori_ori_n743_));
  INV        o721(.A(ori_ori_n743_), .Y(ori_ori_n744_));
  AOI210     o722(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n404_), .Y(ori_ori_n745_));
  AOI210     o723(.A0(ori_ori_n745_), .A1(ori_ori_n744_), .B0(ori_ori_n740_), .Y(ori_ori_n746_));
  NO2        o724(.A(ori_ori_n193_), .B(ori_ori_n129_), .Y(ori_ori_n747_));
  OAI210     o725(.A0(ori_ori_n747_), .A1(ori_ori_n730_), .B0(i_2_), .Y(ori_ori_n748_));
  INV        o726(.A(ori_ori_n177_), .Y(ori_ori_n749_));
  NO3        o727(.A(ori_ori_n599_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n750_));
  AOI210     o728(.A0(ori_ori_n749_), .A1(ori_ori_n89_), .B0(ori_ori_n750_), .Y(ori_ori_n751_));
  AOI210     o729(.A0(ori_ori_n751_), .A1(ori_ori_n748_), .B0(ori_ori_n195_), .Y(ori_ori_n752_));
  OA210      o730(.A0(ori_ori_n600_), .A1(ori_ori_n130_), .B0(i_13_), .Y(ori_ori_n753_));
  NA2        o731(.A(ori_ori_n202_), .B(ori_ori_n205_), .Y(ori_ori_n754_));
  NA2        o732(.A(ori_ori_n156_), .B(ori_ori_n575_), .Y(ori_ori_n755_));
  AOI210     o733(.A0(ori_ori_n755_), .A1(ori_ori_n754_), .B0(ori_ori_n370_), .Y(ori_ori_n756_));
  AOI210     o734(.A0(ori_ori_n211_), .A1(ori_ori_n152_), .B0(ori_ori_n501_), .Y(ori_ori_n757_));
  NA2        o735(.A(ori_ori_n757_), .B(ori_ori_n408_), .Y(ori_ori_n758_));
  NO2        o736(.A(ori_ori_n105_), .B(ori_ori_n44_), .Y(ori_ori_n759_));
  INV        o737(.A(ori_ori_n305_), .Y(ori_ori_n760_));
  NA4        o738(.A(ori_ori_n760_), .B(ori_ori_n307_), .C(ori_ori_n128_), .D(ori_ori_n42_), .Y(ori_ori_n761_));
  OAI210     o739(.A0(ori_ori_n761_), .A1(ori_ori_n759_), .B0(ori_ori_n758_), .Y(ori_ori_n762_));
  NO4        o740(.A(ori_ori_n762_), .B(ori_ori_n756_), .C(ori_ori_n753_), .D(ori_ori_n752_), .Y(ori_ori_n763_));
  NA2        o741(.A(ori_ori_n551_), .B(ori_ori_n28_), .Y(ori_ori_n764_));
  NA2        o742(.A(ori_ori_n729_), .B(ori_ori_n282_), .Y(ori_ori_n765_));
  NA2        o743(.A(ori_ori_n765_), .B(ori_ori_n764_), .Y(ori_ori_n766_));
  NO2        o744(.A(ori_ori_n62_), .B(i_12_), .Y(ori_ori_n767_));
  NO2        o745(.A(ori_ori_n767_), .B(ori_ori_n130_), .Y(ori_ori_n768_));
  NO2        o746(.A(ori_ori_n768_), .B(ori_ori_n575_), .Y(ori_ori_n769_));
  AOI220     o747(.A0(ori_ori_n769_), .A1(ori_ori_n36_), .B0(ori_ori_n766_), .B1(ori_ori_n46_), .Y(ori_ori_n770_));
  NA4        o748(.A(ori_ori_n770_), .B(ori_ori_n763_), .C(ori_ori_n746_), .D(ori_ori_n736_), .Y(ori6));
  NO3        o749(.A(ori_ori_n258_), .B(ori_ori_n309_), .C(i_1_), .Y(ori_ori_n772_));
  NO2        o750(.A(ori_ori_n189_), .B(ori_ori_n143_), .Y(ori_ori_n773_));
  OAI210     o751(.A0(ori_ori_n773_), .A1(ori_ori_n772_), .B0(ori_ori_n717_), .Y(ori_ori_n774_));
  NA4        o752(.A(ori_ori_n384_), .B(ori_ori_n465_), .C(ori_ori_n71_), .D(ori_ori_n104_), .Y(ori_ori_n775_));
  INV        o753(.A(ori_ori_n775_), .Y(ori_ori_n776_));
  NO2        o754(.A(ori_ori_n223_), .B(ori_ori_n470_), .Y(ori_ori_n777_));
  NO2        o755(.A(ori_ori_n776_), .B(ori_ori_n328_), .Y(ori_ori_n778_));
  AO210      o756(.A0(ori_ori_n778_), .A1(ori_ori_n774_), .B0(i_12_), .Y(ori_ori_n779_));
  NA2        o757(.A(ori_ori_n558_), .B(ori_ori_n63_), .Y(ori_ori_n780_));
  BUFFER     o758(.A(ori_ori_n603_), .Y(ori_ori_n781_));
  NA2        o759(.A(ori_ori_n781_), .B(ori_ori_n780_), .Y(ori_ori_n782_));
  NA2        o760(.A(ori_ori_n782_), .B(ori_ori_n73_), .Y(ori_ori_n783_));
  INV        o761(.A(ori_ori_n327_), .Y(ori_ori_n784_));
  NA2        o762(.A(ori_ori_n75_), .B(ori_ori_n135_), .Y(ori_ori_n785_));
  INV        o763(.A(ori_ori_n128_), .Y(ori_ori_n786_));
  NA2        o764(.A(ori_ori_n786_), .B(ori_ori_n46_), .Y(ori_ori_n787_));
  AOI210     o765(.A0(ori_ori_n787_), .A1(ori_ori_n785_), .B0(ori_ori_n784_), .Y(ori_ori_n788_));
  NO3        o766(.A(ori_ori_n254_), .B(ori_ori_n136_), .C(i_9_), .Y(ori_ori_n789_));
  NA2        o767(.A(ori_ori_n789_), .B(ori_ori_n767_), .Y(ori_ori_n790_));
  AOI210     o768(.A0(ori_ori_n790_), .A1(ori_ori_n499_), .B0(ori_ori_n189_), .Y(ori_ori_n791_));
  NO2        o769(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n792_));
  NAi32      o770(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n793_));
  NO2        o771(.A(ori_ori_n701_), .B(ori_ori_n793_), .Y(ori_ori_n794_));
  OAI210     o772(.A0(ori_ori_n666_), .A1(ori_ori_n543_), .B0(ori_ori_n542_), .Y(ori_ori_n795_));
  NAi21      o773(.An(ori_ori_n794_), .B(ori_ori_n795_), .Y(ori_ori_n796_));
  OR3        o774(.A(ori_ori_n796_), .B(ori_ori_n791_), .C(ori_ori_n788_), .Y(ori_ori_n797_));
  NO2        o775(.A(ori_ori_n680_), .B(i_2_), .Y(ori_ori_n798_));
  NA2        o776(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n799_));
  NO2        o777(.A(ori_ori_n799_), .B(ori_ori_n396_), .Y(ori_ori_n800_));
  NA2        o778(.A(ori_ori_n800_), .B(ori_ori_n798_), .Y(ori_ori_n801_));
  AO220      o779(.A0(ori_ori_n356_), .A1(ori_ori_n346_), .B0(ori_ori_n388_), .B1(ori_ori_n575_), .Y(ori_ori_n802_));
  NA3        o780(.A(ori_ori_n802_), .B(ori_ori_n259_), .C(i_7_), .Y(ori_ori_n803_));
  OR2        o781(.A(ori_ori_n600_), .B(ori_ori_n436_), .Y(ori_ori_n804_));
  NA3        o782(.A(ori_ori_n804_), .B(ori_ori_n151_), .C(ori_ori_n69_), .Y(ori_ori_n805_));
  AO210      o783(.A0(ori_ori_n477_), .A1(ori_ori_n733_), .B0(ori_ori_n36_), .Y(ori_ori_n806_));
  NA4        o784(.A(ori_ori_n806_), .B(ori_ori_n805_), .C(ori_ori_n803_), .D(ori_ori_n801_), .Y(ori_ori_n807_));
  OAI210     o785(.A0(ori_ori_n616_), .A1(i_11_), .B0(ori_ori_n87_), .Y(ori_ori_n808_));
  AOI220     o786(.A0(ori_ori_n808_), .A1(ori_ori_n542_), .B0(ori_ori_n777_), .B1(ori_ori_n697_), .Y(ori_ori_n809_));
  NA3        o787(.A(ori_ori_n370_), .B(ori_ori_n242_), .C(ori_ori_n151_), .Y(ori_ori_n810_));
  NA2        o788(.A(ori_ori_n388_), .B(ori_ori_n70_), .Y(ori_ori_n811_));
  NA4        o789(.A(ori_ori_n811_), .B(ori_ori_n810_), .C(ori_ori_n809_), .D(ori_ori_n583_), .Y(ori_ori_n812_));
  AO210      o790(.A0(ori_ori_n501_), .A1(ori_ori_n46_), .B0(ori_ori_n88_), .Y(ori_ori_n813_));
  NA3        o791(.A(ori_ori_n813_), .B(ori_ori_n466_), .C(ori_ori_n220_), .Y(ori_ori_n814_));
  AOI210     o792(.A0(ori_ori_n436_), .A1(ori_ori_n434_), .B0(ori_ori_n541_), .Y(ori_ori_n815_));
  NO2        o793(.A(ori_ori_n591_), .B(ori_ori_n105_), .Y(ori_ori_n816_));
  OAI210     o794(.A0(ori_ori_n816_), .A1(ori_ori_n115_), .B0(ori_ori_n394_), .Y(ori_ori_n817_));
  INV        o795(.A(ori_ori_n565_), .Y(ori_ori_n818_));
  NA3        o796(.A(ori_ori_n818_), .B(ori_ori_n327_), .C(i_7_), .Y(ori_ori_n819_));
  NA4        o797(.A(ori_ori_n819_), .B(ori_ori_n817_), .C(ori_ori_n815_), .D(ori_ori_n814_), .Y(ori_ori_n820_));
  NO4        o798(.A(ori_ori_n820_), .B(ori_ori_n812_), .C(ori_ori_n807_), .D(ori_ori_n797_), .Y(ori_ori_n821_));
  NA4        o799(.A(ori_ori_n821_), .B(ori_ori_n783_), .C(ori_ori_n779_), .D(ori_ori_n378_), .Y(ori3));
  NA2        o800(.A(i_6_), .B(i_7_), .Y(ori_ori_n823_));
  NO2        o801(.A(ori_ori_n823_), .B(i_0_), .Y(ori_ori_n824_));
  NO2        o802(.A(i_11_), .B(ori_ori_n240_), .Y(ori_ori_n825_));
  OAI210     o803(.A0(ori_ori_n824_), .A1(ori_ori_n297_), .B0(ori_ori_n825_), .Y(ori_ori_n826_));
  NO2        o804(.A(ori_ori_n826_), .B(ori_ori_n195_), .Y(ori_ori_n827_));
  NO3        o805(.A(ori_ori_n441_), .B(ori_ori_n92_), .C(ori_ori_n44_), .Y(ori_ori_n828_));
  OA210      o806(.A0(ori_ori_n828_), .A1(ori_ori_n827_), .B0(ori_ori_n178_), .Y(ori_ori_n829_));
  NA3        o807(.A(ori_ori_n810_), .B(ori_ori_n583_), .C(ori_ori_n369_), .Y(ori_ori_n830_));
  NA2        o808(.A(ori_ori_n830_), .B(ori_ori_n40_), .Y(ori_ori_n831_));
  NOi21      o809(.An(ori_ori_n99_), .B(ori_ori_n742_), .Y(ori_ori_n832_));
  NO3        o810(.A(ori_ori_n608_), .B(ori_ori_n445_), .C(ori_ori_n135_), .Y(ori_ori_n833_));
  NA2        o811(.A(ori_ori_n397_), .B(ori_ori_n45_), .Y(ori_ori_n834_));
  AN2        o812(.A(ori_ori_n443_), .B(ori_ori_n55_), .Y(ori_ori_n835_));
  NO3        o813(.A(ori_ori_n835_), .B(ori_ori_n833_), .C(ori_ori_n832_), .Y(ori_ori_n836_));
  AOI210     o814(.A0(ori_ori_n836_), .A1(ori_ori_n831_), .B0(ori_ori_n48_), .Y(ori_ori_n837_));
  NO4        o815(.A(ori_ori_n374_), .B(ori_ori_n381_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n838_));
  NA2        o816(.A(ori_ori_n189_), .B(ori_ori_n549_), .Y(ori_ori_n839_));
  NOi21      o817(.An(ori_ori_n839_), .B(ori_ori_n838_), .Y(ori_ori_n840_));
  NA2        o818(.A(ori_ori_n689_), .B(ori_ori_n656_), .Y(ori_ori_n841_));
  NA2        o819(.A(ori_ori_n331_), .B(i_5_), .Y(ori_ori_n842_));
  OAI220     o820(.A0(ori_ori_n842_), .A1(ori_ori_n841_), .B0(ori_ori_n840_), .B1(ori_ori_n63_), .Y(ori_ori_n843_));
  NOi21      o821(.An(i_5_), .B(i_9_), .Y(ori_ori_n844_));
  NA2        o822(.A(ori_ori_n844_), .B(ori_ori_n432_), .Y(ori_ori_n845_));
  BUFFER     o823(.A(ori_ori_n272_), .Y(ori_ori_n846_));
  AOI210     o824(.A0(ori_ori_n846_), .A1(ori_ori_n463_), .B0(ori_ori_n670_), .Y(ori_ori_n847_));
  NO3        o825(.A(ori_ori_n400_), .B(ori_ori_n272_), .C(ori_ori_n73_), .Y(ori_ori_n848_));
  NO2        o826(.A(ori_ori_n179_), .B(ori_ori_n152_), .Y(ori_ori_n849_));
  AOI210     o827(.A0(ori_ori_n849_), .A1(ori_ori_n248_), .B0(ori_ori_n848_), .Y(ori_ori_n850_));
  OAI220     o828(.A0(ori_ori_n850_), .A1(ori_ori_n184_), .B0(ori_ori_n847_), .B1(ori_ori_n845_), .Y(ori_ori_n851_));
  NO4        o829(.A(ori_ori_n851_), .B(ori_ori_n843_), .C(ori_ori_n837_), .D(ori_ori_n829_), .Y(ori_ori_n852_));
  NA2        o830(.A(ori_ori_n189_), .B(ori_ori_n24_), .Y(ori_ori_n853_));
  NO2        o831(.A(ori_ori_n654_), .B(ori_ori_n572_), .Y(ori_ori_n854_));
  NO2        o832(.A(ori_ori_n854_), .B(ori_ori_n853_), .Y(ori_ori_n855_));
  INV        o833(.A(ori_ori_n855_), .Y(ori_ori_n856_));
  NA2        o834(.A(ori_ori_n550_), .B(i_0_), .Y(ori_ori_n857_));
  NO4        o835(.A(ori_ori_n564_), .B(ori_ori_n217_), .C(ori_ori_n404_), .D(ori_ori_n396_), .Y(ori_ori_n858_));
  NA2        o836(.A(ori_ori_n858_), .B(i_11_), .Y(ori_ori_n859_));
  AN2        o837(.A(ori_ori_n99_), .B(ori_ori_n247_), .Y(ori_ori_n860_));
  NA2        o838(.A(ori_ori_n729_), .B(ori_ori_n328_), .Y(ori_ori_n861_));
  AOI210     o839(.A0(ori_ori_n466_), .A1(ori_ori_n89_), .B0(ori_ori_n58_), .Y(ori_ori_n862_));
  OAI220     o840(.A0(ori_ori_n862_), .A1(ori_ori_n861_), .B0(ori_ori_n639_), .B1(ori_ori_n517_), .Y(ori_ori_n863_));
  NO2        o841(.A(ori_ori_n256_), .B(ori_ori_n158_), .Y(ori_ori_n864_));
  NA2        o842(.A(i_0_), .B(i_10_), .Y(ori_ori_n865_));
  INV        o843(.A(ori_ori_n520_), .Y(ori_ori_n866_));
  NO4        o844(.A(ori_ori_n118_), .B(ori_ori_n58_), .C(ori_ori_n649_), .D(i_5_), .Y(ori_ori_n867_));
  AO220      o845(.A0(ori_ori_n867_), .A1(ori_ori_n866_), .B0(ori_ori_n864_), .B1(i_6_), .Y(ori_ori_n868_));
  AOI220     o846(.A0(ori_ori_n331_), .A1(ori_ori_n101_), .B0(ori_ori_n189_), .B1(ori_ori_n84_), .Y(ori_ori_n869_));
  NA2        o847(.A(ori_ori_n544_), .B(i_4_), .Y(ori_ori_n870_));
  NA2        o848(.A(ori_ori_n191_), .B(ori_ori_n205_), .Y(ori_ori_n871_));
  OAI220     o849(.A0(ori_ori_n871_), .A1(ori_ori_n861_), .B0(ori_ori_n870_), .B1(ori_ori_n869_), .Y(ori_ori_n872_));
  NO4        o850(.A(ori_ori_n872_), .B(ori_ori_n868_), .C(ori_ori_n863_), .D(ori_ori_n860_), .Y(ori_ori_n873_));
  NA3        o851(.A(ori_ori_n873_), .B(ori_ori_n859_), .C(ori_ori_n856_), .Y(ori_ori_n874_));
  NA2        o852(.A(i_11_), .B(i_9_), .Y(ori_ori_n875_));
  NO2        o853(.A(ori_ori_n48_), .B(i_7_), .Y(ori_ori_n876_));
  NA2        o854(.A(ori_ori_n385_), .B(ori_ori_n182_), .Y(ori_ori_n877_));
  NA2        o855(.A(ori_ori_n877_), .B(ori_ori_n165_), .Y(ori_ori_n878_));
  NO2        o856(.A(ori_ori_n179_), .B(i_0_), .Y(ori_ori_n879_));
  INV        o857(.A(ori_ori_n879_), .Y(ori_ori_n880_));
  NA2        o858(.A(ori_ori_n462_), .B(ori_ori_n234_), .Y(ori_ori_n881_));
  INV        o859(.A(ori_ori_n393_), .Y(ori_ori_n882_));
  OAI220     o860(.A0(ori_ori_n882_), .A1(ori_ori_n845_), .B0(ori_ori_n881_), .B1(ori_ori_n880_), .Y(ori_ori_n883_));
  NO2        o861(.A(ori_ori_n883_), .B(ori_ori_n878_), .Y(ori_ori_n884_));
  NA2        o862(.A(ori_ori_n638_), .B(ori_ori_n125_), .Y(ori_ori_n885_));
  NO2        o863(.A(i_6_), .B(ori_ori_n885_), .Y(ori_ori_n886_));
  AOI210     o864(.A0(ori_ori_n435_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n887_));
  NA2        o865(.A(ori_ori_n176_), .B(ori_ori_n106_), .Y(ori_ori_n888_));
  NOi32      o866(.An(ori_ori_n887_), .Bn(ori_ori_n191_), .C(ori_ori_n888_), .Y(ori_ori_n889_));
  NA2        o867(.A(ori_ori_n584_), .B(ori_ori_n328_), .Y(ori_ori_n890_));
  NO2        o868(.A(ori_ori_n890_), .B(ori_ori_n834_), .Y(ori_ori_n891_));
  NO3        o869(.A(ori_ori_n891_), .B(ori_ori_n889_), .C(ori_ori_n886_), .Y(ori_ori_n892_));
  NOi21      o870(.An(i_7_), .B(i_5_), .Y(ori_ori_n893_));
  NOi31      o871(.An(ori_ori_n893_), .B(i_0_), .C(ori_ori_n707_), .Y(ori_ori_n894_));
  NA2        o872(.A(ori_ori_n892_), .B(ori_ori_n884_), .Y(ori_ori_n895_));
  AN2        o873(.A(ori_ori_n330_), .B(ori_ori_n328_), .Y(ori_ori_n896_));
  OA210      o874(.A0(ori_ori_n462_), .A1(ori_ori_n226_), .B0(ori_ori_n461_), .Y(ori_ori_n897_));
  NA3        o875(.A(ori_ori_n799_), .B(ori_ori_n380_), .C(ori_ori_n616_), .Y(ori_ori_n898_));
  NA2        o876(.A(ori_ori_n95_), .B(ori_ori_n44_), .Y(ori_ori_n899_));
  NO2        o877(.A(ori_ori_n75_), .B(ori_ori_n731_), .Y(ori_ori_n900_));
  AOI220     o878(.A0(ori_ori_n900_), .A1(ori_ori_n899_), .B0(ori_ori_n178_), .B1(ori_ori_n572_), .Y(ori_ori_n901_));
  AOI210     o879(.A0(ori_ori_n901_), .A1(ori_ori_n898_), .B0(ori_ori_n47_), .Y(ori_ori_n902_));
  NO3        o880(.A(ori_ori_n564_), .B(ori_ori_n354_), .C(ori_ori_n24_), .Y(ori_ori_n903_));
  INV        o881(.A(ori_ori_n903_), .Y(ori_ori_n904_));
  NO2        o882(.A(ori_ori_n578_), .B(ori_ori_n108_), .Y(ori_ori_n905_));
  NA2        o883(.A(ori_ori_n905_), .B(i_0_), .Y(ori_ori_n906_));
  OAI220     o884(.A0(ori_ori_n906_), .A1(ori_ori_n86_), .B0(ori_ori_n904_), .B1(ori_ori_n177_), .Y(ori_ori_n907_));
  NO3        o885(.A(ori_ori_n907_), .B(ori_ori_n902_), .C(ori_ori_n503_), .Y(ori_ori_n908_));
  INV        o886(.A(ori_ori_n908_), .Y(ori_ori_n909_));
  NO3        o887(.A(ori_ori_n909_), .B(ori_ori_n895_), .C(ori_ori_n874_), .Y(ori_ori_n910_));
  NO2        o888(.A(i_0_), .B(ori_ori_n707_), .Y(ori_ori_n911_));
  AOI210     o889(.A0(ori_ori_n780_), .A1(ori_ori_n668_), .B0(ori_ori_n888_), .Y(ori_ori_n912_));
  INV        o890(.A(ori_ori_n912_), .Y(ori_ori_n913_));
  NO2        o891(.A(ori_ori_n795_), .B(ori_ori_n391_), .Y(ori_ori_n914_));
  NA3        o892(.A(ori_ori_n824_), .B(i_2_), .C(ori_ori_n48_), .Y(ori_ori_n915_));
  NA2        o893(.A(ori_ori_n825_), .B(i_9_), .Y(ori_ori_n916_));
  AOI210     o894(.A0(ori_ori_n915_), .A1(ori_ori_n483_), .B0(ori_ori_n916_), .Y(ori_ori_n917_));
  OAI210     o895(.A0(ori_ori_n248_), .A1(i_9_), .B0(ori_ori_n233_), .Y(ori_ori_n918_));
  AOI210     o896(.A0(ori_ori_n918_), .A1(ori_ori_n857_), .B0(ori_ori_n158_), .Y(ori_ori_n919_));
  NO3        o897(.A(ori_ori_n919_), .B(ori_ori_n917_), .C(ori_ori_n914_), .Y(ori_ori_n920_));
  NA2        o898(.A(ori_ori_n920_), .B(ori_ori_n913_), .Y(ori_ori_n921_));
  NA2        o899(.A(ori_ori_n896_), .B(ori_ori_n370_), .Y(ori_ori_n922_));
  AOI210     o900(.A0(ori_ori_n304_), .A1(ori_ori_n167_), .B0(ori_ori_n922_), .Y(ori_ori_n923_));
  INV        o901(.A(ori_ori_n923_), .Y(ori_ori_n924_));
  NO3        o902(.A(ori_ori_n865_), .B(ori_ori_n844_), .C(ori_ori_n193_), .Y(ori_ori_n925_));
  AOI220     o903(.A0(ori_ori_n925_), .A1(i_11_), .B0(ori_ori_n545_), .B1(ori_ori_n75_), .Y(ori_ori_n926_));
  NO3        o904(.A(ori_ori_n212_), .B(ori_ori_n381_), .C(i_0_), .Y(ori_ori_n927_));
  OAI210     o905(.A0(ori_ori_n927_), .A1(ori_ori_n76_), .B0(i_13_), .Y(ori_ori_n928_));
  INV        o906(.A(ori_ori_n220_), .Y(ori_ori_n929_));
  OAI220     o907(.A0(ori_ori_n514_), .A1(ori_ori_n143_), .B0(ori_ori_n621_), .B1(ori_ori_n594_), .Y(ori_ori_n930_));
  NA3        o908(.A(ori_ori_n930_), .B(ori_ori_n389_), .C(ori_ori_n929_), .Y(ori_ori_n931_));
  NA4        o909(.A(ori_ori_n931_), .B(ori_ori_n928_), .C(ori_ori_n926_), .D(ori_ori_n924_), .Y(ori_ori_n932_));
  NO2        o910(.A(ori_ori_n246_), .B(ori_ori_n95_), .Y(ori_ori_n933_));
  AOI210     o911(.A0(ori_ori_n933_), .A1(ori_ori_n911_), .B0(ori_ori_n112_), .Y(ori_ori_n934_));
  AOI220     o912(.A0(ori_ori_n893_), .A1(ori_ori_n471_), .B0(ori_ori_n824_), .B1(ori_ori_n168_), .Y(ori_ori_n935_));
  NA2        o913(.A(ori_ori_n346_), .B(ori_ori_n180_), .Y(ori_ori_n936_));
  OA220      o914(.A0(ori_ori_n936_), .A1(ori_ori_n935_), .B0(ori_ori_n934_), .B1(i_5_), .Y(ori_ori_n937_));
  AOI210     o915(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n179_), .Y(ori_ori_n938_));
  NA2        o916(.A(ori_ori_n938_), .B(ori_ori_n897_), .Y(ori_ori_n939_));
  NA3        o917(.A(ori_ori_n592_), .B(ori_ori_n189_), .C(ori_ori_n84_), .Y(ori_ori_n940_));
  NA2        o918(.A(ori_ori_n940_), .B(ori_ori_n527_), .Y(ori_ori_n941_));
  NO3        o919(.A(ori_ori_n834_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n942_));
  NA2        o920(.A(ori_ori_n476_), .B(ori_ori_n469_), .Y(ori_ori_n943_));
  NO3        o921(.A(ori_ori_n943_), .B(ori_ori_n942_), .C(ori_ori_n941_), .Y(ori_ori_n944_));
  NA3        o922(.A(ori_ori_n384_), .B(ori_ori_n176_), .C(ori_ori_n175_), .Y(ori_ori_n945_));
  NA3        o923(.A(ori_ori_n876_), .B(ori_ori_n297_), .C(ori_ori_n233_), .Y(ori_ori_n946_));
  NA2        o924(.A(ori_ori_n946_), .B(ori_ori_n945_), .Y(ori_ori_n947_));
  NA3        o925(.A(ori_ori_n384_), .B(ori_ori_n332_), .C(ori_ori_n224_), .Y(ori_ori_n948_));
  INV        o926(.A(ori_ori_n948_), .Y(ori_ori_n949_));
  NO3        o927(.A(ori_ori_n875_), .B(ori_ori_n220_), .C(ori_ori_n193_), .Y(ori_ori_n950_));
  NO3        o928(.A(ori_ori_n950_), .B(ori_ori_n949_), .C(ori_ori_n947_), .Y(ori_ori_n951_));
  NA4        o929(.A(ori_ori_n951_), .B(ori_ori_n944_), .C(ori_ori_n939_), .D(ori_ori_n937_), .Y(ori_ori_n952_));
  NO2        o930(.A(ori_ori_n86_), .B(i_5_), .Y(ori_ori_n953_));
  NA3        o931(.A(ori_ori_n825_), .B(ori_ori_n113_), .C(ori_ori_n128_), .Y(ori_ori_n954_));
  INV        o932(.A(ori_ori_n954_), .Y(ori_ori_n955_));
  NA2        o933(.A(ori_ori_n955_), .B(ori_ori_n953_), .Y(ori_ori_n956_));
  NA3        o934(.A(ori_ori_n307_), .B(i_5_), .C(ori_ori_n195_), .Y(ori_ori_n957_));
  NAi31      o935(.An(ori_ori_n245_), .B(ori_ori_n957_), .C(ori_ori_n246_), .Y(ori_ori_n958_));
  NO4        o936(.A(ori_ori_n243_), .B(ori_ori_n212_), .C(i_0_), .D(i_12_), .Y(ori_ori_n959_));
  AOI220     o937(.A0(ori_ori_n959_), .A1(ori_ori_n958_), .B0(ori_ori_n776_), .B1(ori_ori_n180_), .Y(ori_ori_n960_));
  AN2        o938(.A(ori_ori_n865_), .B(ori_ori_n158_), .Y(ori_ori_n961_));
  NO4        o939(.A(ori_ori_n961_), .B(i_12_), .C(ori_ori_n625_), .D(ori_ori_n135_), .Y(ori_ori_n962_));
  NA2        o940(.A(ori_ori_n962_), .B(ori_ori_n220_), .Y(ori_ori_n963_));
  NA3        o941(.A(ori_ori_n101_), .B(ori_ori_n549_), .C(i_11_), .Y(ori_ori_n964_));
  NO2        o942(.A(ori_ori_n964_), .B(ori_ori_n160_), .Y(ori_ori_n965_));
  NA2        o943(.A(ori_ori_n893_), .B(ori_ori_n459_), .Y(ori_ori_n966_));
  NA2        o944(.A(ori_ori_n64_), .B(ori_ori_n104_), .Y(ori_ori_n967_));
  OAI220     o945(.A0(ori_ori_n967_), .A1(ori_ori_n957_), .B0(ori_ori_n966_), .B1(ori_ori_n657_), .Y(ori_ori_n968_));
  AOI210     o946(.A0(ori_ori_n968_), .A1(ori_ori_n879_), .B0(ori_ori_n965_), .Y(ori_ori_n969_));
  NA4        o947(.A(ori_ori_n969_), .B(ori_ori_n963_), .C(ori_ori_n960_), .D(ori_ori_n956_), .Y(ori_ori_n970_));
  NO4        o948(.A(ori_ori_n970_), .B(ori_ori_n952_), .C(ori_ori_n932_), .D(ori_ori_n921_), .Y(ori_ori_n971_));
  OAI210     o949(.A0(ori_ori_n798_), .A1(ori_ori_n792_), .B0(ori_ori_n37_), .Y(ori_ori_n972_));
  NA3        o950(.A(ori_ori_n887_), .B(ori_ori_n365_), .C(i_5_), .Y(ori_ori_n973_));
  NA3        o951(.A(ori_ori_n973_), .B(ori_ori_n972_), .C(ori_ori_n590_), .Y(ori_ori_n974_));
  NA2        o952(.A(ori_ori_n974_), .B(ori_ori_n210_), .Y(ori_ori_n975_));
  BUFFER     o953(.A(ori_ori_n366_), .Y(ori_ori_n976_));
  NA2        o954(.A(ori_ori_n190_), .B(ori_ori_n191_), .Y(ori_ori_n977_));
  AO210      o955(.A0(ori_ori_n976_), .A1(ori_ori_n33_), .B0(ori_ori_n977_), .Y(ori_ori_n978_));
  NAi31      o956(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n979_));
  AOI210     o957(.A0(ori_ori_n121_), .A1(ori_ori_n70_), .B0(ori_ori_n979_), .Y(ori_ori_n980_));
  NO2        o958(.A(ori_ori_n980_), .B(ori_ori_n622_), .Y(ori_ori_n981_));
  NA2        o959(.A(ori_ori_n981_), .B(ori_ori_n978_), .Y(ori_ori_n982_));
  NO2        o960(.A(ori_ori_n453_), .B(ori_ori_n272_), .Y(ori_ori_n983_));
  NO2        o961(.A(ori_ori_n983_), .B(ori_ori_n858_), .Y(ori_ori_n984_));
  OAI210     o962(.A0(ori_ori_n964_), .A1(ori_ori_n152_), .B0(ori_ori_n984_), .Y(ori_ori_n985_));
  AOI210     o963(.A0(ori_ori_n982_), .A1(ori_ori_n48_), .B0(ori_ori_n985_), .Y(ori_ori_n986_));
  AOI210     o964(.A0(ori_ori_n986_), .A1(ori_ori_n975_), .B0(ori_ori_n73_), .Y(ori_ori_n987_));
  INV        o965(.A(ori_ori_n377_), .Y(ori_ori_n988_));
  NO2        o966(.A(ori_ori_n988_), .B(ori_ori_n737_), .Y(ori_ori_n989_));
  OAI210     o967(.A0(ori_ori_n80_), .A1(ori_ori_n54_), .B0(ori_ori_n111_), .Y(ori_ori_n990_));
  NA2        o968(.A(ori_ori_n990_), .B(ori_ori_n76_), .Y(ori_ori_n991_));
  AOI210     o969(.A0(ori_ori_n938_), .A1(ori_ori_n876_), .B0(ori_ori_n894_), .Y(ori_ori_n992_));
  AOI210     o970(.A0(ori_ori_n992_), .A1(ori_ori_n991_), .B0(ori_ori_n660_), .Y(ori_ori_n993_));
  NA2        o971(.A(ori_ori_n266_), .B(ori_ori_n57_), .Y(ori_ori_n994_));
  AOI220     o972(.A0(ori_ori_n994_), .A1(ori_ori_n76_), .B0(ori_ori_n343_), .B1(ori_ori_n258_), .Y(ori_ori_n995_));
  NO2        o973(.A(ori_ori_n995_), .B(ori_ori_n240_), .Y(ori_ori_n996_));
  NO2        o974(.A(ori_ori_n996_), .B(ori_ori_n993_), .Y(ori_ori_n997_));
  OAI210     o975(.A0(ori_ori_n274_), .A1(ori_ori_n163_), .B0(ori_ori_n89_), .Y(ori_ori_n998_));
  NO2        o976(.A(ori_ori_n998_), .B(i_11_), .Y(ori_ori_n999_));
  NA2        o977(.A(ori_ori_n585_), .B(ori_ori_n217_), .Y(ori_ori_n1000_));
  OAI210     o978(.A0(ori_ori_n1000_), .A1(ori_ori_n887_), .B0(ori_ori_n210_), .Y(ori_ori_n1001_));
  NA2        o979(.A(ori_ori_n169_), .B(i_5_), .Y(ori_ori_n1002_));
  NO2        o980(.A(ori_ori_n1001_), .B(ori_ori_n1002_), .Y(ori_ori_n1003_));
  INV        o981(.A(ori_ori_n360_), .Y(ori_ori_n1004_));
  NO2        o982(.A(ori_ori_n1004_), .B(ori_ori_n41_), .Y(ori_ori_n1005_));
  NO3        o983(.A(ori_ori_n1005_), .B(ori_ori_n1003_), .C(ori_ori_n999_), .Y(ori_ori_n1006_));
  OAI210     o984(.A0(ori_ori_n997_), .A1(i_4_), .B0(ori_ori_n1006_), .Y(ori_ori_n1007_));
  NO3        o985(.A(ori_ori_n1007_), .B(ori_ori_n989_), .C(ori_ori_n987_), .Y(ori_ori_n1008_));
  NA4        o986(.A(ori_ori_n1008_), .B(ori_ori_n971_), .C(ori_ori_n910_), .D(ori_ori_n852_), .Y(ori4));
  INV        o987(.A(ori_ori_n681_), .Y(ori_ori_n1012_));
  INV        o988(.A(ori_ori_n527_), .Y(ori_ori_n1013_));
  INV        o989(.A(ori_ori_n695_), .Y(ori_ori_n1014_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m0033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m0034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m0036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m0037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m0038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m0039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m0040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m0041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m0042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m0043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m0044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m0045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m0046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m0047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m0049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m0050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m0051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m0052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m0053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m0054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m0055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m0057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m0059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m0060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m0062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m0063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m0064(.A(i_6_), .Y(mai_mai_n87_));
  OR4        m0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n88_));
  INV        m0066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m0067(.A(i_2_), .B(i_7_), .Y(mai_mai_n90_));
  NO2        m0068(.A(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  OAI210     m0069(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NAi21      m0070(.An(i_6_), .B(i_10_), .Y(mai_mai_n93_));
  NA2        m0071(.A(i_6_), .B(i_9_), .Y(mai_mai_n94_));
  AOI210     m0072(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n64_), .Y(mai_mai_n95_));
  NA2        m0073(.A(i_2_), .B(i_6_), .Y(mai_mai_n96_));
  NO3        m0074(.A(mai_mai_n96_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n97_));
  NO2        m0075(.A(mai_mai_n97_), .B(mai_mai_n95_), .Y(mai_mai_n98_));
  AOI210     m0076(.A0(mai_mai_n98_), .A1(mai_mai_n92_), .B0(mai_mai_n81_), .Y(mai_mai_n99_));
  AN3        m0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n100_));
  NAi21      m0078(.An(i_6_), .B(i_11_), .Y(mai_mai_n101_));
  NO2        m0079(.A(i_5_), .B(i_8_), .Y(mai_mai_n102_));
  NOi21      m0080(.An(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  AOI220     m0081(.A0(mai_mai_n103_), .A1(mai_mai_n63_), .B0(mai_mai_n100_), .B1(mai_mai_n32_), .Y(mai_mai_n104_));
  INV        m0082(.A(i_7_), .Y(mai_mai_n105_));
  NA2        m0083(.A(mai_mai_n47_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  NO2        m0084(.A(i_0_), .B(i_5_), .Y(mai_mai_n107_));
  NO2        m0085(.A(mai_mai_n107_), .B(mai_mai_n87_), .Y(mai_mai_n108_));
  NA2        m0086(.A(i_12_), .B(i_3_), .Y(mai_mai_n109_));
  INV        m0087(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NA3        m0088(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n106_), .Y(mai_mai_n111_));
  NAi21      m0089(.An(i_7_), .B(i_11_), .Y(mai_mai_n112_));
  NO3        m0090(.A(mai_mai_n112_), .B(mai_mai_n93_), .C(mai_mai_n54_), .Y(mai_mai_n113_));
  AN2        m0091(.A(i_2_), .B(i_10_), .Y(mai_mai_n114_));
  NO2        m0092(.A(mai_mai_n114_), .B(i_7_), .Y(mai_mai_n115_));
  OR2        m0093(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n116_));
  NO2        m0094(.A(i_8_), .B(mai_mai_n105_), .Y(mai_mai_n117_));
  NO3        m0095(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(mai_mai_n115_), .Y(mai_mai_n118_));
  NA2        m0096(.A(i_12_), .B(i_7_), .Y(mai_mai_n119_));
  NO2        m0097(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n120_));
  NA2        m0098(.A(i_11_), .B(i_12_), .Y(mai_mai_n121_));
  INV        m0099(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  NO2        m0100(.A(mai_mai_n122_), .B(mai_mai_n118_), .Y(mai_mai_n123_));
  NAi41      m0101(.An(mai_mai_n113_), .B(mai_mai_n123_), .C(mai_mai_n111_), .D(mai_mai_n104_), .Y(mai_mai_n124_));
  NOi21      m0102(.An(i_1_), .B(i_5_), .Y(mai_mai_n125_));
  NA2        m0103(.A(mai_mai_n125_), .B(i_11_), .Y(mai_mai_n126_));
  NA2        m0104(.A(mai_mai_n105_), .B(mai_mai_n37_), .Y(mai_mai_n127_));
  NA2        m0105(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n128_));
  NA2        m0106(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n129_));
  NO2        m0107(.A(mai_mai_n129_), .B(mai_mai_n47_), .Y(mai_mai_n130_));
  NA2        m0108(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n131_));
  NAi21      m0109(.An(i_3_), .B(i_8_), .Y(mai_mai_n132_));
  NA2        m0110(.A(mai_mai_n132_), .B(mai_mai_n63_), .Y(mai_mai_n133_));
  NOi31      m0111(.An(mai_mai_n133_), .B(mai_mai_n131_), .C(mai_mai_n130_), .Y(mai_mai_n134_));
  NO2        m0112(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n135_));
  NO2        m0113(.A(i_6_), .B(i_5_), .Y(mai_mai_n136_));
  NA2        m0114(.A(mai_mai_n136_), .B(i_3_), .Y(mai_mai_n137_));
  AO210      m0115(.A0(mai_mai_n137_), .A1(mai_mai_n48_), .B0(mai_mai_n135_), .Y(mai_mai_n138_));
  OAI220     m0116(.A0(mai_mai_n138_), .A1(mai_mai_n112_), .B0(mai_mai_n134_), .B1(mai_mai_n126_), .Y(mai_mai_n139_));
  NO3        m0117(.A(mai_mai_n139_), .B(mai_mai_n124_), .C(mai_mai_n99_), .Y(mai_mai_n140_));
  NA3        m0118(.A(mai_mai_n140_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m0119(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n142_));
  NA2        m0120(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n143_));
  NA2        m0121(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NA4        m0122(.A(mai_mai_n144_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0123(.A(i_8_), .B(i_7_), .Y(mai_mai_n146_));
  NA2        m0124(.A(mai_mai_n146_), .B(i_6_), .Y(mai_mai_n147_));
  NO2        m0125(.A(i_12_), .B(i_13_), .Y(mai_mai_n148_));
  NAi21      m0126(.An(i_5_), .B(i_11_), .Y(mai_mai_n149_));
  NOi21      m0127(.An(mai_mai_n148_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  NO2        m0128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NA2        m0129(.A(i_2_), .B(i_3_), .Y(mai_mai_n152_));
  NO2        m0130(.A(mai_mai_n152_), .B(i_4_), .Y(mai_mai_n153_));
  AN2        m0131(.A(mai_mai_n148_), .B(mai_mai_n84_), .Y(mai_mai_n154_));
  NA2        m0132(.A(i_1_), .B(i_5_), .Y(mai_mai_n155_));
  NO2        m0133(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n156_));
  OR2        m0134(.A(i_0_), .B(i_1_), .Y(mai_mai_n157_));
  NO3        m0135(.A(mai_mai_n157_), .B(mai_mai_n81_), .C(i_13_), .Y(mai_mai_n158_));
  NAi32      m0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n159_));
  NAi21      m0137(.An(mai_mai_n159_), .B(mai_mai_n158_), .Y(mai_mai_n160_));
  NOi21      m0138(.An(i_4_), .B(i_10_), .Y(mai_mai_n161_));
  NA2        m0139(.A(mai_mai_n161_), .B(mai_mai_n40_), .Y(mai_mai_n162_));
  NO2        m0140(.A(i_3_), .B(i_5_), .Y(mai_mai_n163_));
  NO3        m0141(.A(mai_mai_n74_), .B(i_2_), .C(i_1_), .Y(mai_mai_n164_));
  NA3        m0142(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n165_));
  NA2        m0143(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n166_));
  NOi21      m0144(.An(i_4_), .B(i_9_), .Y(mai_mai_n167_));
  NOi21      m0145(.An(i_11_), .B(i_13_), .Y(mai_mai_n168_));
  NA2        m0146(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  OR2        m0147(.A(mai_mai_n169_), .B(mai_mai_n166_), .Y(mai_mai_n170_));
  NO2        m0148(.A(i_4_), .B(i_5_), .Y(mai_mai_n171_));
  NAi21      m0149(.An(i_12_), .B(i_11_), .Y(mai_mai_n172_));
  NO2        m0150(.A(mai_mai_n172_), .B(i_13_), .Y(mai_mai_n173_));
  NA3        m0151(.A(mai_mai_n173_), .B(mai_mai_n171_), .C(mai_mai_n84_), .Y(mai_mai_n174_));
  AOI210     m0152(.A0(mai_mai_n174_), .A1(mai_mai_n170_), .B0(mai_mai_n165_), .Y(mai_mai_n175_));
  NO2        m0153(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n176_));
  NA2        m0154(.A(mai_mai_n176_), .B(mai_mai_n47_), .Y(mai_mai_n177_));
  NAi31      m0155(.An(i_4_), .B(mai_mai_n154_), .C(i_11_), .Y(mai_mai_n178_));
  NA2        m0156(.A(i_3_), .B(i_5_), .Y(mai_mai_n179_));
  OR2        m0157(.A(mai_mai_n179_), .B(mai_mai_n169_), .Y(mai_mai_n180_));
  AOI210     m0158(.A0(mai_mai_n180_), .A1(mai_mai_n178_), .B0(mai_mai_n177_), .Y(mai_mai_n181_));
  NO2        m0159(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n182_));
  NO2        m0160(.A(i_13_), .B(i_10_), .Y(mai_mai_n183_));
  NA3        m0161(.A(mai_mai_n183_), .B(mai_mai_n182_), .C(mai_mai_n45_), .Y(mai_mai_n184_));
  NO2        m0162(.A(i_2_), .B(i_1_), .Y(mai_mai_n185_));
  NA2        m0163(.A(mai_mai_n185_), .B(i_3_), .Y(mai_mai_n186_));
  NAi21      m0164(.An(i_4_), .B(i_12_), .Y(mai_mai_n187_));
  NO4        m0165(.A(mai_mai_n187_), .B(mai_mai_n186_), .C(mai_mai_n184_), .D(mai_mai_n25_), .Y(mai_mai_n188_));
  NO3        m0166(.A(mai_mai_n188_), .B(mai_mai_n181_), .C(mai_mai_n175_), .Y(mai_mai_n189_));
  INV        m0167(.A(i_8_), .Y(mai_mai_n190_));
  NO2        m0168(.A(mai_mai_n190_), .B(i_7_), .Y(mai_mai_n191_));
  NA2        m0169(.A(mai_mai_n191_), .B(i_6_), .Y(mai_mai_n192_));
  NO3        m0170(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n193_));
  NA2        m0171(.A(mai_mai_n193_), .B(mai_mai_n117_), .Y(mai_mai_n194_));
  NO3        m0172(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n195_));
  NO3        m0173(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n196_));
  NA2        m0174(.A(i_12_), .B(mai_mai_n196_), .Y(mai_mai_n197_));
  NO2        m0175(.A(mai_mai_n197_), .B(mai_mai_n194_), .Y(mai_mai_n198_));
  NO2        m0176(.A(i_3_), .B(i_8_), .Y(mai_mai_n199_));
  NO3        m0177(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n200_));
  NO2        m0178(.A(mai_mai_n107_), .B(mai_mai_n59_), .Y(mai_mai_n201_));
  NO2        m0179(.A(i_13_), .B(i_9_), .Y(mai_mai_n202_));
  NA3        m0180(.A(mai_mai_n202_), .B(i_6_), .C(mai_mai_n190_), .Y(mai_mai_n203_));
  NAi21      m0181(.An(i_12_), .B(i_3_), .Y(mai_mai_n204_));
  OR2        m0182(.A(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  NO2        m0183(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n206_));
  NO3        m0184(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n207_));
  NA3        m0185(.A(mai_mai_n207_), .B(mai_mai_n206_), .C(i_10_), .Y(mai_mai_n208_));
  NO2        m0186(.A(mai_mai_n208_), .B(mai_mai_n205_), .Y(mai_mai_n209_));
  NO2        m0187(.A(mai_mai_n209_), .B(mai_mai_n198_), .Y(mai_mai_n210_));
  OAI220     m0188(.A0(mai_mai_n210_), .A1(i_4_), .B0(mai_mai_n192_), .B1(mai_mai_n189_), .Y(mai_mai_n211_));
  NAi21      m0189(.An(i_12_), .B(i_7_), .Y(mai_mai_n212_));
  NA3        m0190(.A(i_13_), .B(mai_mai_n190_), .C(i_10_), .Y(mai_mai_n213_));
  NO2        m0191(.A(mai_mai_n213_), .B(mai_mai_n212_), .Y(mai_mai_n214_));
  NA2        m0192(.A(i_0_), .B(i_5_), .Y(mai_mai_n215_));
  NA2        m0193(.A(mai_mai_n215_), .B(mai_mai_n108_), .Y(mai_mai_n216_));
  OAI220     m0194(.A0(mai_mai_n216_), .A1(mai_mai_n186_), .B0(mai_mai_n177_), .B1(mai_mai_n137_), .Y(mai_mai_n217_));
  NAi31      m0195(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n218_));
  NO2        m0196(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n219_));
  NO2        m0197(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n220_));
  NO2        m0198(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n221_));
  INV        m0199(.A(i_13_), .Y(mai_mai_n222_));
  NO2        m0200(.A(i_12_), .B(mai_mai_n222_), .Y(mai_mai_n223_));
  NA2        m0201(.A(mai_mai_n217_), .B(mai_mai_n214_), .Y(mai_mai_n224_));
  NO2        m0202(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n225_));
  NO2        m0203(.A(mai_mai_n179_), .B(i_4_), .Y(mai_mai_n226_));
  NA2        m0204(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n227_));
  OR2        m0205(.A(i_8_), .B(i_7_), .Y(mai_mai_n228_));
  NO2        m0206(.A(mai_mai_n228_), .B(mai_mai_n87_), .Y(mai_mai_n229_));
  NO2        m0207(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n230_));
  NA2        m0208(.A(mai_mai_n230_), .B(mai_mai_n229_), .Y(mai_mai_n231_));
  INV        m0209(.A(i_12_), .Y(mai_mai_n232_));
  NO2        m0210(.A(mai_mai_n45_), .B(mai_mai_n232_), .Y(mai_mai_n233_));
  NO3        m0211(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n234_));
  NA2        m0212(.A(i_2_), .B(i_1_), .Y(mai_mai_n235_));
  NO2        m0213(.A(mai_mai_n231_), .B(mai_mai_n227_), .Y(mai_mai_n236_));
  NO3        m0214(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n237_));
  NAi21      m0215(.An(i_4_), .B(i_3_), .Y(mai_mai_n238_));
  NO2        m0216(.A(mai_mai_n238_), .B(mai_mai_n76_), .Y(mai_mai_n239_));
  NO2        m0217(.A(i_0_), .B(i_6_), .Y(mai_mai_n240_));
  NOi41      m0218(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n241_));
  NA2        m0219(.A(mai_mai_n241_), .B(mai_mai_n240_), .Y(mai_mai_n242_));
  NO2        m0220(.A(mai_mai_n235_), .B(mai_mai_n179_), .Y(mai_mai_n243_));
  NAi21      m0221(.An(mai_mai_n242_), .B(mai_mai_n243_), .Y(mai_mai_n244_));
  INV        m0222(.A(mai_mai_n244_), .Y(mai_mai_n245_));
  AOI220     m0223(.A0(mai_mai_n245_), .A1(mai_mai_n40_), .B0(mai_mai_n236_), .B1(mai_mai_n202_), .Y(mai_mai_n246_));
  NO2        m0224(.A(i_11_), .B(mai_mai_n222_), .Y(mai_mai_n247_));
  NOi21      m0225(.An(i_1_), .B(i_6_), .Y(mai_mai_n248_));
  NAi21      m0226(.An(i_3_), .B(i_7_), .Y(mai_mai_n249_));
  NA2        m0227(.A(mai_mai_n232_), .B(i_9_), .Y(mai_mai_n250_));
  OR4        m0228(.A(mai_mai_n250_), .B(mai_mai_n249_), .C(mai_mai_n248_), .D(mai_mai_n182_), .Y(mai_mai_n251_));
  NO2        m0229(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n252_));
  NO2        m0230(.A(i_12_), .B(i_3_), .Y(mai_mai_n253_));
  NA2        m0231(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n254_));
  NA2        m0232(.A(i_3_), .B(i_9_), .Y(mai_mai_n255_));
  NAi21      m0233(.An(i_7_), .B(i_10_), .Y(mai_mai_n256_));
  NO2        m0234(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n257_));
  NA3        m0235(.A(mai_mai_n257_), .B(mai_mai_n254_), .C(mai_mai_n65_), .Y(mai_mai_n258_));
  NA2        m0236(.A(mai_mai_n258_), .B(mai_mai_n251_), .Y(mai_mai_n259_));
  NA3        m0237(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n260_));
  INV        m0238(.A(mai_mai_n147_), .Y(mai_mai_n261_));
  NA2        m0239(.A(mai_mai_n232_), .B(i_13_), .Y(mai_mai_n262_));
  NO2        m0240(.A(mai_mai_n262_), .B(mai_mai_n76_), .Y(mai_mai_n263_));
  AOI220     m0241(.A0(mai_mai_n263_), .A1(mai_mai_n261_), .B0(mai_mai_n259_), .B1(mai_mai_n247_), .Y(mai_mai_n264_));
  NO2        m0242(.A(mai_mai_n228_), .B(mai_mai_n37_), .Y(mai_mai_n265_));
  NA2        m0243(.A(i_12_), .B(i_6_), .Y(mai_mai_n266_));
  OR2        m0244(.A(i_13_), .B(i_9_), .Y(mai_mai_n267_));
  NO3        m0245(.A(mai_mai_n267_), .B(mai_mai_n266_), .C(mai_mai_n49_), .Y(mai_mai_n268_));
  NO2        m0246(.A(mai_mai_n238_), .B(i_2_), .Y(mai_mai_n269_));
  NA3        m0247(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n45_), .Y(mai_mai_n270_));
  NA2        m0248(.A(mai_mai_n247_), .B(i_9_), .Y(mai_mai_n271_));
  NA2        m0249(.A(mai_mai_n254_), .B(mai_mai_n65_), .Y(mai_mai_n272_));
  OAI210     m0250(.A0(mai_mai_n272_), .A1(mai_mai_n271_), .B0(mai_mai_n270_), .Y(mai_mai_n273_));
  NA2        m0251(.A(mai_mai_n156_), .B(mai_mai_n64_), .Y(mai_mai_n274_));
  NO3        m0252(.A(i_11_), .B(mai_mai_n222_), .C(mai_mai_n25_), .Y(mai_mai_n275_));
  NO2        m0253(.A(mai_mai_n249_), .B(i_8_), .Y(mai_mai_n276_));
  NO2        m0254(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n277_));
  NA3        m0255(.A(mai_mai_n277_), .B(mai_mai_n276_), .C(mai_mai_n275_), .Y(mai_mai_n278_));
  NO3        m0256(.A(mai_mai_n26_), .B(mai_mai_n87_), .C(i_5_), .Y(mai_mai_n279_));
  NA3        m0257(.A(mai_mai_n279_), .B(mai_mai_n265_), .C(mai_mai_n223_), .Y(mai_mai_n280_));
  AOI210     m0258(.A0(mai_mai_n280_), .A1(mai_mai_n278_), .B0(mai_mai_n274_), .Y(mai_mai_n281_));
  AOI210     m0259(.A0(mai_mai_n273_), .A1(mai_mai_n265_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  NA4        m0260(.A(mai_mai_n282_), .B(mai_mai_n264_), .C(mai_mai_n246_), .D(mai_mai_n224_), .Y(mai_mai_n283_));
  NO3        m0261(.A(i_12_), .B(mai_mai_n222_), .C(mai_mai_n37_), .Y(mai_mai_n284_));
  INV        m0262(.A(mai_mai_n284_), .Y(mai_mai_n285_));
  NA2        m0263(.A(i_8_), .B(mai_mai_n105_), .Y(mai_mai_n286_));
  NOi21      m0264(.An(mai_mai_n163_), .B(mai_mai_n87_), .Y(mai_mai_n287_));
  NO3        m0265(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n288_));
  AOI220     m0266(.A0(mai_mai_n288_), .A1(mai_mai_n193_), .B0(mai_mai_n287_), .B1(mai_mai_n230_), .Y(mai_mai_n289_));
  NO2        m0267(.A(mai_mai_n289_), .B(mai_mai_n286_), .Y(mai_mai_n290_));
  NO3        m0268(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n291_));
  NO2        m0269(.A(mai_mai_n235_), .B(i_0_), .Y(mai_mai_n292_));
  AOI220     m0270(.A0(mai_mai_n292_), .A1(mai_mai_n191_), .B0(mai_mai_n291_), .B1(mai_mai_n146_), .Y(mai_mai_n293_));
  NA2        m0271(.A(mai_mai_n277_), .B(mai_mai_n26_), .Y(mai_mai_n294_));
  NO2        m0272(.A(mai_mai_n294_), .B(mai_mai_n293_), .Y(mai_mai_n295_));
  NA2        m0273(.A(i_0_), .B(i_1_), .Y(mai_mai_n296_));
  NO2        m0274(.A(mai_mai_n296_), .B(i_2_), .Y(mai_mai_n297_));
  NO2        m0275(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n298_));
  NA3        m0276(.A(mai_mai_n298_), .B(mai_mai_n297_), .C(mai_mai_n163_), .Y(mai_mai_n299_));
  INV        m0277(.A(mai_mai_n299_), .Y(mai_mai_n300_));
  NO3        m0278(.A(mai_mai_n300_), .B(mai_mai_n295_), .C(mai_mai_n290_), .Y(mai_mai_n301_));
  NO2        m0279(.A(i_3_), .B(i_10_), .Y(mai_mai_n302_));
  NA3        m0280(.A(mai_mai_n302_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n303_));
  NO2        m0281(.A(i_2_), .B(mai_mai_n105_), .Y(mai_mai_n304_));
  NA2        m0282(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n305_));
  NO2        m0283(.A(mai_mai_n305_), .B(i_8_), .Y(mai_mai_n306_));
  NOi21      m0284(.An(mai_mai_n215_), .B(mai_mai_n107_), .Y(mai_mai_n307_));
  NA3        m0285(.A(mai_mai_n307_), .B(mai_mai_n306_), .C(mai_mai_n304_), .Y(mai_mai_n308_));
  AN2        m0286(.A(i_3_), .B(i_10_), .Y(mai_mai_n309_));
  NO2        m0287(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n310_));
  NO2        m0288(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n311_));
  OR2        m0289(.A(mai_mai_n308_), .B(mai_mai_n303_), .Y(mai_mai_n312_));
  OAI220     m0290(.A0(mai_mai_n312_), .A1(i_6_), .B0(mai_mai_n301_), .B1(mai_mai_n285_), .Y(mai_mai_n313_));
  NO3        m0291(.A(mai_mai_n313_), .B(mai_mai_n283_), .C(mai_mai_n211_), .Y(mai_mai_n314_));
  NO3        m0292(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n315_));
  NO2        m0293(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n316_));
  NA2        m0294(.A(mai_mai_n292_), .B(mai_mai_n316_), .Y(mai_mai_n317_));
  NO3        m0295(.A(i_6_), .B(mai_mai_n190_), .C(i_7_), .Y(mai_mai_n318_));
  NA2        m0296(.A(mai_mai_n318_), .B(mai_mai_n195_), .Y(mai_mai_n319_));
  AOI210     m0297(.A0(mai_mai_n319_), .A1(mai_mai_n317_), .B0(mai_mai_n166_), .Y(mai_mai_n320_));
  NO2        m0298(.A(i_2_), .B(i_3_), .Y(mai_mai_n321_));
  OR2        m0299(.A(i_0_), .B(i_5_), .Y(mai_mai_n322_));
  NA2        m0300(.A(mai_mai_n215_), .B(mai_mai_n322_), .Y(mai_mai_n323_));
  NA4        m0301(.A(mai_mai_n323_), .B(mai_mai_n229_), .C(mai_mai_n321_), .D(i_1_), .Y(mai_mai_n324_));
  NA3        m0302(.A(mai_mai_n292_), .B(mai_mai_n287_), .C(mai_mai_n117_), .Y(mai_mai_n325_));
  NAi21      m0303(.An(i_8_), .B(i_7_), .Y(mai_mai_n326_));
  NO2        m0304(.A(mai_mai_n326_), .B(i_6_), .Y(mai_mai_n327_));
  NO2        m0305(.A(mai_mai_n157_), .B(mai_mai_n47_), .Y(mai_mai_n328_));
  NA2        m0306(.A(mai_mai_n325_), .B(mai_mai_n324_), .Y(mai_mai_n329_));
  OAI210     m0307(.A0(mai_mai_n329_), .A1(mai_mai_n320_), .B0(i_4_), .Y(mai_mai_n330_));
  NO2        m0308(.A(i_12_), .B(i_10_), .Y(mai_mai_n331_));
  NOi21      m0309(.An(i_5_), .B(i_0_), .Y(mai_mai_n332_));
  NO3        m0310(.A(mai_mai_n305_), .B(mai_mai_n332_), .C(mai_mai_n132_), .Y(mai_mai_n333_));
  NA4        m0311(.A(mai_mai_n85_), .B(mai_mai_n36_), .C(mai_mai_n87_), .D(i_8_), .Y(mai_mai_n334_));
  NA2        m0312(.A(mai_mai_n333_), .B(mai_mai_n331_), .Y(mai_mai_n335_));
  NO2        m0313(.A(i_6_), .B(i_8_), .Y(mai_mai_n336_));
  NOi21      m0314(.An(i_0_), .B(i_2_), .Y(mai_mai_n337_));
  AN2        m0315(.A(mai_mai_n337_), .B(mai_mai_n336_), .Y(mai_mai_n338_));
  NO2        m0316(.A(i_1_), .B(i_7_), .Y(mai_mai_n339_));
  AO220      m0317(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n327_), .B1(mai_mai_n230_), .Y(mai_mai_n340_));
  NA3        m0318(.A(mai_mai_n340_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n341_));
  NA3        m0319(.A(mai_mai_n341_), .B(mai_mai_n335_), .C(mai_mai_n330_), .Y(mai_mai_n342_));
  NO3        m0320(.A(mai_mai_n228_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n343_));
  NO3        m0321(.A(mai_mai_n326_), .B(i_2_), .C(i_1_), .Y(mai_mai_n344_));
  OAI210     m0322(.A0(mai_mai_n344_), .A1(mai_mai_n343_), .B0(i_6_), .Y(mai_mai_n345_));
  NO2        m0323(.A(mai_mai_n345_), .B(mai_mai_n323_), .Y(mai_mai_n346_));
  NOi21      m0324(.An(mai_mai_n155_), .B(mai_mai_n108_), .Y(mai_mai_n347_));
  NO2        m0325(.A(mai_mai_n347_), .B(mai_mai_n128_), .Y(mai_mai_n348_));
  OAI210     m0326(.A0(mai_mai_n348_), .A1(mai_mai_n346_), .B0(i_3_), .Y(mai_mai_n349_));
  INV        m0327(.A(mai_mai_n85_), .Y(mai_mai_n350_));
  NO2        m0328(.A(mai_mai_n296_), .B(mai_mai_n82_), .Y(mai_mai_n351_));
  NO2        m0329(.A(mai_mai_n96_), .B(mai_mai_n190_), .Y(mai_mai_n352_));
  NA3        m0330(.A(mai_mai_n307_), .B(mai_mai_n352_), .C(mai_mai_n64_), .Y(mai_mai_n353_));
  NO2        m0331(.A(mai_mai_n353_), .B(mai_mai_n350_), .Y(mai_mai_n354_));
  NO2        m0332(.A(mai_mai_n190_), .B(i_9_), .Y(mai_mai_n355_));
  NA2        m0333(.A(mai_mai_n355_), .B(mai_mai_n201_), .Y(mai_mai_n356_));
  NO2        m0334(.A(mai_mai_n356_), .B(mai_mai_n47_), .Y(mai_mai_n357_));
  NO3        m0335(.A(mai_mai_n357_), .B(mai_mai_n354_), .C(mai_mai_n295_), .Y(mai_mai_n358_));
  AOI210     m0336(.A0(mai_mai_n358_), .A1(mai_mai_n349_), .B0(mai_mai_n162_), .Y(mai_mai_n359_));
  AOI210     m0337(.A0(mai_mai_n342_), .A1(mai_mai_n315_), .B0(mai_mai_n359_), .Y(mai_mai_n360_));
  NOi32      m0338(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n361_));
  INV        m0339(.A(mai_mai_n361_), .Y(mai_mai_n362_));
  NAi21      m0340(.An(i_1_), .B(i_5_), .Y(mai_mai_n363_));
  NAi41      m0341(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n364_));
  OAI220     m0342(.A0(mai_mai_n364_), .A1(mai_mai_n363_), .B0(mai_mai_n218_), .B1(mai_mai_n159_), .Y(mai_mai_n365_));
  AOI210     m0343(.A0(mai_mai_n364_), .A1(mai_mai_n159_), .B0(mai_mai_n157_), .Y(mai_mai_n366_));
  NOi32      m0344(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n367_));
  NAi21      m0345(.An(i_6_), .B(i_1_), .Y(mai_mai_n368_));
  NA3        m0346(.A(mai_mai_n368_), .B(mai_mai_n367_), .C(mai_mai_n47_), .Y(mai_mai_n369_));
  NO2        m0347(.A(mai_mai_n369_), .B(i_0_), .Y(mai_mai_n370_));
  OR3        m0348(.A(mai_mai_n370_), .B(mai_mai_n366_), .C(mai_mai_n365_), .Y(mai_mai_n371_));
  NO2        m0349(.A(i_1_), .B(mai_mai_n105_), .Y(mai_mai_n372_));
  NAi21      m0350(.An(i_3_), .B(i_4_), .Y(mai_mai_n373_));
  NO2        m0351(.A(mai_mai_n373_), .B(i_9_), .Y(mai_mai_n374_));
  AN2        m0352(.A(i_6_), .B(i_7_), .Y(mai_mai_n375_));
  OAI210     m0353(.A0(mai_mai_n375_), .A1(mai_mai_n372_), .B0(mai_mai_n374_), .Y(mai_mai_n376_));
  NA2        m0354(.A(i_2_), .B(i_7_), .Y(mai_mai_n377_));
  NO2        m0355(.A(mai_mai_n373_), .B(i_10_), .Y(mai_mai_n378_));
  NA3        m0356(.A(mai_mai_n378_), .B(mai_mai_n377_), .C(mai_mai_n240_), .Y(mai_mai_n379_));
  AOI210     m0357(.A0(mai_mai_n379_), .A1(mai_mai_n376_), .B0(mai_mai_n182_), .Y(mai_mai_n380_));
  AOI210     m0358(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n381_));
  OAI210     m0359(.A0(mai_mai_n381_), .A1(mai_mai_n185_), .B0(mai_mai_n378_), .Y(mai_mai_n382_));
  AOI220     m0360(.A0(mai_mai_n378_), .A1(mai_mai_n339_), .B0(mai_mai_n234_), .B1(mai_mai_n185_), .Y(mai_mai_n383_));
  AOI210     m0361(.A0(mai_mai_n383_), .A1(mai_mai_n382_), .B0(i_5_), .Y(mai_mai_n384_));
  NO3        m0362(.A(mai_mai_n384_), .B(mai_mai_n380_), .C(mai_mai_n371_), .Y(mai_mai_n385_));
  NO2        m0363(.A(mai_mai_n385_), .B(mai_mai_n362_), .Y(mai_mai_n386_));
  NO2        m0364(.A(mai_mai_n60_), .B(mai_mai_n25_), .Y(mai_mai_n387_));
  AN2        m0365(.A(i_12_), .B(i_5_), .Y(mai_mai_n388_));
  NO2        m0366(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n389_));
  NA2        m0367(.A(mai_mai_n389_), .B(mai_mai_n388_), .Y(mai_mai_n390_));
  NO2        m0368(.A(i_11_), .B(i_6_), .Y(mai_mai_n391_));
  NA3        m0369(.A(mai_mai_n391_), .B(mai_mai_n328_), .C(mai_mai_n222_), .Y(mai_mai_n392_));
  NO2        m0370(.A(mai_mai_n392_), .B(mai_mai_n390_), .Y(mai_mai_n393_));
  NO2        m0371(.A(mai_mai_n238_), .B(i_5_), .Y(mai_mai_n394_));
  NO2        m0372(.A(i_5_), .B(i_10_), .Y(mai_mai_n395_));
  AOI220     m0373(.A0(mai_mai_n395_), .A1(mai_mai_n269_), .B0(mai_mai_n394_), .B1(mai_mai_n195_), .Y(mai_mai_n396_));
  NA2        m0374(.A(mai_mai_n148_), .B(mai_mai_n46_), .Y(mai_mai_n397_));
  NO2        m0375(.A(mai_mai_n397_), .B(mai_mai_n396_), .Y(mai_mai_n398_));
  OAI210     m0376(.A0(mai_mai_n398_), .A1(mai_mai_n393_), .B0(mai_mai_n387_), .Y(mai_mai_n399_));
  NO2        m0377(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n400_));
  NA2        m0378(.A(mai_mai_n393_), .B(mai_mai_n400_), .Y(mai_mai_n401_));
  NO3        m0379(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n402_));
  NO2        m0380(.A(i_11_), .B(i_12_), .Y(mai_mai_n403_));
  NA2        m0381(.A(mai_mai_n395_), .B(mai_mai_n232_), .Y(mai_mai_n404_));
  NA3        m0382(.A(mai_mai_n117_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n405_));
  OAI220     m0383(.A0(mai_mai_n405_), .A1(mai_mai_n218_), .B0(mai_mai_n404_), .B1(mai_mai_n334_), .Y(mai_mai_n406_));
  NAi21      m0384(.An(i_13_), .B(i_0_), .Y(mai_mai_n407_));
  NO2        m0385(.A(mai_mai_n407_), .B(mai_mai_n235_), .Y(mai_mai_n408_));
  NA2        m0386(.A(mai_mai_n406_), .B(mai_mai_n408_), .Y(mai_mai_n409_));
  NA3        m0387(.A(mai_mai_n409_), .B(mai_mai_n401_), .C(mai_mai_n399_), .Y(mai_mai_n410_));
  NA2        m0388(.A(mai_mai_n45_), .B(mai_mai_n222_), .Y(mai_mai_n411_));
  NO3        m0389(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n412_));
  NO2        m0390(.A(i_0_), .B(i_11_), .Y(mai_mai_n413_));
  AN2        m0391(.A(i_1_), .B(i_6_), .Y(mai_mai_n414_));
  NOi21      m0392(.An(i_2_), .B(i_12_), .Y(mai_mai_n415_));
  NAi21      m0393(.An(i_9_), .B(i_4_), .Y(mai_mai_n416_));
  OR2        m0394(.A(i_13_), .B(i_10_), .Y(mai_mai_n417_));
  NO3        m0395(.A(mai_mai_n417_), .B(mai_mai_n121_), .C(mai_mai_n416_), .Y(mai_mai_n418_));
  NO2        m0396(.A(mai_mai_n169_), .B(mai_mai_n127_), .Y(mai_mai_n419_));
  NO2        m0397(.A(mai_mai_n105_), .B(mai_mai_n25_), .Y(mai_mai_n420_));
  NA2        m0398(.A(mai_mai_n284_), .B(mai_mai_n420_), .Y(mai_mai_n421_));
  NO2        m0399(.A(mai_mai_n421_), .B(mai_mai_n347_), .Y(mai_mai_n422_));
  INV        m0400(.A(mai_mai_n422_), .Y(mai_mai_n423_));
  NO2        m0401(.A(mai_mai_n423_), .B(mai_mai_n26_), .Y(mai_mai_n424_));
  NA2        m0402(.A(mai_mai_n325_), .B(mai_mai_n324_), .Y(mai_mai_n425_));
  NO2        m0403(.A(mai_mai_n179_), .B(mai_mai_n87_), .Y(mai_mai_n426_));
  AOI220     m0404(.A0(mai_mai_n426_), .A1(mai_mai_n297_), .B0(mai_mai_n279_), .B1(mai_mai_n207_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n427_), .B(mai_mai_n286_), .Y(mai_mai_n428_));
  NO2        m0406(.A(mai_mai_n428_), .B(mai_mai_n425_), .Y(mai_mai_n429_));
  NA2        m0407(.A(mai_mai_n190_), .B(i_10_), .Y(mai_mai_n430_));
  NA3        m0408(.A(mai_mai_n254_), .B(mai_mai_n65_), .C(i_2_), .Y(mai_mai_n431_));
  NA2        m0409(.A(mai_mai_n298_), .B(mai_mai_n230_), .Y(mai_mai_n432_));
  OAI220     m0410(.A0(mai_mai_n432_), .A1(mai_mai_n179_), .B0(mai_mai_n431_), .B1(mai_mai_n430_), .Y(mai_mai_n433_));
  NO2        m0411(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n434_));
  NA3        m0412(.A(mai_mai_n339_), .B(mai_mai_n338_), .C(mai_mai_n434_), .Y(mai_mai_n435_));
  NA2        m0413(.A(mai_mai_n318_), .B(mai_mai_n323_), .Y(mai_mai_n436_));
  OAI210     m0414(.A0(mai_mai_n436_), .A1(mai_mai_n186_), .B0(mai_mai_n435_), .Y(mai_mai_n437_));
  NO2        m0415(.A(mai_mai_n437_), .B(mai_mai_n433_), .Y(mai_mai_n438_));
  AOI210     m0416(.A0(mai_mai_n438_), .A1(mai_mai_n429_), .B0(mai_mai_n271_), .Y(mai_mai_n439_));
  NO4        m0417(.A(mai_mai_n439_), .B(mai_mai_n424_), .C(mai_mai_n410_), .D(mai_mai_n386_), .Y(mai_mai_n440_));
  NO2        m0418(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n441_));
  NO2        m0419(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n442_));
  NA3        m0420(.A(mai_mai_n442_), .B(mai_mai_n441_), .C(i_2_), .Y(mai_mai_n443_));
  NO2        m0421(.A(i_10_), .B(i_9_), .Y(mai_mai_n444_));
  NAi21      m0422(.An(i_12_), .B(i_8_), .Y(mai_mai_n445_));
  NO2        m0423(.A(mai_mai_n445_), .B(i_3_), .Y(mai_mai_n446_));
  NA2        m0424(.A(mai_mai_n446_), .B(mai_mai_n444_), .Y(mai_mai_n447_));
  NO2        m0425(.A(mai_mai_n47_), .B(i_4_), .Y(mai_mai_n448_));
  NO2        m0426(.A(mai_mai_n447_), .B(mai_mai_n443_), .Y(mai_mai_n449_));
  NA2        m0427(.A(mai_mai_n311_), .B(i_0_), .Y(mai_mai_n450_));
  NO3        m0428(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n451_));
  NA2        m0429(.A(mai_mai_n266_), .B(mai_mai_n101_), .Y(mai_mai_n452_));
  NA2        m0430(.A(mai_mai_n452_), .B(mai_mai_n451_), .Y(mai_mai_n453_));
  NA2        m0431(.A(i_8_), .B(i_9_), .Y(mai_mai_n454_));
  AOI210     m0432(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n455_));
  OR2        m0433(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n456_));
  NA2        m0434(.A(mai_mai_n284_), .B(mai_mai_n201_), .Y(mai_mai_n457_));
  OAI220     m0435(.A0(mai_mai_n457_), .A1(mai_mai_n456_), .B0(mai_mai_n453_), .B1(mai_mai_n450_), .Y(mai_mai_n458_));
  NA2        m0436(.A(mai_mai_n247_), .B(mai_mai_n310_), .Y(mai_mai_n459_));
  NO3        m0437(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n460_));
  INV        m0438(.A(mai_mai_n460_), .Y(mai_mai_n461_));
  NA3        m0439(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n462_));
  NA4        m0440(.A(mai_mai_n149_), .B(mai_mai_n120_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n463_));
  OAI220     m0441(.A0(mai_mai_n463_), .A1(mai_mai_n462_), .B0(mai_mai_n461_), .B1(mai_mai_n459_), .Y(mai_mai_n464_));
  NO3        m0442(.A(mai_mai_n464_), .B(mai_mai_n458_), .C(mai_mai_n449_), .Y(mai_mai_n465_));
  NA2        m0443(.A(mai_mai_n297_), .B(mai_mai_n112_), .Y(mai_mai_n466_));
  OR2        m0444(.A(mai_mai_n466_), .B(mai_mai_n203_), .Y(mai_mai_n467_));
  OA210      m0445(.A0(mai_mai_n356_), .A1(mai_mai_n105_), .B0(mai_mai_n299_), .Y(mai_mai_n468_));
  OA220      m0446(.A0(mai_mai_n468_), .A1(mai_mai_n162_), .B0(mai_mai_n467_), .B1(mai_mai_n227_), .Y(mai_mai_n469_));
  NA2        m0447(.A(mai_mai_n100_), .B(i_13_), .Y(mai_mai_n470_));
  NO2        m0448(.A(i_2_), .B(i_13_), .Y(mai_mai_n471_));
  NO3        m0449(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n472_));
  NO2        m0450(.A(i_6_), .B(i_7_), .Y(mai_mai_n473_));
  NA2        m0451(.A(mai_mai_n473_), .B(mai_mai_n472_), .Y(mai_mai_n474_));
  NO2        m0452(.A(i_11_), .B(i_1_), .Y(mai_mai_n475_));
  NO2        m0453(.A(mai_mai_n74_), .B(i_3_), .Y(mai_mai_n476_));
  OR2        m0454(.A(i_11_), .B(i_8_), .Y(mai_mai_n477_));
  NOi21      m0455(.An(i_2_), .B(i_7_), .Y(mai_mai_n478_));
  NAi31      m0456(.An(mai_mai_n477_), .B(mai_mai_n478_), .C(mai_mai_n476_), .Y(mai_mai_n479_));
  NO2        m0457(.A(mai_mai_n417_), .B(i_6_), .Y(mai_mai_n480_));
  NA3        m0458(.A(mai_mai_n480_), .B(mai_mai_n441_), .C(mai_mai_n76_), .Y(mai_mai_n481_));
  NO2        m0459(.A(mai_mai_n481_), .B(mai_mai_n479_), .Y(mai_mai_n482_));
  NO2        m0460(.A(i_6_), .B(i_10_), .Y(mai_mai_n483_));
  NA3        m0461(.A(mai_mai_n241_), .B(mai_mai_n168_), .C(mai_mai_n136_), .Y(mai_mai_n484_));
  NA2        m0462(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n485_));
  NO2        m0463(.A(mai_mai_n157_), .B(i_3_), .Y(mai_mai_n486_));
  NAi31      m0464(.An(mai_mai_n485_), .B(mai_mai_n486_), .C(mai_mai_n223_), .Y(mai_mai_n487_));
  NA3        m0465(.A(mai_mai_n400_), .B(mai_mai_n176_), .C(mai_mai_n153_), .Y(mai_mai_n488_));
  NA3        m0466(.A(mai_mai_n488_), .B(mai_mai_n487_), .C(mai_mai_n484_), .Y(mai_mai_n489_));
  NO2        m0467(.A(mai_mai_n489_), .B(mai_mai_n482_), .Y(mai_mai_n490_));
  NA2        m0468(.A(mai_mai_n451_), .B(mai_mai_n388_), .Y(mai_mai_n491_));
  NA2        m0469(.A(mai_mai_n460_), .B(mai_mai_n395_), .Y(mai_mai_n492_));
  NAi21      m0470(.An(mai_mai_n213_), .B(mai_mai_n403_), .Y(mai_mai_n493_));
  NO2        m0471(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n494_));
  NO2        m0472(.A(i_0_), .B(mai_mai_n87_), .Y(mai_mai_n495_));
  NA3        m0473(.A(mai_mai_n495_), .B(mai_mai_n494_), .C(mai_mai_n146_), .Y(mai_mai_n496_));
  OR3        m0474(.A(mai_mai_n305_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n497_));
  NO2        m0475(.A(mai_mai_n497_), .B(mai_mai_n496_), .Y(mai_mai_n498_));
  NA2        m0476(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n499_));
  NA2        m0477(.A(mai_mai_n315_), .B(mai_mai_n234_), .Y(mai_mai_n500_));
  OAI220     m0478(.A0(mai_mai_n500_), .A1(mai_mai_n431_), .B0(mai_mai_n499_), .B1(mai_mai_n470_), .Y(mai_mai_n501_));
  NA4        m0479(.A(mai_mai_n309_), .B(mai_mai_n221_), .C(mai_mai_n74_), .D(mai_mai_n232_), .Y(mai_mai_n502_));
  NO2        m0480(.A(mai_mai_n502_), .B(mai_mai_n474_), .Y(mai_mai_n503_));
  NO3        m0481(.A(mai_mai_n503_), .B(mai_mai_n501_), .C(mai_mai_n498_), .Y(mai_mai_n504_));
  NA4        m0482(.A(mai_mai_n504_), .B(mai_mai_n490_), .C(mai_mai_n469_), .D(mai_mai_n465_), .Y(mai_mai_n505_));
  NA3        m0483(.A(mai_mai_n309_), .B(mai_mai_n173_), .C(mai_mai_n171_), .Y(mai_mai_n506_));
  OAI210     m0484(.A0(mai_mai_n303_), .A1(i_4_), .B0(mai_mai_n506_), .Y(mai_mai_n507_));
  AN2        m0485(.A(mai_mai_n288_), .B(mai_mai_n229_), .Y(mai_mai_n508_));
  NA2        m0486(.A(mai_mai_n508_), .B(mai_mai_n507_), .Y(mai_mai_n509_));
  NA4        m0487(.A(mai_mai_n442_), .B(mai_mai_n441_), .C(mai_mai_n199_), .D(i_2_), .Y(mai_mai_n510_));
  INV        m0488(.A(mai_mai_n510_), .Y(mai_mai_n511_));
  NA2        m0489(.A(mai_mai_n388_), .B(mai_mai_n222_), .Y(mai_mai_n512_));
  NA2        m0490(.A(mai_mai_n361_), .B(mai_mai_n74_), .Y(mai_mai_n513_));
  NA2        m0491(.A(mai_mai_n375_), .B(mai_mai_n367_), .Y(mai_mai_n514_));
  OR2        m0492(.A(mai_mai_n512_), .B(mai_mai_n514_), .Y(mai_mai_n515_));
  NO2        m0493(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n516_));
  NAi41      m0494(.An(mai_mai_n513_), .B(mai_mai_n483_), .C(mai_mai_n516_), .D(mai_mai_n47_), .Y(mai_mai_n517_));
  AOI210     m0495(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n418_), .Y(mai_mai_n518_));
  NA3        m0496(.A(mai_mai_n518_), .B(mai_mai_n517_), .C(mai_mai_n515_), .Y(mai_mai_n519_));
  AOI210     m0497(.A0(mai_mai_n511_), .A1(mai_mai_n200_), .B0(mai_mai_n519_), .Y(mai_mai_n520_));
  INV        m0498(.A(mai_mai_n138_), .Y(mai_mai_n521_));
  NA2        m0499(.A(mai_mai_n521_), .B(mai_mai_n419_), .Y(mai_mai_n522_));
  NA3        m0500(.A(mai_mai_n522_), .B(mai_mai_n520_), .C(mai_mai_n509_), .Y(mai_mai_n523_));
  NA2        m0501(.A(mai_mai_n394_), .B(mai_mai_n297_), .Y(mai_mai_n524_));
  OAI210     m0502(.A0(mai_mai_n390_), .A1(mai_mai_n165_), .B0(mai_mai_n524_), .Y(mai_mai_n525_));
  NO2        m0503(.A(i_12_), .B(mai_mai_n190_), .Y(mai_mai_n526_));
  NA2        m0504(.A(mai_mai_n526_), .B(mai_mai_n222_), .Y(mai_mai_n527_));
  NA3        m0505(.A(mai_mai_n483_), .B(mai_mai_n171_), .C(mai_mai_n27_), .Y(mai_mai_n528_));
  NO2        m0506(.A(mai_mai_n528_), .B(mai_mai_n527_), .Y(mai_mai_n529_));
  NOi31      m0507(.An(mai_mai_n318_), .B(mai_mai_n417_), .C(mai_mai_n38_), .Y(mai_mai_n530_));
  OAI210     m0508(.A0(mai_mai_n530_), .A1(mai_mai_n529_), .B0(mai_mai_n525_), .Y(mai_mai_n531_));
  NO2        m0509(.A(i_8_), .B(i_7_), .Y(mai_mai_n532_));
  OAI210     m0510(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n533_));
  NA2        m0511(.A(mai_mai_n533_), .B(mai_mai_n221_), .Y(mai_mai_n534_));
  NO2        m0512(.A(mai_mai_n534_), .B(mai_mai_n238_), .Y(mai_mai_n535_));
  NA2        m0513(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n536_));
  NO2        m0514(.A(mai_mai_n536_), .B(i_6_), .Y(mai_mai_n537_));
  NA3        m0515(.A(mai_mai_n537_), .B(mai_mai_n535_), .C(mai_mai_n532_), .Y(mai_mai_n538_));
  AOI220     m0516(.A0(mai_mai_n426_), .A1(mai_mai_n328_), .B0(mai_mai_n243_), .B1(mai_mai_n240_), .Y(mai_mai_n539_));
  OAI220     m0517(.A0(mai_mai_n539_), .A1(mai_mai_n262_), .B0(mai_mai_n470_), .B1(mai_mai_n137_), .Y(mai_mai_n540_));
  NA2        m0518(.A(mai_mai_n540_), .B(mai_mai_n265_), .Y(mai_mai_n541_));
  NO2        m0519(.A(mai_mai_n219_), .B(mai_mai_n45_), .Y(mai_mai_n542_));
  NO2        m0520(.A(mai_mai_n157_), .B(i_5_), .Y(mai_mai_n543_));
  NA3        m0521(.A(mai_mai_n543_), .B(mai_mai_n411_), .C(mai_mai_n321_), .Y(mai_mai_n544_));
  NO2        m0522(.A(mai_mai_n544_), .B(mai_mai_n542_), .Y(mai_mai_n545_));
  NA2        m0523(.A(mai_mai_n545_), .B(mai_mai_n460_), .Y(mai_mai_n546_));
  NA4        m0524(.A(mai_mai_n546_), .B(mai_mai_n541_), .C(mai_mai_n538_), .D(mai_mai_n531_), .Y(mai_mai_n547_));
  NA3        m0525(.A(mai_mai_n215_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n548_));
  NA2        m0526(.A(mai_mai_n284_), .B(mai_mai_n85_), .Y(mai_mai_n549_));
  NO2        m0527(.A(mai_mai_n548_), .B(mai_mai_n549_), .Y(mai_mai_n550_));
  NA2        m0528(.A(mai_mai_n298_), .B(mai_mai_n288_), .Y(mai_mai_n551_));
  NO2        m0529(.A(mai_mai_n551_), .B(mai_mai_n170_), .Y(mai_mai_n552_));
  NA2        m0530(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n553_));
  NA2        m0531(.A(mai_mai_n444_), .B(mai_mai_n219_), .Y(mai_mai_n554_));
  NO2        m0532(.A(mai_mai_n553_), .B(mai_mai_n554_), .Y(mai_mai_n555_));
  AOI210     m0533(.A0(mai_mai_n368_), .A1(mai_mai_n47_), .B0(mai_mai_n372_), .Y(mai_mai_n556_));
  NA2        m0534(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n557_));
  NA3        m0535(.A(mai_mai_n526_), .B(mai_mai_n275_), .C(mai_mai_n557_), .Y(mai_mai_n558_));
  NO2        m0536(.A(mai_mai_n556_), .B(mai_mai_n558_), .Y(mai_mai_n559_));
  NO4        m0537(.A(mai_mai_n559_), .B(mai_mai_n555_), .C(mai_mai_n552_), .D(mai_mai_n550_), .Y(mai_mai_n560_));
  NO4        m0538(.A(mai_mai_n248_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n561_));
  NO3        m0539(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n562_));
  NO2        m0540(.A(mai_mai_n228_), .B(mai_mai_n36_), .Y(mai_mai_n563_));
  AN2        m0541(.A(mai_mai_n563_), .B(mai_mai_n562_), .Y(mai_mai_n564_));
  OA210      m0542(.A0(mai_mai_n564_), .A1(mai_mai_n561_), .B0(mai_mai_n361_), .Y(mai_mai_n565_));
  NO2        m0543(.A(mai_mai_n417_), .B(i_1_), .Y(mai_mai_n566_));
  NOi31      m0544(.An(mai_mai_n566_), .B(mai_mai_n452_), .C(mai_mai_n74_), .Y(mai_mai_n567_));
  INV        m0545(.A(mai_mai_n565_), .Y(mai_mai_n568_));
  NOi21      m0546(.An(i_10_), .B(i_6_), .Y(mai_mai_n569_));
  NO2        m0547(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n570_));
  AOI220     m0548(.A0(mai_mai_n284_), .A1(mai_mai_n570_), .B0(mai_mai_n275_), .B1(mai_mai_n569_), .Y(mai_mai_n571_));
  NO2        m0549(.A(mai_mai_n571_), .B(mai_mai_n450_), .Y(mai_mai_n572_));
  NO2        m0550(.A(mai_mai_n119_), .B(mai_mai_n23_), .Y(mai_mai_n573_));
  NA2        m0551(.A(mai_mai_n318_), .B(mai_mai_n164_), .Y(mai_mai_n574_));
  AOI220     m0552(.A0(mai_mai_n574_), .A1(mai_mai_n432_), .B0(mai_mai_n180_), .B1(mai_mai_n178_), .Y(mai_mai_n575_));
  NO2        m0553(.A(mai_mai_n195_), .B(mai_mai_n37_), .Y(mai_mai_n576_));
  NOi31      m0554(.An(mai_mai_n150_), .B(mai_mai_n576_), .C(mai_mai_n334_), .Y(mai_mai_n577_));
  NO3        m0555(.A(mai_mai_n577_), .B(mai_mai_n575_), .C(mai_mai_n572_), .Y(mai_mai_n578_));
  NO2        m0556(.A(mai_mai_n513_), .B(mai_mai_n383_), .Y(mai_mai_n579_));
  INV        m0557(.A(mai_mai_n321_), .Y(mai_mai_n580_));
  NO2        m0558(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n581_));
  NA2        m0559(.A(mai_mai_n171_), .B(i_0_), .Y(mai_mai_n582_));
  NO3        m0560(.A(mai_mai_n582_), .B(mai_mai_n345_), .C(mai_mai_n303_), .Y(mai_mai_n583_));
  OR2        m0561(.A(i_2_), .B(i_5_), .Y(mai_mai_n584_));
  OR2        m0562(.A(mai_mai_n584_), .B(mai_mai_n414_), .Y(mai_mai_n585_));
  AOI210     m0563(.A0(mai_mai_n377_), .A1(mai_mai_n240_), .B0(mai_mai_n195_), .Y(mai_mai_n586_));
  AOI210     m0564(.A0(mai_mai_n586_), .A1(mai_mai_n585_), .B0(mai_mai_n493_), .Y(mai_mai_n587_));
  NO3        m0565(.A(mai_mai_n587_), .B(mai_mai_n583_), .C(mai_mai_n579_), .Y(mai_mai_n588_));
  NA4        m0566(.A(mai_mai_n588_), .B(mai_mai_n578_), .C(mai_mai_n568_), .D(mai_mai_n560_), .Y(mai_mai_n589_));
  NO4        m0567(.A(mai_mai_n589_), .B(mai_mai_n547_), .C(mai_mai_n523_), .D(mai_mai_n505_), .Y(mai_mai_n590_));
  NA4        m0568(.A(mai_mai_n590_), .B(mai_mai_n440_), .C(mai_mai_n360_), .D(mai_mai_n314_), .Y(mai7));
  NO2        m0569(.A(mai_mai_n96_), .B(mai_mai_n55_), .Y(mai_mai_n592_));
  NO2        m0570(.A(mai_mai_n112_), .B(mai_mai_n93_), .Y(mai_mai_n593_));
  NA2        m0571(.A(mai_mai_n389_), .B(mai_mai_n593_), .Y(mai_mai_n594_));
  NA2        m0572(.A(mai_mai_n483_), .B(mai_mai_n85_), .Y(mai_mai_n595_));
  NA2        m0573(.A(i_11_), .B(mai_mai_n190_), .Y(mai_mai_n596_));
  NA2        m0574(.A(mai_mai_n148_), .B(mai_mai_n596_), .Y(mai_mai_n597_));
  OAI210     m0575(.A0(mai_mai_n597_), .A1(mai_mai_n595_), .B0(mai_mai_n594_), .Y(mai_mai_n598_));
  NA3        m0576(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n599_));
  NO2        m0577(.A(mai_mai_n232_), .B(i_4_), .Y(mai_mai_n600_));
  NA2        m0578(.A(mai_mai_n600_), .B(i_8_), .Y(mai_mai_n601_));
  NO2        m0579(.A(mai_mai_n109_), .B(mai_mai_n599_), .Y(mai_mai_n602_));
  NA2        m0580(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n603_));
  OAI210     m0581(.A0(mai_mai_n90_), .A1(mai_mai_n199_), .B0(mai_mai_n200_), .Y(mai_mai_n604_));
  NO2        m0582(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n605_));
  NA2        m0583(.A(i_4_), .B(i_8_), .Y(mai_mai_n606_));
  AOI210     m0584(.A0(mai_mai_n606_), .A1(mai_mai_n309_), .B0(mai_mai_n605_), .Y(mai_mai_n607_));
  OAI220     m0585(.A0(mai_mai_n607_), .A1(mai_mai_n603_), .B0(mai_mai_n604_), .B1(i_13_), .Y(mai_mai_n608_));
  NO4        m0586(.A(mai_mai_n608_), .B(mai_mai_n602_), .C(mai_mai_n598_), .D(mai_mai_n592_), .Y(mai_mai_n609_));
  AOI210     m0587(.A0(mai_mai_n132_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n610_));
  AOI210     m0588(.A0(mai_mai_n610_), .A1(mai_mai_n232_), .B0(mai_mai_n161_), .Y(mai_mai_n611_));
  OR2        m0589(.A(i_6_), .B(i_10_), .Y(mai_mai_n612_));
  NO2        m0590(.A(mai_mai_n612_), .B(mai_mai_n23_), .Y(mai_mai_n613_));
  OR3        m0591(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n614_));
  NO3        m0592(.A(mai_mai_n614_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n615_));
  INV        m0593(.A(mai_mai_n196_), .Y(mai_mai_n616_));
  NO2        m0594(.A(mai_mai_n615_), .B(mai_mai_n613_), .Y(mai_mai_n617_));
  OA220      m0595(.A0(mai_mai_n617_), .A1(mai_mai_n580_), .B0(mai_mai_n611_), .B1(mai_mai_n267_), .Y(mai_mai_n618_));
  AOI210     m0596(.A0(mai_mai_n618_), .A1(mai_mai_n609_), .B0(mai_mai_n64_), .Y(mai_mai_n619_));
  NOi21      m0597(.An(i_11_), .B(i_7_), .Y(mai_mai_n620_));
  AO210      m0598(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n621_));
  NO2        m0599(.A(mai_mai_n621_), .B(mai_mai_n620_), .Y(mai_mai_n622_));
  NA2        m0600(.A(mai_mai_n622_), .B(mai_mai_n202_), .Y(mai_mai_n623_));
  NA3        m0601(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n624_));
  NAi31      m0602(.An(mai_mai_n624_), .B(mai_mai_n212_), .C(i_11_), .Y(mai_mai_n625_));
  AOI210     m0603(.A0(mai_mai_n625_), .A1(mai_mai_n623_), .B0(mai_mai_n64_), .Y(mai_mai_n626_));
  NA2        m0604(.A(mai_mai_n89_), .B(mai_mai_n64_), .Y(mai_mai_n627_));
  AO210      m0605(.A0(mai_mai_n627_), .A1(mai_mai_n383_), .B0(mai_mai_n41_), .Y(mai_mai_n628_));
  NO3        m0606(.A(mai_mai_n256_), .B(mai_mai_n204_), .C(mai_mai_n596_), .Y(mai_mai_n629_));
  OAI210     m0607(.A0(mai_mai_n629_), .A1(mai_mai_n223_), .B0(mai_mai_n64_), .Y(mai_mai_n630_));
  NA2        m0608(.A(mai_mai_n415_), .B(mai_mai_n31_), .Y(mai_mai_n631_));
  OR2        m0609(.A(mai_mai_n204_), .B(mai_mai_n112_), .Y(mai_mai_n632_));
  NA2        m0610(.A(mai_mai_n632_), .B(mai_mai_n631_), .Y(mai_mai_n633_));
  NO2        m0611(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n634_));
  NO2        m0612(.A(mai_mai_n634_), .B(i_4_), .Y(mai_mai_n635_));
  NA2        m0613(.A(mai_mai_n635_), .B(mai_mai_n633_), .Y(mai_mai_n636_));
  NO2        m0614(.A(i_1_), .B(i_12_), .Y(mai_mai_n637_));
  NA3        m0615(.A(mai_mai_n637_), .B(mai_mai_n114_), .C(mai_mai_n24_), .Y(mai_mai_n638_));
  BUFFER     m0616(.A(mai_mai_n638_), .Y(mai_mai_n639_));
  NA4        m0617(.A(mai_mai_n639_), .B(mai_mai_n636_), .C(mai_mai_n630_), .D(mai_mai_n628_), .Y(mai_mai_n640_));
  OAI210     m0618(.A0(mai_mai_n640_), .A1(mai_mai_n626_), .B0(i_6_), .Y(mai_mai_n641_));
  NO2        m0619(.A(mai_mai_n624_), .B(mai_mai_n112_), .Y(mai_mai_n642_));
  NA2        m0620(.A(mai_mai_n642_), .B(mai_mai_n581_), .Y(mai_mai_n643_));
  NO2        m0621(.A(i_6_), .B(i_11_), .Y(mai_mai_n644_));
  NA2        m0622(.A(mai_mai_n643_), .B(mai_mai_n453_), .Y(mai_mai_n645_));
  NO3        m0623(.A(mai_mai_n612_), .B(mai_mai_n228_), .C(mai_mai_n23_), .Y(mai_mai_n646_));
  AOI210     m0624(.A0(i_1_), .A1(mai_mai_n257_), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  NO2        m0625(.A(mai_mai_n647_), .B(mai_mai_n45_), .Y(mai_mai_n648_));
  INV        m0626(.A(i_2_), .Y(mai_mai_n649_));
  NA2        m0627(.A(mai_mai_n142_), .B(i_9_), .Y(mai_mai_n650_));
  NA3        m0628(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n651_));
  NO2        m0629(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n652_));
  NO2        m0630(.A(mai_mai_n650_), .B(mai_mai_n649_), .Y(mai_mai_n653_));
  NA3        m0631(.A(mai_mai_n634_), .B(mai_mai_n321_), .C(i_6_), .Y(mai_mai_n654_));
  NO2        m0632(.A(mai_mai_n654_), .B(mai_mai_n23_), .Y(mai_mai_n655_));
  AOI210     m0633(.A0(mai_mai_n475_), .A1(mai_mai_n420_), .B0(mai_mai_n237_), .Y(mai_mai_n656_));
  NO2        m0634(.A(mai_mai_n656_), .B(mai_mai_n603_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n652_), .B(mai_mai_n266_), .Y(mai_mai_n658_));
  NO2        m0636(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n659_));
  NA2        m0637(.A(mai_mai_n659_), .B(mai_mai_n24_), .Y(mai_mai_n660_));
  NO2        m0638(.A(mai_mai_n660_), .B(mai_mai_n658_), .Y(mai_mai_n661_));
  OR4        m0639(.A(mai_mai_n661_), .B(mai_mai_n657_), .C(mai_mai_n655_), .D(mai_mai_n653_), .Y(mai_mai_n662_));
  NO3        m0640(.A(mai_mai_n662_), .B(mai_mai_n648_), .C(mai_mai_n645_), .Y(mai_mai_n663_));
  NO2        m0641(.A(mai_mai_n232_), .B(mai_mai_n105_), .Y(mai_mai_n664_));
  NO2        m0642(.A(mai_mai_n664_), .B(mai_mai_n620_), .Y(mai_mai_n665_));
  NA2        m0643(.A(mai_mai_n665_), .B(i_1_), .Y(mai_mai_n666_));
  NO2        m0644(.A(mai_mai_n666_), .B(mai_mai_n614_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n416_), .B(mai_mai_n87_), .Y(mai_mai_n668_));
  NA2        m0646(.A(mai_mai_n667_), .B(mai_mai_n47_), .Y(mai_mai_n669_));
  NO2        m0647(.A(mai_mai_n228_), .B(mai_mai_n45_), .Y(mai_mai_n670_));
  NO3        m0648(.A(mai_mai_n670_), .B(mai_mai_n311_), .C(mai_mai_n233_), .Y(mai_mai_n671_));
  NO2        m0649(.A(mai_mai_n121_), .B(mai_mai_n37_), .Y(mai_mai_n672_));
  NO2        m0650(.A(mai_mai_n672_), .B(i_6_), .Y(mai_mai_n673_));
  NO2        m0651(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n674_));
  NO2        m0652(.A(mai_mai_n674_), .B(mai_mai_n64_), .Y(mai_mai_n675_));
  NO2        m0653(.A(mai_mai_n675_), .B(mai_mai_n637_), .Y(mai_mai_n676_));
  NO4        m0654(.A(mai_mai_n676_), .B(mai_mai_n673_), .C(mai_mai_n671_), .D(i_4_), .Y(mai_mai_n677_));
  NA2        m0655(.A(i_1_), .B(i_3_), .Y(mai_mai_n678_));
  INV        m0656(.A(mai_mai_n677_), .Y(mai_mai_n679_));
  NA4        m0657(.A(mai_mai_n679_), .B(mai_mai_n669_), .C(mai_mai_n663_), .D(mai_mai_n641_), .Y(mai_mai_n680_));
  NO3        m0658(.A(mai_mai_n477_), .B(i_3_), .C(i_7_), .Y(mai_mai_n681_));
  NOi21      m0659(.An(mai_mai_n681_), .B(i_10_), .Y(mai_mai_n682_));
  OA210      m0660(.A0(mai_mai_n682_), .A1(mai_mai_n241_), .B0(mai_mai_n87_), .Y(mai_mai_n683_));
  NA2        m0661(.A(mai_mai_n375_), .B(mai_mai_n374_), .Y(mai_mai_n684_));
  NA3        m0662(.A(mai_mai_n161_), .B(mai_mai_n85_), .C(mai_mai_n87_), .Y(mai_mai_n685_));
  NA2        m0663(.A(mai_mai_n685_), .B(mai_mai_n684_), .Y(mai_mai_n686_));
  OAI210     m0664(.A0(mai_mai_n686_), .A1(mai_mai_n683_), .B0(i_1_), .Y(mai_mai_n687_));
  AOI210     m0665(.A0(mai_mai_n266_), .A1(mai_mai_n101_), .B0(i_1_), .Y(mai_mai_n688_));
  NO2        m0666(.A(mai_mai_n373_), .B(i_2_), .Y(mai_mai_n689_));
  NA2        m0667(.A(mai_mai_n689_), .B(mai_mai_n688_), .Y(mai_mai_n690_));
  OAI210     m0668(.A0(mai_mai_n654_), .A1(mai_mai_n445_), .B0(mai_mai_n690_), .Y(mai_mai_n691_));
  INV        m0669(.A(mai_mai_n691_), .Y(mai_mai_n692_));
  AOI210     m0670(.A0(mai_mai_n692_), .A1(mai_mai_n687_), .B0(i_13_), .Y(mai_mai_n693_));
  OR2        m0671(.A(i_11_), .B(i_7_), .Y(mai_mai_n694_));
  NA3        m0672(.A(mai_mai_n694_), .B(mai_mai_n110_), .C(mai_mai_n142_), .Y(mai_mai_n695_));
  AOI220     m0673(.A0(mai_mai_n471_), .A1(mai_mai_n161_), .B0(mai_mai_n448_), .B1(mai_mai_n142_), .Y(mai_mai_n696_));
  OAI210     m0674(.A0(mai_mai_n696_), .A1(mai_mai_n45_), .B0(mai_mai_n695_), .Y(mai_mai_n697_));
  AOI210     m0675(.A0(mai_mai_n651_), .A1(mai_mai_n55_), .B0(i_12_), .Y(mai_mai_n698_));
  NO2        m0676(.A(mai_mai_n478_), .B(mai_mai_n24_), .Y(mai_mai_n699_));
  AOI220     m0677(.A0(mai_mai_n699_), .A1(mai_mai_n668_), .B0(mai_mai_n241_), .B1(mai_mai_n135_), .Y(mai_mai_n700_));
  OAI220     m0678(.A0(mai_mai_n700_), .A1(mai_mai_n41_), .B0(mai_mai_n1045_), .B1(mai_mai_n96_), .Y(mai_mai_n701_));
  AOI210     m0679(.A0(mai_mai_n697_), .A1(mai_mai_n336_), .B0(mai_mai_n701_), .Y(mai_mai_n702_));
  INV        m0680(.A(mai_mai_n119_), .Y(mai_mai_n703_));
  AOI220     m0681(.A0(mai_mai_n703_), .A1(mai_mai_n73_), .B0(mai_mai_n391_), .B1(mai_mai_n652_), .Y(mai_mai_n704_));
  NO2        m0682(.A(mai_mai_n704_), .B(mai_mai_n238_), .Y(mai_mai_n705_));
  AOI210     m0683(.A0(mai_mai_n445_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n706_));
  NOi31      m0684(.An(mai_mai_n706_), .B(mai_mai_n595_), .C(mai_mai_n45_), .Y(mai_mai_n707_));
  NA2        m0685(.A(mai_mai_n131_), .B(i_13_), .Y(mai_mai_n708_));
  NO2        m0686(.A(mai_mai_n651_), .B(mai_mai_n119_), .Y(mai_mai_n709_));
  INV        m0687(.A(mai_mai_n709_), .Y(mai_mai_n710_));
  OAI220     m0688(.A0(mai_mai_n710_), .A1(mai_mai_n72_), .B0(mai_mai_n708_), .B1(mai_mai_n688_), .Y(mai_mai_n711_));
  NO3        m0689(.A(mai_mai_n72_), .B(mai_mai_n32_), .C(mai_mai_n105_), .Y(mai_mai_n712_));
  NA2        m0690(.A(mai_mai_n26_), .B(mai_mai_n190_), .Y(mai_mai_n713_));
  NA2        m0691(.A(mai_mai_n713_), .B(i_7_), .Y(mai_mai_n714_));
  NO3        m0692(.A(mai_mai_n478_), .B(mai_mai_n232_), .C(mai_mai_n87_), .Y(mai_mai_n715_));
  AOI210     m0693(.A0(mai_mai_n715_), .A1(mai_mai_n714_), .B0(mai_mai_n712_), .Y(mai_mai_n716_));
  AOI220     m0694(.A0(mai_mai_n391_), .A1(mai_mai_n652_), .B0(mai_mai_n95_), .B1(mai_mai_n106_), .Y(mai_mai_n717_));
  OAI220     m0695(.A0(mai_mai_n717_), .A1(mai_mai_n601_), .B0(mai_mai_n716_), .B1(mai_mai_n616_), .Y(mai_mai_n718_));
  NO4        m0696(.A(mai_mai_n718_), .B(mai_mai_n711_), .C(mai_mai_n707_), .D(mai_mai_n705_), .Y(mai_mai_n719_));
  OR2        m0697(.A(i_11_), .B(i_6_), .Y(mai_mai_n720_));
  NA3        m0698(.A(mai_mai_n600_), .B(mai_mai_n713_), .C(i_7_), .Y(mai_mai_n721_));
  AOI210     m0699(.A0(mai_mai_n721_), .A1(mai_mai_n710_), .B0(mai_mai_n720_), .Y(mai_mai_n722_));
  NA3        m0700(.A(mai_mai_n415_), .B(mai_mai_n605_), .C(mai_mai_n101_), .Y(mai_mai_n723_));
  NA2        m0701(.A(mai_mai_n644_), .B(i_13_), .Y(mai_mai_n724_));
  NA2        m0702(.A(mai_mai_n106_), .B(mai_mai_n713_), .Y(mai_mai_n725_));
  NAi21      m0703(.An(i_11_), .B(i_12_), .Y(mai_mai_n726_));
  NOi41      m0704(.An(mai_mai_n115_), .B(mai_mai_n726_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n727_));
  NO3        m0705(.A(mai_mai_n478_), .B(mai_mai_n581_), .C(mai_mai_n606_), .Y(mai_mai_n728_));
  AOI220     m0706(.A0(mai_mai_n728_), .A1(mai_mai_n315_), .B0(mai_mai_n727_), .B1(mai_mai_n725_), .Y(mai_mai_n729_));
  NA3        m0707(.A(mai_mai_n729_), .B(mai_mai_n724_), .C(mai_mai_n723_), .Y(mai_mai_n730_));
  OAI210     m0708(.A0(mai_mai_n730_), .A1(mai_mai_n722_), .B0(mai_mai_n64_), .Y(mai_mai_n731_));
  NO2        m0709(.A(i_2_), .B(i_12_), .Y(mai_mai_n732_));
  NA2        m0710(.A(mai_mai_n372_), .B(mai_mai_n732_), .Y(mai_mai_n733_));
  NA2        m0711(.A(mai_mai_n374_), .B(mai_mai_n372_), .Y(mai_mai_n734_));
  NO2        m0712(.A(mai_mai_n132_), .B(i_2_), .Y(mai_mai_n735_));
  NA2        m0713(.A(mai_mai_n735_), .B(mai_mai_n637_), .Y(mai_mai_n736_));
  NA3        m0714(.A(mai_mai_n736_), .B(mai_mai_n734_), .C(mai_mai_n733_), .Y(mai_mai_n737_));
  NA3        m0715(.A(mai_mai_n737_), .B(mai_mai_n46_), .C(mai_mai_n222_), .Y(mai_mai_n738_));
  NA4        m0716(.A(mai_mai_n738_), .B(mai_mai_n731_), .C(mai_mai_n719_), .D(mai_mai_n702_), .Y(mai_mai_n739_));
  OR4        m0717(.A(mai_mai_n739_), .B(mai_mai_n693_), .C(mai_mai_n680_), .D(mai_mai_n619_), .Y(mai5));
  NA2        m0718(.A(mai_mai_n665_), .B(mai_mai_n269_), .Y(mai_mai_n741_));
  AN2        m0719(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n742_));
  NA3        m0720(.A(mai_mai_n742_), .B(mai_mai_n732_), .C(mai_mai_n112_), .Y(mai_mai_n743_));
  NO2        m0721(.A(mai_mai_n601_), .B(i_11_), .Y(mai_mai_n744_));
  NA2        m0722(.A(mai_mai_n90_), .B(mai_mai_n744_), .Y(mai_mai_n745_));
  NA3        m0723(.A(mai_mai_n745_), .B(mai_mai_n743_), .C(mai_mai_n741_), .Y(mai_mai_n746_));
  NO3        m0724(.A(i_11_), .B(mai_mai_n232_), .C(i_13_), .Y(mai_mai_n747_));
  NO2        m0725(.A(mai_mai_n128_), .B(mai_mai_n23_), .Y(mai_mai_n748_));
  NA2        m0726(.A(i_12_), .B(i_8_), .Y(mai_mai_n749_));
  OAI210     m0727(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n749_), .Y(mai_mai_n750_));
  INV        m0728(.A(mai_mai_n444_), .Y(mai_mai_n751_));
  AOI220     m0729(.A0(mai_mai_n321_), .A1(mai_mai_n573_), .B0(mai_mai_n750_), .B1(mai_mai_n748_), .Y(mai_mai_n752_));
  INV        m0730(.A(mai_mai_n752_), .Y(mai_mai_n753_));
  NO2        m0731(.A(mai_mai_n753_), .B(mai_mai_n746_), .Y(mai_mai_n754_));
  INV        m0732(.A(mai_mai_n168_), .Y(mai_mai_n755_));
  INV        m0733(.A(mai_mai_n241_), .Y(mai_mai_n756_));
  OAI210     m0734(.A0(mai_mai_n689_), .A1(mai_mai_n446_), .B0(mai_mai_n115_), .Y(mai_mai_n757_));
  AOI210     m0735(.A0(mai_mai_n757_), .A1(mai_mai_n756_), .B0(mai_mai_n755_), .Y(mai_mai_n758_));
  NO2        m0736(.A(mai_mai_n454_), .B(mai_mai_n26_), .Y(mai_mai_n759_));
  NO2        m0737(.A(mai_mai_n759_), .B(mai_mai_n420_), .Y(mai_mai_n760_));
  NA2        m0738(.A(mai_mai_n760_), .B(i_2_), .Y(mai_mai_n761_));
  INV        m0739(.A(mai_mai_n761_), .Y(mai_mai_n762_));
  AOI210     m0740(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n417_), .Y(mai_mai_n763_));
  AOI210     m0741(.A0(mai_mai_n763_), .A1(mai_mai_n762_), .B0(mai_mai_n758_), .Y(mai_mai_n764_));
  NO2        m0742(.A(mai_mai_n187_), .B(mai_mai_n129_), .Y(mai_mai_n765_));
  OAI210     m0743(.A0(mai_mai_n765_), .A1(mai_mai_n748_), .B0(i_2_), .Y(mai_mai_n766_));
  INV        m0744(.A(mai_mai_n169_), .Y(mai_mai_n767_));
  NO3        m0745(.A(mai_mai_n621_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n768_));
  AOI210     m0746(.A0(mai_mai_n767_), .A1(mai_mai_n90_), .B0(mai_mai_n768_), .Y(mai_mai_n769_));
  AOI210     m0747(.A0(mai_mai_n769_), .A1(mai_mai_n766_), .B0(mai_mai_n190_), .Y(mai_mai_n770_));
  OA210      m0748(.A0(mai_mai_n622_), .A1(mai_mai_n130_), .B0(i_13_), .Y(mai_mai_n771_));
  NA2        m0749(.A(mai_mai_n196_), .B(mai_mai_n199_), .Y(mai_mai_n772_));
  NA2        m0750(.A(mai_mai_n154_), .B(mai_mai_n596_), .Y(mai_mai_n773_));
  AOI210     m0751(.A0(mai_mai_n773_), .A1(mai_mai_n772_), .B0(mai_mai_n377_), .Y(mai_mai_n774_));
  AOI210     m0752(.A0(mai_mai_n204_), .A1(mai_mai_n152_), .B0(mai_mai_n516_), .Y(mai_mai_n775_));
  NA2        m0753(.A(mai_mai_n775_), .B(mai_mai_n420_), .Y(mai_mai_n776_));
  NO2        m0754(.A(mai_mai_n106_), .B(mai_mai_n45_), .Y(mai_mai_n777_));
  INV        m0755(.A(mai_mai_n304_), .Y(mai_mai_n778_));
  NA4        m0756(.A(mai_mai_n778_), .B(mai_mai_n309_), .C(mai_mai_n128_), .D(mai_mai_n43_), .Y(mai_mai_n779_));
  OAI210     m0757(.A0(mai_mai_n779_), .A1(mai_mai_n777_), .B0(mai_mai_n776_), .Y(mai_mai_n780_));
  NO4        m0758(.A(mai_mai_n780_), .B(mai_mai_n774_), .C(mai_mai_n771_), .D(mai_mai_n770_), .Y(mai_mai_n781_));
  NA2        m0759(.A(mai_mai_n573_), .B(mai_mai_n28_), .Y(mai_mai_n782_));
  NA2        m0760(.A(mai_mai_n747_), .B(mai_mai_n276_), .Y(mai_mai_n783_));
  NA2        m0761(.A(mai_mai_n783_), .B(mai_mai_n782_), .Y(mai_mai_n784_));
  NO2        m0762(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n785_));
  NO2        m0763(.A(mai_mai_n785_), .B(mai_mai_n130_), .Y(mai_mai_n786_));
  NO2        m0764(.A(mai_mai_n786_), .B(mai_mai_n596_), .Y(mai_mai_n787_));
  AOI220     m0765(.A0(mai_mai_n787_), .A1(mai_mai_n36_), .B0(mai_mai_n784_), .B1(mai_mai_n47_), .Y(mai_mai_n788_));
  NA4        m0766(.A(mai_mai_n788_), .B(mai_mai_n781_), .C(mai_mai_n764_), .D(mai_mai_n754_), .Y(mai6));
  NO3        m0767(.A(mai_mai_n252_), .B(mai_mai_n310_), .C(i_1_), .Y(mai_mai_n790_));
  NO2        m0768(.A(mai_mai_n182_), .B(mai_mai_n143_), .Y(mai_mai_n791_));
  OAI210     m0769(.A0(mai_mai_n791_), .A1(mai_mai_n790_), .B0(mai_mai_n735_), .Y(mai_mai_n792_));
  NO2        m0770(.A(mai_mai_n218_), .B(mai_mai_n485_), .Y(mai_mai_n793_));
  NO2        m0771(.A(i_11_), .B(i_9_), .Y(mai_mai_n794_));
  INV        m0772(.A(mai_mai_n332_), .Y(mai_mai_n795_));
  AO210      m0773(.A0(mai_mai_n795_), .A1(mai_mai_n792_), .B0(i_12_), .Y(mai_mai_n796_));
  NA2        m0774(.A(mai_mai_n378_), .B(mai_mai_n339_), .Y(mai_mai_n797_));
  NA2        m0775(.A(mai_mai_n581_), .B(mai_mai_n64_), .Y(mai_mai_n798_));
  NA2        m0776(.A(mai_mai_n682_), .B(mai_mai_n72_), .Y(mai_mai_n799_));
  BUFFER     m0777(.A(mai_mai_n627_), .Y(mai_mai_n800_));
  NA4        m0778(.A(mai_mai_n800_), .B(mai_mai_n799_), .C(mai_mai_n798_), .D(mai_mai_n797_), .Y(mai_mai_n801_));
  INV        m0779(.A(mai_mai_n194_), .Y(mai_mai_n802_));
  AOI220     m0780(.A0(mai_mai_n802_), .A1(mai_mai_n794_), .B0(mai_mai_n801_), .B1(mai_mai_n74_), .Y(mai_mai_n803_));
  INV        m0781(.A(mai_mai_n331_), .Y(mai_mai_n804_));
  NA2        m0782(.A(mai_mai_n76_), .B(mai_mai_n135_), .Y(mai_mai_n805_));
  INV        m0783(.A(mai_mai_n128_), .Y(mai_mai_n806_));
  NA2        m0784(.A(mai_mai_n806_), .B(mai_mai_n47_), .Y(mai_mai_n807_));
  AOI210     m0785(.A0(mai_mai_n807_), .A1(mai_mai_n805_), .B0(mai_mai_n804_), .Y(mai_mai_n808_));
  NO3        m0786(.A(mai_mai_n248_), .B(mai_mai_n136_), .C(i_9_), .Y(mai_mai_n809_));
  NA2        m0787(.A(mai_mai_n809_), .B(mai_mai_n785_), .Y(mai_mai_n810_));
  AOI210     m0788(.A0(mai_mai_n810_), .A1(mai_mai_n514_), .B0(mai_mai_n182_), .Y(mai_mai_n811_));
  NO2        m0789(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n812_));
  NA3        m0790(.A(mai_mai_n812_), .B(mai_mai_n473_), .C(mai_mai_n395_), .Y(mai_mai_n813_));
  NAi32      m0791(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n814_));
  NO2        m0792(.A(mai_mai_n720_), .B(mai_mai_n814_), .Y(mai_mai_n815_));
  OAI210     m0793(.A0(mai_mai_n681_), .A1(mai_mai_n563_), .B0(mai_mai_n562_), .Y(mai_mai_n816_));
  NAi31      m0794(.An(mai_mai_n815_), .B(mai_mai_n816_), .C(mai_mai_n813_), .Y(mai_mai_n817_));
  OR3        m0795(.A(mai_mai_n817_), .B(mai_mai_n811_), .C(mai_mai_n808_), .Y(mai_mai_n818_));
  NO2        m0796(.A(mai_mai_n694_), .B(i_2_), .Y(mai_mai_n819_));
  NA2        m0797(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n820_));
  NO2        m0798(.A(mai_mai_n820_), .B(mai_mai_n414_), .Y(mai_mai_n821_));
  NA2        m0799(.A(mai_mai_n821_), .B(mai_mai_n819_), .Y(mai_mai_n822_));
  OR2        m0800(.A(mai_mai_n622_), .B(mai_mai_n446_), .Y(mai_mai_n823_));
  NA3        m0801(.A(mai_mai_n823_), .B(mai_mai_n151_), .C(mai_mai_n70_), .Y(mai_mai_n824_));
  AO210      m0802(.A0(mai_mai_n492_), .A1(mai_mai_n751_), .B0(mai_mai_n36_), .Y(mai_mai_n825_));
  NA3        m0803(.A(mai_mai_n825_), .B(mai_mai_n824_), .C(mai_mai_n822_), .Y(mai_mai_n826_));
  OAI210     m0804(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n88_), .Y(mai_mai_n827_));
  AOI220     m0805(.A0(mai_mai_n827_), .A1(mai_mai_n562_), .B0(mai_mai_n793_), .B1(mai_mai_n714_), .Y(mai_mai_n828_));
  NA3        m0806(.A(mai_mai_n377_), .B(mai_mai_n234_), .C(mai_mai_n151_), .Y(mai_mai_n829_));
  NA2        m0807(.A(mai_mai_n402_), .B(mai_mai_n71_), .Y(mai_mai_n830_));
  NA4        m0808(.A(mai_mai_n830_), .B(mai_mai_n829_), .C(mai_mai_n828_), .D(mai_mai_n604_), .Y(mai_mai_n831_));
  AO210      m0809(.A0(mai_mai_n516_), .A1(mai_mai_n47_), .B0(mai_mai_n89_), .Y(mai_mai_n832_));
  NA3        m0810(.A(mai_mai_n832_), .B(mai_mai_n483_), .C(mai_mai_n215_), .Y(mai_mai_n833_));
  AOI210     m0811(.A0(mai_mai_n446_), .A1(mai_mai_n444_), .B0(mai_mai_n561_), .Y(mai_mai_n834_));
  NO2        m0812(.A(mai_mai_n612_), .B(mai_mai_n106_), .Y(mai_mai_n835_));
  OAI210     m0813(.A0(mai_mai_n835_), .A1(mai_mai_n116_), .B0(mai_mai_n413_), .Y(mai_mai_n836_));
  NA2        m0814(.A(mai_mai_n240_), .B(mai_mai_n47_), .Y(mai_mai_n837_));
  INV        m0815(.A(mai_mai_n585_), .Y(mai_mai_n838_));
  NA3        m0816(.A(mai_mai_n838_), .B(mai_mai_n331_), .C(i_7_), .Y(mai_mai_n839_));
  NA4        m0817(.A(mai_mai_n839_), .B(mai_mai_n836_), .C(mai_mai_n834_), .D(mai_mai_n833_), .Y(mai_mai_n840_));
  NO4        m0818(.A(mai_mai_n840_), .B(mai_mai_n831_), .C(mai_mai_n826_), .D(mai_mai_n818_), .Y(mai_mai_n841_));
  NA4        m0819(.A(mai_mai_n841_), .B(mai_mai_n803_), .C(mai_mai_n796_), .D(mai_mai_n385_), .Y(mai3));
  NA2        m0820(.A(i_12_), .B(i_10_), .Y(mai_mai_n843_));
  NA2        m0821(.A(i_6_), .B(i_7_), .Y(mai_mai_n844_));
  NO2        m0822(.A(mai_mai_n844_), .B(i_0_), .Y(mai_mai_n845_));
  NO2        m0823(.A(i_11_), .B(mai_mai_n232_), .Y(mai_mai_n846_));
  OAI210     m0824(.A0(mai_mai_n845_), .A1(mai_mai_n292_), .B0(mai_mai_n846_), .Y(mai_mai_n847_));
  NO2        m0825(.A(mai_mai_n847_), .B(mai_mai_n190_), .Y(mai_mai_n848_));
  NO3        m0826(.A(mai_mai_n450_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n849_));
  OA210      m0827(.A0(mai_mai_n849_), .A1(mai_mai_n848_), .B0(mai_mai_n171_), .Y(mai_mai_n850_));
  NA2        m0828(.A(mai_mai_n829_), .B(mai_mai_n376_), .Y(mai_mai_n851_));
  NA2        m0829(.A(mai_mai_n851_), .B(mai_mai_n40_), .Y(mai_mai_n852_));
  NOi21      m0830(.An(mai_mai_n100_), .B(mai_mai_n760_), .Y(mai_mai_n853_));
  NO3        m0831(.A(mai_mai_n632_), .B(mai_mai_n454_), .C(mai_mai_n135_), .Y(mai_mai_n854_));
  NA2        m0832(.A(mai_mai_n415_), .B(mai_mai_n46_), .Y(mai_mai_n855_));
  AN2        m0833(.A(mai_mai_n452_), .B(mai_mai_n56_), .Y(mai_mai_n856_));
  NO3        m0834(.A(mai_mai_n856_), .B(mai_mai_n854_), .C(mai_mai_n853_), .Y(mai_mai_n857_));
  AOI210     m0835(.A0(mai_mai_n857_), .A1(mai_mai_n852_), .B0(mai_mai_n49_), .Y(mai_mai_n858_));
  NO4        m0836(.A(mai_mai_n381_), .B(mai_mai_n388_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n859_));
  NA2        m0837(.A(mai_mai_n182_), .B(mai_mai_n569_), .Y(mai_mai_n860_));
  NOi21      m0838(.An(mai_mai_n860_), .B(mai_mai_n859_), .Y(mai_mai_n861_));
  NA2        m0839(.A(mai_mai_n706_), .B(mai_mai_n674_), .Y(mai_mai_n862_));
  NA2        m0840(.A(mai_mai_n337_), .B(mai_mai_n434_), .Y(mai_mai_n863_));
  OAI220     m0841(.A0(mai_mai_n863_), .A1(mai_mai_n862_), .B0(mai_mai_n861_), .B1(mai_mai_n64_), .Y(mai_mai_n864_));
  NOi21      m0842(.An(i_5_), .B(i_9_), .Y(mai_mai_n865_));
  NA2        m0843(.A(mai_mai_n865_), .B(mai_mai_n442_), .Y(mai_mai_n866_));
  BUFFER     m0844(.A(mai_mai_n266_), .Y(mai_mai_n867_));
  NA2        m0845(.A(mai_mai_n867_), .B(mai_mai_n475_), .Y(mai_mai_n868_));
  NO2        m0846(.A(mai_mai_n172_), .B(mai_mai_n152_), .Y(mai_mai_n869_));
  NO2        m0847(.A(mai_mai_n868_), .B(mai_mai_n866_), .Y(mai_mai_n870_));
  NO4        m0848(.A(mai_mai_n870_), .B(mai_mai_n864_), .C(mai_mai_n858_), .D(mai_mai_n850_), .Y(mai_mai_n871_));
  NA2        m0849(.A(mai_mai_n182_), .B(mai_mai_n24_), .Y(mai_mai_n872_));
  NO2        m0850(.A(mai_mai_n672_), .B(mai_mai_n593_), .Y(mai_mai_n873_));
  NO2        m0851(.A(mai_mai_n873_), .B(mai_mai_n872_), .Y(mai_mai_n874_));
  NA2        m0852(.A(mai_mai_n315_), .B(mai_mai_n133_), .Y(mai_mai_n875_));
  NAi21      m0853(.An(mai_mai_n162_), .B(mai_mai_n434_), .Y(mai_mai_n876_));
  OAI220     m0854(.A0(mai_mai_n876_), .A1(mai_mai_n837_), .B0(mai_mai_n875_), .B1(mai_mai_n404_), .Y(mai_mai_n877_));
  NO2        m0855(.A(mai_mai_n877_), .B(mai_mai_n874_), .Y(mai_mai_n878_));
  NO2        m0856(.A(mai_mai_n395_), .B(mai_mai_n296_), .Y(mai_mai_n879_));
  NA2        m0857(.A(mai_mai_n879_), .B(mai_mai_n709_), .Y(mai_mai_n880_));
  NA2        m0858(.A(mai_mai_n570_), .B(i_0_), .Y(mai_mai_n881_));
  NO3        m0859(.A(mai_mai_n881_), .B(mai_mai_n390_), .C(mai_mai_n90_), .Y(mai_mai_n882_));
  NO4        m0860(.A(mai_mai_n584_), .B(mai_mai_n212_), .C(mai_mai_n417_), .D(mai_mai_n414_), .Y(mai_mai_n883_));
  AOI210     m0861(.A0(mai_mai_n883_), .A1(i_11_), .B0(mai_mai_n882_), .Y(mai_mai_n884_));
  INV        m0862(.A(mai_mai_n473_), .Y(mai_mai_n885_));
  AN2        m0863(.A(mai_mai_n100_), .B(mai_mai_n239_), .Y(mai_mai_n886_));
  NA2        m0864(.A(mai_mai_n747_), .B(mai_mai_n332_), .Y(mai_mai_n887_));
  AOI210     m0865(.A0(mai_mai_n483_), .A1(mai_mai_n90_), .B0(mai_mai_n59_), .Y(mai_mai_n888_));
  OAI220     m0866(.A0(mai_mai_n888_), .A1(mai_mai_n887_), .B0(mai_mai_n660_), .B1(mai_mai_n534_), .Y(mai_mai_n889_));
  NO2        m0867(.A(mai_mai_n250_), .B(mai_mai_n155_), .Y(mai_mai_n890_));
  NA2        m0868(.A(i_0_), .B(i_10_), .Y(mai_mai_n891_));
  AN2        m0869(.A(mai_mai_n890_), .B(i_6_), .Y(mai_mai_n892_));
  NO3        m0870(.A(mai_mai_n892_), .B(mai_mai_n889_), .C(mai_mai_n886_), .Y(mai_mai_n893_));
  NA4        m0871(.A(mai_mai_n893_), .B(mai_mai_n884_), .C(mai_mai_n880_), .D(mai_mai_n878_), .Y(mai_mai_n894_));
  NO2        m0872(.A(mai_mai_n107_), .B(mai_mai_n37_), .Y(mai_mai_n895_));
  NA2        m0873(.A(i_11_), .B(i_9_), .Y(mai_mai_n896_));
  NO3        m0874(.A(i_12_), .B(mai_mai_n896_), .C(mai_mai_n603_), .Y(mai_mai_n897_));
  AN2        m0875(.A(mai_mai_n897_), .B(mai_mai_n895_), .Y(mai_mai_n898_));
  NO2        m0876(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n899_));
  NA2        m0877(.A(mai_mai_n400_), .B(mai_mai_n176_), .Y(mai_mai_n900_));
  NA2        m0878(.A(mai_mai_n900_), .B(mai_mai_n160_), .Y(mai_mai_n901_));
  NO2        m0879(.A(mai_mai_n896_), .B(mai_mai_n74_), .Y(mai_mai_n902_));
  AOI210     m0880(.A0(mai_mai_n375_), .A1(mai_mai_n42_), .B0(mai_mai_n412_), .Y(mai_mai_n903_));
  NO2        m0881(.A(mai_mai_n903_), .B(mai_mai_n866_), .Y(mai_mai_n904_));
  NO3        m0882(.A(mai_mai_n904_), .B(mai_mai_n901_), .C(mai_mai_n898_), .Y(mai_mai_n905_));
  NA2        m0883(.A(mai_mai_n659_), .B(mai_mai_n125_), .Y(mai_mai_n906_));
  NO2        m0884(.A(i_6_), .B(mai_mai_n906_), .Y(mai_mai_n907_));
  AOI210     m0885(.A0(mai_mai_n445_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n908_));
  NA2        m0886(.A(mai_mai_n168_), .B(mai_mai_n107_), .Y(mai_mai_n909_));
  NOi32      m0887(.An(mai_mai_n908_), .Bn(mai_mai_n185_), .C(mai_mai_n909_), .Y(mai_mai_n910_));
  NA2        m0888(.A(mai_mai_n605_), .B(mai_mai_n332_), .Y(mai_mai_n911_));
  NO2        m0889(.A(mai_mai_n911_), .B(mai_mai_n855_), .Y(mai_mai_n912_));
  NO3        m0890(.A(mai_mai_n912_), .B(mai_mai_n910_), .C(mai_mai_n907_), .Y(mai_mai_n913_));
  NOi21      m0891(.An(i_7_), .B(i_5_), .Y(mai_mai_n914_));
  NOi31      m0892(.An(mai_mai_n914_), .B(i_0_), .C(mai_mai_n726_), .Y(mai_mai_n915_));
  NA3        m0893(.A(mai_mai_n915_), .B(mai_mai_n389_), .C(i_6_), .Y(mai_mai_n916_));
  OA210      m0894(.A0(mai_mai_n909_), .A1(mai_mai_n514_), .B0(mai_mai_n916_), .Y(mai_mai_n917_));
  NO3        m0895(.A(mai_mai_n407_), .B(mai_mai_n364_), .C(mai_mai_n363_), .Y(mai_mai_n918_));
  NO2        m0896(.A(mai_mai_n260_), .B(mai_mai_n322_), .Y(mai_mai_n919_));
  NO2        m0897(.A(mai_mai_n726_), .B(mai_mai_n255_), .Y(mai_mai_n920_));
  AOI210     m0898(.A0(mai_mai_n920_), .A1(mai_mai_n919_), .B0(mai_mai_n918_), .Y(mai_mai_n921_));
  NA4        m0899(.A(mai_mai_n921_), .B(mai_mai_n917_), .C(mai_mai_n913_), .D(mai_mai_n905_), .Y(mai_mai_n922_));
  NO2        m0900(.A(mai_mai_n872_), .B(mai_mai_n235_), .Y(mai_mai_n923_));
  AN2        m0901(.A(mai_mai_n336_), .B(mai_mai_n332_), .Y(mai_mai_n924_));
  AN2        m0902(.A(mai_mai_n924_), .B(mai_mai_n869_), .Y(mai_mai_n925_));
  OAI210     m0903(.A0(mai_mai_n925_), .A1(mai_mai_n923_), .B0(i_10_), .Y(mai_mai_n926_));
  NO2        m0904(.A(mai_mai_n843_), .B(mai_mai_n321_), .Y(mai_mai_n927_));
  OA210      m0905(.A0(mai_mai_n473_), .A1(mai_mai_n221_), .B0(mai_mai_n472_), .Y(mai_mai_n928_));
  NA2        m0906(.A(mai_mai_n927_), .B(mai_mai_n902_), .Y(mai_mai_n929_));
  NA3        m0907(.A(mai_mai_n472_), .B(mai_mai_n415_), .C(mai_mai_n46_), .Y(mai_mai_n930_));
  OAI210     m0908(.A0(mai_mai_n876_), .A1(mai_mai_n885_), .B0(mai_mai_n930_), .Y(mai_mai_n931_));
  NO2        m0909(.A(mai_mai_n253_), .B(mai_mai_n47_), .Y(mai_mai_n932_));
  NA2        m0910(.A(mai_mai_n902_), .B(mai_mai_n309_), .Y(mai_mai_n933_));
  OAI210     m0911(.A0(mai_mai_n932_), .A1(mai_mai_n184_), .B0(mai_mai_n933_), .Y(mai_mai_n934_));
  AOI220     m0912(.A0(mai_mai_n934_), .A1(mai_mai_n473_), .B0(mai_mai_n931_), .B1(mai_mai_n74_), .Y(mai_mai_n935_));
  NA2        m0913(.A(mai_mai_n96_), .B(mai_mai_n45_), .Y(mai_mai_n936_));
  NO2        m0914(.A(mai_mai_n76_), .B(mai_mai_n749_), .Y(mai_mai_n937_));
  AOI220     m0915(.A0(mai_mai_n937_), .A1(mai_mai_n936_), .B0(mai_mai_n171_), .B1(mai_mai_n593_), .Y(mai_mai_n938_));
  NO2        m0916(.A(mai_mai_n938_), .B(mai_mai_n48_), .Y(mai_mai_n939_));
  NA2        m0917(.A(mai_mai_n699_), .B(mai_mai_n543_), .Y(mai_mai_n940_));
  NAi21      m0918(.An(i_9_), .B(i_5_), .Y(mai_mai_n941_));
  NO2        m0919(.A(mai_mai_n941_), .B(mai_mai_n407_), .Y(mai_mai_n942_));
  NO2        m0920(.A(mai_mai_n599_), .B(mai_mai_n109_), .Y(mai_mai_n943_));
  AOI220     m0921(.A0(mai_mai_n943_), .A1(i_0_), .B0(mai_mai_n942_), .B1(mai_mai_n622_), .Y(mai_mai_n944_));
  OAI220     m0922(.A0(mai_mai_n944_), .A1(mai_mai_n87_), .B0(mai_mai_n940_), .B1(mai_mai_n169_), .Y(mai_mai_n945_));
  NO3        m0923(.A(mai_mai_n945_), .B(mai_mai_n939_), .C(mai_mai_n519_), .Y(mai_mai_n946_));
  NA4        m0924(.A(mai_mai_n946_), .B(mai_mai_n935_), .C(mai_mai_n929_), .D(mai_mai_n926_), .Y(mai_mai_n947_));
  NO3        m0925(.A(mai_mai_n947_), .B(mai_mai_n922_), .C(mai_mai_n894_), .Y(mai_mai_n948_));
  NO2        m0926(.A(i_0_), .B(mai_mai_n726_), .Y(mai_mai_n949_));
  NA2        m0927(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n950_));
  INV        m0928(.A(mai_mai_n950_), .Y(mai_mai_n951_));
  NO3        m0929(.A(mai_mai_n109_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n952_));
  AO220      m0930(.A0(mai_mai_n952_), .A1(mai_mai_n951_), .B0(mai_mai_n949_), .B1(mai_mai_n171_), .Y(mai_mai_n953_));
  AOI210     m0931(.A0(mai_mai_n798_), .A1(mai_mai_n684_), .B0(mai_mai_n909_), .Y(mai_mai_n954_));
  AOI210     m0932(.A0(mai_mai_n953_), .A1(mai_mai_n352_), .B0(mai_mai_n954_), .Y(mai_mai_n955_));
  NA2        m0933(.A(mai_mai_n735_), .B(mai_mai_n150_), .Y(mai_mai_n956_));
  INV        m0934(.A(mai_mai_n956_), .Y(mai_mai_n957_));
  NA3        m0935(.A(mai_mai_n957_), .B(mai_mai_n674_), .C(mai_mai_n74_), .Y(mai_mai_n958_));
  NO2        m0936(.A(mai_mai_n816_), .B(mai_mai_n407_), .Y(mai_mai_n959_));
  NA3        m0937(.A(mai_mai_n845_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n960_));
  NA2        m0938(.A(mai_mai_n846_), .B(i_9_), .Y(mai_mai_n961_));
  AOI210     m0939(.A0(mai_mai_n960_), .A1(mai_mai_n496_), .B0(mai_mai_n961_), .Y(mai_mai_n962_));
  OAI210     m0940(.A0(mai_mai_n240_), .A1(i_9_), .B0(mai_mai_n225_), .Y(mai_mai_n963_));
  AOI210     m0941(.A0(mai_mai_n963_), .A1(mai_mai_n881_), .B0(mai_mai_n155_), .Y(mai_mai_n964_));
  NO3        m0942(.A(mai_mai_n964_), .B(mai_mai_n962_), .C(mai_mai_n959_), .Y(mai_mai_n965_));
  NA3        m0943(.A(mai_mai_n965_), .B(mai_mai_n958_), .C(mai_mai_n955_), .Y(mai_mai_n966_));
  NA3        m0944(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n967_));
  NA2        m0945(.A(mai_mai_n899_), .B(mai_mai_n486_), .Y(mai_mai_n968_));
  AOI210     m0946(.A0(mai_mai_n967_), .A1(mai_mai_n162_), .B0(mai_mai_n968_), .Y(mai_mai_n969_));
  INV        m0947(.A(mai_mai_n969_), .Y(mai_mai_n970_));
  NO3        m0948(.A(mai_mai_n891_), .B(mai_mai_n865_), .C(mai_mai_n187_), .Y(mai_mai_n971_));
  AOI220     m0949(.A0(mai_mai_n971_), .A1(i_11_), .B0(mai_mai_n567_), .B1(mai_mai_n76_), .Y(mai_mai_n972_));
  NO3        m0950(.A(mai_mai_n206_), .B(mai_mai_n388_), .C(i_0_), .Y(mai_mai_n973_));
  OAI210     m0951(.A0(mai_mai_n973_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n974_));
  NA3        m0952(.A(mai_mai_n974_), .B(mai_mai_n972_), .C(mai_mai_n970_), .Y(mai_mai_n975_));
  NO2        m0953(.A(mai_mai_n238_), .B(mai_mai_n96_), .Y(mai_mai_n976_));
  AOI210     m0954(.A0(mai_mai_n976_), .A1(mai_mai_n949_), .B0(mai_mai_n113_), .Y(mai_mai_n977_));
  OR2        m0955(.A(mai_mai_n977_), .B(i_5_), .Y(mai_mai_n978_));
  AOI210     m0956(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n172_), .Y(mai_mai_n979_));
  NA2        m0957(.A(mai_mai_n979_), .B(mai_mai_n928_), .Y(mai_mai_n980_));
  NO3        m0958(.A(mai_mai_n855_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n981_));
  NA2        m0959(.A(mai_mai_n491_), .B(mai_mai_n484_), .Y(mai_mai_n982_));
  NO2        m0960(.A(mai_mai_n982_), .B(mai_mai_n981_), .Y(mai_mai_n983_));
  NA3        m0961(.A(mai_mai_n395_), .B(mai_mai_n168_), .C(mai_mai_n167_), .Y(mai_mai_n984_));
  NA3        m0962(.A(mai_mai_n899_), .B(mai_mai_n292_), .C(mai_mai_n225_), .Y(mai_mai_n985_));
  NA2        m0963(.A(mai_mai_n985_), .B(mai_mai_n984_), .Y(mai_mai_n986_));
  NOi31      m0964(.An(mai_mai_n394_), .B(mai_mai_n950_), .C(mai_mai_n235_), .Y(mai_mai_n987_));
  NO3        m0965(.A(mai_mai_n896_), .B(mai_mai_n215_), .C(mai_mai_n187_), .Y(mai_mai_n988_));
  NO3        m0966(.A(mai_mai_n988_), .B(mai_mai_n987_), .C(mai_mai_n986_), .Y(mai_mai_n989_));
  NA4        m0967(.A(mai_mai_n989_), .B(mai_mai_n983_), .C(mai_mai_n980_), .D(mai_mai_n978_), .Y(mai_mai_n990_));
  INV        m0968(.A(mai_mai_n615_), .Y(mai_mai_n991_));
  NO3        m0969(.A(mai_mai_n991_), .B(mai_mai_n557_), .C(mai_mai_n350_), .Y(mai_mai_n992_));
  NO2        m0970(.A(mai_mai_n87_), .B(i_5_), .Y(mai_mai_n993_));
  NA3        m0971(.A(mai_mai_n846_), .B(mai_mai_n114_), .C(mai_mai_n128_), .Y(mai_mai_n994_));
  INV        m0972(.A(mai_mai_n994_), .Y(mai_mai_n995_));
  AOI210     m0973(.A0(mai_mai_n995_), .A1(mai_mai_n993_), .B0(mai_mai_n992_), .Y(mai_mai_n996_));
  NAi21      m0974(.An(mai_mai_n237_), .B(mai_mai_n238_), .Y(mai_mai_n997_));
  NO4        m0975(.A(mai_mai_n235_), .B(mai_mai_n206_), .C(i_0_), .D(i_12_), .Y(mai_mai_n998_));
  NA2        m0976(.A(mai_mai_n998_), .B(mai_mai_n997_), .Y(mai_mai_n999_));
  NA2        m0977(.A(mai_mai_n999_), .B(mai_mai_n996_), .Y(mai_mai_n1000_));
  NO4        m0978(.A(mai_mai_n1000_), .B(mai_mai_n990_), .C(mai_mai_n975_), .D(mai_mai_n966_), .Y(mai_mai_n1001_));
  OAI210     m0979(.A0(mai_mai_n819_), .A1(mai_mai_n812_), .B0(mai_mai_n37_), .Y(mai_mai_n1002_));
  NA3        m0980(.A(mai_mai_n908_), .B(mai_mai_n372_), .C(i_5_), .Y(mai_mai_n1003_));
  NA3        m0981(.A(mai_mai_n1003_), .B(mai_mai_n1002_), .C(mai_mai_n611_), .Y(mai_mai_n1004_));
  NA2        m0982(.A(mai_mai_n1004_), .B(mai_mai_n202_), .Y(mai_mai_n1005_));
  NA2        m0983(.A(mai_mai_n183_), .B(mai_mai_n185_), .Y(mai_mai_n1006_));
  AO210      m0984(.A0(mai_mai_n694_), .A1(mai_mai_n33_), .B0(mai_mai_n1006_), .Y(mai_mai_n1007_));
  OAI210     m0985(.A0(mai_mai_n615_), .A1(mai_mai_n613_), .B0(mai_mai_n321_), .Y(mai_mai_n1008_));
  NAi31      m0986(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n1009_));
  NO2        m0987(.A(mai_mai_n71_), .B(mai_mai_n1009_), .Y(mai_mai_n1010_));
  INV        m0988(.A(mai_mai_n1010_), .Y(mai_mai_n1011_));
  NA3        m0989(.A(mai_mai_n1011_), .B(mai_mai_n1008_), .C(mai_mai_n1007_), .Y(mai_mai_n1012_));
  NO4        m0990(.A(mai_mai_n228_), .B(mai_mai_n149_), .C(mai_mai_n678_), .D(mai_mai_n37_), .Y(mai_mai_n1013_));
  NO2        m0991(.A(mai_mai_n1013_), .B(mai_mai_n883_), .Y(mai_mai_n1014_));
  INV        m0992(.A(mai_mai_n1014_), .Y(mai_mai_n1015_));
  AOI210     m0993(.A0(mai_mai_n1012_), .A1(mai_mai_n49_), .B0(mai_mai_n1015_), .Y(mai_mai_n1016_));
  AOI210     m0994(.A0(mai_mai_n1016_), .A1(mai_mai_n1005_), .B0(mai_mai_n74_), .Y(mai_mai_n1017_));
  NO2        m0995(.A(mai_mai_n564_), .B(mai_mai_n384_), .Y(mai_mai_n1018_));
  NO2        m0996(.A(mai_mai_n1018_), .B(mai_mai_n755_), .Y(mai_mai_n1019_));
  OAI210     m0997(.A0(mai_mai_n81_), .A1(mai_mai_n55_), .B0(mai_mai_n112_), .Y(mai_mai_n1020_));
  NA2        m0998(.A(mai_mai_n1020_), .B(mai_mai_n77_), .Y(mai_mai_n1021_));
  AOI210     m0999(.A0(mai_mai_n979_), .A1(mai_mai_n899_), .B0(mai_mai_n915_), .Y(mai_mai_n1022_));
  AOI210     m1000(.A0(mai_mai_n1022_), .A1(mai_mai_n1021_), .B0(mai_mai_n678_), .Y(mai_mai_n1023_));
  NA2        m1001(.A(mai_mai_n260_), .B(mai_mai_n58_), .Y(mai_mai_n1024_));
  AOI220     m1002(.A0(mai_mai_n1024_), .A1(mai_mai_n77_), .B0(mai_mai_n351_), .B1(mai_mai_n252_), .Y(mai_mai_n1025_));
  NO2        m1003(.A(mai_mai_n1025_), .B(mai_mai_n232_), .Y(mai_mai_n1026_));
  NA3        m1004(.A(mai_mai_n100_), .B(mai_mai_n310_), .C(mai_mai_n31_), .Y(mai_mai_n1027_));
  INV        m1005(.A(mai_mai_n1027_), .Y(mai_mai_n1028_));
  NO3        m1006(.A(mai_mai_n1028_), .B(mai_mai_n1026_), .C(mai_mai_n1023_), .Y(mai_mai_n1029_));
  OAI210     m1007(.A0(mai_mai_n268_), .A1(mai_mai_n158_), .B0(mai_mai_n90_), .Y(mai_mai_n1030_));
  NA3        m1008(.A(mai_mai_n759_), .B(mai_mai_n292_), .C(mai_mai_n81_), .Y(mai_mai_n1031_));
  AOI210     m1009(.A0(mai_mai_n1031_), .A1(mai_mai_n1030_), .B0(i_11_), .Y(mai_mai_n1032_));
  NO3        m1010(.A(mai_mai_n60_), .B(mai_mai_n59_), .C(i_4_), .Y(mai_mai_n1033_));
  OAI210     m1011(.A0(mai_mai_n919_), .A1(mai_mai_n310_), .B0(mai_mai_n1033_), .Y(mai_mai_n1034_));
  NO2        m1012(.A(mai_mai_n1034_), .B(mai_mai_n726_), .Y(mai_mai_n1035_));
  NO4        m1013(.A(mai_mai_n941_), .B(mai_mai_n477_), .C(mai_mai_n249_), .D(mai_mai_n248_), .Y(mai_mai_n1036_));
  NO2        m1014(.A(mai_mai_n1036_), .B(mai_mai_n561_), .Y(mai_mai_n1037_));
  NO2        m1015(.A(mai_mai_n1037_), .B(mai_mai_n41_), .Y(mai_mai_n1038_));
  NO3        m1016(.A(mai_mai_n1038_), .B(mai_mai_n1035_), .C(mai_mai_n1032_), .Y(mai_mai_n1039_));
  OAI210     m1017(.A0(mai_mai_n1029_), .A1(i_4_), .B0(mai_mai_n1039_), .Y(mai_mai_n1040_));
  NO3        m1018(.A(mai_mai_n1040_), .B(mai_mai_n1019_), .C(mai_mai_n1017_), .Y(mai_mai_n1041_));
  NA4        m1019(.A(mai_mai_n1041_), .B(mai_mai_n1001_), .C(mai_mai_n948_), .D(mai_mai_n871_), .Y(mai4));
  INV        m1020(.A(mai_mai_n698_), .Y(mai_mai_n1045_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u0033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  NA2        u0034(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n57_));
  NA3        u0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n58_));
  NO2        u0036(.A(i_1_), .B(i_6_), .Y(men_men_n59_));
  NA2        u0037(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  OAI210     u0038(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n58_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_12_), .Y(men_men_n62_));
  NAi21      u0040(.An(i_2_), .B(i_7_), .Y(men_men_n63_));
  INV        u0041(.A(i_1_), .Y(men_men_n64_));
  NA2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NA3        u0043(.A(men_men_n65_), .B(men_men_n63_), .C(men_men_n31_), .Y(men_men_n66_));
  NA2        u0044(.A(i_1_), .B(i_10_), .Y(men_men_n67_));
  NO2        u0045(.A(men_men_n67_), .B(i_6_), .Y(men_men_n68_));
  NAi31      u0046(.An(men_men_n68_), .B(men_men_n66_), .C(men_men_n62_), .Y(men_men_n69_));
  NA2        u0047(.A(men_men_n51_), .B(i_2_), .Y(men_men_n70_));
  AOI210     u0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n71_));
  NA2        u0049(.A(i_1_), .B(i_6_), .Y(men_men_n72_));
  NO2        u0050(.A(men_men_n72_), .B(men_men_n25_), .Y(men_men_n73_));
  INV        u0051(.A(i_0_), .Y(men_men_n74_));
  NAi21      u0052(.An(i_5_), .B(i_10_), .Y(men_men_n75_));
  NA2        u0053(.A(i_5_), .B(i_9_), .Y(men_men_n76_));
  AOI210     u0054(.A0(men_men_n76_), .A1(men_men_n75_), .B0(men_men_n74_), .Y(men_men_n77_));
  NO2        u0055(.A(men_men_n77_), .B(men_men_n73_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n78_), .Y(men_men_n79_));
  OAI210     u0057(.A0(men_men_n79_), .A1(men_men_n69_), .B0(i_0_), .Y(men_men_n80_));
  NA2        u0058(.A(i_12_), .B(i_5_), .Y(men_men_n81_));
  NA2        u0059(.A(i_2_), .B(i_8_), .Y(men_men_n82_));
  NO2        u0060(.A(men_men_n82_), .B(men_men_n59_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_9_), .Y(men_men_n84_));
  NO2        u0062(.A(i_3_), .B(i_7_), .Y(men_men_n85_));
  NO3        u0063(.A(men_men_n85_), .B(men_men_n84_), .C(men_men_n64_), .Y(men_men_n86_));
  INV        u0064(.A(i_6_), .Y(men_men_n87_));
  NO2        u0065(.A(i_2_), .B(i_7_), .Y(men_men_n88_));
  INV        u0066(.A(men_men_n88_), .Y(men_men_n89_));
  OAI210     u0067(.A0(men_men_n86_), .A1(men_men_n83_), .B0(men_men_n89_), .Y(men_men_n90_));
  NAi21      u0068(.An(i_6_), .B(i_10_), .Y(men_men_n91_));
  NA2        u0069(.A(i_6_), .B(i_9_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n64_), .Y(men_men_n93_));
  NA2        u0071(.A(i_2_), .B(i_6_), .Y(men_men_n94_));
  NO3        u0072(.A(men_men_n94_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n95_));
  NO2        u0073(.A(men_men_n95_), .B(men_men_n93_), .Y(men_men_n96_));
  AOI210     u0074(.A0(men_men_n96_), .A1(men_men_n90_), .B0(men_men_n81_), .Y(men_men_n97_));
  AN3        u0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n98_));
  NAi21      u0076(.An(i_6_), .B(i_11_), .Y(men_men_n99_));
  NO2        u0077(.A(i_5_), .B(i_8_), .Y(men_men_n100_));
  NOi21      u0078(.An(men_men_n100_), .B(men_men_n99_), .Y(men_men_n101_));
  AOI220     u0079(.A0(men_men_n101_), .A1(men_men_n63_), .B0(men_men_n98_), .B1(men_men_n32_), .Y(men_men_n102_));
  INV        u0080(.A(i_7_), .Y(men_men_n103_));
  NA2        u0081(.A(men_men_n47_), .B(men_men_n103_), .Y(men_men_n104_));
  NO2        u0082(.A(i_0_), .B(i_5_), .Y(men_men_n105_));
  NO2        u0083(.A(men_men_n105_), .B(men_men_n87_), .Y(men_men_n106_));
  NA2        u0084(.A(i_12_), .B(i_3_), .Y(men_men_n107_));
  INV        u0085(.A(men_men_n107_), .Y(men_men_n108_));
  NA3        u0086(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n104_), .Y(men_men_n109_));
  NAi21      u0087(.An(i_7_), .B(i_11_), .Y(men_men_n110_));
  AN2        u0088(.A(i_2_), .B(i_10_), .Y(men_men_n111_));
  NO2        u0089(.A(men_men_n111_), .B(i_7_), .Y(men_men_n112_));
  OR2        u0090(.A(men_men_n81_), .B(men_men_n59_), .Y(men_men_n113_));
  NO2        u0091(.A(i_8_), .B(men_men_n103_), .Y(men_men_n114_));
  NO3        u0092(.A(men_men_n114_), .B(men_men_n113_), .C(men_men_n112_), .Y(men_men_n115_));
  NA2        u0093(.A(i_12_), .B(i_7_), .Y(men_men_n116_));
  NO2        u0094(.A(men_men_n64_), .B(men_men_n26_), .Y(men_men_n117_));
  NA2        u0095(.A(men_men_n117_), .B(i_0_), .Y(men_men_n118_));
  NA2        u0096(.A(i_11_), .B(i_12_), .Y(men_men_n119_));
  OAI210     u0097(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n119_), .Y(men_men_n120_));
  NO2        u0098(.A(men_men_n120_), .B(men_men_n115_), .Y(men_men_n121_));
  NA3        u0099(.A(men_men_n121_), .B(men_men_n109_), .C(men_men_n102_), .Y(men_men_n122_));
  NOi21      u0100(.An(i_1_), .B(i_5_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n123_), .B(i_11_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n125_));
  NA2        u0103(.A(i_7_), .B(men_men_n25_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n126_), .B(men_men_n125_), .Y(men_men_n127_));
  NO2        u0105(.A(men_men_n127_), .B(men_men_n47_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n129_));
  NAi21      u0107(.An(i_3_), .B(i_8_), .Y(men_men_n130_));
  NA2        u0108(.A(men_men_n130_), .B(men_men_n63_), .Y(men_men_n131_));
  NOi31      u0109(.An(men_men_n131_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n132_));
  NO2        u0110(.A(i_1_), .B(men_men_n87_), .Y(men_men_n133_));
  NO2        u0111(.A(i_6_), .B(i_5_), .Y(men_men_n134_));
  NA2        u0112(.A(men_men_n134_), .B(i_3_), .Y(men_men_n135_));
  AO210      u0113(.A0(men_men_n135_), .A1(men_men_n48_), .B0(men_men_n133_), .Y(men_men_n136_));
  OAI220     u0114(.A0(men_men_n136_), .A1(men_men_n110_), .B0(men_men_n132_), .B1(men_men_n124_), .Y(men_men_n137_));
  NO3        u0115(.A(men_men_n137_), .B(men_men_n122_), .C(men_men_n97_), .Y(men_men_n138_));
  NA3        u0116(.A(men_men_n138_), .B(men_men_n80_), .C(men_men_n57_), .Y(men2));
  NO2        u0117(.A(men_men_n64_), .B(men_men_n37_), .Y(men_men_n140_));
  NA2        u0118(.A(i_6_), .B(men_men_n25_), .Y(men_men_n141_));
  NA2        u0119(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n142_));
  NA4        u0120(.A(men_men_n142_), .B(men_men_n78_), .C(men_men_n70_), .D(men_men_n30_), .Y(men0));
  AN2        u0121(.A(i_8_), .B(i_7_), .Y(men_men_n144_));
  NA2        u0122(.A(men_men_n144_), .B(i_6_), .Y(men_men_n145_));
  NO2        u0123(.A(i_12_), .B(i_13_), .Y(men_men_n146_));
  NAi21      u0124(.An(i_5_), .B(i_11_), .Y(men_men_n147_));
  NOi21      u0125(.An(men_men_n146_), .B(men_men_n147_), .Y(men_men_n148_));
  NO2        u0126(.A(i_0_), .B(i_1_), .Y(men_men_n149_));
  NA2        u0127(.A(i_2_), .B(i_3_), .Y(men_men_n150_));
  NO2        u0128(.A(men_men_n150_), .B(i_4_), .Y(men_men_n151_));
  NA3        u0129(.A(men_men_n151_), .B(men_men_n149_), .C(men_men_n148_), .Y(men_men_n152_));
  AN2        u0130(.A(men_men_n146_), .B(men_men_n84_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n153_), .B(men_men_n27_), .Y(men_men_n154_));
  NA2        u0132(.A(i_1_), .B(i_5_), .Y(men_men_n155_));
  NO2        u0133(.A(men_men_n74_), .B(men_men_n47_), .Y(men_men_n156_));
  NA2        u0134(.A(men_men_n156_), .B(men_men_n36_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n155_), .C(men_men_n154_), .Y(men_men_n158_));
  OR2        u0136(.A(i_0_), .B(i_1_), .Y(men_men_n159_));
  NO3        u0137(.A(men_men_n159_), .B(men_men_n81_), .C(i_13_), .Y(men_men_n160_));
  NAi32      u0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n161_));
  NAi21      u0139(.An(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  NOi21      u0140(.An(i_4_), .B(i_10_), .Y(men_men_n163_));
  NA2        u0141(.A(men_men_n163_), .B(men_men_n40_), .Y(men_men_n164_));
  NO2        u0142(.A(i_3_), .B(i_5_), .Y(men_men_n165_));
  NO3        u0143(.A(men_men_n74_), .B(i_2_), .C(i_1_), .Y(men_men_n166_));
  NA2        u0144(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  OAI210     u0145(.A0(men_men_n167_), .A1(men_men_n164_), .B0(men_men_n162_), .Y(men_men_n168_));
  NO2        u0146(.A(men_men_n168_), .B(men_men_n158_), .Y(men_men_n169_));
  AOI210     u0147(.A0(men_men_n169_), .A1(men_men_n152_), .B0(men_men_n145_), .Y(men_men_n170_));
  NA3        u0148(.A(men_men_n74_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n171_));
  NA2        u0149(.A(i_3_), .B(men_men_n49_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_4_), .B(i_9_), .Y(men_men_n173_));
  NOi21      u0151(.An(i_11_), .B(i_13_), .Y(men_men_n174_));
  NA2        u0152(.A(men_men_n174_), .B(men_men_n173_), .Y(men_men_n175_));
  OR2        u0153(.A(men_men_n175_), .B(men_men_n172_), .Y(men_men_n176_));
  NO2        u0154(.A(i_4_), .B(i_5_), .Y(men_men_n177_));
  NAi21      u0155(.An(i_12_), .B(i_11_), .Y(men_men_n178_));
  NO2        u0156(.A(men_men_n178_), .B(i_13_), .Y(men_men_n179_));
  NA3        u0157(.A(men_men_n179_), .B(men_men_n177_), .C(men_men_n84_), .Y(men_men_n180_));
  AOI210     u0158(.A0(men_men_n180_), .A1(men_men_n176_), .B0(men_men_n171_), .Y(men_men_n181_));
  NO2        u0159(.A(men_men_n74_), .B(men_men_n64_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n36_), .B(i_5_), .Y(men_men_n183_));
  NA2        u0161(.A(i_3_), .B(i_5_), .Y(men_men_n184_));
  NO2        u0162(.A(men_men_n74_), .B(i_5_), .Y(men_men_n185_));
  NO2        u0163(.A(i_13_), .B(i_10_), .Y(men_men_n186_));
  NA3        u0164(.A(men_men_n186_), .B(men_men_n185_), .C(men_men_n45_), .Y(men_men_n187_));
  NO2        u0165(.A(i_2_), .B(i_1_), .Y(men_men_n188_));
  NA2        u0166(.A(men_men_n188_), .B(i_3_), .Y(men_men_n189_));
  NAi21      u0167(.An(i_4_), .B(i_12_), .Y(men_men_n190_));
  NO4        u0168(.A(men_men_n190_), .B(men_men_n189_), .C(men_men_n187_), .D(men_men_n25_), .Y(men_men_n191_));
  NO2        u0169(.A(men_men_n191_), .B(men_men_n181_), .Y(men_men_n192_));
  INV        u0170(.A(i_8_), .Y(men_men_n193_));
  NO2        u0171(.A(men_men_n193_), .B(i_7_), .Y(men_men_n194_));
  NA2        u0172(.A(men_men_n194_), .B(i_6_), .Y(men_men_n195_));
  NO3        u0173(.A(i_3_), .B(men_men_n87_), .C(men_men_n49_), .Y(men_men_n196_));
  NA2        u0174(.A(men_men_n196_), .B(men_men_n114_), .Y(men_men_n197_));
  NO3        u0175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n198_));
  NA3        u0176(.A(men_men_n198_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n199_));
  NO3        u0177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n200_));
  OAI210     u0178(.A0(men_men_n98_), .A1(i_12_), .B0(men_men_n200_), .Y(men_men_n201_));
  AOI210     u0179(.A0(men_men_n201_), .A1(men_men_n199_), .B0(men_men_n197_), .Y(men_men_n202_));
  NO2        u0180(.A(i_3_), .B(i_8_), .Y(men_men_n203_));
  NO3        u0181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n204_));
  NA3        u0182(.A(men_men_n204_), .B(men_men_n203_), .C(men_men_n40_), .Y(men_men_n205_));
  NO2        u0183(.A(men_men_n105_), .B(men_men_n59_), .Y(men_men_n206_));
  INV        u0184(.A(men_men_n206_), .Y(men_men_n207_));
  NO2        u0185(.A(i_13_), .B(i_9_), .Y(men_men_n208_));
  NA3        u0186(.A(men_men_n208_), .B(i_6_), .C(men_men_n193_), .Y(men_men_n209_));
  NAi21      u0187(.An(i_12_), .B(i_3_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n45_), .B(i_5_), .Y(men_men_n211_));
  NO3        u0189(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n212_));
  NA3        u0190(.A(men_men_n212_), .B(men_men_n211_), .C(i_10_), .Y(men_men_n213_));
  OAI220     u0191(.A0(men_men_n213_), .A1(men_men_n209_), .B0(men_men_n207_), .B1(men_men_n205_), .Y(men_men_n214_));
  AOI210     u0192(.A0(men_men_n214_), .A1(i_7_), .B0(men_men_n202_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(i_4_), .B0(men_men_n195_), .B1(men_men_n192_), .Y(men_men_n216_));
  NAi21      u0194(.An(i_12_), .B(i_7_), .Y(men_men_n217_));
  NA3        u0195(.A(i_13_), .B(men_men_n193_), .C(i_10_), .Y(men_men_n218_));
  NA2        u0196(.A(i_0_), .B(i_5_), .Y(men_men_n219_));
  NAi31      u0197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n220_));
  NO2        u0198(.A(men_men_n36_), .B(i_13_), .Y(men_men_n221_));
  NO2        u0199(.A(men_men_n74_), .B(men_men_n26_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n47_), .B(men_men_n64_), .Y(men_men_n223_));
  NA3        u0201(.A(men_men_n223_), .B(men_men_n222_), .C(men_men_n221_), .Y(men_men_n224_));
  INV        u0202(.A(i_13_), .Y(men_men_n225_));
  NO2        u0203(.A(i_12_), .B(men_men_n225_), .Y(men_men_n226_));
  NA3        u0204(.A(men_men_n226_), .B(men_men_n198_), .C(men_men_n196_), .Y(men_men_n227_));
  OAI210     u0205(.A0(men_men_n224_), .A1(men_men_n220_), .B0(men_men_n227_), .Y(men_men_n228_));
  NA2        u0206(.A(men_men_n228_), .B(men_men_n144_), .Y(men_men_n229_));
  NO2        u0207(.A(i_12_), .B(men_men_n37_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n184_), .B(i_4_), .Y(men_men_n231_));
  NA2        u0209(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  OR2        u0210(.A(i_8_), .B(i_7_), .Y(men_men_n233_));
  NO2        u0211(.A(men_men_n233_), .B(men_men_n87_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n54_), .B(i_1_), .Y(men_men_n235_));
  INV        u0213(.A(i_12_), .Y(men_men_n236_));
  NO2        u0214(.A(men_men_n45_), .B(men_men_n236_), .Y(men_men_n237_));
  NO3        u0215(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n238_));
  NA2        u0216(.A(i_2_), .B(i_1_), .Y(men_men_n239_));
  NO3        u0217(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n240_));
  NAi21      u0218(.An(i_4_), .B(i_3_), .Y(men_men_n241_));
  NO2        u0219(.A(i_0_), .B(i_6_), .Y(men_men_n242_));
  NOi41      u0220(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n243_));
  NA2        u0221(.A(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n239_), .B(men_men_n184_), .Y(men_men_n245_));
  NAi21      u0223(.An(men_men_n244_), .B(men_men_n245_), .Y(men_men_n246_));
  INV        u0224(.A(men_men_n246_), .Y(men_men_n247_));
  NA2        u0225(.A(men_men_n247_), .B(men_men_n40_), .Y(men_men_n248_));
  NO2        u0226(.A(i_11_), .B(men_men_n225_), .Y(men_men_n249_));
  NOi21      u0227(.An(i_1_), .B(i_6_), .Y(men_men_n250_));
  NAi21      u0228(.An(i_3_), .B(i_7_), .Y(men_men_n251_));
  NA2        u0229(.A(men_men_n236_), .B(i_9_), .Y(men_men_n252_));
  OR4        u0230(.A(men_men_n252_), .B(men_men_n251_), .C(men_men_n250_), .D(men_men_n185_), .Y(men_men_n253_));
  NO2        u0231(.A(i_12_), .B(i_3_), .Y(men_men_n254_));
  NA2        u0232(.A(men_men_n74_), .B(i_5_), .Y(men_men_n255_));
  NA2        u0233(.A(i_3_), .B(i_9_), .Y(men_men_n256_));
  NAi21      u0234(.An(i_7_), .B(i_10_), .Y(men_men_n257_));
  NO2        u0235(.A(men_men_n257_), .B(men_men_n256_), .Y(men_men_n258_));
  NA3        u0236(.A(men_men_n258_), .B(men_men_n255_), .C(men_men_n65_), .Y(men_men_n259_));
  NA2        u0237(.A(men_men_n259_), .B(men_men_n253_), .Y(men_men_n260_));
  NA3        u0238(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n261_));
  INV        u0239(.A(men_men_n145_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n236_), .B(i_13_), .Y(men_men_n263_));
  NO2        u0241(.A(men_men_n263_), .B(men_men_n76_), .Y(men_men_n264_));
  AOI220     u0242(.A0(men_men_n264_), .A1(men_men_n262_), .B0(men_men_n260_), .B1(men_men_n249_), .Y(men_men_n265_));
  NA2        u0243(.A(i_12_), .B(i_6_), .Y(men_men_n266_));
  OR2        u0244(.A(i_13_), .B(i_9_), .Y(men_men_n267_));
  NO2        u0245(.A(men_men_n241_), .B(i_2_), .Y(men_men_n268_));
  NA2        u0246(.A(men_men_n249_), .B(i_9_), .Y(men_men_n269_));
  NO3        u0247(.A(i_11_), .B(men_men_n225_), .C(men_men_n25_), .Y(men_men_n270_));
  NO2        u0248(.A(men_men_n251_), .B(i_8_), .Y(men_men_n271_));
  NO2        u0249(.A(i_6_), .B(men_men_n49_), .Y(men_men_n272_));
  NA3        u0250(.A(men_men_n265_), .B(men_men_n248_), .C(men_men_n229_), .Y(men_men_n273_));
  NO3        u0251(.A(i_12_), .B(men_men_n225_), .C(men_men_n37_), .Y(men_men_n274_));
  INV        u0252(.A(men_men_n274_), .Y(men_men_n275_));
  NO3        u0253(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n276_));
  NO3        u0254(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n239_), .B(i_0_), .Y(men_men_n278_));
  AOI220     u0256(.A0(men_men_n278_), .A1(men_men_n194_), .B0(men_men_n277_), .B1(men_men_n144_), .Y(men_men_n279_));
  NA2        u0257(.A(men_men_n272_), .B(men_men_n26_), .Y(men_men_n280_));
  NO2        u0258(.A(men_men_n280_), .B(men_men_n279_), .Y(men_men_n281_));
  NA2        u0259(.A(i_0_), .B(i_1_), .Y(men_men_n282_));
  NO2        u0260(.A(men_men_n282_), .B(i_2_), .Y(men_men_n283_));
  NO2        u0261(.A(men_men_n60_), .B(i_6_), .Y(men_men_n284_));
  NA3        u0262(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n165_), .Y(men_men_n285_));
  OAI210     u0263(.A0(men_men_n167_), .A1(men_men_n145_), .B0(men_men_n285_), .Y(men_men_n286_));
  NO2        u0264(.A(men_men_n286_), .B(men_men_n281_), .Y(men_men_n287_));
  NO2        u0265(.A(i_3_), .B(i_10_), .Y(men_men_n288_));
  NA3        u0266(.A(men_men_n288_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n289_));
  NO2        u0267(.A(i_2_), .B(men_men_n103_), .Y(men_men_n290_));
  NA2        u0268(.A(i_1_), .B(men_men_n36_), .Y(men_men_n291_));
  NO2        u0269(.A(men_men_n291_), .B(i_8_), .Y(men_men_n292_));
  NA2        u0270(.A(men_men_n292_), .B(men_men_n290_), .Y(men_men_n293_));
  AN2        u0271(.A(i_3_), .B(i_10_), .Y(men_men_n294_));
  NA4        u0272(.A(men_men_n294_), .B(men_men_n198_), .C(men_men_n179_), .D(men_men_n177_), .Y(men_men_n295_));
  NO2        u0273(.A(i_5_), .B(men_men_n37_), .Y(men_men_n296_));
  NO2        u0274(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n297_));
  OR2        u0275(.A(men_men_n293_), .B(men_men_n289_), .Y(men_men_n298_));
  OAI220     u0276(.A0(men_men_n298_), .A1(i_6_), .B0(men_men_n287_), .B1(men_men_n275_), .Y(men_men_n299_));
  NO4        u0277(.A(men_men_n299_), .B(men_men_n273_), .C(men_men_n216_), .D(men_men_n170_), .Y(men_men_n300_));
  NO3        u0278(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n301_));
  NO2        u0279(.A(men_men_n60_), .B(men_men_n87_), .Y(men_men_n302_));
  NA2        u0280(.A(men_men_n278_), .B(men_men_n302_), .Y(men_men_n303_));
  NO3        u0281(.A(i_6_), .B(men_men_n193_), .C(i_7_), .Y(men_men_n304_));
  NA2        u0282(.A(men_men_n304_), .B(men_men_n198_), .Y(men_men_n305_));
  AOI210     u0283(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n172_), .Y(men_men_n306_));
  NO2        u0284(.A(i_2_), .B(i_3_), .Y(men_men_n307_));
  OR2        u0285(.A(i_0_), .B(i_5_), .Y(men_men_n308_));
  NA2        u0286(.A(men_men_n219_), .B(men_men_n308_), .Y(men_men_n309_));
  NAi21      u0287(.An(i_8_), .B(i_7_), .Y(men_men_n310_));
  NO2        u0288(.A(men_men_n310_), .B(i_6_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n159_), .B(men_men_n47_), .Y(men_men_n312_));
  NA3        u0290(.A(men_men_n312_), .B(men_men_n311_), .C(men_men_n165_), .Y(men_men_n313_));
  INV        u0291(.A(men_men_n313_), .Y(men_men_n314_));
  OAI210     u0292(.A0(men_men_n314_), .A1(men_men_n306_), .B0(i_4_), .Y(men_men_n315_));
  NO2        u0293(.A(i_12_), .B(i_10_), .Y(men_men_n316_));
  NOi21      u0294(.An(i_5_), .B(i_0_), .Y(men_men_n317_));
  AOI210     u0295(.A0(i_2_), .A1(men_men_n49_), .B0(men_men_n103_), .Y(men_men_n318_));
  NO4        u0296(.A(men_men_n318_), .B(men_men_n291_), .C(men_men_n317_), .D(men_men_n130_), .Y(men_men_n319_));
  NA4        u0297(.A(men_men_n85_), .B(men_men_n36_), .C(men_men_n87_), .D(i_8_), .Y(men_men_n320_));
  NA2        u0298(.A(men_men_n319_), .B(men_men_n316_), .Y(men_men_n321_));
  NO2        u0299(.A(i_6_), .B(i_8_), .Y(men_men_n322_));
  NOi21      u0300(.An(i_0_), .B(i_2_), .Y(men_men_n323_));
  AN2        u0301(.A(men_men_n323_), .B(men_men_n322_), .Y(men_men_n324_));
  NO2        u0302(.A(i_1_), .B(i_7_), .Y(men_men_n325_));
  AO220      u0303(.A0(men_men_n325_), .A1(men_men_n324_), .B0(men_men_n311_), .B1(men_men_n235_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n326_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n327_));
  NA3        u0305(.A(men_men_n327_), .B(men_men_n321_), .C(men_men_n315_), .Y(men_men_n328_));
  NA3        u0306(.A(men_men_n250_), .B(men_men_n290_), .C(men_men_n193_), .Y(men_men_n329_));
  NO2        u0307(.A(men_men_n329_), .B(men_men_n309_), .Y(men_men_n330_));
  NOi21      u0308(.An(men_men_n155_), .B(men_men_n106_), .Y(men_men_n331_));
  NO2        u0309(.A(men_men_n331_), .B(men_men_n126_), .Y(men_men_n332_));
  OAI210     u0310(.A0(men_men_n332_), .A1(men_men_n330_), .B0(i_3_), .Y(men_men_n333_));
  INV        u0311(.A(men_men_n85_), .Y(men_men_n334_));
  NO2        u0312(.A(men_men_n282_), .B(men_men_n82_), .Y(men_men_n335_));
  NA2        u0313(.A(men_men_n335_), .B(men_men_n134_), .Y(men_men_n336_));
  NO2        u0314(.A(men_men_n94_), .B(men_men_n193_), .Y(men_men_n337_));
  NA3        u0315(.A(men_men_n219_), .B(men_men_n337_), .C(men_men_n64_), .Y(men_men_n338_));
  AOI210     u0316(.A0(men_men_n338_), .A1(men_men_n336_), .B0(men_men_n334_), .Y(men_men_n339_));
  NO2        u0317(.A(men_men_n193_), .B(i_9_), .Y(men_men_n340_));
  NA2        u0318(.A(men_men_n340_), .B(men_men_n206_), .Y(men_men_n341_));
  NO2        u0319(.A(men_men_n341_), .B(men_men_n47_), .Y(men_men_n342_));
  NO3        u0320(.A(men_men_n342_), .B(men_men_n339_), .C(men_men_n281_), .Y(men_men_n343_));
  AOI210     u0321(.A0(men_men_n343_), .A1(men_men_n333_), .B0(men_men_n164_), .Y(men_men_n344_));
  AOI210     u0322(.A0(men_men_n328_), .A1(men_men_n301_), .B0(men_men_n344_), .Y(men_men_n345_));
  NOi32      u0323(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n346_));
  INV        u0324(.A(men_men_n346_), .Y(men_men_n347_));
  NAi21      u0325(.An(i_0_), .B(i_6_), .Y(men_men_n348_));
  NAi21      u0326(.An(i_1_), .B(i_5_), .Y(men_men_n349_));
  NA2        u0327(.A(men_men_n349_), .B(men_men_n348_), .Y(men_men_n350_));
  NA2        u0328(.A(men_men_n350_), .B(men_men_n25_), .Y(men_men_n351_));
  OAI210     u0329(.A0(men_men_n351_), .A1(men_men_n161_), .B0(men_men_n244_), .Y(men_men_n352_));
  NAi41      u0330(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n353_));
  OAI220     u0331(.A0(men_men_n353_), .A1(men_men_n349_), .B0(men_men_n220_), .B1(men_men_n161_), .Y(men_men_n354_));
  AOI210     u0332(.A0(men_men_n353_), .A1(men_men_n161_), .B0(men_men_n159_), .Y(men_men_n355_));
  NOi32      u0333(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n356_));
  NAi21      u0334(.An(i_6_), .B(i_1_), .Y(men_men_n357_));
  NA3        u0335(.A(men_men_n357_), .B(men_men_n356_), .C(men_men_n47_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n358_), .B(i_0_), .Y(men_men_n359_));
  OR3        u0337(.A(men_men_n359_), .B(men_men_n355_), .C(men_men_n354_), .Y(men_men_n360_));
  NO2        u0338(.A(i_1_), .B(men_men_n103_), .Y(men_men_n361_));
  NAi21      u0339(.An(i_3_), .B(i_4_), .Y(men_men_n362_));
  NO2        u0340(.A(men_men_n362_), .B(i_9_), .Y(men_men_n363_));
  AN2        u0341(.A(i_6_), .B(i_7_), .Y(men_men_n364_));
  OAI210     u0342(.A0(men_men_n364_), .A1(men_men_n361_), .B0(men_men_n363_), .Y(men_men_n365_));
  NA2        u0343(.A(i_2_), .B(i_7_), .Y(men_men_n366_));
  NO2        u0344(.A(men_men_n362_), .B(i_10_), .Y(men_men_n367_));
  NA3        u0345(.A(men_men_n367_), .B(men_men_n366_), .C(men_men_n242_), .Y(men_men_n368_));
  AOI210     u0346(.A0(men_men_n368_), .A1(men_men_n365_), .B0(men_men_n185_), .Y(men_men_n369_));
  AOI210     u0347(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n370_));
  OAI210     u0348(.A0(men_men_n370_), .A1(men_men_n188_), .B0(men_men_n367_), .Y(men_men_n371_));
  AOI220     u0349(.A0(men_men_n367_), .A1(men_men_n325_), .B0(men_men_n238_), .B1(men_men_n188_), .Y(men_men_n372_));
  AOI210     u0350(.A0(men_men_n372_), .A1(men_men_n371_), .B0(i_5_), .Y(men_men_n373_));
  NO4        u0351(.A(men_men_n373_), .B(men_men_n369_), .C(men_men_n360_), .D(men_men_n352_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n374_), .B(men_men_n347_), .Y(men_men_n375_));
  NO2        u0353(.A(men_men_n60_), .B(men_men_n25_), .Y(men_men_n376_));
  AN2        u0354(.A(i_12_), .B(i_5_), .Y(men_men_n377_));
  NO2        u0355(.A(i_4_), .B(men_men_n26_), .Y(men_men_n378_));
  NA2        u0356(.A(men_men_n378_), .B(men_men_n377_), .Y(men_men_n379_));
  NO2        u0357(.A(i_11_), .B(i_6_), .Y(men_men_n380_));
  NA3        u0358(.A(men_men_n380_), .B(men_men_n312_), .C(men_men_n225_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n381_), .B(men_men_n379_), .Y(men_men_n382_));
  NO2        u0360(.A(men_men_n241_), .B(i_5_), .Y(men_men_n383_));
  NO2        u0361(.A(i_5_), .B(i_10_), .Y(men_men_n384_));
  AOI220     u0362(.A0(men_men_n384_), .A1(men_men_n268_), .B0(men_men_n383_), .B1(men_men_n198_), .Y(men_men_n385_));
  NA2        u0363(.A(men_men_n146_), .B(men_men_n46_), .Y(men_men_n386_));
  NO2        u0364(.A(men_men_n386_), .B(men_men_n385_), .Y(men_men_n387_));
  OAI210     u0365(.A0(men_men_n387_), .A1(men_men_n382_), .B0(men_men_n376_), .Y(men_men_n388_));
  NO2        u0366(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n389_));
  NO2        u0367(.A(men_men_n152_), .B(men_men_n87_), .Y(men_men_n390_));
  OAI210     u0368(.A0(men_men_n390_), .A1(men_men_n382_), .B0(men_men_n389_), .Y(men_men_n391_));
  NO3        u0369(.A(men_men_n87_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n392_));
  NO2        u0370(.A(i_3_), .B(men_men_n103_), .Y(men_men_n393_));
  NO2        u0371(.A(i_11_), .B(i_12_), .Y(men_men_n394_));
  NA2        u0372(.A(men_men_n384_), .B(men_men_n236_), .Y(men_men_n395_));
  NA3        u0373(.A(men_men_n114_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n396_));
  OAI220     u0374(.A0(men_men_n396_), .A1(men_men_n220_), .B0(men_men_n395_), .B1(men_men_n320_), .Y(men_men_n397_));
  NAi21      u0375(.An(i_13_), .B(i_0_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n398_), .B(men_men_n239_), .Y(men_men_n399_));
  NA2        u0377(.A(men_men_n397_), .B(men_men_n399_), .Y(men_men_n400_));
  NA3        u0378(.A(men_men_n400_), .B(men_men_n391_), .C(men_men_n388_), .Y(men_men_n401_));
  NA2        u0379(.A(men_men_n45_), .B(men_men_n225_), .Y(men_men_n402_));
  NO3        u0380(.A(i_1_), .B(i_12_), .C(men_men_n87_), .Y(men_men_n403_));
  NO2        u0381(.A(i_0_), .B(i_11_), .Y(men_men_n404_));
  INV        u0382(.A(i_5_), .Y(men_men_n405_));
  AN2        u0383(.A(i_1_), .B(i_6_), .Y(men_men_n406_));
  NOi21      u0384(.An(i_2_), .B(i_12_), .Y(men_men_n407_));
  NA2        u0385(.A(men_men_n407_), .B(men_men_n406_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n408_), .B(men_men_n405_), .Y(men_men_n409_));
  NA2        u0387(.A(men_men_n144_), .B(i_9_), .Y(men_men_n410_));
  NO2        u0388(.A(men_men_n410_), .B(i_4_), .Y(men_men_n411_));
  NA2        u0389(.A(men_men_n409_), .B(men_men_n411_), .Y(men_men_n412_));
  NAi21      u0390(.An(i_9_), .B(i_4_), .Y(men_men_n413_));
  OR2        u0391(.A(i_13_), .B(i_10_), .Y(men_men_n414_));
  NO3        u0392(.A(men_men_n414_), .B(men_men_n119_), .C(men_men_n413_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n175_), .B(men_men_n125_), .Y(men_men_n416_));
  OR2        u0394(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n417_));
  NO2        u0395(.A(men_men_n103_), .B(men_men_n25_), .Y(men_men_n418_));
  NA2        u0396(.A(men_men_n274_), .B(men_men_n418_), .Y(men_men_n419_));
  NA2        u0397(.A(men_men_n272_), .B(men_men_n212_), .Y(men_men_n420_));
  OAI220     u0398(.A0(men_men_n420_), .A1(men_men_n417_), .B0(men_men_n419_), .B1(men_men_n331_), .Y(men_men_n421_));
  INV        u0399(.A(men_men_n421_), .Y(men_men_n422_));
  AOI210     u0400(.A0(men_men_n422_), .A1(men_men_n412_), .B0(men_men_n26_), .Y(men_men_n423_));
  AOI220     u0401(.A0(men_men_n284_), .A1(men_men_n276_), .B0(men_men_n278_), .B1(men_men_n302_), .Y(men_men_n424_));
  NO2        u0402(.A(men_men_n424_), .B(men_men_n172_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n184_), .B(men_men_n87_), .Y(men_men_n426_));
  INV        u0404(.A(men_men_n425_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n196_), .B(men_men_n98_), .Y(men_men_n428_));
  NA3        u0406(.A(men_men_n312_), .B(men_men_n165_), .C(men_men_n87_), .Y(men_men_n429_));
  AOI210     u0407(.A0(men_men_n429_), .A1(men_men_n428_), .B0(men_men_n310_), .Y(men_men_n430_));
  NA2        u0408(.A(men_men_n193_), .B(i_10_), .Y(men_men_n431_));
  NA3        u0409(.A(men_men_n255_), .B(men_men_n65_), .C(i_2_), .Y(men_men_n432_));
  NO2        u0410(.A(men_men_n432_), .B(men_men_n431_), .Y(men_men_n433_));
  NO2        u0411(.A(i_3_), .B(men_men_n49_), .Y(men_men_n434_));
  NA3        u0412(.A(men_men_n325_), .B(men_men_n324_), .C(men_men_n434_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n304_), .B(men_men_n309_), .Y(men_men_n436_));
  OAI210     u0414(.A0(men_men_n436_), .A1(men_men_n189_), .B0(men_men_n435_), .Y(men_men_n437_));
  NO3        u0415(.A(men_men_n437_), .B(men_men_n433_), .C(men_men_n430_), .Y(men_men_n438_));
  AOI210     u0416(.A0(men_men_n438_), .A1(men_men_n427_), .B0(men_men_n269_), .Y(men_men_n439_));
  NO4        u0417(.A(men_men_n439_), .B(men_men_n423_), .C(men_men_n401_), .D(men_men_n375_), .Y(men_men_n440_));
  NO2        u0418(.A(men_men_n64_), .B(i_4_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n74_), .B(i_13_), .Y(men_men_n442_));
  NO2        u0420(.A(i_10_), .B(i_9_), .Y(men_men_n443_));
  NAi21      u0421(.An(i_12_), .B(i_8_), .Y(men_men_n444_));
  NO2        u0422(.A(men_men_n444_), .B(i_3_), .Y(men_men_n445_));
  NO2        u0423(.A(men_men_n47_), .B(i_4_), .Y(men_men_n446_));
  NA2        u0424(.A(men_men_n446_), .B(men_men_n106_), .Y(men_men_n447_));
  NO2        u0425(.A(men_men_n447_), .B(men_men_n205_), .Y(men_men_n448_));
  NA2        u0426(.A(men_men_n297_), .B(i_0_), .Y(men_men_n449_));
  NO3        u0427(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n450_));
  NA2        u0428(.A(men_men_n266_), .B(men_men_n99_), .Y(men_men_n451_));
  NA2        u0429(.A(men_men_n451_), .B(men_men_n450_), .Y(men_men_n452_));
  NA2        u0430(.A(i_8_), .B(i_9_), .Y(men_men_n453_));
  AOI210     u0431(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n454_));
  OR2        u0432(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n274_), .B(men_men_n206_), .Y(men_men_n456_));
  OAI220     u0434(.A0(men_men_n456_), .A1(men_men_n455_), .B0(men_men_n452_), .B1(men_men_n449_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n249_), .B(men_men_n296_), .Y(men_men_n458_));
  NO3        u0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n459_));
  INV        u0437(.A(men_men_n459_), .Y(men_men_n460_));
  NA3        u0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n461_));
  NA4        u0439(.A(men_men_n147_), .B(men_men_n117_), .C(men_men_n81_), .D(men_men_n23_), .Y(men_men_n462_));
  OAI220     u0440(.A0(men_men_n462_), .A1(men_men_n461_), .B0(men_men_n460_), .B1(men_men_n458_), .Y(men_men_n463_));
  NO3        u0441(.A(men_men_n463_), .B(men_men_n457_), .C(men_men_n448_), .Y(men_men_n464_));
  NA2        u0442(.A(men_men_n283_), .B(men_men_n110_), .Y(men_men_n465_));
  OR2        u0443(.A(men_men_n465_), .B(men_men_n209_), .Y(men_men_n466_));
  OA210      u0444(.A0(men_men_n341_), .A1(men_men_n103_), .B0(men_men_n285_), .Y(men_men_n467_));
  OA220      u0445(.A0(men_men_n467_), .A1(men_men_n164_), .B0(men_men_n466_), .B1(men_men_n232_), .Y(men_men_n468_));
  NA2        u0446(.A(men_men_n98_), .B(i_13_), .Y(men_men_n469_));
  NA2        u0447(.A(men_men_n426_), .B(men_men_n376_), .Y(men_men_n470_));
  NO2        u0448(.A(i_2_), .B(i_13_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n470_), .B(men_men_n469_), .Y(men_men_n472_));
  NO3        u0450(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n473_));
  NO2        u0451(.A(i_6_), .B(i_7_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n474_), .B(men_men_n473_), .Y(men_men_n475_));
  NO2        u0453(.A(i_11_), .B(i_1_), .Y(men_men_n476_));
  NO2        u0454(.A(men_men_n74_), .B(i_3_), .Y(men_men_n477_));
  OR2        u0455(.A(i_11_), .B(i_8_), .Y(men_men_n478_));
  NOi21      u0456(.An(i_2_), .B(i_7_), .Y(men_men_n479_));
  NAi31      u0457(.An(men_men_n478_), .B(men_men_n479_), .C(men_men_n477_), .Y(men_men_n480_));
  NO2        u0458(.A(men_men_n414_), .B(i_6_), .Y(men_men_n481_));
  NA3        u0459(.A(men_men_n481_), .B(men_men_n441_), .C(men_men_n76_), .Y(men_men_n482_));
  NO2        u0460(.A(men_men_n482_), .B(men_men_n480_), .Y(men_men_n483_));
  NO2        u0461(.A(i_3_), .B(men_men_n193_), .Y(men_men_n484_));
  NO2        u0462(.A(i_6_), .B(i_10_), .Y(men_men_n485_));
  NA4        u0463(.A(men_men_n485_), .B(men_men_n301_), .C(men_men_n484_), .D(men_men_n236_), .Y(men_men_n486_));
  NO2        u0464(.A(men_men_n486_), .B(men_men_n157_), .Y(men_men_n487_));
  NA3        u0465(.A(men_men_n243_), .B(men_men_n174_), .C(men_men_n134_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n489_));
  NO2        u0467(.A(men_men_n159_), .B(i_3_), .Y(men_men_n490_));
  NAi31      u0468(.An(men_men_n489_), .B(men_men_n490_), .C(men_men_n226_), .Y(men_men_n491_));
  NA3        u0469(.A(men_men_n389_), .B(men_men_n182_), .C(men_men_n151_), .Y(men_men_n492_));
  NA3        u0470(.A(men_men_n492_), .B(men_men_n491_), .C(men_men_n488_), .Y(men_men_n493_));
  NO4        u0471(.A(men_men_n493_), .B(men_men_n487_), .C(men_men_n483_), .D(men_men_n472_), .Y(men_men_n494_));
  NA2        u0472(.A(men_men_n450_), .B(men_men_n377_), .Y(men_men_n495_));
  NA2        u0473(.A(men_men_n459_), .B(men_men_n384_), .Y(men_men_n496_));
  NO2        u0474(.A(men_men_n496_), .B(men_men_n224_), .Y(men_men_n497_));
  NAi21      u0475(.An(men_men_n218_), .B(men_men_n394_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n325_), .B(men_men_n219_), .Y(men_men_n499_));
  NO2        u0477(.A(men_men_n26_), .B(i_5_), .Y(men_men_n500_));
  NO2        u0478(.A(men_men_n499_), .B(men_men_n498_), .Y(men_men_n501_));
  NA2        u0479(.A(men_men_n27_), .B(i_10_), .Y(men_men_n502_));
  NA2        u0480(.A(men_men_n301_), .B(men_men_n238_), .Y(men_men_n503_));
  OAI220     u0481(.A0(men_men_n503_), .A1(men_men_n432_), .B0(men_men_n502_), .B1(men_men_n469_), .Y(men_men_n504_));
  NA4        u0482(.A(men_men_n294_), .B(men_men_n223_), .C(men_men_n74_), .D(men_men_n236_), .Y(men_men_n505_));
  NO2        u0483(.A(men_men_n505_), .B(men_men_n475_), .Y(men_men_n506_));
  NO4        u0484(.A(men_men_n506_), .B(men_men_n504_), .C(men_men_n501_), .D(men_men_n497_), .Y(men_men_n507_));
  NA4        u0485(.A(men_men_n507_), .B(men_men_n494_), .C(men_men_n468_), .D(men_men_n464_), .Y(men_men_n508_));
  NA3        u0486(.A(men_men_n294_), .B(men_men_n179_), .C(men_men_n177_), .Y(men_men_n509_));
  OAI210     u0487(.A0(men_men_n289_), .A1(men_men_n183_), .B0(men_men_n509_), .Y(men_men_n510_));
  AN2        u0488(.A(men_men_n276_), .B(men_men_n234_), .Y(men_men_n511_));
  NA2        u0489(.A(men_men_n511_), .B(men_men_n510_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n124_), .B(men_men_n113_), .Y(men_men_n513_));
  AN2        u0491(.A(men_men_n513_), .B(men_men_n450_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n301_), .B(men_men_n166_), .Y(men_men_n515_));
  OAI210     u0493(.A0(men_men_n515_), .A1(men_men_n232_), .B0(men_men_n295_), .Y(men_men_n516_));
  AOI220     u0494(.A0(men_men_n516_), .A1(men_men_n311_), .B0(men_men_n514_), .B1(men_men_n297_), .Y(men_men_n517_));
  NA2        u0495(.A(men_men_n377_), .B(men_men_n225_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n346_), .B(men_men_n74_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n364_), .B(men_men_n356_), .Y(men_men_n520_));
  OR2        u0498(.A(men_men_n518_), .B(men_men_n520_), .Y(men_men_n521_));
  NO2        u0499(.A(men_men_n36_), .B(i_8_), .Y(men_men_n522_));
  NAi41      u0500(.An(men_men_n519_), .B(men_men_n485_), .C(men_men_n522_), .D(men_men_n47_), .Y(men_men_n523_));
  AOI210     u0501(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n415_), .Y(men_men_n524_));
  NA3        u0502(.A(men_men_n524_), .B(men_men_n523_), .C(men_men_n521_), .Y(men_men_n525_));
  INV        u0503(.A(men_men_n525_), .Y(men_men_n526_));
  NA2        u0504(.A(men_men_n255_), .B(men_men_n65_), .Y(men_men_n527_));
  OAI210     u0505(.A0(i_8_), .A1(men_men_n527_), .B0(men_men_n136_), .Y(men_men_n528_));
  NO2        u0506(.A(i_7_), .B(men_men_n199_), .Y(men_men_n529_));
  OR2        u0507(.A(men_men_n184_), .B(i_4_), .Y(men_men_n530_));
  NO2        u0508(.A(men_men_n530_), .B(men_men_n87_), .Y(men_men_n531_));
  AOI220     u0509(.A0(men_men_n531_), .A1(men_men_n529_), .B0(men_men_n528_), .B1(men_men_n416_), .Y(men_men_n532_));
  NA4        u0510(.A(men_men_n532_), .B(men_men_n526_), .C(men_men_n517_), .D(men_men_n512_), .Y(men_men_n533_));
  NA2        u0511(.A(men_men_n383_), .B(men_men_n283_), .Y(men_men_n534_));
  OAI210     u0512(.A0(men_men_n379_), .A1(men_men_n171_), .B0(men_men_n534_), .Y(men_men_n535_));
  NO2        u0513(.A(i_12_), .B(men_men_n193_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n536_), .B(men_men_n225_), .Y(men_men_n537_));
  NO3        u0515(.A(men_men_n1058_), .B(men_men_n537_), .C(men_men_n465_), .Y(men_men_n538_));
  NOi31      u0516(.An(men_men_n304_), .B(men_men_n414_), .C(men_men_n38_), .Y(men_men_n539_));
  OAI210     u0517(.A0(men_men_n539_), .A1(men_men_n538_), .B0(men_men_n535_), .Y(men_men_n540_));
  NO2        u0518(.A(i_8_), .B(i_7_), .Y(men_men_n541_));
  AOI220     u0519(.A0(men_men_n312_), .A1(men_men_n40_), .B0(men_men_n235_), .B1(men_men_n208_), .Y(men_men_n542_));
  NO2        u0520(.A(men_men_n542_), .B(men_men_n530_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n45_), .B(i_10_), .Y(men_men_n544_));
  NO2        u0522(.A(men_men_n544_), .B(i_6_), .Y(men_men_n545_));
  NA3        u0523(.A(men_men_n545_), .B(men_men_n543_), .C(men_men_n541_), .Y(men_men_n546_));
  NOi31      u0524(.An(men_men_n278_), .B(men_men_n289_), .C(men_men_n183_), .Y(men_men_n547_));
  NA3        u0525(.A(men_men_n294_), .B(men_men_n177_), .C(men_men_n98_), .Y(men_men_n548_));
  NO2        u0526(.A(men_men_n221_), .B(men_men_n45_), .Y(men_men_n549_));
  NO2        u0527(.A(men_men_n159_), .B(i_5_), .Y(men_men_n550_));
  NA3        u0528(.A(men_men_n550_), .B(men_men_n402_), .C(men_men_n307_), .Y(men_men_n551_));
  OAI210     u0529(.A0(men_men_n551_), .A1(men_men_n549_), .B0(men_men_n548_), .Y(men_men_n552_));
  OAI210     u0530(.A0(men_men_n552_), .A1(men_men_n547_), .B0(men_men_n459_), .Y(men_men_n553_));
  NA3        u0531(.A(men_men_n553_), .B(men_men_n546_), .C(men_men_n540_), .Y(men_men_n554_));
  NA3        u0532(.A(men_men_n219_), .B(men_men_n72_), .C(men_men_n45_), .Y(men_men_n555_));
  NA2        u0533(.A(men_men_n274_), .B(men_men_n85_), .Y(men_men_n556_));
  AOI210     u0534(.A0(men_men_n555_), .A1(men_men_n336_), .B0(men_men_n556_), .Y(men_men_n557_));
  NA2        u0535(.A(men_men_n284_), .B(men_men_n276_), .Y(men_men_n558_));
  NO2        u0536(.A(men_men_n558_), .B(men_men_n176_), .Y(men_men_n559_));
  NA2        u0537(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n560_));
  NA2        u0538(.A(men_men_n443_), .B(men_men_n221_), .Y(men_men_n561_));
  NO2        u0539(.A(men_men_n560_), .B(men_men_n561_), .Y(men_men_n562_));
  AOI210     u0540(.A0(men_men_n357_), .A1(men_men_n47_), .B0(men_men_n361_), .Y(men_men_n563_));
  NA2        u0541(.A(i_0_), .B(men_men_n49_), .Y(men_men_n564_));
  NA3        u0542(.A(men_men_n536_), .B(men_men_n270_), .C(men_men_n564_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n563_), .B(men_men_n565_), .Y(men_men_n566_));
  NO4        u0544(.A(men_men_n566_), .B(men_men_n562_), .C(men_men_n559_), .D(men_men_n557_), .Y(men_men_n567_));
  NO4        u0545(.A(men_men_n250_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n568_));
  NO3        u0546(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n569_));
  NO2        u0547(.A(men_men_n233_), .B(men_men_n36_), .Y(men_men_n570_));
  AN2        u0548(.A(men_men_n570_), .B(men_men_n569_), .Y(men_men_n571_));
  OA210      u0549(.A0(men_men_n571_), .A1(men_men_n568_), .B0(men_men_n346_), .Y(men_men_n572_));
  NO2        u0550(.A(men_men_n414_), .B(i_1_), .Y(men_men_n573_));
  NOi31      u0551(.An(men_men_n573_), .B(men_men_n451_), .C(men_men_n74_), .Y(men_men_n574_));
  AN4        u0552(.A(men_men_n574_), .B(men_men_n411_), .C(men_men_n500_), .D(i_2_), .Y(men_men_n575_));
  NO2        u0553(.A(men_men_n424_), .B(men_men_n180_), .Y(men_men_n576_));
  NO3        u0554(.A(men_men_n576_), .B(men_men_n575_), .C(men_men_n572_), .Y(men_men_n577_));
  NOi21      u0555(.An(i_10_), .B(i_6_), .Y(men_men_n578_));
  NO2        u0556(.A(men_men_n87_), .B(men_men_n25_), .Y(men_men_n579_));
  AOI220     u0557(.A0(men_men_n274_), .A1(men_men_n579_), .B0(men_men_n270_), .B1(men_men_n578_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n580_), .B(men_men_n449_), .Y(men_men_n581_));
  NO2        u0559(.A(men_men_n116_), .B(men_men_n23_), .Y(men_men_n582_));
  NOi31      u0560(.An(men_men_n148_), .B(i_10_), .C(men_men_n320_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n583_), .B(men_men_n581_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n519_), .B(men_men_n372_), .Y(men_men_n585_));
  INV        u0563(.A(men_men_n307_), .Y(men_men_n586_));
  NO2        u0564(.A(i_12_), .B(men_men_n87_), .Y(men_men_n587_));
  NA3        u0565(.A(men_men_n587_), .B(men_men_n270_), .C(men_men_n564_), .Y(men_men_n588_));
  NA3        u0566(.A(men_men_n380_), .B(men_men_n274_), .C(men_men_n219_), .Y(men_men_n589_));
  AOI210     u0567(.A0(men_men_n589_), .A1(men_men_n588_), .B0(men_men_n586_), .Y(men_men_n590_));
  OR2        u0568(.A(i_2_), .B(i_5_), .Y(men_men_n591_));
  OR2        u0569(.A(men_men_n591_), .B(men_men_n406_), .Y(men_men_n592_));
  AOI210     u0570(.A0(men_men_n366_), .A1(men_men_n242_), .B0(men_men_n198_), .Y(men_men_n593_));
  AOI210     u0571(.A0(men_men_n593_), .A1(men_men_n592_), .B0(men_men_n498_), .Y(men_men_n594_));
  NO3        u0572(.A(men_men_n594_), .B(men_men_n590_), .C(men_men_n585_), .Y(men_men_n595_));
  NA4        u0573(.A(men_men_n595_), .B(men_men_n584_), .C(men_men_n577_), .D(men_men_n567_), .Y(men_men_n596_));
  NO4        u0574(.A(men_men_n596_), .B(men_men_n554_), .C(men_men_n533_), .D(men_men_n508_), .Y(men_men_n597_));
  NA4        u0575(.A(men_men_n597_), .B(men_men_n440_), .C(men_men_n345_), .D(men_men_n300_), .Y(men7));
  NO2        u0576(.A(men_men_n94_), .B(men_men_n55_), .Y(men_men_n599_));
  NA2        u0577(.A(men_men_n485_), .B(men_men_n85_), .Y(men_men_n600_));
  NA2        u0578(.A(i_11_), .B(men_men_n193_), .Y(men_men_n601_));
  NA3        u0579(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n236_), .B(i_4_), .Y(men_men_n603_));
  NA2        u0581(.A(men_men_n603_), .B(i_8_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n107_), .B(men_men_n602_), .Y(men_men_n605_));
  NA2        u0583(.A(i_2_), .B(men_men_n87_), .Y(men_men_n606_));
  OAI210     u0584(.A0(men_men_n88_), .A1(men_men_n203_), .B0(men_men_n204_), .Y(men_men_n607_));
  NO2        u0585(.A(i_7_), .B(men_men_n37_), .Y(men_men_n608_));
  NA2        u0586(.A(i_4_), .B(i_8_), .Y(men_men_n609_));
  AOI210     u0587(.A0(men_men_n609_), .A1(men_men_n294_), .B0(men_men_n608_), .Y(men_men_n610_));
  OAI220     u0588(.A0(men_men_n610_), .A1(men_men_n606_), .B0(men_men_n607_), .B1(i_13_), .Y(men_men_n611_));
  NO3        u0589(.A(men_men_n611_), .B(men_men_n605_), .C(men_men_n599_), .Y(men_men_n612_));
  AOI210     u0590(.A0(men_men_n130_), .A1(men_men_n63_), .B0(i_10_), .Y(men_men_n613_));
  AOI210     u0591(.A0(men_men_n613_), .A1(men_men_n236_), .B0(men_men_n163_), .Y(men_men_n614_));
  OR2        u0592(.A(i_6_), .B(i_10_), .Y(men_men_n615_));
  NO2        u0593(.A(men_men_n615_), .B(men_men_n23_), .Y(men_men_n616_));
  OR3        u0594(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n617_));
  NO3        u0595(.A(men_men_n617_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n618_));
  INV        u0596(.A(men_men_n200_), .Y(men_men_n619_));
  NO2        u0597(.A(men_men_n618_), .B(men_men_n616_), .Y(men_men_n620_));
  OA220      u0598(.A0(men_men_n620_), .A1(men_men_n586_), .B0(men_men_n614_), .B1(men_men_n267_), .Y(men_men_n621_));
  AOI210     u0599(.A0(men_men_n621_), .A1(men_men_n612_), .B0(men_men_n64_), .Y(men_men_n622_));
  NOi21      u0600(.An(i_11_), .B(i_7_), .Y(men_men_n623_));
  AO210      u0601(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n624_));
  NO2        u0602(.A(men_men_n624_), .B(men_men_n623_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n625_), .B(men_men_n208_), .Y(men_men_n626_));
  NA3        u0604(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n627_));
  NAi31      u0605(.An(men_men_n627_), .B(men_men_n217_), .C(i_11_), .Y(men_men_n628_));
  AOI210     u0606(.A0(men_men_n628_), .A1(men_men_n626_), .B0(men_men_n64_), .Y(men_men_n629_));
  OR2        u0607(.A(men_men_n372_), .B(men_men_n41_), .Y(men_men_n630_));
  NO3        u0608(.A(men_men_n257_), .B(men_men_n210_), .C(men_men_n601_), .Y(men_men_n631_));
  OAI210     u0609(.A0(men_men_n631_), .A1(men_men_n226_), .B0(men_men_n64_), .Y(men_men_n632_));
  NA2        u0610(.A(men_men_n407_), .B(men_men_n31_), .Y(men_men_n633_));
  OR2        u0611(.A(men_men_n210_), .B(men_men_n110_), .Y(men_men_n634_));
  NA2        u0612(.A(men_men_n634_), .B(men_men_n633_), .Y(men_men_n635_));
  NO2        u0613(.A(men_men_n64_), .B(i_9_), .Y(men_men_n636_));
  NO2        u0614(.A(men_men_n636_), .B(i_4_), .Y(men_men_n637_));
  NA2        u0615(.A(men_men_n637_), .B(men_men_n635_), .Y(men_men_n638_));
  NO2        u0616(.A(i_1_), .B(i_12_), .Y(men_men_n639_));
  NA3        u0617(.A(men_men_n639_), .B(men_men_n111_), .C(men_men_n24_), .Y(men_men_n640_));
  BUFFER     u0618(.A(men_men_n640_), .Y(men_men_n641_));
  NA4        u0619(.A(men_men_n641_), .B(men_men_n638_), .C(men_men_n632_), .D(men_men_n630_), .Y(men_men_n642_));
  OAI210     u0620(.A0(men_men_n642_), .A1(men_men_n629_), .B0(i_6_), .Y(men_men_n643_));
  NO2        u0621(.A(men_men_n627_), .B(men_men_n110_), .Y(men_men_n644_));
  NA2        u0622(.A(men_men_n644_), .B(men_men_n587_), .Y(men_men_n645_));
  NO2        u0623(.A(men_men_n236_), .B(men_men_n87_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n646_), .B(i_11_), .Y(men_men_n647_));
  NA2        u0625(.A(men_men_n645_), .B(men_men_n452_), .Y(men_men_n648_));
  NO4        u0626(.A(men_men_n217_), .B(men_men_n130_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n649_));
  NA2        u0627(.A(men_men_n649_), .B(men_men_n636_), .Y(men_men_n650_));
  NA2        u0628(.A(men_men_n236_), .B(i_6_), .Y(men_men_n651_));
  NO3        u0629(.A(men_men_n615_), .B(men_men_n233_), .C(men_men_n23_), .Y(men_men_n652_));
  AOI210     u0630(.A0(i_1_), .A1(men_men_n258_), .B0(men_men_n652_), .Y(men_men_n653_));
  OAI210     u0631(.A0(men_men_n653_), .A1(men_men_n45_), .B0(men_men_n650_), .Y(men_men_n654_));
  NA3        u0632(.A(men_men_n541_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n655_));
  INV        u0633(.A(i_2_), .Y(men_men_n656_));
  NA2        u0634(.A(men_men_n140_), .B(i_9_), .Y(men_men_n657_));
  NA3        u0635(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n47_), .B(i_1_), .Y(men_men_n659_));
  NA3        u0637(.A(men_men_n659_), .B(men_men_n266_), .C(men_men_n45_), .Y(men_men_n660_));
  OAI220     u0638(.A0(men_men_n660_), .A1(men_men_n658_), .B0(men_men_n657_), .B1(men_men_n656_), .Y(men_men_n661_));
  AOI210     u0639(.A0(men_men_n476_), .A1(men_men_n418_), .B0(men_men_n240_), .Y(men_men_n662_));
  NO2        u0640(.A(men_men_n662_), .B(men_men_n606_), .Y(men_men_n663_));
  NAi21      u0641(.An(men_men_n655_), .B(men_men_n93_), .Y(men_men_n664_));
  NO2        u0642(.A(i_11_), .B(men_men_n37_), .Y(men_men_n665_));
  INV        u0643(.A(men_men_n664_), .Y(men_men_n666_));
  OR3        u0644(.A(men_men_n666_), .B(men_men_n663_), .C(men_men_n661_), .Y(men_men_n667_));
  NO3        u0645(.A(men_men_n667_), .B(men_men_n654_), .C(men_men_n648_), .Y(men_men_n668_));
  NO2        u0646(.A(men_men_n236_), .B(men_men_n103_), .Y(men_men_n669_));
  NO2        u0647(.A(men_men_n669_), .B(men_men_n623_), .Y(men_men_n670_));
  NA2        u0648(.A(men_men_n670_), .B(i_1_), .Y(men_men_n671_));
  NO2        u0649(.A(men_men_n671_), .B(men_men_n617_), .Y(men_men_n672_));
  NO2        u0650(.A(men_men_n413_), .B(men_men_n87_), .Y(men_men_n673_));
  NA2        u0651(.A(men_men_n672_), .B(men_men_n47_), .Y(men_men_n674_));
  NA2        u0652(.A(i_3_), .B(men_men_n193_), .Y(men_men_n675_));
  NO2        u0653(.A(men_men_n675_), .B(men_men_n116_), .Y(men_men_n676_));
  AN2        u0654(.A(men_men_n676_), .B(men_men_n545_), .Y(men_men_n677_));
  NO2        u0655(.A(men_men_n233_), .B(men_men_n45_), .Y(men_men_n678_));
  NO3        u0656(.A(men_men_n678_), .B(men_men_n297_), .C(men_men_n237_), .Y(men_men_n679_));
  NO2        u0657(.A(men_men_n119_), .B(men_men_n37_), .Y(men_men_n680_));
  NO2        u0658(.A(men_men_n680_), .B(i_6_), .Y(men_men_n681_));
  NO2        u0659(.A(men_men_n87_), .B(i_9_), .Y(men_men_n682_));
  NO2        u0660(.A(men_men_n682_), .B(men_men_n64_), .Y(men_men_n683_));
  NO2        u0661(.A(men_men_n683_), .B(men_men_n639_), .Y(men_men_n684_));
  NO4        u0662(.A(men_men_n684_), .B(men_men_n681_), .C(men_men_n679_), .D(i_4_), .Y(men_men_n685_));
  NA2        u0663(.A(i_1_), .B(i_3_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n453_), .B(men_men_n94_), .Y(men_men_n687_));
  AOI210     u0665(.A0(men_men_n678_), .A1(men_men_n578_), .B0(men_men_n687_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n688_), .B(men_men_n686_), .Y(men_men_n689_));
  NO3        u0667(.A(men_men_n689_), .B(men_men_n685_), .C(men_men_n677_), .Y(men_men_n690_));
  NA4        u0668(.A(men_men_n690_), .B(men_men_n674_), .C(men_men_n668_), .D(men_men_n643_), .Y(men_men_n691_));
  NO3        u0669(.A(men_men_n478_), .B(i_3_), .C(i_7_), .Y(men_men_n692_));
  NOi21      u0670(.An(men_men_n692_), .B(i_10_), .Y(men_men_n693_));
  OA210      u0671(.A0(men_men_n693_), .A1(men_men_n243_), .B0(men_men_n87_), .Y(men_men_n694_));
  NA2        u0672(.A(men_men_n364_), .B(men_men_n363_), .Y(men_men_n695_));
  NA3        u0673(.A(men_men_n485_), .B(men_men_n522_), .C(men_men_n47_), .Y(men_men_n696_));
  NO3        u0674(.A(men_men_n479_), .B(men_men_n609_), .C(men_men_n87_), .Y(men_men_n697_));
  NA2        u0675(.A(men_men_n697_), .B(men_men_n25_), .Y(men_men_n698_));
  NA3        u0676(.A(men_men_n163_), .B(men_men_n85_), .C(men_men_n87_), .Y(men_men_n699_));
  NA4        u0677(.A(men_men_n699_), .B(men_men_n698_), .C(men_men_n696_), .D(men_men_n695_), .Y(men_men_n700_));
  OAI210     u0678(.A0(men_men_n700_), .A1(men_men_n694_), .B0(i_1_), .Y(men_men_n701_));
  AOI210     u0679(.A0(men_men_n266_), .A1(men_men_n99_), .B0(i_1_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n362_), .B(i_2_), .Y(men_men_n703_));
  NA2        u0681(.A(men_men_n703_), .B(men_men_n702_), .Y(men_men_n704_));
  AOI210     u0682(.A0(men_men_n704_), .A1(men_men_n701_), .B0(i_13_), .Y(men_men_n705_));
  OR2        u0683(.A(i_11_), .B(i_7_), .Y(men_men_n706_));
  NA3        u0684(.A(men_men_n706_), .B(men_men_n108_), .C(men_men_n140_), .Y(men_men_n707_));
  AOI220     u0685(.A0(men_men_n471_), .A1(men_men_n163_), .B0(men_men_n446_), .B1(men_men_n140_), .Y(men_men_n708_));
  OAI210     u0686(.A0(men_men_n708_), .A1(men_men_n45_), .B0(men_men_n707_), .Y(men_men_n709_));
  AOI210     u0687(.A0(men_men_n658_), .A1(men_men_n55_), .B0(i_12_), .Y(men_men_n710_));
  NO2        u0688(.A(men_men_n479_), .B(men_men_n24_), .Y(men_men_n711_));
  AOI220     u0689(.A0(men_men_n711_), .A1(men_men_n673_), .B0(men_men_n243_), .B1(men_men_n133_), .Y(men_men_n712_));
  OAI220     u0690(.A0(men_men_n712_), .A1(men_men_n41_), .B0(men_men_n1057_), .B1(men_men_n94_), .Y(men_men_n713_));
  AOI210     u0691(.A0(men_men_n709_), .A1(men_men_n322_), .B0(men_men_n713_), .Y(men_men_n714_));
  NA2        u0692(.A(men_men_n380_), .B(men_men_n659_), .Y(men_men_n715_));
  NO2        u0693(.A(men_men_n715_), .B(men_men_n241_), .Y(men_men_n716_));
  AOI210     u0694(.A0(men_men_n444_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n717_));
  NOi31      u0695(.An(men_men_n717_), .B(men_men_n600_), .C(men_men_n45_), .Y(men_men_n718_));
  NA2        u0696(.A(men_men_n129_), .B(i_13_), .Y(men_men_n719_));
  NO2        u0697(.A(men_men_n658_), .B(men_men_n116_), .Y(men_men_n720_));
  INV        u0698(.A(men_men_n720_), .Y(men_men_n721_));
  OAI220     u0699(.A0(men_men_n721_), .A1(men_men_n72_), .B0(men_men_n719_), .B1(men_men_n702_), .Y(men_men_n722_));
  NA2        u0700(.A(men_men_n26_), .B(men_men_n193_), .Y(men_men_n723_));
  NA2        u0701(.A(men_men_n723_), .B(i_7_), .Y(men_men_n724_));
  NO3        u0702(.A(men_men_n479_), .B(men_men_n236_), .C(men_men_n87_), .Y(men_men_n725_));
  NA2        u0703(.A(men_men_n725_), .B(men_men_n724_), .Y(men_men_n726_));
  AOI220     u0704(.A0(men_men_n380_), .A1(men_men_n659_), .B0(men_men_n93_), .B1(men_men_n104_), .Y(men_men_n727_));
  OAI220     u0705(.A0(men_men_n727_), .A1(men_men_n604_), .B0(men_men_n726_), .B1(men_men_n619_), .Y(men_men_n728_));
  NO4        u0706(.A(men_men_n728_), .B(men_men_n722_), .C(men_men_n718_), .D(men_men_n716_), .Y(men_men_n729_));
  OR2        u0707(.A(i_11_), .B(i_6_), .Y(men_men_n730_));
  NA3        u0708(.A(men_men_n603_), .B(men_men_n723_), .C(i_7_), .Y(men_men_n731_));
  AOI210     u0709(.A0(men_men_n731_), .A1(men_men_n721_), .B0(men_men_n730_), .Y(men_men_n732_));
  NA3        u0710(.A(men_men_n407_), .B(men_men_n608_), .C(men_men_n99_), .Y(men_men_n733_));
  NA2        u0711(.A(men_men_n647_), .B(i_13_), .Y(men_men_n734_));
  NA2        u0712(.A(men_men_n104_), .B(men_men_n723_), .Y(men_men_n735_));
  NAi21      u0713(.An(i_11_), .B(i_12_), .Y(men_men_n736_));
  NOi41      u0714(.An(men_men_n112_), .B(men_men_n736_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n737_));
  NO3        u0715(.A(men_men_n479_), .B(men_men_n587_), .C(men_men_n609_), .Y(men_men_n738_));
  AOI220     u0716(.A0(men_men_n738_), .A1(men_men_n301_), .B0(men_men_n737_), .B1(men_men_n735_), .Y(men_men_n739_));
  NA3        u0717(.A(men_men_n739_), .B(men_men_n734_), .C(men_men_n733_), .Y(men_men_n740_));
  OAI210     u0718(.A0(men_men_n740_), .A1(men_men_n732_), .B0(men_men_n64_), .Y(men_men_n741_));
  NO2        u0719(.A(i_2_), .B(i_12_), .Y(men_men_n742_));
  NA2        u0720(.A(men_men_n361_), .B(men_men_n742_), .Y(men_men_n743_));
  NA2        u0721(.A(i_8_), .B(men_men_n25_), .Y(men_men_n744_));
  NO3        u0722(.A(men_men_n744_), .B(men_men_n378_), .C(men_men_n603_), .Y(men_men_n745_));
  OAI210     u0723(.A0(men_men_n745_), .A1(men_men_n363_), .B0(men_men_n361_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n130_), .B(i_2_), .Y(men_men_n747_));
  NA2        u0725(.A(men_men_n746_), .B(men_men_n743_), .Y(men_men_n748_));
  NA3        u0726(.A(men_men_n748_), .B(men_men_n46_), .C(men_men_n225_), .Y(men_men_n749_));
  NA4        u0727(.A(men_men_n749_), .B(men_men_n741_), .C(men_men_n729_), .D(men_men_n714_), .Y(men_men_n750_));
  OR4        u0728(.A(men_men_n750_), .B(men_men_n705_), .C(men_men_n691_), .D(men_men_n622_), .Y(men5));
  NA2        u0729(.A(men_men_n670_), .B(men_men_n268_), .Y(men_men_n752_));
  AN2        u0730(.A(men_men_n24_), .B(i_10_), .Y(men_men_n753_));
  NA3        u0731(.A(men_men_n753_), .B(men_men_n742_), .C(men_men_n110_), .Y(men_men_n754_));
  NO2        u0732(.A(men_men_n604_), .B(i_11_), .Y(men_men_n755_));
  NA2        u0733(.A(men_men_n88_), .B(men_men_n755_), .Y(men_men_n756_));
  NA3        u0734(.A(men_men_n756_), .B(men_men_n754_), .C(men_men_n752_), .Y(men_men_n757_));
  NO3        u0735(.A(i_11_), .B(men_men_n236_), .C(i_13_), .Y(men_men_n758_));
  NO2        u0736(.A(men_men_n126_), .B(men_men_n23_), .Y(men_men_n759_));
  NA2        u0737(.A(i_12_), .B(i_8_), .Y(men_men_n760_));
  OAI210     u0738(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n760_), .Y(men_men_n761_));
  INV        u0739(.A(men_men_n443_), .Y(men_men_n762_));
  AOI220     u0740(.A0(men_men_n307_), .A1(men_men_n582_), .B0(men_men_n761_), .B1(men_men_n759_), .Y(men_men_n763_));
  INV        u0741(.A(men_men_n763_), .Y(men_men_n764_));
  NO2        u0742(.A(men_men_n764_), .B(men_men_n757_), .Y(men_men_n765_));
  INV        u0743(.A(men_men_n174_), .Y(men_men_n766_));
  INV        u0744(.A(men_men_n243_), .Y(men_men_n767_));
  OAI210     u0745(.A0(men_men_n703_), .A1(men_men_n445_), .B0(men_men_n112_), .Y(men_men_n768_));
  AOI210     u0746(.A0(men_men_n768_), .A1(men_men_n767_), .B0(men_men_n766_), .Y(men_men_n769_));
  NO2        u0747(.A(men_men_n453_), .B(men_men_n26_), .Y(men_men_n770_));
  NO2        u0748(.A(men_men_n770_), .B(men_men_n418_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n771_), .B(i_2_), .Y(men_men_n772_));
  INV        u0750(.A(men_men_n772_), .Y(men_men_n773_));
  AOI210     u0751(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n414_), .Y(men_men_n774_));
  AOI210     u0752(.A0(men_men_n774_), .A1(men_men_n773_), .B0(men_men_n769_), .Y(men_men_n775_));
  NO2        u0753(.A(men_men_n190_), .B(men_men_n127_), .Y(men_men_n776_));
  OAI210     u0754(.A0(men_men_n776_), .A1(men_men_n759_), .B0(i_2_), .Y(men_men_n777_));
  INV        u0755(.A(men_men_n175_), .Y(men_men_n778_));
  NO3        u0756(.A(men_men_n624_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n779_));
  AOI210     u0757(.A0(men_men_n778_), .A1(men_men_n88_), .B0(men_men_n779_), .Y(men_men_n780_));
  AOI210     u0758(.A0(men_men_n780_), .A1(men_men_n777_), .B0(men_men_n193_), .Y(men_men_n781_));
  OA210      u0759(.A0(men_men_n625_), .A1(men_men_n128_), .B0(i_13_), .Y(men_men_n782_));
  NA2        u0760(.A(men_men_n200_), .B(men_men_n203_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n153_), .B(men_men_n601_), .Y(men_men_n784_));
  AOI210     u0762(.A0(men_men_n784_), .A1(men_men_n783_), .B0(men_men_n366_), .Y(men_men_n785_));
  AOI210     u0763(.A0(men_men_n210_), .A1(men_men_n150_), .B0(men_men_n522_), .Y(men_men_n786_));
  NA2        u0764(.A(men_men_n786_), .B(men_men_n418_), .Y(men_men_n787_));
  NO2        u0765(.A(men_men_n104_), .B(men_men_n45_), .Y(men_men_n788_));
  INV        u0766(.A(men_men_n290_), .Y(men_men_n789_));
  NA4        u0767(.A(men_men_n789_), .B(men_men_n294_), .C(men_men_n126_), .D(men_men_n43_), .Y(men_men_n790_));
  OAI210     u0768(.A0(men_men_n790_), .A1(men_men_n788_), .B0(men_men_n787_), .Y(men_men_n791_));
  NO4        u0769(.A(men_men_n791_), .B(men_men_n785_), .C(men_men_n782_), .D(men_men_n781_), .Y(men_men_n792_));
  NA2        u0770(.A(men_men_n582_), .B(men_men_n28_), .Y(men_men_n793_));
  NA2        u0771(.A(men_men_n758_), .B(men_men_n271_), .Y(men_men_n794_));
  NA2        u0772(.A(men_men_n794_), .B(men_men_n793_), .Y(men_men_n795_));
  NO2        u0773(.A(men_men_n63_), .B(i_12_), .Y(men_men_n796_));
  NO2        u0774(.A(men_men_n796_), .B(men_men_n128_), .Y(men_men_n797_));
  NO2        u0775(.A(men_men_n797_), .B(men_men_n601_), .Y(men_men_n798_));
  AOI220     u0776(.A0(men_men_n798_), .A1(men_men_n36_), .B0(men_men_n795_), .B1(men_men_n47_), .Y(men_men_n799_));
  NA4        u0777(.A(men_men_n799_), .B(men_men_n792_), .C(men_men_n775_), .D(men_men_n765_), .Y(men6));
  NA4        u0778(.A(men_men_n384_), .B(men_men_n484_), .C(men_men_n72_), .D(men_men_n103_), .Y(men_men_n801_));
  INV        u0779(.A(men_men_n801_), .Y(men_men_n802_));
  NO2        u0780(.A(men_men_n220_), .B(men_men_n489_), .Y(men_men_n803_));
  NO2        u0781(.A(i_11_), .B(i_9_), .Y(men_men_n804_));
  NO2        u0782(.A(men_men_n802_), .B(men_men_n317_), .Y(men_men_n805_));
  OR2        u0783(.A(men_men_n805_), .B(i_12_), .Y(men_men_n806_));
  NA2        u0784(.A(men_men_n367_), .B(men_men_n325_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n587_), .B(men_men_n64_), .Y(men_men_n808_));
  NA2        u0786(.A(men_men_n693_), .B(men_men_n72_), .Y(men_men_n809_));
  NA3        u0787(.A(men_men_n809_), .B(men_men_n808_), .C(men_men_n807_), .Y(men_men_n810_));
  INV        u0788(.A(men_men_n197_), .Y(men_men_n811_));
  AOI220     u0789(.A0(men_men_n811_), .A1(men_men_n804_), .B0(men_men_n810_), .B1(men_men_n74_), .Y(men_men_n812_));
  INV        u0790(.A(men_men_n316_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n76_), .B(men_men_n133_), .Y(men_men_n814_));
  INV        u0792(.A(men_men_n126_), .Y(men_men_n815_));
  NA2        u0793(.A(men_men_n815_), .B(men_men_n47_), .Y(men_men_n816_));
  AOI210     u0794(.A0(men_men_n816_), .A1(men_men_n814_), .B0(men_men_n813_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n250_), .B(i_9_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n818_), .B(men_men_n796_), .Y(men_men_n819_));
  AOI210     u0797(.A0(men_men_n819_), .A1(men_men_n520_), .B0(men_men_n185_), .Y(men_men_n820_));
  NO2        u0798(.A(men_men_n32_), .B(i_11_), .Y(men_men_n821_));
  NA3        u0799(.A(men_men_n821_), .B(men_men_n474_), .C(men_men_n384_), .Y(men_men_n822_));
  NAi32      u0800(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n823_));
  NO2        u0801(.A(men_men_n730_), .B(men_men_n823_), .Y(men_men_n824_));
  NAi21      u0802(.An(men_men_n824_), .B(men_men_n822_), .Y(men_men_n825_));
  OR3        u0803(.A(men_men_n825_), .B(men_men_n820_), .C(men_men_n817_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n706_), .B(i_2_), .Y(men_men_n827_));
  NA2        u0805(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n828_));
  NO2        u0806(.A(men_men_n828_), .B(men_men_n406_), .Y(men_men_n829_));
  NA2        u0807(.A(men_men_n829_), .B(men_men_n827_), .Y(men_men_n830_));
  AO220      u0808(.A0(men_men_n350_), .A1(men_men_n340_), .B0(men_men_n392_), .B1(men_men_n601_), .Y(men_men_n831_));
  NA3        u0809(.A(men_men_n831_), .B(men_men_n254_), .C(i_7_), .Y(men_men_n832_));
  BUFFER     u0810(.A(men_men_n625_), .Y(men_men_n833_));
  NA3        u0811(.A(men_men_n833_), .B(men_men_n149_), .C(men_men_n70_), .Y(men_men_n834_));
  AO210      u0812(.A0(men_men_n496_), .A1(men_men_n762_), .B0(men_men_n36_), .Y(men_men_n835_));
  NA4        u0813(.A(men_men_n835_), .B(men_men_n834_), .C(men_men_n832_), .D(men_men_n830_), .Y(men_men_n836_));
  NO2        u0814(.A(men_men_n646_), .B(i_11_), .Y(men_men_n837_));
  AOI220     u0815(.A0(men_men_n837_), .A1(men_men_n569_), .B0(men_men_n803_), .B1(men_men_n724_), .Y(men_men_n838_));
  NA3        u0816(.A(men_men_n366_), .B(men_men_n238_), .C(men_men_n149_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n392_), .B(men_men_n71_), .Y(men_men_n840_));
  NA4        u0818(.A(men_men_n840_), .B(men_men_n839_), .C(men_men_n838_), .D(men_men_n607_), .Y(men_men_n841_));
  AOI210     u0819(.A0(men_men_n445_), .A1(men_men_n443_), .B0(men_men_n568_), .Y(men_men_n842_));
  NO2        u0820(.A(men_men_n615_), .B(men_men_n104_), .Y(men_men_n843_));
  OAI210     u0821(.A0(men_men_n843_), .A1(men_men_n113_), .B0(men_men_n404_), .Y(men_men_n844_));
  NA2        u0822(.A(men_men_n242_), .B(men_men_n47_), .Y(men_men_n845_));
  INV        u0823(.A(men_men_n592_), .Y(men_men_n846_));
  NA3        u0824(.A(men_men_n846_), .B(men_men_n316_), .C(i_7_), .Y(men_men_n847_));
  NA3        u0825(.A(men_men_n847_), .B(men_men_n844_), .C(men_men_n842_), .Y(men_men_n848_));
  NO4        u0826(.A(men_men_n848_), .B(men_men_n841_), .C(men_men_n836_), .D(men_men_n826_), .Y(men_men_n849_));
  NA4        u0827(.A(men_men_n849_), .B(men_men_n812_), .C(men_men_n806_), .D(men_men_n374_), .Y(men3));
  NA2        u0828(.A(i_12_), .B(i_10_), .Y(men_men_n851_));
  NA2        u0829(.A(i_6_), .B(i_7_), .Y(men_men_n852_));
  NO2        u0830(.A(men_men_n852_), .B(i_0_), .Y(men_men_n853_));
  NO2        u0831(.A(i_11_), .B(men_men_n236_), .Y(men_men_n854_));
  NA3        u0832(.A(men_men_n839_), .B(men_men_n607_), .C(men_men_n365_), .Y(men_men_n855_));
  NA2        u0833(.A(men_men_n855_), .B(men_men_n40_), .Y(men_men_n856_));
  NOi21      u0834(.An(men_men_n98_), .B(men_men_n771_), .Y(men_men_n857_));
  NO3        u0835(.A(men_men_n634_), .B(men_men_n453_), .C(men_men_n133_), .Y(men_men_n858_));
  AN2        u0836(.A(men_men_n451_), .B(men_men_n56_), .Y(men_men_n859_));
  NO3        u0837(.A(men_men_n859_), .B(men_men_n858_), .C(men_men_n857_), .Y(men_men_n860_));
  AOI210     u0838(.A0(men_men_n860_), .A1(men_men_n856_), .B0(men_men_n49_), .Y(men_men_n861_));
  NO4        u0839(.A(men_men_n370_), .B(men_men_n377_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n862_));
  NA2        u0840(.A(men_men_n185_), .B(men_men_n578_), .Y(men_men_n863_));
  NOi21      u0841(.An(men_men_n863_), .B(men_men_n862_), .Y(men_men_n864_));
  NO2        u0842(.A(men_men_n864_), .B(men_men_n64_), .Y(men_men_n865_));
  NOi21      u0843(.An(i_5_), .B(i_9_), .Y(men_men_n866_));
  NA2        u0844(.A(men_men_n866_), .B(men_men_n442_), .Y(men_men_n867_));
  BUFFER     u0845(.A(men_men_n266_), .Y(men_men_n868_));
  AOI210     u0846(.A0(men_men_n868_), .A1(men_men_n476_), .B0(men_men_n697_), .Y(men_men_n869_));
  NO3        u0847(.A(men_men_n410_), .B(men_men_n266_), .C(men_men_n74_), .Y(men_men_n870_));
  NO2        u0848(.A(men_men_n178_), .B(men_men_n150_), .Y(men_men_n871_));
  AOI210     u0849(.A0(men_men_n871_), .A1(men_men_n242_), .B0(men_men_n870_), .Y(men_men_n872_));
  OAI220     u0850(.A0(men_men_n872_), .A1(men_men_n183_), .B0(men_men_n869_), .B1(men_men_n867_), .Y(men_men_n873_));
  NO3        u0851(.A(men_men_n873_), .B(men_men_n865_), .C(men_men_n861_), .Y(men_men_n874_));
  NA2        u0852(.A(men_men_n185_), .B(men_men_n24_), .Y(men_men_n875_));
  NA2        u0853(.A(men_men_n301_), .B(men_men_n131_), .Y(men_men_n876_));
  NAi21      u0854(.An(men_men_n164_), .B(men_men_n434_), .Y(men_men_n877_));
  OAI220     u0855(.A0(men_men_n877_), .A1(men_men_n845_), .B0(men_men_n876_), .B1(men_men_n395_), .Y(men_men_n878_));
  INV        u0856(.A(men_men_n878_), .Y(men_men_n879_));
  NO2        u0857(.A(men_men_n384_), .B(men_men_n282_), .Y(men_men_n880_));
  NA2        u0858(.A(men_men_n880_), .B(men_men_n720_), .Y(men_men_n881_));
  NA2        u0859(.A(men_men_n579_), .B(i_0_), .Y(men_men_n882_));
  NO3        u0860(.A(men_men_n882_), .B(men_men_n379_), .C(men_men_n88_), .Y(men_men_n883_));
  NO4        u0861(.A(men_men_n591_), .B(men_men_n217_), .C(men_men_n414_), .D(men_men_n406_), .Y(men_men_n884_));
  AOI210     u0862(.A0(men_men_n884_), .A1(i_11_), .B0(men_men_n883_), .Y(men_men_n885_));
  INV        u0863(.A(men_men_n474_), .Y(men_men_n886_));
  NA2        u0864(.A(men_men_n758_), .B(men_men_n317_), .Y(men_men_n887_));
  AOI210     u0865(.A0(men_men_n485_), .A1(men_men_n88_), .B0(men_men_n59_), .Y(men_men_n888_));
  NO2        u0866(.A(men_men_n888_), .B(men_men_n887_), .Y(men_men_n889_));
  NO2        u0867(.A(men_men_n252_), .B(men_men_n155_), .Y(men_men_n890_));
  NA2        u0868(.A(i_0_), .B(i_10_), .Y(men_men_n891_));
  INV        u0869(.A(men_men_n544_), .Y(men_men_n892_));
  NO4        u0870(.A(men_men_n116_), .B(men_men_n59_), .C(men_men_n675_), .D(i_5_), .Y(men_men_n893_));
  AO220      u0871(.A0(men_men_n893_), .A1(men_men_n892_), .B0(men_men_n890_), .B1(i_6_), .Y(men_men_n894_));
  AOI220     u0872(.A0(men_men_n323_), .A1(men_men_n100_), .B0(men_men_n185_), .B1(men_men_n85_), .Y(men_men_n895_));
  NA2        u0873(.A(men_men_n573_), .B(i_4_), .Y(men_men_n896_));
  NA2        u0874(.A(men_men_n188_), .B(men_men_n203_), .Y(men_men_n897_));
  OAI220     u0875(.A0(men_men_n897_), .A1(men_men_n887_), .B0(men_men_n896_), .B1(men_men_n895_), .Y(men_men_n898_));
  NO3        u0876(.A(men_men_n898_), .B(men_men_n894_), .C(men_men_n889_), .Y(men_men_n899_));
  NA4        u0877(.A(men_men_n899_), .B(men_men_n885_), .C(men_men_n881_), .D(men_men_n879_), .Y(men_men_n900_));
  NO2        u0878(.A(men_men_n105_), .B(men_men_n37_), .Y(men_men_n901_));
  NA2        u0879(.A(i_11_), .B(i_9_), .Y(men_men_n902_));
  NO3        u0880(.A(i_12_), .B(men_men_n902_), .C(men_men_n606_), .Y(men_men_n903_));
  AN2        u0881(.A(men_men_n903_), .B(men_men_n901_), .Y(men_men_n904_));
  NO2        u0882(.A(men_men_n49_), .B(i_7_), .Y(men_men_n905_));
  NA2        u0883(.A(men_men_n389_), .B(men_men_n182_), .Y(men_men_n906_));
  NA2        u0884(.A(men_men_n906_), .B(men_men_n162_), .Y(men_men_n907_));
  NO2        u0885(.A(men_men_n902_), .B(men_men_n74_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n178_), .B(i_0_), .Y(men_men_n909_));
  INV        u0887(.A(men_men_n909_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n474_), .B(men_men_n231_), .Y(men_men_n911_));
  AOI210     u0889(.A0(men_men_n364_), .A1(men_men_n42_), .B0(men_men_n403_), .Y(men_men_n912_));
  OAI220     u0890(.A0(men_men_n912_), .A1(men_men_n867_), .B0(men_men_n911_), .B1(men_men_n910_), .Y(men_men_n913_));
  NO3        u0891(.A(men_men_n913_), .B(men_men_n907_), .C(men_men_n904_), .Y(men_men_n914_));
  NA2        u0892(.A(men_men_n665_), .B(men_men_n123_), .Y(men_men_n915_));
  NO2        u0893(.A(i_6_), .B(men_men_n915_), .Y(men_men_n916_));
  AOI210     u0894(.A0(men_men_n444_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n917_));
  NA2        u0895(.A(men_men_n174_), .B(men_men_n105_), .Y(men_men_n918_));
  NOi32      u0896(.An(men_men_n917_), .Bn(men_men_n188_), .C(men_men_n918_), .Y(men_men_n919_));
  NO2        u0897(.A(men_men_n919_), .B(men_men_n916_), .Y(men_men_n920_));
  NOi21      u0898(.An(i_7_), .B(i_5_), .Y(men_men_n921_));
  NOi31      u0899(.An(men_men_n921_), .B(i_0_), .C(men_men_n736_), .Y(men_men_n922_));
  NA3        u0900(.A(men_men_n922_), .B(men_men_n378_), .C(i_6_), .Y(men_men_n923_));
  OA210      u0901(.A0(men_men_n918_), .A1(men_men_n520_), .B0(men_men_n923_), .Y(men_men_n924_));
  NO3        u0902(.A(men_men_n398_), .B(men_men_n353_), .C(men_men_n349_), .Y(men_men_n925_));
  NO2        u0903(.A(men_men_n261_), .B(men_men_n308_), .Y(men_men_n926_));
  NO2        u0904(.A(men_men_n736_), .B(men_men_n256_), .Y(men_men_n927_));
  AOI210     u0905(.A0(men_men_n927_), .A1(men_men_n926_), .B0(men_men_n925_), .Y(men_men_n928_));
  NA4        u0906(.A(men_men_n928_), .B(men_men_n924_), .C(men_men_n920_), .D(men_men_n914_), .Y(men_men_n929_));
  NO2        u0907(.A(men_men_n875_), .B(men_men_n239_), .Y(men_men_n930_));
  AN2        u0908(.A(men_men_n322_), .B(men_men_n317_), .Y(men_men_n931_));
  AN2        u0909(.A(men_men_n931_), .B(men_men_n871_), .Y(men_men_n932_));
  OAI210     u0910(.A0(men_men_n932_), .A1(men_men_n930_), .B0(i_10_), .Y(men_men_n933_));
  NO2        u0911(.A(men_men_n851_), .B(men_men_n307_), .Y(men_men_n934_));
  NA2        u0912(.A(men_men_n934_), .B(men_men_n908_), .Y(men_men_n935_));
  NA3        u0913(.A(men_men_n473_), .B(men_men_n407_), .C(men_men_n46_), .Y(men_men_n936_));
  OAI210     u0914(.A0(men_men_n877_), .A1(men_men_n886_), .B0(men_men_n936_), .Y(men_men_n937_));
  NO2        u0915(.A(men_men_n254_), .B(men_men_n47_), .Y(men_men_n938_));
  NA2        u0916(.A(men_men_n908_), .B(men_men_n294_), .Y(men_men_n939_));
  OAI210     u0917(.A0(men_men_n938_), .A1(men_men_n187_), .B0(men_men_n939_), .Y(men_men_n940_));
  AOI220     u0918(.A0(men_men_n940_), .A1(men_men_n474_), .B0(men_men_n937_), .B1(men_men_n74_), .Y(men_men_n941_));
  NA3        u0919(.A(men_men_n828_), .B(men_men_n376_), .C(men_men_n646_), .Y(men_men_n942_));
  NO2        u0920(.A(men_men_n942_), .B(men_men_n48_), .Y(men_men_n943_));
  NO3        u0921(.A(men_men_n591_), .B(men_men_n348_), .C(men_men_n24_), .Y(men_men_n944_));
  AOI210     u0922(.A0(men_men_n711_), .A1(men_men_n550_), .B0(men_men_n944_), .Y(men_men_n945_));
  NAi21      u0923(.An(i_9_), .B(i_5_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n946_), .B(men_men_n398_), .Y(men_men_n947_));
  NA2        u0925(.A(men_men_n947_), .B(men_men_n625_), .Y(men_men_n948_));
  OAI220     u0926(.A0(men_men_n948_), .A1(men_men_n87_), .B0(men_men_n945_), .B1(men_men_n175_), .Y(men_men_n949_));
  NO3        u0927(.A(men_men_n949_), .B(men_men_n943_), .C(men_men_n525_), .Y(men_men_n950_));
  NA4        u0928(.A(men_men_n950_), .B(men_men_n941_), .C(men_men_n935_), .D(men_men_n933_), .Y(men_men_n951_));
  NO3        u0929(.A(men_men_n951_), .B(men_men_n929_), .C(men_men_n900_), .Y(men_men_n952_));
  NO2        u0930(.A(i_0_), .B(men_men_n736_), .Y(men_men_n953_));
  NA2        u0931(.A(men_men_n74_), .B(men_men_n45_), .Y(men_men_n954_));
  INV        u0932(.A(men_men_n954_), .Y(men_men_n955_));
  NO3        u0933(.A(men_men_n107_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n956_));
  AO220      u0934(.A0(men_men_n956_), .A1(men_men_n955_), .B0(men_men_n953_), .B1(men_men_n177_), .Y(men_men_n957_));
  NO2        u0935(.A(men_men_n808_), .B(men_men_n918_), .Y(men_men_n958_));
  AOI210     u0936(.A0(men_men_n957_), .A1(men_men_n337_), .B0(men_men_n958_), .Y(men_men_n959_));
  NA2        u0937(.A(men_men_n747_), .B(men_men_n148_), .Y(men_men_n960_));
  INV        u0938(.A(men_men_n960_), .Y(men_men_n961_));
  NA3        u0939(.A(men_men_n961_), .B(men_men_n682_), .C(men_men_n74_), .Y(men_men_n962_));
  OAI210     u0940(.A0(men_men_n242_), .A1(i_9_), .B0(men_men_n230_), .Y(men_men_n963_));
  AOI210     u0941(.A0(men_men_n963_), .A1(men_men_n882_), .B0(men_men_n155_), .Y(men_men_n964_));
  INV        u0942(.A(men_men_n964_), .Y(men_men_n965_));
  NA3        u0943(.A(men_men_n965_), .B(men_men_n962_), .C(men_men_n959_), .Y(men_men_n966_));
  NA2        u0944(.A(men_men_n931_), .B(men_men_n366_), .Y(men_men_n967_));
  AOI210     u0945(.A0(men_men_n289_), .A1(men_men_n164_), .B0(men_men_n967_), .Y(men_men_n968_));
  NA3        u0946(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n969_));
  NA2        u0947(.A(men_men_n905_), .B(men_men_n490_), .Y(men_men_n970_));
  AOI210     u0948(.A0(men_men_n969_), .A1(men_men_n164_), .B0(men_men_n970_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n971_), .B(men_men_n968_), .Y(men_men_n972_));
  NO3        u0950(.A(men_men_n891_), .B(men_men_n866_), .C(men_men_n190_), .Y(men_men_n973_));
  AOI220     u0951(.A0(men_men_n973_), .A1(i_11_), .B0(men_men_n574_), .B1(men_men_n76_), .Y(men_men_n974_));
  NO3        u0952(.A(men_men_n211_), .B(men_men_n377_), .C(i_0_), .Y(men_men_n975_));
  OAI210     u0953(.A0(men_men_n975_), .A1(men_men_n77_), .B0(i_13_), .Y(men_men_n976_));
  INV        u0954(.A(men_men_n219_), .Y(men_men_n977_));
  OAI220     u0955(.A0(men_men_n537_), .A1(men_men_n141_), .B0(men_men_n651_), .B1(men_men_n619_), .Y(men_men_n978_));
  NA3        u0956(.A(men_men_n978_), .B(men_men_n393_), .C(men_men_n977_), .Y(men_men_n979_));
  NA4        u0957(.A(men_men_n979_), .B(men_men_n976_), .C(men_men_n974_), .D(men_men_n972_), .Y(men_men_n980_));
  AOI220     u0958(.A0(men_men_n921_), .A1(men_men_n490_), .B0(men_men_n853_), .B1(men_men_n165_), .Y(men_men_n981_));
  NA2        u0959(.A(men_men_n340_), .B(men_men_n179_), .Y(men_men_n982_));
  OR2        u0960(.A(men_men_n982_), .B(men_men_n981_), .Y(men_men_n983_));
  NA3        u0961(.A(men_men_n616_), .B(men_men_n185_), .C(men_men_n85_), .Y(men_men_n984_));
  NA2        u0962(.A(men_men_n984_), .B(men_men_n548_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n495_), .B(men_men_n488_), .Y(men_men_n986_));
  NO2        u0964(.A(men_men_n986_), .B(men_men_n985_), .Y(men_men_n987_));
  NA3        u0965(.A(men_men_n384_), .B(men_men_n174_), .C(men_men_n173_), .Y(men_men_n988_));
  INV        u0966(.A(men_men_n988_), .Y(men_men_n989_));
  NA3        u0967(.A(men_men_n384_), .B(men_men_n324_), .C(men_men_n221_), .Y(men_men_n990_));
  INV        u0968(.A(men_men_n990_), .Y(men_men_n991_));
  NOi31      u0969(.An(men_men_n383_), .B(men_men_n954_), .C(men_men_n239_), .Y(men_men_n992_));
  NO3        u0970(.A(men_men_n902_), .B(men_men_n219_), .C(men_men_n190_), .Y(men_men_n993_));
  NO4        u0971(.A(men_men_n993_), .B(men_men_n992_), .C(men_men_n991_), .D(men_men_n989_), .Y(men_men_n994_));
  NA3        u0972(.A(men_men_n994_), .B(men_men_n987_), .C(men_men_n983_), .Y(men_men_n995_));
  INV        u0973(.A(men_men_n618_), .Y(men_men_n996_));
  NO3        u0974(.A(men_men_n996_), .B(men_men_n564_), .C(men_men_n334_), .Y(men_men_n997_));
  NO2        u0975(.A(men_men_n87_), .B(i_5_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n854_), .B(men_men_n111_), .C(men_men_n126_), .Y(men_men_n999_));
  INV        u0977(.A(men_men_n999_), .Y(men_men_n1000_));
  AOI210     u0978(.A0(men_men_n1000_), .A1(men_men_n998_), .B0(men_men_n997_), .Y(men_men_n1001_));
  NA3        u0979(.A(men_men_n294_), .B(i_5_), .C(men_men_n193_), .Y(men_men_n1002_));
  NAi31      u0980(.An(men_men_n240_), .B(men_men_n1002_), .C(men_men_n241_), .Y(men_men_n1003_));
  NO4        u0981(.A(men_men_n239_), .B(men_men_n211_), .C(i_0_), .D(i_12_), .Y(men_men_n1004_));
  AOI220     u0982(.A0(men_men_n1004_), .A1(men_men_n1003_), .B0(men_men_n802_), .B1(men_men_n179_), .Y(men_men_n1005_));
  AN2        u0983(.A(men_men_n891_), .B(men_men_n155_), .Y(men_men_n1006_));
  NO4        u0984(.A(men_men_n1006_), .B(i_12_), .C(men_men_n655_), .D(men_men_n133_), .Y(men_men_n1007_));
  NA2        u0985(.A(men_men_n1007_), .B(men_men_n219_), .Y(men_men_n1008_));
  NA3        u0986(.A(men_men_n100_), .B(men_men_n578_), .C(i_11_), .Y(men_men_n1009_));
  NO2        u0987(.A(men_men_n1009_), .B(men_men_n157_), .Y(men_men_n1010_));
  NA2        u0988(.A(men_men_n921_), .B(men_men_n471_), .Y(men_men_n1011_));
  NA2        u0989(.A(men_men_n65_), .B(men_men_n103_), .Y(men_men_n1012_));
  OAI220     u0990(.A0(men_men_n1012_), .A1(men_men_n1002_), .B0(men_men_n1011_), .B1(men_men_n683_), .Y(men_men_n1013_));
  AOI210     u0991(.A0(men_men_n1013_), .A1(men_men_n909_), .B0(men_men_n1010_), .Y(men_men_n1014_));
  NA4        u0992(.A(men_men_n1014_), .B(men_men_n1008_), .C(men_men_n1005_), .D(men_men_n1001_), .Y(men_men_n1015_));
  NO4        u0993(.A(men_men_n1015_), .B(men_men_n995_), .C(men_men_n980_), .D(men_men_n966_), .Y(men_men_n1016_));
  OAI210     u0994(.A0(men_men_n827_), .A1(men_men_n821_), .B0(men_men_n37_), .Y(men_men_n1017_));
  NA2        u0995(.A(men_men_n1017_), .B(men_men_n614_), .Y(men_men_n1018_));
  NA2        u0996(.A(men_men_n1018_), .B(men_men_n208_), .Y(men_men_n1019_));
  AN2        u0997(.A(men_men_n706_), .B(men_men_n362_), .Y(men_men_n1020_));
  NA2        u0998(.A(men_men_n186_), .B(men_men_n188_), .Y(men_men_n1021_));
  AO210      u0999(.A0(men_men_n1020_), .A1(men_men_n33_), .B0(men_men_n1021_), .Y(men_men_n1022_));
  OAI210     u1000(.A0(men_men_n618_), .A1(men_men_n616_), .B0(men_men_n307_), .Y(men_men_n1023_));
  NAi31      u1001(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1024_));
  AOI210     u1002(.A0(men_men_n119_), .A1(men_men_n71_), .B0(men_men_n1024_), .Y(men_men_n1025_));
  NO2        u1003(.A(men_men_n1025_), .B(men_men_n652_), .Y(men_men_n1026_));
  NA3        u1004(.A(men_men_n1026_), .B(men_men_n1023_), .C(men_men_n1022_), .Y(men_men_n1027_));
  NO2        u1005(.A(men_men_n461_), .B(men_men_n266_), .Y(men_men_n1028_));
  NO4        u1006(.A(men_men_n233_), .B(men_men_n147_), .C(men_men_n686_), .D(men_men_n37_), .Y(men_men_n1029_));
  NO3        u1007(.A(men_men_n1029_), .B(men_men_n1028_), .C(men_men_n884_), .Y(men_men_n1030_));
  OAI210     u1008(.A0(men_men_n1009_), .A1(men_men_n150_), .B0(men_men_n1030_), .Y(men_men_n1031_));
  AOI210     u1009(.A0(men_men_n1027_), .A1(men_men_n49_), .B0(men_men_n1031_), .Y(men_men_n1032_));
  AOI210     u1010(.A0(men_men_n1032_), .A1(men_men_n1019_), .B0(men_men_n74_), .Y(men_men_n1033_));
  NO2        u1011(.A(men_men_n571_), .B(men_men_n373_), .Y(men_men_n1034_));
  NO2        u1012(.A(men_men_n1034_), .B(men_men_n766_), .Y(men_men_n1035_));
  NA3        u1013(.A(men_men_n98_), .B(men_men_n296_), .C(men_men_n31_), .Y(men_men_n1036_));
  NA2        u1014(.A(men_men_n160_), .B(men_men_n88_), .Y(men_men_n1037_));
  NA3        u1015(.A(men_men_n770_), .B(men_men_n278_), .C(men_men_n81_), .Y(men_men_n1038_));
  AOI210     u1016(.A0(men_men_n1038_), .A1(men_men_n1037_), .B0(i_11_), .Y(men_men_n1039_));
  NA2        u1017(.A(men_men_n609_), .B(men_men_n217_), .Y(men_men_n1040_));
  OAI210     u1018(.A0(men_men_n1040_), .A1(men_men_n917_), .B0(men_men_n208_), .Y(men_men_n1041_));
  NA2        u1019(.A(men_men_n166_), .B(i_5_), .Y(men_men_n1042_));
  NO2        u1020(.A(men_men_n1041_), .B(men_men_n1042_), .Y(men_men_n1043_));
  NO3        u1021(.A(men_men_n60_), .B(men_men_n59_), .C(i_4_), .Y(men_men_n1044_));
  OAI210     u1022(.A0(men_men_n926_), .A1(men_men_n296_), .B0(men_men_n1044_), .Y(men_men_n1045_));
  NO2        u1023(.A(men_men_n1045_), .B(men_men_n736_), .Y(men_men_n1046_));
  NO4        u1024(.A(men_men_n946_), .B(men_men_n478_), .C(men_men_n251_), .D(men_men_n250_), .Y(men_men_n1047_));
  NO2        u1025(.A(men_men_n1047_), .B(men_men_n568_), .Y(men_men_n1048_));
  INV        u1026(.A(men_men_n354_), .Y(men_men_n1049_));
  AOI210     u1027(.A0(men_men_n1049_), .A1(men_men_n1048_), .B0(men_men_n41_), .Y(men_men_n1050_));
  NO4        u1028(.A(men_men_n1050_), .B(men_men_n1046_), .C(men_men_n1043_), .D(men_men_n1039_), .Y(men_men_n1051_));
  OAI210     u1029(.A0(men_men_n1036_), .A1(i_4_), .B0(men_men_n1051_), .Y(men_men_n1052_));
  NO3        u1030(.A(men_men_n1052_), .B(men_men_n1035_), .C(men_men_n1033_), .Y(men_men_n1053_));
  NA4        u1031(.A(men_men_n1053_), .B(men_men_n1016_), .C(men_men_n952_), .D(men_men_n874_), .Y(men4));
  INV        u1032(.A(men_men_n710_), .Y(men_men_n1057_));
  INV        u1033(.A(men_men_n485_), .Y(men_men_n1058_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule