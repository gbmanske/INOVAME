//Benchmark atmr_max1024_476_0.125

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n354_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n451_, men_men_n452_, men_men_n453_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  INV        o005(.A(ori_ori_n19_), .Y(ori_ori_n22_));
  NA2        o006(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n23_));
  INV        o007(.A(x5), .Y(ori_ori_n24_));
  NA2        o008(.A(x7), .B(x6), .Y(ori_ori_n25_));
  NA2        o009(.A(x4), .B(x2), .Y(ori_ori_n26_));
  INV        o010(.A(ori_ori_n23_), .Y(ori_ori_n27_));
  NO2        o011(.A(x4), .B(x3), .Y(ori_ori_n28_));
  INV        o012(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  NOi21      o013(.An(ori_ori_n22_), .B(ori_ori_n27_), .Y(ori00));
  NO2        o014(.A(x1), .B(x0), .Y(ori_ori_n31_));
  INV        o015(.A(x6), .Y(ori_ori_n32_));
  NO2        o016(.A(ori_ori_n32_), .B(ori_ori_n24_), .Y(ori_ori_n33_));
  NA2        o017(.A(x4), .B(x3), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n22_), .B(ori_ori_n34_), .Y(ori_ori_n35_));
  NO2        o019(.A(x2), .B(x0), .Y(ori_ori_n36_));
  INV        o020(.A(x3), .Y(ori_ori_n37_));
  NO2        o021(.A(ori_ori_n37_), .B(ori_ori_n18_), .Y(ori_ori_n38_));
  INV        o022(.A(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o023(.A(ori_ori_n33_), .B(x4), .Y(ori_ori_n40_));
  OAI210     o024(.A0(ori_ori_n40_), .A1(ori_ori_n39_), .B0(ori_ori_n36_), .Y(ori_ori_n41_));
  INV        o025(.A(x4), .Y(ori_ori_n42_));
  NO2        o026(.A(ori_ori_n42_), .B(ori_ori_n17_), .Y(ori_ori_n43_));
  NA2        o027(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n44_), .A1(ori_ori_n20_), .B0(ori_ori_n41_), .Y(ori_ori_n45_));
  INV        o029(.A(ori_ori_n31_), .Y(ori_ori_n46_));
  INV        o030(.A(x2), .Y(ori_ori_n47_));
  NO2        o031(.A(ori_ori_n47_), .B(ori_ori_n17_), .Y(ori_ori_n48_));
  NA2        o032(.A(ori_ori_n37_), .B(ori_ori_n18_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(ori_ori_n48_), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n46_), .A1(ori_ori_n29_), .B0(ori_ori_n50_), .Y(ori_ori_n51_));
  NO3        o035(.A(ori_ori_n51_), .B(ori_ori_n45_), .C(ori_ori_n35_), .Y(ori01));
  NA2        o036(.A(x8), .B(x7), .Y(ori_ori_n53_));
  NA2        o037(.A(ori_ori_n37_), .B(x1), .Y(ori_ori_n54_));
  INV        o038(.A(x6), .Y(ori_ori_n55_));
  NO2        o039(.A(ori_ori_n54_), .B(x5), .Y(ori_ori_n56_));
  NO2        o040(.A(x8), .B(x2), .Y(ori_ori_n57_));
  INV        o041(.A(ori_ori_n57_), .Y(ori_ori_n58_));
  OAI210     o042(.A0(ori_ori_n38_), .A1(ori_ori_n24_), .B0(ori_ori_n47_), .Y(ori_ori_n59_));
  OAI210     o043(.A0(ori_ori_n49_), .A1(ori_ori_n20_), .B0(ori_ori_n59_), .Y(ori_ori_n60_));
  INV        o044(.A(ori_ori_n60_), .Y(ori_ori_n61_));
  NA2        o045(.A(ori_ori_n61_), .B(x4), .Y(ori_ori_n62_));
  NA2        o046(.A(ori_ori_n42_), .B(x2), .Y(ori_ori_n63_));
  OAI210     o047(.A0(ori_ori_n63_), .A1(ori_ori_n49_), .B0(x0), .Y(ori_ori_n64_));
  NA2        o048(.A(x5), .B(x3), .Y(ori_ori_n65_));
  NO2        o049(.A(x8), .B(x6), .Y(ori_ori_n66_));
  NO3        o050(.A(ori_ori_n65_), .B(ori_ori_n55_), .C(ori_ori_n47_), .Y(ori_ori_n67_));
  NAi21      o051(.An(x4), .B(x3), .Y(ori_ori_n68_));
  INV        o052(.A(ori_ori_n68_), .Y(ori_ori_n69_));
  NO2        o053(.A(x4), .B(x2), .Y(ori_ori_n70_));
  NO2        o054(.A(ori_ori_n68_), .B(ori_ori_n18_), .Y(ori_ori_n71_));
  NO3        o055(.A(ori_ori_n71_), .B(ori_ori_n67_), .C(ori_ori_n64_), .Y(ori_ori_n72_));
  NA2        o056(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n74_));
  INV        o058(.A(x8), .Y(ori_ori_n75_));
  NA2        o059(.A(x2), .B(x1), .Y(ori_ori_n76_));
  INV        o060(.A(ori_ori_n74_), .Y(ori_ori_n77_));
  NO2        o061(.A(ori_ori_n77_), .B(ori_ori_n25_), .Y(ori_ori_n78_));
  AOI210     o062(.A0(ori_ori_n49_), .A1(ori_ori_n24_), .B0(ori_ori_n47_), .Y(ori_ori_n79_));
  OAI210     o063(.A0(ori_ori_n39_), .A1(ori_ori_n33_), .B0(ori_ori_n42_), .Y(ori_ori_n80_));
  NO3        o064(.A(ori_ori_n80_), .B(ori_ori_n79_), .C(ori_ori_n78_), .Y(ori_ori_n81_));
  NA2        o065(.A(x4), .B(ori_ori_n37_), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n42_), .B(ori_ori_n47_), .Y(ori_ori_n83_));
  NO2        o067(.A(ori_ori_n82_), .B(x1), .Y(ori_ori_n84_));
  NO2        o068(.A(x3), .B(x2), .Y(ori_ori_n85_));
  NA3        o069(.A(ori_ori_n85_), .B(ori_ori_n25_), .C(ori_ori_n24_), .Y(ori_ori_n86_));
  INV        o070(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  NA2        o071(.A(ori_ori_n47_), .B(x1), .Y(ori_ori_n88_));
  OAI210     o072(.A0(ori_ori_n88_), .A1(ori_ori_n34_), .B0(ori_ori_n17_), .Y(ori_ori_n89_));
  NO4        o073(.A(ori_ori_n89_), .B(ori_ori_n87_), .C(ori_ori_n84_), .D(ori_ori_n81_), .Y(ori_ori_n90_));
  AO210      o074(.A0(ori_ori_n72_), .A1(ori_ori_n62_), .B0(ori_ori_n90_), .Y(ori02));
  NO2        o075(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n92_));
  NA2        o076(.A(ori_ori_n37_), .B(x0), .Y(ori_ori_n93_));
  BUFFER     o077(.A(x0), .Y(ori_ori_n94_));
  INV        o078(.A(ori_ori_n94_), .Y(ori_ori_n95_));
  NO2        o079(.A(x4), .B(x1), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n96_), .B(x2), .Y(ori_ori_n97_));
  NOi21      o081(.An(x0), .B(x1), .Y(ori_ori_n98_));
  NOi21      o082(.An(x0), .B(x4), .Y(ori_ori_n99_));
  NO2        o083(.A(ori_ori_n97_), .B(ori_ori_n65_), .Y(ori_ori_n100_));
  NO2        o084(.A(x5), .B(ori_ori_n42_), .Y(ori_ori_n101_));
  NA2        o085(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n102_));
  AOI210     o086(.A0(ori_ori_n102_), .A1(ori_ori_n88_), .B0(ori_ori_n93_), .Y(ori_ori_n103_));
  OAI210     o087(.A0(ori_ori_n103_), .A1(ori_ori_n31_), .B0(ori_ori_n101_), .Y(ori_ori_n104_));
  NAi21      o088(.An(x0), .B(x4), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n105_), .B(x1), .Y(ori_ori_n106_));
  NO2        o090(.A(x7), .B(x0), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n70_), .B(ori_ori_n83_), .Y(ori_ori_n108_));
  NO2        o092(.A(ori_ori_n108_), .B(x3), .Y(ori_ori_n109_));
  OAI210     o093(.A0(ori_ori_n107_), .A1(ori_ori_n106_), .B0(ori_ori_n109_), .Y(ori_ori_n110_));
  NA2        o094(.A(x5), .B(x0), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n42_), .B(x2), .Y(ori_ori_n112_));
  NA3        o096(.A(ori_ori_n110_), .B(ori_ori_n104_), .C(ori_ori_n32_), .Y(ori_ori_n113_));
  NO2        o097(.A(ori_ori_n113_), .B(ori_ori_n100_), .Y(ori_ori_n114_));
  NO3        o098(.A(ori_ori_n65_), .B(ori_ori_n63_), .C(ori_ori_n23_), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n26_), .B(ori_ori_n24_), .Y(ori_ori_n116_));
  NA2        o100(.A(x7), .B(x3), .Y(ori_ori_n117_));
  NO2        o101(.A(ori_ori_n82_), .B(x5), .Y(ori_ori_n118_));
  NO2        o102(.A(ori_ori_n37_), .B(x2), .Y(ori_ori_n119_));
  INV        o103(.A(x7), .Y(ori_ori_n120_));
  NA2        o104(.A(ori_ori_n120_), .B(ori_ori_n18_), .Y(ori_ori_n121_));
  NA2        o105(.A(ori_ori_n121_), .B(ori_ori_n119_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n24_), .B(x4), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n123_), .B(ori_ori_n99_), .Y(ori_ori_n124_));
  NO2        o108(.A(ori_ori_n124_), .B(ori_ori_n122_), .Y(ori_ori_n125_));
  INV        o109(.A(ori_ori_n125_), .Y(ori_ori_n126_));
  OAI210     o110(.A0(ori_ori_n117_), .A1(ori_ori_n44_), .B0(ori_ori_n126_), .Y(ori_ori_n127_));
  NA2        o111(.A(x5), .B(x1), .Y(ori_ori_n128_));
  INV        o112(.A(ori_ori_n128_), .Y(ori_ori_n129_));
  AOI210     o113(.A0(ori_ori_n129_), .A1(ori_ori_n99_), .B0(ori_ori_n32_), .Y(ori_ori_n130_));
  NAi21      o114(.An(x2), .B(x7), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n131_), .B(ori_ori_n42_), .Y(ori_ori_n132_));
  NA2        o116(.A(ori_ori_n132_), .B(ori_ori_n56_), .Y(ori_ori_n133_));
  NA2        o117(.A(ori_ori_n133_), .B(ori_ori_n130_), .Y(ori_ori_n134_));
  NO3        o118(.A(ori_ori_n134_), .B(ori_ori_n127_), .C(ori_ori_n115_), .Y(ori_ori_n135_));
  NO2        o119(.A(ori_ori_n135_), .B(ori_ori_n114_), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n111_), .B(ori_ori_n108_), .Y(ori_ori_n137_));
  NA2        o121(.A(ori_ori_n24_), .B(ori_ori_n18_), .Y(ori_ori_n138_));
  NA2        o122(.A(ori_ori_n24_), .B(ori_ori_n17_), .Y(ori_ori_n139_));
  NA3        o123(.A(ori_ori_n139_), .B(ori_ori_n138_), .C(ori_ori_n23_), .Y(ori_ori_n140_));
  AN2        o124(.A(ori_ori_n140_), .B(ori_ori_n112_), .Y(ori_ori_n141_));
  NA2        o125(.A(x8), .B(x0), .Y(ori_ori_n142_));
  NO2        o126(.A(ori_ori_n120_), .B(ori_ori_n24_), .Y(ori_ori_n143_));
  NA2        o127(.A(x2), .B(x0), .Y(ori_ori_n144_));
  NA2        o128(.A(x4), .B(x1), .Y(ori_ori_n145_));
  NAi21      o129(.An(ori_ori_n96_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NOi31      o130(.An(ori_ori_n146_), .B(ori_ori_n123_), .C(ori_ori_n144_), .Y(ori_ori_n147_));
  NO3        o131(.A(ori_ori_n147_), .B(ori_ori_n141_), .C(ori_ori_n137_), .Y(ori_ori_n148_));
  NO2        o132(.A(ori_ori_n148_), .B(ori_ori_n37_), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n140_), .B(ori_ori_n63_), .Y(ori_ori_n150_));
  INV        o134(.A(ori_ori_n101_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n88_), .B(ori_ori_n17_), .Y(ori_ori_n152_));
  AOI210     o136(.A0(ori_ori_n31_), .A1(ori_ori_n75_), .B0(ori_ori_n152_), .Y(ori_ori_n153_));
  NO3        o137(.A(ori_ori_n153_), .B(ori_ori_n151_), .C(x7), .Y(ori_ori_n154_));
  NA3        o138(.A(ori_ori_n146_), .B(ori_ori_n151_), .C(ori_ori_n36_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n139_), .A1(ori_ori_n108_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NO3        o140(.A(ori_ori_n156_), .B(ori_ori_n154_), .C(ori_ori_n150_), .Y(ori_ori_n157_));
  NO2        o141(.A(ori_ori_n157_), .B(x3), .Y(ori_ori_n158_));
  NO3        o142(.A(ori_ori_n158_), .B(ori_ori_n149_), .C(ori_ori_n136_), .Y(ori03));
  NO2        o143(.A(ori_ori_n42_), .B(x3), .Y(ori_ori_n160_));
  NO2        o144(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n161_));
  NA2        o145(.A(x6), .B(ori_ori_n24_), .Y(ori_ori_n162_));
  NO2        o146(.A(ori_ori_n162_), .B(x4), .Y(ori_ori_n163_));
  NO2        o147(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n164_));
  NA2        o148(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n165_));
  NO3        o149(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n166_));
  NO2        o150(.A(x5), .B(x1), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n165_), .B(ori_ori_n138_), .Y(ori_ori_n168_));
  NO3        o152(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  INV        o154(.A(ori_ori_n170_), .Y(ori_ori_n171_));
  AOI220     o155(.A0(ori_ori_n171_), .A1(ori_ori_n42_), .B0(ori_ori_n166_), .B1(ori_ori_n101_), .Y(ori_ori_n172_));
  INV        o156(.A(ori_ori_n172_), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n42_), .B(ori_ori_n37_), .Y(ori_ori_n174_));
  NA2        o158(.A(ori_ori_n174_), .B(ori_ori_n19_), .Y(ori_ori_n175_));
  NO2        o159(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n176_));
  NO2        o160(.A(ori_ori_n176_), .B(x6), .Y(ori_ori_n177_));
  NOi21      o161(.An(ori_ori_n70_), .B(ori_ori_n177_), .Y(ori_ori_n178_));
  NA2        o162(.A(ori_ori_n176_), .B(x6), .Y(ori_ori_n179_));
  AOI210     o163(.A0(ori_ori_n179_), .A1(ori_ori_n178_), .B0(ori_ori_n120_), .Y(ori_ori_n180_));
  OR2        o164(.A(ori_ori_n180_), .B(ori_ori_n143_), .Y(ori_ori_n181_));
  NA2        o165(.A(ori_ori_n37_), .B(ori_ori_n47_), .Y(ori_ori_n182_));
  NA2        o166(.A(ori_ori_n112_), .B(ori_ori_n74_), .Y(ori_ori_n183_));
  NA2        o167(.A(x6), .B(ori_ori_n42_), .Y(ori_ori_n184_));
  OAI210     o168(.A0(ori_ori_n95_), .A1(ori_ori_n66_), .B0(x4), .Y(ori_ori_n185_));
  AOI210     o169(.A0(ori_ori_n185_), .A1(ori_ori_n184_), .B0(ori_ori_n65_), .Y(ori_ori_n186_));
  NA2        o170(.A(ori_ori_n161_), .B(ori_ori_n106_), .Y(ori_ori_n187_));
  NA3        o171(.A(ori_ori_n165_), .B(ori_ori_n101_), .C(x6), .Y(ori_ori_n188_));
  INV        o172(.A(ori_ori_n56_), .Y(ori_ori_n189_));
  NA3        o173(.A(ori_ori_n189_), .B(ori_ori_n188_), .C(ori_ori_n187_), .Y(ori_ori_n190_));
  OAI210     o174(.A0(ori_ori_n190_), .A1(ori_ori_n186_), .B0(x2), .Y(ori_ori_n191_));
  NA3        o175(.A(ori_ori_n191_), .B(ori_ori_n183_), .C(ori_ori_n181_), .Y(ori_ori_n192_));
  AOI210     o176(.A0(ori_ori_n173_), .A1(x8), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  NO2        o177(.A(ori_ori_n75_), .B(x3), .Y(ori_ori_n194_));
  NA2        o178(.A(ori_ori_n194_), .B(ori_ori_n163_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n196_));
  AOI210     o180(.A0(ori_ori_n177_), .A1(ori_ori_n123_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  AOI210     o181(.A0(ori_ori_n197_), .A1(ori_ori_n195_), .B0(x2), .Y(ori_ori_n198_));
  AOI220     o182(.A0(ori_ori_n163_), .A1(ori_ori_n152_), .B0(x2), .B1(ori_ori_n56_), .Y(ori_ori_n199_));
  NA2        o183(.A(ori_ori_n37_), .B(ori_ori_n17_), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n200_), .B(ori_ori_n24_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n201_), .B(ori_ori_n96_), .Y(ori_ori_n202_));
  NA2        o186(.A(ori_ori_n165_), .B(x6), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n165_), .B(x6), .Y(ori_ori_n204_));
  INV        o188(.A(ori_ori_n204_), .Y(ori_ori_n205_));
  NA3        o189(.A(ori_ori_n205_), .B(ori_ori_n203_), .C(ori_ori_n116_), .Y(ori_ori_n206_));
  NA4        o190(.A(ori_ori_n206_), .B(ori_ori_n202_), .C(ori_ori_n199_), .D(ori_ori_n120_), .Y(ori_ori_n207_));
  NA2        o191(.A(ori_ori_n161_), .B(ori_ori_n176_), .Y(ori_ori_n208_));
  NAi21      o192(.An(x1), .B(x4), .Y(ori_ori_n209_));
  AOI210     o193(.A0(x3), .A1(x2), .B0(ori_ori_n42_), .Y(ori_ori_n210_));
  OAI210     o194(.A0(ori_ori_n111_), .A1(x3), .B0(ori_ori_n210_), .Y(ori_ori_n211_));
  NA2        o195(.A(ori_ori_n211_), .B(ori_ori_n209_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n212_), .B(ori_ori_n208_), .Y(ori_ori_n213_));
  NA2        o197(.A(x6), .B(x2), .Y(ori_ori_n214_));
  NA2        o198(.A(x4), .B(ori_ori_n213_), .Y(ori_ori_n215_));
  NO2        o199(.A(x3), .B(ori_ori_n162_), .Y(ori_ori_n216_));
  BUFFER     o200(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  NA2        o201(.A(x4), .B(x0), .Y(ori_ori_n218_));
  NA2        o202(.A(ori_ori_n217_), .B(ori_ori_n36_), .Y(ori_ori_n219_));
  AOI210     o203(.A0(ori_ori_n219_), .A1(ori_ori_n215_), .B0(x8), .Y(ori_ori_n220_));
  OAI210     o204(.A0(x0), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n221_));
  NO2        o205(.A(ori_ori_n221_), .B(ori_ori_n182_), .Y(ori_ori_n222_));
  NO4        o206(.A(ori_ori_n222_), .B(ori_ori_n220_), .C(ori_ori_n207_), .D(ori_ori_n198_), .Y(ori_ori_n223_));
  OAI210     o207(.A0(x1), .A1(ori_ori_n204_), .B0(x2), .Y(ori_ori_n224_));
  OAI210     o208(.A0(x0), .A1(x6), .B0(ori_ori_n38_), .Y(ori_ori_n225_));
  AOI210     o209(.A0(ori_ori_n225_), .A1(ori_ori_n224_), .B0(ori_ori_n151_), .Y(ori_ori_n226_));
  NOi21      o210(.An(ori_ori_n214_), .B(ori_ori_n17_), .Y(ori_ori_n227_));
  NA3        o211(.A(ori_ori_n227_), .B(ori_ori_n167_), .C(ori_ori_n34_), .Y(ori_ori_n228_));
  AOI210     o212(.A0(ori_ori_n32_), .A1(ori_ori_n47_), .B0(x0), .Y(ori_ori_n229_));
  NA3        o213(.A(ori_ori_n229_), .B(ori_ori_n129_), .C(ori_ori_n29_), .Y(ori_ori_n230_));
  NA2        o214(.A(x3), .B(x2), .Y(ori_ori_n231_));
  AOI220     o215(.A0(ori_ori_n231_), .A1(ori_ori_n182_), .B0(ori_ori_n230_), .B1(ori_ori_n228_), .Y(ori_ori_n232_));
  NAi21      o216(.An(x4), .B(x0), .Y(ori_ori_n233_));
  NO3        o217(.A(ori_ori_n233_), .B(ori_ori_n38_), .C(x2), .Y(ori_ori_n234_));
  OAI210     o218(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  OAI220     o219(.A0(ori_ori_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n236_));
  NO2        o220(.A(ori_ori_n229_), .B(ori_ori_n227_), .Y(ori_ori_n237_));
  AOI220     o221(.A0(ori_ori_n237_), .A1(ori_ori_n69_), .B0(ori_ori_n236_), .B1(ori_ori_n28_), .Y(ori_ori_n238_));
  AOI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n235_), .B0(ori_ori_n24_), .Y(ori_ori_n239_));
  NO2        o223(.A(ori_ori_n229_), .B(ori_ori_n227_), .Y(ori_ori_n240_));
  INV        o224(.A(ori_ori_n168_), .Y(ori_ori_n241_));
  NA2        o225(.A(ori_ori_n32_), .B(ori_ori_n37_), .Y(ori_ori_n242_));
  OR2        o226(.A(ori_ori_n242_), .B(ori_ori_n218_), .Y(ori_ori_n243_));
  OAI220     o227(.A0(ori_ori_n243_), .A1(ori_ori_n128_), .B0(ori_ori_n184_), .B1(ori_ori_n241_), .Y(ori_ori_n244_));
  AO210      o228(.A0(ori_ori_n240_), .A1(ori_ori_n118_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NO4        o229(.A(ori_ori_n245_), .B(ori_ori_n239_), .C(ori_ori_n232_), .D(ori_ori_n226_), .Y(ori_ori_n246_));
  OAI210     o230(.A0(ori_ori_n223_), .A1(ori_ori_n193_), .B0(ori_ori_n246_), .Y(ori04));
  NO2        o231(.A(x2), .B(x1), .Y(ori_ori_n248_));
  OAI210     o232(.A0(ori_ori_n200_), .A1(ori_ori_n248_), .B0(ori_ori_n32_), .Y(ori_ori_n249_));
  INV        o233(.A(ori_ori_n233_), .Y(ori_ori_n250_));
  OAI210     o234(.A0(ori_ori_n47_), .A1(ori_ori_n250_), .B0(ori_ori_n194_), .Y(ori_ori_n251_));
  NO2        o235(.A(ori_ori_n231_), .B(ori_ori_n164_), .Y(ori_ori_n252_));
  NA2        o236(.A(ori_ori_n252_), .B(ori_ori_n75_), .Y(ori_ori_n253_));
  NA3        o237(.A(ori_ori_n253_), .B(x6), .C(ori_ori_n251_), .Y(ori_ori_n254_));
  NA2        o238(.A(ori_ori_n254_), .B(ori_ori_n249_), .Y(ori_ori_n255_));
  OAI210     o239(.A0(ori_ori_n94_), .A1(ori_ori_n88_), .B0(ori_ori_n142_), .Y(ori_ori_n256_));
  NA3        o240(.A(ori_ori_n256_), .B(x6), .C(x3), .Y(ori_ori_n257_));
  AOI210     o241(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n258_));
  NO2        o242(.A(ori_ori_n258_), .B(ori_ori_n242_), .Y(ori_ori_n259_));
  INV        o243(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NA2        o244(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n261_));
  INV        o245(.A(ori_ori_n261_), .Y(ori_ori_n262_));
  NA2        o246(.A(ori_ori_n262_), .B(ori_ori_n66_), .Y(ori_ori_n263_));
  NA3        o247(.A(ori_ori_n263_), .B(ori_ori_n260_), .C(ori_ori_n257_), .Y(ori_ori_n264_));
  OAI210     o248(.A0(ori_ori_n92_), .A1(x3), .B0(ori_ori_n234_), .Y(ori_ori_n265_));
  NA2        o249(.A(ori_ori_n166_), .B(ori_ori_n70_), .Y(ori_ori_n266_));
  NA3        o250(.A(ori_ori_n266_), .B(ori_ori_n265_), .C(ori_ori_n120_), .Y(ori_ori_n267_));
  AOI210     o251(.A0(ori_ori_n264_), .A1(x4), .B0(ori_ori_n267_), .Y(ori_ori_n268_));
  NOi21      o252(.An(x4), .B(x0), .Y(ori_ori_n269_));
  XO2        o253(.A(x4), .B(x0), .Y(ori_ori_n270_));
  INV        o254(.A(ori_ori_n209_), .Y(ori_ori_n271_));
  AOI220     o255(.A0(ori_ori_n271_), .A1(x8), .B0(ori_ori_n269_), .B1(ori_ori_n76_), .Y(ori_ori_n272_));
  NO2        o256(.A(ori_ori_n272_), .B(x3), .Y(ori_ori_n273_));
  INV        o257(.A(ori_ori_n76_), .Y(ori_ori_n274_));
  NO2        o258(.A(ori_ori_n75_), .B(x4), .Y(ori_ori_n275_));
  AOI220     o259(.A0(ori_ori_n275_), .A1(ori_ori_n38_), .B0(ori_ori_n99_), .B1(ori_ori_n274_), .Y(ori_ori_n276_));
  NO2        o260(.A(ori_ori_n270_), .B(x2), .Y(ori_ori_n277_));
  INV        o261(.A(ori_ori_n277_), .Y(ori_ori_n278_));
  NA4        o262(.A(ori_ori_n278_), .B(ori_ori_n276_), .C(ori_ori_n175_), .D(x6), .Y(ori_ori_n279_));
  NO2        o263(.A(ori_ori_n144_), .B(ori_ori_n75_), .Y(ori_ori_n280_));
  NA2        o264(.A(ori_ori_n280_), .B(ori_ori_n54_), .Y(ori_ori_n281_));
  NO2        o265(.A(x8), .B(ori_ori_n68_), .Y(ori_ori_n282_));
  NO2        o266(.A(ori_ori_n31_), .B(x2), .Y(ori_ori_n283_));
  NA2        o267(.A(ori_ori_n283_), .B(ori_ori_n282_), .Y(ori_ori_n284_));
  NA2        o268(.A(ori_ori_n281_), .B(ori_ori_n284_), .Y(ori_ori_n285_));
  OAI220     o269(.A0(ori_ori_n285_), .A1(x6), .B0(ori_ori_n279_), .B1(ori_ori_n273_), .Y(ori_ori_n286_));
  NA2        o270(.A(ori_ori_n42_), .B(ori_ori_n36_), .Y(ori_ori_n287_));
  OAI210     o271(.A0(ori_ori_n287_), .A1(ori_ori_n75_), .B0(ori_ori_n243_), .Y(ori_ori_n288_));
  AOI210     o272(.A0(ori_ori_n288_), .A1(ori_ori_n18_), .B0(ori_ori_n120_), .Y(ori_ori_n289_));
  AO220      o273(.A0(ori_ori_n289_), .A1(ori_ori_n286_), .B0(ori_ori_n268_), .B1(ori_ori_n255_), .Y(ori_ori_n290_));
  NA2        o274(.A(ori_ori_n283_), .B(x6), .Y(ori_ori_n291_));
  AOI210     o275(.A0(x6), .A1(x1), .B0(ori_ori_n119_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n275_), .B(x0), .Y(ori_ori_n293_));
  NA2        o277(.A(ori_ori_n70_), .B(x6), .Y(ori_ori_n294_));
  OAI210     o278(.A0(ori_ori_n293_), .A1(ori_ori_n292_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  AOI220     o279(.A0(ori_ori_n295_), .A1(ori_ori_n291_), .B0(ori_ori_n169_), .B1(ori_ori_n43_), .Y(ori_ori_n296_));
  NA2        o280(.A(ori_ori_n296_), .B(ori_ori_n290_), .Y(ori_ori_n297_));
  INV        o281(.A(ori_ori_n92_), .Y(ori_ori_n298_));
  NA2        o282(.A(ori_ori_n298_), .B(ori_ori_n261_), .Y(ori_ori_n299_));
  NA3        o283(.A(ori_ori_n299_), .B(ori_ori_n160_), .C(ori_ori_n120_), .Y(ori_ori_n300_));
  NA3        o284(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n301_));
  NA2        o285(.A(ori_ori_n174_), .B(x0), .Y(ori_ori_n302_));
  OAI220     o286(.A0(ori_ori_n302_), .A1(x2), .B0(ori_ori_n301_), .B1(ori_ori_n274_), .Y(ori_ori_n303_));
  INV        o287(.A(ori_ori_n303_), .Y(ori_ori_n304_));
  AOI210     o288(.A0(ori_ori_n304_), .A1(ori_ori_n300_), .B0(ori_ori_n24_), .Y(ori_ori_n305_));
  NA2        o289(.A(ori_ori_n305_), .B(x6), .Y(ori_ori_n306_));
  NO2        o290(.A(ori_ori_n29_), .B(x0), .Y(ori_ori_n307_));
  NA2        o291(.A(ori_ori_n160_), .B(ori_ori_n120_), .Y(ori_ori_n308_));
  OAI210     o292(.A0(ori_ori_n308_), .A1(x8), .B0(ori_ori_n354_), .Y(ori_ori_n309_));
  NAi31      o293(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n310_));
  OAI210     o294(.A0(ori_ori_n310_), .A1(x4), .B0(ori_ori_n131_), .Y(ori_ori_n311_));
  NA3        o295(.A(ori_ori_n311_), .B(ori_ori_n117_), .C(x9), .Y(ori_ori_n312_));
  NA2        o296(.A(ori_ori_n282_), .B(ori_ori_n120_), .Y(ori_ori_n313_));
  NA4        o297(.A(ori_ori_n313_), .B(x1), .C(ori_ori_n312_), .D(ori_ori_n44_), .Y(ori_ori_n314_));
  OAI210     o298(.A0(ori_ori_n309_), .A1(ori_ori_n307_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  INV        o299(.A(ori_ori_n105_), .Y(ori_ori_n316_));
  NO2        o300(.A(ori_ori_n316_), .B(ori_ori_n37_), .Y(ori_ori_n317_));
  AOI210     o301(.A0(ori_ori_n209_), .A1(ori_ori_n53_), .B0(ori_ori_n98_), .Y(ori_ori_n318_));
  NO2        o302(.A(ori_ori_n318_), .B(x3), .Y(ori_ori_n319_));
  NO3        o303(.A(ori_ori_n319_), .B(ori_ori_n317_), .C(x2), .Y(ori_ori_n320_));
  OAI210     o304(.A0(ori_ori_n233_), .A1(ori_ori_n37_), .B0(ori_ori_n270_), .Y(ori_ori_n321_));
  INV        o305(.A(ori_ori_n301_), .Y(ori_ori_n322_));
  AOI220     o306(.A0(ori_ori_n322_), .A1(ori_ori_n75_), .B0(ori_ori_n321_), .B1(ori_ori_n120_), .Y(ori_ori_n323_));
  NO2        o307(.A(ori_ori_n323_), .B(ori_ori_n47_), .Y(ori_ori_n324_));
  NO2        o308(.A(ori_ori_n324_), .B(ori_ori_n320_), .Y(ori_ori_n325_));
  AOI210     o309(.A0(ori_ori_n325_), .A1(ori_ori_n315_), .B0(ori_ori_n24_), .Y(ori_ori_n326_));
  NA4        o310(.A(ori_ori_n28_), .B(ori_ori_n75_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n327_));
  NO3        o311(.A(ori_ori_n57_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n328_));
  NA2        o312(.A(ori_ori_n328_), .B(ori_ori_n210_), .Y(ori_ori_n329_));
  NO2        o313(.A(ori_ori_n329_), .B(ori_ori_n85_), .Y(ori_ori_n330_));
  NA2        o314(.A(ori_ori_n330_), .B(x7), .Y(ori_ori_n331_));
  INV        o315(.A(x7), .Y(ori_ori_n332_));
  NA3        o316(.A(ori_ori_n332_), .B(ori_ori_n119_), .C(ori_ori_n106_), .Y(ori_ori_n333_));
  NA3        o317(.A(ori_ori_n333_), .B(ori_ori_n331_), .C(ori_ori_n327_), .Y(ori_ori_n334_));
  OAI210     o318(.A0(ori_ori_n334_), .A1(ori_ori_n326_), .B0(ori_ori_n32_), .Y(ori_ori_n335_));
  INV        o319(.A(ori_ori_n164_), .Y(ori_ori_n336_));
  NO4        o320(.A(ori_ori_n336_), .B(ori_ori_n65_), .C(x4), .D(ori_ori_n47_), .Y(ori_ori_n337_));
  NA2        o321(.A(ori_ori_n200_), .B(ori_ori_n21_), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n128_), .B(ori_ori_n107_), .Y(ori_ori_n339_));
  NA2        o323(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  NO2        o324(.A(ori_ori_n340_), .B(ori_ori_n26_), .Y(ori_ori_n341_));
  NA2        o325(.A(ori_ori_n310_), .B(ori_ori_n73_), .Y(ori_ori_n342_));
  NA2        o326(.A(ori_ori_n342_), .B(ori_ori_n143_), .Y(ori_ori_n343_));
  OAI220     o327(.A0(x3), .A1(ori_ori_n58_), .B0(ori_ori_n128_), .B1(ori_ori_n37_), .Y(ori_ori_n344_));
  NA2        o328(.A(x3), .B(ori_ori_n47_), .Y(ori_ori_n345_));
  NO2        o329(.A(ori_ori_n121_), .B(ori_ori_n345_), .Y(ori_ori_n346_));
  AOI220     o330(.A0(ori_ori_n346_), .A1(x0), .B0(ori_ori_n344_), .B1(ori_ori_n107_), .Y(ori_ori_n347_));
  AOI210     o331(.A0(ori_ori_n347_), .A1(ori_ori_n343_), .B0(ori_ori_n184_), .Y(ori_ori_n348_));
  NO3        o332(.A(ori_ori_n348_), .B(ori_ori_n341_), .C(ori_ori_n337_), .Y(ori_ori_n349_));
  NA3        o333(.A(ori_ori_n349_), .B(ori_ori_n335_), .C(ori_ori_n306_), .Y(ori_ori_n350_));
  AOI210     o334(.A0(ori_ori_n297_), .A1(ori_ori_n24_), .B0(ori_ori_n350_), .Y(ori05));
  INV        o335(.A(x1), .Y(ori_ori_n354_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  INV        m047(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  NO3        m048(.A(mai_mai_n64_), .B(mai_mai_n61_), .C(mai_mai_n60_), .Y(mai_mai_n65_));
  NO2        m049(.A(x7), .B(x6), .Y(mai_mai_n66_));
  NO2        m050(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n67_));
  NO2        m051(.A(x8), .B(x2), .Y(mai_mai_n68_));
  OA210      m052(.A0(mai_mai_n68_), .A1(mai_mai_n67_), .B0(mai_mai_n66_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n70_), .Y(mai_mai_n71_));
  NAi31      m055(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n72_));
  NO2        m056(.A(mai_mai_n71_), .B(mai_mai_n69_), .Y(mai_mai_n73_));
  OAI210     m057(.A0(mai_mai_n73_), .A1(mai_mai_n65_), .B0(x4), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n75_));
  OAI210     m059(.A0(mai_mai_n75_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n76_));
  NA2        m060(.A(x5), .B(x3), .Y(mai_mai_n77_));
  NO2        m061(.A(x8), .B(x6), .Y(mai_mai_n78_));
  NO3        m062(.A(mai_mai_n78_), .B(mai_mai_n77_), .C(mai_mai_n54_), .Y(mai_mai_n79_));
  NAi21      m063(.An(x4), .B(x3), .Y(mai_mai_n80_));
  INV        m064(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m065(.A(mai_mai_n81_), .B(mai_mai_n22_), .Y(mai_mai_n82_));
  NO2        m066(.A(x4), .B(x2), .Y(mai_mai_n83_));
  NO2        m067(.A(mai_mai_n83_), .B(x3), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n82_), .C(mai_mai_n18_), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n79_), .C(mai_mai_n76_), .Y(mai_mai_n86_));
  NO3        m070(.A(mai_mai_n21_), .B(mai_mai_n43_), .C(x1), .Y(mai_mai_n87_));
  INV        m071(.A(x4), .Y(mai_mai_n88_));
  NA2        m072(.A(mai_mai_n87_), .B(mai_mai_n88_), .Y(mai_mai_n89_));
  NA2        m073(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n25_), .Y(mai_mai_n91_));
  INV        m075(.A(x8), .Y(mai_mai_n92_));
  NA2        m076(.A(x2), .B(x1), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n92_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n91_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n26_), .Y(mai_mai_n96_));
  AOI210     m080(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n97_));
  OAI210     m081(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n98_));
  NO3        m082(.A(mai_mai_n98_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n99_));
  NA2        m083(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n100_));
  NO2        m084(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n101_));
  OAI210     m085(.A0(mai_mai_n101_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n102_));
  AOI210     m086(.A0(mai_mai_n100_), .A1(mai_mai_n52_), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m087(.A(x3), .B(x2), .Y(mai_mai_n104_));
  NA2        m088(.A(mai_mai_n104_), .B(mai_mai_n25_), .Y(mai_mai_n105_));
  NO2        m089(.A(x6), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  NA2        m090(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n107_));
  OAI210     m091(.A0(mai_mai_n107_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n108_));
  NO4        m092(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n103_), .D(mai_mai_n99_), .Y(mai_mai_n109_));
  AO220      m093(.A0(mai_mai_n109_), .A1(mai_mai_n89_), .B0(mai_mai_n86_), .B1(mai_mai_n74_), .Y(mai02));
  NO2        m094(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n111_));
  NO2        m095(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n112_));
  NA2        m096(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n113_));
  AOI220     m097(.A0(mai_mai_n54_), .A1(mai_mai_n112_), .B0(mai_mai_n111_), .B1(x4), .Y(mai_mai_n114_));
  NO3        m098(.A(mai_mai_n114_), .B(x7), .C(x5), .Y(mai_mai_n115_));
  NA2        m099(.A(x9), .B(x2), .Y(mai_mai_n116_));
  OR2        m100(.A(x8), .B(x0), .Y(mai_mai_n117_));
  INV        m101(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NAi21      m102(.An(x2), .B(x8), .Y(mai_mai_n119_));
  NO2        m103(.A(x4), .B(x1), .Y(mai_mai_n120_));
  NOi21      m104(.An(x0), .B(x1), .Y(mai_mai_n121_));
  NO3        m105(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n122_));
  NOi21      m106(.An(x0), .B(x4), .Y(mai_mai_n123_));
  NO2        m107(.A(x8), .B(mai_mai_n62_), .Y(mai_mai_n124_));
  AOI220     m108(.A0(mai_mai_n124_), .A1(mai_mai_n123_), .B0(mai_mai_n122_), .B1(mai_mai_n121_), .Y(mai_mai_n125_));
  NO2        m109(.A(mai_mai_n125_), .B(mai_mai_n77_), .Y(mai_mai_n126_));
  NO2        m110(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n127_));
  NA2        m111(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n128_));
  AOI210     m112(.A0(mai_mai_n128_), .A1(mai_mai_n107_), .B0(mai_mai_n113_), .Y(mai_mai_n129_));
  OAI210     m113(.A0(mai_mai_n129_), .A1(mai_mai_n35_), .B0(mai_mai_n127_), .Y(mai_mai_n130_));
  NAi21      m114(.An(x0), .B(x4), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n131_), .B(x1), .Y(mai_mai_n132_));
  NO2        m116(.A(x7), .B(x0), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n83_), .B(mai_mai_n101_), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n134_), .B(x3), .Y(mai_mai_n135_));
  OAI210     m119(.A0(mai_mai_n133_), .A1(mai_mai_n132_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NO2        m120(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n137_));
  NA2        m121(.A(x5), .B(x0), .Y(mai_mai_n138_));
  NO2        m122(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n139_));
  NA3        m123(.A(mai_mai_n139_), .B(mai_mai_n138_), .C(mai_mai_n137_), .Y(mai_mai_n140_));
  NA4        m124(.A(mai_mai_n140_), .B(mai_mai_n136_), .C(mai_mai_n130_), .D(mai_mai_n36_), .Y(mai_mai_n141_));
  NO3        m125(.A(mai_mai_n141_), .B(mai_mai_n126_), .C(mai_mai_n115_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n143_));
  AOI220     m127(.A0(mai_mai_n121_), .A1(mai_mai_n143_), .B0(mai_mai_n67_), .B1(mai_mai_n17_), .Y(mai_mai_n144_));
  NO3        m128(.A(mai_mai_n144_), .B(mai_mai_n60_), .C(mai_mai_n62_), .Y(mai_mai_n145_));
  NO2        m129(.A(mai_mai_n100_), .B(x5), .Y(mai_mai_n146_));
  NO2        m130(.A(x9), .B(x7), .Y(mai_mai_n147_));
  NOi21      m131(.An(x8), .B(x0), .Y(mai_mai_n148_));
  NO2        m132(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n149_));
  INV        m133(.A(x7), .Y(mai_mai_n150_));
  NA2        m134(.A(mai_mai_n150_), .B(mai_mai_n18_), .Y(mai_mai_n151_));
  AOI220     m135(.A0(mai_mai_n151_), .A1(mai_mai_n149_), .B0(mai_mai_n111_), .B1(mai_mai_n38_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n153_), .B(mai_mai_n123_), .Y(mai_mai_n154_));
  NO2        m138(.A(mai_mai_n154_), .B(mai_mai_n152_), .Y(mai_mai_n155_));
  AOI210     m139(.A0(mai_mai_n148_), .A1(mai_mai_n146_), .B0(mai_mai_n155_), .Y(mai_mai_n156_));
  INV        m140(.A(mai_mai_n156_), .Y(mai_mai_n157_));
  NA2        m141(.A(x5), .B(x1), .Y(mai_mai_n158_));
  INV        m142(.A(mai_mai_n158_), .Y(mai_mai_n159_));
  AOI210     m143(.A0(mai_mai_n159_), .A1(mai_mai_n123_), .B0(mai_mai_n36_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n62_), .B(mai_mai_n92_), .Y(mai_mai_n161_));
  NO3        m145(.A(x2), .B(mai_mai_n161_), .C(mai_mai_n48_), .Y(mai_mai_n162_));
  NA2        m146(.A(mai_mai_n162_), .B(mai_mai_n67_), .Y(mai_mai_n163_));
  NAi31      m147(.An(mai_mai_n77_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n164_));
  NA3        m148(.A(mai_mai_n164_), .B(mai_mai_n163_), .C(mai_mai_n160_), .Y(mai_mai_n165_));
  NO3        m149(.A(mai_mai_n165_), .B(mai_mai_n157_), .C(mai_mai_n145_), .Y(mai_mai_n166_));
  NO2        m150(.A(mai_mai_n166_), .B(mai_mai_n142_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n138_), .B(mai_mai_n134_), .Y(mai_mai_n168_));
  NA2        m152(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n169_));
  NA2        m153(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n170_));
  NA3        m154(.A(mai_mai_n170_), .B(mai_mai_n169_), .C(mai_mai_n24_), .Y(mai_mai_n171_));
  AN2        m155(.A(mai_mai_n171_), .B(mai_mai_n139_), .Y(mai_mai_n172_));
  NA2        m156(.A(x8), .B(x0), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n150_), .B(mai_mai_n25_), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n121_), .B(x4), .Y(mai_mai_n175_));
  NA2        m159(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  AOI210     m160(.A0(mai_mai_n173_), .A1(mai_mai_n128_), .B0(mai_mai_n176_), .Y(mai_mai_n177_));
  NA2        m161(.A(x2), .B(x0), .Y(mai_mai_n178_));
  NA2        m162(.A(x4), .B(x1), .Y(mai_mai_n179_));
  NAi21      m163(.An(mai_mai_n120_), .B(mai_mai_n179_), .Y(mai_mai_n180_));
  NOi31      m164(.An(mai_mai_n180_), .B(mai_mai_n153_), .C(mai_mai_n178_), .Y(mai_mai_n181_));
  NO4        m165(.A(mai_mai_n181_), .B(mai_mai_n177_), .C(mai_mai_n172_), .D(mai_mai_n168_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n182_), .B(mai_mai_n43_), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n171_), .B(mai_mai_n75_), .Y(mai_mai_n184_));
  INV        m168(.A(mai_mai_n127_), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n107_), .B(mai_mai_n17_), .Y(mai_mai_n186_));
  NA3        m170(.A(mai_mai_n180_), .B(mai_mai_n185_), .C(mai_mai_n42_), .Y(mai_mai_n187_));
  OAI210     m171(.A0(mai_mai_n170_), .A1(mai_mai_n134_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  NO2        m172(.A(mai_mai_n188_), .B(mai_mai_n184_), .Y(mai_mai_n189_));
  NO2        m173(.A(mai_mai_n189_), .B(x3), .Y(mai_mai_n190_));
  NO3        m174(.A(mai_mai_n190_), .B(mai_mai_n183_), .C(mai_mai_n167_), .Y(mai03));
  NO2        m175(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n192_));
  NO2        m176(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n193_));
  INV        m177(.A(mai_mai_n193_), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n195_));
  OAI210     m179(.A0(mai_mai_n195_), .A1(mai_mai_n25_), .B0(mai_mai_n63_), .Y(mai_mai_n196_));
  OAI220     m180(.A0(mai_mai_n196_), .A1(mai_mai_n17_), .B0(mai_mai_n194_), .B1(mai_mai_n107_), .Y(mai_mai_n197_));
  NA2        m181(.A(mai_mai_n197_), .B(mai_mai_n192_), .Y(mai_mai_n198_));
  NO2        m182(.A(mai_mai_n77_), .B(x6), .Y(mai_mai_n199_));
  NA2        m183(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n200_));
  NO2        m184(.A(mai_mai_n200_), .B(x4), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n202_));
  AN2        m186(.A(mai_mai_n199_), .B(mai_mai_n55_), .Y(mai_mai_n203_));
  NA2        m187(.A(mai_mai_n203_), .B(mai_mai_n62_), .Y(mai_mai_n204_));
  NA2        m188(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n205_), .B(mai_mai_n200_), .Y(mai_mai_n206_));
  NA2        m190(.A(x9), .B(mai_mai_n54_), .Y(mai_mai_n207_));
  NA2        m191(.A(mai_mai_n207_), .B(x4), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n200_), .B(mai_mai_n80_), .Y(mai_mai_n209_));
  AOI210     m193(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n178_), .Y(mai_mai_n210_));
  AOI220     m194(.A0(mai_mai_n210_), .A1(mai_mai_n209_), .B0(mai_mai_n208_), .B1(mai_mai_n206_), .Y(mai_mai_n211_));
  NO2        m195(.A(x5), .B(x1), .Y(mai_mai_n212_));
  AOI220     m196(.A0(mai_mai_n212_), .A1(mai_mai_n17_), .B0(mai_mai_n104_), .B1(x5), .Y(mai_mai_n213_));
  NO2        m197(.A(mai_mai_n205_), .B(mai_mai_n169_), .Y(mai_mai_n214_));
  INV        m198(.A(mai_mai_n214_), .Y(mai_mai_n215_));
  OAI210     m199(.A0(mai_mai_n213_), .A1(mai_mai_n64_), .B0(mai_mai_n215_), .Y(mai_mai_n216_));
  NA2        m200(.A(mai_mai_n216_), .B(mai_mai_n48_), .Y(mai_mai_n217_));
  NA4        m201(.A(mai_mai_n217_), .B(mai_mai_n211_), .C(mai_mai_n204_), .D(mai_mai_n198_), .Y(mai_mai_n218_));
  NO2        m202(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n219_));
  NA2        m203(.A(mai_mai_n219_), .B(mai_mai_n19_), .Y(mai_mai_n220_));
  NO2        m204(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n221_), .B(x6), .Y(mai_mai_n222_));
  NOi21      m206(.An(mai_mai_n83_), .B(mai_mai_n222_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n62_), .B(mai_mai_n92_), .Y(mai_mai_n224_));
  NO2        m208(.A(mai_mai_n223_), .B(mai_mai_n150_), .Y(mai_mai_n225_));
  AO210      m209(.A0(mai_mai_n225_), .A1(mai_mai_n220_), .B0(mai_mai_n174_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n227_));
  NO3        m211(.A(mai_mai_n179_), .B(mai_mai_n62_), .C(x6), .Y(mai_mai_n228_));
  AOI220     m212(.A0(mai_mai_n228_), .A1(mai_mai_n17_), .B0(mai_mai_n139_), .B1(mai_mai_n91_), .Y(mai_mai_n229_));
  NA2        m213(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n230_));
  NO2        m214(.A(mai_mai_n230_), .B(mai_mai_n77_), .Y(mai_mai_n231_));
  NO2        m215(.A(mai_mai_n158_), .B(mai_mai_n43_), .Y(mai_mai_n232_));
  OAI210     m216(.A0(mai_mai_n232_), .A1(mai_mai_n214_), .B0(mai_mai_n436_), .Y(mai_mai_n233_));
  NA2        m217(.A(mai_mai_n193_), .B(mai_mai_n132_), .Y(mai_mai_n234_));
  OAI210     m218(.A0(mai_mai_n92_), .A1(mai_mai_n36_), .B0(mai_mai_n67_), .Y(mai_mai_n235_));
  NA3        m219(.A(mai_mai_n235_), .B(mai_mai_n234_), .C(mai_mai_n233_), .Y(mai_mai_n236_));
  OAI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n231_), .B0(x2), .Y(mai_mai_n237_));
  NA3        m221(.A(mai_mai_n237_), .B(mai_mai_n229_), .C(mai_mai_n226_), .Y(mai_mai_n238_));
  AOI210     m222(.A0(mai_mai_n218_), .A1(x8), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NO2        m223(.A(mai_mai_n92_), .B(x3), .Y(mai_mai_n240_));
  NO3        m224(.A(mai_mai_n90_), .B(mai_mai_n78_), .C(mai_mai_n25_), .Y(mai_mai_n241_));
  AOI210     m225(.A0(mai_mai_n222_), .A1(mai_mai_n153_), .B0(mai_mai_n241_), .Y(mai_mai_n242_));
  NO2        m226(.A(mai_mai_n242_), .B(x2), .Y(mai_mai_n243_));
  NO2        m227(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n244_));
  AOI220     m228(.A0(mai_mai_n201_), .A1(mai_mai_n186_), .B0(mai_mai_n244_), .B1(mai_mai_n67_), .Y(mai_mai_n245_));
  NA2        m229(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n246_));
  NA3        m230(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n247_));
  AOI210     m231(.A0(mai_mai_n247_), .A1(mai_mai_n138_), .B0(mai_mai_n246_), .Y(mai_mai_n248_));
  NA2        m232(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n249_));
  NO2        m233(.A(mai_mai_n249_), .B(mai_mai_n25_), .Y(mai_mai_n250_));
  OAI210     m234(.A0(mai_mai_n250_), .A1(mai_mai_n248_), .B0(mai_mai_n120_), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n205_), .B(x6), .Y(mai_mai_n252_));
  NO2        m236(.A(mai_mai_n205_), .B(x6), .Y(mai_mai_n253_));
  NA2        m237(.A(mai_mai_n252_), .B(mai_mai_n143_), .Y(mai_mai_n254_));
  NA4        m238(.A(mai_mai_n254_), .B(mai_mai_n251_), .C(mai_mai_n245_), .D(mai_mai_n150_), .Y(mai_mai_n255_));
  NA2        m239(.A(mai_mai_n193_), .B(mai_mai_n221_), .Y(mai_mai_n256_));
  NO2        m240(.A(x9), .B(x6), .Y(mai_mai_n257_));
  NO2        m241(.A(mai_mai_n138_), .B(mai_mai_n18_), .Y(mai_mai_n258_));
  NAi21      m242(.An(mai_mai_n258_), .B(mai_mai_n247_), .Y(mai_mai_n259_));
  NAi21      m243(.An(x1), .B(x4), .Y(mai_mai_n260_));
  AOI220     m244(.A0(mai_mai_n48_), .A1(mai_mai_n260_), .B0(mai_mai_n259_), .B1(mai_mai_n257_), .Y(mai_mai_n261_));
  NA2        m245(.A(mai_mai_n261_), .B(mai_mai_n256_), .Y(mai_mai_n262_));
  NA2        m246(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n263_));
  NO2        m247(.A(mai_mai_n263_), .B(mai_mai_n256_), .Y(mai_mai_n264_));
  NO3        m248(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n265_));
  NA2        m249(.A(mai_mai_n107_), .B(mai_mai_n25_), .Y(mai_mai_n266_));
  NA2        m250(.A(x6), .B(x2), .Y(mai_mai_n267_));
  NO2        m251(.A(mai_mai_n267_), .B(mai_mai_n169_), .Y(mai_mai_n268_));
  AOI210     m252(.A0(mai_mai_n266_), .A1(mai_mai_n265_), .B0(mai_mai_n268_), .Y(mai_mai_n269_));
  OAI220     m253(.A0(mai_mai_n269_), .A1(mai_mai_n43_), .B0(mai_mai_n175_), .B1(mai_mai_n46_), .Y(mai_mai_n270_));
  OAI210     m254(.A0(mai_mai_n270_), .A1(mai_mai_n264_), .B0(mai_mai_n262_), .Y(mai_mai_n271_));
  NA2        m255(.A(x4), .B(x0), .Y(mai_mai_n272_));
  NA2        m256(.A(mai_mai_n199_), .B(mai_mai_n42_), .Y(mai_mai_n273_));
  AOI210     m257(.A0(mai_mai_n273_), .A1(mai_mai_n271_), .B0(x8), .Y(mai_mai_n274_));
  OAI210     m258(.A0(mai_mai_n258_), .A1(mai_mai_n212_), .B0(x6), .Y(mai_mai_n275_));
  INV        m259(.A(mai_mai_n173_), .Y(mai_mai_n276_));
  OAI210     m260(.A0(mai_mai_n276_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n277_));
  AOI210     m261(.A0(mai_mai_n277_), .A1(mai_mai_n275_), .B0(mai_mai_n227_), .Y(mai_mai_n278_));
  NO4        m262(.A(mai_mai_n278_), .B(mai_mai_n274_), .C(mai_mai_n255_), .D(mai_mai_n243_), .Y(mai_mai_n279_));
  NO2        m263(.A(mai_mai_n161_), .B(x1), .Y(mai_mai_n280_));
  NO2        m264(.A(x3), .B(mai_mai_n36_), .Y(mai_mai_n281_));
  OAI210     m265(.A0(mai_mai_n281_), .A1(mai_mai_n253_), .B0(x2), .Y(mai_mai_n282_));
  OAI210     m266(.A0(mai_mai_n276_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n283_));
  AOI210     m267(.A0(mai_mai_n283_), .A1(mai_mai_n282_), .B0(mai_mai_n185_), .Y(mai_mai_n284_));
  NOi21      m268(.An(mai_mai_n267_), .B(mai_mai_n17_), .Y(mai_mai_n285_));
  NA3        m269(.A(mai_mai_n285_), .B(mai_mai_n212_), .C(mai_mai_n40_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n287_));
  NA3        m271(.A(mai_mai_n287_), .B(mai_mai_n159_), .C(mai_mai_n32_), .Y(mai_mai_n288_));
  NA2        m272(.A(x3), .B(x2), .Y(mai_mai_n289_));
  AOI220     m273(.A0(mai_mai_n289_), .A1(mai_mai_n227_), .B0(mai_mai_n288_), .B1(mai_mai_n286_), .Y(mai_mai_n290_));
  NAi21      m274(.An(x4), .B(x0), .Y(mai_mai_n291_));
  NO3        m275(.A(mai_mai_n291_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n292_));
  OAI210     m276(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n292_), .Y(mai_mai_n293_));
  OAI220     m277(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n294_));
  NA2        m278(.A(mai_mai_n36_), .B(mai_mai_n54_), .Y(mai_mai_n295_));
  OAI210     m279(.A0(mai_mai_n287_), .A1(mai_mai_n285_), .B0(mai_mai_n295_), .Y(mai_mai_n296_));
  AOI220     m280(.A0(mai_mai_n296_), .A1(mai_mai_n81_), .B0(mai_mai_n294_), .B1(mai_mai_n31_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n297_), .A1(mai_mai_n293_), .B0(mai_mai_n25_), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n299_));
  OAI210     m283(.A0(mai_mai_n287_), .A1(mai_mai_n285_), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  INV        m284(.A(mai_mai_n214_), .Y(mai_mai_n301_));
  NA2        m285(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n302_));
  OR2        m286(.A(mai_mai_n302_), .B(mai_mai_n272_), .Y(mai_mai_n303_));
  OAI220     m287(.A0(mai_mai_n303_), .A1(mai_mai_n158_), .B0(mai_mai_n230_), .B1(mai_mai_n301_), .Y(mai_mai_n304_));
  AO210      m288(.A0(mai_mai_n300_), .A1(mai_mai_n146_), .B0(mai_mai_n304_), .Y(mai_mai_n305_));
  NO4        m289(.A(mai_mai_n305_), .B(mai_mai_n298_), .C(mai_mai_n290_), .D(mai_mai_n284_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n279_), .A1(mai_mai_n239_), .B0(mai_mai_n306_), .Y(mai04));
  OAI210     m291(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n308_));
  NA3        m292(.A(mai_mai_n308_), .B(mai_mai_n265_), .C(mai_mai_n84_), .Y(mai_mai_n309_));
  NO2        m293(.A(x2), .B(x1), .Y(mai_mai_n310_));
  OAI210     m294(.A0(mai_mai_n249_), .A1(mai_mai_n310_), .B0(mai_mai_n36_), .Y(mai_mai_n311_));
  NO2        m295(.A(mai_mai_n310_), .B(mai_mai_n291_), .Y(mai_mai_n312_));
  NA2        m296(.A(mai_mai_n312_), .B(mai_mai_n240_), .Y(mai_mai_n313_));
  NO2        m297(.A(mai_mai_n263_), .B(mai_mai_n90_), .Y(mai_mai_n314_));
  NO2        m298(.A(mai_mai_n314_), .B(mai_mai_n36_), .Y(mai_mai_n315_));
  NO2        m299(.A(mai_mai_n289_), .B(mai_mai_n202_), .Y(mai_mai_n316_));
  NA2        m300(.A(x9), .B(x0), .Y(mai_mai_n317_));
  AOI210     m301(.A0(mai_mai_n90_), .A1(mai_mai_n75_), .B0(mai_mai_n317_), .Y(mai_mai_n318_));
  OAI210     m302(.A0(mai_mai_n318_), .A1(mai_mai_n316_), .B0(mai_mai_n92_), .Y(mai_mai_n319_));
  NA3        m303(.A(mai_mai_n319_), .B(mai_mai_n315_), .C(mai_mai_n313_), .Y(mai_mai_n320_));
  NA2        m304(.A(mai_mai_n320_), .B(mai_mai_n311_), .Y(mai_mai_n321_));
  NO2        m305(.A(mai_mai_n207_), .B(mai_mai_n113_), .Y(mai_mai_n322_));
  INV        m306(.A(mai_mai_n322_), .Y(mai_mai_n323_));
  OAI210     m307(.A0(mai_mai_n117_), .A1(mai_mai_n107_), .B0(mai_mai_n173_), .Y(mai_mai_n324_));
  NA3        m308(.A(mai_mai_n324_), .B(x6), .C(x3), .Y(mai_mai_n325_));
  NOi21      m309(.An(mai_mai_n148_), .B(mai_mai_n128_), .Y(mai_mai_n326_));
  AOI210     m310(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n327_));
  OAI220     m311(.A0(mai_mai_n327_), .A1(mai_mai_n302_), .B0(mai_mai_n263_), .B1(mai_mai_n299_), .Y(mai_mai_n328_));
  AOI210     m312(.A0(mai_mai_n326_), .A1(mai_mai_n63_), .B0(mai_mai_n328_), .Y(mai_mai_n329_));
  NO2        m313(.A(mai_mai_n107_), .B(mai_mai_n17_), .Y(mai_mai_n330_));
  AOI220     m314(.A0(mai_mai_n330_), .A1(mai_mai_n78_), .B0(mai_mai_n314_), .B1(mai_mai_n92_), .Y(mai_mai_n331_));
  NA4        m315(.A(mai_mai_n331_), .B(mai_mai_n329_), .C(mai_mai_n325_), .D(mai_mai_n323_), .Y(mai_mai_n332_));
  OAI210     m316(.A0(mai_mai_n112_), .A1(x3), .B0(mai_mai_n292_), .Y(mai_mai_n333_));
  NA2        m317(.A(mai_mai_n333_), .B(mai_mai_n150_), .Y(mai_mai_n334_));
  AOI210     m318(.A0(mai_mai_n332_), .A1(x4), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  NA3        m319(.A(mai_mai_n312_), .B(mai_mai_n207_), .C(mai_mai_n92_), .Y(mai_mai_n336_));
  NOi21      m320(.An(x4), .B(x0), .Y(mai_mai_n337_));
  XO2        m321(.A(x4), .B(x0), .Y(mai_mai_n338_));
  OAI210     m322(.A0(mai_mai_n338_), .A1(mai_mai_n116_), .B0(mai_mai_n260_), .Y(mai_mai_n339_));
  AOI220     m323(.A0(mai_mai_n339_), .A1(x8), .B0(mai_mai_n337_), .B1(mai_mai_n93_), .Y(mai_mai_n340_));
  AOI210     m324(.A0(mai_mai_n340_), .A1(mai_mai_n336_), .B0(x3), .Y(mai_mai_n341_));
  INV        m325(.A(mai_mai_n93_), .Y(mai_mai_n342_));
  NO2        m326(.A(mai_mai_n92_), .B(x4), .Y(mai_mai_n343_));
  AOI220     m327(.A0(mai_mai_n343_), .A1(mai_mai_n44_), .B0(mai_mai_n123_), .B1(mai_mai_n342_), .Y(mai_mai_n344_));
  NO3        m328(.A(mai_mai_n338_), .B(mai_mai_n161_), .C(x2), .Y(mai_mai_n345_));
  NO3        m329(.A(mai_mai_n224_), .B(mai_mai_n28_), .C(mai_mai_n24_), .Y(mai_mai_n346_));
  NO2        m330(.A(mai_mai_n346_), .B(mai_mai_n345_), .Y(mai_mai_n347_));
  NA4        m331(.A(mai_mai_n347_), .B(mai_mai_n344_), .C(mai_mai_n220_), .D(x6), .Y(mai_mai_n348_));
  OAI220     m332(.A0(mai_mai_n291_), .A1(mai_mai_n90_), .B0(mai_mai_n178_), .B1(mai_mai_n92_), .Y(mai_mai_n349_));
  NO2        m333(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n350_));
  OR2        m334(.A(mai_mai_n343_), .B(mai_mai_n350_), .Y(mai_mai_n351_));
  NO2        m335(.A(mai_mai_n148_), .B(mai_mai_n107_), .Y(mai_mai_n352_));
  AOI220     m336(.A0(mai_mai_n352_), .A1(mai_mai_n351_), .B0(mai_mai_n349_), .B1(mai_mai_n61_), .Y(mai_mai_n353_));
  NO2        m337(.A(mai_mai_n148_), .B(mai_mai_n80_), .Y(mai_mai_n354_));
  NO2        m338(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n355_));
  NOi21      m339(.An(mai_mai_n120_), .B(mai_mai_n27_), .Y(mai_mai_n356_));
  AOI210     m340(.A0(mai_mai_n355_), .A1(mai_mai_n354_), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  OAI210     m341(.A0(mai_mai_n353_), .A1(mai_mai_n62_), .B0(mai_mai_n357_), .Y(mai_mai_n358_));
  OAI220     m342(.A0(mai_mai_n358_), .A1(x6), .B0(mai_mai_n348_), .B1(mai_mai_n341_), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n63_), .A1(mai_mai_n48_), .B0(mai_mai_n42_), .Y(mai_mai_n360_));
  OAI210     m344(.A0(mai_mai_n360_), .A1(mai_mai_n92_), .B0(mai_mai_n303_), .Y(mai_mai_n361_));
  AOI210     m345(.A0(mai_mai_n361_), .A1(mai_mai_n18_), .B0(mai_mai_n150_), .Y(mai_mai_n362_));
  AO220      m346(.A0(mai_mai_n362_), .A1(mai_mai_n359_), .B0(mai_mai_n335_), .B1(mai_mai_n321_), .Y(mai_mai_n363_));
  NA2        m347(.A(mai_mai_n83_), .B(x6), .Y(mai_mai_n364_));
  NA2        m348(.A(mai_mai_n435_), .B(mai_mai_n35_), .Y(mai_mai_n365_));
  NA3        m349(.A(mai_mai_n365_), .B(mai_mai_n363_), .C(mai_mai_n309_), .Y(mai_mai_n366_));
  AOI210     m350(.A0(mai_mai_n195_), .A1(x8), .B0(mai_mai_n112_), .Y(mai_mai_n367_));
  INV        m351(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  NA3        m352(.A(mai_mai_n368_), .B(mai_mai_n192_), .C(mai_mai_n150_), .Y(mai_mai_n369_));
  AO220      m353(.A0(x4), .A1(mai_mai_n147_), .B0(mai_mai_n111_), .B1(x4), .Y(mai_mai_n370_));
  NA3        m354(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n371_));
  NO2        m355(.A(mai_mai_n371_), .B(mai_mai_n342_), .Y(mai_mai_n372_));
  AOI210     m356(.A0(mai_mai_n370_), .A1(mai_mai_n118_), .B0(mai_mai_n372_), .Y(mai_mai_n373_));
  AOI210     m357(.A0(mai_mai_n373_), .A1(mai_mai_n369_), .B0(mai_mai_n25_), .Y(mai_mai_n374_));
  OAI210     m358(.A0(mai_mai_n192_), .A1(mai_mai_n68_), .B0(mai_mai_n202_), .Y(mai_mai_n375_));
  NA3        m359(.A(mai_mai_n195_), .B(mai_mai_n221_), .C(x8), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n376_), .A1(mai_mai_n375_), .B0(mai_mai_n25_), .Y(mai_mai_n377_));
  AOI210     m361(.A0(mai_mai_n119_), .A1(mai_mai_n117_), .B0(mai_mai_n42_), .Y(mai_mai_n378_));
  NOi31      m362(.An(mai_mai_n378_), .B(mai_mai_n350_), .C(mai_mai_n179_), .Y(mai_mai_n379_));
  OAI210     m363(.A0(mai_mai_n379_), .A1(mai_mai_n377_), .B0(mai_mai_n147_), .Y(mai_mai_n380_));
  NAi31      m364(.An(mai_mai_n50_), .B(mai_mai_n280_), .C(mai_mai_n174_), .Y(mai_mai_n381_));
  NA2        m365(.A(mai_mai_n381_), .B(mai_mai_n380_), .Y(mai_mai_n382_));
  OAI210     m366(.A0(mai_mai_n382_), .A1(mai_mai_n374_), .B0(x6), .Y(mai_mai_n383_));
  INV        m367(.A(mai_mai_n133_), .Y(mai_mai_n384_));
  NA3        m368(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n385_));
  AOI220     m369(.A0(mai_mai_n385_), .A1(mai_mai_n384_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n386_));
  AOI220     m370(.A0(mai_mai_n437_), .A1(mai_mai_n219_), .B0(mai_mai_n192_), .B1(mai_mai_n150_), .Y(mai_mai_n387_));
  AOI210     m371(.A0(mai_mai_n124_), .A1(mai_mai_n244_), .B0(x1), .Y(mai_mai_n388_));
  OAI210     m372(.A0(mai_mai_n387_), .A1(x8), .B0(mai_mai_n388_), .Y(mai_mai_n389_));
  NO4        m373(.A(x8), .B(mai_mai_n291_), .C(x9), .D(x2), .Y(mai_mai_n390_));
  NOi21      m374(.An(mai_mai_n122_), .B(mai_mai_n178_), .Y(mai_mai_n391_));
  NO3        m375(.A(mai_mai_n391_), .B(mai_mai_n390_), .C(mai_mai_n18_), .Y(mai_mai_n392_));
  NO3        m376(.A(x9), .B(mai_mai_n150_), .C(x0), .Y(mai_mai_n393_));
  AOI220     m377(.A0(mai_mai_n393_), .A1(mai_mai_n240_), .B0(mai_mai_n354_), .B1(mai_mai_n150_), .Y(mai_mai_n394_));
  NA3        m378(.A(mai_mai_n394_), .B(mai_mai_n392_), .C(mai_mai_n50_), .Y(mai_mai_n395_));
  OAI210     m379(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n395_), .Y(mai_mai_n396_));
  NOi31      m380(.An(mai_mai_n437_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n397_));
  AOI210     m381(.A0(mai_mai_n38_), .A1(x9), .B0(mai_mai_n131_), .Y(mai_mai_n398_));
  NO3        m382(.A(mai_mai_n398_), .B(mai_mai_n122_), .C(mai_mai_n43_), .Y(mai_mai_n399_));
  NOi31      m383(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n400_));
  AOI220     m384(.A0(mai_mai_n400_), .A1(mai_mai_n337_), .B0(mai_mai_n123_), .B1(x3), .Y(mai_mai_n401_));
  AOI210     m385(.A0(mai_mai_n260_), .A1(mai_mai_n60_), .B0(mai_mai_n121_), .Y(mai_mai_n402_));
  OAI210     m386(.A0(mai_mai_n402_), .A1(x3), .B0(mai_mai_n401_), .Y(mai_mai_n403_));
  NO3        m387(.A(mai_mai_n403_), .B(mai_mai_n399_), .C(x2), .Y(mai_mai_n404_));
  NO2        m388(.A(mai_mai_n404_), .B(mai_mai_n397_), .Y(mai_mai_n405_));
  AOI210     m389(.A0(mai_mai_n405_), .A1(mai_mai_n396_), .B0(mai_mai_n25_), .Y(mai_mai_n406_));
  NA2        m390(.A(mai_mai_n438_), .B(mai_mai_n378_), .Y(mai_mai_n407_));
  NO2        m391(.A(mai_mai_n407_), .B(mai_mai_n104_), .Y(mai_mai_n408_));
  NO3        m392(.A(mai_mai_n263_), .B(mai_mai_n173_), .C(mai_mai_n40_), .Y(mai_mai_n409_));
  OAI210     m393(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(x7), .Y(mai_mai_n410_));
  NA2        m394(.A(mai_mai_n224_), .B(x7), .Y(mai_mai_n411_));
  NA3        m395(.A(mai_mai_n411_), .B(mai_mai_n149_), .C(mai_mai_n132_), .Y(mai_mai_n412_));
  NA2        m396(.A(mai_mai_n412_), .B(mai_mai_n410_), .Y(mai_mai_n413_));
  OAI210     m397(.A0(mai_mai_n413_), .A1(mai_mai_n406_), .B0(mai_mai_n36_), .Y(mai_mai_n414_));
  NO2        m398(.A(mai_mai_n393_), .B(mai_mai_n202_), .Y(mai_mai_n415_));
  NO4        m399(.A(mai_mai_n415_), .B(mai_mai_n77_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n416_));
  NO2        m400(.A(mai_mai_n164_), .B(mai_mai_n28_), .Y(mai_mai_n417_));
  AOI220     m401(.A0(mai_mai_n350_), .A1(mai_mai_n92_), .B0(mai_mai_n148_), .B1(mai_mai_n195_), .Y(mai_mai_n418_));
  NA2        m402(.A(mai_mai_n418_), .B(mai_mai_n90_), .Y(mai_mai_n419_));
  NA2        m403(.A(mai_mai_n419_), .B(mai_mai_n174_), .Y(mai_mai_n420_));
  AOI210     m404(.A0(x2), .A1(mai_mai_n27_), .B0(mai_mai_n72_), .Y(mai_mai_n421_));
  OAI210     m405(.A0(mai_mai_n147_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n422_));
  NO3        m406(.A(mai_mai_n400_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n423_));
  AOI210     m407(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n421_), .Y(mai_mai_n424_));
  INV        m408(.A(mai_mai_n424_), .Y(mai_mai_n425_));
  NA2        m409(.A(mai_mai_n425_), .B(x0), .Y(mai_mai_n426_));
  AOI210     m410(.A0(mai_mai_n426_), .A1(mai_mai_n420_), .B0(mai_mai_n230_), .Y(mai_mai_n427_));
  INV        m411(.A(x5), .Y(mai_mai_n428_));
  NO4        m412(.A(mai_mai_n107_), .B(mai_mai_n428_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n429_));
  NO4        m413(.A(mai_mai_n429_), .B(mai_mai_n427_), .C(mai_mai_n417_), .D(mai_mai_n416_), .Y(mai_mai_n430_));
  NA3        m414(.A(mai_mai_n430_), .B(mai_mai_n414_), .C(mai_mai_n383_), .Y(mai_mai_n431_));
  AOI210     m415(.A0(mai_mai_n366_), .A1(mai_mai_n25_), .B0(mai_mai_n431_), .Y(mai05));
  INV        m416(.A(mai_mai_n364_), .Y(mai_mai_n435_));
  INV        m417(.A(x6), .Y(mai_mai_n436_));
  INV        m418(.A(x0), .Y(mai_mai_n437_));
  INV        m419(.A(x4), .Y(mai_mai_n438_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO3        u012(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n63_));
  INV        u047(.A(men_men_n63_), .Y(men_men_n64_));
  NO3        u048(.A(men_men_n64_), .B(men_men_n61_), .C(men_men_n60_), .Y(men_men_n65_));
  NO2        u049(.A(x7), .B(x6), .Y(men_men_n66_));
  NO2        u050(.A(men_men_n61_), .B(x5), .Y(men_men_n67_));
  NO2        u051(.A(x8), .B(x2), .Y(men_men_n68_));
  INV        u052(.A(men_men_n68_), .Y(men_men_n69_));
  NO2        u053(.A(men_men_n69_), .B(x1), .Y(men_men_n70_));
  OA210      u054(.A0(men_men_n70_), .A1(men_men_n67_), .B0(men_men_n66_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n72_), .Y(men_men_n73_));
  NAi31      u057(.An(x1), .B(x9), .C(x5), .Y(men_men_n74_));
  OAI220     u058(.A0(men_men_n74_), .A1(men_men_n43_), .B0(men_men_n73_), .B1(men_men_n71_), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n65_), .B0(x4), .Y(men_men_n76_));
  NA2        u060(.A(men_men_n48_), .B(x2), .Y(men_men_n77_));
  OAI210     u061(.A0(men_men_n77_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n78_));
  NA2        u062(.A(x5), .B(x3), .Y(men_men_n79_));
  NO2        u063(.A(x8), .B(x6), .Y(men_men_n80_));
  NO4        u064(.A(men_men_n80_), .B(men_men_n79_), .C(men_men_n66_), .D(men_men_n54_), .Y(men_men_n81_));
  NAi21      u065(.An(x4), .B(x3), .Y(men_men_n82_));
  INV        u066(.A(men_men_n82_), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(men_men_n22_), .Y(men_men_n84_));
  NO2        u068(.A(x4), .B(x2), .Y(men_men_n85_));
  NO2        u069(.A(men_men_n85_), .B(x3), .Y(men_men_n86_));
  NO3        u070(.A(men_men_n86_), .B(men_men_n84_), .C(men_men_n18_), .Y(men_men_n87_));
  NO3        u071(.A(men_men_n87_), .B(men_men_n81_), .C(men_men_n78_), .Y(men_men_n88_));
  NO4        u072(.A(men_men_n21_), .B(x6), .C(men_men_n43_), .D(x1), .Y(men_men_n89_));
  NA2        u073(.A(men_men_n62_), .B(men_men_n48_), .Y(men_men_n90_));
  INV        u074(.A(men_men_n90_), .Y(men_men_n91_));
  OAI210     u075(.A0(men_men_n89_), .A1(men_men_n67_), .B0(men_men_n91_), .Y(men_men_n92_));
  NA2        u076(.A(x3), .B(men_men_n18_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n25_), .Y(men_men_n94_));
  INV        u078(.A(x8), .Y(men_men_n95_));
  NA2        u079(.A(x2), .B(x1), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n26_), .Y(men_men_n97_));
  AOI210     u081(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n98_));
  OAI210     u082(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n99_));
  NO3        u083(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n100_));
  NA2        u084(.A(x4), .B(men_men_n43_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n102_));
  AOI210     u086(.A0(men_men_n101_), .A1(men_men_n52_), .B0(x1), .Y(men_men_n103_));
  NO2        u087(.A(x3), .B(x2), .Y(men_men_n104_));
  NA2        u088(.A(men_men_n104_), .B(men_men_n25_), .Y(men_men_n105_));
  AOI210     u089(.A0(x8), .A1(x6), .B0(men_men_n105_), .Y(men_men_n106_));
  NA2        u090(.A(men_men_n54_), .B(x1), .Y(men_men_n107_));
  OAI210     u091(.A0(men_men_n107_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n108_));
  NO4        u092(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n103_), .D(men_men_n100_), .Y(men_men_n109_));
  AO220      u093(.A0(men_men_n109_), .A1(men_men_n92_), .B0(men_men_n88_), .B1(men_men_n76_), .Y(men02));
  NO2        u094(.A(x3), .B(men_men_n54_), .Y(men_men_n111_));
  NA2        u095(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n43_), .B(x0), .Y(men_men_n113_));
  OAI210     u097(.A0(men_men_n90_), .A1(men_men_n112_), .B0(men_men_n113_), .Y(men_men_n114_));
  NA2        u098(.A(men_men_n114_), .B(x1), .Y(men_men_n115_));
  NO3        u099(.A(men_men_n115_), .B(x7), .C(x5), .Y(men_men_n116_));
  NA2        u100(.A(x9), .B(x2), .Y(men_men_n117_));
  OR2        u101(.A(x8), .B(x0), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  NAi21      u103(.An(x2), .B(x8), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  OAI220     u105(.A0(men_men_n121_), .A1(men_men_n119_), .B0(men_men_n117_), .B1(x7), .Y(men_men_n122_));
  NO2        u106(.A(x4), .B(x1), .Y(men_men_n123_));
  NA3        u107(.A(men_men_n123_), .B(men_men_n122_), .C(men_men_n60_), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x1), .Y(men_men_n125_));
  NO3        u109(.A(x9), .B(x8), .C(x7), .Y(men_men_n126_));
  NOi21      u110(.An(x0), .B(x4), .Y(men_men_n127_));
  NAi21      u111(.An(x8), .B(x7), .Y(men_men_n128_));
  NO2        u112(.A(men_men_n128_), .B(men_men_n62_), .Y(men_men_n129_));
  AOI220     u113(.A0(men_men_n129_), .A1(men_men_n127_), .B0(men_men_n126_), .B1(men_men_n125_), .Y(men_men_n130_));
  AOI210     u114(.A0(men_men_n130_), .A1(men_men_n124_), .B0(men_men_n79_), .Y(men_men_n131_));
  NO2        u115(.A(x5), .B(men_men_n48_), .Y(men_men_n132_));
  NA2        u116(.A(x2), .B(men_men_n18_), .Y(men_men_n133_));
  AOI210     u117(.A0(men_men_n133_), .A1(men_men_n107_), .B0(men_men_n113_), .Y(men_men_n134_));
  OAI210     u118(.A0(men_men_n134_), .A1(men_men_n35_), .B0(men_men_n132_), .Y(men_men_n135_));
  NAi21      u119(.An(x0), .B(x4), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n136_), .B(x1), .Y(men_men_n137_));
  NO2        u121(.A(x7), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n85_), .B(men_men_n102_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n139_), .B(x3), .Y(men_men_n140_));
  OAI210     u124(.A0(men_men_n138_), .A1(men_men_n137_), .B0(men_men_n140_), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n21_), .B(men_men_n43_), .Y(men_men_n142_));
  NA2        u126(.A(x5), .B(x0), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n48_), .B(x2), .Y(men_men_n144_));
  NA3        u128(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n142_), .Y(men_men_n145_));
  NA4        u129(.A(men_men_n145_), .B(men_men_n141_), .C(men_men_n135_), .D(men_men_n36_), .Y(men_men_n146_));
  NO3        u130(.A(men_men_n146_), .B(men_men_n131_), .C(men_men_n116_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n79_), .B(men_men_n77_), .C(men_men_n24_), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n149_));
  AOI220     u133(.A0(men_men_n125_), .A1(men_men_n149_), .B0(men_men_n67_), .B1(men_men_n17_), .Y(men_men_n150_));
  NO3        u134(.A(men_men_n150_), .B(men_men_n60_), .C(men_men_n62_), .Y(men_men_n151_));
  NA2        u135(.A(x7), .B(x3), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n101_), .B(x5), .Y(men_men_n153_));
  NO2        u137(.A(x9), .B(x7), .Y(men_men_n154_));
  NOi21      u138(.An(x8), .B(x0), .Y(men_men_n155_));
  OA210      u139(.A0(men_men_n154_), .A1(x1), .B0(men_men_n155_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n43_), .B(x2), .Y(men_men_n157_));
  INV        u141(.A(x7), .Y(men_men_n158_));
  NA2        u142(.A(men_men_n158_), .B(men_men_n18_), .Y(men_men_n159_));
  AOI220     u143(.A0(men_men_n159_), .A1(men_men_n157_), .B0(men_men_n111_), .B1(men_men_n38_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n25_), .B(x4), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n161_), .B(men_men_n127_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n160_), .Y(men_men_n163_));
  AOI210     u147(.A0(men_men_n156_), .A1(men_men_n153_), .B0(men_men_n163_), .Y(men_men_n164_));
  OAI210     u148(.A0(men_men_n152_), .A1(men_men_n50_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u149(.A(x5), .B(x1), .Y(men_men_n166_));
  INV        u150(.A(men_men_n166_), .Y(men_men_n167_));
  AOI210     u151(.A0(men_men_n167_), .A1(men_men_n127_), .B0(men_men_n36_), .Y(men_men_n168_));
  NO2        u152(.A(men_men_n62_), .B(men_men_n95_), .Y(men_men_n169_));
  NAi21      u153(.An(x2), .B(x7), .Y(men_men_n170_));
  NAi31      u154(.An(men_men_n79_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n171_), .B(men_men_n168_), .Y(men_men_n172_));
  NO4        u156(.A(men_men_n172_), .B(men_men_n165_), .C(men_men_n151_), .D(men_men_n148_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n173_), .B(men_men_n147_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n143_), .B(men_men_n139_), .Y(men_men_n175_));
  NA2        u159(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n176_));
  NA2        u160(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n177_));
  NA3        u161(.A(men_men_n177_), .B(men_men_n176_), .C(men_men_n24_), .Y(men_men_n178_));
  AN2        u162(.A(men_men_n178_), .B(men_men_n144_), .Y(men_men_n179_));
  NA2        u163(.A(x8), .B(x0), .Y(men_men_n180_));
  NO2        u164(.A(men_men_n158_), .B(men_men_n25_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n125_), .B(x4), .Y(men_men_n182_));
  NA2        u166(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  AOI210     u167(.A0(men_men_n180_), .A1(men_men_n133_), .B0(men_men_n183_), .Y(men_men_n184_));
  NA2        u168(.A(x2), .B(x0), .Y(men_men_n185_));
  NA2        u169(.A(x4), .B(x1), .Y(men_men_n186_));
  NAi21      u170(.An(men_men_n123_), .B(men_men_n186_), .Y(men_men_n187_));
  NOi31      u171(.An(men_men_n187_), .B(men_men_n161_), .C(men_men_n185_), .Y(men_men_n188_));
  NO4        u172(.A(men_men_n188_), .B(men_men_n184_), .C(men_men_n179_), .D(men_men_n175_), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n189_), .B(men_men_n43_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n178_), .B(men_men_n77_), .Y(men_men_n191_));
  INV        u175(.A(men_men_n132_), .Y(men_men_n192_));
  NO2        u176(.A(men_men_n107_), .B(men_men_n17_), .Y(men_men_n193_));
  AOI210     u177(.A0(men_men_n35_), .A1(men_men_n95_), .B0(men_men_n193_), .Y(men_men_n194_));
  NO3        u178(.A(men_men_n194_), .B(men_men_n192_), .C(x7), .Y(men_men_n195_));
  NA3        u179(.A(men_men_n187_), .B(men_men_n192_), .C(men_men_n42_), .Y(men_men_n196_));
  OAI210     u180(.A0(men_men_n177_), .A1(men_men_n139_), .B0(men_men_n196_), .Y(men_men_n197_));
  NO3        u181(.A(men_men_n197_), .B(men_men_n195_), .C(men_men_n191_), .Y(men_men_n198_));
  NO2        u182(.A(men_men_n198_), .B(x3), .Y(men_men_n199_));
  NO3        u183(.A(men_men_n199_), .B(men_men_n190_), .C(men_men_n174_), .Y(men03));
  NO2        u184(.A(men_men_n48_), .B(x3), .Y(men_men_n201_));
  NO2        u185(.A(x6), .B(men_men_n25_), .Y(men_men_n202_));
  NO2        u186(.A(men_men_n54_), .B(x1), .Y(men_men_n203_));
  OAI210     u187(.A0(men_men_n203_), .A1(men_men_n25_), .B0(men_men_n63_), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n204_), .B(men_men_n17_), .Y(men_men_n205_));
  NA2        u189(.A(men_men_n205_), .B(men_men_n201_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n79_), .B(x6), .Y(men_men_n207_));
  NA2        u191(.A(x6), .B(men_men_n25_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n208_), .B(x4), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n18_), .B(x0), .Y(men_men_n210_));
  AO220      u194(.A0(men_men_n210_), .A1(men_men_n209_), .B0(men_men_n207_), .B1(men_men_n55_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n211_), .B(men_men_n62_), .Y(men_men_n212_));
  NA2        u196(.A(x3), .B(men_men_n17_), .Y(men_men_n213_));
  NO2        u197(.A(men_men_n213_), .B(men_men_n208_), .Y(men_men_n214_));
  NA2        u198(.A(x9), .B(men_men_n54_), .Y(men_men_n215_));
  NA2        u199(.A(men_men_n208_), .B(men_men_n82_), .Y(men_men_n216_));
  AOI210     u200(.A0(men_men_n25_), .A1(x3), .B0(men_men_n185_), .Y(men_men_n217_));
  AOI220     u201(.A0(men_men_n217_), .A1(men_men_n216_), .B0(x9), .B1(men_men_n214_), .Y(men_men_n218_));
  NO3        u202(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n219_));
  NO2        u203(.A(x5), .B(x1), .Y(men_men_n220_));
  AOI220     u204(.A0(men_men_n220_), .A1(men_men_n17_), .B0(men_men_n104_), .B1(x5), .Y(men_men_n221_));
  NO2        u205(.A(men_men_n213_), .B(men_men_n176_), .Y(men_men_n222_));
  NO3        u206(.A(x3), .B(x2), .C(x1), .Y(men_men_n223_));
  NO2        u207(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  OAI210     u208(.A0(men_men_n221_), .A1(men_men_n64_), .B0(men_men_n224_), .Y(men_men_n225_));
  NA2        u209(.A(men_men_n225_), .B(men_men_n48_), .Y(men_men_n226_));
  NA4        u210(.A(men_men_n226_), .B(men_men_n218_), .C(men_men_n212_), .D(men_men_n206_), .Y(men_men_n227_));
  NO2        u211(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n228_));
  NA2        u212(.A(men_men_n228_), .B(men_men_n19_), .Y(men_men_n229_));
  NO2        u213(.A(x3), .B(men_men_n17_), .Y(men_men_n230_));
  NO2        u214(.A(men_men_n230_), .B(x6), .Y(men_men_n231_));
  NOi21      u215(.An(men_men_n85_), .B(men_men_n231_), .Y(men_men_n232_));
  NA2        u216(.A(men_men_n62_), .B(men_men_n95_), .Y(men_men_n233_));
  NA3        u217(.A(men_men_n233_), .B(men_men_n230_), .C(x6), .Y(men_men_n234_));
  AOI210     u218(.A0(men_men_n234_), .A1(men_men_n232_), .B0(men_men_n158_), .Y(men_men_n235_));
  AO210      u219(.A0(men_men_n235_), .A1(men_men_n229_), .B0(men_men_n181_), .Y(men_men_n236_));
  NA2        u220(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n237_));
  OAI210     u221(.A0(men_men_n237_), .A1(men_men_n25_), .B0(men_men_n177_), .Y(men_men_n238_));
  NO2        u222(.A(men_men_n186_), .B(x6), .Y(men_men_n239_));
  AOI220     u223(.A0(men_men_n239_), .A1(men_men_n238_), .B0(men_men_n144_), .B1(men_men_n94_), .Y(men_men_n240_));
  NA2        u224(.A(x6), .B(men_men_n48_), .Y(men_men_n241_));
  OAI210     u225(.A0(men_men_n119_), .A1(men_men_n80_), .B0(x4), .Y(men_men_n242_));
  AOI210     u226(.A0(men_men_n242_), .A1(men_men_n241_), .B0(men_men_n79_), .Y(men_men_n243_));
  NO2        u227(.A(men_men_n166_), .B(men_men_n43_), .Y(men_men_n244_));
  OAI210     u228(.A0(men_men_n244_), .A1(men_men_n222_), .B0(x9), .Y(men_men_n245_));
  NA2        u229(.A(men_men_n202_), .B(men_men_n137_), .Y(men_men_n246_));
  NA3        u230(.A(men_men_n213_), .B(men_men_n132_), .C(x6), .Y(men_men_n247_));
  OAI210     u231(.A0(men_men_n95_), .A1(men_men_n36_), .B0(men_men_n67_), .Y(men_men_n248_));
  NA4        u232(.A(men_men_n248_), .B(men_men_n247_), .C(men_men_n246_), .D(men_men_n245_), .Y(men_men_n249_));
  OAI210     u233(.A0(men_men_n249_), .A1(men_men_n243_), .B0(x2), .Y(men_men_n250_));
  NA3        u234(.A(men_men_n250_), .B(men_men_n240_), .C(men_men_n236_), .Y(men_men_n251_));
  AOI210     u235(.A0(men_men_n227_), .A1(x8), .B0(men_men_n251_), .Y(men_men_n252_));
  NO2        u236(.A(men_men_n95_), .B(x3), .Y(men_men_n253_));
  NA2        u237(.A(men_men_n253_), .B(men_men_n209_), .Y(men_men_n254_));
  NO3        u238(.A(men_men_n93_), .B(men_men_n80_), .C(men_men_n25_), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n231_), .A1(men_men_n161_), .B0(men_men_n255_), .Y(men_men_n256_));
  AOI210     u240(.A0(men_men_n256_), .A1(men_men_n254_), .B0(x2), .Y(men_men_n257_));
  NO2        u241(.A(x4), .B(men_men_n54_), .Y(men_men_n258_));
  AOI220     u242(.A0(men_men_n209_), .A1(men_men_n193_), .B0(men_men_n258_), .B1(men_men_n67_), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n62_), .B(x6), .Y(men_men_n260_));
  NA3        u244(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n261_));
  NO2        u245(.A(men_men_n261_), .B(men_men_n260_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n263_));
  NA2        u247(.A(men_men_n262_), .B(men_men_n123_), .Y(men_men_n264_));
  NA2        u248(.A(men_men_n213_), .B(x6), .Y(men_men_n265_));
  NO2        u249(.A(men_men_n213_), .B(x6), .Y(men_men_n266_));
  NAi21      u250(.An(men_men_n169_), .B(men_men_n266_), .Y(men_men_n267_));
  NA3        u251(.A(men_men_n267_), .B(men_men_n265_), .C(men_men_n149_), .Y(men_men_n268_));
  NA4        u252(.A(men_men_n268_), .B(men_men_n264_), .C(men_men_n259_), .D(men_men_n158_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n202_), .B(men_men_n230_), .Y(men_men_n270_));
  NO2        u254(.A(x9), .B(x6), .Y(men_men_n271_));
  NO2        u255(.A(men_men_n143_), .B(men_men_n18_), .Y(men_men_n272_));
  NAi21      u256(.An(men_men_n272_), .B(men_men_n261_), .Y(men_men_n273_));
  NAi21      u257(.An(x1), .B(x4), .Y(men_men_n274_));
  AOI210     u258(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n275_));
  OAI210     u259(.A0(men_men_n143_), .A1(x3), .B0(men_men_n275_), .Y(men_men_n276_));
  AOI220     u260(.A0(men_men_n276_), .A1(men_men_n274_), .B0(men_men_n273_), .B1(men_men_n271_), .Y(men_men_n277_));
  INV        u261(.A(men_men_n277_), .Y(men_men_n278_));
  NA2        u262(.A(men_men_n62_), .B(x2), .Y(men_men_n279_));
  NO2        u263(.A(men_men_n279_), .B(men_men_n270_), .Y(men_men_n280_));
  NO3        u264(.A(x9), .B(x6), .C(x0), .Y(men_men_n281_));
  NA2        u265(.A(x6), .B(x2), .Y(men_men_n282_));
  NO2        u266(.A(men_men_n282_), .B(men_men_n176_), .Y(men_men_n283_));
  NO2        u267(.A(men_men_n281_), .B(men_men_n283_), .Y(men_men_n284_));
  OAI220     u268(.A0(men_men_n284_), .A1(men_men_n43_), .B0(men_men_n182_), .B1(men_men_n46_), .Y(men_men_n285_));
  OAI210     u269(.A0(men_men_n285_), .A1(men_men_n280_), .B0(men_men_n278_), .Y(men_men_n286_));
  NO2        u270(.A(men_men_n453_), .B(men_men_n208_), .Y(men_men_n287_));
  OR3        u271(.A(men_men_n287_), .B(men_men_n207_), .C(men_men_n153_), .Y(men_men_n288_));
  NA2        u272(.A(x4), .B(x0), .Y(men_men_n289_));
  NO3        u273(.A(men_men_n74_), .B(men_men_n289_), .C(x6), .Y(men_men_n290_));
  AOI210     u274(.A0(men_men_n288_), .A1(men_men_n42_), .B0(men_men_n290_), .Y(men_men_n291_));
  AOI210     u275(.A0(men_men_n291_), .A1(men_men_n286_), .B0(x8), .Y(men_men_n292_));
  INV        u276(.A(men_men_n260_), .Y(men_men_n293_));
  OAI210     u277(.A0(men_men_n272_), .A1(men_men_n220_), .B0(men_men_n293_), .Y(men_men_n294_));
  INV        u278(.A(men_men_n180_), .Y(men_men_n295_));
  NO2        u279(.A(men_men_n294_), .B(men_men_n237_), .Y(men_men_n296_));
  NO4        u280(.A(men_men_n296_), .B(men_men_n292_), .C(men_men_n269_), .D(men_men_n257_), .Y(men_men_n297_));
  NO2        u281(.A(men_men_n169_), .B(x1), .Y(men_men_n298_));
  NO3        u282(.A(men_men_n298_), .B(x3), .C(men_men_n36_), .Y(men_men_n299_));
  OAI210     u283(.A0(men_men_n299_), .A1(men_men_n266_), .B0(x2), .Y(men_men_n300_));
  OAI210     u284(.A0(men_men_n295_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n301_));
  AOI210     u285(.A0(men_men_n301_), .A1(men_men_n300_), .B0(men_men_n192_), .Y(men_men_n302_));
  NOi21      u286(.An(men_men_n282_), .B(men_men_n17_), .Y(men_men_n303_));
  NA3        u287(.A(men_men_n303_), .B(men_men_n220_), .C(men_men_n40_), .Y(men_men_n304_));
  AOI210     u288(.A0(men_men_n36_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n305_));
  NA3        u289(.A(men_men_n305_), .B(men_men_n167_), .C(men_men_n32_), .Y(men_men_n306_));
  NA2        u290(.A(x3), .B(x2), .Y(men_men_n307_));
  AOI220     u291(.A0(men_men_n307_), .A1(men_men_n237_), .B0(men_men_n306_), .B1(men_men_n304_), .Y(men_men_n308_));
  NAi21      u292(.An(x4), .B(x0), .Y(men_men_n309_));
  NO3        u293(.A(men_men_n309_), .B(men_men_n44_), .C(x2), .Y(men_men_n310_));
  OAI210     u294(.A0(x6), .A1(men_men_n18_), .B0(men_men_n310_), .Y(men_men_n311_));
  NO2        u295(.A(x9), .B(x8), .Y(men_men_n312_));
  NA3        u296(.A(men_men_n312_), .B(men_men_n36_), .C(men_men_n54_), .Y(men_men_n313_));
  OAI210     u297(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n313_), .Y(men_men_n314_));
  AOI220     u298(.A0(men_men_n314_), .A1(men_men_n83_), .B0(men_men_n18_), .B1(men_men_n31_), .Y(men_men_n315_));
  AOI210     u299(.A0(men_men_n315_), .A1(men_men_n311_), .B0(men_men_n25_), .Y(men_men_n316_));
  NA3        u300(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n317_));
  OAI210     u301(.A0(men_men_n305_), .A1(men_men_n303_), .B0(men_men_n317_), .Y(men_men_n318_));
  AN2        u302(.A(men_men_n318_), .B(men_men_n153_), .Y(men_men_n319_));
  NO4        u303(.A(men_men_n319_), .B(men_men_n316_), .C(men_men_n308_), .D(men_men_n302_), .Y(men_men_n320_));
  OAI210     u304(.A0(men_men_n297_), .A1(men_men_n252_), .B0(men_men_n320_), .Y(men04));
  OAI210     u305(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n322_));
  NA3        u306(.A(men_men_n322_), .B(men_men_n281_), .C(men_men_n86_), .Y(men_men_n323_));
  NO2        u307(.A(x2), .B(x1), .Y(men_men_n324_));
  OAI210     u308(.A0(men_men_n263_), .A1(men_men_n324_), .B0(men_men_n36_), .Y(men_men_n325_));
  NO2        u309(.A(men_men_n324_), .B(men_men_n309_), .Y(men_men_n326_));
  AOI210     u310(.A0(men_men_n62_), .A1(x4), .B0(men_men_n112_), .Y(men_men_n327_));
  NA2        u311(.A(men_men_n327_), .B(men_men_n253_), .Y(men_men_n328_));
  NA3        u312(.A(men_men_n93_), .B(x6), .C(men_men_n328_), .Y(men_men_n329_));
  NA2        u313(.A(men_men_n329_), .B(men_men_n325_), .Y(men_men_n330_));
  NO2        u314(.A(men_men_n215_), .B(men_men_n113_), .Y(men_men_n331_));
  NO3        u315(.A(men_men_n260_), .B(men_men_n120_), .C(men_men_n18_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n332_), .B(men_men_n331_), .Y(men_men_n333_));
  NO2        u317(.A(men_men_n279_), .B(men_men_n317_), .Y(men_men_n334_));
  AOI210     u318(.A0(men_men_n18_), .A1(men_men_n63_), .B0(men_men_n334_), .Y(men_men_n335_));
  NA3        u319(.A(men_men_n452_), .B(men_men_n335_), .C(men_men_n333_), .Y(men_men_n336_));
  OAI210     u320(.A0(x1), .A1(x3), .B0(men_men_n310_), .Y(men_men_n337_));
  NA3        u321(.A(men_men_n233_), .B(men_men_n219_), .C(men_men_n85_), .Y(men_men_n338_));
  NA3        u322(.A(men_men_n338_), .B(men_men_n337_), .C(men_men_n158_), .Y(men_men_n339_));
  AOI210     u323(.A0(men_men_n336_), .A1(x4), .B0(men_men_n339_), .Y(men_men_n340_));
  NA2        u324(.A(men_men_n326_), .B(men_men_n95_), .Y(men_men_n341_));
  NOi21      u325(.An(x4), .B(x0), .Y(men_men_n342_));
  XO2        u326(.A(x4), .B(x0), .Y(men_men_n343_));
  NA2        u327(.A(men_men_n117_), .B(men_men_n274_), .Y(men_men_n344_));
  AOI220     u328(.A0(men_men_n344_), .A1(x8), .B0(men_men_n342_), .B1(men_men_n96_), .Y(men_men_n345_));
  AOI210     u329(.A0(men_men_n345_), .A1(men_men_n341_), .B0(x3), .Y(men_men_n346_));
  NO2        u330(.A(men_men_n95_), .B(x4), .Y(men_men_n347_));
  NA2        u331(.A(men_men_n347_), .B(men_men_n44_), .Y(men_men_n348_));
  NO3        u332(.A(men_men_n343_), .B(men_men_n169_), .C(x2), .Y(men_men_n349_));
  NO3        u333(.A(men_men_n233_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n350_));
  NO2        u334(.A(men_men_n350_), .B(men_men_n349_), .Y(men_men_n351_));
  NA4        u335(.A(men_men_n351_), .B(men_men_n348_), .C(men_men_n229_), .D(x6), .Y(men_men_n352_));
  NO2        u336(.A(men_men_n43_), .B(x0), .Y(men_men_n353_));
  OR2        u337(.A(men_men_n347_), .B(men_men_n353_), .Y(men_men_n354_));
  NO2        u338(.A(men_men_n155_), .B(men_men_n107_), .Y(men_men_n355_));
  AOI220     u339(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n451_), .B1(men_men_n61_), .Y(men_men_n356_));
  NO2        u340(.A(men_men_n155_), .B(men_men_n82_), .Y(men_men_n357_));
  NO2        u341(.A(men_men_n35_), .B(x2), .Y(men_men_n358_));
  NOi21      u342(.An(men_men_n123_), .B(men_men_n27_), .Y(men_men_n359_));
  AOI210     u343(.A0(men_men_n358_), .A1(men_men_n357_), .B0(men_men_n359_), .Y(men_men_n360_));
  OAI210     u344(.A0(men_men_n356_), .A1(men_men_n62_), .B0(men_men_n360_), .Y(men_men_n361_));
  OAI220     u345(.A0(men_men_n361_), .A1(x6), .B0(men_men_n352_), .B1(men_men_n346_), .Y(men_men_n362_));
  OAI210     u346(.A0(men_men_n63_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n363_), .B(men_men_n95_), .Y(men_men_n364_));
  AOI210     u348(.A0(men_men_n364_), .A1(men_men_n18_), .B0(men_men_n158_), .Y(men_men_n365_));
  AO220      u349(.A0(men_men_n365_), .A1(men_men_n362_), .B0(men_men_n340_), .B1(men_men_n330_), .Y(men_men_n366_));
  NA2        u350(.A(men_men_n358_), .B(x6), .Y(men_men_n367_));
  AOI210     u351(.A0(x6), .A1(x1), .B0(men_men_n157_), .Y(men_men_n368_));
  NA2        u352(.A(men_men_n347_), .B(x0), .Y(men_men_n369_));
  NO2        u353(.A(men_men_n369_), .B(men_men_n368_), .Y(men_men_n370_));
  AOI220     u354(.A0(men_men_n370_), .A1(men_men_n367_), .B0(men_men_n223_), .B1(men_men_n49_), .Y(men_men_n371_));
  NA3        u355(.A(men_men_n371_), .B(men_men_n366_), .C(men_men_n323_), .Y(men_men_n372_));
  NA3        u356(.A(x2), .B(men_men_n201_), .C(men_men_n158_), .Y(men_men_n373_));
  OAI210     u357(.A0(men_men_n28_), .A1(x1), .B0(men_men_n237_), .Y(men_men_n374_));
  AO220      u358(.A0(men_men_n374_), .A1(men_men_n154_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n375_));
  NA3        u359(.A(x7), .B(x3), .C(x0), .Y(men_men_n376_));
  NA2        u360(.A(men_men_n228_), .B(x0), .Y(men_men_n377_));
  OAI220     u361(.A0(men_men_n377_), .A1(men_men_n215_), .B0(men_men_n376_), .B1(x2), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n375_), .A1(men_men_n119_), .B0(men_men_n378_), .Y(men_men_n379_));
  AOI210     u363(.A0(men_men_n379_), .A1(men_men_n373_), .B0(men_men_n25_), .Y(men_men_n380_));
  NA3        u364(.A(men_men_n121_), .B(men_men_n228_), .C(x0), .Y(men_men_n381_));
  OAI210     u365(.A0(men_men_n201_), .A1(men_men_n68_), .B0(men_men_n210_), .Y(men_men_n382_));
  NO2        u366(.A(men_men_n382_), .B(men_men_n25_), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n120_), .A1(men_men_n118_), .B0(men_men_n42_), .Y(men_men_n384_));
  NOi31      u368(.An(men_men_n384_), .B(men_men_n353_), .C(men_men_n186_), .Y(men_men_n385_));
  OAI210     u369(.A0(men_men_n385_), .A1(men_men_n383_), .B0(men_men_n154_), .Y(men_men_n386_));
  NAi31      u370(.An(men_men_n50_), .B(men_men_n298_), .C(men_men_n181_), .Y(men_men_n387_));
  NA3        u371(.A(men_men_n387_), .B(men_men_n386_), .C(men_men_n381_), .Y(men_men_n388_));
  OAI210     u372(.A0(men_men_n388_), .A1(men_men_n380_), .B0(x6), .Y(men_men_n389_));
  OAI210     u373(.A0(men_men_n169_), .A1(men_men_n48_), .B0(men_men_n138_), .Y(men_men_n390_));
  NA3        u374(.A(men_men_n55_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n391_));
  AOI220     u375(.A0(men_men_n391_), .A1(men_men_n390_), .B0(men_men_n40_), .B1(men_men_n32_), .Y(men_men_n392_));
  NO2        u376(.A(men_men_n158_), .B(x0), .Y(men_men_n393_));
  AOI220     u377(.A0(men_men_n393_), .A1(men_men_n228_), .B0(men_men_n201_), .B1(men_men_n158_), .Y(men_men_n394_));
  AOI210     u378(.A0(men_men_n129_), .A1(men_men_n258_), .B0(x1), .Y(men_men_n395_));
  OAI210     u379(.A0(men_men_n394_), .A1(x8), .B0(men_men_n395_), .Y(men_men_n396_));
  NAi31      u380(.An(x2), .B(x8), .C(x0), .Y(men_men_n397_));
  OAI210     u381(.A0(men_men_n397_), .A1(x4), .B0(men_men_n170_), .Y(men_men_n398_));
  NA3        u382(.A(men_men_n398_), .B(men_men_n152_), .C(x9), .Y(men_men_n399_));
  NO4        u383(.A(men_men_n128_), .B(men_men_n309_), .C(x9), .D(x2), .Y(men_men_n400_));
  NOi21      u384(.An(men_men_n126_), .B(men_men_n185_), .Y(men_men_n401_));
  NO3        u385(.A(men_men_n401_), .B(men_men_n400_), .C(men_men_n18_), .Y(men_men_n402_));
  NO3        u386(.A(x9), .B(men_men_n158_), .C(x0), .Y(men_men_n403_));
  AOI220     u387(.A0(men_men_n403_), .A1(men_men_n253_), .B0(men_men_n357_), .B1(men_men_n158_), .Y(men_men_n404_));
  NA4        u388(.A(men_men_n404_), .B(men_men_n402_), .C(men_men_n399_), .D(men_men_n50_), .Y(men_men_n405_));
  OAI210     u389(.A0(men_men_n396_), .A1(men_men_n392_), .B0(men_men_n405_), .Y(men_men_n406_));
  NOi31      u390(.An(men_men_n393_), .B(men_men_n32_), .C(x8), .Y(men_men_n407_));
  NO2        u391(.A(men_men_n126_), .B(men_men_n43_), .Y(men_men_n408_));
  AOI210     u392(.A0(men_men_n127_), .A1(x3), .B0(men_men_n342_), .Y(men_men_n409_));
  NA2        u393(.A(x3), .B(men_men_n409_), .Y(men_men_n410_));
  NO3        u394(.A(men_men_n410_), .B(men_men_n408_), .C(x2), .Y(men_men_n411_));
  OAI220     u395(.A0(men_men_n343_), .A1(men_men_n312_), .B0(men_men_n309_), .B1(men_men_n43_), .Y(men_men_n412_));
  AOI210     u396(.A0(x9), .A1(men_men_n48_), .B0(men_men_n376_), .Y(men_men_n413_));
  AOI220     u397(.A0(men_men_n413_), .A1(men_men_n95_), .B0(men_men_n412_), .B1(men_men_n158_), .Y(men_men_n414_));
  NO2        u398(.A(men_men_n414_), .B(men_men_n54_), .Y(men_men_n415_));
  NO3        u399(.A(men_men_n415_), .B(men_men_n411_), .C(men_men_n407_), .Y(men_men_n416_));
  AOI210     u400(.A0(men_men_n416_), .A1(men_men_n406_), .B0(men_men_n25_), .Y(men_men_n417_));
  NO3        u401(.A(men_men_n62_), .B(x4), .C(x1), .Y(men_men_n418_));
  NO3        u402(.A(men_men_n68_), .B(men_men_n18_), .C(x0), .Y(men_men_n419_));
  AOI220     u403(.A0(men_men_n419_), .A1(men_men_n275_), .B0(men_men_n418_), .B1(men_men_n384_), .Y(men_men_n420_));
  NO2        u404(.A(men_men_n420_), .B(men_men_n104_), .Y(men_men_n421_));
  NO3        u405(.A(men_men_n279_), .B(men_men_n180_), .C(men_men_n40_), .Y(men_men_n422_));
  OAI210     u406(.A0(men_men_n422_), .A1(men_men_n421_), .B0(x7), .Y(men_men_n423_));
  NA3        u407(.A(men_men_n62_), .B(men_men_n157_), .C(men_men_n137_), .Y(men_men_n424_));
  NA2        u408(.A(men_men_n424_), .B(men_men_n423_), .Y(men_men_n425_));
  OAI210     u409(.A0(men_men_n425_), .A1(men_men_n417_), .B0(men_men_n36_), .Y(men_men_n426_));
  NO2        u410(.A(men_men_n403_), .B(men_men_n210_), .Y(men_men_n427_));
  NO4        u411(.A(men_men_n427_), .B(men_men_n79_), .C(x4), .D(men_men_n54_), .Y(men_men_n428_));
  NA2        u412(.A(men_men_n263_), .B(men_men_n21_), .Y(men_men_n429_));
  NO2        u413(.A(men_men_n166_), .B(men_men_n138_), .Y(men_men_n430_));
  NA2        u414(.A(men_men_n430_), .B(men_men_n429_), .Y(men_men_n431_));
  AOI210     u415(.A0(men_men_n431_), .A1(men_men_n171_), .B0(men_men_n28_), .Y(men_men_n432_));
  AOI220     u416(.A0(men_men_n353_), .A1(men_men_n95_), .B0(men_men_n155_), .B1(men_men_n203_), .Y(men_men_n433_));
  NA3        u417(.A(men_men_n433_), .B(men_men_n397_), .C(men_men_n93_), .Y(men_men_n434_));
  NA2        u418(.A(men_men_n434_), .B(men_men_n181_), .Y(men_men_n435_));
  OAI220     u419(.A0(men_men_n453_), .A1(men_men_n69_), .B0(men_men_n166_), .B1(men_men_n43_), .Y(men_men_n436_));
  NA2        u420(.A(x3), .B(men_men_n54_), .Y(men_men_n437_));
  AOI210     u421(.A0(men_men_n170_), .A1(men_men_n27_), .B0(men_men_n74_), .Y(men_men_n438_));
  NO2        u422(.A(x3), .B(men_men_n54_), .Y(men_men_n439_));
  NO2        u423(.A(men_men_n439_), .B(men_men_n438_), .Y(men_men_n440_));
  OAI210     u424(.A0(men_men_n159_), .A1(men_men_n437_), .B0(men_men_n440_), .Y(men_men_n441_));
  AOI220     u425(.A0(men_men_n441_), .A1(x0), .B0(men_men_n436_), .B1(men_men_n138_), .Y(men_men_n442_));
  AOI210     u426(.A0(men_men_n442_), .A1(men_men_n435_), .B0(men_men_n241_), .Y(men_men_n443_));
  NA2        u427(.A(x9), .B(x5), .Y(men_men_n444_));
  NO4        u428(.A(men_men_n107_), .B(men_men_n444_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n445_));
  NO4        u429(.A(men_men_n445_), .B(men_men_n443_), .C(men_men_n432_), .D(men_men_n428_), .Y(men_men_n446_));
  NA3        u430(.A(men_men_n446_), .B(men_men_n426_), .C(men_men_n389_), .Y(men_men_n447_));
  AOI210     u431(.A0(men_men_n372_), .A1(men_men_n25_), .B0(men_men_n447_), .Y(men05));
  INV        u432(.A(men_men_n185_), .Y(men_men_n451_));
  INV        u433(.A(men_men_n80_), .Y(men_men_n452_));
  INV        u434(.A(x9), .Y(men_men_n453_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule