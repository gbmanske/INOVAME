//Benchmark atmr_alu4_1266_0.0156

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n973_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1048_, mai_mai_n1049_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1092_, men_men_n1093_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NA3        o034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n57_));
  NO2        o035(.A(i_1_), .B(i_6_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  OAI210     o037(.A0(ori_ori_n59_), .A1(ori_ori_n58_), .B0(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n61_));
  NAi21      o039(.An(i_2_), .B(i_7_), .Y(ori_ori_n62_));
  INV        o040(.A(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NA3        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .C(ori_ori_n31_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_1_), .B(i_10_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(i_6_), .Y(ori_ori_n67_));
  NAi31      o045(.An(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n61_), .Y(ori_ori_n68_));
  NA2        o046(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_1_), .B(i_6_), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n71_), .B(ori_ori_n25_), .Y(ori_ori_n72_));
  INV        o050(.A(i_0_), .Y(ori_ori_n73_));
  NAi21      o051(.An(i_5_), .B(i_10_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_5_), .B(i_9_), .Y(ori_ori_n75_));
  AOI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n73_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  OAI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n68_), .B0(i_0_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_12_), .B(i_5_), .Y(ori_ori_n80_));
  NA2        o058(.A(i_2_), .B(i_8_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n81_), .B(ori_ori_n58_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_9_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_3_), .B(i_7_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(ori_ori_n63_), .Y(ori_ori_n85_));
  INV        o063(.A(i_6_), .Y(ori_ori_n86_));
  OR4        o064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NO2        o066(.A(i_2_), .B(i_7_), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n88_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  OAI210     o068(.A0(ori_ori_n85_), .A1(ori_ori_n82_), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NAi21      o069(.An(i_6_), .B(i_10_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_6_), .B(i_9_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n93_), .A1(ori_ori_n92_), .B0(ori_ori_n63_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_2_), .B(i_6_), .Y(ori_ori_n95_));
  NO3        o073(.A(ori_ori_n95_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n96_), .B(ori_ori_n94_), .Y(ori_ori_n97_));
  AOI210     o075(.A0(ori_ori_n97_), .A1(ori_ori_n91_), .B0(ori_ori_n80_), .Y(ori_ori_n98_));
  AN3        o076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n99_));
  NAi21      o077(.An(i_6_), .B(i_11_), .Y(ori_ori_n100_));
  NO2        o078(.A(i_5_), .B(i_8_), .Y(ori_ori_n101_));
  NOi21      o079(.An(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  AOI220     o080(.A0(ori_ori_n102_), .A1(ori_ori_n62_), .B0(ori_ori_n99_), .B1(ori_ori_n32_), .Y(ori_ori_n103_));
  INV        o081(.A(i_7_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n46_), .B(ori_ori_n104_), .Y(ori_ori_n105_));
  NO2        o083(.A(i_0_), .B(i_5_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(ori_ori_n86_), .Y(ori_ori_n107_));
  NA2        o085(.A(i_12_), .B(i_3_), .Y(ori_ori_n108_));
  INV        o086(.A(ori_ori_n108_), .Y(ori_ori_n109_));
  NA3        o087(.A(ori_ori_n109_), .B(ori_ori_n107_), .C(ori_ori_n105_), .Y(ori_ori_n110_));
  NAi21      o088(.An(i_7_), .B(i_11_), .Y(ori_ori_n111_));
  AN2        o089(.A(i_2_), .B(i_10_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n112_), .B(i_7_), .Y(ori_ori_n113_));
  OR2        o091(.A(ori_ori_n80_), .B(ori_ori_n58_), .Y(ori_ori_n114_));
  NO2        o092(.A(i_8_), .B(ori_ori_n104_), .Y(ori_ori_n115_));
  NO3        o093(.A(ori_ori_n115_), .B(ori_ori_n114_), .C(ori_ori_n113_), .Y(ori_ori_n116_));
  NA2        o094(.A(i_12_), .B(i_7_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n63_), .B(ori_ori_n26_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(i_0_), .Y(ori_ori_n119_));
  NA2        o097(.A(i_11_), .B(i_12_), .Y(ori_ori_n120_));
  OAI210     o098(.A0(ori_ori_n119_), .A1(ori_ori_n117_), .B0(ori_ori_n120_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n121_), .B(ori_ori_n116_), .Y(ori_ori_n122_));
  NA3        o100(.A(ori_ori_n122_), .B(ori_ori_n110_), .C(ori_ori_n103_), .Y(ori_ori_n123_));
  NOi21      o101(.An(i_1_), .B(i_5_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(i_11_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n126_));
  NA2        o104(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(ori_ori_n126_), .Y(ori_ori_n128_));
  NO2        o106(.A(ori_ori_n128_), .B(ori_ori_n46_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n93_), .B(ori_ori_n92_), .Y(ori_ori_n130_));
  NAi21      o108(.An(i_3_), .B(i_8_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n131_), .B(ori_ori_n62_), .Y(ori_ori_n132_));
  NOi31      o110(.An(ori_ori_n132_), .B(ori_ori_n130_), .C(ori_ori_n129_), .Y(ori_ori_n133_));
  NO2        o111(.A(i_1_), .B(ori_ori_n86_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_6_), .B(i_5_), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n135_), .B(i_3_), .Y(ori_ori_n136_));
  AO210      o114(.A0(ori_ori_n136_), .A1(ori_ori_n47_), .B0(ori_ori_n134_), .Y(ori_ori_n137_));
  OAI220     o115(.A0(ori_ori_n137_), .A1(ori_ori_n111_), .B0(ori_ori_n133_), .B1(ori_ori_n125_), .Y(ori_ori_n138_));
  NO3        o116(.A(ori_ori_n138_), .B(ori_ori_n123_), .C(ori_ori_n98_), .Y(ori_ori_n139_));
  NA3        o117(.A(ori_ori_n139_), .B(ori_ori_n79_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o118(.A(ori_ori_n63_), .B(ori_ori_n37_), .Y(ori_ori_n141_));
  INV        o119(.A(i_6_), .Y(ori_ori_n142_));
  NA2        o120(.A(ori_ori_n142_), .B(ori_ori_n141_), .Y(ori_ori_n143_));
  NA4        o121(.A(ori_ori_n143_), .B(ori_ori_n77_), .C(ori_ori_n69_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o122(.A(i_8_), .B(i_7_), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n145_), .B(i_6_), .Y(ori_ori_n146_));
  NO2        o124(.A(i_12_), .B(i_13_), .Y(ori_ori_n147_));
  NAi21      o125(.An(i_5_), .B(i_11_), .Y(ori_ori_n148_));
  NOi21      o126(.An(ori_ori_n147_), .B(ori_ori_n148_), .Y(ori_ori_n149_));
  NO2        o127(.A(i_0_), .B(i_1_), .Y(ori_ori_n150_));
  NA2        o128(.A(i_2_), .B(i_3_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n151_), .B(i_4_), .Y(ori_ori_n152_));
  NA3        o130(.A(ori_ori_n152_), .B(ori_ori_n150_), .C(ori_ori_n149_), .Y(ori_ori_n153_));
  AN2        o131(.A(ori_ori_n147_), .B(ori_ori_n83_), .Y(ori_ori_n154_));
  NA2        o132(.A(i_1_), .B(i_5_), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n73_), .B(ori_ori_n46_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n156_), .B(ori_ori_n36_), .Y(ori_ori_n157_));
  OR2        o135(.A(i_0_), .B(i_1_), .Y(ori_ori_n158_));
  NO3        o136(.A(ori_ori_n158_), .B(ori_ori_n80_), .C(i_13_), .Y(ori_ori_n159_));
  NAi32      o137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n160_));
  NAi21      o138(.An(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NOi21      o139(.An(i_4_), .B(i_10_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n162_), .B(ori_ori_n40_), .Y(ori_ori_n163_));
  NO2        o141(.A(i_3_), .B(i_5_), .Y(ori_ori_n164_));
  NO3        o142(.A(ori_ori_n73_), .B(i_2_), .C(i_1_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n165_), .B(ori_ori_n164_), .Y(ori_ori_n166_));
  OAI210     o144(.A0(ori_ori_n166_), .A1(ori_ori_n163_), .B0(ori_ori_n161_), .Y(ori_ori_n167_));
  INV        o145(.A(ori_ori_n167_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n168_), .B(ori_ori_n146_), .Y(ori_ori_n169_));
  NA2        o147(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n170_));
  NOi21      o148(.An(i_4_), .B(i_9_), .Y(ori_ori_n171_));
  NOi21      o149(.An(i_11_), .B(i_13_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(ori_ori_n171_), .Y(ori_ori_n173_));
  NO2        o151(.A(i_4_), .B(i_5_), .Y(ori_ori_n174_));
  NAi21      o152(.An(i_12_), .B(i_11_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n73_), .B(ori_ori_n63_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(ori_ori_n46_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n36_), .B(i_5_), .Y(ori_ori_n178_));
  NAi31      o156(.An(ori_ori_n178_), .B(ori_ori_n154_), .C(i_11_), .Y(ori_ori_n179_));
  NA2        o157(.A(i_3_), .B(i_5_), .Y(ori_ori_n180_));
  OR2        o158(.A(ori_ori_n180_), .B(ori_ori_n173_), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n181_), .A1(ori_ori_n179_), .B0(ori_ori_n177_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n183_));
  NO2        o161(.A(i_13_), .B(i_10_), .Y(ori_ori_n184_));
  NA3        o162(.A(ori_ori_n184_), .B(ori_ori_n183_), .C(ori_ori_n44_), .Y(ori_ori_n185_));
  NO2        o163(.A(i_2_), .B(i_1_), .Y(ori_ori_n186_));
  NAi21      o164(.An(i_4_), .B(i_12_), .Y(ori_ori_n187_));
  INV        o165(.A(ori_ori_n182_), .Y(ori_ori_n188_));
  INV        o166(.A(i_8_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n189_), .B(i_7_), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n190_), .B(i_6_), .Y(ori_ori_n191_));
  NO3        o169(.A(i_3_), .B(ori_ori_n86_), .C(ori_ori_n48_), .Y(ori_ori_n192_));
  NO3        o170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n193_));
  NO3        o171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n194_));
  NO2        o172(.A(i_3_), .B(i_8_), .Y(ori_ori_n195_));
  NO3        o173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n196_));
  NA3        o174(.A(ori_ori_n196_), .B(ori_ori_n195_), .C(ori_ori_n40_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n106_), .B(ori_ori_n58_), .Y(ori_ori_n198_));
  INV        o176(.A(ori_ori_n198_), .Y(ori_ori_n199_));
  NO2        o177(.A(i_13_), .B(i_9_), .Y(ori_ori_n200_));
  NAi21      o178(.An(i_12_), .B(i_3_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n202_));
  NO3        o180(.A(i_0_), .B(i_2_), .C(ori_ori_n63_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n199_), .B(ori_ori_n197_), .Y(ori_ori_n204_));
  NA2        o182(.A(ori_ori_n204_), .B(i_7_), .Y(ori_ori_n205_));
  OAI220     o183(.A0(ori_ori_n205_), .A1(i_4_), .B0(ori_ori_n191_), .B1(ori_ori_n188_), .Y(ori_ori_n206_));
  NAi21      o184(.An(i_12_), .B(i_7_), .Y(ori_ori_n207_));
  NA3        o185(.A(i_13_), .B(ori_ori_n189_), .C(i_10_), .Y(ori_ori_n208_));
  NA2        o186(.A(i_0_), .B(i_5_), .Y(ori_ori_n209_));
  NAi31      o187(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n73_), .B(ori_ori_n26_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n46_), .B(ori_ori_n63_), .Y(ori_ori_n213_));
  NA3        o191(.A(ori_ori_n213_), .B(ori_ori_n212_), .C(ori_ori_n211_), .Y(ori_ori_n214_));
  INV        o192(.A(i_13_), .Y(ori_ori_n215_));
  NO2        o193(.A(i_12_), .B(ori_ori_n215_), .Y(ori_ori_n216_));
  NA3        o194(.A(ori_ori_n216_), .B(ori_ori_n193_), .C(ori_ori_n192_), .Y(ori_ori_n217_));
  OAI210     o195(.A0(ori_ori_n214_), .A1(ori_ori_n210_), .B0(ori_ori_n217_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n145_), .Y(ori_ori_n219_));
  NO2        o197(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n220_));
  OR2        o198(.A(i_8_), .B(i_7_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n53_), .B(i_1_), .Y(ori_ori_n222_));
  INV        o200(.A(i_12_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n44_), .B(ori_ori_n223_), .Y(ori_ori_n224_));
  NO3        o202(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n225_));
  NA2        o203(.A(i_2_), .B(i_1_), .Y(ori_ori_n226_));
  NO3        o204(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n227_));
  NAi21      o205(.An(i_4_), .B(i_3_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n228_), .B(ori_ori_n75_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_0_), .B(i_6_), .Y(ori_ori_n230_));
  NOi41      o208(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n226_), .B(ori_ori_n180_), .Y(ori_ori_n232_));
  NO2        o210(.A(i_11_), .B(ori_ori_n215_), .Y(ori_ori_n233_));
  NOi21      o211(.An(i_1_), .B(i_6_), .Y(ori_ori_n234_));
  NAi21      o212(.An(i_3_), .B(i_7_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n223_), .B(i_9_), .Y(ori_ori_n236_));
  OR4        o214(.A(ori_ori_n236_), .B(ori_ori_n235_), .C(ori_ori_n234_), .D(ori_ori_n183_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n238_));
  NA2        o216(.A(i_3_), .B(i_9_), .Y(ori_ori_n239_));
  NAi21      o217(.An(i_7_), .B(i_10_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n240_), .B(ori_ori_n239_), .Y(ori_ori_n241_));
  NA3        o219(.A(ori_ori_n241_), .B(ori_ori_n238_), .C(ori_ori_n64_), .Y(ori_ori_n242_));
  NA2        o220(.A(ori_ori_n242_), .B(ori_ori_n237_), .Y(ori_ori_n243_));
  INV        o221(.A(ori_ori_n146_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n223_), .B(i_13_), .Y(ori_ori_n245_));
  NO2        o223(.A(ori_ori_n245_), .B(ori_ori_n75_), .Y(ori_ori_n246_));
  AOI220     o224(.A0(ori_ori_n246_), .A1(ori_ori_n244_), .B0(ori_ori_n243_), .B1(ori_ori_n233_), .Y(ori_ori_n247_));
  NO2        o225(.A(ori_ori_n221_), .B(ori_ori_n37_), .Y(ori_ori_n248_));
  NA2        o226(.A(i_12_), .B(i_6_), .Y(ori_ori_n249_));
  OR2        o227(.A(i_13_), .B(i_9_), .Y(ori_ori_n250_));
  NO3        o228(.A(ori_ori_n250_), .B(ori_ori_n249_), .C(ori_ori_n48_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n228_), .B(i_2_), .Y(ori_ori_n252_));
  NA3        o230(.A(ori_ori_n252_), .B(ori_ori_n251_), .C(ori_ori_n44_), .Y(ori_ori_n253_));
  NA2        o231(.A(ori_ori_n233_), .B(i_9_), .Y(ori_ori_n254_));
  NA2        o232(.A(ori_ori_n238_), .B(ori_ori_n64_), .Y(ori_ori_n255_));
  OAI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n254_), .B0(ori_ori_n253_), .Y(ori_ori_n256_));
  NA2        o234(.A(ori_ori_n156_), .B(ori_ori_n63_), .Y(ori_ori_n257_));
  NO3        o235(.A(i_11_), .B(ori_ori_n215_), .C(ori_ori_n25_), .Y(ori_ori_n258_));
  NO2        o236(.A(ori_ori_n235_), .B(i_8_), .Y(ori_ori_n259_));
  NO2        o237(.A(i_6_), .B(ori_ori_n48_), .Y(ori_ori_n260_));
  NA3        o238(.A(ori_ori_n260_), .B(ori_ori_n259_), .C(ori_ori_n258_), .Y(ori_ori_n261_));
  NO3        o239(.A(ori_ori_n26_), .B(ori_ori_n86_), .C(i_5_), .Y(ori_ori_n262_));
  NA3        o240(.A(ori_ori_n262_), .B(ori_ori_n248_), .C(ori_ori_n216_), .Y(ori_ori_n263_));
  AOI210     o241(.A0(ori_ori_n263_), .A1(ori_ori_n261_), .B0(ori_ori_n257_), .Y(ori_ori_n264_));
  AOI210     o242(.A0(ori_ori_n256_), .A1(ori_ori_n248_), .B0(ori_ori_n264_), .Y(ori_ori_n265_));
  NA3        o243(.A(ori_ori_n265_), .B(ori_ori_n247_), .C(ori_ori_n219_), .Y(ori_ori_n266_));
  NO3        o244(.A(i_12_), .B(ori_ori_n215_), .C(ori_ori_n37_), .Y(ori_ori_n267_));
  INV        o245(.A(ori_ori_n267_), .Y(ori_ori_n268_));
  NA2        o246(.A(i_8_), .B(ori_ori_n104_), .Y(ori_ori_n269_));
  NOi21      o247(.An(ori_ori_n164_), .B(ori_ori_n86_), .Y(ori_ori_n270_));
  NO3        o248(.A(i_0_), .B(ori_ori_n46_), .C(i_1_), .Y(ori_ori_n271_));
  AOI220     o249(.A0(ori_ori_n271_), .A1(ori_ori_n192_), .B0(ori_ori_n270_), .B1(ori_ori_n222_), .Y(ori_ori_n272_));
  NO2        o250(.A(ori_ori_n272_), .B(ori_ori_n269_), .Y(ori_ori_n273_));
  NO3        o251(.A(i_0_), .B(i_2_), .C(ori_ori_n63_), .Y(ori_ori_n274_));
  NO2        o252(.A(ori_ori_n226_), .B(i_0_), .Y(ori_ori_n275_));
  AOI220     o253(.A0(ori_ori_n275_), .A1(ori_ori_n190_), .B0(ori_ori_n274_), .B1(ori_ori_n145_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n260_), .B(ori_ori_n26_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n277_), .B(ori_ori_n276_), .Y(ori_ori_n278_));
  NA2        o256(.A(i_0_), .B(i_1_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n279_), .B(i_2_), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n59_), .B(i_6_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n166_), .B(ori_ori_n146_), .Y(ori_ori_n282_));
  NO3        o260(.A(ori_ori_n282_), .B(ori_ori_n278_), .C(ori_ori_n273_), .Y(ori_ori_n283_));
  NO2        o261(.A(i_2_), .B(ori_ori_n104_), .Y(ori_ori_n284_));
  NA2        o262(.A(i_1_), .B(ori_ori_n36_), .Y(ori_ori_n285_));
  AN2        o263(.A(i_3_), .B(i_10_), .Y(ori_ori_n286_));
  NO2        o264(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n287_));
  NO2        o265(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n283_), .B(ori_ori_n268_), .Y(ori_ori_n289_));
  NO4        o267(.A(ori_ori_n289_), .B(ori_ori_n266_), .C(ori_ori_n206_), .D(ori_ori_n169_), .Y(ori_ori_n290_));
  NO3        o268(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n291_));
  NO2        o269(.A(ori_ori_n59_), .B(ori_ori_n86_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n275_), .B(ori_ori_n292_), .Y(ori_ori_n293_));
  NO3        o271(.A(i_6_), .B(ori_ori_n189_), .C(i_7_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n294_), .B(ori_ori_n193_), .Y(ori_ori_n295_));
  AOI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n293_), .B0(ori_ori_n170_), .Y(ori_ori_n296_));
  NO2        o274(.A(i_2_), .B(i_3_), .Y(ori_ori_n297_));
  OR2        o275(.A(i_0_), .B(i_5_), .Y(ori_ori_n298_));
  NA3        o276(.A(ori_ori_n275_), .B(ori_ori_n270_), .C(ori_ori_n115_), .Y(ori_ori_n299_));
  NAi21      o277(.An(i_8_), .B(i_7_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n158_), .B(ori_ori_n46_), .Y(ori_ori_n301_));
  INV        o279(.A(ori_ori_n299_), .Y(ori_ori_n302_));
  OAI210     o280(.A0(ori_ori_n302_), .A1(ori_ori_n296_), .B0(i_4_), .Y(ori_ori_n303_));
  NO2        o281(.A(i_12_), .B(i_10_), .Y(ori_ori_n304_));
  NOi21      o282(.An(i_5_), .B(i_0_), .Y(ori_ori_n305_));
  AOI210     o283(.A0(i_2_), .A1(ori_ori_n48_), .B0(ori_ori_n104_), .Y(ori_ori_n306_));
  NO4        o284(.A(ori_ori_n306_), .B(ori_ori_n285_), .C(ori_ori_n305_), .D(ori_ori_n131_), .Y(ori_ori_n307_));
  NA4        o285(.A(ori_ori_n84_), .B(ori_ori_n36_), .C(ori_ori_n86_), .D(i_8_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n307_), .B(ori_ori_n304_), .Y(ori_ori_n309_));
  NO2        o287(.A(i_6_), .B(i_8_), .Y(ori_ori_n310_));
  NOi21      o288(.An(i_0_), .B(i_2_), .Y(ori_ori_n311_));
  AN2        o289(.A(ori_ori_n311_), .B(ori_ori_n310_), .Y(ori_ori_n312_));
  NO2        o290(.A(i_1_), .B(i_7_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n309_), .B(ori_ori_n303_), .Y(ori_ori_n314_));
  NOi21      o292(.An(ori_ori_n155_), .B(ori_ori_n107_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n315_), .B(ori_ori_n127_), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n316_), .B(i_3_), .Y(ori_ori_n317_));
  NO2        o295(.A(ori_ori_n189_), .B(i_9_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n318_), .B(ori_ori_n198_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n319_), .B(ori_ori_n46_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n320_), .B(ori_ori_n278_), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n321_), .A1(ori_ori_n317_), .B0(ori_ori_n163_), .Y(ori_ori_n322_));
  AOI210     o300(.A0(ori_ori_n314_), .A1(ori_ori_n291_), .B0(ori_ori_n322_), .Y(ori_ori_n323_));
  NOi32      o301(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n324_));
  INV        o302(.A(ori_ori_n324_), .Y(ori_ori_n325_));
  NAi21      o303(.An(i_1_), .B(i_5_), .Y(ori_ori_n326_));
  NAi41      o304(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n327_));
  OAI220     o305(.A0(ori_ori_n327_), .A1(ori_ori_n326_), .B0(ori_ori_n210_), .B1(ori_ori_n160_), .Y(ori_ori_n328_));
  AOI210     o306(.A0(ori_ori_n327_), .A1(ori_ori_n160_), .B0(ori_ori_n158_), .Y(ori_ori_n329_));
  NOi32      o307(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n330_));
  NAi21      o308(.An(i_6_), .B(i_1_), .Y(ori_ori_n331_));
  NA3        o309(.A(ori_ori_n331_), .B(ori_ori_n330_), .C(ori_ori_n46_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n332_), .B(i_0_), .Y(ori_ori_n333_));
  OR3        o311(.A(ori_ori_n333_), .B(ori_ori_n329_), .C(ori_ori_n328_), .Y(ori_ori_n334_));
  NO2        o312(.A(i_1_), .B(ori_ori_n104_), .Y(ori_ori_n335_));
  NAi21      o313(.An(i_3_), .B(i_4_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n336_), .B(i_9_), .Y(ori_ori_n337_));
  AN2        o315(.A(i_6_), .B(i_7_), .Y(ori_ori_n338_));
  OAI210     o316(.A0(ori_ori_n338_), .A1(ori_ori_n335_), .B0(ori_ori_n337_), .Y(ori_ori_n339_));
  NA2        o317(.A(i_2_), .B(i_7_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n336_), .B(i_10_), .Y(ori_ori_n341_));
  NA3        o319(.A(ori_ori_n341_), .B(ori_ori_n340_), .C(ori_ori_n230_), .Y(ori_ori_n342_));
  AOI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n339_), .B0(ori_ori_n183_), .Y(ori_ori_n343_));
  AOI210     o321(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n344_));
  OAI210     o322(.A0(ori_ori_n344_), .A1(ori_ori_n186_), .B0(ori_ori_n341_), .Y(ori_ori_n345_));
  AOI220     o323(.A0(ori_ori_n341_), .A1(ori_ori_n313_), .B0(ori_ori_n225_), .B1(ori_ori_n186_), .Y(ori_ori_n346_));
  AOI210     o324(.A0(ori_ori_n346_), .A1(ori_ori_n345_), .B0(i_5_), .Y(ori_ori_n347_));
  NO3        o325(.A(ori_ori_n347_), .B(ori_ori_n343_), .C(ori_ori_n334_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(ori_ori_n325_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n59_), .B(ori_ori_n25_), .Y(ori_ori_n350_));
  AN2        o328(.A(i_12_), .B(i_5_), .Y(ori_ori_n351_));
  NO2        o329(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n352_), .B(ori_ori_n351_), .Y(ori_ori_n353_));
  NO2        o331(.A(i_11_), .B(i_6_), .Y(ori_ori_n354_));
  NA3        o332(.A(ori_ori_n354_), .B(ori_ori_n301_), .C(ori_ori_n215_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n355_), .B(ori_ori_n353_), .Y(ori_ori_n356_));
  NO2        o334(.A(ori_ori_n228_), .B(i_5_), .Y(ori_ori_n357_));
  NO2        o335(.A(i_5_), .B(i_10_), .Y(ori_ori_n358_));
  AOI220     o336(.A0(ori_ori_n358_), .A1(ori_ori_n252_), .B0(ori_ori_n357_), .B1(ori_ori_n193_), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n147_), .B(ori_ori_n45_), .Y(ori_ori_n360_));
  NO2        o338(.A(ori_ori_n360_), .B(ori_ori_n359_), .Y(ori_ori_n361_));
  OAI210     o339(.A0(ori_ori_n361_), .A1(ori_ori_n356_), .B0(ori_ori_n350_), .Y(ori_ori_n362_));
  NO2        o340(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n363_));
  NO2        o341(.A(ori_ori_n153_), .B(ori_ori_n86_), .Y(ori_ori_n364_));
  OAI210     o342(.A0(ori_ori_n364_), .A1(ori_ori_n356_), .B0(ori_ori_n363_), .Y(ori_ori_n365_));
  NO3        o343(.A(ori_ori_n86_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n366_));
  NO2        o344(.A(i_11_), .B(i_12_), .Y(ori_ori_n367_));
  NA2        o345(.A(ori_ori_n358_), .B(ori_ori_n223_), .Y(ori_ori_n368_));
  NAi21      o346(.An(i_13_), .B(i_0_), .Y(ori_ori_n369_));
  NA2        o347(.A(ori_ori_n365_), .B(ori_ori_n362_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n44_), .B(ori_ori_n215_), .Y(ori_ori_n371_));
  NO3        o349(.A(i_1_), .B(i_12_), .C(ori_ori_n86_), .Y(ori_ori_n372_));
  NO2        o350(.A(i_0_), .B(i_11_), .Y(ori_ori_n373_));
  AN2        o351(.A(i_1_), .B(i_6_), .Y(ori_ori_n374_));
  NOi21      o352(.An(i_2_), .B(i_12_), .Y(ori_ori_n375_));
  NA2        o353(.A(ori_ori_n145_), .B(i_9_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n376_), .B(i_4_), .Y(ori_ori_n377_));
  NAi21      o355(.An(i_9_), .B(i_4_), .Y(ori_ori_n378_));
  OR2        o356(.A(i_13_), .B(i_10_), .Y(ori_ori_n379_));
  NO3        o357(.A(ori_ori_n379_), .B(ori_ori_n120_), .C(ori_ori_n378_), .Y(ori_ori_n380_));
  NO2        o358(.A(ori_ori_n173_), .B(ori_ori_n126_), .Y(ori_ori_n381_));
  NO2        o359(.A(ori_ori_n104_), .B(ori_ori_n25_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n267_), .B(ori_ori_n382_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n383_), .B(ori_ori_n315_), .Y(ori_ori_n384_));
  INV        o362(.A(ori_ori_n384_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n385_), .B(ori_ori_n26_), .Y(ori_ori_n386_));
  INV        o364(.A(ori_ori_n299_), .Y(ori_ori_n387_));
  NO2        o365(.A(ori_ori_n180_), .B(ori_ori_n86_), .Y(ori_ori_n388_));
  AOI220     o366(.A0(ori_ori_n388_), .A1(ori_ori_n280_), .B0(ori_ori_n262_), .B1(ori_ori_n203_), .Y(ori_ori_n389_));
  NO2        o367(.A(ori_ori_n389_), .B(ori_ori_n269_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n390_), .B(ori_ori_n387_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n192_), .B(ori_ori_n99_), .Y(ori_ori_n392_));
  NA3        o370(.A(ori_ori_n301_), .B(ori_ori_n164_), .C(ori_ori_n86_), .Y(ori_ori_n393_));
  AOI210     o371(.A0(ori_ori_n393_), .A1(ori_ori_n392_), .B0(ori_ori_n300_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n189_), .B(i_10_), .Y(ori_ori_n395_));
  NA3        o373(.A(ori_ori_n238_), .B(ori_ori_n64_), .C(i_2_), .Y(ori_ori_n396_));
  NA2        o374(.A(ori_ori_n281_), .B(ori_ori_n222_), .Y(ori_ori_n397_));
  OAI220     o375(.A0(ori_ori_n397_), .A1(ori_ori_n180_), .B0(ori_ori_n396_), .B1(ori_ori_n395_), .Y(ori_ori_n398_));
  NO2        o376(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n399_));
  NA3        o377(.A(ori_ori_n313_), .B(ori_ori_n312_), .C(ori_ori_n399_), .Y(ori_ori_n400_));
  INV        o378(.A(ori_ori_n400_), .Y(ori_ori_n401_));
  NO3        o379(.A(ori_ori_n401_), .B(ori_ori_n398_), .C(ori_ori_n394_), .Y(ori_ori_n402_));
  AOI210     o380(.A0(ori_ori_n402_), .A1(ori_ori_n391_), .B0(ori_ori_n254_), .Y(ori_ori_n403_));
  NO4        o381(.A(ori_ori_n403_), .B(ori_ori_n386_), .C(ori_ori_n370_), .D(ori_ori_n349_), .Y(ori_ori_n404_));
  NO2        o382(.A(ori_ori_n63_), .B(i_4_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n73_), .B(i_13_), .Y(ori_ori_n406_));
  NA3        o384(.A(ori_ori_n406_), .B(ori_ori_n405_), .C(i_2_), .Y(ori_ori_n407_));
  NO2        o385(.A(i_10_), .B(i_9_), .Y(ori_ori_n408_));
  NAi21      o386(.An(i_12_), .B(i_8_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n409_), .B(i_3_), .Y(ori_ori_n410_));
  NA2        o388(.A(ori_ori_n410_), .B(ori_ori_n408_), .Y(ori_ori_n411_));
  NO2        o389(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n412_), .B(ori_ori_n107_), .Y(ori_ori_n413_));
  OAI220     o391(.A0(ori_ori_n413_), .A1(ori_ori_n197_), .B0(ori_ori_n411_), .B1(ori_ori_n407_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n288_), .B(i_0_), .Y(ori_ori_n415_));
  NO3        o393(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n249_), .B(ori_ori_n100_), .Y(ori_ori_n417_));
  NA2        o395(.A(ori_ori_n417_), .B(ori_ori_n416_), .Y(ori_ori_n418_));
  NA2        o396(.A(i_8_), .B(i_9_), .Y(ori_ori_n419_));
  AOI210     o397(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n420_));
  OR2        o398(.A(ori_ori_n420_), .B(ori_ori_n419_), .Y(ori_ori_n421_));
  NA2        o399(.A(ori_ori_n267_), .B(ori_ori_n198_), .Y(ori_ori_n422_));
  OAI220     o400(.A0(ori_ori_n422_), .A1(ori_ori_n421_), .B0(ori_ori_n418_), .B1(ori_ori_n415_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n233_), .B(ori_ori_n287_), .Y(ori_ori_n424_));
  NO3        o402(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n425_));
  INV        o403(.A(ori_ori_n425_), .Y(ori_ori_n426_));
  NA3        o404(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n427_));
  NA4        o405(.A(ori_ori_n148_), .B(ori_ori_n118_), .C(ori_ori_n80_), .D(ori_ori_n23_), .Y(ori_ori_n428_));
  OAI220     o406(.A0(ori_ori_n428_), .A1(ori_ori_n427_), .B0(ori_ori_n426_), .B1(ori_ori_n424_), .Y(ori_ori_n429_));
  NO3        o407(.A(ori_ori_n429_), .B(ori_ori_n423_), .C(ori_ori_n414_), .Y(ori_ori_n430_));
  NA2        o408(.A(ori_ori_n99_), .B(i_13_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n388_), .B(ori_ori_n350_), .Y(ori_ori_n432_));
  NO2        o410(.A(i_2_), .B(i_13_), .Y(ori_ori_n433_));
  NO2        o411(.A(ori_ori_n432_), .B(ori_ori_n431_), .Y(ori_ori_n434_));
  NO3        o412(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n435_));
  NO2        o413(.A(i_6_), .B(i_7_), .Y(ori_ori_n436_));
  NO2        o414(.A(i_11_), .B(i_1_), .Y(ori_ori_n437_));
  OR2        o415(.A(i_11_), .B(i_8_), .Y(ori_ori_n438_));
  NOi21      o416(.An(i_2_), .B(i_7_), .Y(ori_ori_n439_));
  NO2        o417(.A(i_6_), .B(i_10_), .Y(ori_ori_n440_));
  NA3        o418(.A(ori_ori_n231_), .B(ori_ori_n172_), .C(ori_ori_n135_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n442_));
  NO2        o420(.A(ori_ori_n158_), .B(i_3_), .Y(ori_ori_n443_));
  NAi31      o421(.An(ori_ori_n442_), .B(ori_ori_n443_), .C(ori_ori_n216_), .Y(ori_ori_n444_));
  NA3        o422(.A(ori_ori_n363_), .B(ori_ori_n176_), .C(ori_ori_n152_), .Y(ori_ori_n445_));
  NA3        o423(.A(ori_ori_n445_), .B(ori_ori_n444_), .C(ori_ori_n441_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n446_), .B(ori_ori_n434_), .Y(ori_ori_n447_));
  NA2        o425(.A(ori_ori_n416_), .B(ori_ori_n351_), .Y(ori_ori_n448_));
  NA2        o426(.A(ori_ori_n425_), .B(ori_ori_n358_), .Y(ori_ori_n449_));
  NO2        o427(.A(ori_ori_n449_), .B(ori_ori_n214_), .Y(ori_ori_n450_));
  NAi21      o428(.An(ori_ori_n208_), .B(ori_ori_n367_), .Y(ori_ori_n451_));
  NA2        o429(.A(ori_ori_n313_), .B(ori_ori_n209_), .Y(ori_ori_n452_));
  NO2        o430(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n453_));
  NO2        o431(.A(i_0_), .B(ori_ori_n86_), .Y(ori_ori_n454_));
  NA3        o432(.A(ori_ori_n454_), .B(ori_ori_n453_), .C(ori_ori_n145_), .Y(ori_ori_n455_));
  OR3        o433(.A(ori_ori_n285_), .B(ori_ori_n38_), .C(ori_ori_n46_), .Y(ori_ori_n456_));
  OAI220     o434(.A0(ori_ori_n456_), .A1(ori_ori_n455_), .B0(ori_ori_n452_), .B1(ori_ori_n451_), .Y(ori_ori_n457_));
  NA2        o435(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n458_));
  NA2        o436(.A(ori_ori_n291_), .B(ori_ori_n225_), .Y(ori_ori_n459_));
  OAI220     o437(.A0(ori_ori_n459_), .A1(ori_ori_n396_), .B0(ori_ori_n458_), .B1(ori_ori_n431_), .Y(ori_ori_n460_));
  NO3        o438(.A(ori_ori_n460_), .B(ori_ori_n457_), .C(ori_ori_n450_), .Y(ori_ori_n461_));
  NA3        o439(.A(ori_ori_n461_), .B(ori_ori_n447_), .C(ori_ori_n430_), .Y(ori_ori_n462_));
  NA2        o440(.A(ori_ori_n125_), .B(ori_ori_n114_), .Y(ori_ori_n463_));
  AN2        o441(.A(ori_ori_n463_), .B(ori_ori_n416_), .Y(ori_ori_n464_));
  NA2        o442(.A(ori_ori_n464_), .B(ori_ori_n288_), .Y(ori_ori_n465_));
  NA4        o443(.A(ori_ori_n406_), .B(ori_ori_n405_), .C(ori_ori_n195_), .D(i_2_), .Y(ori_ori_n466_));
  INV        o444(.A(ori_ori_n466_), .Y(ori_ori_n467_));
  NA2        o445(.A(ori_ori_n351_), .B(ori_ori_n215_), .Y(ori_ori_n468_));
  NA2        o446(.A(ori_ori_n324_), .B(ori_ori_n73_), .Y(ori_ori_n469_));
  NA2        o447(.A(ori_ori_n338_), .B(ori_ori_n330_), .Y(ori_ori_n470_));
  OR2        o448(.A(ori_ori_n468_), .B(ori_ori_n470_), .Y(ori_ori_n471_));
  NO2        o449(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n472_));
  AOI210     o450(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n380_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n473_), .B(ori_ori_n471_), .Y(ori_ori_n474_));
  AOI210     o452(.A0(ori_ori_n467_), .A1(ori_ori_n196_), .B0(ori_ori_n474_), .Y(ori_ori_n475_));
  NA2        o453(.A(ori_ori_n238_), .B(ori_ori_n64_), .Y(ori_ori_n476_));
  OAI210     o454(.A0(i_8_), .A1(ori_ori_n476_), .B0(ori_ori_n137_), .Y(ori_ori_n477_));
  NA2        o455(.A(ori_ori_n477_), .B(ori_ori_n381_), .Y(ori_ori_n478_));
  NA3        o456(.A(ori_ori_n478_), .B(ori_ori_n475_), .C(ori_ori_n465_), .Y(ori_ori_n479_));
  NO2        o457(.A(i_12_), .B(ori_ori_n189_), .Y(ori_ori_n480_));
  NO2        o458(.A(i_8_), .B(i_7_), .Y(ori_ori_n481_));
  OAI210     o459(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(ori_ori_n482_));
  NA2        o460(.A(ori_ori_n482_), .B(ori_ori_n213_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n483_), .B(ori_ori_n228_), .Y(ori_ori_n484_));
  NA2        o462(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n485_));
  NO2        o463(.A(ori_ori_n485_), .B(i_6_), .Y(ori_ori_n486_));
  NA3        o464(.A(ori_ori_n486_), .B(ori_ori_n484_), .C(ori_ori_n481_), .Y(ori_ori_n487_));
  AOI220     o465(.A0(ori_ori_n388_), .A1(ori_ori_n301_), .B0(ori_ori_n232_), .B1(ori_ori_n230_), .Y(ori_ori_n488_));
  OAI220     o466(.A0(ori_ori_n488_), .A1(ori_ori_n245_), .B0(ori_ori_n431_), .B1(ori_ori_n136_), .Y(ori_ori_n489_));
  NA2        o467(.A(ori_ori_n489_), .B(ori_ori_n248_), .Y(ori_ori_n490_));
  NA3        o468(.A(ori_ori_n286_), .B(ori_ori_n174_), .C(ori_ori_n99_), .Y(ori_ori_n491_));
  NO2        o469(.A(ori_ori_n211_), .B(ori_ori_n44_), .Y(ori_ori_n492_));
  NO2        o470(.A(ori_ori_n158_), .B(i_5_), .Y(ori_ori_n493_));
  NA3        o471(.A(ori_ori_n493_), .B(ori_ori_n371_), .C(ori_ori_n297_), .Y(ori_ori_n494_));
  OAI210     o472(.A0(ori_ori_n494_), .A1(ori_ori_n492_), .B0(ori_ori_n491_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n495_), .B(ori_ori_n425_), .Y(ori_ori_n496_));
  NA3        o474(.A(ori_ori_n496_), .B(ori_ori_n490_), .C(ori_ori_n487_), .Y(ori_ori_n497_));
  NA3        o475(.A(ori_ori_n209_), .B(ori_ori_n71_), .C(ori_ori_n44_), .Y(ori_ori_n498_));
  NA2        o476(.A(ori_ori_n267_), .B(ori_ori_n84_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n498_), .B(ori_ori_n499_), .Y(ori_ori_n500_));
  NA2        o478(.A(ori_ori_n213_), .B(ori_ori_n212_), .Y(ori_ori_n501_));
  NA2        o479(.A(ori_ori_n408_), .B(ori_ori_n211_), .Y(ori_ori_n502_));
  NO2        o480(.A(ori_ori_n501_), .B(ori_ori_n502_), .Y(ori_ori_n503_));
  AOI210     o481(.A0(ori_ori_n331_), .A1(ori_ori_n46_), .B0(ori_ori_n335_), .Y(ori_ori_n504_));
  NA2        o482(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n505_));
  NA3        o483(.A(ori_ori_n480_), .B(ori_ori_n258_), .C(ori_ori_n505_), .Y(ori_ori_n506_));
  NO2        o484(.A(ori_ori_n504_), .B(ori_ori_n506_), .Y(ori_ori_n507_));
  NO3        o485(.A(ori_ori_n507_), .B(ori_ori_n503_), .C(ori_ori_n500_), .Y(ori_ori_n508_));
  NO4        o486(.A(ori_ori_n234_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n509_));
  NO3        o487(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n510_));
  NO2        o488(.A(ori_ori_n221_), .B(ori_ori_n36_), .Y(ori_ori_n511_));
  NO2        o489(.A(ori_ori_n379_), .B(i_1_), .Y(ori_ori_n512_));
  NOi31      o490(.An(ori_ori_n512_), .B(ori_ori_n417_), .C(ori_ori_n73_), .Y(ori_ori_n513_));
  AN4        o491(.A(ori_ori_n513_), .B(ori_ori_n377_), .C(ori_ori_n453_), .D(i_2_), .Y(ori_ori_n514_));
  INV        o492(.A(ori_ori_n514_), .Y(ori_ori_n515_));
  NOi21      o493(.An(i_10_), .B(i_6_), .Y(ori_ori_n516_));
  NO2        o494(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n517_));
  AOI220     o495(.A0(ori_ori_n267_), .A1(ori_ori_n517_), .B0(ori_ori_n258_), .B1(ori_ori_n516_), .Y(ori_ori_n518_));
  NO2        o496(.A(ori_ori_n518_), .B(ori_ori_n415_), .Y(ori_ori_n519_));
  NO2        o497(.A(ori_ori_n117_), .B(ori_ori_n23_), .Y(ori_ori_n520_));
  NA2        o498(.A(ori_ori_n294_), .B(ori_ori_n165_), .Y(ori_ori_n521_));
  AOI220     o499(.A0(ori_ori_n521_), .A1(ori_ori_n397_), .B0(ori_ori_n181_), .B1(ori_ori_n179_), .Y(ori_ori_n522_));
  NO2        o500(.A(ori_ori_n193_), .B(ori_ori_n37_), .Y(ori_ori_n523_));
  NOi31      o501(.An(ori_ori_n149_), .B(ori_ori_n523_), .C(ori_ori_n308_), .Y(ori_ori_n524_));
  NO3        o502(.A(ori_ori_n524_), .B(ori_ori_n522_), .C(ori_ori_n519_), .Y(ori_ori_n525_));
  NO2        o503(.A(ori_ori_n469_), .B(ori_ori_n346_), .Y(ori_ori_n526_));
  INV        o504(.A(ori_ori_n297_), .Y(ori_ori_n527_));
  NO2        o505(.A(i_12_), .B(ori_ori_n86_), .Y(ori_ori_n528_));
  NA3        o506(.A(ori_ori_n528_), .B(ori_ori_n258_), .C(ori_ori_n505_), .Y(ori_ori_n529_));
  NA3        o507(.A(ori_ori_n354_), .B(ori_ori_n267_), .C(ori_ori_n209_), .Y(ori_ori_n530_));
  AOI210     o508(.A0(ori_ori_n530_), .A1(ori_ori_n529_), .B0(ori_ori_n527_), .Y(ori_ori_n531_));
  OR2        o509(.A(i_2_), .B(i_5_), .Y(ori_ori_n532_));
  OR2        o510(.A(ori_ori_n532_), .B(ori_ori_n374_), .Y(ori_ori_n533_));
  AOI210     o511(.A0(ori_ori_n340_), .A1(ori_ori_n230_), .B0(ori_ori_n193_), .Y(ori_ori_n534_));
  AOI210     o512(.A0(ori_ori_n534_), .A1(ori_ori_n533_), .B0(ori_ori_n451_), .Y(ori_ori_n535_));
  NO3        o513(.A(ori_ori_n535_), .B(ori_ori_n531_), .C(ori_ori_n526_), .Y(ori_ori_n536_));
  NA4        o514(.A(ori_ori_n536_), .B(ori_ori_n525_), .C(ori_ori_n515_), .D(ori_ori_n508_), .Y(ori_ori_n537_));
  NO4        o515(.A(ori_ori_n537_), .B(ori_ori_n497_), .C(ori_ori_n479_), .D(ori_ori_n462_), .Y(ori_ori_n538_));
  NA4        o516(.A(ori_ori_n538_), .B(ori_ori_n404_), .C(ori_ori_n323_), .D(ori_ori_n290_), .Y(ori7));
  NO2        o517(.A(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n540_));
  NO2        o518(.A(ori_ori_n111_), .B(ori_ori_n92_), .Y(ori_ori_n541_));
  NA2        o519(.A(ori_ori_n352_), .B(ori_ori_n541_), .Y(ori_ori_n542_));
  NA2        o520(.A(ori_ori_n440_), .B(ori_ori_n84_), .Y(ori_ori_n543_));
  NA2        o521(.A(i_11_), .B(ori_ori_n189_), .Y(ori_ori_n544_));
  NA2        o522(.A(ori_ori_n147_), .B(ori_ori_n544_), .Y(ori_ori_n545_));
  OAI210     o523(.A0(ori_ori_n545_), .A1(ori_ori_n543_), .B0(ori_ori_n542_), .Y(ori_ori_n546_));
  NA3        o524(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n547_));
  NO2        o525(.A(ori_ori_n223_), .B(i_4_), .Y(ori_ori_n548_));
  NA2        o526(.A(ori_ori_n548_), .B(i_8_), .Y(ori_ori_n549_));
  NO2        o527(.A(ori_ori_n108_), .B(ori_ori_n547_), .Y(ori_ori_n550_));
  NA2        o528(.A(i_2_), .B(ori_ori_n86_), .Y(ori_ori_n551_));
  OAI210     o529(.A0(ori_ori_n89_), .A1(ori_ori_n195_), .B0(ori_ori_n196_), .Y(ori_ori_n552_));
  NO2        o530(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n553_));
  NA2        o531(.A(i_4_), .B(i_8_), .Y(ori_ori_n554_));
  AOI210     o532(.A0(ori_ori_n554_), .A1(ori_ori_n286_), .B0(ori_ori_n553_), .Y(ori_ori_n555_));
  OAI220     o533(.A0(ori_ori_n555_), .A1(ori_ori_n551_), .B0(ori_ori_n552_), .B1(i_13_), .Y(ori_ori_n556_));
  NO4        o534(.A(ori_ori_n556_), .B(ori_ori_n550_), .C(ori_ori_n546_), .D(ori_ori_n540_), .Y(ori_ori_n557_));
  AOI210     o535(.A0(ori_ori_n131_), .A1(ori_ori_n62_), .B0(i_10_), .Y(ori_ori_n558_));
  AOI210     o536(.A0(ori_ori_n558_), .A1(ori_ori_n223_), .B0(ori_ori_n162_), .Y(ori_ori_n559_));
  OR2        o537(.A(i_6_), .B(i_10_), .Y(ori_ori_n560_));
  NO2        o538(.A(ori_ori_n560_), .B(ori_ori_n23_), .Y(ori_ori_n561_));
  OR3        o539(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n562_));
  INV        o540(.A(ori_ori_n194_), .Y(ori_ori_n563_));
  INV        o541(.A(ori_ori_n561_), .Y(ori_ori_n564_));
  OA220      o542(.A0(ori_ori_n564_), .A1(ori_ori_n527_), .B0(ori_ori_n559_), .B1(ori_ori_n250_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n565_), .A1(ori_ori_n557_), .B0(ori_ori_n63_), .Y(ori_ori_n566_));
  NOi21      o544(.An(i_11_), .B(i_7_), .Y(ori_ori_n567_));
  AO210      o545(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n568_));
  NO2        o546(.A(ori_ori_n568_), .B(ori_ori_n567_), .Y(ori_ori_n569_));
  NA2        o547(.A(ori_ori_n569_), .B(ori_ori_n200_), .Y(ori_ori_n570_));
  NA3        o548(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n571_));
  NAi31      o549(.An(ori_ori_n571_), .B(ori_ori_n207_), .C(i_11_), .Y(ori_ori_n572_));
  AOI210     o550(.A0(ori_ori_n572_), .A1(ori_ori_n570_), .B0(ori_ori_n63_), .Y(ori_ori_n573_));
  NA2        o551(.A(ori_ori_n88_), .B(ori_ori_n63_), .Y(ori_ori_n574_));
  AO210      o552(.A0(ori_ori_n574_), .A1(ori_ori_n346_), .B0(ori_ori_n41_), .Y(ori_ori_n575_));
  NO3        o553(.A(ori_ori_n240_), .B(ori_ori_n201_), .C(ori_ori_n544_), .Y(ori_ori_n576_));
  OAI210     o554(.A0(ori_ori_n576_), .A1(ori_ori_n216_), .B0(ori_ori_n63_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n375_), .B(ori_ori_n31_), .Y(ori_ori_n578_));
  OR2        o556(.A(ori_ori_n201_), .B(ori_ori_n111_), .Y(ori_ori_n579_));
  NA2        o557(.A(ori_ori_n579_), .B(ori_ori_n578_), .Y(ori_ori_n580_));
  NO2        o558(.A(i_1_), .B(i_4_), .Y(ori_ori_n581_));
  NA2        o559(.A(ori_ori_n581_), .B(ori_ori_n580_), .Y(ori_ori_n582_));
  NO2        o560(.A(i_1_), .B(i_12_), .Y(ori_ori_n583_));
  NA3        o561(.A(ori_ori_n583_), .B(ori_ori_n112_), .C(ori_ori_n24_), .Y(ori_ori_n584_));
  BUFFER     o562(.A(ori_ori_n584_), .Y(ori_ori_n585_));
  NA4        o563(.A(ori_ori_n585_), .B(ori_ori_n582_), .C(ori_ori_n577_), .D(ori_ori_n575_), .Y(ori_ori_n586_));
  OAI210     o564(.A0(ori_ori_n586_), .A1(ori_ori_n573_), .B0(i_6_), .Y(ori_ori_n587_));
  NO2        o565(.A(ori_ori_n571_), .B(ori_ori_n111_), .Y(ori_ori_n588_));
  NA2        o566(.A(ori_ori_n588_), .B(ori_ori_n528_), .Y(ori_ori_n589_));
  NO2        o567(.A(ori_ori_n223_), .B(ori_ori_n86_), .Y(ori_ori_n590_));
  NO2        o568(.A(ori_ori_n590_), .B(i_11_), .Y(ori_ori_n591_));
  NA2        o569(.A(ori_ori_n589_), .B(ori_ori_n418_), .Y(ori_ori_n592_));
  NO3        o570(.A(ori_ori_n560_), .B(ori_ori_n221_), .C(ori_ori_n23_), .Y(ori_ori_n593_));
  AOI210     o571(.A0(i_1_), .A1(ori_ori_n241_), .B0(ori_ori_n593_), .Y(ori_ori_n594_));
  NO2        o572(.A(ori_ori_n594_), .B(ori_ori_n44_), .Y(ori_ori_n595_));
  NA3        o573(.A(ori_ori_n481_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n596_));
  INV        o574(.A(i_2_), .Y(ori_ori_n597_));
  NA2        o575(.A(ori_ori_n141_), .B(i_9_), .Y(ori_ori_n598_));
  NA3        o576(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n599_));
  NO2        o577(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n600_));
  NA3        o578(.A(ori_ori_n600_), .B(ori_ori_n249_), .C(ori_ori_n44_), .Y(ori_ori_n601_));
  OAI220     o579(.A0(ori_ori_n601_), .A1(ori_ori_n599_), .B0(ori_ori_n598_), .B1(ori_ori_n597_), .Y(ori_ori_n602_));
  AOI210     o580(.A0(ori_ori_n437_), .A1(ori_ori_n382_), .B0(ori_ori_n227_), .Y(ori_ori_n603_));
  NO2        o581(.A(ori_ori_n603_), .B(ori_ori_n551_), .Y(ori_ori_n604_));
  NAi21      o582(.An(ori_ori_n596_), .B(ori_ori_n94_), .Y(ori_ori_n605_));
  NA2        o583(.A(ori_ori_n600_), .B(ori_ori_n249_), .Y(ori_ori_n606_));
  NO2        o584(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n607_));
  NA2        o585(.A(ori_ori_n607_), .B(ori_ori_n24_), .Y(ori_ori_n608_));
  OAI210     o586(.A0(ori_ori_n608_), .A1(ori_ori_n606_), .B0(ori_ori_n605_), .Y(ori_ori_n609_));
  OR3        o587(.A(ori_ori_n609_), .B(ori_ori_n604_), .C(ori_ori_n602_), .Y(ori_ori_n610_));
  NO3        o588(.A(ori_ori_n610_), .B(ori_ori_n595_), .C(ori_ori_n592_), .Y(ori_ori_n611_));
  NO2        o589(.A(ori_ori_n223_), .B(ori_ori_n104_), .Y(ori_ori_n612_));
  NO2        o590(.A(ori_ori_n612_), .B(ori_ori_n567_), .Y(ori_ori_n613_));
  NA2        o591(.A(ori_ori_n613_), .B(i_1_), .Y(ori_ori_n614_));
  NO2        o592(.A(ori_ori_n614_), .B(ori_ori_n562_), .Y(ori_ori_n615_));
  NO2        o593(.A(ori_ori_n378_), .B(ori_ori_n86_), .Y(ori_ori_n616_));
  NA2        o594(.A(ori_ori_n615_), .B(ori_ori_n46_), .Y(ori_ori_n617_));
  NA2        o595(.A(i_3_), .B(ori_ori_n189_), .Y(ori_ori_n618_));
  NO2        o596(.A(ori_ori_n618_), .B(ori_ori_n117_), .Y(ori_ori_n619_));
  AN2        o597(.A(ori_ori_n619_), .B(ori_ori_n486_), .Y(ori_ori_n620_));
  NO2        o598(.A(ori_ori_n221_), .B(ori_ori_n44_), .Y(ori_ori_n621_));
  NO3        o599(.A(ori_ori_n621_), .B(ori_ori_n288_), .C(ori_ori_n224_), .Y(ori_ori_n622_));
  NO2        o600(.A(ori_ori_n120_), .B(ori_ori_n37_), .Y(ori_ori_n623_));
  NO2        o601(.A(ori_ori_n623_), .B(i_6_), .Y(ori_ori_n624_));
  NO2        o602(.A(ori_ori_n86_), .B(i_9_), .Y(ori_ori_n625_));
  NO2        o603(.A(ori_ori_n625_), .B(ori_ori_n63_), .Y(ori_ori_n626_));
  NO2        o604(.A(ori_ori_n626_), .B(ori_ori_n583_), .Y(ori_ori_n627_));
  NO4        o605(.A(ori_ori_n627_), .B(ori_ori_n624_), .C(ori_ori_n622_), .D(i_4_), .Y(ori_ori_n628_));
  NA2        o606(.A(i_1_), .B(i_3_), .Y(ori_ori_n629_));
  NO2        o607(.A(ori_ori_n419_), .B(ori_ori_n95_), .Y(ori_ori_n630_));
  AOI210     o608(.A0(ori_ori_n621_), .A1(ori_ori_n516_), .B0(ori_ori_n630_), .Y(ori_ori_n631_));
  NO2        o609(.A(ori_ori_n631_), .B(ori_ori_n629_), .Y(ori_ori_n632_));
  NO3        o610(.A(ori_ori_n632_), .B(ori_ori_n628_), .C(ori_ori_n620_), .Y(ori_ori_n633_));
  NA4        o611(.A(ori_ori_n633_), .B(ori_ori_n617_), .C(ori_ori_n611_), .D(ori_ori_n587_), .Y(ori_ori_n634_));
  NO3        o612(.A(ori_ori_n438_), .B(i_3_), .C(i_7_), .Y(ori_ori_n635_));
  NOi21      o613(.An(ori_ori_n635_), .B(i_10_), .Y(ori_ori_n636_));
  OA210      o614(.A0(ori_ori_n636_), .A1(ori_ori_n231_), .B0(ori_ori_n86_), .Y(ori_ori_n637_));
  NO3        o615(.A(ori_ori_n439_), .B(ori_ori_n554_), .C(ori_ori_n86_), .Y(ori_ori_n638_));
  NA2        o616(.A(ori_ori_n638_), .B(ori_ori_n25_), .Y(ori_ori_n639_));
  INV        o617(.A(ori_ori_n639_), .Y(ori_ori_n640_));
  OAI210     o618(.A0(ori_ori_n640_), .A1(ori_ori_n637_), .B0(i_1_), .Y(ori_ori_n641_));
  AOI210     o619(.A0(ori_ori_n249_), .A1(ori_ori_n100_), .B0(i_1_), .Y(ori_ori_n642_));
  NO2        o620(.A(ori_ori_n336_), .B(i_2_), .Y(ori_ori_n643_));
  NA2        o621(.A(ori_ori_n643_), .B(ori_ori_n642_), .Y(ori_ori_n644_));
  AOI210     o622(.A0(ori_ori_n644_), .A1(ori_ori_n641_), .B0(i_13_), .Y(ori_ori_n645_));
  OR2        o623(.A(i_11_), .B(i_7_), .Y(ori_ori_n646_));
  NA3        o624(.A(ori_ori_n646_), .B(ori_ori_n109_), .C(ori_ori_n141_), .Y(ori_ori_n647_));
  AOI220     o625(.A0(ori_ori_n433_), .A1(ori_ori_n162_), .B0(ori_ori_n412_), .B1(ori_ori_n141_), .Y(ori_ori_n648_));
  OAI210     o626(.A0(ori_ori_n648_), .A1(ori_ori_n44_), .B0(ori_ori_n647_), .Y(ori_ori_n649_));
  AOI210     o627(.A0(ori_ori_n599_), .A1(ori_ori_n54_), .B0(i_12_), .Y(ori_ori_n650_));
  NO2        o628(.A(ori_ori_n439_), .B(ori_ori_n24_), .Y(ori_ori_n651_));
  NA2        o629(.A(ori_ori_n651_), .B(ori_ori_n616_), .Y(ori_ori_n652_));
  OAI220     o630(.A0(ori_ori_n652_), .A1(ori_ori_n41_), .B0(ori_ori_n973_), .B1(ori_ori_n95_), .Y(ori_ori_n653_));
  AOI210     o631(.A0(ori_ori_n649_), .A1(ori_ori_n310_), .B0(ori_ori_n653_), .Y(ori_ori_n654_));
  NA2        o632(.A(ori_ori_n354_), .B(ori_ori_n600_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n655_), .B(ori_ori_n228_), .Y(ori_ori_n656_));
  AOI210     o634(.A0(ori_ori_n409_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n657_));
  NOi31      o635(.An(ori_ori_n657_), .B(ori_ori_n543_), .C(ori_ori_n44_), .Y(ori_ori_n658_));
  NA2        o636(.A(ori_ori_n130_), .B(i_13_), .Y(ori_ori_n659_));
  NO2        o637(.A(ori_ori_n599_), .B(ori_ori_n117_), .Y(ori_ori_n660_));
  INV        o638(.A(ori_ori_n660_), .Y(ori_ori_n661_));
  OAI220     o639(.A0(ori_ori_n661_), .A1(ori_ori_n71_), .B0(ori_ori_n659_), .B1(ori_ori_n642_), .Y(ori_ori_n662_));
  NO3        o640(.A(ori_ori_n71_), .B(ori_ori_n32_), .C(ori_ori_n104_), .Y(ori_ori_n663_));
  NA2        o641(.A(ori_ori_n26_), .B(ori_ori_n189_), .Y(ori_ori_n664_));
  NA2        o642(.A(ori_ori_n664_), .B(i_7_), .Y(ori_ori_n665_));
  INV        o643(.A(ori_ori_n663_), .Y(ori_ori_n666_));
  AOI220     o644(.A0(ori_ori_n354_), .A1(ori_ori_n600_), .B0(ori_ori_n94_), .B1(ori_ori_n105_), .Y(ori_ori_n667_));
  OAI220     o645(.A0(ori_ori_n667_), .A1(ori_ori_n549_), .B0(ori_ori_n666_), .B1(ori_ori_n563_), .Y(ori_ori_n668_));
  NO4        o646(.A(ori_ori_n668_), .B(ori_ori_n662_), .C(ori_ori_n658_), .D(ori_ori_n656_), .Y(ori_ori_n669_));
  OR2        o647(.A(i_11_), .B(i_6_), .Y(ori_ori_n670_));
  NA3        o648(.A(ori_ori_n548_), .B(ori_ori_n664_), .C(i_7_), .Y(ori_ori_n671_));
  AOI210     o649(.A0(ori_ori_n671_), .A1(ori_ori_n661_), .B0(ori_ori_n670_), .Y(ori_ori_n672_));
  NA3        o650(.A(ori_ori_n375_), .B(ori_ori_n553_), .C(ori_ori_n100_), .Y(ori_ori_n673_));
  NA2        o651(.A(ori_ori_n591_), .B(i_13_), .Y(ori_ori_n674_));
  NA2        o652(.A(ori_ori_n105_), .B(ori_ori_n664_), .Y(ori_ori_n675_));
  NAi21      o653(.An(i_11_), .B(i_12_), .Y(ori_ori_n676_));
  NOi41      o654(.An(ori_ori_n113_), .B(ori_ori_n676_), .C(i_13_), .D(ori_ori_n86_), .Y(ori_ori_n677_));
  NO3        o655(.A(ori_ori_n439_), .B(ori_ori_n528_), .C(ori_ori_n554_), .Y(ori_ori_n678_));
  AOI220     o656(.A0(ori_ori_n678_), .A1(ori_ori_n291_), .B0(ori_ori_n677_), .B1(ori_ori_n675_), .Y(ori_ori_n679_));
  NA3        o657(.A(ori_ori_n679_), .B(ori_ori_n674_), .C(ori_ori_n673_), .Y(ori_ori_n680_));
  OAI210     o658(.A0(ori_ori_n680_), .A1(ori_ori_n672_), .B0(ori_ori_n63_), .Y(ori_ori_n681_));
  NO2        o659(.A(i_2_), .B(i_12_), .Y(ori_ori_n682_));
  NA2        o660(.A(ori_ori_n335_), .B(ori_ori_n682_), .Y(ori_ori_n683_));
  NA2        o661(.A(ori_ori_n337_), .B(ori_ori_n335_), .Y(ori_ori_n684_));
  NO2        o662(.A(ori_ori_n131_), .B(i_2_), .Y(ori_ori_n685_));
  NA2        o663(.A(ori_ori_n685_), .B(ori_ori_n583_), .Y(ori_ori_n686_));
  NA3        o664(.A(ori_ori_n686_), .B(ori_ori_n684_), .C(ori_ori_n683_), .Y(ori_ori_n687_));
  NA3        o665(.A(ori_ori_n687_), .B(ori_ori_n45_), .C(ori_ori_n215_), .Y(ori_ori_n688_));
  NA4        o666(.A(ori_ori_n688_), .B(ori_ori_n681_), .C(ori_ori_n669_), .D(ori_ori_n654_), .Y(ori_ori_n689_));
  OR4        o667(.A(ori_ori_n689_), .B(ori_ori_n645_), .C(ori_ori_n634_), .D(ori_ori_n566_), .Y(ori5));
  NA2        o668(.A(ori_ori_n613_), .B(ori_ori_n252_), .Y(ori_ori_n691_));
  AN2        o669(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n692_));
  NA3        o670(.A(ori_ori_n692_), .B(ori_ori_n682_), .C(ori_ori_n111_), .Y(ori_ori_n693_));
  NO2        o671(.A(ori_ori_n549_), .B(i_11_), .Y(ori_ori_n694_));
  NA2        o672(.A(ori_ori_n89_), .B(ori_ori_n694_), .Y(ori_ori_n695_));
  NA3        o673(.A(ori_ori_n695_), .B(ori_ori_n693_), .C(ori_ori_n691_), .Y(ori_ori_n696_));
  NO3        o674(.A(i_11_), .B(ori_ori_n223_), .C(i_13_), .Y(ori_ori_n697_));
  NO2        o675(.A(ori_ori_n127_), .B(ori_ori_n23_), .Y(ori_ori_n698_));
  NA2        o676(.A(i_12_), .B(i_8_), .Y(ori_ori_n699_));
  OAI210     o677(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n699_), .Y(ori_ori_n700_));
  INV        o678(.A(ori_ori_n408_), .Y(ori_ori_n701_));
  AOI220     o679(.A0(ori_ori_n297_), .A1(ori_ori_n520_), .B0(ori_ori_n700_), .B1(ori_ori_n698_), .Y(ori_ori_n702_));
  INV        o680(.A(ori_ori_n702_), .Y(ori_ori_n703_));
  NO2        o681(.A(ori_ori_n703_), .B(ori_ori_n696_), .Y(ori_ori_n704_));
  INV        o682(.A(ori_ori_n172_), .Y(ori_ori_n705_));
  INV        o683(.A(ori_ori_n231_), .Y(ori_ori_n706_));
  OAI210     o684(.A0(ori_ori_n643_), .A1(ori_ori_n410_), .B0(ori_ori_n113_), .Y(ori_ori_n707_));
  AOI210     o685(.A0(ori_ori_n707_), .A1(ori_ori_n706_), .B0(ori_ori_n705_), .Y(ori_ori_n708_));
  NO2        o686(.A(ori_ori_n419_), .B(ori_ori_n26_), .Y(ori_ori_n709_));
  NO2        o687(.A(ori_ori_n709_), .B(ori_ori_n382_), .Y(ori_ori_n710_));
  NA2        o688(.A(ori_ori_n710_), .B(i_2_), .Y(ori_ori_n711_));
  INV        o689(.A(ori_ori_n711_), .Y(ori_ori_n712_));
  AOI210     o690(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n379_), .Y(ori_ori_n713_));
  AOI210     o691(.A0(ori_ori_n713_), .A1(ori_ori_n712_), .B0(ori_ori_n708_), .Y(ori_ori_n714_));
  NO2        o692(.A(ori_ori_n187_), .B(ori_ori_n128_), .Y(ori_ori_n715_));
  OAI210     o693(.A0(ori_ori_n715_), .A1(ori_ori_n698_), .B0(i_2_), .Y(ori_ori_n716_));
  INV        o694(.A(ori_ori_n173_), .Y(ori_ori_n717_));
  NO3        o695(.A(ori_ori_n568_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n718_));
  AOI210     o696(.A0(ori_ori_n717_), .A1(ori_ori_n89_), .B0(ori_ori_n718_), .Y(ori_ori_n719_));
  AOI210     o697(.A0(ori_ori_n719_), .A1(ori_ori_n716_), .B0(ori_ori_n189_), .Y(ori_ori_n720_));
  OA210      o698(.A0(ori_ori_n569_), .A1(ori_ori_n129_), .B0(i_13_), .Y(ori_ori_n721_));
  NA2        o699(.A(ori_ori_n194_), .B(ori_ori_n195_), .Y(ori_ori_n722_));
  NA2        o700(.A(ori_ori_n154_), .B(ori_ori_n544_), .Y(ori_ori_n723_));
  AOI210     o701(.A0(ori_ori_n723_), .A1(ori_ori_n722_), .B0(ori_ori_n340_), .Y(ori_ori_n724_));
  AOI210     o702(.A0(ori_ori_n201_), .A1(ori_ori_n151_), .B0(ori_ori_n472_), .Y(ori_ori_n725_));
  NA2        o703(.A(ori_ori_n725_), .B(ori_ori_n382_), .Y(ori_ori_n726_));
  NO2        o704(.A(ori_ori_n105_), .B(ori_ori_n44_), .Y(ori_ori_n727_));
  INV        o705(.A(ori_ori_n284_), .Y(ori_ori_n728_));
  NA4        o706(.A(ori_ori_n728_), .B(ori_ori_n286_), .C(ori_ori_n127_), .D(ori_ori_n42_), .Y(ori_ori_n729_));
  OAI210     o707(.A0(ori_ori_n729_), .A1(ori_ori_n727_), .B0(ori_ori_n726_), .Y(ori_ori_n730_));
  NO4        o708(.A(ori_ori_n730_), .B(ori_ori_n724_), .C(ori_ori_n721_), .D(ori_ori_n720_), .Y(ori_ori_n731_));
  NA2        o709(.A(ori_ori_n520_), .B(ori_ori_n28_), .Y(ori_ori_n732_));
  NA2        o710(.A(ori_ori_n697_), .B(ori_ori_n259_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n733_), .B(ori_ori_n732_), .Y(ori_ori_n734_));
  NO2        o712(.A(ori_ori_n62_), .B(i_12_), .Y(ori_ori_n735_));
  NO2        o713(.A(ori_ori_n735_), .B(ori_ori_n129_), .Y(ori_ori_n736_));
  NO2        o714(.A(ori_ori_n736_), .B(ori_ori_n544_), .Y(ori_ori_n737_));
  AOI220     o715(.A0(ori_ori_n737_), .A1(ori_ori_n36_), .B0(ori_ori_n734_), .B1(ori_ori_n46_), .Y(ori_ori_n738_));
  NA4        o716(.A(ori_ori_n738_), .B(ori_ori_n731_), .C(ori_ori_n714_), .D(ori_ori_n704_), .Y(ori6));
  NO3        o717(.A(i_9_), .B(ori_ori_n287_), .C(i_1_), .Y(ori_ori_n740_));
  NA2        o718(.A(ori_ori_n740_), .B(ori_ori_n685_), .Y(ori_ori_n741_));
  NO2        o719(.A(ori_ori_n210_), .B(ori_ori_n442_), .Y(ori_ori_n742_));
  INV        o720(.A(ori_ori_n305_), .Y(ori_ori_n743_));
  AO210      o721(.A0(ori_ori_n743_), .A1(ori_ori_n741_), .B0(i_12_), .Y(ori_ori_n744_));
  NA2        o722(.A(ori_ori_n528_), .B(ori_ori_n63_), .Y(ori_ori_n745_));
  NA2        o723(.A(ori_ori_n636_), .B(ori_ori_n71_), .Y(ori_ori_n746_));
  BUFFER     o724(.A(ori_ori_n574_), .Y(ori_ori_n747_));
  NA3        o725(.A(ori_ori_n747_), .B(ori_ori_n746_), .C(ori_ori_n745_), .Y(ori_ori_n748_));
  NA2        o726(.A(ori_ori_n748_), .B(ori_ori_n73_), .Y(ori_ori_n749_));
  INV        o727(.A(ori_ori_n304_), .Y(ori_ori_n750_));
  NA2        o728(.A(ori_ori_n75_), .B(ori_ori_n134_), .Y(ori_ori_n751_));
  INV        o729(.A(ori_ori_n127_), .Y(ori_ori_n752_));
  NA2        o730(.A(ori_ori_n752_), .B(ori_ori_n46_), .Y(ori_ori_n753_));
  AOI210     o731(.A0(ori_ori_n753_), .A1(ori_ori_n751_), .B0(ori_ori_n750_), .Y(ori_ori_n754_));
  NO3        o732(.A(ori_ori_n234_), .B(ori_ori_n135_), .C(i_9_), .Y(ori_ori_n755_));
  NA2        o733(.A(ori_ori_n755_), .B(ori_ori_n735_), .Y(ori_ori_n756_));
  AOI210     o734(.A0(ori_ori_n756_), .A1(ori_ori_n470_), .B0(ori_ori_n183_), .Y(ori_ori_n757_));
  NO2        o735(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n758_));
  NA3        o736(.A(ori_ori_n758_), .B(ori_ori_n436_), .C(ori_ori_n358_), .Y(ori_ori_n759_));
  NAi32      o737(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n760_));
  NO2        o738(.A(ori_ori_n670_), .B(ori_ori_n760_), .Y(ori_ori_n761_));
  OAI210     o739(.A0(ori_ori_n635_), .A1(ori_ori_n511_), .B0(ori_ori_n510_), .Y(ori_ori_n762_));
  NAi31      o740(.An(ori_ori_n761_), .B(ori_ori_n762_), .C(ori_ori_n759_), .Y(ori_ori_n763_));
  OR3        o741(.A(ori_ori_n763_), .B(ori_ori_n757_), .C(ori_ori_n754_), .Y(ori_ori_n764_));
  NO2        o742(.A(ori_ori_n646_), .B(i_2_), .Y(ori_ori_n765_));
  NA2        o743(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n766_));
  NO2        o744(.A(ori_ori_n766_), .B(ori_ori_n374_), .Y(ori_ori_n767_));
  NA2        o745(.A(ori_ori_n767_), .B(ori_ori_n765_), .Y(ori_ori_n768_));
  OR2        o746(.A(ori_ori_n569_), .B(ori_ori_n410_), .Y(ori_ori_n769_));
  NA3        o747(.A(ori_ori_n769_), .B(ori_ori_n150_), .C(ori_ori_n69_), .Y(ori_ori_n770_));
  AO210      o748(.A0(ori_ori_n449_), .A1(ori_ori_n701_), .B0(ori_ori_n36_), .Y(ori_ori_n771_));
  NA3        o749(.A(ori_ori_n771_), .B(ori_ori_n770_), .C(ori_ori_n768_), .Y(ori_ori_n772_));
  OAI210     o750(.A0(ori_ori_n590_), .A1(i_11_), .B0(ori_ori_n87_), .Y(ori_ori_n773_));
  AOI220     o751(.A0(ori_ori_n773_), .A1(ori_ori_n510_), .B0(ori_ori_n742_), .B1(ori_ori_n665_), .Y(ori_ori_n774_));
  NA3        o752(.A(ori_ori_n340_), .B(ori_ori_n225_), .C(ori_ori_n150_), .Y(ori_ori_n775_));
  NA2        o753(.A(ori_ori_n366_), .B(ori_ori_n70_), .Y(ori_ori_n776_));
  NA4        o754(.A(ori_ori_n776_), .B(ori_ori_n775_), .C(ori_ori_n774_), .D(ori_ori_n552_), .Y(ori_ori_n777_));
  AO210      o755(.A0(ori_ori_n472_), .A1(ori_ori_n46_), .B0(ori_ori_n88_), .Y(ori_ori_n778_));
  NA3        o756(.A(ori_ori_n778_), .B(ori_ori_n440_), .C(ori_ori_n209_), .Y(ori_ori_n779_));
  AOI210     o757(.A0(ori_ori_n410_), .A1(ori_ori_n408_), .B0(ori_ori_n509_), .Y(ori_ori_n780_));
  NO2        o758(.A(ori_ori_n560_), .B(ori_ori_n105_), .Y(ori_ori_n781_));
  OAI210     o759(.A0(ori_ori_n781_), .A1(ori_ori_n114_), .B0(ori_ori_n373_), .Y(ori_ori_n782_));
  NA2        o760(.A(ori_ori_n230_), .B(ori_ori_n46_), .Y(ori_ori_n783_));
  INV        o761(.A(ori_ori_n533_), .Y(ori_ori_n784_));
  NA3        o762(.A(ori_ori_n784_), .B(ori_ori_n304_), .C(i_7_), .Y(ori_ori_n785_));
  NA4        o763(.A(ori_ori_n785_), .B(ori_ori_n782_), .C(ori_ori_n780_), .D(ori_ori_n779_), .Y(ori_ori_n786_));
  NO4        o764(.A(ori_ori_n786_), .B(ori_ori_n777_), .C(ori_ori_n772_), .D(ori_ori_n764_), .Y(ori_ori_n787_));
  NA4        o765(.A(ori_ori_n787_), .B(ori_ori_n749_), .C(ori_ori_n744_), .D(ori_ori_n348_), .Y(ori3));
  NA2        o766(.A(i_12_), .B(i_10_), .Y(ori_ori_n789_));
  NO2        o767(.A(i_11_), .B(ori_ori_n223_), .Y(ori_ori_n790_));
  NA3        o768(.A(ori_ori_n775_), .B(ori_ori_n552_), .C(ori_ori_n339_), .Y(ori_ori_n791_));
  NA2        o769(.A(ori_ori_n791_), .B(ori_ori_n40_), .Y(ori_ori_n792_));
  NOi21      o770(.An(ori_ori_n99_), .B(ori_ori_n710_), .Y(ori_ori_n793_));
  NO3        o771(.A(ori_ori_n579_), .B(ori_ori_n419_), .C(ori_ori_n134_), .Y(ori_ori_n794_));
  NA2        o772(.A(ori_ori_n375_), .B(ori_ori_n45_), .Y(ori_ori_n795_));
  AN2        o773(.A(ori_ori_n417_), .B(ori_ori_n55_), .Y(ori_ori_n796_));
  NO3        o774(.A(ori_ori_n796_), .B(ori_ori_n794_), .C(ori_ori_n793_), .Y(ori_ori_n797_));
  AOI210     o775(.A0(ori_ori_n797_), .A1(ori_ori_n792_), .B0(ori_ori_n48_), .Y(ori_ori_n798_));
  NO4        o776(.A(ori_ori_n344_), .B(ori_ori_n351_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n799_));
  NA2        o777(.A(ori_ori_n183_), .B(ori_ori_n516_), .Y(ori_ori_n800_));
  NOi21      o778(.An(ori_ori_n800_), .B(ori_ori_n799_), .Y(ori_ori_n801_));
  NA2        o779(.A(ori_ori_n657_), .B(ori_ori_n625_), .Y(ori_ori_n802_));
  NA2        o780(.A(ori_ori_n311_), .B(ori_ori_n399_), .Y(ori_ori_n803_));
  OAI220     o781(.A0(ori_ori_n803_), .A1(ori_ori_n802_), .B0(ori_ori_n801_), .B1(ori_ori_n63_), .Y(ori_ori_n804_));
  NOi21      o782(.An(i_5_), .B(i_9_), .Y(ori_ori_n805_));
  NA2        o783(.A(ori_ori_n805_), .B(ori_ori_n406_), .Y(ori_ori_n806_));
  BUFFER     o784(.A(ori_ori_n249_), .Y(ori_ori_n807_));
  AOI210     o785(.A0(ori_ori_n807_), .A1(ori_ori_n437_), .B0(ori_ori_n638_), .Y(ori_ori_n808_));
  NO3        o786(.A(ori_ori_n376_), .B(ori_ori_n249_), .C(ori_ori_n73_), .Y(ori_ori_n809_));
  NO2        o787(.A(ori_ori_n175_), .B(ori_ori_n151_), .Y(ori_ori_n810_));
  AOI210     o788(.A0(ori_ori_n810_), .A1(ori_ori_n230_), .B0(ori_ori_n809_), .Y(ori_ori_n811_));
  OAI220     o789(.A0(ori_ori_n811_), .A1(ori_ori_n178_), .B0(ori_ori_n808_), .B1(ori_ori_n806_), .Y(ori_ori_n812_));
  NO3        o790(.A(ori_ori_n812_), .B(ori_ori_n804_), .C(ori_ori_n798_), .Y(ori_ori_n813_));
  NA2        o791(.A(ori_ori_n183_), .B(ori_ori_n24_), .Y(ori_ori_n814_));
  NO2        o792(.A(ori_ori_n623_), .B(ori_ori_n541_), .Y(ori_ori_n815_));
  NO2        o793(.A(ori_ori_n815_), .B(ori_ori_n814_), .Y(ori_ori_n816_));
  NA2        o794(.A(ori_ori_n291_), .B(ori_ori_n132_), .Y(ori_ori_n817_));
  NAi21      o795(.An(ori_ori_n163_), .B(ori_ori_n399_), .Y(ori_ori_n818_));
  OAI220     o796(.A0(ori_ori_n818_), .A1(ori_ori_n783_), .B0(ori_ori_n817_), .B1(ori_ori_n368_), .Y(ori_ori_n819_));
  NO2        o797(.A(ori_ori_n819_), .B(ori_ori_n816_), .Y(ori_ori_n820_));
  NA2        o798(.A(ori_ori_n517_), .B(i_0_), .Y(ori_ori_n821_));
  NO3        o799(.A(ori_ori_n821_), .B(ori_ori_n353_), .C(ori_ori_n89_), .Y(ori_ori_n822_));
  NO4        o800(.A(ori_ori_n532_), .B(ori_ori_n207_), .C(ori_ori_n379_), .D(ori_ori_n374_), .Y(ori_ori_n823_));
  AOI210     o801(.A0(ori_ori_n823_), .A1(i_11_), .B0(ori_ori_n822_), .Y(ori_ori_n824_));
  INV        o802(.A(ori_ori_n436_), .Y(ori_ori_n825_));
  AN2        o803(.A(ori_ori_n99_), .B(ori_ori_n229_), .Y(ori_ori_n826_));
  NA2        o804(.A(ori_ori_n697_), .B(ori_ori_n305_), .Y(ori_ori_n827_));
  AOI210     o805(.A0(ori_ori_n440_), .A1(ori_ori_n89_), .B0(ori_ori_n58_), .Y(ori_ori_n828_));
  OAI220     o806(.A0(ori_ori_n828_), .A1(ori_ori_n827_), .B0(ori_ori_n608_), .B1(ori_ori_n483_), .Y(ori_ori_n829_));
  NO2        o807(.A(ori_ori_n236_), .B(ori_ori_n155_), .Y(ori_ori_n830_));
  NA2        o808(.A(i_0_), .B(i_10_), .Y(ori_ori_n831_));
  INV        o809(.A(ori_ori_n485_), .Y(ori_ori_n832_));
  NO4        o810(.A(ori_ori_n117_), .B(ori_ori_n58_), .C(ori_ori_n618_), .D(i_5_), .Y(ori_ori_n833_));
  AO220      o811(.A0(ori_ori_n833_), .A1(ori_ori_n832_), .B0(ori_ori_n830_), .B1(i_6_), .Y(ori_ori_n834_));
  NA2        o812(.A(ori_ori_n186_), .B(ori_ori_n195_), .Y(ori_ori_n835_));
  NO2        o813(.A(ori_ori_n835_), .B(ori_ori_n827_), .Y(ori_ori_n836_));
  NO4        o814(.A(ori_ori_n836_), .B(ori_ori_n834_), .C(ori_ori_n829_), .D(ori_ori_n826_), .Y(ori_ori_n837_));
  NA3        o815(.A(ori_ori_n837_), .B(ori_ori_n824_), .C(ori_ori_n820_), .Y(ori_ori_n838_));
  NO2        o816(.A(ori_ori_n106_), .B(ori_ori_n37_), .Y(ori_ori_n839_));
  NA2        o817(.A(i_11_), .B(i_9_), .Y(ori_ori_n840_));
  NO3        o818(.A(i_12_), .B(ori_ori_n840_), .C(ori_ori_n551_), .Y(ori_ori_n841_));
  AN2        o819(.A(ori_ori_n841_), .B(ori_ori_n839_), .Y(ori_ori_n842_));
  NO2        o820(.A(ori_ori_n48_), .B(i_7_), .Y(ori_ori_n843_));
  NA2        o821(.A(ori_ori_n363_), .B(ori_ori_n176_), .Y(ori_ori_n844_));
  NA2        o822(.A(ori_ori_n844_), .B(ori_ori_n161_), .Y(ori_ori_n845_));
  NO2        o823(.A(ori_ori_n840_), .B(ori_ori_n73_), .Y(ori_ori_n846_));
  NO2        o824(.A(ori_ori_n175_), .B(i_0_), .Y(ori_ori_n847_));
  INV        o825(.A(ori_ori_n372_), .Y(ori_ori_n848_));
  NO2        o826(.A(ori_ori_n848_), .B(ori_ori_n806_), .Y(ori_ori_n849_));
  NO3        o827(.A(ori_ori_n849_), .B(ori_ori_n845_), .C(ori_ori_n842_), .Y(ori_ori_n850_));
  NA2        o828(.A(ori_ori_n607_), .B(ori_ori_n124_), .Y(ori_ori_n851_));
  NO2        o829(.A(i_6_), .B(ori_ori_n851_), .Y(ori_ori_n852_));
  AOI210     o830(.A0(ori_ori_n409_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n853_));
  NA2        o831(.A(ori_ori_n172_), .B(ori_ori_n106_), .Y(ori_ori_n854_));
  NOi32      o832(.An(ori_ori_n853_), .Bn(ori_ori_n186_), .C(ori_ori_n854_), .Y(ori_ori_n855_));
  NA2        o833(.A(ori_ori_n553_), .B(ori_ori_n305_), .Y(ori_ori_n856_));
  NO2        o834(.A(ori_ori_n856_), .B(ori_ori_n795_), .Y(ori_ori_n857_));
  NO3        o835(.A(ori_ori_n857_), .B(ori_ori_n855_), .C(ori_ori_n852_), .Y(ori_ori_n858_));
  NOi21      o836(.An(i_7_), .B(i_5_), .Y(ori_ori_n859_));
  OR2        o837(.A(ori_ori_n854_), .B(ori_ori_n470_), .Y(ori_ori_n860_));
  INV        o838(.A(ori_ori_n298_), .Y(ori_ori_n861_));
  NA3        o839(.A(ori_ori_n860_), .B(ori_ori_n858_), .C(ori_ori_n850_), .Y(ori_ori_n862_));
  NO2        o840(.A(ori_ori_n789_), .B(ori_ori_n297_), .Y(ori_ori_n863_));
  OA210      o841(.A0(ori_ori_n436_), .A1(ori_ori_n213_), .B0(ori_ori_n435_), .Y(ori_ori_n864_));
  NA2        o842(.A(ori_ori_n863_), .B(ori_ori_n846_), .Y(ori_ori_n865_));
  NA3        o843(.A(ori_ori_n435_), .B(ori_ori_n375_), .C(ori_ori_n45_), .Y(ori_ori_n866_));
  OAI210     o844(.A0(ori_ori_n818_), .A1(ori_ori_n825_), .B0(ori_ori_n866_), .Y(ori_ori_n867_));
  NO2        o845(.A(i_2_), .B(ori_ori_n185_), .Y(ori_ori_n868_));
  AOI220     o846(.A0(ori_ori_n868_), .A1(ori_ori_n436_), .B0(ori_ori_n867_), .B1(ori_ori_n73_), .Y(ori_ori_n869_));
  NA3        o847(.A(ori_ori_n766_), .B(ori_ori_n350_), .C(ori_ori_n590_), .Y(ori_ori_n870_));
  NA2        o848(.A(ori_ori_n95_), .B(ori_ori_n44_), .Y(ori_ori_n871_));
  NO2        o849(.A(ori_ori_n75_), .B(ori_ori_n699_), .Y(ori_ori_n872_));
  AOI220     o850(.A0(ori_ori_n872_), .A1(ori_ori_n871_), .B0(ori_ori_n174_), .B1(ori_ori_n541_), .Y(ori_ori_n873_));
  AOI210     o851(.A0(ori_ori_n873_), .A1(ori_ori_n870_), .B0(ori_ori_n47_), .Y(ori_ori_n874_));
  NA2        o852(.A(ori_ori_n651_), .B(ori_ori_n493_), .Y(ori_ori_n875_));
  NO2        o853(.A(ori_ori_n875_), .B(ori_ori_n173_), .Y(ori_ori_n876_));
  NO3        o854(.A(ori_ori_n876_), .B(ori_ori_n874_), .C(ori_ori_n474_), .Y(ori_ori_n877_));
  NA3        o855(.A(ori_ori_n877_), .B(ori_ori_n869_), .C(ori_ori_n865_), .Y(ori_ori_n878_));
  NO3        o856(.A(ori_ori_n878_), .B(ori_ori_n862_), .C(ori_ori_n838_), .Y(ori_ori_n879_));
  NO2        o857(.A(i_0_), .B(ori_ori_n676_), .Y(ori_ori_n880_));
  NA2        o858(.A(ori_ori_n73_), .B(ori_ori_n44_), .Y(ori_ori_n881_));
  NO2        o859(.A(ori_ori_n745_), .B(ori_ori_n854_), .Y(ori_ori_n882_));
  INV        o860(.A(ori_ori_n882_), .Y(ori_ori_n883_));
  NO2        o861(.A(ori_ori_n762_), .B(ori_ori_n369_), .Y(ori_ori_n884_));
  NA2        o862(.A(ori_ori_n790_), .B(i_9_), .Y(ori_ori_n885_));
  NO2        o863(.A(ori_ori_n455_), .B(ori_ori_n885_), .Y(ori_ori_n886_));
  OAI210     o864(.A0(ori_ori_n230_), .A1(i_9_), .B0(ori_ori_n220_), .Y(ori_ori_n887_));
  AOI210     o865(.A0(ori_ori_n887_), .A1(ori_ori_n821_), .B0(ori_ori_n155_), .Y(ori_ori_n888_));
  NO3        o866(.A(ori_ori_n888_), .B(ori_ori_n886_), .C(ori_ori_n884_), .Y(ori_ori_n889_));
  NA2        o867(.A(ori_ori_n889_), .B(ori_ori_n883_), .Y(ori_ori_n890_));
  NO3        o868(.A(ori_ori_n831_), .B(ori_ori_n805_), .C(ori_ori_n187_), .Y(ori_ori_n891_));
  AOI220     o869(.A0(ori_ori_n891_), .A1(i_11_), .B0(ori_ori_n513_), .B1(ori_ori_n75_), .Y(ori_ori_n892_));
  NO3        o870(.A(ori_ori_n202_), .B(ori_ori_n351_), .C(i_0_), .Y(ori_ori_n893_));
  OAI210     o871(.A0(ori_ori_n893_), .A1(ori_ori_n76_), .B0(i_13_), .Y(ori_ori_n894_));
  NA2        o872(.A(ori_ori_n894_), .B(ori_ori_n892_), .Y(ori_ori_n895_));
  NO2        o873(.A(ori_ori_n228_), .B(ori_ori_n95_), .Y(ori_ori_n896_));
  NA2        o874(.A(ori_ori_n896_), .B(ori_ori_n880_), .Y(ori_ori_n897_));
  OR2        o875(.A(ori_ori_n897_), .B(i_5_), .Y(ori_ori_n898_));
  AOI210     o876(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n175_), .Y(ori_ori_n899_));
  NA2        o877(.A(ori_ori_n899_), .B(ori_ori_n864_), .Y(ori_ori_n900_));
  INV        o878(.A(ori_ori_n491_), .Y(ori_ori_n901_));
  NO3        o879(.A(ori_ori_n795_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n902_));
  NA2        o880(.A(ori_ori_n448_), .B(ori_ori_n441_), .Y(ori_ori_n903_));
  NO3        o881(.A(ori_ori_n903_), .B(ori_ori_n902_), .C(ori_ori_n901_), .Y(ori_ori_n904_));
  NA3        o882(.A(ori_ori_n358_), .B(ori_ori_n172_), .C(ori_ori_n171_), .Y(ori_ori_n905_));
  INV        o883(.A(ori_ori_n905_), .Y(ori_ori_n906_));
  NA3        o884(.A(ori_ori_n358_), .B(ori_ori_n312_), .C(ori_ori_n211_), .Y(ori_ori_n907_));
  INV        o885(.A(ori_ori_n907_), .Y(ori_ori_n908_));
  NOi31      o886(.An(ori_ori_n357_), .B(ori_ori_n881_), .C(ori_ori_n226_), .Y(ori_ori_n909_));
  NO3        o887(.A(ori_ori_n840_), .B(ori_ori_n209_), .C(ori_ori_n187_), .Y(ori_ori_n910_));
  NO4        o888(.A(ori_ori_n910_), .B(ori_ori_n909_), .C(ori_ori_n908_), .D(ori_ori_n906_), .Y(ori_ori_n911_));
  NA4        o889(.A(ori_ori_n911_), .B(ori_ori_n904_), .C(ori_ori_n900_), .D(ori_ori_n898_), .Y(ori_ori_n912_));
  NO2        o890(.A(ori_ori_n86_), .B(i_5_), .Y(ori_ori_n913_));
  NA3        o891(.A(ori_ori_n790_), .B(ori_ori_n112_), .C(ori_ori_n127_), .Y(ori_ori_n914_));
  INV        o892(.A(ori_ori_n914_), .Y(ori_ori_n915_));
  NA2        o893(.A(ori_ori_n915_), .B(ori_ori_n913_), .Y(ori_ori_n916_));
  NA3        o894(.A(ori_ori_n286_), .B(i_5_), .C(ori_ori_n189_), .Y(ori_ori_n917_));
  NAi31      o895(.An(ori_ori_n227_), .B(ori_ori_n917_), .C(ori_ori_n228_), .Y(ori_ori_n918_));
  NO4        o896(.A(ori_ori_n226_), .B(ori_ori_n202_), .C(i_0_), .D(i_12_), .Y(ori_ori_n919_));
  NA2        o897(.A(ori_ori_n919_), .B(ori_ori_n918_), .Y(ori_ori_n920_));
  AN2        o898(.A(ori_ori_n831_), .B(ori_ori_n155_), .Y(ori_ori_n921_));
  NO4        o899(.A(ori_ori_n921_), .B(i_12_), .C(ori_ori_n596_), .D(ori_ori_n134_), .Y(ori_ori_n922_));
  NA2        o900(.A(ori_ori_n922_), .B(ori_ori_n209_), .Y(ori_ori_n923_));
  NA3        o901(.A(ori_ori_n101_), .B(ori_ori_n516_), .C(i_11_), .Y(ori_ori_n924_));
  NO2        o902(.A(ori_ori_n924_), .B(ori_ori_n157_), .Y(ori_ori_n925_));
  NA2        o903(.A(ori_ori_n859_), .B(ori_ori_n433_), .Y(ori_ori_n926_));
  NA2        o904(.A(ori_ori_n64_), .B(ori_ori_n104_), .Y(ori_ori_n927_));
  OAI220     o905(.A0(ori_ori_n927_), .A1(ori_ori_n917_), .B0(ori_ori_n926_), .B1(ori_ori_n626_), .Y(ori_ori_n928_));
  AOI210     o906(.A0(ori_ori_n928_), .A1(ori_ori_n847_), .B0(ori_ori_n925_), .Y(ori_ori_n929_));
  NA4        o907(.A(ori_ori_n929_), .B(ori_ori_n923_), .C(ori_ori_n920_), .D(ori_ori_n916_), .Y(ori_ori_n930_));
  NO4        o908(.A(ori_ori_n930_), .B(ori_ori_n912_), .C(ori_ori_n895_), .D(ori_ori_n890_), .Y(ori_ori_n931_));
  OAI210     o909(.A0(ori_ori_n765_), .A1(ori_ori_n758_), .B0(ori_ori_n37_), .Y(ori_ori_n932_));
  NA3        o910(.A(ori_ori_n853_), .B(ori_ori_n335_), .C(i_5_), .Y(ori_ori_n933_));
  NA3        o911(.A(ori_ori_n933_), .B(ori_ori_n932_), .C(ori_ori_n559_), .Y(ori_ori_n934_));
  NA2        o912(.A(ori_ori_n934_), .B(ori_ori_n200_), .Y(ori_ori_n935_));
  AN2        o913(.A(ori_ori_n646_), .B(ori_ori_n336_), .Y(ori_ori_n936_));
  NA2        o914(.A(ori_ori_n184_), .B(ori_ori_n186_), .Y(ori_ori_n937_));
  AO210      o915(.A0(ori_ori_n936_), .A1(ori_ori_n33_), .B0(ori_ori_n937_), .Y(ori_ori_n938_));
  NAi31      o916(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n939_));
  AOI210     o917(.A0(ori_ori_n120_), .A1(ori_ori_n70_), .B0(ori_ori_n939_), .Y(ori_ori_n940_));
  NO2        o918(.A(ori_ori_n940_), .B(ori_ori_n593_), .Y(ori_ori_n941_));
  NA2        o919(.A(ori_ori_n941_), .B(ori_ori_n938_), .Y(ori_ori_n942_));
  NO2        o920(.A(ori_ori_n427_), .B(ori_ori_n249_), .Y(ori_ori_n943_));
  NO2        o921(.A(ori_ori_n943_), .B(ori_ori_n823_), .Y(ori_ori_n944_));
  OAI210     o922(.A0(ori_ori_n924_), .A1(ori_ori_n151_), .B0(ori_ori_n944_), .Y(ori_ori_n945_));
  AOI210     o923(.A0(ori_ori_n942_), .A1(ori_ori_n48_), .B0(ori_ori_n945_), .Y(ori_ori_n946_));
  AOI210     o924(.A0(ori_ori_n946_), .A1(ori_ori_n935_), .B0(ori_ori_n73_), .Y(ori_ori_n947_));
  INV        o925(.A(ori_ori_n347_), .Y(ori_ori_n948_));
  NO2        o926(.A(ori_ori_n948_), .B(ori_ori_n705_), .Y(ori_ori_n949_));
  OAI210     o927(.A0(ori_ori_n80_), .A1(ori_ori_n54_), .B0(ori_ori_n111_), .Y(ori_ori_n950_));
  NA2        o928(.A(ori_ori_n950_), .B(ori_ori_n76_), .Y(ori_ori_n951_));
  NA2        o929(.A(ori_ori_n899_), .B(ori_ori_n843_), .Y(ori_ori_n952_));
  AOI210     o930(.A0(ori_ori_n952_), .A1(ori_ori_n951_), .B0(ori_ori_n629_), .Y(ori_ori_n953_));
  INV        o931(.A(ori_ori_n953_), .Y(ori_ori_n954_));
  OAI210     o932(.A0(ori_ori_n251_), .A1(ori_ori_n159_), .B0(ori_ori_n89_), .Y(ori_ori_n955_));
  NO2        o933(.A(ori_ori_n955_), .B(i_11_), .Y(ori_ori_n956_));
  NA2        o934(.A(ori_ori_n554_), .B(ori_ori_n207_), .Y(ori_ori_n957_));
  OAI210     o935(.A0(ori_ori_n957_), .A1(ori_ori_n853_), .B0(ori_ori_n200_), .Y(ori_ori_n958_));
  NA2        o936(.A(ori_ori_n165_), .B(i_5_), .Y(ori_ori_n959_));
  NO2        o937(.A(ori_ori_n958_), .B(ori_ori_n959_), .Y(ori_ori_n960_));
  NO3        o938(.A(ori_ori_n59_), .B(ori_ori_n58_), .C(i_4_), .Y(ori_ori_n961_));
  OAI210     o939(.A0(ori_ori_n861_), .A1(ori_ori_n287_), .B0(ori_ori_n961_), .Y(ori_ori_n962_));
  NO2        o940(.A(ori_ori_n962_), .B(ori_ori_n676_), .Y(ori_ori_n963_));
  INV        o941(.A(ori_ori_n509_), .Y(ori_ori_n964_));
  INV        o942(.A(ori_ori_n328_), .Y(ori_ori_n965_));
  AOI210     o943(.A0(ori_ori_n965_), .A1(ori_ori_n964_), .B0(ori_ori_n41_), .Y(ori_ori_n966_));
  NO4        o944(.A(ori_ori_n966_), .B(ori_ori_n963_), .C(ori_ori_n960_), .D(ori_ori_n956_), .Y(ori_ori_n967_));
  OAI210     o945(.A0(ori_ori_n954_), .A1(i_4_), .B0(ori_ori_n967_), .Y(ori_ori_n968_));
  NO3        o946(.A(ori_ori_n968_), .B(ori_ori_n949_), .C(ori_ori_n947_), .Y(ori_ori_n969_));
  NA4        o947(.A(ori_ori_n969_), .B(ori_ori_n931_), .C(ori_ori_n879_), .D(ori_ori_n813_), .Y(ori4));
  INV        o948(.A(ori_ori_n650_), .Y(ori_ori_n973_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m0033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m0034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m0036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m0037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m0038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m0039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m0040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m0041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m0042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m0043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m0044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m0045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m0046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m0047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m0049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m0050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m0051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m0052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m0053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m0054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m0055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m0057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m0059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m0060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m0062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m0063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m0064(.A(i_6_), .Y(mai_mai_n87_));
  OR4        m0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n88_));
  INV        m0066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m0067(.A(i_2_), .B(i_7_), .Y(mai_mai_n90_));
  NO2        m0068(.A(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  OAI210     m0069(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NAi21      m0070(.An(i_6_), .B(i_10_), .Y(mai_mai_n93_));
  NA2        m0071(.A(i_6_), .B(i_9_), .Y(mai_mai_n94_));
  AOI210     m0072(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n64_), .Y(mai_mai_n95_));
  NA2        m0073(.A(i_2_), .B(i_6_), .Y(mai_mai_n96_));
  NO3        m0074(.A(mai_mai_n96_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n97_));
  NO2        m0075(.A(mai_mai_n97_), .B(mai_mai_n95_), .Y(mai_mai_n98_));
  AOI210     m0076(.A0(mai_mai_n98_), .A1(mai_mai_n92_), .B0(mai_mai_n81_), .Y(mai_mai_n99_));
  AN3        m0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n100_));
  NAi21      m0078(.An(i_6_), .B(i_11_), .Y(mai_mai_n101_));
  NO2        m0079(.A(i_5_), .B(i_8_), .Y(mai_mai_n102_));
  NOi21      m0080(.An(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  AOI220     m0081(.A0(mai_mai_n103_), .A1(mai_mai_n63_), .B0(mai_mai_n100_), .B1(mai_mai_n32_), .Y(mai_mai_n104_));
  INV        m0082(.A(i_7_), .Y(mai_mai_n105_));
  NA2        m0083(.A(mai_mai_n47_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  NO2        m0084(.A(i_0_), .B(i_5_), .Y(mai_mai_n107_));
  NO2        m0085(.A(mai_mai_n107_), .B(mai_mai_n87_), .Y(mai_mai_n108_));
  NA2        m0086(.A(i_12_), .B(i_3_), .Y(mai_mai_n109_));
  INV        m0087(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NA3        m0088(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n106_), .Y(mai_mai_n111_));
  NAi21      m0089(.An(i_7_), .B(i_11_), .Y(mai_mai_n112_));
  NO3        m0090(.A(mai_mai_n112_), .B(mai_mai_n93_), .C(mai_mai_n54_), .Y(mai_mai_n113_));
  AN2        m0091(.A(i_2_), .B(i_10_), .Y(mai_mai_n114_));
  NO2        m0092(.A(mai_mai_n114_), .B(i_7_), .Y(mai_mai_n115_));
  OR2        m0093(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n116_));
  NO2        m0094(.A(i_8_), .B(mai_mai_n105_), .Y(mai_mai_n117_));
  NO3        m0095(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(mai_mai_n115_), .Y(mai_mai_n118_));
  NA2        m0096(.A(i_12_), .B(i_7_), .Y(mai_mai_n119_));
  NO2        m0097(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n120_));
  NA2        m0098(.A(mai_mai_n120_), .B(i_0_), .Y(mai_mai_n121_));
  NA2        m0099(.A(i_11_), .B(i_12_), .Y(mai_mai_n122_));
  OAI210     m0100(.A0(mai_mai_n121_), .A1(mai_mai_n119_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NO2        m0101(.A(mai_mai_n123_), .B(mai_mai_n118_), .Y(mai_mai_n124_));
  NAi41      m0102(.An(mai_mai_n113_), .B(mai_mai_n124_), .C(mai_mai_n111_), .D(mai_mai_n104_), .Y(mai_mai_n125_));
  NOi21      m0103(.An(i_1_), .B(i_5_), .Y(mai_mai_n126_));
  NA2        m0104(.A(mai_mai_n126_), .B(i_11_), .Y(mai_mai_n127_));
  NA2        m0105(.A(mai_mai_n105_), .B(mai_mai_n37_), .Y(mai_mai_n128_));
  NA2        m0106(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n129_));
  NA2        m0107(.A(mai_mai_n129_), .B(mai_mai_n128_), .Y(mai_mai_n130_));
  NO2        m0108(.A(mai_mai_n130_), .B(mai_mai_n47_), .Y(mai_mai_n131_));
  NA2        m0109(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n132_));
  NAi21      m0110(.An(i_3_), .B(i_8_), .Y(mai_mai_n133_));
  NA2        m0111(.A(mai_mai_n133_), .B(mai_mai_n63_), .Y(mai_mai_n134_));
  NOi31      m0112(.An(mai_mai_n134_), .B(mai_mai_n132_), .C(mai_mai_n131_), .Y(mai_mai_n135_));
  NO2        m0113(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n136_));
  NO2        m0114(.A(i_6_), .B(i_5_), .Y(mai_mai_n137_));
  NA2        m0115(.A(mai_mai_n137_), .B(i_3_), .Y(mai_mai_n138_));
  AO210      m0116(.A0(mai_mai_n138_), .A1(mai_mai_n48_), .B0(mai_mai_n136_), .Y(mai_mai_n139_));
  OAI220     m0117(.A0(mai_mai_n139_), .A1(mai_mai_n112_), .B0(mai_mai_n135_), .B1(mai_mai_n127_), .Y(mai_mai_n140_));
  NO3        m0118(.A(mai_mai_n140_), .B(mai_mai_n125_), .C(mai_mai_n99_), .Y(mai_mai_n141_));
  NA3        m0119(.A(mai_mai_n141_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m0120(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n143_));
  NA2        m0121(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n144_));
  NA2        m0122(.A(mai_mai_n144_), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  NA4        m0123(.A(mai_mai_n145_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0124(.A(i_8_), .B(i_7_), .Y(mai_mai_n147_));
  NA2        m0125(.A(mai_mai_n147_), .B(i_6_), .Y(mai_mai_n148_));
  NO2        m0126(.A(i_12_), .B(i_13_), .Y(mai_mai_n149_));
  NAi21      m0127(.An(i_5_), .B(i_11_), .Y(mai_mai_n150_));
  NOi21      m0128(.An(mai_mai_n149_), .B(mai_mai_n150_), .Y(mai_mai_n151_));
  NO2        m0129(.A(i_0_), .B(i_1_), .Y(mai_mai_n152_));
  NA2        m0130(.A(i_2_), .B(i_3_), .Y(mai_mai_n153_));
  NO2        m0131(.A(mai_mai_n153_), .B(i_4_), .Y(mai_mai_n154_));
  NA3        m0132(.A(mai_mai_n154_), .B(mai_mai_n152_), .C(mai_mai_n151_), .Y(mai_mai_n155_));
  OR2        m0133(.A(mai_mai_n155_), .B(mai_mai_n25_), .Y(mai_mai_n156_));
  AN2        m0134(.A(mai_mai_n149_), .B(mai_mai_n84_), .Y(mai_mai_n157_));
  NO2        m0135(.A(mai_mai_n157_), .B(mai_mai_n27_), .Y(mai_mai_n158_));
  NA2        m0136(.A(i_1_), .B(i_5_), .Y(mai_mai_n159_));
  NO2        m0137(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n160_));
  NA2        m0138(.A(mai_mai_n160_), .B(mai_mai_n36_), .Y(mai_mai_n161_));
  NO3        m0139(.A(mai_mai_n161_), .B(mai_mai_n159_), .C(mai_mai_n158_), .Y(mai_mai_n162_));
  OR2        m0140(.A(i_0_), .B(i_1_), .Y(mai_mai_n163_));
  NO3        m0141(.A(mai_mai_n163_), .B(mai_mai_n81_), .C(i_13_), .Y(mai_mai_n164_));
  NAi32      m0142(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n165_));
  NAi21      m0143(.An(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  NOi21      m0144(.An(i_4_), .B(i_10_), .Y(mai_mai_n167_));
  NA2        m0145(.A(mai_mai_n167_), .B(mai_mai_n40_), .Y(mai_mai_n168_));
  NO2        m0146(.A(i_3_), .B(i_5_), .Y(mai_mai_n169_));
  INV        m0147(.A(mai_mai_n162_), .Y(mai_mai_n170_));
  AOI210     m0148(.A0(mai_mai_n170_), .A1(mai_mai_n156_), .B0(mai_mai_n148_), .Y(mai_mai_n171_));
  NA3        m0149(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n172_));
  NA2        m0150(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n173_));
  NOi21      m0151(.An(i_4_), .B(i_9_), .Y(mai_mai_n174_));
  NOi21      m0152(.An(i_11_), .B(i_13_), .Y(mai_mai_n175_));
  NA2        m0153(.A(mai_mai_n175_), .B(mai_mai_n174_), .Y(mai_mai_n176_));
  OR2        m0154(.A(mai_mai_n176_), .B(mai_mai_n173_), .Y(mai_mai_n177_));
  NO2        m0155(.A(i_4_), .B(i_5_), .Y(mai_mai_n178_));
  NAi21      m0156(.An(i_12_), .B(i_11_), .Y(mai_mai_n179_));
  NO2        m0157(.A(mai_mai_n179_), .B(i_13_), .Y(mai_mai_n180_));
  NA3        m0158(.A(mai_mai_n180_), .B(mai_mai_n178_), .C(mai_mai_n84_), .Y(mai_mai_n181_));
  AOI210     m0159(.A0(mai_mai_n181_), .A1(mai_mai_n177_), .B0(mai_mai_n172_), .Y(mai_mai_n182_));
  NO2        m0160(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n183_));
  NA2        m0161(.A(mai_mai_n183_), .B(mai_mai_n47_), .Y(mai_mai_n184_));
  NA2        m0162(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n185_));
  NA2        m0163(.A(i_3_), .B(i_5_), .Y(mai_mai_n186_));
  NO2        m0164(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n187_));
  NO2        m0165(.A(i_13_), .B(i_10_), .Y(mai_mai_n188_));
  NA3        m0166(.A(mai_mai_n188_), .B(mai_mai_n187_), .C(mai_mai_n45_), .Y(mai_mai_n189_));
  NO2        m0167(.A(i_2_), .B(i_1_), .Y(mai_mai_n190_));
  NA2        m0168(.A(mai_mai_n190_), .B(i_3_), .Y(mai_mai_n191_));
  NAi21      m0169(.An(i_4_), .B(i_12_), .Y(mai_mai_n192_));
  NO4        m0170(.A(mai_mai_n192_), .B(mai_mai_n191_), .C(mai_mai_n189_), .D(mai_mai_n25_), .Y(mai_mai_n193_));
  NO2        m0171(.A(mai_mai_n193_), .B(mai_mai_n182_), .Y(mai_mai_n194_));
  INV        m0172(.A(i_8_), .Y(mai_mai_n195_));
  NO2        m0173(.A(mai_mai_n195_), .B(i_7_), .Y(mai_mai_n196_));
  NA2        m0174(.A(mai_mai_n196_), .B(i_6_), .Y(mai_mai_n197_));
  NO3        m0175(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n198_));
  NA2        m0176(.A(mai_mai_n198_), .B(mai_mai_n117_), .Y(mai_mai_n199_));
  NO3        m0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n200_));
  NA3        m0178(.A(mai_mai_n200_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n201_));
  NO3        m0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n202_));
  OAI210     m0180(.A0(mai_mai_n100_), .A1(i_12_), .B0(mai_mai_n202_), .Y(mai_mai_n203_));
  AOI210     m0181(.A0(mai_mai_n203_), .A1(mai_mai_n201_), .B0(mai_mai_n199_), .Y(mai_mai_n204_));
  NO2        m0182(.A(i_3_), .B(i_8_), .Y(mai_mai_n205_));
  NO3        m0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n206_));
  NA3        m0184(.A(mai_mai_n206_), .B(mai_mai_n205_), .C(mai_mai_n40_), .Y(mai_mai_n207_));
  NO2        m0185(.A(mai_mai_n107_), .B(mai_mai_n59_), .Y(mai_mai_n208_));
  INV        m0186(.A(mai_mai_n208_), .Y(mai_mai_n209_));
  NO2        m0187(.A(i_13_), .B(i_9_), .Y(mai_mai_n210_));
  NA3        m0188(.A(mai_mai_n210_), .B(i_6_), .C(mai_mai_n195_), .Y(mai_mai_n211_));
  NAi21      m0189(.An(i_12_), .B(i_3_), .Y(mai_mai_n212_));
  OR2        m0190(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n213_));
  NO2        m0191(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n214_));
  NO3        m0192(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n215_));
  NA3        m0193(.A(mai_mai_n215_), .B(mai_mai_n214_), .C(i_10_), .Y(mai_mai_n216_));
  OAI220     m0194(.A0(mai_mai_n216_), .A1(mai_mai_n213_), .B0(mai_mai_n209_), .B1(mai_mai_n207_), .Y(mai_mai_n217_));
  AOI210     m0195(.A0(mai_mai_n217_), .A1(i_7_), .B0(mai_mai_n204_), .Y(mai_mai_n218_));
  OAI220     m0196(.A0(mai_mai_n218_), .A1(i_4_), .B0(mai_mai_n197_), .B1(mai_mai_n194_), .Y(mai_mai_n219_));
  NAi21      m0197(.An(i_12_), .B(i_7_), .Y(mai_mai_n220_));
  NA3        m0198(.A(i_13_), .B(mai_mai_n195_), .C(i_10_), .Y(mai_mai_n221_));
  NO2        m0199(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  NA2        m0200(.A(i_0_), .B(i_5_), .Y(mai_mai_n223_));
  NA2        m0201(.A(mai_mai_n223_), .B(mai_mai_n108_), .Y(mai_mai_n224_));
  OAI220     m0202(.A0(mai_mai_n224_), .A1(mai_mai_n191_), .B0(mai_mai_n184_), .B1(mai_mai_n138_), .Y(mai_mai_n225_));
  NAi31      m0203(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n226_));
  NO2        m0204(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n227_));
  NO2        m0205(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n228_));
  NO2        m0206(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n229_));
  INV        m0207(.A(i_13_), .Y(mai_mai_n230_));
  NO2        m0208(.A(i_12_), .B(mai_mai_n230_), .Y(mai_mai_n231_));
  NA2        m0209(.A(mai_mai_n225_), .B(mai_mai_n222_), .Y(mai_mai_n232_));
  NO2        m0210(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n233_));
  NO2        m0211(.A(mai_mai_n186_), .B(i_4_), .Y(mai_mai_n234_));
  NA2        m0212(.A(mai_mai_n234_), .B(mai_mai_n233_), .Y(mai_mai_n235_));
  OR2        m0213(.A(i_8_), .B(i_7_), .Y(mai_mai_n236_));
  NO2        m0214(.A(mai_mai_n236_), .B(mai_mai_n87_), .Y(mai_mai_n237_));
  NO2        m0215(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n238_));
  NA2        m0216(.A(mai_mai_n238_), .B(mai_mai_n237_), .Y(mai_mai_n239_));
  INV        m0217(.A(i_12_), .Y(mai_mai_n240_));
  NO2        m0218(.A(mai_mai_n45_), .B(mai_mai_n240_), .Y(mai_mai_n241_));
  NO3        m0219(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n242_));
  NA2        m0220(.A(i_2_), .B(i_1_), .Y(mai_mai_n243_));
  NO2        m0221(.A(mai_mai_n239_), .B(mai_mai_n235_), .Y(mai_mai_n244_));
  NO3        m0222(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n245_));
  NAi21      m0223(.An(i_4_), .B(i_3_), .Y(mai_mai_n246_));
  NO2        m0224(.A(i_0_), .B(i_6_), .Y(mai_mai_n247_));
  NOi41      m0225(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n248_));
  NA2        m0226(.A(mai_mai_n248_), .B(mai_mai_n247_), .Y(mai_mai_n249_));
  NO2        m0227(.A(mai_mai_n243_), .B(mai_mai_n186_), .Y(mai_mai_n250_));
  NAi21      m0228(.An(mai_mai_n249_), .B(mai_mai_n250_), .Y(mai_mai_n251_));
  INV        m0229(.A(mai_mai_n251_), .Y(mai_mai_n252_));
  AOI220     m0230(.A0(mai_mai_n252_), .A1(mai_mai_n40_), .B0(mai_mai_n244_), .B1(mai_mai_n210_), .Y(mai_mai_n253_));
  NO2        m0231(.A(i_11_), .B(mai_mai_n230_), .Y(mai_mai_n254_));
  NOi21      m0232(.An(i_1_), .B(i_6_), .Y(mai_mai_n255_));
  NAi21      m0233(.An(i_3_), .B(i_7_), .Y(mai_mai_n256_));
  NA2        m0234(.A(mai_mai_n240_), .B(i_9_), .Y(mai_mai_n257_));
  OR4        m0235(.A(mai_mai_n257_), .B(mai_mai_n256_), .C(mai_mai_n255_), .D(mai_mai_n187_), .Y(mai_mai_n258_));
  NO2        m0236(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n259_));
  NO2        m0237(.A(i_12_), .B(i_3_), .Y(mai_mai_n260_));
  NA2        m0238(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n261_));
  NA2        m0239(.A(i_3_), .B(i_9_), .Y(mai_mai_n262_));
  NAi21      m0240(.An(i_7_), .B(i_10_), .Y(mai_mai_n263_));
  NO2        m0241(.A(mai_mai_n263_), .B(mai_mai_n262_), .Y(mai_mai_n264_));
  NA3        m0242(.A(mai_mai_n264_), .B(mai_mai_n261_), .C(mai_mai_n65_), .Y(mai_mai_n265_));
  NA2        m0243(.A(mai_mai_n265_), .B(mai_mai_n258_), .Y(mai_mai_n266_));
  NA3        m0244(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n267_));
  INV        m0245(.A(mai_mai_n148_), .Y(mai_mai_n268_));
  NA2        m0246(.A(mai_mai_n240_), .B(i_13_), .Y(mai_mai_n269_));
  NO2        m0247(.A(mai_mai_n269_), .B(mai_mai_n76_), .Y(mai_mai_n270_));
  AOI220     m0248(.A0(mai_mai_n270_), .A1(mai_mai_n268_), .B0(mai_mai_n266_), .B1(mai_mai_n254_), .Y(mai_mai_n271_));
  NO2        m0249(.A(mai_mai_n236_), .B(mai_mai_n37_), .Y(mai_mai_n272_));
  NA2        m0250(.A(i_12_), .B(i_6_), .Y(mai_mai_n273_));
  OR2        m0251(.A(i_13_), .B(i_9_), .Y(mai_mai_n274_));
  NO3        m0252(.A(mai_mai_n274_), .B(mai_mai_n273_), .C(mai_mai_n49_), .Y(mai_mai_n275_));
  NO2        m0253(.A(mai_mai_n246_), .B(i_2_), .Y(mai_mai_n276_));
  NA3        m0254(.A(mai_mai_n276_), .B(mai_mai_n275_), .C(mai_mai_n45_), .Y(mai_mai_n277_));
  NA2        m0255(.A(mai_mai_n254_), .B(i_9_), .Y(mai_mai_n278_));
  NA2        m0256(.A(mai_mai_n261_), .B(mai_mai_n65_), .Y(mai_mai_n279_));
  OAI210     m0257(.A0(mai_mai_n279_), .A1(mai_mai_n278_), .B0(mai_mai_n277_), .Y(mai_mai_n280_));
  NO3        m0258(.A(i_11_), .B(mai_mai_n230_), .C(mai_mai_n25_), .Y(mai_mai_n281_));
  NO2        m0259(.A(mai_mai_n256_), .B(i_8_), .Y(mai_mai_n282_));
  NO2        m0260(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n283_));
  NA2        m0261(.A(mai_mai_n280_), .B(mai_mai_n272_), .Y(mai_mai_n284_));
  NA4        m0262(.A(mai_mai_n284_), .B(mai_mai_n271_), .C(mai_mai_n253_), .D(mai_mai_n232_), .Y(mai_mai_n285_));
  NO3        m0263(.A(i_12_), .B(mai_mai_n230_), .C(mai_mai_n37_), .Y(mai_mai_n286_));
  INV        m0264(.A(mai_mai_n286_), .Y(mai_mai_n287_));
  NO3        m0265(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n288_));
  NO2        m0266(.A(mai_mai_n243_), .B(i_0_), .Y(mai_mai_n289_));
  NA2        m0267(.A(i_0_), .B(i_1_), .Y(mai_mai_n290_));
  NO2        m0268(.A(mai_mai_n290_), .B(i_2_), .Y(mai_mai_n291_));
  NO2        m0269(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n292_));
  NA3        m0270(.A(mai_mai_n292_), .B(mai_mai_n291_), .C(mai_mai_n169_), .Y(mai_mai_n293_));
  NO2        m0271(.A(i_3_), .B(i_10_), .Y(mai_mai_n294_));
  NA3        m0272(.A(mai_mai_n294_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n295_));
  NO2        m0273(.A(i_2_), .B(mai_mai_n105_), .Y(mai_mai_n296_));
  NA2        m0274(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n297_));
  NO2        m0275(.A(mai_mai_n297_), .B(i_8_), .Y(mai_mai_n298_));
  NOi21      m0276(.An(mai_mai_n223_), .B(mai_mai_n107_), .Y(mai_mai_n299_));
  NA3        m0277(.A(mai_mai_n299_), .B(mai_mai_n298_), .C(mai_mai_n296_), .Y(mai_mai_n300_));
  AN2        m0278(.A(i_3_), .B(i_10_), .Y(mai_mai_n301_));
  NA4        m0279(.A(mai_mai_n301_), .B(mai_mai_n200_), .C(mai_mai_n180_), .D(mai_mai_n178_), .Y(mai_mai_n302_));
  NO2        m0280(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n303_));
  NO2        m0281(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n304_));
  OR2        m0282(.A(mai_mai_n300_), .B(mai_mai_n295_), .Y(mai_mai_n305_));
  OAI220     m0283(.A0(mai_mai_n305_), .A1(i_6_), .B0(mai_mai_n293_), .B1(mai_mai_n287_), .Y(mai_mai_n306_));
  NO4        m0284(.A(mai_mai_n306_), .B(mai_mai_n285_), .C(mai_mai_n219_), .D(mai_mai_n171_), .Y(mai_mai_n307_));
  NO3        m0285(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n308_));
  NO2        m0286(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n309_));
  NO3        m0287(.A(i_6_), .B(mai_mai_n195_), .C(i_7_), .Y(mai_mai_n310_));
  NO2        m0288(.A(i_2_), .B(i_3_), .Y(mai_mai_n311_));
  OR2        m0289(.A(i_0_), .B(i_5_), .Y(mai_mai_n312_));
  NA2        m0290(.A(mai_mai_n223_), .B(mai_mai_n312_), .Y(mai_mai_n313_));
  NA4        m0291(.A(mai_mai_n313_), .B(mai_mai_n237_), .C(mai_mai_n311_), .D(i_1_), .Y(mai_mai_n314_));
  NAi21      m0292(.An(i_8_), .B(i_7_), .Y(mai_mai_n315_));
  NO2        m0293(.A(mai_mai_n315_), .B(i_6_), .Y(mai_mai_n316_));
  NO2        m0294(.A(mai_mai_n163_), .B(mai_mai_n47_), .Y(mai_mai_n317_));
  NA3        m0295(.A(mai_mai_n317_), .B(mai_mai_n316_), .C(mai_mai_n169_), .Y(mai_mai_n318_));
  NA2        m0296(.A(mai_mai_n318_), .B(mai_mai_n314_), .Y(mai_mai_n319_));
  NA2        m0297(.A(mai_mai_n319_), .B(i_4_), .Y(mai_mai_n320_));
  NO2        m0298(.A(i_12_), .B(i_10_), .Y(mai_mai_n321_));
  NOi21      m0299(.An(i_5_), .B(i_0_), .Y(mai_mai_n322_));
  NA4        m0300(.A(mai_mai_n85_), .B(mai_mai_n36_), .C(mai_mai_n87_), .D(i_8_), .Y(mai_mai_n323_));
  NO2        m0301(.A(i_6_), .B(i_8_), .Y(mai_mai_n324_));
  NOi21      m0302(.An(i_0_), .B(i_2_), .Y(mai_mai_n325_));
  AN2        m0303(.A(mai_mai_n325_), .B(mai_mai_n324_), .Y(mai_mai_n326_));
  NO2        m0304(.A(i_1_), .B(i_7_), .Y(mai_mai_n327_));
  AO220      m0305(.A0(mai_mai_n327_), .A1(mai_mai_n326_), .B0(mai_mai_n316_), .B1(mai_mai_n238_), .Y(mai_mai_n328_));
  NA3        m0306(.A(mai_mai_n328_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n329_));
  NA2        m0307(.A(mai_mai_n329_), .B(mai_mai_n320_), .Y(mai_mai_n330_));
  NO3        m0308(.A(mai_mai_n236_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n331_));
  NO3        m0309(.A(mai_mai_n315_), .B(i_2_), .C(i_1_), .Y(mai_mai_n332_));
  OAI210     m0310(.A0(mai_mai_n332_), .A1(mai_mai_n331_), .B0(i_6_), .Y(mai_mai_n333_));
  NA3        m0311(.A(mai_mai_n255_), .B(mai_mai_n296_), .C(mai_mai_n195_), .Y(mai_mai_n334_));
  AOI210     m0312(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n313_), .Y(mai_mai_n335_));
  NOi21      m0313(.An(mai_mai_n159_), .B(mai_mai_n108_), .Y(mai_mai_n336_));
  NO2        m0314(.A(mai_mai_n336_), .B(mai_mai_n129_), .Y(mai_mai_n337_));
  OAI210     m0315(.A0(mai_mai_n337_), .A1(mai_mai_n335_), .B0(i_3_), .Y(mai_mai_n338_));
  INV        m0316(.A(mai_mai_n85_), .Y(mai_mai_n339_));
  NO2        m0317(.A(mai_mai_n290_), .B(mai_mai_n82_), .Y(mai_mai_n340_));
  NA2        m0318(.A(mai_mai_n340_), .B(mai_mai_n137_), .Y(mai_mai_n341_));
  NO2        m0319(.A(mai_mai_n96_), .B(mai_mai_n195_), .Y(mai_mai_n342_));
  NA3        m0320(.A(mai_mai_n299_), .B(mai_mai_n342_), .C(mai_mai_n64_), .Y(mai_mai_n343_));
  AOI210     m0321(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(mai_mai_n339_), .Y(mai_mai_n344_));
  NO2        m0322(.A(mai_mai_n195_), .B(i_9_), .Y(mai_mai_n345_));
  NA2        m0323(.A(mai_mai_n345_), .B(mai_mai_n208_), .Y(mai_mai_n346_));
  NO2        m0324(.A(mai_mai_n346_), .B(mai_mai_n47_), .Y(mai_mai_n347_));
  NO2        m0325(.A(mai_mai_n347_), .B(mai_mai_n344_), .Y(mai_mai_n348_));
  AOI210     m0326(.A0(mai_mai_n348_), .A1(mai_mai_n338_), .B0(mai_mai_n168_), .Y(mai_mai_n349_));
  AOI210     m0327(.A0(mai_mai_n330_), .A1(mai_mai_n308_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NOi32      m0328(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n351_));
  INV        m0329(.A(mai_mai_n351_), .Y(mai_mai_n352_));
  NAi21      m0330(.An(i_0_), .B(i_6_), .Y(mai_mai_n353_));
  NAi21      m0331(.An(i_1_), .B(i_5_), .Y(mai_mai_n354_));
  NA2        m0332(.A(mai_mai_n354_), .B(mai_mai_n353_), .Y(mai_mai_n355_));
  NA2        m0333(.A(mai_mai_n355_), .B(mai_mai_n25_), .Y(mai_mai_n356_));
  OAI210     m0334(.A0(mai_mai_n356_), .A1(mai_mai_n165_), .B0(mai_mai_n249_), .Y(mai_mai_n357_));
  NAi41      m0335(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n358_));
  OAI220     m0336(.A0(mai_mai_n358_), .A1(mai_mai_n354_), .B0(mai_mai_n226_), .B1(mai_mai_n165_), .Y(mai_mai_n359_));
  AOI210     m0337(.A0(mai_mai_n358_), .A1(mai_mai_n165_), .B0(mai_mai_n163_), .Y(mai_mai_n360_));
  NOi32      m0338(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n361_));
  OR2        m0339(.A(mai_mai_n360_), .B(mai_mai_n359_), .Y(mai_mai_n362_));
  NO2        m0340(.A(i_1_), .B(mai_mai_n105_), .Y(mai_mai_n363_));
  NAi21      m0341(.An(i_3_), .B(i_4_), .Y(mai_mai_n364_));
  NO2        m0342(.A(mai_mai_n364_), .B(i_9_), .Y(mai_mai_n365_));
  AN2        m0343(.A(i_6_), .B(i_7_), .Y(mai_mai_n366_));
  OAI210     m0344(.A0(mai_mai_n366_), .A1(mai_mai_n363_), .B0(mai_mai_n365_), .Y(mai_mai_n367_));
  NA2        m0345(.A(i_2_), .B(i_7_), .Y(mai_mai_n368_));
  NO2        m0346(.A(mai_mai_n364_), .B(i_10_), .Y(mai_mai_n369_));
  NA3        m0347(.A(mai_mai_n369_), .B(mai_mai_n368_), .C(mai_mai_n247_), .Y(mai_mai_n370_));
  AOI210     m0348(.A0(mai_mai_n370_), .A1(mai_mai_n367_), .B0(mai_mai_n187_), .Y(mai_mai_n371_));
  AOI210     m0349(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n372_));
  OAI210     m0350(.A0(mai_mai_n372_), .A1(mai_mai_n190_), .B0(mai_mai_n369_), .Y(mai_mai_n373_));
  AOI220     m0351(.A0(mai_mai_n369_), .A1(mai_mai_n327_), .B0(mai_mai_n242_), .B1(mai_mai_n190_), .Y(mai_mai_n374_));
  AOI210     m0352(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(i_5_), .Y(mai_mai_n375_));
  NO4        m0353(.A(mai_mai_n375_), .B(mai_mai_n371_), .C(mai_mai_n362_), .D(mai_mai_n357_), .Y(mai_mai_n376_));
  NO2        m0354(.A(mai_mai_n376_), .B(mai_mai_n352_), .Y(mai_mai_n377_));
  AN2        m0355(.A(i_12_), .B(i_5_), .Y(mai_mai_n378_));
  NO2        m0356(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n379_));
  NA2        m0357(.A(mai_mai_n379_), .B(mai_mai_n378_), .Y(mai_mai_n380_));
  NO2        m0358(.A(i_11_), .B(i_6_), .Y(mai_mai_n381_));
  NO2        m0359(.A(mai_mai_n246_), .B(i_5_), .Y(mai_mai_n382_));
  NO2        m0360(.A(i_5_), .B(i_10_), .Y(mai_mai_n383_));
  NO2        m0361(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n384_));
  NO3        m0362(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n385_));
  NO2        m0363(.A(i_3_), .B(mai_mai_n105_), .Y(mai_mai_n386_));
  NA4        m0364(.A(mai_mai_n294_), .B(mai_mai_n94_), .C(mai_mai_n76_), .D(mai_mai_n55_), .Y(mai_mai_n387_));
  NO2        m0365(.A(i_11_), .B(i_12_), .Y(mai_mai_n388_));
  NA2        m0366(.A(mai_mai_n388_), .B(mai_mai_n36_), .Y(mai_mai_n389_));
  NO2        m0367(.A(mai_mai_n387_), .B(mai_mai_n389_), .Y(mai_mai_n390_));
  NA3        m0368(.A(mai_mai_n117_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n391_));
  NO2        m0369(.A(mai_mai_n391_), .B(mai_mai_n226_), .Y(mai_mai_n392_));
  NAi21      m0370(.An(i_13_), .B(i_0_), .Y(mai_mai_n393_));
  NO2        m0371(.A(mai_mai_n393_), .B(mai_mai_n243_), .Y(mai_mai_n394_));
  OAI210     m0372(.A0(mai_mai_n392_), .A1(mai_mai_n390_), .B0(mai_mai_n394_), .Y(mai_mai_n395_));
  INV        m0373(.A(mai_mai_n395_), .Y(mai_mai_n396_));
  NA2        m0374(.A(mai_mai_n45_), .B(mai_mai_n230_), .Y(mai_mai_n397_));
  NO3        m0375(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n398_));
  NO2        m0376(.A(i_0_), .B(i_11_), .Y(mai_mai_n399_));
  INV        m0377(.A(i_5_), .Y(mai_mai_n400_));
  AN2        m0378(.A(i_1_), .B(i_6_), .Y(mai_mai_n401_));
  NOi21      m0379(.An(i_2_), .B(i_12_), .Y(mai_mai_n402_));
  NA2        m0380(.A(mai_mai_n402_), .B(mai_mai_n401_), .Y(mai_mai_n403_));
  NO2        m0381(.A(mai_mai_n403_), .B(mai_mai_n400_), .Y(mai_mai_n404_));
  NA2        m0382(.A(mai_mai_n147_), .B(i_9_), .Y(mai_mai_n405_));
  NO2        m0383(.A(mai_mai_n405_), .B(i_4_), .Y(mai_mai_n406_));
  NA2        m0384(.A(mai_mai_n404_), .B(mai_mai_n406_), .Y(mai_mai_n407_));
  NAi21      m0385(.An(i_9_), .B(i_4_), .Y(mai_mai_n408_));
  OR2        m0386(.A(i_13_), .B(i_10_), .Y(mai_mai_n409_));
  NO3        m0387(.A(mai_mai_n409_), .B(mai_mai_n122_), .C(mai_mai_n408_), .Y(mai_mai_n410_));
  NO2        m0388(.A(mai_mai_n176_), .B(mai_mai_n128_), .Y(mai_mai_n411_));
  OR2        m0389(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n412_));
  NO2        m0390(.A(mai_mai_n105_), .B(mai_mai_n25_), .Y(mai_mai_n413_));
  NA2        m0391(.A(mai_mai_n286_), .B(mai_mai_n413_), .Y(mai_mai_n414_));
  NA2        m0392(.A(mai_mai_n283_), .B(mai_mai_n215_), .Y(mai_mai_n415_));
  OAI220     m0393(.A0(mai_mai_n415_), .A1(mai_mai_n412_), .B0(mai_mai_n414_), .B1(mai_mai_n336_), .Y(mai_mai_n416_));
  INV        m0394(.A(mai_mai_n416_), .Y(mai_mai_n417_));
  AOI210     m0395(.A0(mai_mai_n417_), .A1(mai_mai_n407_), .B0(mai_mai_n26_), .Y(mai_mai_n418_));
  INV        m0396(.A(mai_mai_n314_), .Y(mai_mai_n419_));
  AOI220     m0397(.A0(mai_mai_n292_), .A1(mai_mai_n288_), .B0(mai_mai_n289_), .B1(mai_mai_n309_), .Y(mai_mai_n420_));
  NO2        m0398(.A(mai_mai_n420_), .B(mai_mai_n173_), .Y(mai_mai_n421_));
  NO2        m0399(.A(mai_mai_n186_), .B(mai_mai_n87_), .Y(mai_mai_n422_));
  NO2        m0400(.A(mai_mai_n421_), .B(mai_mai_n419_), .Y(mai_mai_n423_));
  NA2        m0401(.A(mai_mai_n195_), .B(i_10_), .Y(mai_mai_n424_));
  NA3        m0402(.A(mai_mai_n261_), .B(mai_mai_n65_), .C(i_2_), .Y(mai_mai_n425_));
  NO2        m0403(.A(mai_mai_n425_), .B(mai_mai_n424_), .Y(mai_mai_n426_));
  NA2        m0404(.A(mai_mai_n310_), .B(mai_mai_n313_), .Y(mai_mai_n427_));
  NO2        m0405(.A(mai_mai_n427_), .B(mai_mai_n191_), .Y(mai_mai_n428_));
  NO2        m0406(.A(mai_mai_n428_), .B(mai_mai_n426_), .Y(mai_mai_n429_));
  AOI210     m0407(.A0(mai_mai_n429_), .A1(mai_mai_n423_), .B0(mai_mai_n278_), .Y(mai_mai_n430_));
  NO4        m0408(.A(mai_mai_n430_), .B(mai_mai_n418_), .C(mai_mai_n396_), .D(mai_mai_n377_), .Y(mai_mai_n431_));
  NO2        m0409(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n432_));
  NO2        m0410(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n433_));
  NO2        m0411(.A(i_10_), .B(i_9_), .Y(mai_mai_n434_));
  NAi21      m0412(.An(i_12_), .B(i_8_), .Y(mai_mai_n435_));
  NO2        m0413(.A(mai_mai_n435_), .B(i_3_), .Y(mai_mai_n436_));
  NO2        m0414(.A(mai_mai_n47_), .B(i_4_), .Y(mai_mai_n437_));
  NA2        m0415(.A(mai_mai_n437_), .B(mai_mai_n108_), .Y(mai_mai_n438_));
  NO2        m0416(.A(mai_mai_n438_), .B(mai_mai_n207_), .Y(mai_mai_n439_));
  NA2        m0417(.A(mai_mai_n304_), .B(i_0_), .Y(mai_mai_n440_));
  NO3        m0418(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n441_));
  NA2        m0419(.A(mai_mai_n273_), .B(mai_mai_n101_), .Y(mai_mai_n442_));
  NA2        m0420(.A(mai_mai_n442_), .B(mai_mai_n441_), .Y(mai_mai_n443_));
  NA2        m0421(.A(i_8_), .B(i_9_), .Y(mai_mai_n444_));
  AOI210     m0422(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n445_));
  OR2        m0423(.A(mai_mai_n445_), .B(mai_mai_n444_), .Y(mai_mai_n446_));
  NA2        m0424(.A(mai_mai_n286_), .B(mai_mai_n208_), .Y(mai_mai_n447_));
  OAI220     m0425(.A0(mai_mai_n447_), .A1(mai_mai_n446_), .B0(mai_mai_n443_), .B1(mai_mai_n440_), .Y(mai_mai_n448_));
  NA2        m0426(.A(mai_mai_n254_), .B(mai_mai_n303_), .Y(mai_mai_n449_));
  NO3        m0427(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n450_));
  INV        m0428(.A(mai_mai_n450_), .Y(mai_mai_n451_));
  NA3        m0429(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n452_));
  NA4        m0430(.A(mai_mai_n150_), .B(mai_mai_n120_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n453_));
  OAI220     m0431(.A0(mai_mai_n453_), .A1(mai_mai_n452_), .B0(mai_mai_n451_), .B1(mai_mai_n449_), .Y(mai_mai_n454_));
  NO3        m0432(.A(mai_mai_n454_), .B(mai_mai_n448_), .C(mai_mai_n439_), .Y(mai_mai_n455_));
  NA2        m0433(.A(mai_mai_n291_), .B(mai_mai_n112_), .Y(mai_mai_n456_));
  OR2        m0434(.A(mai_mai_n456_), .B(mai_mai_n211_), .Y(mai_mai_n457_));
  OA210      m0435(.A0(mai_mai_n346_), .A1(mai_mai_n105_), .B0(mai_mai_n293_), .Y(mai_mai_n458_));
  OA220      m0436(.A0(mai_mai_n458_), .A1(mai_mai_n168_), .B0(mai_mai_n457_), .B1(mai_mai_n235_), .Y(mai_mai_n459_));
  NA2        m0437(.A(mai_mai_n100_), .B(i_13_), .Y(mai_mai_n460_));
  NO2        m0438(.A(i_2_), .B(i_13_), .Y(mai_mai_n461_));
  NA3        m0439(.A(mai_mai_n461_), .B(mai_mai_n167_), .C(mai_mai_n103_), .Y(mai_mai_n462_));
  NO2        m0440(.A(mai_mai_n462_), .B(mai_mai_n240_), .Y(mai_mai_n463_));
  NO3        m0441(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n464_));
  NO2        m0442(.A(i_6_), .B(i_7_), .Y(mai_mai_n465_));
  NA2        m0443(.A(mai_mai_n465_), .B(mai_mai_n464_), .Y(mai_mai_n466_));
  NO2        m0444(.A(i_11_), .B(i_1_), .Y(mai_mai_n467_));
  NO2        m0445(.A(mai_mai_n74_), .B(i_3_), .Y(mai_mai_n468_));
  OR2        m0446(.A(i_11_), .B(i_8_), .Y(mai_mai_n469_));
  NOi21      m0447(.An(i_2_), .B(i_7_), .Y(mai_mai_n470_));
  NAi31      m0448(.An(mai_mai_n469_), .B(mai_mai_n470_), .C(mai_mai_n468_), .Y(mai_mai_n471_));
  NO2        m0449(.A(mai_mai_n409_), .B(i_6_), .Y(mai_mai_n472_));
  NA3        m0450(.A(mai_mai_n472_), .B(mai_mai_n432_), .C(mai_mai_n76_), .Y(mai_mai_n473_));
  NO2        m0451(.A(mai_mai_n473_), .B(mai_mai_n471_), .Y(mai_mai_n474_));
  NO2        m0452(.A(i_3_), .B(mai_mai_n195_), .Y(mai_mai_n475_));
  NO2        m0453(.A(i_6_), .B(i_10_), .Y(mai_mai_n476_));
  NA4        m0454(.A(mai_mai_n476_), .B(mai_mai_n308_), .C(mai_mai_n475_), .D(mai_mai_n240_), .Y(mai_mai_n477_));
  NO2        m0455(.A(mai_mai_n477_), .B(mai_mai_n161_), .Y(mai_mai_n478_));
  NA3        m0456(.A(mai_mai_n248_), .B(mai_mai_n175_), .C(mai_mai_n137_), .Y(mai_mai_n479_));
  NA2        m0457(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n480_));
  NO2        m0458(.A(mai_mai_n163_), .B(i_3_), .Y(mai_mai_n481_));
  NAi31      m0459(.An(mai_mai_n480_), .B(mai_mai_n481_), .C(mai_mai_n231_), .Y(mai_mai_n482_));
  NA3        m0460(.A(mai_mai_n384_), .B(mai_mai_n183_), .C(mai_mai_n154_), .Y(mai_mai_n483_));
  NA3        m0461(.A(mai_mai_n483_), .B(mai_mai_n482_), .C(mai_mai_n479_), .Y(mai_mai_n484_));
  NO4        m0462(.A(mai_mai_n484_), .B(mai_mai_n478_), .C(mai_mai_n474_), .D(mai_mai_n463_), .Y(mai_mai_n485_));
  NA2        m0463(.A(mai_mai_n441_), .B(mai_mai_n378_), .Y(mai_mai_n486_));
  NA2        m0464(.A(mai_mai_n450_), .B(mai_mai_n383_), .Y(mai_mai_n487_));
  NAi21      m0465(.An(mai_mai_n221_), .B(mai_mai_n388_), .Y(mai_mai_n488_));
  NA2        m0466(.A(mai_mai_n327_), .B(mai_mai_n223_), .Y(mai_mai_n489_));
  NO2        m0467(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n490_));
  NO2        m0468(.A(mai_mai_n489_), .B(mai_mai_n488_), .Y(mai_mai_n491_));
  NA2        m0469(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n492_));
  NA2        m0470(.A(mai_mai_n308_), .B(mai_mai_n242_), .Y(mai_mai_n493_));
  OAI220     m0471(.A0(mai_mai_n493_), .A1(mai_mai_n425_), .B0(mai_mai_n492_), .B1(mai_mai_n460_), .Y(mai_mai_n494_));
  NA4        m0472(.A(mai_mai_n301_), .B(mai_mai_n229_), .C(mai_mai_n74_), .D(mai_mai_n240_), .Y(mai_mai_n495_));
  NO2        m0473(.A(mai_mai_n495_), .B(mai_mai_n466_), .Y(mai_mai_n496_));
  NO3        m0474(.A(mai_mai_n496_), .B(mai_mai_n494_), .C(mai_mai_n491_), .Y(mai_mai_n497_));
  NA4        m0475(.A(mai_mai_n497_), .B(mai_mai_n485_), .C(mai_mai_n459_), .D(mai_mai_n455_), .Y(mai_mai_n498_));
  NA3        m0476(.A(mai_mai_n301_), .B(mai_mai_n180_), .C(mai_mai_n178_), .Y(mai_mai_n499_));
  OAI210     m0477(.A0(mai_mai_n295_), .A1(mai_mai_n185_), .B0(mai_mai_n499_), .Y(mai_mai_n500_));
  AN2        m0478(.A(mai_mai_n288_), .B(mai_mai_n237_), .Y(mai_mai_n501_));
  NA2        m0479(.A(mai_mai_n501_), .B(mai_mai_n500_), .Y(mai_mai_n502_));
  NA2        m0480(.A(mai_mai_n127_), .B(mai_mai_n116_), .Y(mai_mai_n503_));
  AN2        m0481(.A(mai_mai_n503_), .B(mai_mai_n441_), .Y(mai_mai_n504_));
  NA2        m0482(.A(mai_mai_n308_), .B(i_0_), .Y(mai_mai_n505_));
  OAI210     m0483(.A0(mai_mai_n505_), .A1(mai_mai_n235_), .B0(mai_mai_n302_), .Y(mai_mai_n506_));
  AOI220     m0484(.A0(mai_mai_n506_), .A1(mai_mai_n316_), .B0(mai_mai_n504_), .B1(mai_mai_n304_), .Y(mai_mai_n507_));
  NA2        m0485(.A(mai_mai_n378_), .B(mai_mai_n230_), .Y(mai_mai_n508_));
  NA2        m0486(.A(mai_mai_n351_), .B(mai_mai_n74_), .Y(mai_mai_n509_));
  NA2        m0487(.A(mai_mai_n366_), .B(mai_mai_n361_), .Y(mai_mai_n510_));
  OR2        m0488(.A(mai_mai_n508_), .B(mai_mai_n510_), .Y(mai_mai_n511_));
  NO2        m0489(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n512_));
  AOI210     m0490(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n410_), .Y(mai_mai_n513_));
  NA2        m0491(.A(mai_mai_n513_), .B(mai_mai_n511_), .Y(mai_mai_n514_));
  INV        m0492(.A(mai_mai_n514_), .Y(mai_mai_n515_));
  INV        m0493(.A(mai_mai_n139_), .Y(mai_mai_n516_));
  NO2        m0494(.A(i_7_), .B(mai_mai_n201_), .Y(mai_mai_n517_));
  OR2        m0495(.A(mai_mai_n186_), .B(i_4_), .Y(mai_mai_n518_));
  NO2        m0496(.A(mai_mai_n518_), .B(mai_mai_n87_), .Y(mai_mai_n519_));
  AOI220     m0497(.A0(mai_mai_n519_), .A1(mai_mai_n517_), .B0(mai_mai_n516_), .B1(mai_mai_n411_), .Y(mai_mai_n520_));
  NA4        m0498(.A(mai_mai_n520_), .B(mai_mai_n515_), .C(mai_mai_n507_), .D(mai_mai_n502_), .Y(mai_mai_n521_));
  NA2        m0499(.A(mai_mai_n382_), .B(mai_mai_n291_), .Y(mai_mai_n522_));
  OAI210     m0500(.A0(mai_mai_n380_), .A1(mai_mai_n172_), .B0(mai_mai_n522_), .Y(mai_mai_n523_));
  NO2        m0501(.A(i_12_), .B(mai_mai_n195_), .Y(mai_mai_n524_));
  NA2        m0502(.A(mai_mai_n524_), .B(mai_mai_n230_), .Y(mai_mai_n525_));
  NO3        m0503(.A(mai_mai_n1049_), .B(mai_mai_n525_), .C(mai_mai_n456_), .Y(mai_mai_n526_));
  NOi31      m0504(.An(mai_mai_n310_), .B(mai_mai_n409_), .C(mai_mai_n38_), .Y(mai_mai_n527_));
  OAI210     m0505(.A0(mai_mai_n527_), .A1(mai_mai_n526_), .B0(mai_mai_n523_), .Y(mai_mai_n528_));
  NO2        m0506(.A(i_8_), .B(i_7_), .Y(mai_mai_n529_));
  AOI220     m0507(.A0(mai_mai_n317_), .A1(mai_mai_n40_), .B0(mai_mai_n238_), .B1(mai_mai_n210_), .Y(mai_mai_n530_));
  NO2        m0508(.A(mai_mai_n530_), .B(mai_mai_n518_), .Y(mai_mai_n531_));
  NA2        m0509(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n532_));
  NO2        m0510(.A(mai_mai_n532_), .B(i_6_), .Y(mai_mai_n533_));
  NA3        m0511(.A(mai_mai_n533_), .B(mai_mai_n531_), .C(mai_mai_n529_), .Y(mai_mai_n534_));
  AOI220     m0512(.A0(mai_mai_n422_), .A1(mai_mai_n317_), .B0(mai_mai_n250_), .B1(mai_mai_n247_), .Y(mai_mai_n535_));
  OAI220     m0513(.A0(mai_mai_n535_), .A1(mai_mai_n269_), .B0(mai_mai_n460_), .B1(mai_mai_n138_), .Y(mai_mai_n536_));
  NA2        m0514(.A(mai_mai_n536_), .B(mai_mai_n272_), .Y(mai_mai_n537_));
  NOi31      m0515(.An(mai_mai_n289_), .B(mai_mai_n295_), .C(mai_mai_n185_), .Y(mai_mai_n538_));
  NA3        m0516(.A(mai_mai_n301_), .B(mai_mai_n178_), .C(mai_mai_n100_), .Y(mai_mai_n539_));
  NO2        m0517(.A(mai_mai_n227_), .B(mai_mai_n45_), .Y(mai_mai_n540_));
  NO2        m0518(.A(mai_mai_n163_), .B(i_5_), .Y(mai_mai_n541_));
  NA3        m0519(.A(mai_mai_n541_), .B(mai_mai_n397_), .C(mai_mai_n311_), .Y(mai_mai_n542_));
  OAI210     m0520(.A0(mai_mai_n542_), .A1(mai_mai_n540_), .B0(mai_mai_n539_), .Y(mai_mai_n543_));
  OAI210     m0521(.A0(mai_mai_n543_), .A1(mai_mai_n538_), .B0(mai_mai_n450_), .Y(mai_mai_n544_));
  NA4        m0522(.A(mai_mai_n544_), .B(mai_mai_n537_), .C(mai_mai_n534_), .D(mai_mai_n528_), .Y(mai_mai_n545_));
  NA3        m0523(.A(mai_mai_n223_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n546_));
  NA2        m0524(.A(mai_mai_n286_), .B(mai_mai_n85_), .Y(mai_mai_n547_));
  AOI210     m0525(.A0(mai_mai_n546_), .A1(mai_mai_n341_), .B0(mai_mai_n547_), .Y(mai_mai_n548_));
  NA2        m0526(.A(mai_mai_n292_), .B(mai_mai_n288_), .Y(mai_mai_n549_));
  NO2        m0527(.A(mai_mai_n549_), .B(mai_mai_n177_), .Y(mai_mai_n550_));
  NA2        m0528(.A(mai_mai_n229_), .B(mai_mai_n228_), .Y(mai_mai_n551_));
  NA2        m0529(.A(mai_mai_n434_), .B(mai_mai_n227_), .Y(mai_mai_n552_));
  NO2        m0530(.A(mai_mai_n551_), .B(mai_mai_n552_), .Y(mai_mai_n553_));
  AOI210     m0531(.A0(i_6_), .A1(mai_mai_n47_), .B0(mai_mai_n363_), .Y(mai_mai_n554_));
  NA2        m0532(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n555_));
  NA3        m0533(.A(mai_mai_n524_), .B(mai_mai_n281_), .C(mai_mai_n555_), .Y(mai_mai_n556_));
  NO2        m0534(.A(mai_mai_n554_), .B(mai_mai_n556_), .Y(mai_mai_n557_));
  NO4        m0535(.A(mai_mai_n557_), .B(mai_mai_n553_), .C(mai_mai_n550_), .D(mai_mai_n548_), .Y(mai_mai_n558_));
  NO4        m0536(.A(mai_mai_n255_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n559_));
  NO3        m0537(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n560_));
  NO2        m0538(.A(mai_mai_n236_), .B(mai_mai_n36_), .Y(mai_mai_n561_));
  AN2        m0539(.A(mai_mai_n561_), .B(mai_mai_n560_), .Y(mai_mai_n562_));
  OA210      m0540(.A0(mai_mai_n562_), .A1(mai_mai_n559_), .B0(mai_mai_n351_), .Y(mai_mai_n563_));
  NO2        m0541(.A(mai_mai_n409_), .B(i_1_), .Y(mai_mai_n564_));
  NOi31      m0542(.An(mai_mai_n564_), .B(mai_mai_n442_), .C(mai_mai_n74_), .Y(mai_mai_n565_));
  AN4        m0543(.A(mai_mai_n565_), .B(mai_mai_n406_), .C(mai_mai_n490_), .D(i_2_), .Y(mai_mai_n566_));
  NO2        m0544(.A(mai_mai_n420_), .B(mai_mai_n181_), .Y(mai_mai_n567_));
  NO3        m0545(.A(mai_mai_n567_), .B(mai_mai_n566_), .C(mai_mai_n563_), .Y(mai_mai_n568_));
  NOi21      m0546(.An(i_10_), .B(i_6_), .Y(mai_mai_n569_));
  NO2        m0547(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n570_));
  AOI220     m0548(.A0(mai_mai_n286_), .A1(mai_mai_n570_), .B0(mai_mai_n281_), .B1(mai_mai_n569_), .Y(mai_mai_n571_));
  NO2        m0549(.A(mai_mai_n571_), .B(mai_mai_n440_), .Y(mai_mai_n572_));
  NO2        m0550(.A(mai_mai_n119_), .B(mai_mai_n23_), .Y(mai_mai_n573_));
  NO2        m0551(.A(mai_mai_n200_), .B(mai_mai_n37_), .Y(mai_mai_n574_));
  NOi31      m0552(.An(mai_mai_n151_), .B(mai_mai_n574_), .C(mai_mai_n323_), .Y(mai_mai_n575_));
  NO2        m0553(.A(mai_mai_n575_), .B(mai_mai_n572_), .Y(mai_mai_n576_));
  NO2        m0554(.A(mai_mai_n509_), .B(mai_mai_n374_), .Y(mai_mai_n577_));
  INV        m0555(.A(mai_mai_n311_), .Y(mai_mai_n578_));
  NO2        m0556(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n579_));
  NA2        m0557(.A(mai_mai_n178_), .B(i_0_), .Y(mai_mai_n580_));
  NO3        m0558(.A(mai_mai_n580_), .B(mai_mai_n333_), .C(mai_mai_n295_), .Y(mai_mai_n581_));
  OR2        m0559(.A(i_2_), .B(i_5_), .Y(mai_mai_n582_));
  OR2        m0560(.A(mai_mai_n582_), .B(mai_mai_n401_), .Y(mai_mai_n583_));
  NO2        m0561(.A(mai_mai_n583_), .B(mai_mai_n488_), .Y(mai_mai_n584_));
  NO3        m0562(.A(mai_mai_n584_), .B(mai_mai_n581_), .C(mai_mai_n577_), .Y(mai_mai_n585_));
  NA4        m0563(.A(mai_mai_n585_), .B(mai_mai_n576_), .C(mai_mai_n568_), .D(mai_mai_n558_), .Y(mai_mai_n586_));
  NO4        m0564(.A(mai_mai_n586_), .B(mai_mai_n545_), .C(mai_mai_n521_), .D(mai_mai_n498_), .Y(mai_mai_n587_));
  NA4        m0565(.A(mai_mai_n587_), .B(mai_mai_n431_), .C(mai_mai_n350_), .D(mai_mai_n307_), .Y(mai7));
  NO2        m0566(.A(mai_mai_n96_), .B(mai_mai_n55_), .Y(mai_mai_n589_));
  NO2        m0567(.A(mai_mai_n112_), .B(mai_mai_n93_), .Y(mai_mai_n590_));
  NA2        m0568(.A(mai_mai_n476_), .B(mai_mai_n85_), .Y(mai_mai_n591_));
  NA2        m0569(.A(i_11_), .B(mai_mai_n195_), .Y(mai_mai_n592_));
  NA3        m0570(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n593_));
  NO2        m0571(.A(mai_mai_n240_), .B(i_4_), .Y(mai_mai_n594_));
  NA2        m0572(.A(mai_mai_n594_), .B(i_8_), .Y(mai_mai_n595_));
  NO2        m0573(.A(mai_mai_n109_), .B(mai_mai_n593_), .Y(mai_mai_n596_));
  NA2        m0574(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n597_));
  OAI210     m0575(.A0(mai_mai_n90_), .A1(mai_mai_n205_), .B0(mai_mai_n206_), .Y(mai_mai_n598_));
  NO2        m0576(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n599_));
  NA2        m0577(.A(i_4_), .B(i_8_), .Y(mai_mai_n600_));
  AOI210     m0578(.A0(mai_mai_n600_), .A1(mai_mai_n301_), .B0(mai_mai_n599_), .Y(mai_mai_n601_));
  OAI220     m0579(.A0(mai_mai_n601_), .A1(mai_mai_n597_), .B0(mai_mai_n598_), .B1(i_13_), .Y(mai_mai_n602_));
  NO3        m0580(.A(mai_mai_n602_), .B(mai_mai_n596_), .C(mai_mai_n589_), .Y(mai_mai_n603_));
  AOI210     m0581(.A0(mai_mai_n133_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n604_));
  AOI210     m0582(.A0(mai_mai_n604_), .A1(mai_mai_n240_), .B0(mai_mai_n167_), .Y(mai_mai_n605_));
  OR2        m0583(.A(i_6_), .B(i_10_), .Y(mai_mai_n606_));
  NO2        m0584(.A(mai_mai_n606_), .B(mai_mai_n23_), .Y(mai_mai_n607_));
  OR3        m0585(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n608_));
  NO3        m0586(.A(mai_mai_n608_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n609_));
  INV        m0587(.A(mai_mai_n202_), .Y(mai_mai_n610_));
  NO2        m0588(.A(mai_mai_n609_), .B(mai_mai_n607_), .Y(mai_mai_n611_));
  OA220      m0589(.A0(mai_mai_n611_), .A1(mai_mai_n578_), .B0(mai_mai_n605_), .B1(mai_mai_n274_), .Y(mai_mai_n612_));
  AOI210     m0590(.A0(mai_mai_n612_), .A1(mai_mai_n603_), .B0(mai_mai_n64_), .Y(mai_mai_n613_));
  NOi21      m0591(.An(i_11_), .B(i_7_), .Y(mai_mai_n614_));
  AO210      m0592(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n615_));
  NO2        m0593(.A(mai_mai_n615_), .B(mai_mai_n614_), .Y(mai_mai_n616_));
  NA2        m0594(.A(mai_mai_n616_), .B(mai_mai_n210_), .Y(mai_mai_n617_));
  NO2        m0595(.A(mai_mai_n617_), .B(mai_mai_n64_), .Y(mai_mai_n618_));
  NA2        m0596(.A(mai_mai_n89_), .B(mai_mai_n64_), .Y(mai_mai_n619_));
  AO210      m0597(.A0(mai_mai_n619_), .A1(mai_mai_n374_), .B0(mai_mai_n41_), .Y(mai_mai_n620_));
  NO3        m0598(.A(mai_mai_n263_), .B(mai_mai_n212_), .C(mai_mai_n592_), .Y(mai_mai_n621_));
  OAI210     m0599(.A0(mai_mai_n621_), .A1(mai_mai_n231_), .B0(mai_mai_n64_), .Y(mai_mai_n622_));
  NA2        m0600(.A(mai_mai_n402_), .B(mai_mai_n31_), .Y(mai_mai_n623_));
  OR2        m0601(.A(mai_mai_n212_), .B(mai_mai_n112_), .Y(mai_mai_n624_));
  NA2        m0602(.A(mai_mai_n624_), .B(mai_mai_n623_), .Y(mai_mai_n625_));
  NO2        m0603(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n626_));
  NO2        m0604(.A(mai_mai_n626_), .B(i_4_), .Y(mai_mai_n627_));
  NA2        m0605(.A(mai_mai_n627_), .B(mai_mai_n625_), .Y(mai_mai_n628_));
  NO2        m0606(.A(i_1_), .B(i_12_), .Y(mai_mai_n629_));
  NA3        m0607(.A(mai_mai_n629_), .B(mai_mai_n114_), .C(mai_mai_n24_), .Y(mai_mai_n630_));
  BUFFER     m0608(.A(mai_mai_n630_), .Y(mai_mai_n631_));
  NA4        m0609(.A(mai_mai_n631_), .B(mai_mai_n628_), .C(mai_mai_n622_), .D(mai_mai_n620_), .Y(mai_mai_n632_));
  OAI210     m0610(.A0(mai_mai_n632_), .A1(mai_mai_n618_), .B0(i_6_), .Y(mai_mai_n633_));
  NO2        m0611(.A(i_6_), .B(i_11_), .Y(mai_mai_n634_));
  INV        m0612(.A(mai_mai_n443_), .Y(mai_mai_n635_));
  NO4        m0613(.A(mai_mai_n220_), .B(mai_mai_n133_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n636_));
  NA2        m0614(.A(mai_mai_n636_), .B(mai_mai_n626_), .Y(mai_mai_n637_));
  NA2        m0615(.A(mai_mai_n240_), .B(i_6_), .Y(mai_mai_n638_));
  NO3        m0616(.A(mai_mai_n606_), .B(mai_mai_n236_), .C(mai_mai_n23_), .Y(mai_mai_n639_));
  AOI210     m0617(.A0(i_1_), .A1(mai_mai_n264_), .B0(mai_mai_n639_), .Y(mai_mai_n640_));
  OAI210     m0618(.A0(mai_mai_n640_), .A1(mai_mai_n45_), .B0(mai_mai_n637_), .Y(mai_mai_n641_));
  INV        m0619(.A(i_2_), .Y(mai_mai_n642_));
  NA2        m0620(.A(mai_mai_n143_), .B(i_9_), .Y(mai_mai_n643_));
  NA3        m0621(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n644_));
  NO2        m0622(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n645_));
  NA3        m0623(.A(mai_mai_n645_), .B(mai_mai_n273_), .C(mai_mai_n45_), .Y(mai_mai_n646_));
  OAI220     m0624(.A0(mai_mai_n646_), .A1(mai_mai_n644_), .B0(mai_mai_n643_), .B1(mai_mai_n642_), .Y(mai_mai_n647_));
  NA3        m0625(.A(mai_mai_n626_), .B(mai_mai_n311_), .C(i_6_), .Y(mai_mai_n648_));
  NO2        m0626(.A(mai_mai_n648_), .B(mai_mai_n23_), .Y(mai_mai_n649_));
  AOI210     m0627(.A0(mai_mai_n467_), .A1(mai_mai_n413_), .B0(mai_mai_n245_), .Y(mai_mai_n650_));
  NO2        m0628(.A(mai_mai_n650_), .B(mai_mai_n597_), .Y(mai_mai_n651_));
  NO2        m0629(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n652_));
  OR3        m0630(.A(mai_mai_n651_), .B(mai_mai_n649_), .C(mai_mai_n647_), .Y(mai_mai_n653_));
  NO3        m0631(.A(mai_mai_n653_), .B(mai_mai_n641_), .C(mai_mai_n635_), .Y(mai_mai_n654_));
  NO2        m0632(.A(mai_mai_n240_), .B(mai_mai_n105_), .Y(mai_mai_n655_));
  NO2        m0633(.A(mai_mai_n655_), .B(mai_mai_n614_), .Y(mai_mai_n656_));
  NA2        m0634(.A(mai_mai_n656_), .B(i_1_), .Y(mai_mai_n657_));
  NO2        m0635(.A(mai_mai_n657_), .B(mai_mai_n608_), .Y(mai_mai_n658_));
  NO2        m0636(.A(mai_mai_n408_), .B(mai_mai_n87_), .Y(mai_mai_n659_));
  NA2        m0637(.A(mai_mai_n658_), .B(mai_mai_n47_), .Y(mai_mai_n660_));
  NA2        m0638(.A(i_3_), .B(mai_mai_n195_), .Y(mai_mai_n661_));
  NO2        m0639(.A(mai_mai_n661_), .B(mai_mai_n119_), .Y(mai_mai_n662_));
  AN2        m0640(.A(mai_mai_n662_), .B(mai_mai_n533_), .Y(mai_mai_n663_));
  NO2        m0641(.A(mai_mai_n236_), .B(mai_mai_n45_), .Y(mai_mai_n664_));
  NO3        m0642(.A(mai_mai_n664_), .B(mai_mai_n304_), .C(mai_mai_n241_), .Y(mai_mai_n665_));
  NO2        m0643(.A(mai_mai_n122_), .B(mai_mai_n37_), .Y(mai_mai_n666_));
  NO2        m0644(.A(mai_mai_n666_), .B(i_6_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n668_));
  NO2        m0646(.A(mai_mai_n668_), .B(mai_mai_n64_), .Y(mai_mai_n669_));
  NO2        m0647(.A(mai_mai_n669_), .B(mai_mai_n629_), .Y(mai_mai_n670_));
  NO4        m0648(.A(mai_mai_n670_), .B(mai_mai_n667_), .C(mai_mai_n665_), .D(i_4_), .Y(mai_mai_n671_));
  NA2        m0649(.A(i_1_), .B(i_3_), .Y(mai_mai_n672_));
  NO2        m0650(.A(mai_mai_n444_), .B(mai_mai_n96_), .Y(mai_mai_n673_));
  AOI210     m0651(.A0(mai_mai_n664_), .A1(mai_mai_n569_), .B0(mai_mai_n673_), .Y(mai_mai_n674_));
  NO2        m0652(.A(mai_mai_n674_), .B(mai_mai_n672_), .Y(mai_mai_n675_));
  NO3        m0653(.A(mai_mai_n675_), .B(mai_mai_n671_), .C(mai_mai_n663_), .Y(mai_mai_n676_));
  NA4        m0654(.A(mai_mai_n676_), .B(mai_mai_n660_), .C(mai_mai_n654_), .D(mai_mai_n633_), .Y(mai_mai_n677_));
  NO3        m0655(.A(mai_mai_n469_), .B(i_3_), .C(i_7_), .Y(mai_mai_n678_));
  NOi21      m0656(.An(mai_mai_n678_), .B(i_10_), .Y(mai_mai_n679_));
  OA210      m0657(.A0(mai_mai_n679_), .A1(mai_mai_n248_), .B0(mai_mai_n87_), .Y(mai_mai_n680_));
  NA2        m0658(.A(mai_mai_n366_), .B(mai_mai_n365_), .Y(mai_mai_n681_));
  NA3        m0659(.A(mai_mai_n476_), .B(mai_mai_n512_), .C(mai_mai_n47_), .Y(mai_mai_n682_));
  NA3        m0660(.A(mai_mai_n167_), .B(mai_mai_n85_), .C(mai_mai_n87_), .Y(mai_mai_n683_));
  NA3        m0661(.A(mai_mai_n683_), .B(mai_mai_n682_), .C(mai_mai_n681_), .Y(mai_mai_n684_));
  OAI210     m0662(.A0(mai_mai_n684_), .A1(mai_mai_n680_), .B0(i_1_), .Y(mai_mai_n685_));
  AOI210     m0663(.A0(mai_mai_n273_), .A1(mai_mai_n101_), .B0(i_1_), .Y(mai_mai_n686_));
  NO2        m0664(.A(mai_mai_n364_), .B(i_2_), .Y(mai_mai_n687_));
  NA2        m0665(.A(mai_mai_n687_), .B(mai_mai_n686_), .Y(mai_mai_n688_));
  OAI210     m0666(.A0(mai_mai_n648_), .A1(mai_mai_n435_), .B0(mai_mai_n688_), .Y(mai_mai_n689_));
  INV        m0667(.A(mai_mai_n689_), .Y(mai_mai_n690_));
  AOI210     m0668(.A0(mai_mai_n690_), .A1(mai_mai_n685_), .B0(i_13_), .Y(mai_mai_n691_));
  OR2        m0669(.A(i_11_), .B(i_7_), .Y(mai_mai_n692_));
  AOI210     m0670(.A0(mai_mai_n644_), .A1(mai_mai_n55_), .B0(i_12_), .Y(mai_mai_n693_));
  NO2        m0671(.A(mai_mai_n470_), .B(mai_mai_n24_), .Y(mai_mai_n694_));
  AOI220     m0672(.A0(mai_mai_n694_), .A1(mai_mai_n659_), .B0(mai_mai_n248_), .B1(mai_mai_n136_), .Y(mai_mai_n695_));
  OAI220     m0673(.A0(mai_mai_n695_), .A1(mai_mai_n41_), .B0(mai_mai_n1048_), .B1(mai_mai_n96_), .Y(mai_mai_n696_));
  INV        m0674(.A(mai_mai_n696_), .Y(mai_mai_n697_));
  INV        m0675(.A(mai_mai_n119_), .Y(mai_mai_n698_));
  AOI220     m0676(.A0(mai_mai_n698_), .A1(mai_mai_n73_), .B0(mai_mai_n381_), .B1(mai_mai_n645_), .Y(mai_mai_n699_));
  NO2        m0677(.A(mai_mai_n699_), .B(mai_mai_n246_), .Y(mai_mai_n700_));
  AOI210     m0678(.A0(mai_mai_n435_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n701_));
  NOi31      m0679(.An(mai_mai_n701_), .B(mai_mai_n591_), .C(mai_mai_n45_), .Y(mai_mai_n702_));
  NA2        m0680(.A(mai_mai_n132_), .B(i_13_), .Y(mai_mai_n703_));
  NO2        m0681(.A(mai_mai_n644_), .B(mai_mai_n119_), .Y(mai_mai_n704_));
  INV        m0682(.A(mai_mai_n704_), .Y(mai_mai_n705_));
  OAI220     m0683(.A0(mai_mai_n705_), .A1(mai_mai_n72_), .B0(mai_mai_n703_), .B1(mai_mai_n686_), .Y(mai_mai_n706_));
  NO3        m0684(.A(mai_mai_n72_), .B(mai_mai_n32_), .C(mai_mai_n105_), .Y(mai_mai_n707_));
  NA2        m0685(.A(mai_mai_n26_), .B(mai_mai_n195_), .Y(mai_mai_n708_));
  NA2        m0686(.A(mai_mai_n708_), .B(i_7_), .Y(mai_mai_n709_));
  NO3        m0687(.A(mai_mai_n470_), .B(mai_mai_n240_), .C(mai_mai_n87_), .Y(mai_mai_n710_));
  AOI210     m0688(.A0(mai_mai_n710_), .A1(mai_mai_n709_), .B0(mai_mai_n707_), .Y(mai_mai_n711_));
  AOI220     m0689(.A0(mai_mai_n381_), .A1(mai_mai_n645_), .B0(mai_mai_n95_), .B1(mai_mai_n106_), .Y(mai_mai_n712_));
  OAI220     m0690(.A0(mai_mai_n712_), .A1(mai_mai_n595_), .B0(mai_mai_n711_), .B1(mai_mai_n610_), .Y(mai_mai_n713_));
  NO4        m0691(.A(mai_mai_n713_), .B(mai_mai_n706_), .C(mai_mai_n702_), .D(mai_mai_n700_), .Y(mai_mai_n714_));
  OR2        m0692(.A(i_11_), .B(i_6_), .Y(mai_mai_n715_));
  NA3        m0693(.A(mai_mai_n594_), .B(mai_mai_n708_), .C(i_7_), .Y(mai_mai_n716_));
  AOI210     m0694(.A0(mai_mai_n716_), .A1(mai_mai_n705_), .B0(mai_mai_n715_), .Y(mai_mai_n717_));
  NA3        m0695(.A(mai_mai_n402_), .B(mai_mai_n599_), .C(mai_mai_n101_), .Y(mai_mai_n718_));
  NA2        m0696(.A(mai_mai_n634_), .B(i_13_), .Y(mai_mai_n719_));
  NA2        m0697(.A(mai_mai_n106_), .B(mai_mai_n708_), .Y(mai_mai_n720_));
  NAi21      m0698(.An(i_11_), .B(i_12_), .Y(mai_mai_n721_));
  NOi41      m0699(.An(mai_mai_n115_), .B(mai_mai_n721_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n722_));
  NA2        m0700(.A(mai_mai_n722_), .B(mai_mai_n720_), .Y(mai_mai_n723_));
  NA3        m0701(.A(mai_mai_n723_), .B(mai_mai_n719_), .C(mai_mai_n718_), .Y(mai_mai_n724_));
  OAI210     m0702(.A0(mai_mai_n724_), .A1(mai_mai_n717_), .B0(mai_mai_n64_), .Y(mai_mai_n725_));
  NO2        m0703(.A(i_2_), .B(i_12_), .Y(mai_mai_n726_));
  NA2        m0704(.A(mai_mai_n363_), .B(mai_mai_n726_), .Y(mai_mai_n727_));
  NA2        m0705(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n728_));
  NO3        m0706(.A(mai_mai_n728_), .B(mai_mai_n379_), .C(mai_mai_n594_), .Y(mai_mai_n729_));
  OAI210     m0707(.A0(mai_mai_n729_), .A1(mai_mai_n365_), .B0(mai_mai_n363_), .Y(mai_mai_n730_));
  NO2        m0708(.A(mai_mai_n133_), .B(i_2_), .Y(mai_mai_n731_));
  NA2        m0709(.A(mai_mai_n731_), .B(mai_mai_n629_), .Y(mai_mai_n732_));
  NA3        m0710(.A(mai_mai_n732_), .B(mai_mai_n730_), .C(mai_mai_n727_), .Y(mai_mai_n733_));
  NA3        m0711(.A(mai_mai_n733_), .B(mai_mai_n46_), .C(mai_mai_n230_), .Y(mai_mai_n734_));
  NA4        m0712(.A(mai_mai_n734_), .B(mai_mai_n725_), .C(mai_mai_n714_), .D(mai_mai_n697_), .Y(mai_mai_n735_));
  OR4        m0713(.A(mai_mai_n735_), .B(mai_mai_n691_), .C(mai_mai_n677_), .D(mai_mai_n613_), .Y(mai5));
  NA2        m0714(.A(mai_mai_n656_), .B(mai_mai_n276_), .Y(mai_mai_n737_));
  AN2        m0715(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n738_));
  NA3        m0716(.A(mai_mai_n738_), .B(mai_mai_n726_), .C(mai_mai_n112_), .Y(mai_mai_n739_));
  NO2        m0717(.A(mai_mai_n595_), .B(i_11_), .Y(mai_mai_n740_));
  NA2        m0718(.A(mai_mai_n90_), .B(mai_mai_n740_), .Y(mai_mai_n741_));
  NA3        m0719(.A(mai_mai_n741_), .B(mai_mai_n739_), .C(mai_mai_n737_), .Y(mai_mai_n742_));
  NO3        m0720(.A(i_11_), .B(mai_mai_n240_), .C(i_13_), .Y(mai_mai_n743_));
  NO2        m0721(.A(mai_mai_n129_), .B(mai_mai_n23_), .Y(mai_mai_n744_));
  NA2        m0722(.A(i_12_), .B(i_8_), .Y(mai_mai_n745_));
  OAI210     m0723(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n745_), .Y(mai_mai_n746_));
  INV        m0724(.A(mai_mai_n434_), .Y(mai_mai_n747_));
  AOI220     m0725(.A0(mai_mai_n311_), .A1(mai_mai_n573_), .B0(mai_mai_n746_), .B1(mai_mai_n744_), .Y(mai_mai_n748_));
  INV        m0726(.A(mai_mai_n748_), .Y(mai_mai_n749_));
  NO2        m0727(.A(mai_mai_n749_), .B(mai_mai_n742_), .Y(mai_mai_n750_));
  INV        m0728(.A(mai_mai_n175_), .Y(mai_mai_n751_));
  INV        m0729(.A(mai_mai_n248_), .Y(mai_mai_n752_));
  OAI210     m0730(.A0(mai_mai_n687_), .A1(mai_mai_n436_), .B0(mai_mai_n115_), .Y(mai_mai_n753_));
  AOI210     m0731(.A0(mai_mai_n753_), .A1(mai_mai_n752_), .B0(mai_mai_n751_), .Y(mai_mai_n754_));
  NO2        m0732(.A(mai_mai_n444_), .B(mai_mai_n26_), .Y(mai_mai_n755_));
  NO2        m0733(.A(mai_mai_n755_), .B(mai_mai_n413_), .Y(mai_mai_n756_));
  NA2        m0734(.A(mai_mai_n756_), .B(i_2_), .Y(mai_mai_n757_));
  INV        m0735(.A(mai_mai_n757_), .Y(mai_mai_n758_));
  AOI210     m0736(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n409_), .Y(mai_mai_n759_));
  AOI210     m0737(.A0(mai_mai_n759_), .A1(mai_mai_n758_), .B0(mai_mai_n754_), .Y(mai_mai_n760_));
  NO2        m0738(.A(mai_mai_n192_), .B(mai_mai_n130_), .Y(mai_mai_n761_));
  OAI210     m0739(.A0(mai_mai_n761_), .A1(mai_mai_n744_), .B0(i_2_), .Y(mai_mai_n762_));
  INV        m0740(.A(mai_mai_n176_), .Y(mai_mai_n763_));
  NO3        m0741(.A(mai_mai_n615_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n764_));
  AOI210     m0742(.A0(mai_mai_n763_), .A1(mai_mai_n90_), .B0(mai_mai_n764_), .Y(mai_mai_n765_));
  AOI210     m0743(.A0(mai_mai_n765_), .A1(mai_mai_n762_), .B0(mai_mai_n195_), .Y(mai_mai_n766_));
  OA210      m0744(.A0(mai_mai_n616_), .A1(mai_mai_n131_), .B0(i_13_), .Y(mai_mai_n767_));
  NA2        m0745(.A(mai_mai_n202_), .B(mai_mai_n205_), .Y(mai_mai_n768_));
  NA2        m0746(.A(mai_mai_n157_), .B(mai_mai_n592_), .Y(mai_mai_n769_));
  AOI210     m0747(.A0(mai_mai_n769_), .A1(mai_mai_n768_), .B0(mai_mai_n368_), .Y(mai_mai_n770_));
  AOI210     m0748(.A0(mai_mai_n212_), .A1(mai_mai_n153_), .B0(mai_mai_n512_), .Y(mai_mai_n771_));
  NA2        m0749(.A(mai_mai_n771_), .B(mai_mai_n413_), .Y(mai_mai_n772_));
  NO2        m0750(.A(mai_mai_n106_), .B(mai_mai_n45_), .Y(mai_mai_n773_));
  INV        m0751(.A(mai_mai_n296_), .Y(mai_mai_n774_));
  NA4        m0752(.A(mai_mai_n774_), .B(mai_mai_n301_), .C(mai_mai_n129_), .D(mai_mai_n43_), .Y(mai_mai_n775_));
  OAI210     m0753(.A0(mai_mai_n775_), .A1(mai_mai_n773_), .B0(mai_mai_n772_), .Y(mai_mai_n776_));
  NO4        m0754(.A(mai_mai_n776_), .B(mai_mai_n770_), .C(mai_mai_n767_), .D(mai_mai_n766_), .Y(mai_mai_n777_));
  NA2        m0755(.A(mai_mai_n573_), .B(mai_mai_n28_), .Y(mai_mai_n778_));
  NA2        m0756(.A(mai_mai_n743_), .B(mai_mai_n282_), .Y(mai_mai_n779_));
  NA2        m0757(.A(mai_mai_n779_), .B(mai_mai_n778_), .Y(mai_mai_n780_));
  NO2        m0758(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n781_));
  NO2        m0759(.A(mai_mai_n781_), .B(mai_mai_n131_), .Y(mai_mai_n782_));
  NO2        m0760(.A(mai_mai_n782_), .B(mai_mai_n592_), .Y(mai_mai_n783_));
  AOI220     m0761(.A0(mai_mai_n783_), .A1(mai_mai_n36_), .B0(mai_mai_n780_), .B1(mai_mai_n47_), .Y(mai_mai_n784_));
  NA4        m0762(.A(mai_mai_n784_), .B(mai_mai_n777_), .C(mai_mai_n760_), .D(mai_mai_n750_), .Y(mai6));
  NO2        m0763(.A(mai_mai_n187_), .B(mai_mai_n144_), .Y(mai_mai_n786_));
  NA2        m0764(.A(mai_mai_n786_), .B(mai_mai_n731_), .Y(mai_mai_n787_));
  NA4        m0765(.A(mai_mai_n383_), .B(mai_mai_n475_), .C(mai_mai_n72_), .D(mai_mai_n105_), .Y(mai_mai_n788_));
  INV        m0766(.A(mai_mai_n788_), .Y(mai_mai_n789_));
  NO2        m0767(.A(mai_mai_n226_), .B(mai_mai_n480_), .Y(mai_mai_n790_));
  NO2        m0768(.A(i_11_), .B(i_9_), .Y(mai_mai_n791_));
  NO2        m0769(.A(mai_mai_n789_), .B(mai_mai_n322_), .Y(mai_mai_n792_));
  AO210      m0770(.A0(mai_mai_n792_), .A1(mai_mai_n787_), .B0(i_12_), .Y(mai_mai_n793_));
  NA2        m0771(.A(mai_mai_n369_), .B(mai_mai_n327_), .Y(mai_mai_n794_));
  NA2        m0772(.A(mai_mai_n579_), .B(mai_mai_n64_), .Y(mai_mai_n795_));
  NA2        m0773(.A(mai_mai_n679_), .B(mai_mai_n72_), .Y(mai_mai_n796_));
  BUFFER     m0774(.A(mai_mai_n619_), .Y(mai_mai_n797_));
  NA4        m0775(.A(mai_mai_n797_), .B(mai_mai_n796_), .C(mai_mai_n795_), .D(mai_mai_n794_), .Y(mai_mai_n798_));
  INV        m0776(.A(mai_mai_n199_), .Y(mai_mai_n799_));
  AOI220     m0777(.A0(mai_mai_n799_), .A1(mai_mai_n791_), .B0(mai_mai_n798_), .B1(mai_mai_n74_), .Y(mai_mai_n800_));
  INV        m0778(.A(mai_mai_n321_), .Y(mai_mai_n801_));
  NA2        m0779(.A(mai_mai_n76_), .B(mai_mai_n136_), .Y(mai_mai_n802_));
  INV        m0780(.A(mai_mai_n129_), .Y(mai_mai_n803_));
  NA2        m0781(.A(mai_mai_n803_), .B(mai_mai_n47_), .Y(mai_mai_n804_));
  AOI210     m0782(.A0(mai_mai_n804_), .A1(mai_mai_n802_), .B0(mai_mai_n801_), .Y(mai_mai_n805_));
  NO3        m0783(.A(mai_mai_n255_), .B(mai_mai_n137_), .C(i_9_), .Y(mai_mai_n806_));
  NA2        m0784(.A(mai_mai_n806_), .B(mai_mai_n781_), .Y(mai_mai_n807_));
  AOI210     m0785(.A0(mai_mai_n807_), .A1(mai_mai_n510_), .B0(mai_mai_n187_), .Y(mai_mai_n808_));
  NO2        m0786(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n809_));
  NA3        m0787(.A(mai_mai_n809_), .B(mai_mai_n465_), .C(mai_mai_n383_), .Y(mai_mai_n810_));
  NAi32      m0788(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n811_));
  NO2        m0789(.A(mai_mai_n715_), .B(mai_mai_n811_), .Y(mai_mai_n812_));
  OAI210     m0790(.A0(mai_mai_n678_), .A1(mai_mai_n561_), .B0(mai_mai_n560_), .Y(mai_mai_n813_));
  NAi31      m0791(.An(mai_mai_n812_), .B(mai_mai_n813_), .C(mai_mai_n810_), .Y(mai_mai_n814_));
  OR3        m0792(.A(mai_mai_n814_), .B(mai_mai_n808_), .C(mai_mai_n805_), .Y(mai_mai_n815_));
  NO2        m0793(.A(mai_mai_n692_), .B(i_2_), .Y(mai_mai_n816_));
  NA2        m0794(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n817_));
  NO2        m0795(.A(mai_mai_n817_), .B(mai_mai_n401_), .Y(mai_mai_n818_));
  NA2        m0796(.A(mai_mai_n818_), .B(mai_mai_n816_), .Y(mai_mai_n819_));
  AO220      m0797(.A0(mai_mai_n355_), .A1(mai_mai_n345_), .B0(mai_mai_n385_), .B1(mai_mai_n592_), .Y(mai_mai_n820_));
  NA3        m0798(.A(mai_mai_n820_), .B(mai_mai_n260_), .C(i_7_), .Y(mai_mai_n821_));
  NA3        m0799(.A(mai_mai_n616_), .B(mai_mai_n152_), .C(mai_mai_n70_), .Y(mai_mai_n822_));
  AO210      m0800(.A0(mai_mai_n487_), .A1(mai_mai_n747_), .B0(mai_mai_n36_), .Y(mai_mai_n823_));
  NA4        m0801(.A(mai_mai_n823_), .B(mai_mai_n822_), .C(mai_mai_n821_), .D(mai_mai_n819_), .Y(mai_mai_n824_));
  OAI210     m0802(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n88_), .Y(mai_mai_n825_));
  AOI220     m0803(.A0(mai_mai_n825_), .A1(mai_mai_n560_), .B0(mai_mai_n790_), .B1(mai_mai_n709_), .Y(mai_mai_n826_));
  NA3        m0804(.A(mai_mai_n368_), .B(mai_mai_n242_), .C(mai_mai_n152_), .Y(mai_mai_n827_));
  NA2        m0805(.A(mai_mai_n385_), .B(mai_mai_n71_), .Y(mai_mai_n828_));
  NA4        m0806(.A(mai_mai_n828_), .B(mai_mai_n827_), .C(mai_mai_n826_), .D(mai_mai_n598_), .Y(mai_mai_n829_));
  AO210      m0807(.A0(mai_mai_n512_), .A1(mai_mai_n47_), .B0(mai_mai_n89_), .Y(mai_mai_n830_));
  NA3        m0808(.A(mai_mai_n830_), .B(mai_mai_n476_), .C(mai_mai_n223_), .Y(mai_mai_n831_));
  AOI210     m0809(.A0(mai_mai_n436_), .A1(mai_mai_n434_), .B0(mai_mai_n559_), .Y(mai_mai_n832_));
  NO2        m0810(.A(mai_mai_n606_), .B(mai_mai_n106_), .Y(mai_mai_n833_));
  OAI210     m0811(.A0(mai_mai_n833_), .A1(mai_mai_n116_), .B0(mai_mai_n399_), .Y(mai_mai_n834_));
  INV        m0812(.A(mai_mai_n583_), .Y(mai_mai_n835_));
  NA3        m0813(.A(mai_mai_n835_), .B(mai_mai_n321_), .C(i_7_), .Y(mai_mai_n836_));
  NA4        m0814(.A(mai_mai_n836_), .B(mai_mai_n834_), .C(mai_mai_n832_), .D(mai_mai_n831_), .Y(mai_mai_n837_));
  NO4        m0815(.A(mai_mai_n837_), .B(mai_mai_n829_), .C(mai_mai_n824_), .D(mai_mai_n815_), .Y(mai_mai_n838_));
  NA4        m0816(.A(mai_mai_n838_), .B(mai_mai_n800_), .C(mai_mai_n793_), .D(mai_mai_n376_), .Y(mai3));
  NA2        m0817(.A(i_6_), .B(i_7_), .Y(mai_mai_n840_));
  NO2        m0818(.A(mai_mai_n840_), .B(i_0_), .Y(mai_mai_n841_));
  NO2        m0819(.A(i_11_), .B(mai_mai_n240_), .Y(mai_mai_n842_));
  OAI210     m0820(.A0(mai_mai_n841_), .A1(mai_mai_n289_), .B0(mai_mai_n842_), .Y(mai_mai_n843_));
  NO2        m0821(.A(mai_mai_n843_), .B(mai_mai_n195_), .Y(mai_mai_n844_));
  NO3        m0822(.A(mai_mai_n440_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n845_));
  OA210      m0823(.A0(mai_mai_n845_), .A1(mai_mai_n844_), .B0(mai_mai_n178_), .Y(mai_mai_n846_));
  NA3        m0824(.A(mai_mai_n827_), .B(mai_mai_n598_), .C(mai_mai_n367_), .Y(mai_mai_n847_));
  NA2        m0825(.A(mai_mai_n847_), .B(mai_mai_n40_), .Y(mai_mai_n848_));
  NOi21      m0826(.An(mai_mai_n100_), .B(mai_mai_n756_), .Y(mai_mai_n849_));
  NO3        m0827(.A(mai_mai_n624_), .B(mai_mai_n444_), .C(mai_mai_n136_), .Y(mai_mai_n850_));
  NA2        m0828(.A(mai_mai_n402_), .B(mai_mai_n46_), .Y(mai_mai_n851_));
  AN2        m0829(.A(mai_mai_n442_), .B(mai_mai_n56_), .Y(mai_mai_n852_));
  NO3        m0830(.A(mai_mai_n852_), .B(mai_mai_n850_), .C(mai_mai_n849_), .Y(mai_mai_n853_));
  AOI210     m0831(.A0(mai_mai_n853_), .A1(mai_mai_n848_), .B0(mai_mai_n49_), .Y(mai_mai_n854_));
  NO4        m0832(.A(mai_mai_n372_), .B(mai_mai_n378_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n855_));
  NA2        m0833(.A(mai_mai_n187_), .B(mai_mai_n569_), .Y(mai_mai_n856_));
  NOi21      m0834(.An(mai_mai_n856_), .B(mai_mai_n855_), .Y(mai_mai_n857_));
  NO2        m0835(.A(mai_mai_n857_), .B(mai_mai_n64_), .Y(mai_mai_n858_));
  NOi21      m0836(.An(i_5_), .B(i_9_), .Y(mai_mai_n859_));
  NA2        m0837(.A(mai_mai_n859_), .B(mai_mai_n433_), .Y(mai_mai_n860_));
  BUFFER     m0838(.A(mai_mai_n273_), .Y(mai_mai_n861_));
  NA2        m0839(.A(mai_mai_n861_), .B(mai_mai_n467_), .Y(mai_mai_n862_));
  NO3        m0840(.A(mai_mai_n405_), .B(mai_mai_n273_), .C(mai_mai_n74_), .Y(mai_mai_n863_));
  NO2        m0841(.A(mai_mai_n179_), .B(mai_mai_n153_), .Y(mai_mai_n864_));
  AOI210     m0842(.A0(mai_mai_n864_), .A1(mai_mai_n247_), .B0(mai_mai_n863_), .Y(mai_mai_n865_));
  OAI220     m0843(.A0(mai_mai_n865_), .A1(mai_mai_n185_), .B0(mai_mai_n862_), .B1(mai_mai_n860_), .Y(mai_mai_n866_));
  NO4        m0844(.A(mai_mai_n866_), .B(mai_mai_n858_), .C(mai_mai_n854_), .D(mai_mai_n846_), .Y(mai_mai_n867_));
  NA2        m0845(.A(mai_mai_n187_), .B(mai_mai_n24_), .Y(mai_mai_n868_));
  NO2        m0846(.A(mai_mai_n666_), .B(mai_mai_n590_), .Y(mai_mai_n869_));
  NO2        m0847(.A(mai_mai_n869_), .B(mai_mai_n868_), .Y(mai_mai_n870_));
  INV        m0848(.A(mai_mai_n870_), .Y(mai_mai_n871_));
  NO2        m0849(.A(mai_mai_n383_), .B(mai_mai_n290_), .Y(mai_mai_n872_));
  NA2        m0850(.A(mai_mai_n872_), .B(mai_mai_n704_), .Y(mai_mai_n873_));
  NA2        m0851(.A(mai_mai_n570_), .B(i_0_), .Y(mai_mai_n874_));
  NO3        m0852(.A(mai_mai_n874_), .B(mai_mai_n380_), .C(mai_mai_n90_), .Y(mai_mai_n875_));
  NO4        m0853(.A(mai_mai_n582_), .B(mai_mai_n220_), .C(mai_mai_n409_), .D(mai_mai_n401_), .Y(mai_mai_n876_));
  AOI210     m0854(.A0(mai_mai_n876_), .A1(i_11_), .B0(mai_mai_n875_), .Y(mai_mai_n877_));
  NA2        m0855(.A(mai_mai_n743_), .B(mai_mai_n322_), .Y(mai_mai_n878_));
  AOI210     m0856(.A0(mai_mai_n476_), .A1(mai_mai_n90_), .B0(mai_mai_n59_), .Y(mai_mai_n879_));
  NO2        m0857(.A(mai_mai_n879_), .B(mai_mai_n878_), .Y(mai_mai_n880_));
  NO2        m0858(.A(mai_mai_n257_), .B(mai_mai_n159_), .Y(mai_mai_n881_));
  NA2        m0859(.A(i_0_), .B(i_10_), .Y(mai_mai_n882_));
  INV        m0860(.A(mai_mai_n532_), .Y(mai_mai_n883_));
  NO4        m0861(.A(mai_mai_n119_), .B(mai_mai_n59_), .C(mai_mai_n661_), .D(i_5_), .Y(mai_mai_n884_));
  AO220      m0862(.A0(mai_mai_n884_), .A1(mai_mai_n883_), .B0(mai_mai_n881_), .B1(i_6_), .Y(mai_mai_n885_));
  AOI220     m0863(.A0(mai_mai_n325_), .A1(mai_mai_n102_), .B0(mai_mai_n187_), .B1(mai_mai_n85_), .Y(mai_mai_n886_));
  NA2        m0864(.A(mai_mai_n564_), .B(i_4_), .Y(mai_mai_n887_));
  NA2        m0865(.A(mai_mai_n190_), .B(mai_mai_n205_), .Y(mai_mai_n888_));
  OAI220     m0866(.A0(mai_mai_n888_), .A1(mai_mai_n878_), .B0(mai_mai_n887_), .B1(mai_mai_n886_), .Y(mai_mai_n889_));
  NO3        m0867(.A(mai_mai_n889_), .B(mai_mai_n885_), .C(mai_mai_n880_), .Y(mai_mai_n890_));
  NA4        m0868(.A(mai_mai_n890_), .B(mai_mai_n877_), .C(mai_mai_n873_), .D(mai_mai_n871_), .Y(mai_mai_n891_));
  NO2        m0869(.A(mai_mai_n107_), .B(mai_mai_n37_), .Y(mai_mai_n892_));
  NA2        m0870(.A(i_11_), .B(i_9_), .Y(mai_mai_n893_));
  NO3        m0871(.A(i_12_), .B(mai_mai_n893_), .C(mai_mai_n597_), .Y(mai_mai_n894_));
  AN2        m0872(.A(mai_mai_n894_), .B(mai_mai_n892_), .Y(mai_mai_n895_));
  NO2        m0873(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n896_));
  NA2        m0874(.A(mai_mai_n384_), .B(mai_mai_n183_), .Y(mai_mai_n897_));
  NA2        m0875(.A(mai_mai_n897_), .B(mai_mai_n166_), .Y(mai_mai_n898_));
  NO2        m0876(.A(mai_mai_n893_), .B(mai_mai_n74_), .Y(mai_mai_n899_));
  NO2        m0877(.A(mai_mai_n179_), .B(i_0_), .Y(mai_mai_n900_));
  INV        m0878(.A(mai_mai_n900_), .Y(mai_mai_n901_));
  NA2        m0879(.A(mai_mai_n465_), .B(mai_mai_n234_), .Y(mai_mai_n902_));
  AOI210     m0880(.A0(mai_mai_n366_), .A1(mai_mai_n42_), .B0(mai_mai_n398_), .Y(mai_mai_n903_));
  OAI220     m0881(.A0(mai_mai_n903_), .A1(mai_mai_n860_), .B0(mai_mai_n902_), .B1(mai_mai_n901_), .Y(mai_mai_n904_));
  NO3        m0882(.A(mai_mai_n904_), .B(mai_mai_n898_), .C(mai_mai_n895_), .Y(mai_mai_n905_));
  NA2        m0883(.A(mai_mai_n652_), .B(mai_mai_n126_), .Y(mai_mai_n906_));
  NO2        m0884(.A(i_6_), .B(mai_mai_n906_), .Y(mai_mai_n907_));
  NA2        m0885(.A(mai_mai_n175_), .B(mai_mai_n107_), .Y(mai_mai_n908_));
  INV        m0886(.A(mai_mai_n907_), .Y(mai_mai_n909_));
  NOi21      m0887(.An(i_7_), .B(i_5_), .Y(mai_mai_n910_));
  NOi31      m0888(.An(mai_mai_n910_), .B(i_0_), .C(mai_mai_n721_), .Y(mai_mai_n911_));
  NA3        m0889(.A(mai_mai_n911_), .B(mai_mai_n379_), .C(i_6_), .Y(mai_mai_n912_));
  BUFFER     m0890(.A(mai_mai_n912_), .Y(mai_mai_n913_));
  NO3        m0891(.A(mai_mai_n393_), .B(mai_mai_n358_), .C(mai_mai_n354_), .Y(mai_mai_n914_));
  NO2        m0892(.A(mai_mai_n267_), .B(mai_mai_n312_), .Y(mai_mai_n915_));
  NO2        m0893(.A(mai_mai_n721_), .B(mai_mai_n262_), .Y(mai_mai_n916_));
  AOI210     m0894(.A0(mai_mai_n916_), .A1(mai_mai_n915_), .B0(mai_mai_n914_), .Y(mai_mai_n917_));
  NA4        m0895(.A(mai_mai_n917_), .B(mai_mai_n913_), .C(mai_mai_n909_), .D(mai_mai_n905_), .Y(mai_mai_n918_));
  NO2        m0896(.A(mai_mai_n868_), .B(mai_mai_n243_), .Y(mai_mai_n919_));
  AN2        m0897(.A(mai_mai_n324_), .B(mai_mai_n322_), .Y(mai_mai_n920_));
  AN2        m0898(.A(mai_mai_n920_), .B(mai_mai_n864_), .Y(mai_mai_n921_));
  OAI210     m0899(.A0(mai_mai_n921_), .A1(mai_mai_n919_), .B0(i_10_), .Y(mai_mai_n922_));
  OA210      m0900(.A0(mai_mai_n465_), .A1(mai_mai_n229_), .B0(mai_mai_n464_), .Y(mai_mai_n923_));
  NO2        m0901(.A(mai_mai_n260_), .B(mai_mai_n47_), .Y(mai_mai_n924_));
  NA2        m0902(.A(mai_mai_n899_), .B(mai_mai_n301_), .Y(mai_mai_n925_));
  OAI210     m0903(.A0(mai_mai_n924_), .A1(mai_mai_n189_), .B0(mai_mai_n925_), .Y(mai_mai_n926_));
  NA2        m0904(.A(mai_mai_n926_), .B(mai_mai_n465_), .Y(mai_mai_n927_));
  NA2        m0905(.A(mai_mai_n96_), .B(mai_mai_n45_), .Y(mai_mai_n928_));
  NO2        m0906(.A(mai_mai_n76_), .B(mai_mai_n745_), .Y(mai_mai_n929_));
  AOI220     m0907(.A0(mai_mai_n929_), .A1(mai_mai_n928_), .B0(mai_mai_n178_), .B1(mai_mai_n590_), .Y(mai_mai_n930_));
  NO2        m0908(.A(mai_mai_n930_), .B(mai_mai_n48_), .Y(mai_mai_n931_));
  NO3        m0909(.A(mai_mai_n582_), .B(mai_mai_n353_), .C(mai_mai_n24_), .Y(mai_mai_n932_));
  AOI210     m0910(.A0(mai_mai_n694_), .A1(mai_mai_n541_), .B0(mai_mai_n932_), .Y(mai_mai_n933_));
  NAi21      m0911(.An(i_9_), .B(i_5_), .Y(mai_mai_n934_));
  NO2        m0912(.A(mai_mai_n934_), .B(mai_mai_n393_), .Y(mai_mai_n935_));
  NO2        m0913(.A(mai_mai_n593_), .B(mai_mai_n109_), .Y(mai_mai_n936_));
  AOI220     m0914(.A0(mai_mai_n936_), .A1(i_0_), .B0(mai_mai_n935_), .B1(mai_mai_n616_), .Y(mai_mai_n937_));
  OAI220     m0915(.A0(mai_mai_n937_), .A1(mai_mai_n87_), .B0(mai_mai_n933_), .B1(mai_mai_n176_), .Y(mai_mai_n938_));
  NO3        m0916(.A(mai_mai_n938_), .B(mai_mai_n931_), .C(mai_mai_n514_), .Y(mai_mai_n939_));
  NA3        m0917(.A(mai_mai_n939_), .B(mai_mai_n927_), .C(mai_mai_n922_), .Y(mai_mai_n940_));
  NO3        m0918(.A(mai_mai_n940_), .B(mai_mai_n918_), .C(mai_mai_n891_), .Y(mai_mai_n941_));
  NO2        m0919(.A(i_0_), .B(mai_mai_n721_), .Y(mai_mai_n942_));
  NA2        m0920(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n943_));
  INV        m0921(.A(mai_mai_n943_), .Y(mai_mai_n944_));
  NO3        m0922(.A(mai_mai_n109_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n945_));
  AO220      m0923(.A0(mai_mai_n945_), .A1(mai_mai_n944_), .B0(mai_mai_n942_), .B1(mai_mai_n178_), .Y(mai_mai_n946_));
  AOI210     m0924(.A0(mai_mai_n795_), .A1(mai_mai_n681_), .B0(mai_mai_n908_), .Y(mai_mai_n947_));
  AOI210     m0925(.A0(mai_mai_n946_), .A1(mai_mai_n342_), .B0(mai_mai_n947_), .Y(mai_mai_n948_));
  NA2        m0926(.A(mai_mai_n731_), .B(mai_mai_n151_), .Y(mai_mai_n949_));
  INV        m0927(.A(mai_mai_n949_), .Y(mai_mai_n950_));
  NA3        m0928(.A(mai_mai_n950_), .B(mai_mai_n668_), .C(mai_mai_n74_), .Y(mai_mai_n951_));
  NO2        m0929(.A(mai_mai_n813_), .B(mai_mai_n393_), .Y(mai_mai_n952_));
  NA3        m0930(.A(mai_mai_n841_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n953_));
  NA2        m0931(.A(mai_mai_n842_), .B(i_9_), .Y(mai_mai_n954_));
  NO2        m0932(.A(mai_mai_n953_), .B(mai_mai_n954_), .Y(mai_mai_n955_));
  OAI210     m0933(.A0(mai_mai_n247_), .A1(i_9_), .B0(mai_mai_n233_), .Y(mai_mai_n956_));
  AOI210     m0934(.A0(mai_mai_n956_), .A1(mai_mai_n874_), .B0(mai_mai_n159_), .Y(mai_mai_n957_));
  NO3        m0935(.A(mai_mai_n957_), .B(mai_mai_n955_), .C(mai_mai_n952_), .Y(mai_mai_n958_));
  NA3        m0936(.A(mai_mai_n958_), .B(mai_mai_n951_), .C(mai_mai_n948_), .Y(mai_mai_n959_));
  NA2        m0937(.A(mai_mai_n920_), .B(mai_mai_n368_), .Y(mai_mai_n960_));
  AOI210     m0938(.A0(mai_mai_n295_), .A1(mai_mai_n168_), .B0(mai_mai_n960_), .Y(mai_mai_n961_));
  NA3        m0939(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n962_));
  NA2        m0940(.A(mai_mai_n896_), .B(mai_mai_n481_), .Y(mai_mai_n963_));
  AOI210     m0941(.A0(mai_mai_n962_), .A1(mai_mai_n168_), .B0(mai_mai_n963_), .Y(mai_mai_n964_));
  NO2        m0942(.A(mai_mai_n964_), .B(mai_mai_n961_), .Y(mai_mai_n965_));
  NO3        m0943(.A(mai_mai_n882_), .B(mai_mai_n859_), .C(mai_mai_n192_), .Y(mai_mai_n966_));
  AOI220     m0944(.A0(mai_mai_n966_), .A1(i_11_), .B0(mai_mai_n565_), .B1(mai_mai_n76_), .Y(mai_mai_n967_));
  NO3        m0945(.A(mai_mai_n214_), .B(mai_mai_n378_), .C(i_0_), .Y(mai_mai_n968_));
  OAI210     m0946(.A0(mai_mai_n968_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n969_));
  INV        m0947(.A(mai_mai_n223_), .Y(mai_mai_n970_));
  OAI220     m0948(.A0(mai_mai_n525_), .A1(mai_mai_n144_), .B0(mai_mai_n638_), .B1(mai_mai_n610_), .Y(mai_mai_n971_));
  NA3        m0949(.A(mai_mai_n971_), .B(mai_mai_n386_), .C(mai_mai_n970_), .Y(mai_mai_n972_));
  NA4        m0950(.A(mai_mai_n972_), .B(mai_mai_n969_), .C(mai_mai_n967_), .D(mai_mai_n965_), .Y(mai_mai_n973_));
  NO2        m0951(.A(mai_mai_n246_), .B(mai_mai_n96_), .Y(mai_mai_n974_));
  AOI210     m0952(.A0(mai_mai_n974_), .A1(mai_mai_n942_), .B0(mai_mai_n113_), .Y(mai_mai_n975_));
  AOI220     m0953(.A0(mai_mai_n910_), .A1(mai_mai_n481_), .B0(mai_mai_n841_), .B1(mai_mai_n169_), .Y(mai_mai_n976_));
  NA2        m0954(.A(mai_mai_n345_), .B(mai_mai_n180_), .Y(mai_mai_n977_));
  OA220      m0955(.A0(mai_mai_n977_), .A1(mai_mai_n976_), .B0(mai_mai_n975_), .B1(i_5_), .Y(mai_mai_n978_));
  AOI210     m0956(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n179_), .Y(mai_mai_n979_));
  NA2        m0957(.A(mai_mai_n979_), .B(mai_mai_n923_), .Y(mai_mai_n980_));
  NA3        m0958(.A(mai_mai_n607_), .B(mai_mai_n187_), .C(mai_mai_n85_), .Y(mai_mai_n981_));
  NA2        m0959(.A(mai_mai_n981_), .B(mai_mai_n539_), .Y(mai_mai_n982_));
  NO3        m0960(.A(mai_mai_n851_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n983_));
  NA3        m0961(.A(mai_mai_n486_), .B(mai_mai_n479_), .C(mai_mai_n462_), .Y(mai_mai_n984_));
  NO3        m0962(.A(mai_mai_n984_), .B(mai_mai_n983_), .C(mai_mai_n982_), .Y(mai_mai_n985_));
  NA3        m0963(.A(mai_mai_n383_), .B(mai_mai_n175_), .C(mai_mai_n174_), .Y(mai_mai_n986_));
  NA3        m0964(.A(mai_mai_n896_), .B(mai_mai_n289_), .C(mai_mai_n233_), .Y(mai_mai_n987_));
  NA2        m0965(.A(mai_mai_n987_), .B(mai_mai_n986_), .Y(mai_mai_n988_));
  NO3        m0966(.A(mai_mai_n893_), .B(mai_mai_n223_), .C(mai_mai_n192_), .Y(mai_mai_n989_));
  NO2        m0967(.A(mai_mai_n989_), .B(mai_mai_n988_), .Y(mai_mai_n990_));
  NA4        m0968(.A(mai_mai_n990_), .B(mai_mai_n985_), .C(mai_mai_n980_), .D(mai_mai_n978_), .Y(mai_mai_n991_));
  INV        m0969(.A(mai_mai_n609_), .Y(mai_mai_n992_));
  NO3        m0970(.A(mai_mai_n992_), .B(mai_mai_n555_), .C(mai_mai_n339_), .Y(mai_mai_n993_));
  NO2        m0971(.A(mai_mai_n87_), .B(i_5_), .Y(mai_mai_n994_));
  NA3        m0972(.A(mai_mai_n842_), .B(mai_mai_n114_), .C(mai_mai_n129_), .Y(mai_mai_n995_));
  INV        m0973(.A(mai_mai_n995_), .Y(mai_mai_n996_));
  AOI210     m0974(.A0(mai_mai_n996_), .A1(mai_mai_n994_), .B0(mai_mai_n993_), .Y(mai_mai_n997_));
  NA3        m0975(.A(mai_mai_n301_), .B(i_5_), .C(mai_mai_n195_), .Y(mai_mai_n998_));
  NAi31      m0976(.An(mai_mai_n245_), .B(mai_mai_n998_), .C(mai_mai_n246_), .Y(mai_mai_n999_));
  NO4        m0977(.A(mai_mai_n243_), .B(mai_mai_n214_), .C(i_0_), .D(i_12_), .Y(mai_mai_n1000_));
  AOI220     m0978(.A0(mai_mai_n1000_), .A1(mai_mai_n999_), .B0(mai_mai_n789_), .B1(mai_mai_n180_), .Y(mai_mai_n1001_));
  NA2        m0979(.A(mai_mai_n910_), .B(mai_mai_n461_), .Y(mai_mai_n1002_));
  NA2        m0980(.A(mai_mai_n65_), .B(mai_mai_n105_), .Y(mai_mai_n1003_));
  OAI220     m0981(.A0(mai_mai_n1003_), .A1(mai_mai_n998_), .B0(mai_mai_n1002_), .B1(mai_mai_n669_), .Y(mai_mai_n1004_));
  NA2        m0982(.A(mai_mai_n1004_), .B(mai_mai_n900_), .Y(mai_mai_n1005_));
  NA3        m0983(.A(mai_mai_n1005_), .B(mai_mai_n1001_), .C(mai_mai_n997_), .Y(mai_mai_n1006_));
  NO4        m0984(.A(mai_mai_n1006_), .B(mai_mai_n991_), .C(mai_mai_n973_), .D(mai_mai_n959_), .Y(mai_mai_n1007_));
  OAI210     m0985(.A0(mai_mai_n816_), .A1(mai_mai_n809_), .B0(mai_mai_n37_), .Y(mai_mai_n1008_));
  NA2        m0986(.A(mai_mai_n1008_), .B(mai_mai_n605_), .Y(mai_mai_n1009_));
  NA2        m0987(.A(mai_mai_n1009_), .B(mai_mai_n210_), .Y(mai_mai_n1010_));
  OAI210     m0988(.A0(mai_mai_n609_), .A1(mai_mai_n607_), .B0(mai_mai_n311_), .Y(mai_mai_n1011_));
  NAi31      m0989(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n1012_));
  AOI210     m0990(.A0(mai_mai_n122_), .A1(mai_mai_n71_), .B0(mai_mai_n1012_), .Y(mai_mai_n1013_));
  INV        m0991(.A(mai_mai_n1013_), .Y(mai_mai_n1014_));
  NA2        m0992(.A(mai_mai_n1014_), .B(mai_mai_n1011_), .Y(mai_mai_n1015_));
  NO2        m0993(.A(mai_mai_n452_), .B(mai_mai_n273_), .Y(mai_mai_n1016_));
  NO4        m0994(.A(mai_mai_n236_), .B(mai_mai_n150_), .C(mai_mai_n672_), .D(mai_mai_n37_), .Y(mai_mai_n1017_));
  NO3        m0995(.A(mai_mai_n1017_), .B(mai_mai_n1016_), .C(mai_mai_n876_), .Y(mai_mai_n1018_));
  INV        m0996(.A(mai_mai_n1018_), .Y(mai_mai_n1019_));
  AOI210     m0997(.A0(mai_mai_n1015_), .A1(mai_mai_n49_), .B0(mai_mai_n1019_), .Y(mai_mai_n1020_));
  AOI210     m0998(.A0(mai_mai_n1020_), .A1(mai_mai_n1010_), .B0(mai_mai_n74_), .Y(mai_mai_n1021_));
  NO2        m0999(.A(mai_mai_n562_), .B(mai_mai_n375_), .Y(mai_mai_n1022_));
  NO2        m1000(.A(mai_mai_n1022_), .B(mai_mai_n751_), .Y(mai_mai_n1023_));
  AOI210     m1001(.A0(mai_mai_n979_), .A1(mai_mai_n896_), .B0(mai_mai_n911_), .Y(mai_mai_n1024_));
  NO2        m1002(.A(mai_mai_n1024_), .B(mai_mai_n672_), .Y(mai_mai_n1025_));
  NA2        m1003(.A(mai_mai_n267_), .B(mai_mai_n58_), .Y(mai_mai_n1026_));
  AOI220     m1004(.A0(mai_mai_n1026_), .A1(mai_mai_n77_), .B0(mai_mai_n340_), .B1(mai_mai_n259_), .Y(mai_mai_n1027_));
  NO2        m1005(.A(mai_mai_n1027_), .B(mai_mai_n240_), .Y(mai_mai_n1028_));
  NA3        m1006(.A(mai_mai_n100_), .B(mai_mai_n303_), .C(mai_mai_n31_), .Y(mai_mai_n1029_));
  INV        m1007(.A(mai_mai_n1029_), .Y(mai_mai_n1030_));
  NO3        m1008(.A(mai_mai_n1030_), .B(mai_mai_n1028_), .C(mai_mai_n1025_), .Y(mai_mai_n1031_));
  OAI210     m1009(.A0(mai_mai_n275_), .A1(mai_mai_n164_), .B0(mai_mai_n90_), .Y(mai_mai_n1032_));
  NA3        m1010(.A(mai_mai_n755_), .B(mai_mai_n289_), .C(mai_mai_n81_), .Y(mai_mai_n1033_));
  AOI210     m1011(.A0(mai_mai_n1033_), .A1(mai_mai_n1032_), .B0(i_11_), .Y(mai_mai_n1034_));
  NO3        m1012(.A(mai_mai_n60_), .B(mai_mai_n59_), .C(i_4_), .Y(mai_mai_n1035_));
  OAI210     m1013(.A0(mai_mai_n915_), .A1(mai_mai_n303_), .B0(mai_mai_n1035_), .Y(mai_mai_n1036_));
  NO2        m1014(.A(mai_mai_n1036_), .B(mai_mai_n721_), .Y(mai_mai_n1037_));
  NO4        m1015(.A(mai_mai_n934_), .B(mai_mai_n469_), .C(mai_mai_n256_), .D(mai_mai_n255_), .Y(mai_mai_n1038_));
  NO2        m1016(.A(mai_mai_n1038_), .B(mai_mai_n559_), .Y(mai_mai_n1039_));
  INV        m1017(.A(mai_mai_n359_), .Y(mai_mai_n1040_));
  AOI210     m1018(.A0(mai_mai_n1040_), .A1(mai_mai_n1039_), .B0(mai_mai_n41_), .Y(mai_mai_n1041_));
  NO3        m1019(.A(mai_mai_n1041_), .B(mai_mai_n1037_), .C(mai_mai_n1034_), .Y(mai_mai_n1042_));
  OAI210     m1020(.A0(mai_mai_n1031_), .A1(i_4_), .B0(mai_mai_n1042_), .Y(mai_mai_n1043_));
  NO3        m1021(.A(mai_mai_n1043_), .B(mai_mai_n1023_), .C(mai_mai_n1021_), .Y(mai_mai_n1044_));
  NA4        m1022(.A(mai_mai_n1044_), .B(mai_mai_n1007_), .C(mai_mai_n941_), .D(mai_mai_n867_), .Y(mai4));
  INV        m1023(.A(mai_mai_n693_), .Y(mai_mai_n1048_));
  INV        m1024(.A(mai_mai_n476_), .Y(mai_mai_n1049_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u0033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  NA2        u0034(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n57_));
  NA3        u0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n58_));
  NO2        u0036(.A(i_1_), .B(i_6_), .Y(men_men_n59_));
  NA2        u0037(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  OAI210     u0038(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n58_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_12_), .Y(men_men_n62_));
  NAi21      u0040(.An(i_2_), .B(i_7_), .Y(men_men_n63_));
  INV        u0041(.A(i_1_), .Y(men_men_n64_));
  NA2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NA3        u0043(.A(men_men_n65_), .B(men_men_n63_), .C(men_men_n31_), .Y(men_men_n66_));
  NA2        u0044(.A(i_1_), .B(i_10_), .Y(men_men_n67_));
  NO2        u0045(.A(men_men_n67_), .B(i_6_), .Y(men_men_n68_));
  NAi31      u0046(.An(men_men_n68_), .B(men_men_n66_), .C(men_men_n62_), .Y(men_men_n69_));
  NA2        u0047(.A(men_men_n51_), .B(i_2_), .Y(men_men_n70_));
  AOI210     u0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n71_));
  NA2        u0049(.A(i_1_), .B(i_6_), .Y(men_men_n72_));
  NO2        u0050(.A(men_men_n72_), .B(men_men_n25_), .Y(men_men_n73_));
  INV        u0051(.A(i_0_), .Y(men_men_n74_));
  NAi21      u0052(.An(i_5_), .B(i_10_), .Y(men_men_n75_));
  NA2        u0053(.A(i_5_), .B(i_9_), .Y(men_men_n76_));
  AOI210     u0054(.A0(men_men_n76_), .A1(men_men_n75_), .B0(men_men_n74_), .Y(men_men_n77_));
  NO2        u0055(.A(men_men_n77_), .B(men_men_n73_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n78_), .Y(men_men_n79_));
  OAI210     u0057(.A0(men_men_n79_), .A1(men_men_n69_), .B0(i_0_), .Y(men_men_n80_));
  NA2        u0058(.A(i_12_), .B(i_5_), .Y(men_men_n81_));
  NA2        u0059(.A(i_2_), .B(i_8_), .Y(men_men_n82_));
  NO2        u0060(.A(men_men_n82_), .B(men_men_n59_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_9_), .Y(men_men_n84_));
  NO2        u0062(.A(i_3_), .B(i_7_), .Y(men_men_n85_));
  NO3        u0063(.A(men_men_n85_), .B(men_men_n84_), .C(men_men_n64_), .Y(men_men_n86_));
  INV        u0064(.A(i_6_), .Y(men_men_n87_));
  NO2        u0065(.A(i_2_), .B(i_7_), .Y(men_men_n88_));
  INV        u0066(.A(men_men_n88_), .Y(men_men_n89_));
  OAI210     u0067(.A0(men_men_n86_), .A1(men_men_n83_), .B0(men_men_n89_), .Y(men_men_n90_));
  NAi21      u0068(.An(i_6_), .B(i_10_), .Y(men_men_n91_));
  NA2        u0069(.A(i_6_), .B(i_9_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n64_), .Y(men_men_n93_));
  NA2        u0071(.A(i_2_), .B(i_6_), .Y(men_men_n94_));
  NO3        u0072(.A(men_men_n94_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n95_));
  NO2        u0073(.A(men_men_n95_), .B(men_men_n93_), .Y(men_men_n96_));
  AOI210     u0074(.A0(men_men_n96_), .A1(men_men_n90_), .B0(men_men_n81_), .Y(men_men_n97_));
  AN3        u0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n98_));
  NAi21      u0076(.An(i_6_), .B(i_11_), .Y(men_men_n99_));
  NO2        u0077(.A(i_5_), .B(i_8_), .Y(men_men_n100_));
  NOi21      u0078(.An(men_men_n100_), .B(men_men_n99_), .Y(men_men_n101_));
  AOI220     u0079(.A0(men_men_n101_), .A1(men_men_n63_), .B0(men_men_n98_), .B1(men_men_n32_), .Y(men_men_n102_));
  INV        u0080(.A(i_7_), .Y(men_men_n103_));
  NA2        u0081(.A(men_men_n47_), .B(men_men_n103_), .Y(men_men_n104_));
  NO2        u0082(.A(i_0_), .B(i_5_), .Y(men_men_n105_));
  NO2        u0083(.A(men_men_n105_), .B(men_men_n87_), .Y(men_men_n106_));
  NA2        u0084(.A(i_12_), .B(i_3_), .Y(men_men_n107_));
  INV        u0085(.A(men_men_n107_), .Y(men_men_n108_));
  NA3        u0086(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n104_), .Y(men_men_n109_));
  NAi21      u0087(.An(i_7_), .B(i_11_), .Y(men_men_n110_));
  NO3        u0088(.A(men_men_n110_), .B(men_men_n91_), .C(men_men_n54_), .Y(men_men_n111_));
  AN2        u0089(.A(i_2_), .B(i_10_), .Y(men_men_n112_));
  NO2        u0090(.A(men_men_n112_), .B(i_7_), .Y(men_men_n113_));
  OR2        u0091(.A(men_men_n81_), .B(men_men_n59_), .Y(men_men_n114_));
  NO2        u0092(.A(i_8_), .B(men_men_n103_), .Y(men_men_n115_));
  NO3        u0093(.A(men_men_n115_), .B(men_men_n114_), .C(men_men_n113_), .Y(men_men_n116_));
  NA2        u0094(.A(i_12_), .B(i_7_), .Y(men_men_n117_));
  NO2        u0095(.A(men_men_n64_), .B(men_men_n26_), .Y(men_men_n118_));
  NA2        u0096(.A(i_11_), .B(i_12_), .Y(men_men_n119_));
  NO2        u0097(.A(men_men_n1093_), .B(men_men_n116_), .Y(men_men_n120_));
  NAi41      u0098(.An(men_men_n111_), .B(men_men_n120_), .C(men_men_n109_), .D(men_men_n102_), .Y(men_men_n121_));
  NOi21      u0099(.An(i_1_), .B(i_5_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n122_), .B(i_11_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n124_));
  NA2        u0102(.A(i_7_), .B(men_men_n25_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n126_));
  NO2        u0104(.A(men_men_n126_), .B(men_men_n47_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n128_));
  NAi21      u0106(.An(i_3_), .B(i_8_), .Y(men_men_n129_));
  NA2        u0107(.A(men_men_n129_), .B(men_men_n63_), .Y(men_men_n130_));
  NOi31      u0108(.An(men_men_n130_), .B(men_men_n128_), .C(men_men_n127_), .Y(men_men_n131_));
  NO2        u0109(.A(i_1_), .B(men_men_n87_), .Y(men_men_n132_));
  NO2        u0110(.A(i_6_), .B(i_5_), .Y(men_men_n133_));
  NA2        u0111(.A(men_men_n133_), .B(i_3_), .Y(men_men_n134_));
  AO210      u0112(.A0(men_men_n134_), .A1(men_men_n48_), .B0(men_men_n132_), .Y(men_men_n135_));
  OAI220     u0113(.A0(men_men_n135_), .A1(men_men_n110_), .B0(men_men_n131_), .B1(men_men_n123_), .Y(men_men_n136_));
  NO3        u0114(.A(men_men_n136_), .B(men_men_n121_), .C(men_men_n97_), .Y(men_men_n137_));
  NA3        u0115(.A(men_men_n137_), .B(men_men_n80_), .C(men_men_n57_), .Y(men2));
  NO2        u0116(.A(men_men_n64_), .B(men_men_n37_), .Y(men_men_n139_));
  NA2        u0117(.A(i_6_), .B(men_men_n25_), .Y(men_men_n140_));
  NA2        u0118(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n141_));
  NA4        u0119(.A(men_men_n141_), .B(men_men_n78_), .C(men_men_n70_), .D(men_men_n30_), .Y(men0));
  AN2        u0120(.A(i_8_), .B(i_7_), .Y(men_men_n143_));
  NA2        u0121(.A(men_men_n143_), .B(i_6_), .Y(men_men_n144_));
  NO2        u0122(.A(i_12_), .B(i_13_), .Y(men_men_n145_));
  NAi21      u0123(.An(i_5_), .B(i_11_), .Y(men_men_n146_));
  NOi21      u0124(.An(men_men_n145_), .B(men_men_n146_), .Y(men_men_n147_));
  NO2        u0125(.A(i_0_), .B(i_1_), .Y(men_men_n148_));
  NA2        u0126(.A(i_2_), .B(i_3_), .Y(men_men_n149_));
  NO2        u0127(.A(men_men_n149_), .B(i_4_), .Y(men_men_n150_));
  NA3        u0128(.A(men_men_n150_), .B(men_men_n148_), .C(men_men_n147_), .Y(men_men_n151_));
  AN2        u0129(.A(men_men_n145_), .B(men_men_n84_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n152_), .B(men_men_n27_), .Y(men_men_n153_));
  NA2        u0131(.A(i_1_), .B(i_5_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n74_), .B(men_men_n47_), .Y(men_men_n155_));
  NA2        u0133(.A(men_men_n155_), .B(men_men_n36_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n156_), .B(men_men_n154_), .C(men_men_n153_), .Y(men_men_n157_));
  OR2        u0135(.A(i_0_), .B(i_1_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n81_), .C(i_13_), .Y(men_men_n159_));
  NAi32      u0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n160_));
  NAi21      u0138(.An(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0139(.An(i_4_), .B(i_10_), .Y(men_men_n162_));
  NA2        u0140(.A(men_men_n162_), .B(men_men_n40_), .Y(men_men_n163_));
  NO2        u0141(.A(i_3_), .B(i_5_), .Y(men_men_n164_));
  NO3        u0142(.A(men_men_n74_), .B(i_2_), .C(i_1_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  OAI210     u0144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n167_));
  NO2        u0145(.A(men_men_n167_), .B(men_men_n157_), .Y(men_men_n168_));
  AOI210     u0146(.A0(men_men_n168_), .A1(men_men_n151_), .B0(men_men_n144_), .Y(men_men_n169_));
  NA3        u0147(.A(men_men_n74_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n170_));
  NA2        u0148(.A(i_3_), .B(men_men_n49_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_4_), .B(i_9_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_11_), .B(i_13_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OR2        u0152(.A(men_men_n174_), .B(men_men_n171_), .Y(men_men_n175_));
  NO2        u0153(.A(i_4_), .B(i_5_), .Y(men_men_n176_));
  NAi21      u0154(.An(i_12_), .B(i_11_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n177_), .B(i_13_), .Y(men_men_n178_));
  NA3        u0156(.A(men_men_n178_), .B(men_men_n176_), .C(men_men_n84_), .Y(men_men_n179_));
  AOI210     u0157(.A0(men_men_n179_), .A1(men_men_n175_), .B0(men_men_n170_), .Y(men_men_n180_));
  NO2        u0158(.A(men_men_n74_), .B(men_men_n64_), .Y(men_men_n181_));
  NA2        u0159(.A(men_men_n181_), .B(men_men_n47_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n36_), .B(i_5_), .Y(men_men_n183_));
  NAi31      u0161(.An(men_men_n183_), .B(men_men_n152_), .C(i_11_), .Y(men_men_n184_));
  NA2        u0162(.A(i_3_), .B(i_5_), .Y(men_men_n185_));
  OR2        u0163(.A(men_men_n185_), .B(men_men_n174_), .Y(men_men_n186_));
  AOI210     u0164(.A0(men_men_n186_), .A1(men_men_n184_), .B0(men_men_n182_), .Y(men_men_n187_));
  NO2        u0165(.A(men_men_n74_), .B(i_5_), .Y(men_men_n188_));
  NO2        u0166(.A(i_13_), .B(i_10_), .Y(men_men_n189_));
  NA3        u0167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n45_), .Y(men_men_n190_));
  NO2        u0168(.A(i_2_), .B(i_1_), .Y(men_men_n191_));
  NA2        u0169(.A(men_men_n191_), .B(i_3_), .Y(men_men_n192_));
  NAi21      u0170(.An(i_4_), .B(i_12_), .Y(men_men_n193_));
  NO4        u0171(.A(men_men_n193_), .B(men_men_n192_), .C(men_men_n190_), .D(men_men_n25_), .Y(men_men_n194_));
  NO3        u0172(.A(men_men_n194_), .B(men_men_n187_), .C(men_men_n180_), .Y(men_men_n195_));
  INV        u0173(.A(i_8_), .Y(men_men_n196_));
  NO2        u0174(.A(men_men_n196_), .B(i_7_), .Y(men_men_n197_));
  NA2        u0175(.A(men_men_n197_), .B(i_6_), .Y(men_men_n198_));
  NO3        u0176(.A(i_3_), .B(men_men_n87_), .C(men_men_n49_), .Y(men_men_n199_));
  NA2        u0177(.A(men_men_n199_), .B(men_men_n115_), .Y(men_men_n200_));
  NO3        u0178(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n201_));
  NA3        u0179(.A(men_men_n201_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n202_));
  NO3        u0180(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n203_));
  OAI210     u0181(.A0(men_men_n98_), .A1(i_12_), .B0(men_men_n203_), .Y(men_men_n204_));
  AOI210     u0182(.A0(men_men_n204_), .A1(men_men_n202_), .B0(men_men_n200_), .Y(men_men_n205_));
  NO2        u0183(.A(i_3_), .B(i_8_), .Y(men_men_n206_));
  NO3        u0184(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n207_));
  NO2        u0185(.A(men_men_n105_), .B(men_men_n59_), .Y(men_men_n208_));
  NO2        u0186(.A(i_13_), .B(i_9_), .Y(men_men_n209_));
  NA3        u0187(.A(men_men_n209_), .B(i_6_), .C(men_men_n196_), .Y(men_men_n210_));
  NAi21      u0188(.An(i_12_), .B(i_3_), .Y(men_men_n211_));
  NO2        u0189(.A(men_men_n45_), .B(i_5_), .Y(men_men_n212_));
  NO3        u0190(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n213_));
  NA3        u0191(.A(men_men_n213_), .B(men_men_n212_), .C(i_10_), .Y(men_men_n214_));
  NO2        u0192(.A(men_men_n214_), .B(men_men_n210_), .Y(men_men_n215_));
  AOI210     u0193(.A0(men_men_n215_), .A1(i_7_), .B0(men_men_n205_), .Y(men_men_n216_));
  OAI220     u0194(.A0(men_men_n216_), .A1(i_4_), .B0(men_men_n198_), .B1(men_men_n195_), .Y(men_men_n217_));
  NAi21      u0195(.An(i_12_), .B(i_7_), .Y(men_men_n218_));
  NA3        u0196(.A(i_13_), .B(men_men_n196_), .C(i_10_), .Y(men_men_n219_));
  NO2        u0197(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n220_));
  NA2        u0198(.A(i_0_), .B(i_5_), .Y(men_men_n221_));
  NA2        u0199(.A(men_men_n221_), .B(men_men_n106_), .Y(men_men_n222_));
  OAI220     u0200(.A0(men_men_n222_), .A1(men_men_n192_), .B0(men_men_n182_), .B1(men_men_n134_), .Y(men_men_n223_));
  NAi31      u0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n224_));
  NO2        u0202(.A(men_men_n36_), .B(i_13_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n74_), .B(men_men_n26_), .Y(men_men_n226_));
  NO2        u0204(.A(men_men_n47_), .B(men_men_n64_), .Y(men_men_n227_));
  NA3        u0205(.A(men_men_n227_), .B(men_men_n226_), .C(men_men_n225_), .Y(men_men_n228_));
  INV        u0206(.A(i_13_), .Y(men_men_n229_));
  NO2        u0207(.A(i_12_), .B(men_men_n229_), .Y(men_men_n230_));
  NA3        u0208(.A(men_men_n230_), .B(men_men_n201_), .C(men_men_n199_), .Y(men_men_n231_));
  OAI210     u0209(.A0(men_men_n228_), .A1(men_men_n224_), .B0(men_men_n231_), .Y(men_men_n232_));
  AOI220     u0210(.A0(men_men_n232_), .A1(men_men_n143_), .B0(men_men_n223_), .B1(men_men_n220_), .Y(men_men_n233_));
  NO2        u0211(.A(i_12_), .B(men_men_n37_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n185_), .B(i_4_), .Y(men_men_n235_));
  NA2        u0213(.A(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  OR2        u0214(.A(i_8_), .B(i_7_), .Y(men_men_n237_));
  NO2        u0215(.A(men_men_n237_), .B(men_men_n87_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n54_), .B(i_1_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  INV        u0218(.A(i_12_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n45_), .B(men_men_n241_), .Y(men_men_n242_));
  NO3        u0220(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n243_));
  NA2        u0221(.A(i_2_), .B(i_1_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n240_), .B(men_men_n236_), .Y(men_men_n245_));
  NO3        u0223(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n246_));
  NAi21      u0224(.An(i_4_), .B(i_3_), .Y(men_men_n247_));
  NO2        u0225(.A(men_men_n247_), .B(men_men_n76_), .Y(men_men_n248_));
  NO2        u0226(.A(i_0_), .B(i_6_), .Y(men_men_n249_));
  NOi41      u0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n250_));
  NA2        u0228(.A(men_men_n250_), .B(men_men_n249_), .Y(men_men_n251_));
  NO2        u0229(.A(men_men_n244_), .B(men_men_n185_), .Y(men_men_n252_));
  NAi21      u0230(.An(men_men_n251_), .B(men_men_n252_), .Y(men_men_n253_));
  INV        u0231(.A(men_men_n253_), .Y(men_men_n254_));
  AOI220     u0232(.A0(men_men_n254_), .A1(men_men_n40_), .B0(men_men_n245_), .B1(men_men_n209_), .Y(men_men_n255_));
  NO2        u0233(.A(i_11_), .B(men_men_n229_), .Y(men_men_n256_));
  NOi21      u0234(.An(i_1_), .B(i_6_), .Y(men_men_n257_));
  NAi21      u0235(.An(i_3_), .B(i_7_), .Y(men_men_n258_));
  NA2        u0236(.A(men_men_n241_), .B(i_9_), .Y(men_men_n259_));
  OR4        u0237(.A(men_men_n259_), .B(men_men_n258_), .C(men_men_n257_), .D(men_men_n188_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n261_));
  NO2        u0239(.A(i_12_), .B(i_3_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n74_), .B(i_5_), .Y(men_men_n263_));
  NA2        u0241(.A(i_3_), .B(i_9_), .Y(men_men_n264_));
  NAi21      u0242(.An(i_7_), .B(i_10_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA3        u0244(.A(men_men_n266_), .B(men_men_n263_), .C(men_men_n65_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n267_), .B(men_men_n260_), .Y(men_men_n268_));
  NA3        u0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n269_));
  INV        u0247(.A(men_men_n144_), .Y(men_men_n270_));
  NA2        u0248(.A(men_men_n241_), .B(i_13_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n271_), .B(men_men_n76_), .Y(men_men_n272_));
  AOI220     u0250(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n268_), .B1(men_men_n256_), .Y(men_men_n273_));
  NO2        u0251(.A(men_men_n237_), .B(men_men_n37_), .Y(men_men_n274_));
  NA2        u0252(.A(i_12_), .B(i_6_), .Y(men_men_n275_));
  OR2        u0253(.A(i_13_), .B(i_9_), .Y(men_men_n276_));
  NO3        u0254(.A(men_men_n276_), .B(men_men_n275_), .C(men_men_n49_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n247_), .B(i_2_), .Y(men_men_n278_));
  NA2        u0256(.A(men_men_n256_), .B(i_9_), .Y(men_men_n279_));
  NA2        u0257(.A(men_men_n155_), .B(men_men_n64_), .Y(men_men_n280_));
  NO3        u0258(.A(i_11_), .B(men_men_n229_), .C(men_men_n25_), .Y(men_men_n281_));
  NO2        u0259(.A(men_men_n258_), .B(i_8_), .Y(men_men_n282_));
  NO2        u0260(.A(i_6_), .B(men_men_n49_), .Y(men_men_n283_));
  NA3        u0261(.A(men_men_n283_), .B(men_men_n282_), .C(men_men_n281_), .Y(men_men_n284_));
  NO3        u0262(.A(men_men_n26_), .B(men_men_n87_), .C(i_5_), .Y(men_men_n285_));
  NA3        u0263(.A(men_men_n285_), .B(men_men_n274_), .C(men_men_n230_), .Y(men_men_n286_));
  AOI210     u0264(.A0(men_men_n286_), .A1(men_men_n284_), .B0(men_men_n280_), .Y(men_men_n287_));
  INV        u0265(.A(men_men_n287_), .Y(men_men_n288_));
  NA4        u0266(.A(men_men_n288_), .B(men_men_n273_), .C(men_men_n255_), .D(men_men_n233_), .Y(men_men_n289_));
  NO3        u0267(.A(i_12_), .B(men_men_n229_), .C(men_men_n37_), .Y(men_men_n290_));
  INV        u0268(.A(men_men_n290_), .Y(men_men_n291_));
  NA2        u0269(.A(i_8_), .B(men_men_n103_), .Y(men_men_n292_));
  NOi21      u0270(.An(men_men_n164_), .B(men_men_n87_), .Y(men_men_n293_));
  NO3        u0271(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n294_));
  AOI220     u0272(.A0(men_men_n294_), .A1(men_men_n199_), .B0(men_men_n293_), .B1(men_men_n239_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n295_), .B(men_men_n292_), .Y(men_men_n296_));
  NO3        u0274(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n244_), .B(i_0_), .Y(men_men_n298_));
  AOI220     u0276(.A0(men_men_n298_), .A1(men_men_n197_), .B0(men_men_n297_), .B1(men_men_n143_), .Y(men_men_n299_));
  NA2        u0277(.A(men_men_n283_), .B(men_men_n26_), .Y(men_men_n300_));
  NO2        u0278(.A(men_men_n300_), .B(men_men_n299_), .Y(men_men_n301_));
  NA2        u0279(.A(i_0_), .B(i_1_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n302_), .B(i_2_), .Y(men_men_n303_));
  NO2        u0281(.A(men_men_n60_), .B(i_6_), .Y(men_men_n304_));
  NA3        u0282(.A(men_men_n304_), .B(men_men_n303_), .C(men_men_n164_), .Y(men_men_n305_));
  OAI210     u0283(.A0(men_men_n166_), .A1(men_men_n144_), .B0(men_men_n305_), .Y(men_men_n306_));
  NO3        u0284(.A(men_men_n306_), .B(men_men_n301_), .C(men_men_n296_), .Y(men_men_n307_));
  NO2        u0285(.A(i_3_), .B(i_10_), .Y(men_men_n308_));
  NA3        u0286(.A(men_men_n308_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n309_));
  NO2        u0287(.A(i_2_), .B(men_men_n103_), .Y(men_men_n310_));
  NA2        u0288(.A(i_1_), .B(men_men_n36_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n311_), .B(i_8_), .Y(men_men_n312_));
  NA2        u0290(.A(men_men_n312_), .B(men_men_n310_), .Y(men_men_n313_));
  AN2        u0291(.A(i_3_), .B(i_10_), .Y(men_men_n314_));
  NA4        u0292(.A(men_men_n314_), .B(men_men_n201_), .C(men_men_n178_), .D(men_men_n176_), .Y(men_men_n315_));
  NO2        u0293(.A(i_5_), .B(men_men_n37_), .Y(men_men_n316_));
  NO2        u0294(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n317_));
  OR2        u0295(.A(men_men_n313_), .B(men_men_n309_), .Y(men_men_n318_));
  OAI220     u0296(.A0(men_men_n318_), .A1(i_6_), .B0(men_men_n307_), .B1(men_men_n291_), .Y(men_men_n319_));
  NO4        u0297(.A(men_men_n319_), .B(men_men_n289_), .C(men_men_n217_), .D(men_men_n169_), .Y(men_men_n320_));
  NO3        u0298(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n321_));
  NO2        u0299(.A(men_men_n60_), .B(men_men_n87_), .Y(men_men_n322_));
  NA2        u0300(.A(men_men_n298_), .B(men_men_n322_), .Y(men_men_n323_));
  NO3        u0301(.A(i_6_), .B(men_men_n196_), .C(i_7_), .Y(men_men_n324_));
  NA2        u0302(.A(men_men_n324_), .B(men_men_n201_), .Y(men_men_n325_));
  AOI210     u0303(.A0(men_men_n325_), .A1(men_men_n323_), .B0(men_men_n171_), .Y(men_men_n326_));
  NO2        u0304(.A(i_2_), .B(i_3_), .Y(men_men_n327_));
  OR2        u0305(.A(i_0_), .B(i_5_), .Y(men_men_n328_));
  NA2        u0306(.A(men_men_n221_), .B(men_men_n328_), .Y(men_men_n329_));
  NA4        u0307(.A(men_men_n329_), .B(men_men_n238_), .C(men_men_n327_), .D(i_1_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n298_), .B(men_men_n293_), .C(men_men_n115_), .Y(men_men_n331_));
  NAi21      u0309(.An(i_8_), .B(i_7_), .Y(men_men_n332_));
  NO2        u0310(.A(men_men_n332_), .B(i_6_), .Y(men_men_n333_));
  NO2        u0311(.A(men_men_n158_), .B(men_men_n47_), .Y(men_men_n334_));
  NA3        u0312(.A(men_men_n334_), .B(men_men_n333_), .C(men_men_n164_), .Y(men_men_n335_));
  NA3        u0313(.A(men_men_n335_), .B(men_men_n331_), .C(men_men_n330_), .Y(men_men_n336_));
  OAI210     u0314(.A0(men_men_n336_), .A1(men_men_n326_), .B0(i_4_), .Y(men_men_n337_));
  NO2        u0315(.A(i_12_), .B(i_10_), .Y(men_men_n338_));
  NOi21      u0316(.An(i_5_), .B(i_0_), .Y(men_men_n339_));
  NO3        u0317(.A(men_men_n311_), .B(men_men_n339_), .C(men_men_n129_), .Y(men_men_n340_));
  NA4        u0318(.A(men_men_n85_), .B(men_men_n36_), .C(men_men_n87_), .D(i_8_), .Y(men_men_n341_));
  NA2        u0319(.A(men_men_n340_), .B(men_men_n338_), .Y(men_men_n342_));
  NO2        u0320(.A(i_6_), .B(i_8_), .Y(men_men_n343_));
  NOi21      u0321(.An(i_0_), .B(i_2_), .Y(men_men_n344_));
  AN2        u0322(.A(men_men_n344_), .B(men_men_n343_), .Y(men_men_n345_));
  NO2        u0323(.A(i_1_), .B(i_7_), .Y(men_men_n346_));
  AO220      u0324(.A0(men_men_n346_), .A1(men_men_n345_), .B0(men_men_n333_), .B1(men_men_n239_), .Y(men_men_n347_));
  NA3        u0325(.A(men_men_n347_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n348_));
  NA3        u0326(.A(men_men_n348_), .B(men_men_n342_), .C(men_men_n337_), .Y(men_men_n349_));
  NO3        u0327(.A(men_men_n237_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n350_));
  NO3        u0328(.A(men_men_n332_), .B(i_2_), .C(i_1_), .Y(men_men_n351_));
  OAI210     u0329(.A0(men_men_n351_), .A1(men_men_n350_), .B0(i_6_), .Y(men_men_n352_));
  NA3        u0330(.A(men_men_n257_), .B(men_men_n310_), .C(men_men_n196_), .Y(men_men_n353_));
  AOI210     u0331(.A0(men_men_n353_), .A1(men_men_n352_), .B0(men_men_n329_), .Y(men_men_n354_));
  NOi21      u0332(.An(men_men_n154_), .B(men_men_n106_), .Y(men_men_n355_));
  NO2        u0333(.A(men_men_n355_), .B(men_men_n125_), .Y(men_men_n356_));
  OAI210     u0334(.A0(men_men_n356_), .A1(men_men_n354_), .B0(i_3_), .Y(men_men_n357_));
  INV        u0335(.A(men_men_n85_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n302_), .B(men_men_n82_), .Y(men_men_n359_));
  NA2        u0337(.A(men_men_n359_), .B(men_men_n133_), .Y(men_men_n360_));
  NO2        u0338(.A(men_men_n94_), .B(men_men_n196_), .Y(men_men_n361_));
  NA2        u0339(.A(men_men_n361_), .B(men_men_n64_), .Y(men_men_n362_));
  AOI210     u0340(.A0(men_men_n362_), .A1(men_men_n360_), .B0(men_men_n358_), .Y(men_men_n363_));
  NO2        u0341(.A(men_men_n196_), .B(i_9_), .Y(men_men_n364_));
  NA2        u0342(.A(men_men_n364_), .B(men_men_n208_), .Y(men_men_n365_));
  NO2        u0343(.A(men_men_n365_), .B(men_men_n47_), .Y(men_men_n366_));
  NO3        u0344(.A(men_men_n366_), .B(men_men_n363_), .C(men_men_n301_), .Y(men_men_n367_));
  AOI210     u0345(.A0(men_men_n367_), .A1(men_men_n357_), .B0(men_men_n163_), .Y(men_men_n368_));
  AOI210     u0346(.A0(men_men_n349_), .A1(men_men_n321_), .B0(men_men_n368_), .Y(men_men_n369_));
  NOi32      u0347(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n370_));
  INV        u0348(.A(men_men_n370_), .Y(men_men_n371_));
  NAi21      u0349(.An(i_0_), .B(i_6_), .Y(men_men_n372_));
  NAi21      u0350(.An(i_1_), .B(i_5_), .Y(men_men_n373_));
  NA2        u0351(.A(men_men_n373_), .B(men_men_n372_), .Y(men_men_n374_));
  NA2        u0352(.A(men_men_n374_), .B(men_men_n25_), .Y(men_men_n375_));
  OAI210     u0353(.A0(men_men_n375_), .A1(men_men_n160_), .B0(men_men_n251_), .Y(men_men_n376_));
  NAi41      u0354(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n377_));
  AOI210     u0355(.A0(men_men_n377_), .A1(men_men_n160_), .B0(men_men_n158_), .Y(men_men_n378_));
  NOi32      u0356(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n379_));
  NAi21      u0357(.An(i_6_), .B(i_1_), .Y(men_men_n380_));
  NA3        u0358(.A(men_men_n380_), .B(men_men_n379_), .C(men_men_n47_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n381_), .B(i_0_), .Y(men_men_n382_));
  OR2        u0360(.A(men_men_n382_), .B(men_men_n378_), .Y(men_men_n383_));
  NO2        u0361(.A(i_1_), .B(men_men_n103_), .Y(men_men_n384_));
  NAi21      u0362(.An(i_3_), .B(i_4_), .Y(men_men_n385_));
  NO2        u0363(.A(men_men_n385_), .B(i_9_), .Y(men_men_n386_));
  AN2        u0364(.A(i_6_), .B(i_7_), .Y(men_men_n387_));
  OAI210     u0365(.A0(men_men_n387_), .A1(men_men_n384_), .B0(men_men_n386_), .Y(men_men_n388_));
  NA2        u0366(.A(i_2_), .B(i_7_), .Y(men_men_n389_));
  NO2        u0367(.A(men_men_n385_), .B(i_10_), .Y(men_men_n390_));
  NA3        u0368(.A(men_men_n390_), .B(men_men_n389_), .C(men_men_n249_), .Y(men_men_n391_));
  AOI210     u0369(.A0(men_men_n391_), .A1(men_men_n388_), .B0(men_men_n188_), .Y(men_men_n392_));
  AOI210     u0370(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n393_));
  OAI210     u0371(.A0(men_men_n393_), .A1(men_men_n191_), .B0(men_men_n390_), .Y(men_men_n394_));
  AOI220     u0372(.A0(men_men_n390_), .A1(men_men_n346_), .B0(men_men_n243_), .B1(men_men_n191_), .Y(men_men_n395_));
  AOI210     u0373(.A0(men_men_n395_), .A1(men_men_n394_), .B0(i_5_), .Y(men_men_n396_));
  NO4        u0374(.A(men_men_n396_), .B(men_men_n392_), .C(men_men_n383_), .D(men_men_n376_), .Y(men_men_n397_));
  NO2        u0375(.A(men_men_n397_), .B(men_men_n371_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n60_), .B(men_men_n25_), .Y(men_men_n399_));
  AN2        u0377(.A(i_12_), .B(i_5_), .Y(men_men_n400_));
  NO2        u0378(.A(i_4_), .B(men_men_n26_), .Y(men_men_n401_));
  NA2        u0379(.A(men_men_n401_), .B(men_men_n400_), .Y(men_men_n402_));
  NO2        u0380(.A(i_11_), .B(i_6_), .Y(men_men_n403_));
  NA3        u0381(.A(men_men_n403_), .B(men_men_n334_), .C(men_men_n229_), .Y(men_men_n404_));
  NO2        u0382(.A(men_men_n404_), .B(men_men_n402_), .Y(men_men_n405_));
  NO2        u0383(.A(men_men_n247_), .B(i_5_), .Y(men_men_n406_));
  NO2        u0384(.A(i_5_), .B(i_10_), .Y(men_men_n407_));
  AOI220     u0385(.A0(men_men_n407_), .A1(men_men_n278_), .B0(men_men_n406_), .B1(men_men_n201_), .Y(men_men_n408_));
  NA2        u0386(.A(men_men_n145_), .B(men_men_n46_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n409_), .B(men_men_n408_), .Y(men_men_n410_));
  OAI210     u0388(.A0(men_men_n410_), .A1(men_men_n405_), .B0(men_men_n399_), .Y(men_men_n411_));
  NO2        u0389(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n412_));
  NO2        u0390(.A(men_men_n151_), .B(men_men_n87_), .Y(men_men_n413_));
  OAI210     u0391(.A0(men_men_n413_), .A1(men_men_n405_), .B0(men_men_n412_), .Y(men_men_n414_));
  NO3        u0392(.A(men_men_n87_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n415_));
  NO2        u0393(.A(i_3_), .B(men_men_n103_), .Y(men_men_n416_));
  NO2        u0394(.A(i_11_), .B(i_12_), .Y(men_men_n417_));
  NA2        u0395(.A(men_men_n407_), .B(men_men_n241_), .Y(men_men_n418_));
  NA3        u0396(.A(men_men_n115_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n419_));
  OAI220     u0397(.A0(men_men_n419_), .A1(men_men_n224_), .B0(men_men_n418_), .B1(men_men_n341_), .Y(men_men_n420_));
  NAi21      u0398(.An(i_13_), .B(i_0_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n421_), .B(men_men_n244_), .Y(men_men_n422_));
  NA2        u0400(.A(men_men_n420_), .B(men_men_n422_), .Y(men_men_n423_));
  NA3        u0401(.A(men_men_n423_), .B(men_men_n414_), .C(men_men_n411_), .Y(men_men_n424_));
  NO3        u0402(.A(i_1_), .B(i_12_), .C(men_men_n87_), .Y(men_men_n425_));
  NO2        u0403(.A(i_0_), .B(i_11_), .Y(men_men_n426_));
  INV        u0404(.A(i_5_), .Y(men_men_n427_));
  AN2        u0405(.A(i_1_), .B(i_6_), .Y(men_men_n428_));
  NOi21      u0406(.An(i_2_), .B(i_12_), .Y(men_men_n429_));
  NA2        u0407(.A(men_men_n429_), .B(men_men_n428_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n430_), .B(men_men_n427_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n143_), .B(i_9_), .Y(men_men_n432_));
  NO2        u0410(.A(men_men_n432_), .B(i_4_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n431_), .B(men_men_n433_), .Y(men_men_n434_));
  NAi21      u0412(.An(i_9_), .B(i_4_), .Y(men_men_n435_));
  OR2        u0413(.A(i_13_), .B(i_10_), .Y(men_men_n436_));
  NO3        u0414(.A(men_men_n436_), .B(men_men_n119_), .C(men_men_n435_), .Y(men_men_n437_));
  NO2        u0415(.A(men_men_n174_), .B(men_men_n124_), .Y(men_men_n438_));
  OR2        u0416(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n439_));
  NO2        u0417(.A(men_men_n103_), .B(men_men_n25_), .Y(men_men_n440_));
  NA2        u0418(.A(men_men_n290_), .B(men_men_n440_), .Y(men_men_n441_));
  NA2        u0419(.A(men_men_n283_), .B(men_men_n213_), .Y(men_men_n442_));
  OAI220     u0420(.A0(men_men_n442_), .A1(men_men_n439_), .B0(men_men_n441_), .B1(men_men_n355_), .Y(men_men_n443_));
  INV        u0421(.A(men_men_n443_), .Y(men_men_n444_));
  AOI210     u0422(.A0(men_men_n444_), .A1(men_men_n434_), .B0(men_men_n26_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n331_), .B(men_men_n330_), .Y(men_men_n446_));
  AOI220     u0424(.A0(men_men_n304_), .A1(men_men_n294_), .B0(men_men_n298_), .B1(men_men_n322_), .Y(men_men_n447_));
  NO2        u0425(.A(men_men_n447_), .B(men_men_n171_), .Y(men_men_n448_));
  NO2        u0426(.A(men_men_n185_), .B(men_men_n87_), .Y(men_men_n449_));
  AOI220     u0427(.A0(men_men_n449_), .A1(men_men_n303_), .B0(men_men_n285_), .B1(men_men_n213_), .Y(men_men_n450_));
  NO2        u0428(.A(men_men_n450_), .B(men_men_n292_), .Y(men_men_n451_));
  NO3        u0429(.A(men_men_n451_), .B(men_men_n448_), .C(men_men_n446_), .Y(men_men_n452_));
  NA2        u0430(.A(men_men_n199_), .B(men_men_n98_), .Y(men_men_n453_));
  NA3        u0431(.A(men_men_n334_), .B(men_men_n164_), .C(men_men_n87_), .Y(men_men_n454_));
  AOI210     u0432(.A0(men_men_n454_), .A1(men_men_n453_), .B0(men_men_n332_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n196_), .B(i_10_), .Y(men_men_n456_));
  NA3        u0434(.A(men_men_n263_), .B(men_men_n65_), .C(i_2_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n304_), .B(men_men_n239_), .Y(men_men_n458_));
  OAI220     u0436(.A0(men_men_n458_), .A1(men_men_n185_), .B0(men_men_n457_), .B1(men_men_n456_), .Y(men_men_n459_));
  NO2        u0437(.A(i_3_), .B(men_men_n49_), .Y(men_men_n460_));
  NA3        u0438(.A(men_men_n346_), .B(men_men_n345_), .C(men_men_n460_), .Y(men_men_n461_));
  NA2        u0439(.A(men_men_n324_), .B(men_men_n329_), .Y(men_men_n462_));
  OAI210     u0440(.A0(men_men_n462_), .A1(men_men_n192_), .B0(men_men_n461_), .Y(men_men_n463_));
  NO3        u0441(.A(men_men_n463_), .B(men_men_n459_), .C(men_men_n455_), .Y(men_men_n464_));
  AOI210     u0442(.A0(men_men_n464_), .A1(men_men_n452_), .B0(men_men_n279_), .Y(men_men_n465_));
  NO4        u0443(.A(men_men_n465_), .B(men_men_n445_), .C(men_men_n424_), .D(men_men_n398_), .Y(men_men_n466_));
  NO2        u0444(.A(men_men_n64_), .B(i_4_), .Y(men_men_n467_));
  NO2        u0445(.A(men_men_n74_), .B(i_13_), .Y(men_men_n468_));
  NO2        u0446(.A(i_10_), .B(i_9_), .Y(men_men_n469_));
  NAi21      u0447(.An(i_12_), .B(i_8_), .Y(men_men_n470_));
  NO2        u0448(.A(men_men_n470_), .B(i_3_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n47_), .B(i_4_), .Y(men_men_n472_));
  NA2        u0450(.A(men_men_n317_), .B(i_0_), .Y(men_men_n473_));
  NO3        u0451(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n275_), .B(men_men_n99_), .Y(men_men_n475_));
  NA2        u0453(.A(men_men_n475_), .B(men_men_n474_), .Y(men_men_n476_));
  NA2        u0454(.A(i_8_), .B(i_9_), .Y(men_men_n477_));
  AOI210     u0455(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n478_));
  OR2        u0456(.A(men_men_n478_), .B(men_men_n477_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n290_), .B(men_men_n208_), .Y(men_men_n480_));
  NO2        u0458(.A(men_men_n480_), .B(men_men_n479_), .Y(men_men_n481_));
  NA2        u0459(.A(men_men_n256_), .B(men_men_n316_), .Y(men_men_n482_));
  NO3        u0460(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n483_));
  INV        u0461(.A(men_men_n483_), .Y(men_men_n484_));
  NA3        u0462(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n485_));
  NA4        u0463(.A(men_men_n146_), .B(men_men_n118_), .C(men_men_n81_), .D(men_men_n23_), .Y(men_men_n486_));
  OAI220     u0464(.A0(men_men_n486_), .A1(men_men_n485_), .B0(men_men_n484_), .B1(men_men_n482_), .Y(men_men_n487_));
  NO2        u0465(.A(men_men_n487_), .B(men_men_n481_), .Y(men_men_n488_));
  INV        u0466(.A(men_men_n303_), .Y(men_men_n489_));
  OR2        u0467(.A(men_men_n489_), .B(men_men_n210_), .Y(men_men_n490_));
  OA210      u0468(.A0(men_men_n365_), .A1(men_men_n103_), .B0(men_men_n305_), .Y(men_men_n491_));
  OA220      u0469(.A0(men_men_n491_), .A1(men_men_n163_), .B0(men_men_n490_), .B1(men_men_n236_), .Y(men_men_n492_));
  NA2        u0470(.A(men_men_n98_), .B(i_13_), .Y(men_men_n493_));
  NA2        u0471(.A(men_men_n449_), .B(men_men_n399_), .Y(men_men_n494_));
  NO2        u0472(.A(i_2_), .B(i_13_), .Y(men_men_n495_));
  NO2        u0473(.A(men_men_n494_), .B(men_men_n493_), .Y(men_men_n496_));
  NO3        u0474(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n497_));
  NO2        u0475(.A(i_6_), .B(i_7_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n498_), .B(men_men_n497_), .Y(men_men_n499_));
  NO2        u0477(.A(i_11_), .B(i_1_), .Y(men_men_n500_));
  NO2        u0478(.A(men_men_n74_), .B(i_3_), .Y(men_men_n501_));
  OR2        u0479(.A(i_11_), .B(i_8_), .Y(men_men_n502_));
  NOi21      u0480(.An(i_2_), .B(i_7_), .Y(men_men_n503_));
  NAi31      u0481(.An(men_men_n502_), .B(men_men_n503_), .C(men_men_n501_), .Y(men_men_n504_));
  NO2        u0482(.A(men_men_n436_), .B(i_6_), .Y(men_men_n505_));
  NA2        u0483(.A(men_men_n505_), .B(men_men_n467_), .Y(men_men_n506_));
  NO2        u0484(.A(men_men_n506_), .B(men_men_n504_), .Y(men_men_n507_));
  NO2        u0485(.A(i_3_), .B(men_men_n196_), .Y(men_men_n508_));
  NO2        u0486(.A(i_6_), .B(i_10_), .Y(men_men_n509_));
  NA4        u0487(.A(men_men_n509_), .B(men_men_n321_), .C(men_men_n508_), .D(men_men_n241_), .Y(men_men_n510_));
  NO2        u0488(.A(men_men_n510_), .B(men_men_n156_), .Y(men_men_n511_));
  NA3        u0489(.A(men_men_n250_), .B(men_men_n173_), .C(men_men_n133_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n513_));
  NO2        u0491(.A(men_men_n158_), .B(i_3_), .Y(men_men_n514_));
  NAi31      u0492(.An(men_men_n513_), .B(men_men_n514_), .C(men_men_n230_), .Y(men_men_n515_));
  NA3        u0493(.A(men_men_n412_), .B(men_men_n181_), .C(men_men_n150_), .Y(men_men_n516_));
  NA3        u0494(.A(men_men_n516_), .B(men_men_n515_), .C(men_men_n512_), .Y(men_men_n517_));
  NO4        u0495(.A(men_men_n517_), .B(men_men_n511_), .C(men_men_n507_), .D(men_men_n496_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n474_), .B(men_men_n400_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n483_), .B(men_men_n407_), .Y(men_men_n520_));
  NO2        u0498(.A(men_men_n520_), .B(men_men_n228_), .Y(men_men_n521_));
  NAi21      u0499(.An(men_men_n219_), .B(men_men_n417_), .Y(men_men_n522_));
  NO2        u0500(.A(men_men_n26_), .B(i_5_), .Y(men_men_n523_));
  NO2        u0501(.A(i_0_), .B(men_men_n87_), .Y(men_men_n524_));
  NA3        u0502(.A(men_men_n524_), .B(men_men_n523_), .C(men_men_n143_), .Y(men_men_n525_));
  OR3        u0503(.A(men_men_n311_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n526_));
  NO2        u0504(.A(men_men_n526_), .B(men_men_n525_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n27_), .B(i_10_), .Y(men_men_n528_));
  NA2        u0506(.A(men_men_n321_), .B(men_men_n243_), .Y(men_men_n529_));
  OAI220     u0507(.A0(men_men_n529_), .A1(men_men_n457_), .B0(men_men_n528_), .B1(men_men_n493_), .Y(men_men_n530_));
  NA4        u0508(.A(men_men_n314_), .B(men_men_n227_), .C(men_men_n74_), .D(men_men_n241_), .Y(men_men_n531_));
  NO2        u0509(.A(men_men_n531_), .B(men_men_n499_), .Y(men_men_n532_));
  NO4        u0510(.A(men_men_n532_), .B(men_men_n530_), .C(men_men_n527_), .D(men_men_n521_), .Y(men_men_n533_));
  NA4        u0511(.A(men_men_n533_), .B(men_men_n518_), .C(men_men_n492_), .D(men_men_n488_), .Y(men_men_n534_));
  NA3        u0512(.A(men_men_n314_), .B(men_men_n178_), .C(men_men_n176_), .Y(men_men_n535_));
  OAI210     u0513(.A0(men_men_n309_), .A1(men_men_n183_), .B0(men_men_n535_), .Y(men_men_n536_));
  AN2        u0514(.A(men_men_n294_), .B(men_men_n238_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n537_), .B(men_men_n536_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n321_), .B(men_men_n165_), .Y(men_men_n539_));
  OAI210     u0517(.A0(men_men_n539_), .A1(men_men_n236_), .B0(men_men_n315_), .Y(men_men_n540_));
  NA2        u0518(.A(men_men_n540_), .B(men_men_n333_), .Y(men_men_n541_));
  NA2        u0519(.A(men_men_n400_), .B(men_men_n229_), .Y(men_men_n542_));
  NA2        u0520(.A(men_men_n370_), .B(men_men_n74_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n387_), .B(men_men_n379_), .Y(men_men_n544_));
  AO210      u0522(.A0(men_men_n543_), .A1(men_men_n542_), .B0(men_men_n544_), .Y(men_men_n545_));
  NO2        u0523(.A(men_men_n36_), .B(i_8_), .Y(men_men_n546_));
  NAi41      u0524(.An(men_men_n543_), .B(men_men_n509_), .C(men_men_n546_), .D(men_men_n47_), .Y(men_men_n547_));
  AOI210     u0525(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n437_), .Y(men_men_n548_));
  NA3        u0526(.A(men_men_n548_), .B(men_men_n547_), .C(men_men_n545_), .Y(men_men_n549_));
  INV        u0527(.A(men_men_n549_), .Y(men_men_n550_));
  NA2        u0528(.A(men_men_n263_), .B(men_men_n65_), .Y(men_men_n551_));
  OAI210     u0529(.A0(i_8_), .A1(men_men_n551_), .B0(men_men_n135_), .Y(men_men_n552_));
  AOI210     u0530(.A0(men_men_n197_), .A1(i_9_), .B0(men_men_n274_), .Y(men_men_n553_));
  NO2        u0531(.A(men_men_n553_), .B(men_men_n202_), .Y(men_men_n554_));
  OR2        u0532(.A(men_men_n185_), .B(i_4_), .Y(men_men_n555_));
  NO2        u0533(.A(men_men_n555_), .B(men_men_n87_), .Y(men_men_n556_));
  AOI220     u0534(.A0(men_men_n556_), .A1(men_men_n554_), .B0(men_men_n552_), .B1(men_men_n438_), .Y(men_men_n557_));
  NA4        u0535(.A(men_men_n557_), .B(men_men_n550_), .C(men_men_n541_), .D(men_men_n538_), .Y(men_men_n558_));
  NA2        u0536(.A(men_men_n406_), .B(men_men_n303_), .Y(men_men_n559_));
  OAI210     u0537(.A0(men_men_n402_), .A1(men_men_n170_), .B0(men_men_n559_), .Y(men_men_n560_));
  NO2        u0538(.A(i_12_), .B(men_men_n196_), .Y(men_men_n561_));
  NA2        u0539(.A(men_men_n561_), .B(men_men_n229_), .Y(men_men_n562_));
  NA3        u0540(.A(men_men_n509_), .B(men_men_n176_), .C(men_men_n27_), .Y(men_men_n563_));
  NO2        u0541(.A(men_men_n563_), .B(men_men_n562_), .Y(men_men_n564_));
  NOi31      u0542(.An(men_men_n324_), .B(men_men_n436_), .C(men_men_n38_), .Y(men_men_n565_));
  OAI210     u0543(.A0(men_men_n565_), .A1(men_men_n564_), .B0(men_men_n560_), .Y(men_men_n566_));
  NO2        u0544(.A(i_8_), .B(i_7_), .Y(men_men_n567_));
  OAI210     u0545(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n568_));
  NA2        u0546(.A(men_men_n568_), .B(men_men_n227_), .Y(men_men_n569_));
  AOI220     u0547(.A0(men_men_n334_), .A1(men_men_n40_), .B0(men_men_n239_), .B1(men_men_n209_), .Y(men_men_n570_));
  OAI220     u0548(.A0(men_men_n570_), .A1(men_men_n555_), .B0(men_men_n569_), .B1(men_men_n247_), .Y(men_men_n571_));
  NA2        u0549(.A(men_men_n45_), .B(i_10_), .Y(men_men_n572_));
  NO2        u0550(.A(men_men_n572_), .B(i_6_), .Y(men_men_n573_));
  NA3        u0551(.A(men_men_n573_), .B(men_men_n571_), .C(men_men_n567_), .Y(men_men_n574_));
  NOi31      u0552(.An(men_men_n298_), .B(men_men_n309_), .C(men_men_n183_), .Y(men_men_n575_));
  NO2        u0553(.A(men_men_n158_), .B(i_5_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n575_), .B(men_men_n483_), .Y(men_men_n577_));
  NA3        u0555(.A(men_men_n577_), .B(men_men_n574_), .C(men_men_n566_), .Y(men_men_n578_));
  NA3        u0556(.A(men_men_n221_), .B(men_men_n72_), .C(men_men_n45_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n290_), .B(men_men_n85_), .Y(men_men_n580_));
  AOI210     u0558(.A0(men_men_n579_), .A1(men_men_n360_), .B0(men_men_n580_), .Y(men_men_n581_));
  NA2        u0559(.A(men_men_n304_), .B(men_men_n294_), .Y(men_men_n582_));
  NO2        u0560(.A(men_men_n582_), .B(men_men_n175_), .Y(men_men_n583_));
  NA2        u0561(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n584_));
  NA2        u0562(.A(men_men_n469_), .B(men_men_n225_), .Y(men_men_n585_));
  NO2        u0563(.A(men_men_n584_), .B(men_men_n585_), .Y(men_men_n586_));
  AOI210     u0564(.A0(men_men_n380_), .A1(men_men_n47_), .B0(men_men_n384_), .Y(men_men_n587_));
  NA2        u0565(.A(i_0_), .B(men_men_n49_), .Y(men_men_n588_));
  NA3        u0566(.A(men_men_n561_), .B(men_men_n281_), .C(men_men_n588_), .Y(men_men_n589_));
  NO2        u0567(.A(men_men_n587_), .B(men_men_n589_), .Y(men_men_n590_));
  NO4        u0568(.A(men_men_n590_), .B(men_men_n586_), .C(men_men_n583_), .D(men_men_n581_), .Y(men_men_n591_));
  NO4        u0569(.A(men_men_n257_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n592_));
  NO3        u0570(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n237_), .B(men_men_n36_), .Y(men_men_n594_));
  AN2        u0572(.A(men_men_n594_), .B(men_men_n593_), .Y(men_men_n595_));
  OA210      u0573(.A0(men_men_n595_), .A1(men_men_n592_), .B0(men_men_n370_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n436_), .B(i_1_), .Y(men_men_n597_));
  NOi31      u0575(.An(men_men_n597_), .B(men_men_n475_), .C(men_men_n74_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n447_), .B(men_men_n179_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n599_), .B(men_men_n596_), .Y(men_men_n600_));
  NOi21      u0578(.An(i_10_), .B(i_6_), .Y(men_men_n601_));
  NO2        u0579(.A(men_men_n87_), .B(men_men_n25_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n117_), .B(men_men_n23_), .Y(men_men_n603_));
  NA2        u0581(.A(men_men_n324_), .B(men_men_n165_), .Y(men_men_n604_));
  AOI220     u0582(.A0(men_men_n604_), .A1(men_men_n458_), .B0(men_men_n186_), .B1(men_men_n184_), .Y(men_men_n605_));
  NOi31      u0583(.An(men_men_n147_), .B(i_10_), .C(men_men_n341_), .Y(men_men_n606_));
  NO2        u0584(.A(men_men_n606_), .B(men_men_n605_), .Y(men_men_n607_));
  INV        u0585(.A(men_men_n327_), .Y(men_men_n608_));
  NO2        u0586(.A(i_12_), .B(men_men_n87_), .Y(men_men_n609_));
  NA3        u0587(.A(men_men_n609_), .B(men_men_n281_), .C(men_men_n588_), .Y(men_men_n610_));
  NA3        u0588(.A(men_men_n403_), .B(men_men_n290_), .C(men_men_n221_), .Y(men_men_n611_));
  AOI210     u0589(.A0(men_men_n611_), .A1(men_men_n610_), .B0(men_men_n608_), .Y(men_men_n612_));
  NA2        u0590(.A(men_men_n176_), .B(i_0_), .Y(men_men_n613_));
  NO3        u0591(.A(men_men_n613_), .B(men_men_n352_), .C(men_men_n309_), .Y(men_men_n614_));
  OR2        u0592(.A(i_2_), .B(i_5_), .Y(men_men_n615_));
  OR2        u0593(.A(men_men_n615_), .B(men_men_n428_), .Y(men_men_n616_));
  AOI210     u0594(.A0(men_men_n389_), .A1(men_men_n249_), .B0(men_men_n201_), .Y(men_men_n617_));
  AOI210     u0595(.A0(men_men_n617_), .A1(men_men_n616_), .B0(men_men_n522_), .Y(men_men_n618_));
  NO3        u0596(.A(men_men_n618_), .B(men_men_n614_), .C(men_men_n612_), .Y(men_men_n619_));
  NA4        u0597(.A(men_men_n619_), .B(men_men_n607_), .C(men_men_n600_), .D(men_men_n591_), .Y(men_men_n620_));
  NO4        u0598(.A(men_men_n620_), .B(men_men_n578_), .C(men_men_n558_), .D(men_men_n534_), .Y(men_men_n621_));
  NA4        u0599(.A(men_men_n621_), .B(men_men_n466_), .C(men_men_n369_), .D(men_men_n320_), .Y(men7));
  NO2        u0600(.A(men_men_n94_), .B(men_men_n55_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n110_), .B(men_men_n91_), .Y(men_men_n624_));
  NA2        u0602(.A(men_men_n401_), .B(men_men_n624_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n509_), .B(men_men_n85_), .Y(men_men_n626_));
  NA2        u0604(.A(i_11_), .B(men_men_n196_), .Y(men_men_n627_));
  NA2        u0605(.A(men_men_n145_), .B(men_men_n627_), .Y(men_men_n628_));
  OAI210     u0606(.A0(men_men_n628_), .A1(men_men_n626_), .B0(men_men_n625_), .Y(men_men_n629_));
  NA3        u0607(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n630_));
  NO2        u0608(.A(men_men_n241_), .B(i_4_), .Y(men_men_n631_));
  NA2        u0609(.A(men_men_n631_), .B(i_8_), .Y(men_men_n632_));
  NO2        u0610(.A(men_men_n107_), .B(men_men_n630_), .Y(men_men_n633_));
  NA2        u0611(.A(i_2_), .B(men_men_n87_), .Y(men_men_n634_));
  OAI210     u0612(.A0(men_men_n88_), .A1(men_men_n206_), .B0(men_men_n207_), .Y(men_men_n635_));
  NO2        u0613(.A(i_7_), .B(men_men_n37_), .Y(men_men_n636_));
  NA2        u0614(.A(i_4_), .B(i_8_), .Y(men_men_n637_));
  AOI210     u0615(.A0(men_men_n637_), .A1(men_men_n314_), .B0(men_men_n636_), .Y(men_men_n638_));
  OAI220     u0616(.A0(men_men_n638_), .A1(men_men_n634_), .B0(men_men_n635_), .B1(i_13_), .Y(men_men_n639_));
  NO4        u0617(.A(men_men_n639_), .B(men_men_n633_), .C(men_men_n629_), .D(men_men_n623_), .Y(men_men_n640_));
  AOI210     u0618(.A0(men_men_n129_), .A1(men_men_n63_), .B0(i_10_), .Y(men_men_n641_));
  AOI210     u0619(.A0(men_men_n641_), .A1(men_men_n241_), .B0(men_men_n162_), .Y(men_men_n642_));
  OR2        u0620(.A(i_6_), .B(i_10_), .Y(men_men_n643_));
  NO2        u0621(.A(men_men_n643_), .B(men_men_n23_), .Y(men_men_n644_));
  OR3        u0622(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n645_));
  NO3        u0623(.A(men_men_n645_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n646_));
  INV        u0624(.A(men_men_n203_), .Y(men_men_n647_));
  NO2        u0625(.A(men_men_n646_), .B(men_men_n644_), .Y(men_men_n648_));
  OA220      u0626(.A0(men_men_n648_), .A1(men_men_n608_), .B0(men_men_n642_), .B1(men_men_n276_), .Y(men_men_n649_));
  AOI210     u0627(.A0(men_men_n649_), .A1(men_men_n640_), .B0(men_men_n64_), .Y(men_men_n650_));
  NOi21      u0628(.An(i_11_), .B(i_7_), .Y(men_men_n651_));
  AO210      u0629(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n652_), .B(men_men_n651_), .Y(men_men_n653_));
  NA2        u0631(.A(men_men_n653_), .B(men_men_n209_), .Y(men_men_n654_));
  NA3        u0632(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n655_));
  NAi31      u0633(.An(men_men_n655_), .B(men_men_n218_), .C(i_11_), .Y(men_men_n656_));
  AOI210     u0634(.A0(men_men_n656_), .A1(men_men_n654_), .B0(men_men_n64_), .Y(men_men_n657_));
  OR2        u0635(.A(men_men_n395_), .B(men_men_n41_), .Y(men_men_n658_));
  NO3        u0636(.A(men_men_n265_), .B(men_men_n211_), .C(men_men_n627_), .Y(men_men_n659_));
  OAI210     u0637(.A0(men_men_n659_), .A1(men_men_n230_), .B0(men_men_n64_), .Y(men_men_n660_));
  NA2        u0638(.A(men_men_n429_), .B(men_men_n31_), .Y(men_men_n661_));
  OR2        u0639(.A(men_men_n211_), .B(men_men_n110_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(men_men_n661_), .Y(men_men_n663_));
  NO2        u0641(.A(men_men_n64_), .B(i_9_), .Y(men_men_n664_));
  NO2        u0642(.A(men_men_n664_), .B(i_4_), .Y(men_men_n665_));
  NA2        u0643(.A(men_men_n665_), .B(men_men_n663_), .Y(men_men_n666_));
  NO2        u0644(.A(i_1_), .B(i_12_), .Y(men_men_n667_));
  NA3        u0645(.A(men_men_n666_), .B(men_men_n660_), .C(men_men_n658_), .Y(men_men_n668_));
  OAI210     u0646(.A0(men_men_n668_), .A1(men_men_n657_), .B0(i_6_), .Y(men_men_n669_));
  NO2        u0647(.A(men_men_n655_), .B(men_men_n110_), .Y(men_men_n670_));
  NA2        u0648(.A(men_men_n670_), .B(men_men_n609_), .Y(men_men_n671_));
  NO2        u0649(.A(men_men_n241_), .B(men_men_n87_), .Y(men_men_n672_));
  NO2        u0650(.A(men_men_n672_), .B(i_11_), .Y(men_men_n673_));
  NA2        u0651(.A(men_men_n671_), .B(men_men_n476_), .Y(men_men_n674_));
  NO4        u0652(.A(men_men_n218_), .B(men_men_n129_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n675_), .B(men_men_n664_), .Y(men_men_n676_));
  NA2        u0654(.A(men_men_n241_), .B(i_6_), .Y(men_men_n677_));
  NO3        u0655(.A(men_men_n643_), .B(men_men_n237_), .C(men_men_n23_), .Y(men_men_n678_));
  AOI210     u0656(.A0(i_1_), .A1(men_men_n266_), .B0(men_men_n678_), .Y(men_men_n679_));
  OAI210     u0657(.A0(men_men_n679_), .A1(men_men_n45_), .B0(men_men_n676_), .Y(men_men_n680_));
  NA3        u0658(.A(men_men_n567_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n681_));
  NA2        u0659(.A(men_men_n139_), .B(i_9_), .Y(men_men_n682_));
  NA3        u0660(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n683_));
  NO2        u0661(.A(men_men_n47_), .B(i_1_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n682_), .B(men_men_n1092_), .Y(men_men_n685_));
  NA3        u0663(.A(men_men_n664_), .B(men_men_n327_), .C(i_6_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n686_), .B(men_men_n23_), .Y(men_men_n687_));
  AOI210     u0665(.A0(men_men_n500_), .A1(men_men_n440_), .B0(men_men_n246_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n688_), .B(men_men_n634_), .Y(men_men_n689_));
  NAi21      u0667(.An(men_men_n681_), .B(men_men_n93_), .Y(men_men_n690_));
  NA2        u0668(.A(men_men_n684_), .B(men_men_n275_), .Y(men_men_n691_));
  NO2        u0669(.A(i_11_), .B(men_men_n37_), .Y(men_men_n692_));
  NA2        u0670(.A(men_men_n692_), .B(men_men_n24_), .Y(men_men_n693_));
  OAI210     u0671(.A0(men_men_n693_), .A1(men_men_n691_), .B0(men_men_n690_), .Y(men_men_n694_));
  OR4        u0672(.A(men_men_n694_), .B(men_men_n689_), .C(men_men_n687_), .D(men_men_n685_), .Y(men_men_n695_));
  NO3        u0673(.A(men_men_n695_), .B(men_men_n680_), .C(men_men_n674_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n241_), .B(men_men_n103_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n697_), .B(men_men_n651_), .Y(men_men_n698_));
  NA2        u0676(.A(men_men_n698_), .B(i_1_), .Y(men_men_n699_));
  NO2        u0677(.A(men_men_n699_), .B(men_men_n645_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n435_), .B(men_men_n87_), .Y(men_men_n701_));
  NA2        u0679(.A(men_men_n700_), .B(men_men_n47_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n237_), .B(men_men_n45_), .Y(men_men_n703_));
  NO3        u0681(.A(men_men_n703_), .B(men_men_n317_), .C(men_men_n242_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n119_), .B(men_men_n37_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(i_6_), .Y(men_men_n706_));
  NO2        u0684(.A(men_men_n87_), .B(i_9_), .Y(men_men_n707_));
  NO2        u0685(.A(men_men_n707_), .B(men_men_n64_), .Y(men_men_n708_));
  NO2        u0686(.A(men_men_n708_), .B(men_men_n667_), .Y(men_men_n709_));
  NO4        u0687(.A(men_men_n709_), .B(men_men_n706_), .C(men_men_n704_), .D(i_4_), .Y(men_men_n710_));
  NA2        u0688(.A(i_1_), .B(i_3_), .Y(men_men_n711_));
  INV        u0689(.A(men_men_n710_), .Y(men_men_n712_));
  NA4        u0690(.A(men_men_n712_), .B(men_men_n702_), .C(men_men_n696_), .D(men_men_n669_), .Y(men_men_n713_));
  AN2        u0691(.A(men_men_n250_), .B(men_men_n87_), .Y(men_men_n714_));
  NA2        u0692(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n715_));
  NA3        u0693(.A(men_men_n509_), .B(men_men_n546_), .C(men_men_n47_), .Y(men_men_n716_));
  NO3        u0694(.A(men_men_n503_), .B(men_men_n637_), .C(men_men_n87_), .Y(men_men_n717_));
  NA2        u0695(.A(men_men_n717_), .B(men_men_n25_), .Y(men_men_n718_));
  NA3        u0696(.A(men_men_n162_), .B(men_men_n85_), .C(men_men_n87_), .Y(men_men_n719_));
  NA4        u0697(.A(men_men_n719_), .B(men_men_n718_), .C(men_men_n716_), .D(men_men_n715_), .Y(men_men_n720_));
  OAI210     u0698(.A0(men_men_n720_), .A1(men_men_n714_), .B0(i_1_), .Y(men_men_n721_));
  AOI210     u0699(.A0(men_men_n275_), .A1(men_men_n99_), .B0(i_1_), .Y(men_men_n722_));
  NO2        u0700(.A(men_men_n385_), .B(i_2_), .Y(men_men_n723_));
  NA2        u0701(.A(men_men_n723_), .B(men_men_n722_), .Y(men_men_n724_));
  OAI210     u0702(.A0(men_men_n686_), .A1(men_men_n470_), .B0(men_men_n724_), .Y(men_men_n725_));
  INV        u0703(.A(men_men_n725_), .Y(men_men_n726_));
  AOI210     u0704(.A0(men_men_n726_), .A1(men_men_n721_), .B0(i_13_), .Y(men_men_n727_));
  OR2        u0705(.A(i_11_), .B(i_7_), .Y(men_men_n728_));
  NA3        u0706(.A(men_men_n728_), .B(men_men_n108_), .C(men_men_n139_), .Y(men_men_n729_));
  AOI220     u0707(.A0(men_men_n495_), .A1(men_men_n162_), .B0(men_men_n472_), .B1(men_men_n139_), .Y(men_men_n730_));
  OAI210     u0708(.A0(men_men_n730_), .A1(men_men_n45_), .B0(men_men_n729_), .Y(men_men_n731_));
  AOI210     u0709(.A0(men_men_n683_), .A1(men_men_n55_), .B0(i_12_), .Y(men_men_n732_));
  INV        u0710(.A(men_men_n732_), .Y(men_men_n733_));
  NO2        u0711(.A(men_men_n503_), .B(men_men_n24_), .Y(men_men_n734_));
  AOI220     u0712(.A0(men_men_n734_), .A1(men_men_n701_), .B0(men_men_n250_), .B1(men_men_n132_), .Y(men_men_n735_));
  OAI220     u0713(.A0(men_men_n735_), .A1(men_men_n41_), .B0(men_men_n733_), .B1(men_men_n94_), .Y(men_men_n736_));
  AOI210     u0714(.A0(men_men_n731_), .A1(men_men_n343_), .B0(men_men_n736_), .Y(men_men_n737_));
  INV        u0715(.A(men_men_n117_), .Y(men_men_n738_));
  AOI220     u0716(.A0(men_men_n738_), .A1(men_men_n73_), .B0(men_men_n403_), .B1(men_men_n684_), .Y(men_men_n739_));
  NO2        u0717(.A(men_men_n739_), .B(men_men_n247_), .Y(men_men_n740_));
  AOI210     u0718(.A0(men_men_n470_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n741_));
  NOi31      u0719(.An(men_men_n741_), .B(men_men_n626_), .C(men_men_n45_), .Y(men_men_n742_));
  NA2        u0720(.A(men_men_n128_), .B(i_13_), .Y(men_men_n743_));
  NO2        u0721(.A(men_men_n683_), .B(men_men_n117_), .Y(men_men_n744_));
  INV        u0722(.A(men_men_n744_), .Y(men_men_n745_));
  OAI220     u0723(.A0(men_men_n745_), .A1(men_men_n72_), .B0(men_men_n743_), .B1(men_men_n722_), .Y(men_men_n746_));
  NA2        u0724(.A(men_men_n26_), .B(men_men_n196_), .Y(men_men_n747_));
  NA2        u0725(.A(men_men_n747_), .B(i_7_), .Y(men_men_n748_));
  NO3        u0726(.A(men_men_n503_), .B(men_men_n241_), .C(men_men_n87_), .Y(men_men_n749_));
  NA2        u0727(.A(men_men_n749_), .B(men_men_n748_), .Y(men_men_n750_));
  AOI220     u0728(.A0(men_men_n403_), .A1(men_men_n684_), .B0(men_men_n93_), .B1(men_men_n104_), .Y(men_men_n751_));
  OAI220     u0729(.A0(men_men_n751_), .A1(men_men_n632_), .B0(men_men_n750_), .B1(men_men_n647_), .Y(men_men_n752_));
  NO4        u0730(.A(men_men_n752_), .B(men_men_n746_), .C(men_men_n742_), .D(men_men_n740_), .Y(men_men_n753_));
  OR2        u0731(.A(i_11_), .B(i_6_), .Y(men_men_n754_));
  NA3        u0732(.A(men_men_n631_), .B(men_men_n747_), .C(i_7_), .Y(men_men_n755_));
  AOI210     u0733(.A0(men_men_n755_), .A1(men_men_n745_), .B0(men_men_n754_), .Y(men_men_n756_));
  NA3        u0734(.A(men_men_n429_), .B(men_men_n636_), .C(men_men_n99_), .Y(men_men_n757_));
  NA2        u0735(.A(men_men_n673_), .B(i_13_), .Y(men_men_n758_));
  NA2        u0736(.A(men_men_n104_), .B(men_men_n747_), .Y(men_men_n759_));
  NAi21      u0737(.An(i_11_), .B(i_12_), .Y(men_men_n760_));
  NOi41      u0738(.An(men_men_n113_), .B(men_men_n760_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n761_));
  NO3        u0739(.A(men_men_n503_), .B(men_men_n609_), .C(men_men_n637_), .Y(men_men_n762_));
  AOI220     u0740(.A0(men_men_n762_), .A1(men_men_n321_), .B0(men_men_n761_), .B1(men_men_n759_), .Y(men_men_n763_));
  NA3        u0741(.A(men_men_n763_), .B(men_men_n758_), .C(men_men_n757_), .Y(men_men_n764_));
  OAI210     u0742(.A0(men_men_n764_), .A1(men_men_n756_), .B0(men_men_n64_), .Y(men_men_n765_));
  NO2        u0743(.A(i_2_), .B(i_12_), .Y(men_men_n766_));
  NA2        u0744(.A(men_men_n384_), .B(men_men_n766_), .Y(men_men_n767_));
  NA2        u0745(.A(i_8_), .B(men_men_n25_), .Y(men_men_n768_));
  NO3        u0746(.A(men_men_n768_), .B(men_men_n401_), .C(men_men_n631_), .Y(men_men_n769_));
  OAI210     u0747(.A0(men_men_n769_), .A1(men_men_n386_), .B0(men_men_n384_), .Y(men_men_n770_));
  NO2        u0748(.A(men_men_n129_), .B(i_2_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n771_), .B(men_men_n667_), .Y(men_men_n772_));
  NA3        u0750(.A(men_men_n772_), .B(men_men_n770_), .C(men_men_n767_), .Y(men_men_n773_));
  NA3        u0751(.A(men_men_n773_), .B(men_men_n46_), .C(men_men_n229_), .Y(men_men_n774_));
  NA4        u0752(.A(men_men_n774_), .B(men_men_n765_), .C(men_men_n753_), .D(men_men_n737_), .Y(men_men_n775_));
  OR4        u0753(.A(men_men_n775_), .B(men_men_n727_), .C(men_men_n713_), .D(men_men_n650_), .Y(men5));
  NA2        u0754(.A(men_men_n698_), .B(men_men_n278_), .Y(men_men_n777_));
  AN2        u0755(.A(men_men_n24_), .B(i_10_), .Y(men_men_n778_));
  NA3        u0756(.A(men_men_n778_), .B(men_men_n766_), .C(men_men_n110_), .Y(men_men_n779_));
  NO2        u0757(.A(men_men_n632_), .B(i_11_), .Y(men_men_n780_));
  NA2        u0758(.A(men_men_n88_), .B(men_men_n780_), .Y(men_men_n781_));
  NA3        u0759(.A(men_men_n781_), .B(men_men_n779_), .C(men_men_n777_), .Y(men_men_n782_));
  NO3        u0760(.A(i_11_), .B(men_men_n241_), .C(i_13_), .Y(men_men_n783_));
  NO2        u0761(.A(men_men_n125_), .B(men_men_n23_), .Y(men_men_n784_));
  NA2        u0762(.A(i_12_), .B(i_8_), .Y(men_men_n785_));
  OAI210     u0763(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n785_), .Y(men_men_n786_));
  INV        u0764(.A(men_men_n469_), .Y(men_men_n787_));
  AOI220     u0765(.A0(men_men_n327_), .A1(men_men_n603_), .B0(men_men_n786_), .B1(men_men_n784_), .Y(men_men_n788_));
  INV        u0766(.A(men_men_n788_), .Y(men_men_n789_));
  NO2        u0767(.A(men_men_n789_), .B(men_men_n782_), .Y(men_men_n790_));
  INV        u0768(.A(men_men_n173_), .Y(men_men_n791_));
  INV        u0769(.A(men_men_n250_), .Y(men_men_n792_));
  OAI210     u0770(.A0(men_men_n723_), .A1(men_men_n471_), .B0(men_men_n113_), .Y(men_men_n793_));
  AOI210     u0771(.A0(men_men_n793_), .A1(men_men_n792_), .B0(men_men_n791_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n477_), .B(men_men_n26_), .Y(men_men_n795_));
  NO2        u0773(.A(men_men_n795_), .B(men_men_n440_), .Y(men_men_n796_));
  NA2        u0774(.A(men_men_n796_), .B(i_2_), .Y(men_men_n797_));
  INV        u0775(.A(men_men_n797_), .Y(men_men_n798_));
  AOI210     u0776(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n436_), .Y(men_men_n799_));
  AOI210     u0777(.A0(men_men_n799_), .A1(men_men_n798_), .B0(men_men_n794_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n193_), .B(men_men_n126_), .Y(men_men_n801_));
  OAI210     u0779(.A0(men_men_n801_), .A1(men_men_n784_), .B0(i_2_), .Y(men_men_n802_));
  INV        u0780(.A(men_men_n174_), .Y(men_men_n803_));
  NO3        u0781(.A(men_men_n652_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n804_));
  AOI210     u0782(.A0(men_men_n803_), .A1(men_men_n88_), .B0(men_men_n804_), .Y(men_men_n805_));
  AOI210     u0783(.A0(men_men_n805_), .A1(men_men_n802_), .B0(men_men_n196_), .Y(men_men_n806_));
  OA210      u0784(.A0(men_men_n653_), .A1(men_men_n127_), .B0(i_13_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n203_), .B(men_men_n206_), .Y(men_men_n808_));
  NA2        u0786(.A(men_men_n152_), .B(men_men_n627_), .Y(men_men_n809_));
  AOI210     u0787(.A0(men_men_n809_), .A1(men_men_n808_), .B0(men_men_n389_), .Y(men_men_n810_));
  AOI210     u0788(.A0(men_men_n211_), .A1(men_men_n149_), .B0(men_men_n546_), .Y(men_men_n811_));
  NA2        u0789(.A(men_men_n811_), .B(men_men_n440_), .Y(men_men_n812_));
  NO2        u0790(.A(men_men_n104_), .B(men_men_n45_), .Y(men_men_n813_));
  INV        u0791(.A(men_men_n310_), .Y(men_men_n814_));
  NA4        u0792(.A(men_men_n814_), .B(men_men_n314_), .C(men_men_n125_), .D(men_men_n43_), .Y(men_men_n815_));
  OAI210     u0793(.A0(men_men_n815_), .A1(men_men_n813_), .B0(men_men_n812_), .Y(men_men_n816_));
  NO4        u0794(.A(men_men_n816_), .B(men_men_n810_), .C(men_men_n807_), .D(men_men_n806_), .Y(men_men_n817_));
  NA2        u0795(.A(men_men_n603_), .B(men_men_n28_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n783_), .B(men_men_n282_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n819_), .B(men_men_n818_), .Y(men_men_n820_));
  NO2        u0798(.A(men_men_n63_), .B(i_12_), .Y(men_men_n821_));
  NO2        u0799(.A(men_men_n821_), .B(men_men_n127_), .Y(men_men_n822_));
  NO2        u0800(.A(men_men_n822_), .B(men_men_n627_), .Y(men_men_n823_));
  AOI220     u0801(.A0(men_men_n823_), .A1(men_men_n36_), .B0(men_men_n820_), .B1(men_men_n47_), .Y(men_men_n824_));
  NA4        u0802(.A(men_men_n824_), .B(men_men_n817_), .C(men_men_n800_), .D(men_men_n790_), .Y(men6));
  NO3        u0803(.A(men_men_n261_), .B(men_men_n316_), .C(i_1_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n188_), .B(men_men_n140_), .Y(men_men_n827_));
  OAI210     u0805(.A0(men_men_n827_), .A1(men_men_n826_), .B0(men_men_n771_), .Y(men_men_n828_));
  NA4        u0806(.A(men_men_n407_), .B(men_men_n508_), .C(men_men_n72_), .D(men_men_n103_), .Y(men_men_n829_));
  INV        u0807(.A(men_men_n829_), .Y(men_men_n830_));
  NO2        u0808(.A(men_men_n224_), .B(men_men_n513_), .Y(men_men_n831_));
  NO2        u0809(.A(i_11_), .B(i_9_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n830_), .B(men_men_n339_), .Y(men_men_n833_));
  AO210      u0811(.A0(men_men_n833_), .A1(men_men_n828_), .B0(i_12_), .Y(men_men_n834_));
  NA2        u0812(.A(men_men_n390_), .B(men_men_n346_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n609_), .B(men_men_n64_), .Y(men_men_n836_));
  NA2        u0814(.A(men_men_n836_), .B(men_men_n835_), .Y(men_men_n837_));
  INV        u0815(.A(men_men_n200_), .Y(men_men_n838_));
  AOI220     u0816(.A0(men_men_n838_), .A1(men_men_n832_), .B0(men_men_n837_), .B1(men_men_n74_), .Y(men_men_n839_));
  INV        u0817(.A(men_men_n338_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n76_), .B(men_men_n132_), .Y(men_men_n841_));
  INV        u0819(.A(men_men_n125_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n842_), .B(men_men_n47_), .Y(men_men_n843_));
  AOI210     u0821(.A0(men_men_n843_), .A1(men_men_n841_), .B0(men_men_n840_), .Y(men_men_n844_));
  NO3        u0822(.A(men_men_n257_), .B(men_men_n133_), .C(i_9_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n845_), .B(men_men_n821_), .Y(men_men_n846_));
  AOI210     u0824(.A0(men_men_n846_), .A1(men_men_n544_), .B0(men_men_n188_), .Y(men_men_n847_));
  NAi32      u0825(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n848_));
  NO2        u0826(.A(men_men_n754_), .B(men_men_n848_), .Y(men_men_n849_));
  OR3        u0827(.A(men_men_n849_), .B(men_men_n847_), .C(men_men_n844_), .Y(men_men_n850_));
  NO2        u0828(.A(men_men_n728_), .B(i_2_), .Y(men_men_n851_));
  NA2        u0829(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n852_));
  NO2        u0830(.A(men_men_n852_), .B(men_men_n428_), .Y(men_men_n853_));
  NA2        u0831(.A(men_men_n853_), .B(men_men_n851_), .Y(men_men_n854_));
  AO220      u0832(.A0(men_men_n374_), .A1(men_men_n364_), .B0(men_men_n415_), .B1(men_men_n627_), .Y(men_men_n855_));
  NA3        u0833(.A(men_men_n855_), .B(men_men_n262_), .C(i_7_), .Y(men_men_n856_));
  OR2        u0834(.A(men_men_n653_), .B(men_men_n471_), .Y(men_men_n857_));
  NA3        u0835(.A(men_men_n857_), .B(men_men_n148_), .C(men_men_n70_), .Y(men_men_n858_));
  AO210      u0836(.A0(men_men_n520_), .A1(men_men_n787_), .B0(men_men_n36_), .Y(men_men_n859_));
  NA4        u0837(.A(men_men_n859_), .B(men_men_n858_), .C(men_men_n856_), .D(men_men_n854_), .Y(men_men_n860_));
  NO2        u0838(.A(men_men_n672_), .B(i_11_), .Y(men_men_n861_));
  AOI220     u0839(.A0(men_men_n861_), .A1(men_men_n593_), .B0(men_men_n831_), .B1(men_men_n748_), .Y(men_men_n862_));
  NA3        u0840(.A(men_men_n389_), .B(men_men_n243_), .C(men_men_n148_), .Y(men_men_n863_));
  NA2        u0841(.A(men_men_n415_), .B(men_men_n71_), .Y(men_men_n864_));
  NA4        u0842(.A(men_men_n864_), .B(men_men_n863_), .C(men_men_n862_), .D(men_men_n635_), .Y(men_men_n865_));
  AOI210     u0843(.A0(men_men_n471_), .A1(men_men_n469_), .B0(men_men_n592_), .Y(men_men_n866_));
  NO2        u0844(.A(men_men_n643_), .B(men_men_n104_), .Y(men_men_n867_));
  OAI210     u0845(.A0(men_men_n867_), .A1(men_men_n114_), .B0(men_men_n426_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n249_), .B(men_men_n47_), .Y(men_men_n869_));
  INV        u0847(.A(men_men_n616_), .Y(men_men_n870_));
  NA3        u0848(.A(men_men_n870_), .B(men_men_n338_), .C(i_7_), .Y(men_men_n871_));
  NA3        u0849(.A(men_men_n871_), .B(men_men_n868_), .C(men_men_n866_), .Y(men_men_n872_));
  NO4        u0850(.A(men_men_n872_), .B(men_men_n865_), .C(men_men_n860_), .D(men_men_n850_), .Y(men_men_n873_));
  NA4        u0851(.A(men_men_n873_), .B(men_men_n839_), .C(men_men_n834_), .D(men_men_n397_), .Y(men3));
  NA2        u0852(.A(i_12_), .B(i_10_), .Y(men_men_n875_));
  NA2        u0853(.A(i_6_), .B(i_7_), .Y(men_men_n876_));
  NO2        u0854(.A(men_men_n876_), .B(i_0_), .Y(men_men_n877_));
  NO2        u0855(.A(i_11_), .B(men_men_n241_), .Y(men_men_n878_));
  OAI210     u0856(.A0(men_men_n877_), .A1(men_men_n298_), .B0(men_men_n878_), .Y(men_men_n879_));
  NO2        u0857(.A(men_men_n879_), .B(men_men_n196_), .Y(men_men_n880_));
  NO3        u0858(.A(men_men_n473_), .B(men_men_n91_), .C(men_men_n45_), .Y(men_men_n881_));
  OA210      u0859(.A0(men_men_n881_), .A1(men_men_n880_), .B0(men_men_n176_), .Y(men_men_n882_));
  NA2        u0860(.A(men_men_n863_), .B(men_men_n388_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n883_), .B(men_men_n40_), .Y(men_men_n884_));
  NOi21      u0862(.An(men_men_n98_), .B(men_men_n796_), .Y(men_men_n885_));
  NO3        u0863(.A(men_men_n662_), .B(men_men_n477_), .C(men_men_n132_), .Y(men_men_n886_));
  NA2        u0864(.A(men_men_n429_), .B(men_men_n46_), .Y(men_men_n887_));
  AN2        u0865(.A(men_men_n475_), .B(men_men_n56_), .Y(men_men_n888_));
  NO3        u0866(.A(men_men_n888_), .B(men_men_n886_), .C(men_men_n885_), .Y(men_men_n889_));
  AOI210     u0867(.A0(men_men_n889_), .A1(men_men_n884_), .B0(men_men_n49_), .Y(men_men_n890_));
  NO4        u0868(.A(men_men_n393_), .B(men_men_n400_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n188_), .B(men_men_n601_), .Y(men_men_n892_));
  NOi21      u0870(.An(men_men_n892_), .B(men_men_n891_), .Y(men_men_n893_));
  NA2        u0871(.A(men_men_n741_), .B(men_men_n707_), .Y(men_men_n894_));
  NA2        u0872(.A(men_men_n344_), .B(men_men_n460_), .Y(men_men_n895_));
  OAI220     u0873(.A0(men_men_n895_), .A1(men_men_n894_), .B0(men_men_n893_), .B1(men_men_n64_), .Y(men_men_n896_));
  NOi21      u0874(.An(i_5_), .B(i_9_), .Y(men_men_n897_));
  NA2        u0875(.A(men_men_n897_), .B(men_men_n468_), .Y(men_men_n898_));
  BUFFER     u0876(.A(men_men_n275_), .Y(men_men_n899_));
  AOI210     u0877(.A0(men_men_n899_), .A1(men_men_n500_), .B0(men_men_n717_), .Y(men_men_n900_));
  NO2        u0878(.A(men_men_n177_), .B(men_men_n149_), .Y(men_men_n901_));
  NO2        u0879(.A(men_men_n900_), .B(men_men_n898_), .Y(men_men_n902_));
  NO4        u0880(.A(men_men_n902_), .B(men_men_n896_), .C(men_men_n890_), .D(men_men_n882_), .Y(men_men_n903_));
  NA2        u0881(.A(men_men_n188_), .B(men_men_n24_), .Y(men_men_n904_));
  NA2        u0882(.A(men_men_n321_), .B(men_men_n130_), .Y(men_men_n905_));
  NAi21      u0883(.An(men_men_n163_), .B(men_men_n460_), .Y(men_men_n906_));
  OAI220     u0884(.A0(men_men_n906_), .A1(men_men_n869_), .B0(men_men_n905_), .B1(men_men_n418_), .Y(men_men_n907_));
  INV        u0885(.A(men_men_n907_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n407_), .B(men_men_n302_), .Y(men_men_n909_));
  NA2        u0887(.A(men_men_n909_), .B(men_men_n744_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n602_), .B(i_0_), .Y(men_men_n911_));
  NO4        u0889(.A(men_men_n615_), .B(men_men_n218_), .C(men_men_n436_), .D(men_men_n428_), .Y(men_men_n912_));
  NA2        u0890(.A(men_men_n912_), .B(i_11_), .Y(men_men_n913_));
  INV        u0891(.A(men_men_n498_), .Y(men_men_n914_));
  AN2        u0892(.A(men_men_n98_), .B(men_men_n248_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n783_), .B(men_men_n339_), .Y(men_men_n916_));
  AOI210     u0894(.A0(men_men_n509_), .A1(men_men_n88_), .B0(men_men_n59_), .Y(men_men_n917_));
  OAI220     u0895(.A0(men_men_n917_), .A1(men_men_n916_), .B0(men_men_n693_), .B1(men_men_n569_), .Y(men_men_n918_));
  NO2        u0896(.A(men_men_n259_), .B(men_men_n154_), .Y(men_men_n919_));
  NA2        u0897(.A(i_0_), .B(i_10_), .Y(men_men_n920_));
  AN2        u0898(.A(men_men_n919_), .B(i_6_), .Y(men_men_n921_));
  AOI220     u0899(.A0(men_men_n344_), .A1(men_men_n100_), .B0(men_men_n188_), .B1(men_men_n85_), .Y(men_men_n922_));
  NA2        u0900(.A(men_men_n597_), .B(i_4_), .Y(men_men_n923_));
  NO2        u0901(.A(men_men_n923_), .B(men_men_n922_), .Y(men_men_n924_));
  NO4        u0902(.A(men_men_n924_), .B(men_men_n921_), .C(men_men_n918_), .D(men_men_n915_), .Y(men_men_n925_));
  NA4        u0903(.A(men_men_n925_), .B(men_men_n913_), .C(men_men_n910_), .D(men_men_n908_), .Y(men_men_n926_));
  NA2        u0904(.A(i_11_), .B(i_9_), .Y(men_men_n927_));
  NO2        u0905(.A(men_men_n49_), .B(i_7_), .Y(men_men_n928_));
  NA2        u0906(.A(men_men_n412_), .B(men_men_n181_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n929_), .B(men_men_n161_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n927_), .B(men_men_n74_), .Y(men_men_n931_));
  NO2        u0909(.A(men_men_n177_), .B(i_0_), .Y(men_men_n932_));
  INV        u0910(.A(men_men_n932_), .Y(men_men_n933_));
  NA2        u0911(.A(men_men_n498_), .B(men_men_n235_), .Y(men_men_n934_));
  AOI210     u0912(.A0(men_men_n387_), .A1(men_men_n42_), .B0(men_men_n425_), .Y(men_men_n935_));
  OAI220     u0913(.A0(men_men_n935_), .A1(men_men_n898_), .B0(men_men_n934_), .B1(men_men_n933_), .Y(men_men_n936_));
  NO2        u0914(.A(men_men_n936_), .B(men_men_n930_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n692_), .B(men_men_n122_), .Y(men_men_n938_));
  NO2        u0916(.A(i_6_), .B(men_men_n938_), .Y(men_men_n939_));
  AOI210     u0917(.A0(men_men_n470_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n173_), .B(men_men_n105_), .Y(men_men_n941_));
  NOi32      u0919(.An(men_men_n940_), .Bn(men_men_n191_), .C(men_men_n941_), .Y(men_men_n942_));
  NA2        u0920(.A(men_men_n636_), .B(men_men_n339_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n943_), .B(men_men_n887_), .Y(men_men_n944_));
  NO3        u0922(.A(men_men_n944_), .B(men_men_n942_), .C(men_men_n939_), .Y(men_men_n945_));
  NOi21      u0923(.An(i_7_), .B(i_5_), .Y(men_men_n946_));
  NOi31      u0924(.An(men_men_n946_), .B(i_0_), .C(men_men_n760_), .Y(men_men_n947_));
  NA3        u0925(.A(men_men_n947_), .B(men_men_n401_), .C(i_6_), .Y(men_men_n948_));
  OA210      u0926(.A0(men_men_n941_), .A1(men_men_n544_), .B0(men_men_n948_), .Y(men_men_n949_));
  NO3        u0927(.A(men_men_n421_), .B(men_men_n377_), .C(men_men_n373_), .Y(men_men_n950_));
  NO2        u0928(.A(men_men_n269_), .B(men_men_n328_), .Y(men_men_n951_));
  NO2        u0929(.A(men_men_n760_), .B(men_men_n264_), .Y(men_men_n952_));
  AOI210     u0930(.A0(men_men_n952_), .A1(men_men_n951_), .B0(men_men_n950_), .Y(men_men_n953_));
  NA4        u0931(.A(men_men_n953_), .B(men_men_n949_), .C(men_men_n945_), .D(men_men_n937_), .Y(men_men_n954_));
  NO2        u0932(.A(men_men_n904_), .B(men_men_n244_), .Y(men_men_n955_));
  AN2        u0933(.A(men_men_n343_), .B(men_men_n339_), .Y(men_men_n956_));
  AN2        u0934(.A(men_men_n956_), .B(men_men_n901_), .Y(men_men_n957_));
  OAI210     u0935(.A0(men_men_n957_), .A1(men_men_n955_), .B0(i_10_), .Y(men_men_n958_));
  NO2        u0936(.A(men_men_n875_), .B(men_men_n327_), .Y(men_men_n959_));
  NA2        u0937(.A(men_men_n959_), .B(men_men_n931_), .Y(men_men_n960_));
  NA3        u0938(.A(men_men_n497_), .B(men_men_n429_), .C(men_men_n46_), .Y(men_men_n961_));
  OAI210     u0939(.A0(men_men_n906_), .A1(men_men_n914_), .B0(men_men_n961_), .Y(men_men_n962_));
  NO2        u0940(.A(men_men_n262_), .B(men_men_n47_), .Y(men_men_n963_));
  NA2        u0941(.A(men_men_n931_), .B(men_men_n314_), .Y(men_men_n964_));
  OAI210     u0942(.A0(men_men_n963_), .A1(men_men_n190_), .B0(men_men_n964_), .Y(men_men_n965_));
  AOI220     u0943(.A0(men_men_n965_), .A1(men_men_n498_), .B0(men_men_n962_), .B1(men_men_n74_), .Y(men_men_n966_));
  NA3        u0944(.A(men_men_n852_), .B(men_men_n399_), .C(men_men_n672_), .Y(men_men_n967_));
  NO2        u0945(.A(men_men_n967_), .B(men_men_n48_), .Y(men_men_n968_));
  NO3        u0946(.A(men_men_n615_), .B(men_men_n372_), .C(men_men_n24_), .Y(men_men_n969_));
  AOI210     u0947(.A0(men_men_n734_), .A1(men_men_n576_), .B0(men_men_n969_), .Y(men_men_n970_));
  NAi21      u0948(.An(i_9_), .B(i_5_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n971_), .B(men_men_n421_), .Y(men_men_n972_));
  NO2        u0950(.A(men_men_n630_), .B(men_men_n107_), .Y(men_men_n973_));
  AOI220     u0951(.A0(men_men_n973_), .A1(i_0_), .B0(men_men_n972_), .B1(men_men_n653_), .Y(men_men_n974_));
  OAI220     u0952(.A0(men_men_n974_), .A1(men_men_n87_), .B0(men_men_n970_), .B1(men_men_n174_), .Y(men_men_n975_));
  NO3        u0953(.A(men_men_n975_), .B(men_men_n968_), .C(men_men_n549_), .Y(men_men_n976_));
  NA4        u0954(.A(men_men_n976_), .B(men_men_n966_), .C(men_men_n960_), .D(men_men_n958_), .Y(men_men_n977_));
  NO3        u0955(.A(men_men_n977_), .B(men_men_n954_), .C(men_men_n926_), .Y(men_men_n978_));
  NO2        u0956(.A(i_0_), .B(men_men_n760_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n74_), .B(men_men_n45_), .Y(men_men_n980_));
  NA2        u0958(.A(men_men_n920_), .B(men_men_n980_), .Y(men_men_n981_));
  NO3        u0959(.A(men_men_n107_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n982_));
  AO220      u0960(.A0(men_men_n982_), .A1(men_men_n981_), .B0(men_men_n979_), .B1(men_men_n176_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n836_), .A1(men_men_n715_), .B0(men_men_n941_), .Y(men_men_n984_));
  AOI210     u0962(.A0(men_men_n983_), .A1(men_men_n361_), .B0(men_men_n984_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n771_), .B(men_men_n147_), .Y(men_men_n986_));
  INV        u0964(.A(men_men_n986_), .Y(men_men_n987_));
  NA3        u0965(.A(men_men_n987_), .B(men_men_n707_), .C(men_men_n74_), .Y(men_men_n988_));
  NA3        u0966(.A(men_men_n877_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n989_));
  NA2        u0967(.A(men_men_n878_), .B(i_9_), .Y(men_men_n990_));
  AOI210     u0968(.A0(men_men_n989_), .A1(men_men_n525_), .B0(men_men_n990_), .Y(men_men_n991_));
  OAI210     u0969(.A0(men_men_n249_), .A1(i_9_), .B0(men_men_n234_), .Y(men_men_n992_));
  AOI210     u0970(.A0(men_men_n992_), .A1(men_men_n911_), .B0(men_men_n154_), .Y(men_men_n993_));
  NO2        u0971(.A(men_men_n993_), .B(men_men_n991_), .Y(men_men_n994_));
  NA3        u0972(.A(men_men_n994_), .B(men_men_n988_), .C(men_men_n985_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n956_), .B(men_men_n389_), .Y(men_men_n996_));
  AOI210     u0974(.A0(men_men_n309_), .A1(men_men_n163_), .B0(men_men_n996_), .Y(men_men_n997_));
  NA3        u0975(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n998_));
  NA2        u0976(.A(men_men_n928_), .B(men_men_n514_), .Y(men_men_n999_));
  AOI210     u0977(.A0(men_men_n998_), .A1(men_men_n163_), .B0(men_men_n999_), .Y(men_men_n1000_));
  NO2        u0978(.A(men_men_n1000_), .B(men_men_n997_), .Y(men_men_n1001_));
  NO3        u0979(.A(men_men_n920_), .B(men_men_n897_), .C(men_men_n193_), .Y(men_men_n1002_));
  AOI220     u0980(.A0(men_men_n1002_), .A1(i_11_), .B0(men_men_n598_), .B1(men_men_n76_), .Y(men_men_n1003_));
  NO3        u0981(.A(men_men_n212_), .B(men_men_n400_), .C(i_0_), .Y(men_men_n1004_));
  OAI210     u0982(.A0(men_men_n1004_), .A1(men_men_n77_), .B0(i_13_), .Y(men_men_n1005_));
  INV        u0983(.A(men_men_n221_), .Y(men_men_n1006_));
  OAI220     u0984(.A0(men_men_n562_), .A1(men_men_n140_), .B0(men_men_n677_), .B1(men_men_n647_), .Y(men_men_n1007_));
  NA3        u0985(.A(men_men_n1007_), .B(men_men_n416_), .C(men_men_n1006_), .Y(men_men_n1008_));
  NA4        u0986(.A(men_men_n1008_), .B(men_men_n1005_), .C(men_men_n1003_), .D(men_men_n1001_), .Y(men_men_n1009_));
  INV        u0987(.A(men_men_n111_), .Y(men_men_n1010_));
  AOI220     u0988(.A0(men_men_n946_), .A1(men_men_n514_), .B0(men_men_n877_), .B1(men_men_n164_), .Y(men_men_n1011_));
  NA2        u0989(.A(men_men_n364_), .B(men_men_n178_), .Y(men_men_n1012_));
  OA220      u0990(.A0(men_men_n1012_), .A1(men_men_n1011_), .B0(men_men_n1010_), .B1(i_5_), .Y(men_men_n1013_));
  NA3        u0991(.A(men_men_n644_), .B(men_men_n188_), .C(men_men_n85_), .Y(men_men_n1014_));
  INV        u0992(.A(men_men_n1014_), .Y(men_men_n1015_));
  NO3        u0993(.A(men_men_n887_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n1016_));
  NA2        u0994(.A(men_men_n519_), .B(men_men_n512_), .Y(men_men_n1017_));
  NO3        u0995(.A(men_men_n1017_), .B(men_men_n1016_), .C(men_men_n1015_), .Y(men_men_n1018_));
  NA3        u0996(.A(men_men_n407_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n1019_));
  NA3        u0997(.A(men_men_n928_), .B(men_men_n298_), .C(men_men_n234_), .Y(men_men_n1020_));
  NA2        u0998(.A(men_men_n1020_), .B(men_men_n1019_), .Y(men_men_n1021_));
  NA3        u0999(.A(men_men_n407_), .B(men_men_n345_), .C(men_men_n225_), .Y(men_men_n1022_));
  INV        u1000(.A(men_men_n1022_), .Y(men_men_n1023_));
  NOi31      u1001(.An(men_men_n406_), .B(men_men_n980_), .C(men_men_n244_), .Y(men_men_n1024_));
  NO3        u1002(.A(men_men_n927_), .B(men_men_n221_), .C(men_men_n193_), .Y(men_men_n1025_));
  NO4        u1003(.A(men_men_n1025_), .B(men_men_n1024_), .C(men_men_n1023_), .D(men_men_n1021_), .Y(men_men_n1026_));
  NA3        u1004(.A(men_men_n1026_), .B(men_men_n1018_), .C(men_men_n1013_), .Y(men_men_n1027_));
  INV        u1005(.A(men_men_n646_), .Y(men_men_n1028_));
  NO3        u1006(.A(men_men_n1028_), .B(men_men_n588_), .C(men_men_n358_), .Y(men_men_n1029_));
  NO2        u1007(.A(men_men_n87_), .B(i_5_), .Y(men_men_n1030_));
  NA3        u1008(.A(men_men_n878_), .B(men_men_n112_), .C(men_men_n125_), .Y(men_men_n1031_));
  INV        u1009(.A(men_men_n1031_), .Y(men_men_n1032_));
  AOI210     u1010(.A0(men_men_n1032_), .A1(men_men_n1030_), .B0(men_men_n1029_), .Y(men_men_n1033_));
  NAi21      u1011(.An(men_men_n246_), .B(men_men_n247_), .Y(men_men_n1034_));
  NO4        u1012(.A(men_men_n244_), .B(men_men_n212_), .C(i_0_), .D(i_12_), .Y(men_men_n1035_));
  AOI220     u1013(.A0(men_men_n1035_), .A1(men_men_n1034_), .B0(men_men_n830_), .B1(men_men_n178_), .Y(men_men_n1036_));
  AN2        u1014(.A(men_men_n920_), .B(men_men_n154_), .Y(men_men_n1037_));
  NO4        u1015(.A(men_men_n1037_), .B(i_12_), .C(men_men_n681_), .D(men_men_n132_), .Y(men_men_n1038_));
  NA2        u1016(.A(men_men_n1038_), .B(men_men_n221_), .Y(men_men_n1039_));
  NA3        u1017(.A(men_men_n100_), .B(men_men_n601_), .C(i_11_), .Y(men_men_n1040_));
  NO2        u1018(.A(men_men_n1040_), .B(men_men_n156_), .Y(men_men_n1041_));
  NA2        u1019(.A(men_men_n946_), .B(men_men_n495_), .Y(men_men_n1042_));
  NO2        u1020(.A(men_men_n1042_), .B(men_men_n708_), .Y(men_men_n1043_));
  AOI210     u1021(.A0(men_men_n1043_), .A1(men_men_n932_), .B0(men_men_n1041_), .Y(men_men_n1044_));
  NA4        u1022(.A(men_men_n1044_), .B(men_men_n1039_), .C(men_men_n1036_), .D(men_men_n1033_), .Y(men_men_n1045_));
  NO4        u1023(.A(men_men_n1045_), .B(men_men_n1027_), .C(men_men_n1009_), .D(men_men_n995_), .Y(men_men_n1046_));
  NA2        u1024(.A(men_men_n851_), .B(men_men_n37_), .Y(men_men_n1047_));
  NA3        u1025(.A(men_men_n940_), .B(men_men_n384_), .C(i_5_), .Y(men_men_n1048_));
  NA3        u1026(.A(men_men_n1048_), .B(men_men_n1047_), .C(men_men_n642_), .Y(men_men_n1049_));
  NA2        u1027(.A(men_men_n1049_), .B(men_men_n209_), .Y(men_men_n1050_));
  AN2        u1028(.A(men_men_n728_), .B(men_men_n385_), .Y(men_men_n1051_));
  NA2        u1029(.A(men_men_n189_), .B(men_men_n191_), .Y(men_men_n1052_));
  AO210      u1030(.A0(men_men_n1051_), .A1(men_men_n33_), .B0(men_men_n1052_), .Y(men_men_n1053_));
  OAI210     u1031(.A0(men_men_n646_), .A1(men_men_n644_), .B0(men_men_n327_), .Y(men_men_n1054_));
  NAi31      u1032(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1055_));
  NO2        u1033(.A(men_men_n71_), .B(men_men_n1055_), .Y(men_men_n1056_));
  NO2        u1034(.A(men_men_n1056_), .B(men_men_n678_), .Y(men_men_n1057_));
  NA3        u1035(.A(men_men_n1057_), .B(men_men_n1054_), .C(men_men_n1053_), .Y(men_men_n1058_));
  NO4        u1036(.A(men_men_n237_), .B(men_men_n146_), .C(men_men_n711_), .D(men_men_n37_), .Y(men_men_n1059_));
  NO2        u1037(.A(men_men_n1059_), .B(men_men_n912_), .Y(men_men_n1060_));
  OAI210     u1038(.A0(men_men_n1040_), .A1(men_men_n149_), .B0(men_men_n1060_), .Y(men_men_n1061_));
  AOI210     u1039(.A0(men_men_n1058_), .A1(men_men_n49_), .B0(men_men_n1061_), .Y(men_men_n1062_));
  AOI210     u1040(.A0(men_men_n1062_), .A1(men_men_n1050_), .B0(men_men_n74_), .Y(men_men_n1063_));
  NO2        u1041(.A(men_men_n595_), .B(men_men_n396_), .Y(men_men_n1064_));
  NO2        u1042(.A(men_men_n1064_), .B(men_men_n791_), .Y(men_men_n1065_));
  OAI210     u1043(.A0(men_men_n81_), .A1(men_men_n55_), .B0(men_men_n110_), .Y(men_men_n1066_));
  NA2        u1044(.A(men_men_n1066_), .B(men_men_n77_), .Y(men_men_n1067_));
  INV        u1045(.A(men_men_n947_), .Y(men_men_n1068_));
  AOI210     u1046(.A0(men_men_n1068_), .A1(men_men_n1067_), .B0(men_men_n711_), .Y(men_men_n1069_));
  NA2        u1047(.A(men_men_n269_), .B(men_men_n58_), .Y(men_men_n1070_));
  AOI220     u1048(.A0(men_men_n1070_), .A1(men_men_n77_), .B0(men_men_n359_), .B1(men_men_n261_), .Y(men_men_n1071_));
  NO2        u1049(.A(men_men_n1071_), .B(men_men_n241_), .Y(men_men_n1072_));
  NA3        u1050(.A(men_men_n98_), .B(men_men_n316_), .C(men_men_n31_), .Y(men_men_n1073_));
  INV        u1051(.A(men_men_n1073_), .Y(men_men_n1074_));
  NO3        u1052(.A(men_men_n1074_), .B(men_men_n1072_), .C(men_men_n1069_), .Y(men_men_n1075_));
  OAI210     u1053(.A0(men_men_n277_), .A1(men_men_n159_), .B0(men_men_n88_), .Y(men_men_n1076_));
  NA3        u1054(.A(men_men_n795_), .B(men_men_n298_), .C(men_men_n81_), .Y(men_men_n1077_));
  AOI210     u1055(.A0(men_men_n1077_), .A1(men_men_n1076_), .B0(i_11_), .Y(men_men_n1078_));
  NA2        u1056(.A(men_men_n637_), .B(men_men_n218_), .Y(men_men_n1079_));
  OAI210     u1057(.A0(men_men_n1079_), .A1(men_men_n940_), .B0(men_men_n209_), .Y(men_men_n1080_));
  NA2        u1058(.A(men_men_n165_), .B(i_5_), .Y(men_men_n1081_));
  NO2        u1059(.A(men_men_n1080_), .B(men_men_n1081_), .Y(men_men_n1082_));
  NO4        u1060(.A(men_men_n971_), .B(men_men_n502_), .C(men_men_n258_), .D(men_men_n257_), .Y(men_men_n1083_));
  NO2        u1061(.A(men_men_n1083_), .B(men_men_n592_), .Y(men_men_n1084_));
  NO2        u1062(.A(men_men_n1084_), .B(men_men_n41_), .Y(men_men_n1085_));
  NO3        u1063(.A(men_men_n1085_), .B(men_men_n1082_), .C(men_men_n1078_), .Y(men_men_n1086_));
  OAI210     u1064(.A0(men_men_n1075_), .A1(i_4_), .B0(men_men_n1086_), .Y(men_men_n1087_));
  NO3        u1065(.A(men_men_n1087_), .B(men_men_n1065_), .C(men_men_n1063_), .Y(men_men_n1088_));
  NA4        u1066(.A(men_men_n1088_), .B(men_men_n1046_), .C(men_men_n978_), .D(men_men_n903_), .Y(men4));
  INV        u1067(.A(i_2_), .Y(men_men_n1092_));
  INV        u1068(.A(men_men_n119_), .Y(men_men_n1093_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule