//Benchmark atmr_alu4_1266_0.125

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n130_, ori_ori_n131_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n621_, ori_ori_n622_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  INV        o019(.A(ori_ori_n35_), .Y(ori1));
  INV        o020(.A(i_11_), .Y(ori_ori_n43_));
  NO2        o021(.A(ori_ori_n43_), .B(i_6_), .Y(ori_ori_n44_));
  INV        o022(.A(i_2_), .Y(ori_ori_n45_));
  NA2        o023(.A(i_0_), .B(i_3_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  NO2        o027(.A(i_5_), .B(ori_ori_n45_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_0_), .B(i_2_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NA2        o031(.A(ori_ori_n50_), .B(ori_ori_n44_), .Y(ori_ori_n54_));
  NA3        o032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n55_));
  NO2        o033(.A(i_1_), .B(i_6_), .Y(ori_ori_n56_));
  NA2        o034(.A(i_8_), .B(i_7_), .Y(ori_ori_n57_));
  OAI210     o035(.A0(ori_ori_n57_), .A1(ori_ori_n56_), .B0(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(i_12_), .Y(ori_ori_n59_));
  NAi21      o037(.An(i_2_), .B(i_7_), .Y(ori_ori_n60_));
  INV        o038(.A(i_1_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n61_), .B(i_6_), .Y(ori_ori_n62_));
  NA3        o040(.A(ori_ori_n62_), .B(ori_ori_n60_), .C(ori_ori_n31_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_1_), .B(i_10_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(i_6_), .Y(ori_ori_n65_));
  NAi31      o043(.An(ori_ori_n65_), .B(ori_ori_n63_), .C(ori_ori_n59_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n67_));
  AOI210     o045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n68_));
  NA2        o046(.A(i_1_), .B(i_6_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n25_), .Y(ori_ori_n70_));
  INV        o048(.A(i_0_), .Y(ori_ori_n71_));
  NAi21      o049(.An(i_5_), .B(i_10_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_5_), .B(i_9_), .Y(ori_ori_n73_));
  AOI210     o051(.A0(ori_ori_n73_), .A1(ori_ori_n72_), .B0(ori_ori_n71_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n74_), .B(ori_ori_n70_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n68_), .A1(ori_ori_n67_), .B0(ori_ori_n75_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n76_), .A1(ori_ori_n66_), .B0(i_0_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_12_), .B(i_5_), .Y(ori_ori_n78_));
  INV        o056(.A(i_8_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n56_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_3_), .B(i_9_), .Y(ori_ori_n81_));
  NO2        o059(.A(i_3_), .B(i_7_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n81_), .B(ori_ori_n61_), .Y(ori_ori_n83_));
  INV        o061(.A(i_6_), .Y(ori_ori_n84_));
  NO2        o062(.A(i_2_), .B(i_7_), .Y(ori_ori_n85_));
  INV        o063(.A(ori_ori_n85_), .Y(ori_ori_n86_));
  OAI210     o064(.A0(ori_ori_n83_), .A1(ori_ori_n80_), .B0(ori_ori_n86_), .Y(ori_ori_n87_));
  NAi21      o065(.An(i_6_), .B(i_10_), .Y(ori_ori_n88_));
  NA2        o066(.A(i_6_), .B(i_9_), .Y(ori_ori_n89_));
  AOI210     o067(.A0(ori_ori_n89_), .A1(ori_ori_n88_), .B0(ori_ori_n61_), .Y(ori_ori_n90_));
  NA2        o068(.A(i_2_), .B(i_6_), .Y(ori_ori_n91_));
  NO3        o069(.A(ori_ori_n91_), .B(ori_ori_n48_), .C(ori_ori_n25_), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(ori_ori_n90_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n93_), .A1(ori_ori_n87_), .B0(ori_ori_n78_), .Y(ori_ori_n94_));
  AN3        o072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n95_), .B(ori_ori_n32_), .Y(ori_ori_n96_));
  INV        o074(.A(i_7_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n45_), .B(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o076(.A(i_0_), .B(i_5_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n84_), .Y(ori_ori_n100_));
  NA2        o078(.A(i_12_), .B(i_3_), .Y(ori_ori_n101_));
  INV        o079(.A(ori_ori_n101_), .Y(ori_ori_n102_));
  NA3        o080(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n98_), .Y(ori_ori_n103_));
  NAi21      o081(.An(i_7_), .B(i_11_), .Y(ori_ori_n104_));
  NO3        o082(.A(ori_ori_n104_), .B(ori_ori_n88_), .C(ori_ori_n51_), .Y(ori_ori_n105_));
  AN2        o083(.A(i_2_), .B(i_10_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(i_7_), .Y(ori_ori_n107_));
  OR2        o085(.A(ori_ori_n78_), .B(ori_ori_n56_), .Y(ori_ori_n108_));
  NA2        o086(.A(i_12_), .B(i_7_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n61_), .B(ori_ori_n26_), .Y(ori_ori_n110_));
  NA2        o088(.A(i_11_), .B(i_12_), .Y(ori_ori_n111_));
  NAi41      o089(.An(ori_ori_n105_), .B(ori_ori_n111_), .C(ori_ori_n103_), .D(ori_ori_n96_), .Y(ori_ori_n112_));
  NOi21      o090(.An(i_1_), .B(i_5_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n113_), .B(i_11_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n97_), .B(ori_ori_n37_), .Y(ori_ori_n115_));
  NA2        o093(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n117_), .B(ori_ori_n45_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n89_), .B(ori_ori_n88_), .Y(ori_ori_n119_));
  NAi21      o097(.An(i_3_), .B(i_8_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n60_), .Y(ori_ori_n121_));
  NOi31      o099(.An(ori_ori_n121_), .B(ori_ori_n119_), .C(ori_ori_n118_), .Y(ori_ori_n122_));
  NO2        o100(.A(i_1_), .B(ori_ori_n84_), .Y(ori_ori_n123_));
  NO2        o101(.A(i_6_), .B(i_5_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(i_3_), .Y(ori_ori_n125_));
  AO210      o103(.A0(ori_ori_n125_), .A1(ori_ori_n46_), .B0(ori_ori_n123_), .Y(ori_ori_n126_));
  OAI220     o104(.A0(ori_ori_n126_), .A1(ori_ori_n104_), .B0(ori_ori_n122_), .B1(ori_ori_n114_), .Y(ori_ori_n127_));
  NO3        o105(.A(ori_ori_n127_), .B(ori_ori_n112_), .C(ori_ori_n94_), .Y(ori_ori_n128_));
  NA3        o106(.A(ori_ori_n128_), .B(ori_ori_n77_), .C(ori_ori_n54_), .Y(ori2));
  NO2        o107(.A(ori_ori_n61_), .B(ori_ori_n37_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n621_), .B(ori_ori_n130_), .Y(ori_ori_n131_));
  NA4        o109(.A(ori_ori_n131_), .B(ori_ori_n75_), .C(ori_ori_n67_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o110(.A(i_12_), .B(i_13_), .Y(ori_ori_n133_));
  NAi21      o111(.An(i_5_), .B(i_11_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_0_), .B(i_1_), .Y(ori_ori_n135_));
  NA2        o113(.A(i_2_), .B(i_3_), .Y(ori_ori_n136_));
  NA2        o114(.A(i_1_), .B(i_5_), .Y(ori_ori_n137_));
  NOi21      o115(.An(i_4_), .B(i_10_), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n138_), .B(ori_ori_n40_), .Y(ori_ori_n139_));
  NOi21      o117(.An(i_4_), .B(i_9_), .Y(ori_ori_n140_));
  NOi21      o118(.An(i_11_), .B(i_13_), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n142_));
  NAi21      o120(.An(i_12_), .B(i_11_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n71_), .B(ori_ori_n61_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n71_), .B(i_5_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_2_), .B(i_1_), .Y(ori_ori_n146_));
  NAi21      o124(.An(i_4_), .B(i_12_), .Y(ori_ori_n147_));
  INV        o125(.A(i_8_), .Y(ori_ori_n148_));
  NO3        o126(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n149_));
  NO2        o127(.A(i_3_), .B(i_8_), .Y(ori_ori_n150_));
  NO3        o128(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n99_), .B(ori_ori_n56_), .Y(ori_ori_n152_));
  NO2        o130(.A(i_13_), .B(i_9_), .Y(ori_ori_n153_));
  NAi21      o131(.An(i_12_), .B(i_3_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n43_), .B(i_5_), .Y(ori_ori_n155_));
  NA3        o133(.A(i_13_), .B(ori_ori_n148_), .C(i_10_), .Y(ori_ori_n156_));
  NA2        o134(.A(i_0_), .B(i_5_), .Y(ori_ori_n157_));
  NAi31      o135(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n71_), .B(ori_ori_n26_), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n45_), .B(ori_ori_n61_), .Y(ori_ori_n161_));
  INV        o139(.A(i_13_), .Y(ori_ori_n162_));
  NO2        o140(.A(i_12_), .B(ori_ori_n162_), .Y(ori_ori_n163_));
  NO2        o141(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n164_));
  INV        o142(.A(i_12_), .Y(ori_ori_n165_));
  NO3        o143(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n166_));
  NA2        o144(.A(i_2_), .B(i_1_), .Y(ori_ori_n167_));
  NO3        o145(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n168_));
  NAi21      o146(.An(i_4_), .B(i_3_), .Y(ori_ori_n169_));
  NO2        o147(.A(i_0_), .B(i_6_), .Y(ori_ori_n170_));
  NOi41      o148(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n171_));
  NO2        o149(.A(i_11_), .B(ori_ori_n162_), .Y(ori_ori_n172_));
  NOi21      o150(.An(i_1_), .B(i_6_), .Y(ori_ori_n173_));
  NAi21      o151(.An(i_3_), .B(i_7_), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n165_), .B(i_9_), .Y(ori_ori_n175_));
  OR4        o153(.A(ori_ori_n175_), .B(ori_ori_n174_), .C(ori_ori_n173_), .D(ori_ori_n145_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n71_), .B(i_5_), .Y(ori_ori_n177_));
  NA2        o155(.A(i_3_), .B(i_9_), .Y(ori_ori_n178_));
  NAi21      o156(.An(i_7_), .B(i_10_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n179_), .B(ori_ori_n178_), .Y(ori_ori_n180_));
  NA3        o158(.A(ori_ori_n180_), .B(ori_ori_n177_), .C(ori_ori_n62_), .Y(ori_ori_n181_));
  NA2        o159(.A(ori_ori_n181_), .B(ori_ori_n176_), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n182_), .B(ori_ori_n172_), .Y(ori_ori_n183_));
  NA2        o161(.A(i_12_), .B(i_6_), .Y(ori_ori_n184_));
  OR2        o162(.A(i_13_), .B(i_9_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n169_), .B(i_2_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n172_), .B(i_9_), .Y(ori_ori_n187_));
  NO3        o165(.A(i_11_), .B(ori_ori_n162_), .C(ori_ori_n25_), .Y(ori_ori_n188_));
  NO3        o166(.A(i_12_), .B(ori_ori_n162_), .C(ori_ori_n37_), .Y(ori_ori_n189_));
  AN2        o167(.A(i_3_), .B(i_10_), .Y(ori_ori_n190_));
  NO2        o168(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n191_));
  NO3        o169(.A(ori_ori_n43_), .B(i_13_), .C(i_9_), .Y(ori_ori_n192_));
  NO2        o170(.A(i_2_), .B(i_3_), .Y(ori_ori_n193_));
  OR2        o171(.A(i_0_), .B(i_5_), .Y(ori_ori_n194_));
  NO2        o172(.A(i_12_), .B(i_10_), .Y(ori_ori_n195_));
  NOi21      o173(.An(i_5_), .B(i_0_), .Y(ori_ori_n196_));
  NO2        o174(.A(i_1_), .B(i_7_), .Y(ori_ori_n197_));
  NOi21      o175(.An(ori_ori_n137_), .B(ori_ori_n100_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n198_), .B(ori_ori_n116_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n199_), .B(i_3_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n148_), .B(i_9_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n201_), .B(ori_ori_n152_), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n202_), .B(ori_ori_n45_), .Y(ori_ori_n203_));
  INV        o181(.A(ori_ori_n203_), .Y(ori_ori_n204_));
  AOI210     o182(.A0(ori_ori_n204_), .A1(ori_ori_n200_), .B0(ori_ori_n139_), .Y(ori_ori_n205_));
  INV        o183(.A(ori_ori_n205_), .Y(ori_ori_n206_));
  NOi32      o184(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n207_));
  INV        o185(.A(ori_ori_n207_), .Y(ori_ori_n208_));
  NOi32      o186(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n209_));
  NAi21      o187(.An(i_6_), .B(i_1_), .Y(ori_ori_n210_));
  NA3        o188(.A(ori_ori_n210_), .B(ori_ori_n209_), .C(ori_ori_n45_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(i_0_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_1_), .B(ori_ori_n97_), .Y(ori_ori_n213_));
  NAi21      o191(.An(i_3_), .B(i_4_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n214_), .B(i_9_), .Y(ori_ori_n215_));
  AN2        o193(.A(i_6_), .B(i_7_), .Y(ori_ori_n216_));
  OAI210     o194(.A0(ori_ori_n216_), .A1(ori_ori_n213_), .B0(ori_ori_n215_), .Y(ori_ori_n217_));
  NA2        o195(.A(i_2_), .B(i_7_), .Y(ori_ori_n218_));
  NO2        o196(.A(ori_ori_n214_), .B(i_10_), .Y(ori_ori_n219_));
  NA3        o197(.A(ori_ori_n219_), .B(ori_ori_n218_), .C(ori_ori_n170_), .Y(ori_ori_n220_));
  AOI210     o198(.A0(ori_ori_n220_), .A1(ori_ori_n217_), .B0(ori_ori_n145_), .Y(ori_ori_n221_));
  AOI210     o199(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n222_));
  OAI210     o200(.A0(ori_ori_n222_), .A1(ori_ori_n146_), .B0(ori_ori_n219_), .Y(ori_ori_n223_));
  AOI220     o201(.A0(ori_ori_n219_), .A1(ori_ori_n197_), .B0(ori_ori_n166_), .B1(ori_ori_n146_), .Y(ori_ori_n224_));
  AOI210     o202(.A0(ori_ori_n224_), .A1(ori_ori_n223_), .B0(i_5_), .Y(ori_ori_n225_));
  NO3        o203(.A(ori_ori_n225_), .B(ori_ori_n221_), .C(ori_ori_n212_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n226_), .B(ori_ori_n208_), .Y(ori_ori_n227_));
  AN2        o205(.A(i_12_), .B(i_5_), .Y(ori_ori_n228_));
  INV        o206(.A(ori_ori_n228_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_11_), .B(i_6_), .Y(ori_ori_n230_));
  NO2        o208(.A(i_5_), .B(i_10_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n232_));
  NO3        o210(.A(ori_ori_n84_), .B(ori_ori_n47_), .C(i_9_), .Y(ori_ori_n233_));
  NO2        o211(.A(i_11_), .B(i_12_), .Y(ori_ori_n234_));
  NAi21      o212(.An(i_13_), .B(i_0_), .Y(ori_ori_n235_));
  NO3        o213(.A(i_1_), .B(i_12_), .C(ori_ori_n84_), .Y(ori_ori_n236_));
  NO2        o214(.A(i_0_), .B(i_11_), .Y(ori_ori_n237_));
  AN2        o215(.A(i_1_), .B(i_6_), .Y(ori_ori_n238_));
  NOi21      o216(.An(i_2_), .B(i_12_), .Y(ori_ori_n239_));
  NAi21      o217(.An(i_9_), .B(i_4_), .Y(ori_ori_n240_));
  OR2        o218(.A(i_13_), .B(i_10_), .Y(ori_ori_n241_));
  NO3        o219(.A(ori_ori_n241_), .B(ori_ori_n111_), .C(ori_ori_n240_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n142_), .B(ori_ori_n115_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n97_), .B(ori_ori_n25_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n189_), .B(ori_ori_n244_), .Y(ori_ori_n245_));
  NO2        o223(.A(ori_ori_n245_), .B(ori_ori_n198_), .Y(ori_ori_n246_));
  INV        o224(.A(ori_ori_n246_), .Y(ori_ori_n247_));
  NO2        o225(.A(ori_ori_n247_), .B(ori_ori_n26_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n148_), .B(i_10_), .Y(ori_ori_n249_));
  NA3        o227(.A(ori_ori_n177_), .B(ori_ori_n62_), .C(i_2_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n250_), .B(ori_ori_n249_), .Y(ori_ori_n251_));
  INV        o229(.A(ori_ori_n251_), .Y(ori_ori_n252_));
  NO2        o230(.A(ori_ori_n252_), .B(ori_ori_n187_), .Y(ori_ori_n253_));
  NO3        o231(.A(ori_ori_n253_), .B(ori_ori_n248_), .C(ori_ori_n227_), .Y(ori_ori_n254_));
  NO2        o232(.A(ori_ori_n71_), .B(i_13_), .Y(ori_ori_n255_));
  NO2        o233(.A(i_10_), .B(i_9_), .Y(ori_ori_n256_));
  NAi21      o234(.An(i_12_), .B(i_8_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n257_), .B(i_3_), .Y(ori_ori_n258_));
  NA2        o236(.A(i_8_), .B(i_9_), .Y(ori_ori_n259_));
  NA2        o237(.A(ori_ori_n189_), .B(ori_ori_n152_), .Y(ori_ori_n260_));
  NO2        o238(.A(ori_ori_n260_), .B(ori_ori_n259_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n172_), .B(ori_ori_n191_), .Y(ori_ori_n262_));
  NO3        o240(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n263_));
  INV        o241(.A(ori_ori_n263_), .Y(ori_ori_n264_));
  NA3        o242(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n265_));
  NA4        o243(.A(ori_ori_n134_), .B(ori_ori_n110_), .C(ori_ori_n78_), .D(ori_ori_n23_), .Y(ori_ori_n266_));
  OAI220     o244(.A0(ori_ori_n266_), .A1(ori_ori_n265_), .B0(ori_ori_n264_), .B1(ori_ori_n262_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n267_), .B(ori_ori_n261_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n95_), .B(i_13_), .Y(ori_ori_n269_));
  NO3        o247(.A(i_4_), .B(ori_ori_n47_), .C(i_8_), .Y(ori_ori_n270_));
  NO2        o248(.A(i_6_), .B(i_7_), .Y(ori_ori_n271_));
  NO2        o249(.A(i_11_), .B(i_1_), .Y(ori_ori_n272_));
  NOi21      o250(.An(i_2_), .B(i_7_), .Y(ori_ori_n273_));
  NO2        o251(.A(i_6_), .B(i_10_), .Y(ori_ori_n274_));
  NA3        o252(.A(ori_ori_n171_), .B(ori_ori_n141_), .C(ori_ori_n124_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n45_), .B(ori_ori_n43_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n263_), .B(ori_ori_n231_), .Y(ori_ori_n277_));
  NAi21      o255(.An(ori_ori_n156_), .B(ori_ori_n234_), .Y(ori_ori_n278_));
  NA2        o256(.A(ori_ori_n197_), .B(ori_ori_n157_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n279_), .B(ori_ori_n278_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n192_), .B(ori_ori_n166_), .Y(ori_ori_n282_));
  OAI220     o260(.A0(ori_ori_n282_), .A1(ori_ori_n250_), .B0(ori_ori_n281_), .B1(ori_ori_n269_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n283_), .B(ori_ori_n280_), .Y(ori_ori_n284_));
  NA3        o262(.A(ori_ori_n284_), .B(ori_ori_n275_), .C(ori_ori_n268_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n228_), .B(ori_ori_n162_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n216_), .B(ori_ori_n209_), .Y(ori_ori_n287_));
  OR2        o265(.A(ori_ori_n286_), .B(ori_ori_n287_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n289_));
  AOI210     o267(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n242_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n290_), .B(ori_ori_n288_), .Y(ori_ori_n291_));
  INV        o269(.A(ori_ori_n291_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n177_), .B(ori_ori_n62_), .Y(ori_ori_n293_));
  OAI210     o271(.A0(i_8_), .A1(ori_ori_n293_), .B0(ori_ori_n126_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n294_), .B(ori_ori_n243_), .Y(ori_ori_n295_));
  NA2        o273(.A(ori_ori_n295_), .B(ori_ori_n292_), .Y(ori_ori_n296_));
  NO2        o274(.A(i_12_), .B(ori_ori_n148_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n43_), .B(i_10_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(i_6_), .Y(ori_ori_n299_));
  NO2        o277(.A(i_0_), .B(i_5_), .Y(ori_ori_n300_));
  NA3        o278(.A(ori_ori_n157_), .B(ori_ori_n69_), .C(ori_ori_n43_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n189_), .B(ori_ori_n82_), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n301_), .B(ori_ori_n302_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n161_), .B(ori_ori_n160_), .Y(ori_ori_n304_));
  NA2        o282(.A(ori_ori_n256_), .B(ori_ori_n159_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n304_), .B(ori_ori_n305_), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n210_), .A1(ori_ori_n45_), .B0(ori_ori_n213_), .Y(ori_ori_n307_));
  NA2        o285(.A(i_0_), .B(ori_ori_n47_), .Y(ori_ori_n308_));
  NA3        o286(.A(ori_ori_n297_), .B(ori_ori_n188_), .C(ori_ori_n308_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n307_), .B(ori_ori_n309_), .Y(ori_ori_n310_));
  NO3        o288(.A(ori_ori_n310_), .B(ori_ori_n306_), .C(ori_ori_n303_), .Y(ori_ori_n311_));
  NOi21      o289(.An(i_10_), .B(i_6_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n84_), .B(ori_ori_n25_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n109_), .B(ori_ori_n23_), .Y(ori_ori_n314_));
  INV        o292(.A(ori_ori_n193_), .Y(ori_ori_n315_));
  NO2        o293(.A(i_12_), .B(ori_ori_n84_), .Y(ori_ori_n316_));
  NA3        o294(.A(ori_ori_n316_), .B(ori_ori_n188_), .C(ori_ori_n308_), .Y(ori_ori_n317_));
  NA3        o295(.A(ori_ori_n230_), .B(ori_ori_n189_), .C(ori_ori_n157_), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n318_), .A1(ori_ori_n317_), .B0(ori_ori_n315_), .Y(ori_ori_n319_));
  OR2        o297(.A(i_2_), .B(i_5_), .Y(ori_ori_n320_));
  OR2        o298(.A(ori_ori_n320_), .B(ori_ori_n238_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n218_), .B(ori_ori_n170_), .Y(ori_ori_n322_));
  AOI210     o300(.A0(ori_ori_n322_), .A1(ori_ori_n321_), .B0(ori_ori_n278_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n323_), .B(ori_ori_n319_), .Y(ori_ori_n324_));
  NA2        o302(.A(ori_ori_n324_), .B(ori_ori_n311_), .Y(ori_ori_n325_));
  NO3        o303(.A(ori_ori_n325_), .B(ori_ori_n296_), .C(ori_ori_n285_), .Y(ori_ori_n326_));
  NA4        o304(.A(ori_ori_n326_), .B(ori_ori_n254_), .C(ori_ori_n206_), .D(ori_ori_n183_), .Y(ori7));
  NO2        o305(.A(ori_ori_n91_), .B(ori_ori_n52_), .Y(ori_ori_n328_));
  NA2        o306(.A(ori_ori_n274_), .B(ori_ori_n82_), .Y(ori_ori_n329_));
  NA2        o307(.A(i_11_), .B(ori_ori_n148_), .Y(ori_ori_n330_));
  INV        o308(.A(ori_ori_n133_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n331_), .B(ori_ori_n329_), .Y(ori_ori_n332_));
  NA3        o310(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n333_));
  NO2        o311(.A(ori_ori_n165_), .B(i_4_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n334_), .B(i_8_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n101_), .B(ori_ori_n333_), .Y(ori_ori_n336_));
  NA2        o314(.A(i_2_), .B(ori_ori_n84_), .Y(ori_ori_n337_));
  OAI210     o315(.A0(ori_ori_n85_), .A1(ori_ori_n150_), .B0(ori_ori_n151_), .Y(ori_ori_n338_));
  NO2        o316(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n339_));
  NA2        o317(.A(i_4_), .B(i_8_), .Y(ori_ori_n340_));
  AOI210     o318(.A0(ori_ori_n340_), .A1(ori_ori_n190_), .B0(ori_ori_n339_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n337_), .Y(ori_ori_n342_));
  NO4        o320(.A(ori_ori_n342_), .B(ori_ori_n336_), .C(ori_ori_n332_), .D(ori_ori_n328_), .Y(ori_ori_n343_));
  AOI210     o321(.A0(ori_ori_n120_), .A1(ori_ori_n60_), .B0(i_10_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n344_), .A1(ori_ori_n165_), .B0(ori_ori_n138_), .Y(ori_ori_n345_));
  OR2        o323(.A(i_6_), .B(i_10_), .Y(ori_ori_n346_));
  OR3        o324(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n347_));
  INV        o325(.A(ori_ori_n149_), .Y(ori_ori_n348_));
  OR2        o326(.A(ori_ori_n345_), .B(ori_ori_n185_), .Y(ori_ori_n349_));
  AOI210     o327(.A0(ori_ori_n349_), .A1(ori_ori_n343_), .B0(ori_ori_n61_), .Y(ori_ori_n350_));
  NOi21      o328(.An(i_11_), .B(i_7_), .Y(ori_ori_n351_));
  AO210      o329(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n351_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n353_), .B(ori_ori_n153_), .Y(ori_ori_n354_));
  NA3        o332(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n354_), .B(ori_ori_n61_), .Y(ori_ori_n356_));
  NO3        o334(.A(ori_ori_n179_), .B(ori_ori_n154_), .C(ori_ori_n330_), .Y(ori_ori_n357_));
  OAI210     o335(.A0(ori_ori_n357_), .A1(ori_ori_n163_), .B0(ori_ori_n61_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n239_), .B(ori_ori_n31_), .Y(ori_ori_n359_));
  OR2        o337(.A(ori_ori_n154_), .B(ori_ori_n104_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n360_), .B(ori_ori_n359_), .Y(ori_ori_n361_));
  NO2        o339(.A(i_1_), .B(i_4_), .Y(ori_ori_n362_));
  NA2        o340(.A(ori_ori_n362_), .B(ori_ori_n361_), .Y(ori_ori_n363_));
  NO2        o341(.A(i_1_), .B(i_12_), .Y(ori_ori_n364_));
  NA3        o342(.A(ori_ori_n364_), .B(ori_ori_n106_), .C(ori_ori_n24_), .Y(ori_ori_n365_));
  BUFFER     o343(.A(ori_ori_n365_), .Y(ori_ori_n366_));
  NA3        o344(.A(ori_ori_n366_), .B(ori_ori_n363_), .C(ori_ori_n358_), .Y(ori_ori_n367_));
  OAI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n356_), .B0(i_6_), .Y(ori_ori_n368_));
  NO2        o346(.A(ori_ori_n355_), .B(ori_ori_n104_), .Y(ori_ori_n369_));
  NA2        o347(.A(ori_ori_n369_), .B(ori_ori_n316_), .Y(ori_ori_n370_));
  NO2        o348(.A(i_6_), .B(i_11_), .Y(ori_ori_n371_));
  INV        o349(.A(ori_ori_n370_), .Y(ori_ori_n372_));
  NO3        o350(.A(ori_ori_n346_), .B(i_8_), .C(ori_ori_n23_), .Y(ori_ori_n373_));
  AOI210     o351(.A0(i_1_), .A1(ori_ori_n180_), .B0(ori_ori_n373_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n374_), .B(ori_ori_n43_), .Y(ori_ori_n375_));
  INV        o353(.A(i_2_), .Y(ori_ori_n376_));
  NA2        o354(.A(ori_ori_n130_), .B(i_9_), .Y(ori_ori_n377_));
  NA3        o355(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n45_), .B(i_1_), .Y(ori_ori_n379_));
  NA3        o357(.A(ori_ori_n379_), .B(ori_ori_n184_), .C(ori_ori_n43_), .Y(ori_ori_n380_));
  OAI220     o358(.A0(ori_ori_n380_), .A1(ori_ori_n378_), .B0(ori_ori_n377_), .B1(ori_ori_n376_), .Y(ori_ori_n381_));
  AOI210     o359(.A0(ori_ori_n272_), .A1(ori_ori_n244_), .B0(ori_ori_n168_), .Y(ori_ori_n382_));
  NO2        o360(.A(ori_ori_n382_), .B(ori_ori_n337_), .Y(ori_ori_n383_));
  OR2        o361(.A(ori_ori_n383_), .B(ori_ori_n381_), .Y(ori_ori_n384_));
  NO3        o362(.A(ori_ori_n384_), .B(ori_ori_n375_), .C(ori_ori_n372_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n165_), .B(ori_ori_n97_), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n386_), .B(ori_ori_n351_), .Y(ori_ori_n387_));
  NA2        o365(.A(ori_ori_n387_), .B(i_1_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n388_), .B(ori_ori_n347_), .Y(ori_ori_n389_));
  NO2        o367(.A(ori_ori_n240_), .B(ori_ori_n84_), .Y(ori_ori_n390_));
  NA2        o368(.A(ori_ori_n389_), .B(ori_ori_n45_), .Y(ori_ori_n391_));
  NA2        o369(.A(i_3_), .B(ori_ori_n148_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n392_), .B(ori_ori_n109_), .Y(ori_ori_n393_));
  AN2        o371(.A(ori_ori_n393_), .B(ori_ori_n299_), .Y(ori_ori_n394_));
  NO2        o372(.A(i_8_), .B(ori_ori_n43_), .Y(ori_ori_n395_));
  NA2        o373(.A(i_1_), .B(i_3_), .Y(ori_ori_n396_));
  NO2        o374(.A(ori_ori_n259_), .B(ori_ori_n91_), .Y(ori_ori_n397_));
  AOI210     o375(.A0(ori_ori_n395_), .A1(ori_ori_n312_), .B0(ori_ori_n397_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n396_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n399_), .B(ori_ori_n394_), .Y(ori_ori_n400_));
  NA4        o378(.A(ori_ori_n400_), .B(ori_ori_n391_), .C(ori_ori_n385_), .D(ori_ori_n368_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n216_), .B(ori_ori_n215_), .Y(ori_ori_n402_));
  NO3        o380(.A(ori_ori_n273_), .B(ori_ori_n340_), .C(ori_ori_n84_), .Y(ori_ori_n403_));
  NA2        o381(.A(ori_ori_n403_), .B(ori_ori_n25_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n404_), .B(ori_ori_n402_), .Y(ori_ori_n405_));
  NA2        o383(.A(ori_ori_n405_), .B(i_1_), .Y(ori_ori_n406_));
  INV        o384(.A(i_1_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n214_), .B(i_2_), .Y(ori_ori_n408_));
  NO2        o386(.A(ori_ori_n406_), .B(i_13_), .Y(ori_ori_n409_));
  OR2        o387(.A(i_11_), .B(i_7_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n411_));
  INV        o389(.A(ori_ori_n411_), .Y(ori_ori_n412_));
  NO2        o390(.A(ori_ori_n273_), .B(ori_ori_n24_), .Y(ori_ori_n413_));
  AOI220     o391(.A0(ori_ori_n413_), .A1(ori_ori_n390_), .B0(ori_ori_n171_), .B1(ori_ori_n123_), .Y(ori_ori_n414_));
  OAI220     o392(.A0(ori_ori_n414_), .A1(ori_ori_n41_), .B0(ori_ori_n412_), .B1(ori_ori_n91_), .Y(ori_ori_n415_));
  INV        o393(.A(ori_ori_n415_), .Y(ori_ori_n416_));
  AOI210     o394(.A0(ori_ori_n257_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n417_));
  NOi31      o395(.An(ori_ori_n417_), .B(ori_ori_n329_), .C(ori_ori_n43_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n119_), .B(i_13_), .Y(ori_ori_n419_));
  NO2        o397(.A(ori_ori_n378_), .B(ori_ori_n109_), .Y(ori_ori_n420_));
  INV        o398(.A(ori_ori_n420_), .Y(ori_ori_n421_));
  OAI220     o399(.A0(ori_ori_n421_), .A1(ori_ori_n69_), .B0(ori_ori_n419_), .B1(ori_ori_n407_), .Y(ori_ori_n422_));
  NO3        o400(.A(ori_ori_n69_), .B(ori_ori_n32_), .C(ori_ori_n97_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n26_), .B(ori_ori_n148_), .Y(ori_ori_n424_));
  NA2        o402(.A(ori_ori_n424_), .B(i_7_), .Y(ori_ori_n425_));
  NO3        o403(.A(ori_ori_n273_), .B(ori_ori_n165_), .C(ori_ori_n84_), .Y(ori_ori_n426_));
  AOI210     o404(.A0(ori_ori_n426_), .A1(ori_ori_n425_), .B0(ori_ori_n423_), .Y(ori_ori_n427_));
  AOI210     o405(.A0(ori_ori_n230_), .A1(ori_ori_n379_), .B0(ori_ori_n90_), .Y(ori_ori_n428_));
  OAI220     o406(.A0(ori_ori_n428_), .A1(ori_ori_n335_), .B0(ori_ori_n427_), .B1(ori_ori_n348_), .Y(ori_ori_n429_));
  NO3        o407(.A(ori_ori_n429_), .B(ori_ori_n422_), .C(ori_ori_n418_), .Y(ori_ori_n430_));
  OR2        o408(.A(i_11_), .B(i_6_), .Y(ori_ori_n431_));
  NA3        o409(.A(ori_ori_n239_), .B(ori_ori_n339_), .C(i_6_), .Y(ori_ori_n432_));
  NA2        o410(.A(ori_ori_n371_), .B(i_13_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n98_), .B(ori_ori_n424_), .Y(ori_ori_n434_));
  NAi21      o412(.An(i_11_), .B(i_12_), .Y(ori_ori_n435_));
  NOi41      o413(.An(ori_ori_n107_), .B(ori_ori_n435_), .C(i_13_), .D(ori_ori_n84_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n316_), .B(ori_ori_n340_), .Y(ori_ori_n437_));
  AOI220     o415(.A0(ori_ori_n437_), .A1(ori_ori_n192_), .B0(ori_ori_n436_), .B1(ori_ori_n434_), .Y(ori_ori_n438_));
  NA3        o416(.A(ori_ori_n438_), .B(ori_ori_n433_), .C(ori_ori_n432_), .Y(ori_ori_n439_));
  NA2        o417(.A(ori_ori_n439_), .B(ori_ori_n61_), .Y(ori_ori_n440_));
  NO2        o418(.A(i_2_), .B(i_12_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n213_), .B(ori_ori_n441_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n215_), .B(ori_ori_n213_), .Y(ori_ori_n443_));
  NA2        o421(.A(ori_ori_n443_), .B(ori_ori_n442_), .Y(ori_ori_n444_));
  NA3        o422(.A(ori_ori_n444_), .B(ori_ori_n44_), .C(ori_ori_n162_), .Y(ori_ori_n445_));
  NA4        o423(.A(ori_ori_n445_), .B(ori_ori_n440_), .C(ori_ori_n430_), .D(ori_ori_n416_), .Y(ori_ori_n446_));
  OR4        o424(.A(ori_ori_n446_), .B(ori_ori_n409_), .C(ori_ori_n401_), .D(ori_ori_n350_), .Y(ori5));
  NA2        o425(.A(ori_ori_n387_), .B(ori_ori_n186_), .Y(ori_ori_n448_));
  AN2        o426(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n449_));
  NA3        o427(.A(ori_ori_n449_), .B(ori_ori_n441_), .C(ori_ori_n104_), .Y(ori_ori_n450_));
  NO2        o428(.A(ori_ori_n335_), .B(i_11_), .Y(ori_ori_n451_));
  NA2        o429(.A(ori_ori_n85_), .B(ori_ori_n451_), .Y(ori_ori_n452_));
  NA3        o430(.A(ori_ori_n452_), .B(ori_ori_n450_), .C(ori_ori_n448_), .Y(ori_ori_n453_));
  NO3        o431(.A(i_11_), .B(ori_ori_n165_), .C(i_13_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n116_), .B(ori_ori_n23_), .Y(ori_ori_n455_));
  INV        o433(.A(ori_ori_n256_), .Y(ori_ori_n456_));
  AOI220     o434(.A0(ori_ori_n193_), .A1(ori_ori_n314_), .B0(i_12_), .B1(ori_ori_n455_), .Y(ori_ori_n457_));
  INV        o435(.A(ori_ori_n457_), .Y(ori_ori_n458_));
  NO2        o436(.A(ori_ori_n458_), .B(ori_ori_n453_), .Y(ori_ori_n459_));
  INV        o437(.A(ori_ori_n141_), .Y(ori_ori_n460_));
  INV        o438(.A(ori_ori_n171_), .Y(ori_ori_n461_));
  OAI210     o439(.A0(ori_ori_n408_), .A1(ori_ori_n258_), .B0(ori_ori_n107_), .Y(ori_ori_n462_));
  AOI210     o440(.A0(ori_ori_n462_), .A1(ori_ori_n461_), .B0(ori_ori_n460_), .Y(ori_ori_n463_));
  NO2        o441(.A(ori_ori_n259_), .B(ori_ori_n26_), .Y(ori_ori_n464_));
  NO2        o442(.A(ori_ori_n464_), .B(ori_ori_n244_), .Y(ori_ori_n465_));
  NA2        o443(.A(ori_ori_n465_), .B(i_2_), .Y(ori_ori_n466_));
  INV        o444(.A(ori_ori_n466_), .Y(ori_ori_n467_));
  AOI210     o445(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n241_), .Y(ori_ori_n468_));
  AOI210     o446(.A0(ori_ori_n468_), .A1(ori_ori_n467_), .B0(ori_ori_n463_), .Y(ori_ori_n469_));
  NO2        o447(.A(ori_ori_n147_), .B(ori_ori_n117_), .Y(ori_ori_n470_));
  OAI210     o448(.A0(ori_ori_n470_), .A1(ori_ori_n455_), .B0(i_2_), .Y(ori_ori_n471_));
  INV        o449(.A(ori_ori_n142_), .Y(ori_ori_n472_));
  NO3        o450(.A(ori_ori_n352_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n473_));
  AOI210     o451(.A0(ori_ori_n472_), .A1(ori_ori_n85_), .B0(ori_ori_n473_), .Y(ori_ori_n474_));
  AOI210     o452(.A0(ori_ori_n474_), .A1(ori_ori_n471_), .B0(ori_ori_n148_), .Y(ori_ori_n475_));
  OA210      o453(.A0(ori_ori_n353_), .A1(ori_ori_n118_), .B0(i_13_), .Y(ori_ori_n476_));
  NA2        o454(.A(ori_ori_n149_), .B(ori_ori_n150_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n477_), .B(ori_ori_n218_), .Y(ori_ori_n478_));
  AOI210     o456(.A0(ori_ori_n154_), .A1(ori_ori_n136_), .B0(ori_ori_n289_), .Y(ori_ori_n479_));
  NA2        o457(.A(ori_ori_n479_), .B(ori_ori_n244_), .Y(ori_ori_n480_));
  NA3        o458(.A(i_2_), .B(ori_ori_n190_), .C(ori_ori_n116_), .Y(ori_ori_n481_));
  NA2        o459(.A(ori_ori_n481_), .B(ori_ori_n480_), .Y(ori_ori_n482_));
  NO4        o460(.A(ori_ori_n482_), .B(ori_ori_n478_), .C(ori_ori_n476_), .D(ori_ori_n475_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n484_));
  NO2        o462(.A(ori_ori_n484_), .B(ori_ori_n118_), .Y(ori_ori_n485_));
  NO2        o463(.A(ori_ori_n485_), .B(ori_ori_n330_), .Y(ori_ori_n486_));
  NA2        o464(.A(ori_ori_n486_), .B(ori_ori_n36_), .Y(ori_ori_n487_));
  NA4        o465(.A(ori_ori_n487_), .B(ori_ori_n483_), .C(ori_ori_n469_), .D(ori_ori_n459_), .Y(ori6));
  NO2        o466(.A(ori_ori_n158_), .B(ori_ori_n276_), .Y(ori_ori_n489_));
  INV        o467(.A(ori_ori_n196_), .Y(ori_ori_n490_));
  OR2        o468(.A(ori_ori_n490_), .B(i_12_), .Y(ori_ori_n491_));
  INV        o469(.A(ori_ori_n195_), .Y(ori_ori_n492_));
  NA2        o470(.A(ori_ori_n73_), .B(ori_ori_n123_), .Y(ori_ori_n493_));
  INV        o471(.A(ori_ori_n116_), .Y(ori_ori_n494_));
  NA2        o472(.A(ori_ori_n494_), .B(ori_ori_n45_), .Y(ori_ori_n495_));
  AOI210     o473(.A0(ori_ori_n495_), .A1(ori_ori_n493_), .B0(ori_ori_n492_), .Y(ori_ori_n496_));
  NO2        o474(.A(ori_ori_n287_), .B(ori_ori_n145_), .Y(ori_ori_n497_));
  NO2        o475(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n498_));
  NAi32      o476(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n431_), .B(ori_ori_n499_), .Y(ori_ori_n500_));
  OR3        o478(.A(ori_ori_n500_), .B(ori_ori_n497_), .C(ori_ori_n496_), .Y(ori_ori_n501_));
  NO2        o479(.A(ori_ori_n410_), .B(i_2_), .Y(ori_ori_n502_));
  NA2        o480(.A(ori_ori_n47_), .B(ori_ori_n37_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n503_), .B(ori_ori_n238_), .Y(ori_ori_n504_));
  NA2        o482(.A(ori_ori_n504_), .B(ori_ori_n502_), .Y(ori_ori_n505_));
  BUFFER     o483(.A(ori_ori_n353_), .Y(ori_ori_n506_));
  NA2        o484(.A(ori_ori_n506_), .B(ori_ori_n135_), .Y(ori_ori_n507_));
  AO210      o485(.A0(ori_ori_n277_), .A1(ori_ori_n456_), .B0(ori_ori_n36_), .Y(ori_ori_n508_));
  NA3        o486(.A(ori_ori_n508_), .B(ori_ori_n507_), .C(ori_ori_n505_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n489_), .B(ori_ori_n425_), .Y(ori_ori_n510_));
  NA3        o488(.A(ori_ori_n218_), .B(ori_ori_n166_), .C(ori_ori_n135_), .Y(ori_ori_n511_));
  NA2        o489(.A(ori_ori_n233_), .B(ori_ori_n68_), .Y(ori_ori_n512_));
  NA4        o490(.A(ori_ori_n512_), .B(ori_ori_n511_), .C(ori_ori_n510_), .D(ori_ori_n338_), .Y(ori_ori_n513_));
  NA2        o491(.A(ori_ori_n258_), .B(ori_ori_n256_), .Y(ori_ori_n514_));
  NO2        o492(.A(ori_ori_n346_), .B(ori_ori_n98_), .Y(ori_ori_n515_));
  OAI210     o493(.A0(ori_ori_n515_), .A1(ori_ori_n108_), .B0(ori_ori_n237_), .Y(ori_ori_n516_));
  INV        o494(.A(ori_ori_n321_), .Y(ori_ori_n517_));
  NA3        o495(.A(ori_ori_n517_), .B(ori_ori_n195_), .C(i_7_), .Y(ori_ori_n518_));
  NA3        o496(.A(ori_ori_n518_), .B(ori_ori_n516_), .C(ori_ori_n514_), .Y(ori_ori_n519_));
  NO4        o497(.A(ori_ori_n519_), .B(ori_ori_n513_), .C(ori_ori_n509_), .D(ori_ori_n501_), .Y(ori_ori_n520_));
  NA3        o498(.A(ori_ori_n520_), .B(ori_ori_n491_), .C(ori_ori_n226_), .Y(ori3));
  NA2        o499(.A(i_12_), .B(i_10_), .Y(ori_ori_n522_));
  NO2        o500(.A(i_11_), .B(ori_ori_n165_), .Y(ori_ori_n523_));
  NA3        o501(.A(ori_ori_n511_), .B(ori_ori_n338_), .C(ori_ori_n217_), .Y(ori_ori_n524_));
  NA2        o502(.A(ori_ori_n524_), .B(ori_ori_n40_), .Y(ori_ori_n525_));
  NOi21      o503(.An(ori_ori_n95_), .B(ori_ori_n465_), .Y(ori_ori_n526_));
  NO3        o504(.A(ori_ori_n360_), .B(ori_ori_n259_), .C(ori_ori_n123_), .Y(ori_ori_n527_));
  NA2        o505(.A(ori_ori_n239_), .B(ori_ori_n44_), .Y(ori_ori_n528_));
  AN2        o506(.A(i_11_), .B(ori_ori_n53_), .Y(ori_ori_n529_));
  NO3        o507(.A(ori_ori_n529_), .B(ori_ori_n527_), .C(ori_ori_n526_), .Y(ori_ori_n530_));
  AOI210     o508(.A0(ori_ori_n530_), .A1(ori_ori_n525_), .B0(ori_ori_n47_), .Y(ori_ori_n531_));
  NO4        o509(.A(ori_ori_n222_), .B(ori_ori_n228_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n532_));
  NA2        o510(.A(ori_ori_n145_), .B(ori_ori_n312_), .Y(ori_ori_n533_));
  NOi21      o511(.An(ori_ori_n533_), .B(ori_ori_n532_), .Y(ori_ori_n534_));
  NO2        o512(.A(ori_ori_n534_), .B(ori_ori_n61_), .Y(ori_ori_n535_));
  NOi21      o513(.An(i_5_), .B(i_9_), .Y(ori_ori_n536_));
  NA2        o514(.A(ori_ori_n536_), .B(ori_ori_n255_), .Y(ori_ori_n537_));
  BUFFER     o515(.A(ori_ori_n184_), .Y(ori_ori_n538_));
  AOI210     o516(.A0(ori_ori_n538_), .A1(ori_ori_n272_), .B0(ori_ori_n403_), .Y(ori_ori_n539_));
  NO2        o517(.A(ori_ori_n539_), .B(ori_ori_n537_), .Y(ori_ori_n540_));
  NO3        o518(.A(ori_ori_n540_), .B(ori_ori_n535_), .C(ori_ori_n531_), .Y(ori_ori_n541_));
  NA2        o519(.A(ori_ori_n313_), .B(i_0_), .Y(ori_ori_n542_));
  NO3        o520(.A(ori_ori_n542_), .B(ori_ori_n229_), .C(ori_ori_n85_), .Y(ori_ori_n543_));
  NO4        o521(.A(ori_ori_n320_), .B(i_12_), .C(ori_ori_n241_), .D(ori_ori_n238_), .Y(ori_ori_n544_));
  AOI210     o522(.A0(ori_ori_n544_), .A1(i_11_), .B0(ori_ori_n543_), .Y(ori_ori_n545_));
  NA2        o523(.A(ori_ori_n454_), .B(ori_ori_n196_), .Y(ori_ori_n546_));
  NO2        o524(.A(ori_ori_n85_), .B(ori_ori_n56_), .Y(ori_ori_n547_));
  NO2        o525(.A(ori_ori_n547_), .B(ori_ori_n546_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n175_), .B(ori_ori_n137_), .Y(ori_ori_n549_));
  INV        o527(.A(ori_ori_n298_), .Y(ori_ori_n550_));
  NO4        o528(.A(ori_ori_n109_), .B(ori_ori_n56_), .C(ori_ori_n392_), .D(i_5_), .Y(ori_ori_n551_));
  AO220      o529(.A0(ori_ori_n551_), .A1(ori_ori_n550_), .B0(ori_ori_n549_), .B1(i_6_), .Y(ori_ori_n552_));
  NO2        o530(.A(ori_ori_n552_), .B(ori_ori_n548_), .Y(ori_ori_n553_));
  NA2        o531(.A(ori_ori_n553_), .B(ori_ori_n545_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n99_), .B(ori_ori_n37_), .Y(ori_ori_n555_));
  NA2        o533(.A(i_11_), .B(i_9_), .Y(ori_ori_n556_));
  NO3        o534(.A(i_12_), .B(ori_ori_n556_), .C(ori_ori_n337_), .Y(ori_ori_n557_));
  AN2        o535(.A(ori_ori_n557_), .B(ori_ori_n555_), .Y(ori_ori_n558_));
  NA2        o536(.A(ori_ori_n232_), .B(ori_ori_n144_), .Y(ori_ori_n559_));
  INV        o537(.A(ori_ori_n559_), .Y(ori_ori_n560_));
  NO2        o538(.A(ori_ori_n556_), .B(ori_ori_n71_), .Y(ori_ori_n561_));
  INV        o539(.A(ori_ori_n236_), .Y(ori_ori_n562_));
  NO2        o540(.A(ori_ori_n562_), .B(ori_ori_n537_), .Y(ori_ori_n563_));
  NO3        o541(.A(ori_ori_n563_), .B(ori_ori_n560_), .C(ori_ori_n558_), .Y(ori_ori_n564_));
  INV        o542(.A(ori_ori_n194_), .Y(ori_ori_n565_));
  INV        o543(.A(ori_ori_n564_), .Y(ori_ori_n566_));
  INV        o544(.A(ori_ori_n522_), .Y(ori_ori_n567_));
  OA210      o545(.A0(ori_ori_n271_), .A1(ori_ori_n161_), .B0(ori_ori_n270_), .Y(ori_ori_n568_));
  NA2        o546(.A(ori_ori_n567_), .B(ori_ori_n561_), .Y(ori_ori_n569_));
  NA2        o547(.A(ori_ori_n413_), .B(ori_ori_n300_), .Y(ori_ori_n570_));
  NAi21      o548(.An(i_9_), .B(i_5_), .Y(ori_ori_n571_));
  NO2        o549(.A(ori_ori_n571_), .B(ori_ori_n235_), .Y(ori_ori_n572_));
  NA2        o550(.A(ori_ori_n572_), .B(ori_ori_n353_), .Y(ori_ori_n573_));
  OAI220     o551(.A0(ori_ori_n573_), .A1(ori_ori_n84_), .B0(ori_ori_n570_), .B1(ori_ori_n142_), .Y(ori_ori_n574_));
  NO2        o552(.A(ori_ori_n574_), .B(ori_ori_n291_), .Y(ori_ori_n575_));
  NA2        o553(.A(ori_ori_n575_), .B(ori_ori_n569_), .Y(ori_ori_n576_));
  NO3        o554(.A(ori_ori_n576_), .B(ori_ori_n566_), .C(ori_ori_n554_), .Y(ori_ori_n577_));
  NO2        o555(.A(i_0_), .B(ori_ori_n435_), .Y(ori_ori_n578_));
  NA2        o556(.A(ori_ori_n170_), .B(ori_ori_n164_), .Y(ori_ori_n579_));
  AOI210     o557(.A0(ori_ori_n579_), .A1(ori_ori_n542_), .B0(ori_ori_n137_), .Y(ori_ori_n580_));
  NO3        o558(.A(ori_ori_n155_), .B(ori_ori_n228_), .C(i_0_), .Y(ori_ori_n581_));
  OAI210     o559(.A0(ori_ori_n581_), .A1(ori_ori_n74_), .B0(i_13_), .Y(ori_ori_n582_));
  INV        o560(.A(ori_ori_n582_), .Y(ori_ori_n583_));
  NO2        o561(.A(ori_ori_n169_), .B(ori_ori_n91_), .Y(ori_ori_n584_));
  AOI210     o562(.A0(ori_ori_n584_), .A1(ori_ori_n578_), .B0(ori_ori_n105_), .Y(ori_ori_n585_));
  OR2        o563(.A(ori_ori_n585_), .B(i_5_), .Y(ori_ori_n586_));
  AOI210     o564(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n143_), .Y(ori_ori_n587_));
  NA2        o565(.A(ori_ori_n587_), .B(ori_ori_n568_), .Y(ori_ori_n588_));
  NO3        o566(.A(ori_ori_n528_), .B(ori_ori_n52_), .C(ori_ori_n47_), .Y(ori_ori_n589_));
  NO2        o567(.A(ori_ori_n622_), .B(ori_ori_n589_), .Y(ori_ori_n590_));
  NA3        o568(.A(ori_ori_n231_), .B(ori_ori_n141_), .C(ori_ori_n140_), .Y(ori_ori_n591_));
  INV        o569(.A(ori_ori_n591_), .Y(ori_ori_n592_));
  NO3        o570(.A(ori_ori_n556_), .B(ori_ori_n157_), .C(ori_ori_n147_), .Y(ori_ori_n593_));
  NO2        o571(.A(ori_ori_n593_), .B(ori_ori_n592_), .Y(ori_ori_n594_));
  NA4        o572(.A(ori_ori_n594_), .B(ori_ori_n590_), .C(ori_ori_n588_), .D(ori_ori_n586_), .Y(ori_ori_n595_));
  NO2        o573(.A(ori_ori_n84_), .B(i_5_), .Y(ori_ori_n596_));
  NA3        o574(.A(ori_ori_n523_), .B(ori_ori_n106_), .C(ori_ori_n116_), .Y(ori_ori_n597_));
  INV        o575(.A(ori_ori_n597_), .Y(ori_ori_n598_));
  NA2        o576(.A(ori_ori_n598_), .B(ori_ori_n596_), .Y(ori_ori_n599_));
  NAi21      o577(.An(ori_ori_n168_), .B(ori_ori_n169_), .Y(ori_ori_n600_));
  NO4        o578(.A(ori_ori_n167_), .B(ori_ori_n155_), .C(i_0_), .D(i_12_), .Y(ori_ori_n601_));
  NA2        o579(.A(ori_ori_n601_), .B(ori_ori_n600_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n602_), .B(ori_ori_n599_), .Y(ori_ori_n603_));
  NO4        o581(.A(ori_ori_n603_), .B(ori_ori_n595_), .C(ori_ori_n583_), .D(ori_ori_n580_), .Y(ori_ori_n604_));
  OAI210     o582(.A0(ori_ori_n502_), .A1(ori_ori_n498_), .B0(ori_ori_n37_), .Y(ori_ori_n605_));
  NA2        o583(.A(ori_ori_n605_), .B(ori_ori_n345_), .Y(ori_ori_n606_));
  NA2        o584(.A(ori_ori_n606_), .B(ori_ori_n153_), .Y(ori_ori_n607_));
  NAi31      o585(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n608_));
  NO2        o586(.A(ori_ori_n68_), .B(ori_ori_n608_), .Y(ori_ori_n609_));
  AOI210     o587(.A0(ori_ori_n609_), .A1(ori_ori_n47_), .B0(ori_ori_n544_), .Y(ori_ori_n610_));
  AOI210     o588(.A0(ori_ori_n610_), .A1(ori_ori_n607_), .B0(ori_ori_n71_), .Y(ori_ori_n611_));
  INV        o589(.A(ori_ori_n225_), .Y(ori_ori_n612_));
  NO2        o590(.A(ori_ori_n612_), .B(ori_ori_n460_), .Y(ori_ori_n613_));
  NO3        o591(.A(ori_ori_n57_), .B(ori_ori_n56_), .C(i_4_), .Y(ori_ori_n614_));
  OAI210     o592(.A0(ori_ori_n565_), .A1(ori_ori_n191_), .B0(ori_ori_n614_), .Y(ori_ori_n615_));
  NO2        o593(.A(ori_ori_n615_), .B(ori_ori_n435_), .Y(ori_ori_n616_));
  NO3        o594(.A(ori_ori_n616_), .B(ori_ori_n613_), .C(ori_ori_n611_), .Y(ori_ori_n617_));
  NA4        o595(.A(ori_ori_n617_), .B(ori_ori_n604_), .C(ori_ori_n577_), .D(ori_ori_n541_), .Y(ori4));
  INV        o596(.A(i_6_), .Y(ori_ori_n621_));
  INV        o597(.A(ori_ori_n275_), .Y(ori_ori_n622_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NO2        m028(.A(mai_mai_n47_), .B(mai_mai_n46_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_0_), .B(i_2_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_7_), .B(i_9_), .Y(mai_mai_n53_));
  NA2        m031(.A(mai_mai_n51_), .B(mai_mai_n45_), .Y(mai_mai_n54_));
  NO2        m032(.A(i_1_), .B(i_6_), .Y(mai_mai_n55_));
  NA2        m033(.A(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  NAi21      m034(.An(i_2_), .B(i_7_), .Y(mai_mai_n57_));
  INV        m035(.A(i_1_), .Y(mai_mai_n58_));
  NA2        m036(.A(i_1_), .B(i_10_), .Y(mai_mai_n59_));
  NO2        m037(.A(mai_mai_n59_), .B(i_6_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n61_));
  AOI210     m039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_1_), .B(i_6_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(mai_mai_n25_), .Y(mai_mai_n64_));
  INV        m042(.A(i_0_), .Y(mai_mai_n65_));
  NAi21      m043(.An(i_5_), .B(i_10_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_5_), .B(i_9_), .Y(mai_mai_n67_));
  AOI210     m045(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n65_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n64_), .Y(mai_mai_n69_));
  OAI210     m047(.A0(mai_mai_n62_), .A1(mai_mai_n61_), .B0(mai_mai_n69_), .Y(mai_mai_n70_));
  OAI210     m048(.A0(mai_mai_n70_), .A1(mai_mai_n60_), .B0(i_0_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_12_), .B(i_5_), .Y(mai_mai_n72_));
  NO2        m050(.A(i_3_), .B(i_9_), .Y(mai_mai_n73_));
  NO2        m051(.A(i_3_), .B(i_7_), .Y(mai_mai_n74_));
  NO3        m052(.A(mai_mai_n74_), .B(mai_mai_n73_), .C(mai_mai_n58_), .Y(mai_mai_n75_));
  INV        m053(.A(i_6_), .Y(mai_mai_n76_));
  OR4        m054(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n77_));
  INV        m055(.A(mai_mai_n77_), .Y(mai_mai_n78_));
  NO2        m056(.A(i_2_), .B(i_7_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n78_), .B(mai_mai_n79_), .Y(mai_mai_n80_));
  NA2        m058(.A(mai_mai_n75_), .B(mai_mai_n80_), .Y(mai_mai_n81_));
  NAi21      m059(.An(i_6_), .B(i_10_), .Y(mai_mai_n82_));
  NA2        m060(.A(i_6_), .B(i_9_), .Y(mai_mai_n83_));
  AOI210     m061(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n58_), .Y(mai_mai_n84_));
  NA2        m062(.A(i_2_), .B(i_6_), .Y(mai_mai_n85_));
  INV        m063(.A(mai_mai_n84_), .Y(mai_mai_n86_));
  AOI210     m064(.A0(mai_mai_n86_), .A1(mai_mai_n81_), .B0(mai_mai_n72_), .Y(mai_mai_n87_));
  AN3        m065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n88_));
  NAi21      m066(.An(i_6_), .B(i_11_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_5_), .B(i_8_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  AOI220     m069(.A0(mai_mai_n91_), .A1(mai_mai_n57_), .B0(mai_mai_n88_), .B1(mai_mai_n32_), .Y(mai_mai_n92_));
  INV        m070(.A(i_7_), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n46_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_0_), .B(i_5_), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n95_), .B(mai_mai_n76_), .Y(mai_mai_n96_));
  NA2        m074(.A(i_12_), .B(i_3_), .Y(mai_mai_n97_));
  INV        m075(.A(mai_mai_n97_), .Y(mai_mai_n98_));
  NA3        m076(.A(mai_mai_n98_), .B(mai_mai_n96_), .C(mai_mai_n94_), .Y(mai_mai_n99_));
  NAi21      m077(.An(i_7_), .B(i_11_), .Y(mai_mai_n100_));
  AN2        m078(.A(i_2_), .B(i_10_), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n101_), .B(i_7_), .Y(mai_mai_n102_));
  OR2        m080(.A(mai_mai_n72_), .B(mai_mai_n55_), .Y(mai_mai_n103_));
  NO2        m081(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n104_));
  NO3        m082(.A(mai_mai_n104_), .B(mai_mai_n103_), .C(mai_mai_n102_), .Y(mai_mai_n105_));
  NA2        m083(.A(i_12_), .B(i_7_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n58_), .B(mai_mai_n26_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n107_), .B(i_0_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_11_), .B(i_12_), .Y(mai_mai_n109_));
  OAI210     m087(.A0(mai_mai_n108_), .A1(mai_mai_n106_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n110_), .B(mai_mai_n105_), .Y(mai_mai_n111_));
  NA3        m089(.A(mai_mai_n111_), .B(mai_mai_n99_), .C(mai_mai_n92_), .Y(mai_mai_n112_));
  NOi21      m090(.An(i_1_), .B(i_5_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n113_), .B(i_11_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n93_), .B(mai_mai_n37_), .Y(mai_mai_n115_));
  NA2        m093(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n117_), .B(mai_mai_n46_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n119_));
  NAi21      m097(.An(i_3_), .B(i_8_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n120_), .B(mai_mai_n57_), .Y(mai_mai_n121_));
  NOi31      m099(.An(mai_mai_n121_), .B(mai_mai_n119_), .C(mai_mai_n118_), .Y(mai_mai_n122_));
  NO2        m100(.A(i_1_), .B(mai_mai_n76_), .Y(mai_mai_n123_));
  NO2        m101(.A(i_6_), .B(i_5_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(i_3_), .Y(mai_mai_n125_));
  OAI220     m103(.A0(mai_mai_n125_), .A1(mai_mai_n100_), .B0(mai_mai_n122_), .B1(mai_mai_n114_), .Y(mai_mai_n126_));
  NO3        m104(.A(mai_mai_n126_), .B(mai_mai_n112_), .C(mai_mai_n87_), .Y(mai_mai_n127_));
  NA3        m105(.A(mai_mai_n127_), .B(mai_mai_n71_), .C(mai_mai_n54_), .Y(mai2));
  NO2        m106(.A(mai_mai_n58_), .B(mai_mai_n37_), .Y(mai_mai_n129_));
  NA2        m107(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n129_), .Y(mai_mai_n131_));
  NA4        m109(.A(mai_mai_n131_), .B(mai_mai_n69_), .C(mai_mai_n61_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m110(.A(i_8_), .B(i_7_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(i_6_), .Y(mai_mai_n134_));
  NO2        m112(.A(i_12_), .B(i_13_), .Y(mai_mai_n135_));
  NAi21      m113(.An(i_5_), .B(i_11_), .Y(mai_mai_n136_));
  NOi21      m114(.An(mai_mai_n135_), .B(mai_mai_n136_), .Y(mai_mai_n137_));
  NO2        m115(.A(i_0_), .B(i_1_), .Y(mai_mai_n138_));
  NA2        m116(.A(i_2_), .B(i_3_), .Y(mai_mai_n139_));
  NO2        m117(.A(mai_mai_n139_), .B(i_4_), .Y(mai_mai_n140_));
  NA3        m118(.A(mai_mai_n140_), .B(mai_mai_n138_), .C(mai_mai_n137_), .Y(mai_mai_n141_));
  AN2        m119(.A(mai_mai_n135_), .B(mai_mai_n73_), .Y(mai_mai_n142_));
  NA2        m120(.A(i_1_), .B(i_5_), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n65_), .B(mai_mai_n46_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n144_), .B(mai_mai_n36_), .Y(mai_mai_n145_));
  NO3        m123(.A(mai_mai_n145_), .B(mai_mai_n143_), .C(i_13_), .Y(mai_mai_n146_));
  OR2        m124(.A(i_0_), .B(i_1_), .Y(mai_mai_n147_));
  NO3        m125(.A(mai_mai_n147_), .B(mai_mai_n72_), .C(i_13_), .Y(mai_mai_n148_));
  NAi32      m126(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n149_));
  NAi21      m127(.An(mai_mai_n149_), .B(mai_mai_n148_), .Y(mai_mai_n150_));
  NOi21      m128(.An(i_4_), .B(i_10_), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n151_), .B(mai_mai_n40_), .Y(mai_mai_n152_));
  NO2        m130(.A(i_3_), .B(i_5_), .Y(mai_mai_n153_));
  NO3        m131(.A(mai_mai_n65_), .B(i_2_), .C(i_1_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n154_), .B(mai_mai_n153_), .Y(mai_mai_n155_));
  OAI210     m133(.A0(mai_mai_n155_), .A1(mai_mai_n152_), .B0(mai_mai_n150_), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n156_), .B(mai_mai_n146_), .Y(mai_mai_n157_));
  AOI210     m135(.A0(mai_mai_n157_), .A1(mai_mai_n141_), .B0(mai_mai_n134_), .Y(mai_mai_n158_));
  NA2        m136(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n159_));
  NOi21      m137(.An(i_4_), .B(i_9_), .Y(mai_mai_n160_));
  NOi21      m138(.An(i_11_), .B(i_13_), .Y(mai_mai_n161_));
  NA2        m139(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  OR2        m140(.A(mai_mai_n162_), .B(mai_mai_n159_), .Y(mai_mai_n163_));
  NO2        m141(.A(i_4_), .B(i_5_), .Y(mai_mai_n164_));
  NAi21      m142(.An(i_12_), .B(i_11_), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n165_), .B(i_13_), .Y(mai_mai_n166_));
  NA3        m144(.A(mai_mai_n166_), .B(mai_mai_n164_), .C(mai_mai_n73_), .Y(mai_mai_n167_));
  NA2        m145(.A(mai_mai_n167_), .B(mai_mai_n163_), .Y(mai_mai_n168_));
  NO2        m146(.A(mai_mai_n65_), .B(mai_mai_n58_), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n169_), .B(mai_mai_n46_), .Y(mai_mai_n170_));
  NAi31      m148(.An(mai_mai_n965_), .B(mai_mai_n142_), .C(i_11_), .Y(mai_mai_n171_));
  NA2        m149(.A(i_3_), .B(i_5_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(mai_mai_n162_), .A1(mai_mai_n171_), .B0(mai_mai_n170_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n65_), .B(i_5_), .Y(mai_mai_n174_));
  NO2        m152(.A(i_13_), .B(i_10_), .Y(mai_mai_n175_));
  NA3        m153(.A(mai_mai_n175_), .B(mai_mai_n174_), .C(mai_mai_n44_), .Y(mai_mai_n176_));
  NO2        m154(.A(i_2_), .B(i_1_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n177_), .B(i_3_), .Y(mai_mai_n178_));
  NAi21      m156(.An(i_4_), .B(i_12_), .Y(mai_mai_n179_));
  NO3        m157(.A(mai_mai_n179_), .B(mai_mai_n178_), .C(mai_mai_n176_), .Y(mai_mai_n180_));
  NO3        m158(.A(mai_mai_n180_), .B(mai_mai_n173_), .C(mai_mai_n168_), .Y(mai_mai_n181_));
  INV        m159(.A(i_8_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n182_), .B(i_7_), .Y(mai_mai_n183_));
  NA2        m161(.A(mai_mai_n183_), .B(i_6_), .Y(mai_mai_n184_));
  NO3        m162(.A(i_3_), .B(mai_mai_n76_), .C(mai_mai_n48_), .Y(mai_mai_n185_));
  NA2        m163(.A(mai_mai_n185_), .B(mai_mai_n104_), .Y(mai_mai_n186_));
  NO3        m164(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n187_));
  NA3        m165(.A(mai_mai_n187_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n188_));
  NO3        m166(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n189_));
  INV        m167(.A(mai_mai_n189_), .Y(mai_mai_n190_));
  AOI210     m168(.A0(mai_mai_n190_), .A1(mai_mai_n188_), .B0(mai_mai_n186_), .Y(mai_mai_n191_));
  NO2        m169(.A(i_3_), .B(i_8_), .Y(mai_mai_n192_));
  NO3        m170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n193_));
  NA3        m171(.A(mai_mai_n193_), .B(mai_mai_n192_), .C(mai_mai_n40_), .Y(mai_mai_n194_));
  NO2        m172(.A(mai_mai_n95_), .B(mai_mai_n55_), .Y(mai_mai_n195_));
  NO2        m173(.A(i_13_), .B(i_9_), .Y(mai_mai_n196_));
  NA3        m174(.A(mai_mai_n196_), .B(i_6_), .C(mai_mai_n182_), .Y(mai_mai_n197_));
  BUFFER     m175(.A(mai_mai_n197_), .Y(mai_mai_n198_));
  NO2        m176(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n199_));
  NO3        m177(.A(i_0_), .B(i_2_), .C(mai_mai_n58_), .Y(mai_mai_n200_));
  NA3        m178(.A(mai_mai_n200_), .B(mai_mai_n199_), .C(i_10_), .Y(mai_mai_n201_));
  OAI210     m179(.A0(mai_mai_n201_), .A1(mai_mai_n198_), .B0(mai_mai_n194_), .Y(mai_mai_n202_));
  AOI210     m180(.A0(mai_mai_n202_), .A1(i_7_), .B0(mai_mai_n191_), .Y(mai_mai_n203_));
  OAI220     m181(.A0(mai_mai_n203_), .A1(i_4_), .B0(mai_mai_n184_), .B1(mai_mai_n181_), .Y(mai_mai_n204_));
  NA3        m182(.A(i_13_), .B(mai_mai_n182_), .C(i_10_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n205_), .B(i_12_), .Y(mai_mai_n206_));
  NA2        m184(.A(i_0_), .B(i_5_), .Y(mai_mai_n207_));
  OAI220     m185(.A0(mai_mai_n76_), .A1(mai_mai_n178_), .B0(mai_mai_n170_), .B1(mai_mai_n125_), .Y(mai_mai_n208_));
  NAi31      m186(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n46_), .B(mai_mai_n58_), .Y(mai_mai_n211_));
  NA3        m189(.A(mai_mai_n211_), .B(i_3_), .C(mai_mai_n210_), .Y(mai_mai_n212_));
  INV        m190(.A(i_13_), .Y(mai_mai_n213_));
  NO2        m191(.A(i_12_), .B(mai_mai_n213_), .Y(mai_mai_n214_));
  NA3        m192(.A(mai_mai_n214_), .B(mai_mai_n187_), .C(mai_mai_n185_), .Y(mai_mai_n215_));
  OAI210     m193(.A0(mai_mai_n212_), .A1(mai_mai_n209_), .B0(mai_mai_n215_), .Y(mai_mai_n216_));
  AOI220     m194(.A0(mai_mai_n216_), .A1(mai_mai_n133_), .B0(mai_mai_n208_), .B1(mai_mai_n206_), .Y(mai_mai_n217_));
  NO2        m195(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n172_), .B(i_4_), .Y(mai_mai_n219_));
  NA2        m197(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  OR2        m198(.A(i_8_), .B(i_7_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n221_), .B(mai_mai_n76_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n52_), .B(i_1_), .Y(mai_mai_n223_));
  INV        m201(.A(i_12_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n44_), .B(mai_mai_n224_), .Y(mai_mai_n225_));
  NO3        m203(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n226_));
  NA2        m204(.A(i_2_), .B(i_1_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n52_), .B(mai_mai_n220_), .Y(mai_mai_n228_));
  NO3        m206(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n229_));
  NAi21      m207(.An(i_4_), .B(i_3_), .Y(mai_mai_n230_));
  INV        m208(.A(mai_mai_n67_), .Y(mai_mai_n231_));
  NO2        m209(.A(i_0_), .B(i_6_), .Y(mai_mai_n232_));
  NOi41      m210(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n233_), .B(mai_mai_n232_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n227_), .B(mai_mai_n172_), .Y(mai_mai_n235_));
  NAi21      m213(.An(mai_mai_n234_), .B(mai_mai_n235_), .Y(mai_mai_n236_));
  INV        m214(.A(mai_mai_n236_), .Y(mai_mai_n237_));
  AOI220     m215(.A0(mai_mai_n237_), .A1(mai_mai_n40_), .B0(mai_mai_n228_), .B1(mai_mai_n196_), .Y(mai_mai_n238_));
  NO2        m216(.A(i_11_), .B(mai_mai_n213_), .Y(mai_mai_n239_));
  NOi21      m217(.An(i_1_), .B(i_6_), .Y(mai_mai_n240_));
  NAi21      m218(.An(i_3_), .B(i_7_), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n224_), .B(i_9_), .Y(mai_mai_n242_));
  NO2        m220(.A(i_12_), .B(i_3_), .Y(mai_mai_n243_));
  NA3        m221(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n244_));
  INV        m222(.A(mai_mai_n134_), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n224_), .B(i_13_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n246_), .B(mai_mai_n67_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n247_), .B(mai_mai_n245_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n221_), .B(mai_mai_n37_), .Y(mai_mai_n249_));
  NA2        m227(.A(i_12_), .B(i_6_), .Y(mai_mai_n250_));
  OR2        m228(.A(i_13_), .B(i_9_), .Y(mai_mai_n251_));
  NO3        m229(.A(mai_mai_n251_), .B(mai_mai_n250_), .C(mai_mai_n48_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n230_), .B(i_2_), .Y(mai_mai_n253_));
  NA3        m231(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n44_), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n239_), .B(i_9_), .Y(mai_mai_n255_));
  OAI210     m233(.A0(mai_mai_n58_), .A1(mai_mai_n255_), .B0(mai_mai_n254_), .Y(mai_mai_n256_));
  NO3        m234(.A(i_11_), .B(mai_mai_n213_), .C(mai_mai_n25_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n241_), .B(i_8_), .Y(mai_mai_n258_));
  NO2        m236(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n259_));
  NA3        m237(.A(mai_mai_n259_), .B(mai_mai_n258_), .C(mai_mai_n257_), .Y(mai_mai_n260_));
  NO3        m238(.A(mai_mai_n26_), .B(mai_mai_n76_), .C(i_5_), .Y(mai_mai_n261_));
  NA3        m239(.A(mai_mai_n261_), .B(mai_mai_n249_), .C(mai_mai_n214_), .Y(mai_mai_n262_));
  AOI210     m240(.A0(mai_mai_n262_), .A1(mai_mai_n260_), .B0(i_1_), .Y(mai_mai_n263_));
  AOI210     m241(.A0(mai_mai_n256_), .A1(mai_mai_n249_), .B0(mai_mai_n263_), .Y(mai_mai_n264_));
  NA4        m242(.A(mai_mai_n264_), .B(mai_mai_n248_), .C(mai_mai_n238_), .D(mai_mai_n217_), .Y(mai_mai_n265_));
  NO3        m243(.A(i_12_), .B(mai_mai_n213_), .C(mai_mai_n37_), .Y(mai_mai_n266_));
  INV        m244(.A(mai_mai_n266_), .Y(mai_mai_n267_));
  NA2        m245(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n268_));
  NO3        m246(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n269_));
  AOI220     m247(.A0(mai_mai_n269_), .A1(mai_mai_n185_), .B0(mai_mai_n153_), .B1(mai_mai_n223_), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n270_), .B(mai_mai_n268_), .Y(mai_mai_n271_));
  NO3        m249(.A(i_0_), .B(i_2_), .C(mai_mai_n58_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n227_), .B(i_0_), .Y(mai_mai_n273_));
  AOI220     m251(.A0(mai_mai_n273_), .A1(mai_mai_n183_), .B0(mai_mai_n272_), .B1(mai_mai_n133_), .Y(mai_mai_n274_));
  NA2        m252(.A(mai_mai_n259_), .B(mai_mai_n26_), .Y(mai_mai_n275_));
  NO2        m253(.A(mai_mai_n275_), .B(mai_mai_n274_), .Y(mai_mai_n276_));
  NA2        m254(.A(i_0_), .B(i_1_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n277_), .B(i_2_), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n56_), .B(i_6_), .Y(mai_mai_n279_));
  NA3        m257(.A(mai_mai_n279_), .B(mai_mai_n278_), .C(mai_mai_n153_), .Y(mai_mai_n280_));
  OAI210     m258(.A0(mai_mai_n155_), .A1(mai_mai_n134_), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  NO3        m259(.A(mai_mai_n281_), .B(mai_mai_n276_), .C(mai_mai_n271_), .Y(mai_mai_n282_));
  NO2        m260(.A(i_3_), .B(i_10_), .Y(mai_mai_n283_));
  NA3        m261(.A(mai_mai_n283_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n284_));
  NO2        m262(.A(i_2_), .B(mai_mai_n93_), .Y(mai_mai_n285_));
  NA2        m263(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n286_));
  NO2        m264(.A(mai_mai_n286_), .B(i_8_), .Y(mai_mai_n287_));
  INV        m265(.A(mai_mai_n287_), .Y(mai_mai_n288_));
  AN2        m266(.A(i_3_), .B(i_10_), .Y(mai_mai_n289_));
  NA4        m267(.A(mai_mai_n289_), .B(mai_mai_n187_), .C(mai_mai_n166_), .D(mai_mai_n164_), .Y(mai_mai_n290_));
  NO2        m268(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n292_));
  OR2        m270(.A(mai_mai_n288_), .B(mai_mai_n284_), .Y(mai_mai_n293_));
  OAI220     m271(.A0(mai_mai_n293_), .A1(i_6_), .B0(mai_mai_n282_), .B1(mai_mai_n267_), .Y(mai_mai_n294_));
  NO4        m272(.A(mai_mai_n294_), .B(mai_mai_n265_), .C(mai_mai_n204_), .D(mai_mai_n158_), .Y(mai_mai_n295_));
  NO3        m273(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n296_));
  NO3        m274(.A(i_6_), .B(mai_mai_n182_), .C(i_7_), .Y(mai_mai_n297_));
  AOI210     m275(.A0(mai_mai_n967_), .A1(mai_mai_n227_), .B0(mai_mai_n159_), .Y(mai_mai_n298_));
  NO2        m276(.A(i_2_), .B(i_3_), .Y(mai_mai_n299_));
  OR2        m277(.A(i_0_), .B(i_5_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n207_), .B(mai_mai_n300_), .Y(mai_mai_n301_));
  NA4        m279(.A(mai_mai_n301_), .B(mai_mai_n222_), .C(mai_mai_n299_), .D(i_1_), .Y(mai_mai_n302_));
  NA3        m280(.A(mai_mai_n273_), .B(mai_mai_n153_), .C(mai_mai_n104_), .Y(mai_mai_n303_));
  NAi21      m281(.An(i_8_), .B(i_7_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n304_), .B(i_6_), .Y(mai_mai_n305_));
  NO2        m283(.A(mai_mai_n147_), .B(mai_mai_n46_), .Y(mai_mai_n306_));
  NA3        m284(.A(mai_mai_n306_), .B(mai_mai_n305_), .C(mai_mai_n153_), .Y(mai_mai_n307_));
  NA3        m285(.A(mai_mai_n307_), .B(mai_mai_n303_), .C(mai_mai_n302_), .Y(mai_mai_n308_));
  OAI210     m286(.A0(mai_mai_n308_), .A1(mai_mai_n298_), .B0(i_4_), .Y(mai_mai_n309_));
  NO2        m287(.A(i_12_), .B(i_10_), .Y(mai_mai_n310_));
  NOi21      m288(.An(i_5_), .B(i_0_), .Y(mai_mai_n311_));
  NO3        m289(.A(mai_mai_n286_), .B(mai_mai_n311_), .C(mai_mai_n120_), .Y(mai_mai_n312_));
  NA4        m290(.A(mai_mai_n74_), .B(mai_mai_n36_), .C(mai_mai_n76_), .D(i_8_), .Y(mai_mai_n313_));
  NA2        m291(.A(mai_mai_n312_), .B(mai_mai_n310_), .Y(mai_mai_n314_));
  NO2        m292(.A(i_6_), .B(i_8_), .Y(mai_mai_n315_));
  AN2        m293(.A(i_0_), .B(mai_mai_n315_), .Y(mai_mai_n316_));
  NO2        m294(.A(i_1_), .B(i_7_), .Y(mai_mai_n317_));
  AO220      m295(.A0(mai_mai_n317_), .A1(mai_mai_n316_), .B0(mai_mai_n305_), .B1(mai_mai_n223_), .Y(mai_mai_n318_));
  NA2        m296(.A(mai_mai_n318_), .B(i_4_), .Y(mai_mai_n319_));
  NA3        m297(.A(mai_mai_n319_), .B(mai_mai_n314_), .C(mai_mai_n309_), .Y(mai_mai_n320_));
  NO3        m298(.A(mai_mai_n221_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n321_));
  NO3        m299(.A(mai_mai_n304_), .B(i_2_), .C(i_1_), .Y(mai_mai_n322_));
  OAI210     m300(.A0(mai_mai_n322_), .A1(mai_mai_n321_), .B0(i_6_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n240_), .B(mai_mai_n285_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n324_), .B(mai_mai_n323_), .Y(mai_mai_n325_));
  NA2        m303(.A(mai_mai_n325_), .B(i_3_), .Y(mai_mai_n326_));
  INV        m304(.A(mai_mai_n74_), .Y(mai_mai_n327_));
  NA2        m305(.A(i_2_), .B(mai_mai_n124_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n85_), .B(mai_mai_n182_), .Y(mai_mai_n329_));
  AOI210     m307(.A0(mai_mai_n85_), .A1(mai_mai_n328_), .B0(mai_mai_n327_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n182_), .B(i_9_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n331_), .B(mai_mai_n195_), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n330_), .B(mai_mai_n276_), .Y(mai_mai_n333_));
  AOI210     m311(.A0(mai_mai_n333_), .A1(mai_mai_n326_), .B0(mai_mai_n152_), .Y(mai_mai_n334_));
  AOI210     m312(.A0(mai_mai_n320_), .A1(mai_mai_n296_), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  NOi32      m313(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n336_));
  INV        m314(.A(mai_mai_n336_), .Y(mai_mai_n337_));
  NAi21      m315(.An(i_0_), .B(i_6_), .Y(mai_mai_n338_));
  NAi21      m316(.An(i_1_), .B(i_5_), .Y(mai_mai_n339_));
  NA2        m317(.A(mai_mai_n339_), .B(mai_mai_n338_), .Y(mai_mai_n340_));
  NA2        m318(.A(mai_mai_n340_), .B(mai_mai_n25_), .Y(mai_mai_n341_));
  OAI210     m319(.A0(mai_mai_n341_), .A1(mai_mai_n149_), .B0(mai_mai_n234_), .Y(mai_mai_n342_));
  NAi41      m320(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n343_));
  OAI220     m321(.A0(mai_mai_n343_), .A1(mai_mai_n339_), .B0(mai_mai_n209_), .B1(mai_mai_n149_), .Y(mai_mai_n344_));
  AOI210     m322(.A0(mai_mai_n343_), .A1(mai_mai_n149_), .B0(mai_mai_n147_), .Y(mai_mai_n345_));
  OR2        m323(.A(mai_mai_n345_), .B(mai_mai_n344_), .Y(mai_mai_n346_));
  NO2        m324(.A(i_1_), .B(mai_mai_n93_), .Y(mai_mai_n347_));
  NAi21      m325(.An(i_3_), .B(i_4_), .Y(mai_mai_n348_));
  NA2        m326(.A(i_2_), .B(i_7_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n348_), .B(i_10_), .Y(mai_mai_n350_));
  AOI210     m328(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n351_));
  OAI210     m329(.A0(mai_mai_n351_), .A1(mai_mai_n177_), .B0(mai_mai_n350_), .Y(mai_mai_n352_));
  AOI220     m330(.A0(mai_mai_n350_), .A1(mai_mai_n317_), .B0(mai_mai_n226_), .B1(mai_mai_n177_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n352_), .B0(i_5_), .Y(mai_mai_n354_));
  NO3        m332(.A(mai_mai_n354_), .B(mai_mai_n346_), .C(mai_mai_n342_), .Y(mai_mai_n355_));
  NO2        m333(.A(mai_mai_n355_), .B(mai_mai_n337_), .Y(mai_mai_n356_));
  NO2        m334(.A(mai_mai_n56_), .B(mai_mai_n25_), .Y(mai_mai_n357_));
  AN2        m335(.A(i_12_), .B(i_5_), .Y(mai_mai_n358_));
  NO2        m336(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n360_));
  NO2        m338(.A(i_11_), .B(i_6_), .Y(mai_mai_n361_));
  NA3        m339(.A(mai_mai_n361_), .B(mai_mai_n306_), .C(mai_mai_n213_), .Y(mai_mai_n362_));
  NO2        m340(.A(mai_mai_n362_), .B(mai_mai_n360_), .Y(mai_mai_n363_));
  NO2        m341(.A(mai_mai_n230_), .B(i_5_), .Y(mai_mai_n364_));
  NO2        m342(.A(i_5_), .B(i_10_), .Y(mai_mai_n365_));
  AOI220     m343(.A0(mai_mai_n365_), .A1(mai_mai_n253_), .B0(mai_mai_n364_), .B1(mai_mai_n187_), .Y(mai_mai_n366_));
  NA2        m344(.A(mai_mai_n135_), .B(mai_mai_n45_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n367_), .B(mai_mai_n366_), .Y(mai_mai_n368_));
  OAI210     m346(.A0(mai_mai_n368_), .A1(mai_mai_n363_), .B0(mai_mai_n357_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n370_));
  NO2        m348(.A(mai_mai_n141_), .B(mai_mai_n76_), .Y(mai_mai_n371_));
  OAI210     m349(.A0(mai_mai_n371_), .A1(mai_mai_n363_), .B0(mai_mai_n370_), .Y(mai_mai_n372_));
  NO3        m350(.A(mai_mai_n76_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n373_));
  NA3        m351(.A(mai_mai_n283_), .B(mai_mai_n83_), .C(mai_mai_n53_), .Y(mai_mai_n374_));
  NO2        m352(.A(mai_mai_n374_), .B(i_12_), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n365_), .B(mai_mai_n224_), .Y(mai_mai_n376_));
  NO2        m354(.A(mai_mai_n36_), .B(mai_mai_n209_), .Y(mai_mai_n377_));
  NAi21      m355(.An(i_13_), .B(i_0_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(mai_mai_n227_), .Y(mai_mai_n379_));
  OAI210     m357(.A0(mai_mai_n377_), .A1(mai_mai_n375_), .B0(mai_mai_n379_), .Y(mai_mai_n380_));
  NA3        m358(.A(mai_mai_n380_), .B(mai_mai_n372_), .C(mai_mai_n369_), .Y(mai_mai_n381_));
  NA2        m359(.A(mai_mai_n44_), .B(mai_mai_n213_), .Y(mai_mai_n382_));
  NO2        m360(.A(i_0_), .B(i_11_), .Y(mai_mai_n383_));
  INV        m361(.A(i_5_), .Y(mai_mai_n384_));
  AN2        m362(.A(i_1_), .B(i_6_), .Y(mai_mai_n385_));
  NOi21      m363(.An(i_2_), .B(i_12_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n386_), .B(mai_mai_n385_), .Y(mai_mai_n387_));
  NO2        m365(.A(mai_mai_n387_), .B(mai_mai_n384_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n133_), .B(i_9_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n389_), .B(i_4_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n388_), .B(mai_mai_n390_), .Y(mai_mai_n391_));
  NAi21      m369(.An(i_9_), .B(i_4_), .Y(mai_mai_n392_));
  OR2        m370(.A(i_13_), .B(i_10_), .Y(mai_mai_n393_));
  NO3        m371(.A(mai_mai_n393_), .B(mai_mai_n109_), .C(mai_mai_n392_), .Y(mai_mai_n394_));
  BUFFER     m372(.A(mai_mai_n205_), .Y(mai_mai_n395_));
  NO2        m373(.A(mai_mai_n93_), .B(mai_mai_n25_), .Y(mai_mai_n396_));
  NA2        m374(.A(mai_mai_n259_), .B(mai_mai_n200_), .Y(mai_mai_n397_));
  NO2        m375(.A(mai_mai_n397_), .B(mai_mai_n395_), .Y(mai_mai_n398_));
  INV        m376(.A(mai_mai_n398_), .Y(mai_mai_n399_));
  AOI210     m377(.A0(mai_mai_n399_), .A1(mai_mai_n391_), .B0(mai_mai_n26_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n303_), .B(mai_mai_n302_), .Y(mai_mai_n401_));
  AOI220     m379(.A0(mai_mai_n279_), .A1(mai_mai_n269_), .B0(mai_mai_n273_), .B1(i_6_), .Y(mai_mai_n402_));
  NO2        m380(.A(mai_mai_n402_), .B(mai_mai_n159_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n172_), .B(mai_mai_n76_), .Y(mai_mai_n404_));
  AOI220     m382(.A0(mai_mai_n404_), .A1(mai_mai_n278_), .B0(mai_mai_n261_), .B1(mai_mai_n200_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n405_), .B(mai_mai_n268_), .Y(mai_mai_n406_));
  NO3        m384(.A(mai_mai_n406_), .B(mai_mai_n403_), .C(mai_mai_n401_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n185_), .B(mai_mai_n88_), .Y(mai_mai_n408_));
  NA3        m386(.A(mai_mai_n306_), .B(mai_mai_n153_), .C(mai_mai_n76_), .Y(mai_mai_n409_));
  AOI210     m387(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(mai_mai_n304_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n279_), .B(mai_mai_n223_), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n411_), .B(mai_mai_n172_), .Y(mai_mai_n412_));
  NA3        m390(.A(mai_mai_n317_), .B(mai_mai_n316_), .C(i_5_), .Y(mai_mai_n413_));
  INV        m391(.A(mai_mai_n297_), .Y(mai_mai_n414_));
  OAI210     m392(.A0(mai_mai_n414_), .A1(mai_mai_n178_), .B0(mai_mai_n413_), .Y(mai_mai_n415_));
  NO3        m393(.A(mai_mai_n415_), .B(mai_mai_n412_), .C(mai_mai_n410_), .Y(mai_mai_n416_));
  AOI210     m394(.A0(mai_mai_n416_), .A1(mai_mai_n407_), .B0(mai_mai_n255_), .Y(mai_mai_n417_));
  NO4        m395(.A(mai_mai_n417_), .B(mai_mai_n400_), .C(mai_mai_n381_), .D(mai_mai_n356_), .Y(mai_mai_n418_));
  NO2        m396(.A(i_10_), .B(i_9_), .Y(mai_mai_n419_));
  NAi21      m397(.An(i_12_), .B(i_8_), .Y(mai_mai_n420_));
  NO2        m398(.A(mai_mai_n420_), .B(i_3_), .Y(mai_mai_n421_));
  NA2        m399(.A(i_2_), .B(mai_mai_n96_), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n422_), .B(mai_mai_n194_), .Y(mai_mai_n423_));
  NA2        m401(.A(mai_mai_n292_), .B(i_0_), .Y(mai_mai_n424_));
  NO3        m402(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n425_));
  NA2        m403(.A(mai_mai_n250_), .B(mai_mai_n89_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n426_), .B(mai_mai_n425_), .Y(mai_mai_n427_));
  NA2        m405(.A(i_8_), .B(i_9_), .Y(mai_mai_n428_));
  NO2        m406(.A(i_7_), .B(i_2_), .Y(mai_mai_n429_));
  OR2        m407(.A(mai_mai_n429_), .B(mai_mai_n428_), .Y(mai_mai_n430_));
  NA2        m408(.A(mai_mai_n266_), .B(mai_mai_n195_), .Y(mai_mai_n431_));
  NO2        m409(.A(mai_mai_n431_), .B(mai_mai_n430_), .Y(mai_mai_n432_));
  NA2        m410(.A(mai_mai_n239_), .B(mai_mai_n291_), .Y(mai_mai_n433_));
  NO3        m411(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n434_));
  INV        m412(.A(mai_mai_n434_), .Y(mai_mai_n435_));
  NA3        m413(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n436_));
  NA4        m414(.A(mai_mai_n136_), .B(mai_mai_n107_), .C(mai_mai_n72_), .D(mai_mai_n23_), .Y(mai_mai_n437_));
  OAI220     m415(.A0(mai_mai_n437_), .A1(mai_mai_n436_), .B0(mai_mai_n435_), .B1(mai_mai_n433_), .Y(mai_mai_n438_));
  NO3        m416(.A(mai_mai_n438_), .B(mai_mai_n432_), .C(mai_mai_n423_), .Y(mai_mai_n439_));
  OR2        m417(.A(mai_mai_n277_), .B(mai_mai_n197_), .Y(mai_mai_n440_));
  OA210      m418(.A0(mai_mai_n332_), .A1(mai_mai_n93_), .B0(mai_mai_n280_), .Y(mai_mai_n441_));
  OA220      m419(.A0(mai_mai_n441_), .A1(mai_mai_n152_), .B0(mai_mai_n440_), .B1(mai_mai_n220_), .Y(mai_mai_n442_));
  NA2        m420(.A(mai_mai_n88_), .B(i_13_), .Y(mai_mai_n443_));
  NA2        m421(.A(mai_mai_n404_), .B(mai_mai_n357_), .Y(mai_mai_n444_));
  NO2        m422(.A(i_2_), .B(i_13_), .Y(mai_mai_n445_));
  NO2        m423(.A(mai_mai_n444_), .B(mai_mai_n443_), .Y(mai_mai_n446_));
  NO3        m424(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n447_));
  NO2        m425(.A(i_6_), .B(i_7_), .Y(mai_mai_n448_));
  NA2        m426(.A(mai_mai_n448_), .B(mai_mai_n447_), .Y(mai_mai_n449_));
  NO2        m427(.A(i_11_), .B(i_1_), .Y(mai_mai_n450_));
  NOi21      m428(.An(i_2_), .B(i_7_), .Y(mai_mai_n451_));
  NO2        m429(.A(i_3_), .B(mai_mai_n182_), .Y(mai_mai_n452_));
  NO2        m430(.A(i_6_), .B(i_10_), .Y(mai_mai_n453_));
  NA3        m431(.A(mai_mai_n453_), .B(mai_mai_n296_), .C(mai_mai_n452_), .Y(mai_mai_n454_));
  NO2        m432(.A(mai_mai_n454_), .B(mai_mai_n145_), .Y(mai_mai_n455_));
  NA2        m433(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n456_));
  NO2        m434(.A(mai_mai_n147_), .B(i_3_), .Y(mai_mai_n457_));
  NAi31      m435(.An(mai_mai_n456_), .B(mai_mai_n457_), .C(mai_mai_n214_), .Y(mai_mai_n458_));
  NA3        m436(.A(mai_mai_n370_), .B(mai_mai_n169_), .C(mai_mai_n140_), .Y(mai_mai_n459_));
  NA2        m437(.A(mai_mai_n459_), .B(mai_mai_n458_), .Y(mai_mai_n460_));
  NO3        m438(.A(mai_mai_n460_), .B(mai_mai_n455_), .C(mai_mai_n446_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n425_), .B(mai_mai_n358_), .Y(mai_mai_n462_));
  NA2        m440(.A(mai_mai_n434_), .B(mai_mai_n365_), .Y(mai_mai_n463_));
  NO2        m441(.A(mai_mai_n463_), .B(mai_mai_n212_), .Y(mai_mai_n464_));
  NO2        m442(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n465_));
  NA3        m443(.A(mai_mai_n966_), .B(mai_mai_n465_), .C(mai_mai_n133_), .Y(mai_mai_n466_));
  OR3        m444(.A(mai_mai_n286_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n467_));
  NO2        m445(.A(mai_mai_n467_), .B(mai_mai_n466_), .Y(mai_mai_n468_));
  NA2        m446(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n469_));
  NO2        m447(.A(mai_mai_n469_), .B(mai_mai_n443_), .Y(mai_mai_n470_));
  NA3        m448(.A(mai_mai_n289_), .B(mai_mai_n211_), .C(mai_mai_n65_), .Y(mai_mai_n471_));
  NO2        m449(.A(mai_mai_n471_), .B(mai_mai_n449_), .Y(mai_mai_n472_));
  NO4        m450(.A(mai_mai_n472_), .B(mai_mai_n470_), .C(mai_mai_n468_), .D(mai_mai_n464_), .Y(mai_mai_n473_));
  NA4        m451(.A(mai_mai_n473_), .B(mai_mai_n461_), .C(mai_mai_n442_), .D(mai_mai_n439_), .Y(mai_mai_n474_));
  AN2        m452(.A(mai_mai_n269_), .B(mai_mai_n222_), .Y(mai_mai_n475_));
  NA2        m453(.A(mai_mai_n475_), .B(mai_mai_n166_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n114_), .B(mai_mai_n103_), .Y(mai_mai_n477_));
  AN2        m455(.A(mai_mai_n477_), .B(mai_mai_n425_), .Y(mai_mai_n478_));
  NA2        m456(.A(mai_mai_n296_), .B(mai_mai_n154_), .Y(mai_mai_n479_));
  OAI210     m457(.A0(mai_mai_n479_), .A1(mai_mai_n220_), .B0(mai_mai_n290_), .Y(mai_mai_n480_));
  AOI220     m458(.A0(mai_mai_n480_), .A1(mai_mai_n305_), .B0(mai_mai_n478_), .B1(mai_mai_n292_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n336_), .B(mai_mai_n65_), .Y(mai_mai_n482_));
  NO2        m460(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n483_));
  AOI210     m461(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n394_), .Y(mai_mai_n484_));
  NO2        m462(.A(i_7_), .B(mai_mai_n188_), .Y(mai_mai_n485_));
  OR2        m463(.A(mai_mai_n172_), .B(i_4_), .Y(mai_mai_n486_));
  INV        m464(.A(mai_mai_n486_), .Y(mai_mai_n487_));
  NA2        m465(.A(mai_mai_n487_), .B(mai_mai_n485_), .Y(mai_mai_n488_));
  NA4        m466(.A(mai_mai_n488_), .B(mai_mai_n484_), .C(mai_mai_n481_), .D(mai_mai_n476_), .Y(mai_mai_n489_));
  NA2        m467(.A(mai_mai_n364_), .B(mai_mai_n278_), .Y(mai_mai_n490_));
  NA2        m468(.A(mai_mai_n360_), .B(mai_mai_n490_), .Y(mai_mai_n491_));
  NO2        m469(.A(i_12_), .B(mai_mai_n182_), .Y(mai_mai_n492_));
  NA2        m470(.A(mai_mai_n453_), .B(mai_mai_n27_), .Y(mai_mai_n493_));
  NO2        m471(.A(mai_mai_n493_), .B(i_12_), .Y(mai_mai_n494_));
  NOi31      m472(.An(mai_mai_n297_), .B(mai_mai_n393_), .C(mai_mai_n38_), .Y(mai_mai_n495_));
  OAI210     m473(.A0(mai_mai_n495_), .A1(mai_mai_n494_), .B0(mai_mai_n491_), .Y(mai_mai_n496_));
  NO2        m474(.A(i_8_), .B(i_7_), .Y(mai_mai_n497_));
  OAI210     m475(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n498_));
  NA2        m476(.A(mai_mai_n498_), .B(mai_mai_n211_), .Y(mai_mai_n499_));
  OAI220     m477(.A0(mai_mai_n46_), .A1(mai_mai_n486_), .B0(mai_mai_n499_), .B1(mai_mai_n230_), .Y(mai_mai_n500_));
  NA2        m478(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n501_));
  NO2        m479(.A(mai_mai_n501_), .B(i_6_), .Y(mai_mai_n502_));
  NA3        m480(.A(mai_mai_n502_), .B(mai_mai_n500_), .C(mai_mai_n497_), .Y(mai_mai_n503_));
  AOI220     m481(.A0(mai_mai_n404_), .A1(mai_mai_n306_), .B0(mai_mai_n235_), .B1(mai_mai_n232_), .Y(mai_mai_n504_));
  OAI220     m482(.A0(mai_mai_n504_), .A1(mai_mai_n246_), .B0(mai_mai_n443_), .B1(mai_mai_n125_), .Y(mai_mai_n505_));
  NA2        m483(.A(mai_mai_n505_), .B(mai_mai_n249_), .Y(mai_mai_n506_));
  NA3        m484(.A(mai_mai_n289_), .B(mai_mai_n164_), .C(mai_mai_n88_), .Y(mai_mai_n507_));
  NO2        m485(.A(mai_mai_n210_), .B(mai_mai_n44_), .Y(mai_mai_n508_));
  NO2        m486(.A(mai_mai_n147_), .B(i_5_), .Y(mai_mai_n509_));
  NA3        m487(.A(mai_mai_n509_), .B(mai_mai_n382_), .C(mai_mai_n299_), .Y(mai_mai_n510_));
  OAI210     m488(.A0(mai_mai_n510_), .A1(mai_mai_n508_), .B0(mai_mai_n507_), .Y(mai_mai_n511_));
  NA2        m489(.A(mai_mai_n511_), .B(mai_mai_n434_), .Y(mai_mai_n512_));
  NA4        m490(.A(mai_mai_n512_), .B(mai_mai_n506_), .C(mai_mai_n503_), .D(mai_mai_n496_), .Y(mai_mai_n513_));
  NA3        m491(.A(mai_mai_n207_), .B(mai_mai_n63_), .C(mai_mai_n44_), .Y(mai_mai_n514_));
  NA2        m492(.A(mai_mai_n266_), .B(mai_mai_n74_), .Y(mai_mai_n515_));
  AOI210     m493(.A0(mai_mai_n514_), .A1(mai_mai_n328_), .B0(mai_mai_n515_), .Y(mai_mai_n516_));
  NO2        m494(.A(mai_mai_n46_), .B(mai_mai_n163_), .Y(mai_mai_n517_));
  AOI210     m495(.A0(i_6_), .A1(mai_mai_n46_), .B0(mai_mai_n347_), .Y(mai_mai_n518_));
  NA2        m496(.A(i_0_), .B(mai_mai_n48_), .Y(mai_mai_n519_));
  NA3        m497(.A(mai_mai_n492_), .B(mai_mai_n257_), .C(mai_mai_n519_), .Y(mai_mai_n520_));
  NO2        m498(.A(mai_mai_n518_), .B(mai_mai_n520_), .Y(mai_mai_n521_));
  NO3        m499(.A(mai_mai_n521_), .B(mai_mai_n517_), .C(mai_mai_n516_), .Y(mai_mai_n522_));
  NO4        m500(.A(mai_mai_n240_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n523_));
  NO3        m501(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n524_));
  NO2        m502(.A(mai_mai_n221_), .B(mai_mai_n36_), .Y(mai_mai_n525_));
  AN2        m503(.A(mai_mai_n525_), .B(mai_mai_n524_), .Y(mai_mai_n526_));
  OA210      m504(.A0(mai_mai_n526_), .A1(mai_mai_n523_), .B0(mai_mai_n336_), .Y(mai_mai_n527_));
  NO2        m505(.A(mai_mai_n393_), .B(i_1_), .Y(mai_mai_n528_));
  NOi31      m506(.An(mai_mai_n528_), .B(mai_mai_n426_), .C(mai_mai_n65_), .Y(mai_mai_n529_));
  AN4        m507(.A(mai_mai_n529_), .B(mai_mai_n390_), .C(mai_mai_n465_), .D(i_2_), .Y(mai_mai_n530_));
  NO2        m508(.A(mai_mai_n402_), .B(mai_mai_n167_), .Y(mai_mai_n531_));
  NO3        m509(.A(mai_mai_n531_), .B(mai_mai_n530_), .C(mai_mai_n527_), .Y(mai_mai_n532_));
  NOi21      m510(.An(i_10_), .B(i_6_), .Y(mai_mai_n533_));
  NO2        m511(.A(mai_mai_n76_), .B(mai_mai_n25_), .Y(mai_mai_n534_));
  AOI220     m512(.A0(mai_mai_n266_), .A1(mai_mai_n534_), .B0(mai_mai_n257_), .B1(mai_mai_n533_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n535_), .B(mai_mai_n424_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n106_), .B(mai_mai_n23_), .Y(mai_mai_n537_));
  NA2        m515(.A(mai_mai_n297_), .B(mai_mai_n154_), .Y(mai_mai_n538_));
  AOI220     m516(.A0(mai_mai_n538_), .A1(mai_mai_n411_), .B0(mai_mai_n162_), .B1(mai_mai_n171_), .Y(mai_mai_n539_));
  NO2        m517(.A(mai_mai_n187_), .B(mai_mai_n37_), .Y(mai_mai_n540_));
  NOi31      m518(.An(mai_mai_n137_), .B(mai_mai_n540_), .C(mai_mai_n313_), .Y(mai_mai_n541_));
  NO3        m519(.A(mai_mai_n541_), .B(mai_mai_n539_), .C(mai_mai_n536_), .Y(mai_mai_n542_));
  NO2        m520(.A(mai_mai_n482_), .B(mai_mai_n353_), .Y(mai_mai_n543_));
  NO2        m521(.A(i_12_), .B(mai_mai_n76_), .Y(mai_mai_n544_));
  NO3        m522(.A(i_4_), .B(mai_mai_n323_), .C(mai_mai_n284_), .Y(mai_mai_n545_));
  NO2        m523(.A(mai_mai_n545_), .B(mai_mai_n543_), .Y(mai_mai_n546_));
  NA4        m524(.A(mai_mai_n546_), .B(mai_mai_n542_), .C(mai_mai_n532_), .D(mai_mai_n522_), .Y(mai_mai_n547_));
  NO4        m525(.A(mai_mai_n547_), .B(mai_mai_n513_), .C(mai_mai_n489_), .D(mai_mai_n474_), .Y(mai_mai_n548_));
  NA4        m526(.A(mai_mai_n548_), .B(mai_mai_n418_), .C(mai_mai_n335_), .D(mai_mai_n295_), .Y(mai7));
  NO2        m527(.A(mai_mai_n100_), .B(mai_mai_n82_), .Y(mai_mai_n550_));
  NA2        m528(.A(mai_mai_n453_), .B(mai_mai_n74_), .Y(mai_mai_n551_));
  NA2        m529(.A(i_11_), .B(mai_mai_n182_), .Y(mai_mai_n552_));
  NA3        m530(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n224_), .B(i_4_), .Y(mai_mai_n554_));
  NA2        m532(.A(mai_mai_n554_), .B(i_8_), .Y(mai_mai_n555_));
  NO2        m533(.A(mai_mai_n97_), .B(mai_mai_n553_), .Y(mai_mai_n556_));
  NA2        m534(.A(i_2_), .B(mai_mai_n76_), .Y(mai_mai_n557_));
  OAI210     m535(.A0(mai_mai_n79_), .A1(mai_mai_n192_), .B0(mai_mai_n193_), .Y(mai_mai_n558_));
  NO2        m536(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n559_));
  NO2        m537(.A(mai_mai_n558_), .B(i_13_), .Y(mai_mai_n560_));
  NO3        m538(.A(mai_mai_n560_), .B(mai_mai_n556_), .C(mai_mai_n550_), .Y(mai_mai_n561_));
  AOI210     m539(.A0(mai_mai_n120_), .A1(mai_mai_n57_), .B0(i_10_), .Y(mai_mai_n562_));
  AOI210     m540(.A0(mai_mai_n562_), .A1(mai_mai_n224_), .B0(mai_mai_n151_), .Y(mai_mai_n563_));
  OR2        m541(.A(i_6_), .B(i_10_), .Y(mai_mai_n564_));
  NO2        m542(.A(mai_mai_n564_), .B(mai_mai_n23_), .Y(mai_mai_n565_));
  OR3        m543(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n566_));
  NO3        m544(.A(mai_mai_n566_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n567_));
  INV        m545(.A(mai_mai_n189_), .Y(mai_mai_n568_));
  NO2        m546(.A(mai_mai_n567_), .B(mai_mai_n565_), .Y(mai_mai_n569_));
  OA220      m547(.A0(mai_mai_n569_), .A1(i_2_), .B0(mai_mai_n563_), .B1(mai_mai_n251_), .Y(mai_mai_n570_));
  AOI210     m548(.A0(mai_mai_n570_), .A1(mai_mai_n561_), .B0(mai_mai_n58_), .Y(mai_mai_n571_));
  NOi21      m549(.An(i_11_), .B(i_7_), .Y(mai_mai_n572_));
  AO210      m550(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n573_));
  NO2        m551(.A(mai_mai_n573_), .B(mai_mai_n572_), .Y(mai_mai_n574_));
  NA2        m552(.A(mai_mai_n574_), .B(mai_mai_n196_), .Y(mai_mai_n575_));
  NA3        m553(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n576_));
  NAi31      m554(.An(mai_mai_n576_), .B(i_12_), .C(i_11_), .Y(mai_mai_n577_));
  AOI210     m555(.A0(mai_mai_n577_), .A1(mai_mai_n575_), .B0(mai_mai_n58_), .Y(mai_mai_n578_));
  NA2        m556(.A(mai_mai_n78_), .B(mai_mai_n58_), .Y(mai_mai_n579_));
  AO210      m557(.A0(mai_mai_n579_), .A1(mai_mai_n353_), .B0(mai_mai_n41_), .Y(mai_mai_n580_));
  NA2        m558(.A(mai_mai_n214_), .B(mai_mai_n58_), .Y(mai_mai_n581_));
  NO2        m559(.A(mai_mai_n58_), .B(i_9_), .Y(mai_mai_n582_));
  NO2        m560(.A(i_1_), .B(i_12_), .Y(mai_mai_n583_));
  NA2        m561(.A(mai_mai_n581_), .B(mai_mai_n580_), .Y(mai_mai_n584_));
  OAI210     m562(.A0(mai_mai_n584_), .A1(mai_mai_n578_), .B0(i_6_), .Y(mai_mai_n585_));
  NO2        m563(.A(mai_mai_n576_), .B(mai_mai_n100_), .Y(mai_mai_n586_));
  NA2        m564(.A(mai_mai_n586_), .B(mai_mai_n544_), .Y(mai_mai_n587_));
  NO2        m565(.A(mai_mai_n224_), .B(mai_mai_n76_), .Y(mai_mai_n588_));
  NO2        m566(.A(mai_mai_n588_), .B(i_11_), .Y(mai_mai_n589_));
  NA2        m567(.A(mai_mai_n587_), .B(mai_mai_n427_), .Y(mai_mai_n590_));
  NO4        m568(.A(i_12_), .B(mai_mai_n120_), .C(i_13_), .D(mai_mai_n76_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n591_), .B(mai_mai_n582_), .Y(mai_mai_n592_));
  NA2        m570(.A(mai_mai_n224_), .B(i_6_), .Y(mai_mai_n593_));
  INV        m571(.A(mai_mai_n592_), .Y(mai_mai_n594_));
  NA3        m572(.A(mai_mai_n497_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n129_), .B(i_9_), .Y(mai_mai_n596_));
  NA2        m574(.A(i_3_), .B(i_9_), .Y(mai_mai_n597_));
  NO2        m575(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n598_));
  NO2        m576(.A(mai_mai_n596_), .B(mai_mai_n964_), .Y(mai_mai_n599_));
  NA3        m577(.A(mai_mai_n582_), .B(mai_mai_n299_), .C(i_6_), .Y(mai_mai_n600_));
  NO2        m578(.A(mai_mai_n600_), .B(mai_mai_n23_), .Y(mai_mai_n601_));
  AOI210     m579(.A0(mai_mai_n450_), .A1(mai_mai_n396_), .B0(mai_mai_n229_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n602_), .B(mai_mai_n557_), .Y(mai_mai_n603_));
  NA2        m581(.A(mai_mai_n598_), .B(mai_mai_n250_), .Y(mai_mai_n604_));
  NO2        m582(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n605_));
  NA2        m583(.A(mai_mai_n605_), .B(mai_mai_n24_), .Y(mai_mai_n606_));
  NO2        m584(.A(mai_mai_n606_), .B(mai_mai_n604_), .Y(mai_mai_n607_));
  OR4        m585(.A(mai_mai_n607_), .B(mai_mai_n603_), .C(mai_mai_n601_), .D(mai_mai_n599_), .Y(mai_mai_n608_));
  NO3        m586(.A(mai_mai_n608_), .B(mai_mai_n594_), .C(mai_mai_n590_), .Y(mai_mai_n609_));
  NO2        m587(.A(mai_mai_n224_), .B(mai_mai_n93_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n610_), .B(mai_mai_n572_), .Y(mai_mai_n611_));
  NO2        m589(.A(mai_mai_n392_), .B(mai_mai_n76_), .Y(mai_mai_n612_));
  NO2        m590(.A(mai_mai_n221_), .B(mai_mai_n44_), .Y(mai_mai_n613_));
  NO3        m591(.A(mai_mai_n613_), .B(mai_mai_n292_), .C(mai_mai_n225_), .Y(mai_mai_n614_));
  NO2        m592(.A(mai_mai_n109_), .B(mai_mai_n37_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n615_), .B(i_6_), .Y(mai_mai_n616_));
  NO2        m594(.A(mai_mai_n76_), .B(i_9_), .Y(mai_mai_n617_));
  NO2        m595(.A(mai_mai_n617_), .B(mai_mai_n58_), .Y(mai_mai_n618_));
  NO2        m596(.A(mai_mai_n618_), .B(mai_mai_n583_), .Y(mai_mai_n619_));
  NO4        m597(.A(mai_mai_n619_), .B(mai_mai_n616_), .C(mai_mai_n614_), .D(i_4_), .Y(mai_mai_n620_));
  NA2        m598(.A(i_1_), .B(i_3_), .Y(mai_mai_n621_));
  INV        m599(.A(mai_mai_n620_), .Y(mai_mai_n622_));
  NA3        m600(.A(mai_mai_n622_), .B(mai_mai_n609_), .C(mai_mai_n585_), .Y(mai_mai_n623_));
  NO3        m601(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n624_));
  NOi21      m602(.An(mai_mai_n624_), .B(i_10_), .Y(mai_mai_n625_));
  OA210      m603(.A0(mai_mai_n625_), .A1(mai_mai_n233_), .B0(mai_mai_n76_), .Y(mai_mai_n626_));
  NA2        m604(.A(mai_mai_n626_), .B(i_1_), .Y(mai_mai_n627_));
  AOI210     m605(.A0(mai_mai_n250_), .A1(mai_mai_n89_), .B0(i_1_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n348_), .B(i_2_), .Y(mai_mai_n629_));
  NA2        m607(.A(mai_mai_n629_), .B(mai_mai_n628_), .Y(mai_mai_n630_));
  AOI210     m608(.A0(mai_mai_n630_), .A1(mai_mai_n627_), .B0(i_13_), .Y(mai_mai_n631_));
  OR2        m609(.A(i_11_), .B(i_7_), .Y(mai_mai_n632_));
  NA3        m610(.A(mai_mai_n632_), .B(mai_mai_n98_), .C(mai_mai_n129_), .Y(mai_mai_n633_));
  AOI220     m611(.A0(mai_mai_n445_), .A1(mai_mai_n151_), .B0(i_2_), .B1(mai_mai_n129_), .Y(mai_mai_n634_));
  OAI210     m612(.A0(mai_mai_n634_), .A1(mai_mai_n44_), .B0(mai_mai_n633_), .Y(mai_mai_n635_));
  NO2        m613(.A(mai_mai_n53_), .B(i_12_), .Y(mai_mai_n636_));
  INV        m614(.A(mai_mai_n636_), .Y(mai_mai_n637_));
  NO2        m615(.A(mai_mai_n451_), .B(mai_mai_n24_), .Y(mai_mai_n638_));
  NA2        m616(.A(mai_mai_n638_), .B(mai_mai_n612_), .Y(mai_mai_n639_));
  OAI220     m617(.A0(mai_mai_n639_), .A1(mai_mai_n41_), .B0(mai_mai_n637_), .B1(mai_mai_n85_), .Y(mai_mai_n640_));
  AOI210     m618(.A0(mai_mai_n635_), .A1(mai_mai_n315_), .B0(mai_mai_n640_), .Y(mai_mai_n641_));
  INV        m619(.A(mai_mai_n106_), .Y(mai_mai_n642_));
  AOI220     m620(.A0(mai_mai_n642_), .A1(mai_mai_n64_), .B0(mai_mai_n361_), .B1(mai_mai_n598_), .Y(mai_mai_n643_));
  NO2        m621(.A(mai_mai_n643_), .B(mai_mai_n230_), .Y(mai_mai_n644_));
  AOI210     m622(.A0(mai_mai_n420_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n645_));
  NOi31      m623(.An(mai_mai_n645_), .B(mai_mai_n551_), .C(mai_mai_n44_), .Y(mai_mai_n646_));
  NA2        m624(.A(mai_mai_n119_), .B(i_13_), .Y(mai_mai_n647_));
  NO2        m625(.A(mai_mai_n597_), .B(mai_mai_n106_), .Y(mai_mai_n648_));
  INV        m626(.A(mai_mai_n648_), .Y(mai_mai_n649_));
  NO2        m627(.A(mai_mai_n647_), .B(mai_mai_n628_), .Y(mai_mai_n650_));
  AOI220     m628(.A0(mai_mai_n361_), .A1(mai_mai_n598_), .B0(mai_mai_n84_), .B1(mai_mai_n94_), .Y(mai_mai_n651_));
  NO2        m629(.A(mai_mai_n651_), .B(mai_mai_n555_), .Y(mai_mai_n652_));
  NO4        m630(.A(mai_mai_n652_), .B(mai_mai_n650_), .C(mai_mai_n646_), .D(mai_mai_n644_), .Y(mai_mai_n653_));
  OR2        m631(.A(i_11_), .B(i_6_), .Y(mai_mai_n654_));
  NA2        m632(.A(mai_mai_n554_), .B(i_7_), .Y(mai_mai_n655_));
  AOI210     m633(.A0(mai_mai_n655_), .A1(mai_mai_n649_), .B0(mai_mai_n654_), .Y(mai_mai_n656_));
  NA3        m634(.A(mai_mai_n386_), .B(mai_mai_n559_), .C(mai_mai_n89_), .Y(mai_mai_n657_));
  NA2        m635(.A(mai_mai_n589_), .B(i_13_), .Y(mai_mai_n658_));
  NAi21      m636(.An(i_11_), .B(i_12_), .Y(mai_mai_n659_));
  NOi41      m637(.An(mai_mai_n102_), .B(mai_mai_n659_), .C(i_13_), .D(mai_mai_n76_), .Y(mai_mai_n660_));
  NA2        m638(.A(mai_mai_n660_), .B(mai_mai_n46_), .Y(mai_mai_n661_));
  NA3        m639(.A(mai_mai_n661_), .B(mai_mai_n658_), .C(mai_mai_n657_), .Y(mai_mai_n662_));
  OAI210     m640(.A0(mai_mai_n662_), .A1(mai_mai_n656_), .B0(mai_mai_n58_), .Y(mai_mai_n663_));
  NO2        m641(.A(i_2_), .B(i_12_), .Y(mai_mai_n664_));
  NA2        m642(.A(mai_mai_n347_), .B(mai_mai_n664_), .Y(mai_mai_n665_));
  NO3        m643(.A(i_9_), .B(mai_mai_n359_), .C(mai_mai_n554_), .Y(mai_mai_n666_));
  NA2        m644(.A(mai_mai_n666_), .B(mai_mai_n347_), .Y(mai_mai_n667_));
  NO2        m645(.A(mai_mai_n120_), .B(i_2_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n668_), .B(mai_mai_n583_), .Y(mai_mai_n669_));
  NA3        m647(.A(mai_mai_n669_), .B(mai_mai_n667_), .C(mai_mai_n665_), .Y(mai_mai_n670_));
  NA3        m648(.A(mai_mai_n670_), .B(mai_mai_n45_), .C(mai_mai_n213_), .Y(mai_mai_n671_));
  NA4        m649(.A(mai_mai_n671_), .B(mai_mai_n663_), .C(mai_mai_n653_), .D(mai_mai_n641_), .Y(mai_mai_n672_));
  OR4        m650(.A(mai_mai_n672_), .B(mai_mai_n631_), .C(mai_mai_n623_), .D(mai_mai_n571_), .Y(mai5));
  NA2        m651(.A(mai_mai_n611_), .B(mai_mai_n253_), .Y(mai_mai_n674_));
  AN2        m652(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n675_));
  NA3        m653(.A(mai_mai_n675_), .B(mai_mai_n664_), .C(mai_mai_n100_), .Y(mai_mai_n676_));
  NO2        m654(.A(mai_mai_n555_), .B(i_11_), .Y(mai_mai_n677_));
  NA2        m655(.A(mai_mai_n79_), .B(mai_mai_n677_), .Y(mai_mai_n678_));
  NA3        m656(.A(mai_mai_n678_), .B(mai_mai_n676_), .C(mai_mai_n674_), .Y(mai_mai_n679_));
  NO3        m657(.A(i_11_), .B(mai_mai_n224_), .C(i_13_), .Y(mai_mai_n680_));
  NO2        m658(.A(mai_mai_n116_), .B(mai_mai_n23_), .Y(mai_mai_n681_));
  NA2        m659(.A(i_12_), .B(i_8_), .Y(mai_mai_n682_));
  OAI210     m660(.A0(mai_mai_n46_), .A1(i_3_), .B0(mai_mai_n682_), .Y(mai_mai_n683_));
  INV        m661(.A(mai_mai_n419_), .Y(mai_mai_n684_));
  AOI220     m662(.A0(mai_mai_n299_), .A1(mai_mai_n537_), .B0(mai_mai_n683_), .B1(mai_mai_n681_), .Y(mai_mai_n685_));
  INV        m663(.A(mai_mai_n685_), .Y(mai_mai_n686_));
  NO2        m664(.A(mai_mai_n686_), .B(mai_mai_n679_), .Y(mai_mai_n687_));
  INV        m665(.A(mai_mai_n161_), .Y(mai_mai_n688_));
  INV        m666(.A(mai_mai_n233_), .Y(mai_mai_n689_));
  OAI210     m667(.A0(mai_mai_n629_), .A1(mai_mai_n421_), .B0(mai_mai_n102_), .Y(mai_mai_n690_));
  AOI210     m668(.A0(mai_mai_n690_), .A1(mai_mai_n689_), .B0(mai_mai_n688_), .Y(mai_mai_n691_));
  NO2        m669(.A(mai_mai_n428_), .B(mai_mai_n26_), .Y(mai_mai_n692_));
  NO2        m670(.A(mai_mai_n692_), .B(mai_mai_n396_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n693_), .B(i_2_), .Y(mai_mai_n694_));
  INV        m672(.A(mai_mai_n694_), .Y(mai_mai_n695_));
  AOI210     m673(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n393_), .Y(mai_mai_n696_));
  AOI210     m674(.A0(mai_mai_n696_), .A1(mai_mai_n695_), .B0(mai_mai_n691_), .Y(mai_mai_n697_));
  NO2        m675(.A(mai_mai_n179_), .B(mai_mai_n117_), .Y(mai_mai_n698_));
  OAI210     m676(.A0(mai_mai_n698_), .A1(mai_mai_n681_), .B0(i_2_), .Y(mai_mai_n699_));
  INV        m677(.A(mai_mai_n162_), .Y(mai_mai_n700_));
  NO3        m678(.A(mai_mai_n573_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n701_));
  AOI210     m679(.A0(mai_mai_n700_), .A1(mai_mai_n79_), .B0(mai_mai_n701_), .Y(mai_mai_n702_));
  AOI210     m680(.A0(mai_mai_n702_), .A1(mai_mai_n699_), .B0(mai_mai_n182_), .Y(mai_mai_n703_));
  OA210      m681(.A0(mai_mai_n574_), .A1(mai_mai_n118_), .B0(i_13_), .Y(mai_mai_n704_));
  INV        m682(.A(mai_mai_n142_), .Y(mai_mai_n705_));
  NO2        m683(.A(mai_mai_n705_), .B(mai_mai_n349_), .Y(mai_mai_n706_));
  NO2        m684(.A(mai_mai_n139_), .B(mai_mai_n483_), .Y(mai_mai_n707_));
  NA2        m685(.A(mai_mai_n707_), .B(mai_mai_n396_), .Y(mai_mai_n708_));
  NO2        m686(.A(mai_mai_n94_), .B(mai_mai_n44_), .Y(mai_mai_n709_));
  INV        m687(.A(mai_mai_n285_), .Y(mai_mai_n710_));
  NA4        m688(.A(mai_mai_n710_), .B(mai_mai_n289_), .C(mai_mai_n116_), .D(mai_mai_n42_), .Y(mai_mai_n711_));
  OAI210     m689(.A0(mai_mai_n711_), .A1(mai_mai_n709_), .B0(mai_mai_n708_), .Y(mai_mai_n712_));
  NO4        m690(.A(mai_mai_n712_), .B(mai_mai_n706_), .C(mai_mai_n704_), .D(mai_mai_n703_), .Y(mai_mai_n713_));
  NA2        m691(.A(mai_mai_n537_), .B(mai_mai_n28_), .Y(mai_mai_n714_));
  NA2        m692(.A(mai_mai_n680_), .B(mai_mai_n258_), .Y(mai_mai_n715_));
  NA2        m693(.A(mai_mai_n715_), .B(mai_mai_n714_), .Y(mai_mai_n716_));
  NO2        m694(.A(mai_mai_n57_), .B(i_12_), .Y(mai_mai_n717_));
  NO2        m695(.A(mai_mai_n717_), .B(mai_mai_n118_), .Y(mai_mai_n718_));
  NO2        m696(.A(mai_mai_n718_), .B(mai_mai_n552_), .Y(mai_mai_n719_));
  AOI220     m697(.A0(mai_mai_n719_), .A1(mai_mai_n36_), .B0(mai_mai_n716_), .B1(mai_mai_n46_), .Y(mai_mai_n720_));
  NA4        m698(.A(mai_mai_n720_), .B(mai_mai_n713_), .C(mai_mai_n697_), .D(mai_mai_n687_), .Y(mai6));
  NO3        m699(.A(i_9_), .B(mai_mai_n291_), .C(i_1_), .Y(mai_mai_n722_));
  NO2        m700(.A(mai_mai_n174_), .B(mai_mai_n130_), .Y(mai_mai_n723_));
  OAI210     m701(.A0(mai_mai_n723_), .A1(mai_mai_n722_), .B0(mai_mai_n668_), .Y(mai_mai_n724_));
  NA4        m702(.A(mai_mai_n365_), .B(mai_mai_n452_), .C(mai_mai_n63_), .D(mai_mai_n93_), .Y(mai_mai_n725_));
  INV        m703(.A(mai_mai_n725_), .Y(mai_mai_n726_));
  NO2        m704(.A(i_11_), .B(i_9_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n726_), .B(mai_mai_n311_), .Y(mai_mai_n728_));
  AO210      m706(.A0(mai_mai_n728_), .A1(mai_mai_n724_), .B0(i_12_), .Y(mai_mai_n729_));
  NA2        m707(.A(mai_mai_n350_), .B(mai_mai_n317_), .Y(mai_mai_n730_));
  NA2        m708(.A(mai_mai_n544_), .B(mai_mai_n58_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n625_), .B(mai_mai_n63_), .Y(mai_mai_n732_));
  BUFFER     m710(.A(mai_mai_n579_), .Y(mai_mai_n733_));
  NA4        m711(.A(mai_mai_n733_), .B(mai_mai_n732_), .C(mai_mai_n731_), .D(mai_mai_n730_), .Y(mai_mai_n734_));
  INV        m712(.A(mai_mai_n186_), .Y(mai_mai_n735_));
  AOI220     m713(.A0(mai_mai_n735_), .A1(mai_mai_n727_), .B0(mai_mai_n734_), .B1(mai_mai_n65_), .Y(mai_mai_n736_));
  INV        m714(.A(mai_mai_n310_), .Y(mai_mai_n737_));
  NA2        m715(.A(mai_mai_n67_), .B(mai_mai_n123_), .Y(mai_mai_n738_));
  INV        m716(.A(mai_mai_n116_), .Y(mai_mai_n739_));
  NA2        m717(.A(mai_mai_n739_), .B(mai_mai_n46_), .Y(mai_mai_n740_));
  AOI210     m718(.A0(mai_mai_n740_), .A1(mai_mai_n738_), .B0(mai_mai_n737_), .Y(mai_mai_n741_));
  NO2        m719(.A(mai_mai_n240_), .B(i_9_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n742_), .B(mai_mai_n717_), .Y(mai_mai_n743_));
  NO2        m721(.A(mai_mai_n743_), .B(mai_mai_n174_), .Y(mai_mai_n744_));
  NO2        m722(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n745_));
  NA3        m723(.A(mai_mai_n745_), .B(mai_mai_n448_), .C(mai_mai_n365_), .Y(mai_mai_n746_));
  OAI210     m724(.A0(mai_mai_n624_), .A1(mai_mai_n525_), .B0(mai_mai_n524_), .Y(mai_mai_n747_));
  NA2        m725(.A(mai_mai_n747_), .B(mai_mai_n746_), .Y(mai_mai_n748_));
  OR3        m726(.A(mai_mai_n748_), .B(mai_mai_n744_), .C(mai_mai_n741_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n632_), .B(i_2_), .Y(mai_mai_n750_));
  NA2        m728(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n751_));
  OAI210     m729(.A0(mai_mai_n751_), .A1(mai_mai_n385_), .B0(mai_mai_n341_), .Y(mai_mai_n752_));
  NA2        m730(.A(mai_mai_n752_), .B(mai_mai_n750_), .Y(mai_mai_n753_));
  AO210      m731(.A0(mai_mai_n340_), .A1(mai_mai_n331_), .B0(mai_mai_n373_), .Y(mai_mai_n754_));
  NA3        m732(.A(mai_mai_n754_), .B(mai_mai_n243_), .C(i_7_), .Y(mai_mai_n755_));
  OR2        m733(.A(mai_mai_n574_), .B(mai_mai_n421_), .Y(mai_mai_n756_));
  NA3        m734(.A(mai_mai_n756_), .B(mai_mai_n138_), .C(mai_mai_n61_), .Y(mai_mai_n757_));
  AO210      m735(.A0(mai_mai_n463_), .A1(mai_mai_n684_), .B0(mai_mai_n36_), .Y(mai_mai_n758_));
  NA4        m736(.A(mai_mai_n758_), .B(mai_mai_n757_), .C(mai_mai_n755_), .D(mai_mai_n753_), .Y(mai_mai_n759_));
  OAI210     m737(.A0(mai_mai_n588_), .A1(i_11_), .B0(mai_mai_n77_), .Y(mai_mai_n760_));
  NA2        m738(.A(mai_mai_n760_), .B(mai_mai_n524_), .Y(mai_mai_n761_));
  NA2        m739(.A(mai_mai_n373_), .B(mai_mai_n62_), .Y(mai_mai_n762_));
  NA3        m740(.A(mai_mai_n762_), .B(mai_mai_n761_), .C(mai_mai_n558_), .Y(mai_mai_n763_));
  AO210      m741(.A0(mai_mai_n483_), .A1(mai_mai_n46_), .B0(mai_mai_n78_), .Y(mai_mai_n764_));
  NA3        m742(.A(mai_mai_n764_), .B(mai_mai_n453_), .C(mai_mai_n207_), .Y(mai_mai_n765_));
  AOI210     m743(.A0(mai_mai_n421_), .A1(mai_mai_n419_), .B0(mai_mai_n523_), .Y(mai_mai_n766_));
  NA2        m744(.A(mai_mai_n103_), .B(mai_mai_n383_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n232_), .B(mai_mai_n46_), .Y(mai_mai_n768_));
  NA3        m746(.A(mai_mai_n767_), .B(mai_mai_n766_), .C(mai_mai_n765_), .Y(mai_mai_n769_));
  NO4        m747(.A(mai_mai_n769_), .B(mai_mai_n763_), .C(mai_mai_n759_), .D(mai_mai_n749_), .Y(mai_mai_n770_));
  NA4        m748(.A(mai_mai_n770_), .B(mai_mai_n736_), .C(mai_mai_n729_), .D(mai_mai_n355_), .Y(mai3));
  NA2        m749(.A(i_6_), .B(i_7_), .Y(mai_mai_n772_));
  NO2        m750(.A(mai_mai_n772_), .B(i_0_), .Y(mai_mai_n773_));
  NO2        m751(.A(i_11_), .B(mai_mai_n224_), .Y(mai_mai_n774_));
  OAI210     m752(.A0(mai_mai_n773_), .A1(mai_mai_n273_), .B0(mai_mai_n774_), .Y(mai_mai_n775_));
  INV        m753(.A(mai_mai_n775_), .Y(mai_mai_n776_));
  NO3        m754(.A(mai_mai_n424_), .B(mai_mai_n82_), .C(mai_mai_n44_), .Y(mai_mai_n777_));
  OA210      m755(.A0(mai_mai_n777_), .A1(mai_mai_n776_), .B0(mai_mai_n164_), .Y(mai_mai_n778_));
  NA2        m756(.A(mai_mai_n386_), .B(mai_mai_n45_), .Y(mai_mai_n779_));
  NO4        m757(.A(mai_mai_n351_), .B(mai_mai_n358_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n780_));
  INV        m758(.A(mai_mai_n780_), .Y(mai_mai_n781_));
  NA2        m759(.A(mai_mai_n645_), .B(mai_mai_n617_), .Y(mai_mai_n782_));
  NA2        m760(.A(i_0_), .B(i_5_), .Y(mai_mai_n783_));
  OAI220     m761(.A0(mai_mai_n783_), .A1(mai_mai_n782_), .B0(mai_mai_n781_), .B1(mai_mai_n58_), .Y(mai_mai_n784_));
  NO2        m762(.A(mai_mai_n165_), .B(mai_mai_n139_), .Y(mai_mai_n785_));
  NA2        m763(.A(mai_mai_n785_), .B(mai_mai_n232_), .Y(mai_mai_n786_));
  NO2        m764(.A(mai_mai_n786_), .B(mai_mai_n965_), .Y(mai_mai_n787_));
  NO3        m765(.A(mai_mai_n787_), .B(mai_mai_n784_), .C(mai_mai_n778_), .Y(mai_mai_n788_));
  NA2        m766(.A(mai_mai_n174_), .B(mai_mai_n24_), .Y(mai_mai_n789_));
  NO2        m767(.A(mai_mai_n615_), .B(mai_mai_n550_), .Y(mai_mai_n790_));
  NO2        m768(.A(mai_mai_n790_), .B(mai_mai_n789_), .Y(mai_mai_n791_));
  NA2        m769(.A(mai_mai_n296_), .B(mai_mai_n121_), .Y(mai_mai_n792_));
  OAI220     m770(.A0(mai_mai_n152_), .A1(mai_mai_n768_), .B0(mai_mai_n792_), .B1(mai_mai_n376_), .Y(mai_mai_n793_));
  NO2        m771(.A(mai_mai_n793_), .B(mai_mai_n791_), .Y(mai_mai_n794_));
  NO2        m772(.A(mai_mai_n365_), .B(mai_mai_n277_), .Y(mai_mai_n795_));
  NA2        m773(.A(mai_mai_n795_), .B(mai_mai_n648_), .Y(mai_mai_n796_));
  INV        m774(.A(mai_mai_n448_), .Y(mai_mai_n797_));
  AN2        m775(.A(mai_mai_n88_), .B(mai_mai_n231_), .Y(mai_mai_n798_));
  NA2        m776(.A(mai_mai_n680_), .B(mai_mai_n311_), .Y(mai_mai_n799_));
  INV        m777(.A(mai_mai_n55_), .Y(mai_mai_n800_));
  OAI220     m778(.A0(mai_mai_n800_), .A1(mai_mai_n799_), .B0(mai_mai_n606_), .B1(mai_mai_n499_), .Y(mai_mai_n801_));
  NO2        m779(.A(mai_mai_n242_), .B(mai_mai_n143_), .Y(mai_mai_n802_));
  NA2        m780(.A(i_0_), .B(i_10_), .Y(mai_mai_n803_));
  AN2        m781(.A(mai_mai_n802_), .B(i_6_), .Y(mai_mai_n804_));
  NA2        m782(.A(mai_mai_n174_), .B(mai_mai_n74_), .Y(mai_mai_n805_));
  NA2        m783(.A(mai_mai_n528_), .B(i_4_), .Y(mai_mai_n806_));
  NA2        m784(.A(mai_mai_n177_), .B(mai_mai_n192_), .Y(mai_mai_n807_));
  OAI220     m785(.A0(mai_mai_n807_), .A1(mai_mai_n799_), .B0(mai_mai_n806_), .B1(mai_mai_n805_), .Y(mai_mai_n808_));
  NO4        m786(.A(mai_mai_n808_), .B(mai_mai_n804_), .C(mai_mai_n801_), .D(mai_mai_n798_), .Y(mai_mai_n809_));
  NA3        m787(.A(mai_mai_n809_), .B(mai_mai_n796_), .C(mai_mai_n794_), .Y(mai_mai_n810_));
  NA2        m788(.A(i_11_), .B(i_9_), .Y(mai_mai_n811_));
  NO2        m789(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n812_));
  NA2        m790(.A(mai_mai_n370_), .B(mai_mai_n169_), .Y(mai_mai_n813_));
  NA2        m791(.A(mai_mai_n813_), .B(mai_mai_n150_), .Y(mai_mai_n814_));
  NO2        m792(.A(mai_mai_n811_), .B(mai_mai_n65_), .Y(mai_mai_n815_));
  NO2        m793(.A(mai_mai_n165_), .B(i_0_), .Y(mai_mai_n816_));
  INV        m794(.A(mai_mai_n816_), .Y(mai_mai_n817_));
  NA2        m795(.A(mai_mai_n448_), .B(mai_mai_n219_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n818_), .B(mai_mai_n817_), .Y(mai_mai_n819_));
  NO2        m797(.A(mai_mai_n819_), .B(mai_mai_n814_), .Y(mai_mai_n820_));
  NA2        m798(.A(mai_mai_n605_), .B(mai_mai_n113_), .Y(mai_mai_n821_));
  NO2        m799(.A(i_6_), .B(mai_mai_n821_), .Y(mai_mai_n822_));
  AOI210     m800(.A0(mai_mai_n420_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n823_));
  NA2        m801(.A(mai_mai_n161_), .B(mai_mai_n95_), .Y(mai_mai_n824_));
  NOi32      m802(.An(mai_mai_n823_), .Bn(mai_mai_n177_), .C(mai_mai_n824_), .Y(mai_mai_n825_));
  NA2        m803(.A(mai_mai_n559_), .B(mai_mai_n311_), .Y(mai_mai_n826_));
  NO2        m804(.A(mai_mai_n826_), .B(mai_mai_n779_), .Y(mai_mai_n827_));
  NO3        m805(.A(mai_mai_n827_), .B(mai_mai_n825_), .C(mai_mai_n822_), .Y(mai_mai_n828_));
  NOi21      m806(.An(i_7_), .B(i_5_), .Y(mai_mai_n829_));
  NOi31      m807(.An(mai_mai_n829_), .B(i_0_), .C(mai_mai_n659_), .Y(mai_mai_n830_));
  NO3        m808(.A(mai_mai_n378_), .B(mai_mai_n343_), .C(mai_mai_n339_), .Y(mai_mai_n831_));
  NO2        m809(.A(mai_mai_n244_), .B(mai_mai_n300_), .Y(mai_mai_n832_));
  INV        m810(.A(mai_mai_n659_), .Y(mai_mai_n833_));
  AOI210     m811(.A0(mai_mai_n833_), .A1(mai_mai_n832_), .B0(mai_mai_n831_), .Y(mai_mai_n834_));
  NA3        m812(.A(mai_mai_n834_), .B(mai_mai_n828_), .C(mai_mai_n820_), .Y(mai_mai_n835_));
  NO2        m813(.A(mai_mai_n789_), .B(mai_mai_n227_), .Y(mai_mai_n836_));
  AN2        m814(.A(mai_mai_n315_), .B(mai_mai_n311_), .Y(mai_mai_n837_));
  AN2        m815(.A(mai_mai_n837_), .B(mai_mai_n785_), .Y(mai_mai_n838_));
  OAI210     m816(.A0(mai_mai_n838_), .A1(mai_mai_n836_), .B0(i_10_), .Y(mai_mai_n839_));
  NA3        m817(.A(mai_mai_n447_), .B(mai_mai_n386_), .C(mai_mai_n45_), .Y(mai_mai_n840_));
  OAI210     m818(.A0(mai_mai_n152_), .A1(mai_mai_n797_), .B0(mai_mai_n840_), .Y(mai_mai_n841_));
  NO2        m819(.A(mai_mai_n243_), .B(mai_mai_n46_), .Y(mai_mai_n842_));
  NA2        m820(.A(mai_mai_n815_), .B(mai_mai_n289_), .Y(mai_mai_n843_));
  OAI210     m821(.A0(mai_mai_n842_), .A1(mai_mai_n176_), .B0(mai_mai_n843_), .Y(mai_mai_n844_));
  AOI220     m822(.A0(mai_mai_n844_), .A1(mai_mai_n448_), .B0(mai_mai_n841_), .B1(mai_mai_n65_), .Y(mai_mai_n845_));
  NA3        m823(.A(mai_mai_n751_), .B(mai_mai_n357_), .C(mai_mai_n588_), .Y(mai_mai_n846_));
  NA2        m824(.A(mai_mai_n85_), .B(mai_mai_n44_), .Y(mai_mai_n847_));
  NO2        m825(.A(mai_mai_n67_), .B(mai_mai_n682_), .Y(mai_mai_n848_));
  AOI220     m826(.A0(mai_mai_n848_), .A1(mai_mai_n847_), .B0(mai_mai_n164_), .B1(mai_mai_n550_), .Y(mai_mai_n849_));
  AOI210     m827(.A0(mai_mai_n849_), .A1(mai_mai_n846_), .B0(mai_mai_n47_), .Y(mai_mai_n850_));
  NO3        m828(.A(i_5_), .B(mai_mai_n338_), .C(mai_mai_n24_), .Y(mai_mai_n851_));
  AOI210     m829(.A0(mai_mai_n638_), .A1(mai_mai_n509_), .B0(mai_mai_n851_), .Y(mai_mai_n852_));
  NAi21      m830(.An(i_9_), .B(i_5_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n553_), .B(mai_mai_n97_), .Y(mai_mai_n854_));
  NA2        m832(.A(mai_mai_n854_), .B(i_0_), .Y(mai_mai_n855_));
  OAI220     m833(.A0(mai_mai_n855_), .A1(mai_mai_n76_), .B0(mai_mai_n852_), .B1(mai_mai_n162_), .Y(mai_mai_n856_));
  NO3        m834(.A(mai_mai_n856_), .B(mai_mai_n850_), .C(mai_mai_n394_), .Y(mai_mai_n857_));
  NA3        m835(.A(mai_mai_n857_), .B(mai_mai_n845_), .C(mai_mai_n839_), .Y(mai_mai_n858_));
  NO3        m836(.A(mai_mai_n858_), .B(mai_mai_n835_), .C(mai_mai_n810_), .Y(mai_mai_n859_));
  NO2        m837(.A(i_0_), .B(mai_mai_n659_), .Y(mai_mai_n860_));
  NO3        m838(.A(mai_mai_n97_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n861_));
  AO220      m839(.A0(mai_mai_n861_), .A1(mai_mai_n44_), .B0(mai_mai_n860_), .B1(mai_mai_n164_), .Y(mai_mai_n862_));
  NO2        m840(.A(mai_mai_n731_), .B(mai_mai_n824_), .Y(mai_mai_n863_));
  AOI210     m841(.A0(mai_mai_n862_), .A1(mai_mai_n329_), .B0(mai_mai_n863_), .Y(mai_mai_n864_));
  NA3        m842(.A(mai_mai_n137_), .B(mai_mai_n617_), .C(mai_mai_n65_), .Y(mai_mai_n865_));
  NO2        m843(.A(mai_mai_n747_), .B(mai_mai_n378_), .Y(mai_mai_n866_));
  NA3        m844(.A(mai_mai_n773_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n867_));
  NA2        m845(.A(mai_mai_n774_), .B(i_9_), .Y(mai_mai_n868_));
  AOI210     m846(.A0(mai_mai_n867_), .A1(mai_mai_n466_), .B0(mai_mai_n868_), .Y(mai_mai_n869_));
  NO2        m847(.A(mai_mai_n869_), .B(mai_mai_n866_), .Y(mai_mai_n870_));
  NA3        m848(.A(mai_mai_n870_), .B(mai_mai_n865_), .C(mai_mai_n864_), .Y(mai_mai_n871_));
  NA2        m849(.A(mai_mai_n837_), .B(mai_mai_n349_), .Y(mai_mai_n872_));
  AOI210     m850(.A0(mai_mai_n284_), .A1(mai_mai_n152_), .B0(mai_mai_n872_), .Y(mai_mai_n873_));
  NA3        m851(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n874_));
  NA2        m852(.A(mai_mai_n812_), .B(mai_mai_n457_), .Y(mai_mai_n875_));
  AOI210     m853(.A0(mai_mai_n874_), .A1(mai_mai_n152_), .B0(mai_mai_n875_), .Y(mai_mai_n876_));
  NO2        m854(.A(mai_mai_n876_), .B(mai_mai_n873_), .Y(mai_mai_n877_));
  NO2        m855(.A(mai_mai_n803_), .B(mai_mai_n179_), .Y(mai_mai_n878_));
  AOI220     m856(.A0(mai_mai_n878_), .A1(i_11_), .B0(mai_mai_n529_), .B1(mai_mai_n67_), .Y(mai_mai_n879_));
  NO3        m857(.A(mai_mai_n199_), .B(mai_mai_n358_), .C(i_0_), .Y(mai_mai_n880_));
  OAI210     m858(.A0(mai_mai_n880_), .A1(mai_mai_n68_), .B0(i_13_), .Y(mai_mai_n881_));
  INV        m859(.A(mai_mai_n207_), .Y(mai_mai_n882_));
  NO2        m860(.A(mai_mai_n593_), .B(mai_mai_n568_), .Y(mai_mai_n883_));
  NA2        m861(.A(mai_mai_n883_), .B(mai_mai_n882_), .Y(mai_mai_n884_));
  NA4        m862(.A(mai_mai_n884_), .B(mai_mai_n881_), .C(mai_mai_n879_), .D(mai_mai_n877_), .Y(mai_mai_n885_));
  NA2        m863(.A(mai_mai_n829_), .B(mai_mai_n457_), .Y(mai_mai_n886_));
  INV        m864(.A(mai_mai_n166_), .Y(mai_mai_n887_));
  OR2        m865(.A(mai_mai_n887_), .B(mai_mai_n886_), .Y(mai_mai_n888_));
  AOI210     m866(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n165_), .Y(mai_mai_n889_));
  NA3        m867(.A(mai_mai_n565_), .B(mai_mai_n174_), .C(mai_mai_n74_), .Y(mai_mai_n890_));
  NA2        m868(.A(mai_mai_n890_), .B(mai_mai_n507_), .Y(mai_mai_n891_));
  NO3        m869(.A(mai_mai_n779_), .B(mai_mai_n53_), .C(mai_mai_n48_), .Y(mai_mai_n892_));
  INV        m870(.A(mai_mai_n462_), .Y(mai_mai_n893_));
  NO3        m871(.A(mai_mai_n893_), .B(mai_mai_n892_), .C(mai_mai_n891_), .Y(mai_mai_n894_));
  NA3        m872(.A(mai_mai_n812_), .B(mai_mai_n273_), .C(mai_mai_n218_), .Y(mai_mai_n895_));
  INV        m873(.A(mai_mai_n895_), .Y(mai_mai_n896_));
  NA3        m874(.A(mai_mai_n365_), .B(mai_mai_n316_), .C(mai_mai_n210_), .Y(mai_mai_n897_));
  INV        m875(.A(mai_mai_n897_), .Y(mai_mai_n898_));
  NO3        m876(.A(mai_mai_n811_), .B(mai_mai_n207_), .C(mai_mai_n179_), .Y(mai_mai_n899_));
  NO3        m877(.A(mai_mai_n899_), .B(mai_mai_n898_), .C(mai_mai_n896_), .Y(mai_mai_n900_));
  NA3        m878(.A(mai_mai_n900_), .B(mai_mai_n894_), .C(mai_mai_n888_), .Y(mai_mai_n901_));
  INV        m879(.A(mai_mai_n567_), .Y(mai_mai_n902_));
  NO3        m880(.A(mai_mai_n902_), .B(mai_mai_n519_), .C(mai_mai_n327_), .Y(mai_mai_n903_));
  INV        m881(.A(mai_mai_n903_), .Y(mai_mai_n904_));
  NA3        m882(.A(mai_mai_n289_), .B(i_5_), .C(mai_mai_n182_), .Y(mai_mai_n905_));
  NA2        m883(.A(mai_mai_n905_), .B(mai_mai_n230_), .Y(mai_mai_n906_));
  NO4        m884(.A(mai_mai_n227_), .B(mai_mai_n199_), .C(i_0_), .D(i_12_), .Y(mai_mai_n907_));
  AOI220     m885(.A0(mai_mai_n907_), .A1(mai_mai_n906_), .B0(mai_mai_n726_), .B1(mai_mai_n166_), .Y(mai_mai_n908_));
  AN2        m886(.A(mai_mai_n803_), .B(mai_mai_n143_), .Y(mai_mai_n909_));
  NO4        m887(.A(mai_mai_n909_), .B(i_12_), .C(mai_mai_n595_), .D(mai_mai_n123_), .Y(mai_mai_n910_));
  NA2        m888(.A(mai_mai_n910_), .B(mai_mai_n207_), .Y(mai_mai_n911_));
  NA3        m889(.A(mai_mai_n90_), .B(mai_mai_n533_), .C(i_11_), .Y(mai_mai_n912_));
  NO2        m890(.A(mai_mai_n912_), .B(mai_mai_n145_), .Y(mai_mai_n913_));
  NA2        m891(.A(mai_mai_n829_), .B(mai_mai_n445_), .Y(mai_mai_n914_));
  OAI220     m892(.A0(i_7_), .A1(mai_mai_n905_), .B0(mai_mai_n914_), .B1(mai_mai_n618_), .Y(mai_mai_n915_));
  AOI210     m893(.A0(mai_mai_n915_), .A1(mai_mai_n816_), .B0(mai_mai_n913_), .Y(mai_mai_n916_));
  NA4        m894(.A(mai_mai_n916_), .B(mai_mai_n911_), .C(mai_mai_n908_), .D(mai_mai_n904_), .Y(mai_mai_n917_));
  NO4        m895(.A(mai_mai_n917_), .B(mai_mai_n901_), .C(mai_mai_n885_), .D(mai_mai_n871_), .Y(mai_mai_n918_));
  OAI210     m896(.A0(mai_mai_n750_), .A1(mai_mai_n745_), .B0(mai_mai_n37_), .Y(mai_mai_n919_));
  NA3        m897(.A(mai_mai_n823_), .B(mai_mai_n347_), .C(i_5_), .Y(mai_mai_n920_));
  NA3        m898(.A(mai_mai_n920_), .B(mai_mai_n919_), .C(mai_mai_n563_), .Y(mai_mai_n921_));
  NA2        m899(.A(mai_mai_n921_), .B(mai_mai_n196_), .Y(mai_mai_n922_));
  NA2        m900(.A(mai_mai_n175_), .B(mai_mai_n177_), .Y(mai_mai_n923_));
  AO210      m901(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n923_), .Y(mai_mai_n924_));
  OAI210     m902(.A0(mai_mai_n567_), .A1(mai_mai_n565_), .B0(mai_mai_n299_), .Y(mai_mai_n925_));
  NAi31      m903(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n926_));
  NO2        m904(.A(mai_mai_n62_), .B(mai_mai_n926_), .Y(mai_mai_n927_));
  INV        m905(.A(mai_mai_n927_), .Y(mai_mai_n928_));
  NA3        m906(.A(mai_mai_n928_), .B(mai_mai_n925_), .C(mai_mai_n924_), .Y(mai_mai_n929_));
  NO2        m907(.A(mai_mai_n436_), .B(mai_mai_n250_), .Y(mai_mai_n930_));
  NO4        m908(.A(mai_mai_n221_), .B(mai_mai_n136_), .C(mai_mai_n621_), .D(mai_mai_n37_), .Y(mai_mai_n931_));
  NO2        m909(.A(mai_mai_n931_), .B(mai_mai_n930_), .Y(mai_mai_n932_));
  OAI210     m910(.A0(mai_mai_n912_), .A1(mai_mai_n139_), .B0(mai_mai_n932_), .Y(mai_mai_n933_));
  AOI210     m911(.A0(mai_mai_n929_), .A1(mai_mai_n48_), .B0(mai_mai_n933_), .Y(mai_mai_n934_));
  AOI210     m912(.A0(mai_mai_n934_), .A1(mai_mai_n922_), .B0(mai_mai_n65_), .Y(mai_mai_n935_));
  NO2        m913(.A(mai_mai_n526_), .B(mai_mai_n354_), .Y(mai_mai_n936_));
  NO2        m914(.A(mai_mai_n936_), .B(mai_mai_n688_), .Y(mai_mai_n937_));
  INV        m915(.A(mai_mai_n100_), .Y(mai_mai_n938_));
  NA2        m916(.A(mai_mai_n938_), .B(mai_mai_n68_), .Y(mai_mai_n939_));
  AOI210     m917(.A0(mai_mai_n889_), .A1(mai_mai_n812_), .B0(mai_mai_n830_), .Y(mai_mai_n940_));
  AOI210     m918(.A0(mai_mai_n940_), .A1(mai_mai_n939_), .B0(mai_mai_n621_), .Y(mai_mai_n941_));
  INV        m919(.A(mai_mai_n244_), .Y(mai_mai_n942_));
  NA2        m920(.A(mai_mai_n942_), .B(mai_mai_n68_), .Y(mai_mai_n943_));
  NO2        m921(.A(mai_mai_n943_), .B(mai_mai_n224_), .Y(mai_mai_n944_));
  NA3        m922(.A(mai_mai_n88_), .B(mai_mai_n291_), .C(mai_mai_n31_), .Y(mai_mai_n945_));
  INV        m923(.A(mai_mai_n945_), .Y(mai_mai_n946_));
  NO3        m924(.A(mai_mai_n946_), .B(mai_mai_n944_), .C(mai_mai_n941_), .Y(mai_mai_n947_));
  OAI210     m925(.A0(mai_mai_n252_), .A1(mai_mai_n148_), .B0(mai_mai_n79_), .Y(mai_mai_n948_));
  NA3        m926(.A(mai_mai_n692_), .B(mai_mai_n273_), .C(mai_mai_n72_), .Y(mai_mai_n949_));
  AOI210     m927(.A0(mai_mai_n949_), .A1(mai_mai_n948_), .B0(i_11_), .Y(mai_mai_n950_));
  INV        m928(.A(mai_mai_n196_), .Y(mai_mai_n951_));
  NA2        m929(.A(mai_mai_n154_), .B(i_5_), .Y(mai_mai_n952_));
  NO2        m930(.A(mai_mai_n951_), .B(mai_mai_n952_), .Y(mai_mai_n953_));
  NO3        m931(.A(mai_mai_n853_), .B(i_11_), .C(mai_mai_n241_), .Y(mai_mai_n954_));
  NO2        m932(.A(mai_mai_n954_), .B(mai_mai_n523_), .Y(mai_mai_n955_));
  INV        m933(.A(mai_mai_n344_), .Y(mai_mai_n956_));
  AOI210     m934(.A0(mai_mai_n956_), .A1(mai_mai_n955_), .B0(mai_mai_n41_), .Y(mai_mai_n957_));
  NO3        m935(.A(mai_mai_n957_), .B(mai_mai_n953_), .C(mai_mai_n950_), .Y(mai_mai_n958_));
  OAI210     m936(.A0(mai_mai_n947_), .A1(i_4_), .B0(mai_mai_n958_), .Y(mai_mai_n959_));
  NO3        m937(.A(mai_mai_n959_), .B(mai_mai_n937_), .C(mai_mai_n935_), .Y(mai_mai_n960_));
  NA4        m938(.A(mai_mai_n960_), .B(mai_mai_n918_), .C(mai_mai_n859_), .D(mai_mai_n788_), .Y(mai4));
  INV        m939(.A(i_2_), .Y(mai_mai_n964_));
  INV        m940(.A(i_5_), .Y(mai_mai_n965_));
  INV        m941(.A(i_0_), .Y(mai_mai_n966_));
  INV        m942(.A(mai_mai_n187_), .Y(mai_mai_n967_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  OAI210     u0028(.A0(men_men_n50_), .A1(i_3_), .B0(men_men_n48_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(men_men_n65_), .B(men_men_n61_), .Y(men_men_n66_));
  NA2        u0044(.A(men_men_n50_), .B(i_2_), .Y(men_men_n67_));
  NA2        u0045(.A(i_1_), .B(i_6_), .Y(men_men_n68_));
  NO2        u0046(.A(men_men_n68_), .B(men_men_n25_), .Y(men_men_n69_));
  INV        u0047(.A(i_0_), .Y(men_men_n70_));
  NAi21      u0048(.An(i_5_), .B(i_10_), .Y(men_men_n71_));
  NA2        u0049(.A(i_5_), .B(i_9_), .Y(men_men_n72_));
  AOI210     u0050(.A0(men_men_n72_), .A1(men_men_n71_), .B0(men_men_n70_), .Y(men_men_n73_));
  NO2        u0051(.A(men_men_n73_), .B(men_men_n69_), .Y(men_men_n74_));
  INV        u0052(.A(men_men_n74_), .Y(men_men_n75_));
  OAI210     u0053(.A0(men_men_n75_), .A1(men_men_n66_), .B0(i_0_), .Y(men_men_n76_));
  NA2        u0054(.A(i_12_), .B(i_5_), .Y(men_men_n77_));
  NA2        u0055(.A(i_2_), .B(i_8_), .Y(men_men_n78_));
  NO2        u0056(.A(men_men_n78_), .B(men_men_n58_), .Y(men_men_n79_));
  NO2        u0057(.A(i_3_), .B(i_9_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_7_), .Y(men_men_n81_));
  INV        u0059(.A(i_6_), .Y(men_men_n82_));
  OR4        u0060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n83_));
  INV        u0061(.A(men_men_n83_), .Y(men_men_n84_));
  NO2        u0062(.A(i_2_), .B(i_7_), .Y(men_men_n85_));
  INV        u0063(.A(men_men_n79_), .Y(men_men_n86_));
  NAi21      u0064(.An(i_6_), .B(i_10_), .Y(men_men_n87_));
  NA2        u0065(.A(i_6_), .B(i_9_), .Y(men_men_n88_));
  AOI210     u0066(.A0(men_men_n88_), .A1(men_men_n87_), .B0(men_men_n63_), .Y(men_men_n89_));
  NA2        u0067(.A(i_2_), .B(i_6_), .Y(men_men_n90_));
  NO3        u0068(.A(men_men_n90_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n91_));
  NO2        u0069(.A(men_men_n91_), .B(men_men_n89_), .Y(men_men_n92_));
  AOI210     u0070(.A0(men_men_n92_), .A1(men_men_n86_), .B0(men_men_n77_), .Y(men_men_n93_));
  AN3        u0071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n94_));
  NAi21      u0072(.An(i_6_), .B(i_11_), .Y(men_men_n95_));
  NO2        u0073(.A(i_5_), .B(i_8_), .Y(men_men_n96_));
  NOi21      u0074(.An(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  AOI220     u0075(.A0(men_men_n97_), .A1(men_men_n62_), .B0(men_men_n94_), .B1(men_men_n32_), .Y(men_men_n98_));
  INV        u0076(.A(i_7_), .Y(men_men_n99_));
  NA2        u0077(.A(men_men_n46_), .B(men_men_n99_), .Y(men_men_n100_));
  NO2        u0078(.A(i_0_), .B(i_5_), .Y(men_men_n101_));
  NO2        u0079(.A(men_men_n101_), .B(men_men_n82_), .Y(men_men_n102_));
  NA2        u0080(.A(i_12_), .B(i_3_), .Y(men_men_n103_));
  INV        u0081(.A(men_men_n103_), .Y(men_men_n104_));
  NA3        u0082(.A(men_men_n104_), .B(men_men_n102_), .C(men_men_n100_), .Y(men_men_n105_));
  NAi21      u0083(.An(i_7_), .B(i_11_), .Y(men_men_n106_));
  NO3        u0084(.A(men_men_n106_), .B(men_men_n87_), .C(men_men_n53_), .Y(men_men_n107_));
  AN2        u0085(.A(i_2_), .B(i_10_), .Y(men_men_n108_));
  NO2        u0086(.A(men_men_n108_), .B(i_7_), .Y(men_men_n109_));
  OR2        u0087(.A(men_men_n77_), .B(men_men_n58_), .Y(men_men_n110_));
  NO2        u0088(.A(i_8_), .B(men_men_n99_), .Y(men_men_n111_));
  NO3        u0089(.A(men_men_n111_), .B(men_men_n110_), .C(men_men_n109_), .Y(men_men_n112_));
  NA2        u0090(.A(i_12_), .B(i_7_), .Y(men_men_n113_));
  NO2        u0091(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n114_));
  NA2        u0092(.A(men_men_n114_), .B(i_0_), .Y(men_men_n115_));
  NA2        u0093(.A(i_11_), .B(i_12_), .Y(men_men_n116_));
  OAI210     u0094(.A0(men_men_n115_), .A1(men_men_n113_), .B0(men_men_n116_), .Y(men_men_n117_));
  NO2        u0095(.A(men_men_n117_), .B(men_men_n112_), .Y(men_men_n118_));
  NAi41      u0096(.An(men_men_n107_), .B(men_men_n118_), .C(men_men_n105_), .D(men_men_n98_), .Y(men_men_n119_));
  NOi21      u0097(.An(i_1_), .B(i_5_), .Y(men_men_n120_));
  NA2        u0098(.A(men_men_n120_), .B(i_11_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n99_), .B(men_men_n37_), .Y(men_men_n122_));
  NA2        u0100(.A(i_7_), .B(men_men_n25_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n123_), .B(men_men_n122_), .Y(men_men_n124_));
  NO2        u0102(.A(men_men_n124_), .B(men_men_n46_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n88_), .B(men_men_n87_), .Y(men_men_n126_));
  NAi21      u0104(.An(i_3_), .B(i_8_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n127_), .B(men_men_n62_), .Y(men_men_n128_));
  NOi21      u0106(.An(men_men_n128_), .B(men_men_n126_), .Y(men_men_n129_));
  NO2        u0107(.A(i_1_), .B(men_men_n82_), .Y(men_men_n130_));
  NO2        u0108(.A(i_6_), .B(i_5_), .Y(men_men_n131_));
  NA2        u0109(.A(men_men_n131_), .B(i_3_), .Y(men_men_n132_));
  AO210      u0110(.A0(men_men_n132_), .A1(men_men_n47_), .B0(men_men_n130_), .Y(men_men_n133_));
  OAI220     u0111(.A0(men_men_n133_), .A1(men_men_n106_), .B0(men_men_n129_), .B1(men_men_n121_), .Y(men_men_n134_));
  NO3        u0112(.A(men_men_n134_), .B(men_men_n119_), .C(men_men_n93_), .Y(men_men_n135_));
  NA3        u0113(.A(men_men_n135_), .B(men_men_n76_), .C(men_men_n56_), .Y(men2));
  NO2        u0114(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n137_));
  NA2        u0115(.A(i_6_), .B(men_men_n25_), .Y(men_men_n138_));
  NA2        u0116(.A(men_men_n138_), .B(men_men_n137_), .Y(men_men_n139_));
  NA4        u0117(.A(men_men_n139_), .B(men_men_n74_), .C(men_men_n67_), .D(men_men_n30_), .Y(men0));
  AN2        u0118(.A(i_8_), .B(i_7_), .Y(men_men_n141_));
  NA2        u0119(.A(men_men_n141_), .B(i_6_), .Y(men_men_n142_));
  NO2        u0120(.A(i_12_), .B(i_13_), .Y(men_men_n143_));
  NAi21      u0121(.An(i_5_), .B(i_11_), .Y(men_men_n144_));
  NOi21      u0122(.An(men_men_n143_), .B(men_men_n144_), .Y(men_men_n145_));
  NO2        u0123(.A(i_0_), .B(i_1_), .Y(men_men_n146_));
  NA2        u0124(.A(i_2_), .B(i_3_), .Y(men_men_n147_));
  NO2        u0125(.A(men_men_n147_), .B(i_4_), .Y(men_men_n148_));
  NA3        u0126(.A(men_men_n148_), .B(men_men_n146_), .C(men_men_n145_), .Y(men_men_n149_));
  OR2        u0127(.A(men_men_n149_), .B(men_men_n25_), .Y(men_men_n150_));
  AN2        u0128(.A(men_men_n143_), .B(men_men_n80_), .Y(men_men_n151_));
  NO2        u0129(.A(men_men_n151_), .B(men_men_n27_), .Y(men_men_n152_));
  NA2        u0130(.A(i_1_), .B(i_5_), .Y(men_men_n153_));
  NO2        u0131(.A(men_men_n70_), .B(men_men_n46_), .Y(men_men_n154_));
  NA2        u0132(.A(men_men_n154_), .B(men_men_n36_), .Y(men_men_n155_));
  NO3        u0133(.A(men_men_n155_), .B(men_men_n153_), .C(men_men_n152_), .Y(men_men_n156_));
  OR2        u0134(.A(i_0_), .B(i_1_), .Y(men_men_n157_));
  NO3        u0135(.A(men_men_n157_), .B(men_men_n77_), .C(i_13_), .Y(men_men_n158_));
  NAi32      u0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n159_));
  NAi21      u0137(.An(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  NOi21      u0138(.An(i_4_), .B(i_10_), .Y(men_men_n161_));
  NA2        u0139(.A(men_men_n161_), .B(men_men_n39_), .Y(men_men_n162_));
  NO2        u0140(.A(i_3_), .B(i_5_), .Y(men_men_n163_));
  NO3        u0141(.A(men_men_n70_), .B(i_2_), .C(i_1_), .Y(men_men_n164_));
  NA2        u0142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OAI210     u0143(.A0(men_men_n165_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n166_));
  NO2        u0144(.A(men_men_n166_), .B(men_men_n156_), .Y(men_men_n167_));
  AOI210     u0145(.A0(men_men_n167_), .A1(men_men_n150_), .B0(men_men_n142_), .Y(men_men_n168_));
  NA3        u0146(.A(men_men_n70_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n169_));
  NOi21      u0147(.An(i_4_), .B(i_9_), .Y(men_men_n170_));
  NOi21      u0148(.An(i_11_), .B(i_13_), .Y(men_men_n171_));
  NA2        u0149(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  NO2        u0150(.A(i_4_), .B(i_5_), .Y(men_men_n173_));
  NAi21      u0151(.An(i_12_), .B(i_11_), .Y(men_men_n174_));
  NO2        u0152(.A(men_men_n174_), .B(i_13_), .Y(men_men_n175_));
  NA3        u0153(.A(men_men_n175_), .B(men_men_n173_), .C(men_men_n80_), .Y(men_men_n176_));
  AOI210     u0154(.A0(men_men_n176_), .A1(men_men_n172_), .B0(men_men_n169_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n70_), .B(men_men_n63_), .Y(men_men_n178_));
  NA2        u0156(.A(men_men_n36_), .B(i_5_), .Y(men_men_n179_));
  NAi31      u0157(.An(men_men_n179_), .B(men_men_n151_), .C(i_11_), .Y(men_men_n180_));
  NA2        u0158(.A(i_3_), .B(i_5_), .Y(men_men_n181_));
  OR2        u0159(.A(men_men_n181_), .B(men_men_n172_), .Y(men_men_n182_));
  AOI210     u0160(.A0(men_men_n182_), .A1(men_men_n180_), .B0(i_2_), .Y(men_men_n183_));
  NO2        u0161(.A(men_men_n70_), .B(i_5_), .Y(men_men_n184_));
  NO2        u0162(.A(i_13_), .B(i_10_), .Y(men_men_n185_));
  NA3        u0163(.A(men_men_n185_), .B(men_men_n184_), .C(men_men_n44_), .Y(men_men_n186_));
  NO2        u0164(.A(i_2_), .B(i_1_), .Y(men_men_n187_));
  NA2        u0165(.A(men_men_n187_), .B(i_3_), .Y(men_men_n188_));
  NAi21      u0166(.An(i_4_), .B(i_12_), .Y(men_men_n189_));
  NO4        u0167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n186_), .D(men_men_n25_), .Y(men_men_n190_));
  NO3        u0168(.A(men_men_n190_), .B(men_men_n183_), .C(men_men_n177_), .Y(men_men_n191_));
  INV        u0169(.A(i_8_), .Y(men_men_n192_));
  NO2        u0170(.A(men_men_n192_), .B(i_7_), .Y(men_men_n193_));
  NA2        u0171(.A(men_men_n193_), .B(i_6_), .Y(men_men_n194_));
  NO3        u0172(.A(i_3_), .B(men_men_n82_), .C(men_men_n48_), .Y(men_men_n195_));
  NA2        u0173(.A(men_men_n195_), .B(men_men_n111_), .Y(men_men_n196_));
  NO3        u0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n197_));
  NA3        u0175(.A(men_men_n197_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n198_));
  NO3        u0176(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n199_));
  OAI210     u0177(.A0(men_men_n94_), .A1(i_12_), .B0(men_men_n199_), .Y(men_men_n200_));
  AOI210     u0178(.A0(men_men_n200_), .A1(men_men_n198_), .B0(men_men_n196_), .Y(men_men_n201_));
  NO2        u0179(.A(i_3_), .B(i_8_), .Y(men_men_n202_));
  NO3        u0180(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n203_));
  NA3        u0181(.A(men_men_n203_), .B(men_men_n202_), .C(men_men_n39_), .Y(men_men_n204_));
  NO2        u0182(.A(men_men_n101_), .B(men_men_n58_), .Y(men_men_n205_));
  INV        u0183(.A(men_men_n205_), .Y(men_men_n206_));
  NO2        u0184(.A(i_13_), .B(i_9_), .Y(men_men_n207_));
  NAi21      u0185(.An(i_12_), .B(i_3_), .Y(men_men_n208_));
  NO2        u0186(.A(men_men_n44_), .B(i_5_), .Y(men_men_n209_));
  NO3        u0187(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n210_));
  NA2        u0188(.A(men_men_n210_), .B(i_10_), .Y(men_men_n211_));
  OAI220     u0189(.A0(men_men_n211_), .A1(men_men_n208_), .B0(men_men_n206_), .B1(men_men_n204_), .Y(men_men_n212_));
  AOI210     u0190(.A0(men_men_n212_), .A1(i_7_), .B0(men_men_n201_), .Y(men_men_n213_));
  OAI220     u0191(.A0(men_men_n213_), .A1(i_4_), .B0(men_men_n194_), .B1(men_men_n191_), .Y(men_men_n214_));
  NAi21      u0192(.An(i_12_), .B(i_7_), .Y(men_men_n215_));
  NA3        u0193(.A(i_13_), .B(men_men_n192_), .C(i_10_), .Y(men_men_n216_));
  NO2        u0194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NA2        u0195(.A(i_0_), .B(i_5_), .Y(men_men_n218_));
  NA2        u0196(.A(men_men_n218_), .B(men_men_n102_), .Y(men_men_n219_));
  OAI220     u0197(.A0(men_men_n219_), .A1(men_men_n188_), .B0(i_2_), .B1(men_men_n132_), .Y(men_men_n220_));
  NAi31      u0198(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n221_));
  NO2        u0199(.A(men_men_n36_), .B(i_13_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n70_), .B(men_men_n26_), .Y(men_men_n223_));
  NO2        u0201(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n224_));
  NA3        u0202(.A(men_men_n224_), .B(men_men_n223_), .C(men_men_n222_), .Y(men_men_n225_));
  INV        u0203(.A(i_13_), .Y(men_men_n226_));
  NO2        u0204(.A(i_12_), .B(men_men_n226_), .Y(men_men_n227_));
  NA3        u0205(.A(men_men_n227_), .B(men_men_n197_), .C(men_men_n195_), .Y(men_men_n228_));
  OAI210     u0206(.A0(men_men_n225_), .A1(men_men_n221_), .B0(men_men_n228_), .Y(men_men_n229_));
  AOI220     u0207(.A0(men_men_n229_), .A1(men_men_n141_), .B0(men_men_n220_), .B1(men_men_n217_), .Y(men_men_n230_));
  NO2        u0208(.A(i_12_), .B(men_men_n37_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n181_), .B(i_4_), .Y(men_men_n232_));
  NA2        u0210(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  OR2        u0211(.A(i_8_), .B(i_7_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n234_), .B(men_men_n82_), .Y(men_men_n235_));
  NO2        u0213(.A(men_men_n53_), .B(i_1_), .Y(men_men_n236_));
  NA2        u0214(.A(men_men_n236_), .B(men_men_n235_), .Y(men_men_n237_));
  INV        u0215(.A(i_12_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n44_), .B(men_men_n238_), .Y(men_men_n239_));
  NO3        u0217(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n240_));
  NA2        u0218(.A(i_2_), .B(i_1_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n237_), .B(men_men_n233_), .Y(men_men_n242_));
  NO3        u0220(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n243_));
  NAi21      u0221(.An(i_4_), .B(i_3_), .Y(men_men_n244_));
  NO2        u0222(.A(i_0_), .B(i_6_), .Y(men_men_n245_));
  NOi41      u0223(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n246_));
  NA2        u0224(.A(men_men_n246_), .B(men_men_n245_), .Y(men_men_n247_));
  NO2        u0225(.A(men_men_n241_), .B(men_men_n181_), .Y(men_men_n248_));
  NAi21      u0226(.An(men_men_n247_), .B(men_men_n248_), .Y(men_men_n249_));
  INV        u0227(.A(men_men_n249_), .Y(men_men_n250_));
  NO2        u0228(.A(men_men_n250_), .B(men_men_n242_), .Y(men_men_n251_));
  NO2        u0229(.A(i_11_), .B(men_men_n226_), .Y(men_men_n252_));
  NOi21      u0230(.An(i_1_), .B(i_6_), .Y(men_men_n253_));
  NAi21      u0231(.An(i_3_), .B(i_7_), .Y(men_men_n254_));
  NA2        u0232(.A(men_men_n238_), .B(i_9_), .Y(men_men_n255_));
  OR4        u0233(.A(men_men_n255_), .B(men_men_n254_), .C(men_men_n253_), .D(men_men_n184_), .Y(men_men_n256_));
  NO2        u0234(.A(i_12_), .B(i_3_), .Y(men_men_n257_));
  NA2        u0235(.A(men_men_n70_), .B(i_5_), .Y(men_men_n258_));
  NA2        u0236(.A(i_3_), .B(i_9_), .Y(men_men_n259_));
  NAi21      u0237(.An(i_7_), .B(i_10_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n260_), .B(men_men_n259_), .Y(men_men_n261_));
  NA3        u0239(.A(men_men_n261_), .B(men_men_n258_), .C(men_men_n64_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n262_), .B(men_men_n256_), .Y(men_men_n263_));
  NA3        u0241(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n264_));
  INV        u0242(.A(men_men_n142_), .Y(men_men_n265_));
  NA2        u0243(.A(men_men_n238_), .B(i_13_), .Y(men_men_n266_));
  NO2        u0244(.A(men_men_n266_), .B(men_men_n72_), .Y(men_men_n267_));
  AOI220     u0245(.A0(men_men_n267_), .A1(men_men_n265_), .B0(men_men_n263_), .B1(men_men_n252_), .Y(men_men_n268_));
  NO2        u0246(.A(men_men_n234_), .B(men_men_n37_), .Y(men_men_n269_));
  NA2        u0247(.A(i_12_), .B(i_6_), .Y(men_men_n270_));
  OR2        u0248(.A(i_13_), .B(i_9_), .Y(men_men_n271_));
  NO3        u0249(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n48_), .Y(men_men_n272_));
  NO2        u0250(.A(men_men_n244_), .B(i_2_), .Y(men_men_n273_));
  NA3        u0251(.A(men_men_n273_), .B(men_men_n272_), .C(men_men_n44_), .Y(men_men_n274_));
  NA2        u0252(.A(men_men_n252_), .B(i_9_), .Y(men_men_n275_));
  OAI210     u0253(.A0(men_men_n70_), .A1(men_men_n275_), .B0(men_men_n274_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n154_), .B(men_men_n63_), .Y(men_men_n277_));
  NO3        u0255(.A(i_11_), .B(men_men_n226_), .C(men_men_n25_), .Y(men_men_n278_));
  NO2        u0256(.A(men_men_n254_), .B(i_8_), .Y(men_men_n279_));
  NO2        u0257(.A(i_6_), .B(men_men_n48_), .Y(men_men_n280_));
  NA3        u0258(.A(men_men_n280_), .B(men_men_n279_), .C(men_men_n278_), .Y(men_men_n281_));
  NA3        u0259(.A(i_6_), .B(men_men_n269_), .C(men_men_n227_), .Y(men_men_n282_));
  AOI210     u0260(.A0(men_men_n282_), .A1(men_men_n281_), .B0(men_men_n277_), .Y(men_men_n283_));
  AOI210     u0261(.A0(men_men_n276_), .A1(men_men_n269_), .B0(men_men_n283_), .Y(men_men_n284_));
  NA4        u0262(.A(men_men_n284_), .B(men_men_n268_), .C(men_men_n251_), .D(men_men_n230_), .Y(men_men_n285_));
  NO3        u0263(.A(i_12_), .B(men_men_n226_), .C(men_men_n37_), .Y(men_men_n286_));
  INV        u0264(.A(men_men_n286_), .Y(men_men_n287_));
  NA2        u0265(.A(i_8_), .B(men_men_n99_), .Y(men_men_n288_));
  NOi21      u0266(.An(men_men_n163_), .B(men_men_n82_), .Y(men_men_n289_));
  NO3        u0267(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n290_));
  AOI220     u0268(.A0(men_men_n290_), .A1(men_men_n195_), .B0(men_men_n289_), .B1(men_men_n236_), .Y(men_men_n291_));
  NO2        u0269(.A(men_men_n291_), .B(men_men_n288_), .Y(men_men_n292_));
  NO2        u0270(.A(men_men_n241_), .B(i_0_), .Y(men_men_n293_));
  AOI220     u0271(.A0(men_men_n293_), .A1(men_men_n193_), .B0(i_1_), .B1(men_men_n141_), .Y(men_men_n294_));
  NA2        u0272(.A(men_men_n280_), .B(men_men_n26_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n296_));
  NA2        u0274(.A(i_0_), .B(i_1_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n297_), .B(i_2_), .Y(men_men_n298_));
  NO2        u0276(.A(men_men_n59_), .B(i_6_), .Y(men_men_n299_));
  NA3        u0277(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n163_), .Y(men_men_n300_));
  OAI210     u0278(.A0(men_men_n165_), .A1(men_men_n142_), .B0(men_men_n300_), .Y(men_men_n301_));
  NO3        u0279(.A(men_men_n301_), .B(men_men_n296_), .C(men_men_n292_), .Y(men_men_n302_));
  NO2        u0280(.A(i_3_), .B(i_10_), .Y(men_men_n303_));
  NA3        u0281(.A(men_men_n303_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n304_));
  NO2        u0282(.A(i_2_), .B(men_men_n99_), .Y(men_men_n305_));
  NA2        u0283(.A(i_1_), .B(men_men_n36_), .Y(men_men_n306_));
  NOi21      u0284(.An(men_men_n218_), .B(men_men_n101_), .Y(men_men_n307_));
  NA3        u0285(.A(men_men_n307_), .B(i_1_), .C(men_men_n305_), .Y(men_men_n308_));
  AN2        u0286(.A(i_3_), .B(i_10_), .Y(men_men_n309_));
  NA3        u0287(.A(men_men_n309_), .B(men_men_n175_), .C(men_men_n173_), .Y(men_men_n310_));
  NO2        u0288(.A(i_5_), .B(men_men_n37_), .Y(men_men_n311_));
  NO2        u0289(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n312_));
  OR2        u0290(.A(men_men_n308_), .B(men_men_n304_), .Y(men_men_n313_));
  OAI220     u0291(.A0(men_men_n313_), .A1(i_6_), .B0(men_men_n302_), .B1(men_men_n287_), .Y(men_men_n314_));
  NO4        u0292(.A(men_men_n314_), .B(men_men_n285_), .C(men_men_n214_), .D(men_men_n168_), .Y(men_men_n315_));
  NO3        u0293(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n316_));
  NO2        u0294(.A(men_men_n59_), .B(men_men_n82_), .Y(men_men_n317_));
  NA2        u0295(.A(men_men_n293_), .B(men_men_n317_), .Y(men_men_n318_));
  NO3        u0296(.A(i_6_), .B(men_men_n192_), .C(i_7_), .Y(men_men_n319_));
  NA2        u0297(.A(men_men_n319_), .B(men_men_n197_), .Y(men_men_n320_));
  AOI210     u0298(.A0(men_men_n320_), .A1(men_men_n318_), .B0(i_5_), .Y(men_men_n321_));
  NO2        u0299(.A(i_2_), .B(i_3_), .Y(men_men_n322_));
  OR2        u0300(.A(i_0_), .B(i_5_), .Y(men_men_n323_));
  NA2        u0301(.A(men_men_n218_), .B(men_men_n323_), .Y(men_men_n324_));
  NA4        u0302(.A(men_men_n324_), .B(men_men_n235_), .C(men_men_n322_), .D(i_1_), .Y(men_men_n325_));
  NA3        u0303(.A(men_men_n293_), .B(men_men_n289_), .C(men_men_n111_), .Y(men_men_n326_));
  NAi21      u0304(.An(i_8_), .B(i_7_), .Y(men_men_n327_));
  NO2        u0305(.A(men_men_n327_), .B(i_6_), .Y(men_men_n328_));
  NO2        u0306(.A(men_men_n157_), .B(men_men_n46_), .Y(men_men_n329_));
  NA3        u0307(.A(men_men_n329_), .B(men_men_n328_), .C(men_men_n163_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n330_), .B(men_men_n326_), .C(men_men_n325_), .Y(men_men_n331_));
  OAI210     u0309(.A0(men_men_n331_), .A1(men_men_n321_), .B0(i_4_), .Y(men_men_n332_));
  NO2        u0310(.A(i_12_), .B(i_10_), .Y(men_men_n333_));
  NOi21      u0311(.An(i_5_), .B(i_0_), .Y(men_men_n334_));
  AOI210     u0312(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n99_), .Y(men_men_n335_));
  NO3        u0313(.A(men_men_n335_), .B(men_men_n306_), .C(men_men_n127_), .Y(men_men_n336_));
  NA4        u0314(.A(men_men_n81_), .B(men_men_n36_), .C(men_men_n82_), .D(i_8_), .Y(men_men_n337_));
  NA2        u0315(.A(men_men_n336_), .B(men_men_n333_), .Y(men_men_n338_));
  NO2        u0316(.A(i_6_), .B(i_8_), .Y(men_men_n339_));
  NOi21      u0317(.An(i_0_), .B(i_2_), .Y(men_men_n340_));
  AN2        u0318(.A(men_men_n340_), .B(men_men_n339_), .Y(men_men_n341_));
  NO2        u0319(.A(i_1_), .B(i_7_), .Y(men_men_n342_));
  AO220      u0320(.A0(men_men_n342_), .A1(men_men_n341_), .B0(men_men_n328_), .B1(men_men_n236_), .Y(men_men_n343_));
  NA3        u0321(.A(men_men_n343_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n344_));
  NA3        u0322(.A(men_men_n344_), .B(men_men_n338_), .C(men_men_n332_), .Y(men_men_n345_));
  NO2        u0323(.A(i_8_), .B(men_men_n324_), .Y(men_men_n346_));
  NO2        u0324(.A(men_men_n101_), .B(men_men_n123_), .Y(men_men_n347_));
  OAI210     u0325(.A0(men_men_n347_), .A1(men_men_n346_), .B0(i_3_), .Y(men_men_n348_));
  NO2        u0326(.A(men_men_n297_), .B(men_men_n78_), .Y(men_men_n349_));
  NA2        u0327(.A(men_men_n349_), .B(men_men_n131_), .Y(men_men_n350_));
  NO2        u0328(.A(men_men_n90_), .B(men_men_n192_), .Y(men_men_n351_));
  NA3        u0329(.A(men_men_n307_), .B(men_men_n351_), .C(men_men_n63_), .Y(men_men_n352_));
  AOI210     u0330(.A0(men_men_n352_), .A1(men_men_n350_), .B0(i_7_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n192_), .B(i_9_), .Y(men_men_n354_));
  NA2        u0332(.A(men_men_n354_), .B(men_men_n205_), .Y(men_men_n355_));
  NO2        u0333(.A(men_men_n353_), .B(men_men_n296_), .Y(men_men_n356_));
  AOI210     u0334(.A0(men_men_n356_), .A1(men_men_n348_), .B0(men_men_n162_), .Y(men_men_n357_));
  AOI210     u0335(.A0(men_men_n345_), .A1(men_men_n316_), .B0(men_men_n357_), .Y(men_men_n358_));
  NOi32      u0336(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n359_));
  INV        u0337(.A(men_men_n359_), .Y(men_men_n360_));
  NAi21      u0338(.An(i_0_), .B(i_6_), .Y(men_men_n361_));
  NAi21      u0339(.An(i_1_), .B(i_5_), .Y(men_men_n362_));
  NA2        u0340(.A(men_men_n362_), .B(men_men_n361_), .Y(men_men_n363_));
  NA2        u0341(.A(men_men_n363_), .B(men_men_n25_), .Y(men_men_n364_));
  OAI210     u0342(.A0(men_men_n364_), .A1(men_men_n159_), .B0(men_men_n247_), .Y(men_men_n365_));
  NAi41      u0343(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n366_));
  OAI220     u0344(.A0(men_men_n366_), .A1(men_men_n362_), .B0(men_men_n221_), .B1(men_men_n159_), .Y(men_men_n367_));
  AOI210     u0345(.A0(men_men_n366_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n368_));
  NOi32      u0346(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n369_));
  NA2        u0347(.A(men_men_n369_), .B(men_men_n46_), .Y(men_men_n370_));
  NO2        u0348(.A(men_men_n370_), .B(i_0_), .Y(men_men_n371_));
  OR3        u0349(.A(men_men_n371_), .B(men_men_n368_), .C(men_men_n367_), .Y(men_men_n372_));
  NO2        u0350(.A(i_1_), .B(men_men_n99_), .Y(men_men_n373_));
  NAi21      u0351(.An(i_3_), .B(i_4_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n374_), .B(i_9_), .Y(men_men_n375_));
  AN2        u0353(.A(i_6_), .B(i_7_), .Y(men_men_n376_));
  OAI210     u0354(.A0(men_men_n376_), .A1(men_men_n373_), .B0(men_men_n375_), .Y(men_men_n377_));
  NA2        u0355(.A(i_2_), .B(i_7_), .Y(men_men_n378_));
  NO2        u0356(.A(men_men_n374_), .B(i_10_), .Y(men_men_n379_));
  NA3        u0357(.A(men_men_n379_), .B(men_men_n378_), .C(men_men_n245_), .Y(men_men_n380_));
  AOI210     u0358(.A0(men_men_n380_), .A1(men_men_n377_), .B0(men_men_n184_), .Y(men_men_n381_));
  AOI220     u0359(.A0(men_men_n379_), .A1(men_men_n342_), .B0(men_men_n240_), .B1(men_men_n187_), .Y(men_men_n382_));
  NO3        u0360(.A(men_men_n381_), .B(men_men_n372_), .C(men_men_n365_), .Y(men_men_n383_));
  NO2        u0361(.A(men_men_n383_), .B(men_men_n360_), .Y(men_men_n384_));
  NO2        u0362(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n385_));
  AN2        u0363(.A(i_12_), .B(i_5_), .Y(men_men_n386_));
  NO2        u0364(.A(i_4_), .B(men_men_n26_), .Y(men_men_n387_));
  NA2        u0365(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n388_));
  NO2        u0366(.A(i_11_), .B(i_6_), .Y(men_men_n389_));
  NA3        u0367(.A(men_men_n389_), .B(men_men_n329_), .C(men_men_n226_), .Y(men_men_n390_));
  NO2        u0368(.A(men_men_n390_), .B(men_men_n388_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n244_), .B(i_5_), .Y(men_men_n392_));
  NO2        u0370(.A(i_5_), .B(i_10_), .Y(men_men_n393_));
  NA2        u0371(.A(men_men_n143_), .B(men_men_n45_), .Y(men_men_n394_));
  NO2        u0372(.A(men_men_n394_), .B(men_men_n244_), .Y(men_men_n395_));
  OAI210     u0373(.A0(men_men_n395_), .A1(men_men_n391_), .B0(men_men_n385_), .Y(men_men_n396_));
  NO2        u0374(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n397_));
  INV        u0375(.A(men_men_n149_), .Y(men_men_n398_));
  OAI210     u0376(.A0(men_men_n398_), .A1(men_men_n391_), .B0(men_men_n397_), .Y(men_men_n399_));
  NO2        u0377(.A(i_3_), .B(men_men_n99_), .Y(men_men_n400_));
  NA2        u0378(.A(men_men_n303_), .B(men_men_n72_), .Y(men_men_n401_));
  NO2        u0379(.A(i_11_), .B(i_12_), .Y(men_men_n402_));
  NA2        u0380(.A(men_men_n402_), .B(men_men_n36_), .Y(men_men_n403_));
  NO2        u0381(.A(men_men_n401_), .B(men_men_n403_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n393_), .B(men_men_n238_), .Y(men_men_n405_));
  NA3        u0383(.A(men_men_n111_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n406_));
  NO2        u0384(.A(men_men_n406_), .B(men_men_n221_), .Y(men_men_n407_));
  NAi21      u0385(.An(i_13_), .B(i_0_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n408_), .B(men_men_n241_), .Y(men_men_n409_));
  OAI210     u0387(.A0(men_men_n407_), .A1(men_men_n404_), .B0(men_men_n409_), .Y(men_men_n410_));
  NA3        u0388(.A(men_men_n410_), .B(men_men_n399_), .C(men_men_n396_), .Y(men_men_n411_));
  NO3        u0389(.A(i_1_), .B(i_12_), .C(men_men_n82_), .Y(men_men_n412_));
  NO2        u0390(.A(i_0_), .B(i_11_), .Y(men_men_n413_));
  AN2        u0391(.A(i_1_), .B(i_6_), .Y(men_men_n414_));
  NOi21      u0392(.An(i_2_), .B(i_12_), .Y(men_men_n415_));
  NA2        u0393(.A(men_men_n415_), .B(men_men_n414_), .Y(men_men_n416_));
  INV        u0394(.A(men_men_n416_), .Y(men_men_n417_));
  NA2        u0395(.A(men_men_n141_), .B(i_9_), .Y(men_men_n418_));
  NO2        u0396(.A(men_men_n418_), .B(i_4_), .Y(men_men_n419_));
  NA2        u0397(.A(men_men_n417_), .B(men_men_n419_), .Y(men_men_n420_));
  OR2        u0398(.A(i_13_), .B(i_10_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n172_), .B(men_men_n122_), .Y(men_men_n422_));
  OR2        u0400(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n423_));
  NO2        u0401(.A(men_men_n99_), .B(men_men_n25_), .Y(men_men_n424_));
  NA2        u0402(.A(men_men_n286_), .B(men_men_n424_), .Y(men_men_n425_));
  INV        u0403(.A(men_men_n210_), .Y(men_men_n426_));
  OAI220     u0404(.A0(men_men_n426_), .A1(men_men_n423_), .B0(men_men_n425_), .B1(men_men_n101_), .Y(men_men_n427_));
  INV        u0405(.A(men_men_n427_), .Y(men_men_n428_));
  AOI210     u0406(.A0(men_men_n428_), .A1(men_men_n420_), .B0(men_men_n26_), .Y(men_men_n429_));
  NA2        u0407(.A(men_men_n326_), .B(men_men_n325_), .Y(men_men_n430_));
  AOI220     u0408(.A0(men_men_n299_), .A1(men_men_n290_), .B0(men_men_n293_), .B1(men_men_n317_), .Y(men_men_n431_));
  NO2        u0409(.A(men_men_n431_), .B(i_5_), .Y(men_men_n432_));
  NO2        u0410(.A(men_men_n181_), .B(men_men_n82_), .Y(men_men_n433_));
  AOI220     u0411(.A0(men_men_n433_), .A1(men_men_n298_), .B0(i_6_), .B1(men_men_n210_), .Y(men_men_n434_));
  NO2        u0412(.A(men_men_n434_), .B(men_men_n288_), .Y(men_men_n435_));
  NO3        u0413(.A(men_men_n435_), .B(men_men_n432_), .C(men_men_n430_), .Y(men_men_n436_));
  NA2        u0414(.A(men_men_n195_), .B(men_men_n94_), .Y(men_men_n437_));
  NA3        u0415(.A(men_men_n329_), .B(men_men_n163_), .C(men_men_n82_), .Y(men_men_n438_));
  AOI210     u0416(.A0(men_men_n438_), .A1(men_men_n437_), .B0(men_men_n327_), .Y(men_men_n439_));
  NA3        u0417(.A(men_men_n258_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n440_));
  NA2        u0418(.A(men_men_n299_), .B(men_men_n236_), .Y(men_men_n441_));
  OAI220     u0419(.A0(men_men_n441_), .A1(men_men_n181_), .B0(men_men_n440_), .B1(men_men_n1043_), .Y(men_men_n442_));
  NO2        u0420(.A(i_3_), .B(men_men_n48_), .Y(men_men_n443_));
  NA3        u0421(.A(men_men_n342_), .B(men_men_n341_), .C(men_men_n443_), .Y(men_men_n444_));
  NA2        u0422(.A(men_men_n319_), .B(men_men_n324_), .Y(men_men_n445_));
  OAI210     u0423(.A0(men_men_n445_), .A1(men_men_n188_), .B0(men_men_n444_), .Y(men_men_n446_));
  NO3        u0424(.A(men_men_n446_), .B(men_men_n442_), .C(men_men_n439_), .Y(men_men_n447_));
  AOI210     u0425(.A0(men_men_n447_), .A1(men_men_n436_), .B0(men_men_n275_), .Y(men_men_n448_));
  NO4        u0426(.A(men_men_n448_), .B(men_men_n429_), .C(men_men_n411_), .D(men_men_n384_), .Y(men_men_n449_));
  NO2        u0427(.A(men_men_n63_), .B(i_4_), .Y(men_men_n450_));
  NO2        u0428(.A(men_men_n70_), .B(i_13_), .Y(men_men_n451_));
  NO2        u0429(.A(i_10_), .B(i_9_), .Y(men_men_n452_));
  NAi21      u0430(.An(i_12_), .B(i_8_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n453_), .B(i_3_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n46_), .B(i_4_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n455_), .B(men_men_n102_), .Y(men_men_n456_));
  NO2        u0434(.A(men_men_n456_), .B(men_men_n204_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n312_), .B(i_0_), .Y(men_men_n458_));
  NO3        u0436(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n270_), .B(men_men_n95_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  NA2        u0439(.A(i_8_), .B(i_9_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n461_), .B(men_men_n458_), .Y(men_men_n463_));
  NO3        u0441(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n464_));
  NA3        u0442(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n465_));
  NO2        u0443(.A(men_men_n463_), .B(men_men_n457_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n298_), .B(men_men_n106_), .Y(men_men_n467_));
  OA220      u0445(.A0(men_men_n355_), .A1(men_men_n162_), .B0(men_men_n467_), .B1(men_men_n233_), .Y(men_men_n468_));
  NA2        u0446(.A(men_men_n94_), .B(i_13_), .Y(men_men_n469_));
  NA2        u0447(.A(men_men_n433_), .B(men_men_n385_), .Y(men_men_n470_));
  NO2        u0448(.A(i_2_), .B(i_13_), .Y(men_men_n471_));
  NA3        u0449(.A(men_men_n471_), .B(men_men_n161_), .C(men_men_n97_), .Y(men_men_n472_));
  OAI220     u0450(.A0(men_men_n472_), .A1(men_men_n238_), .B0(men_men_n470_), .B1(men_men_n469_), .Y(men_men_n473_));
  NO3        u0451(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n474_));
  NO2        u0452(.A(i_6_), .B(i_7_), .Y(men_men_n475_));
  NA2        u0453(.A(men_men_n475_), .B(men_men_n474_), .Y(men_men_n476_));
  NO2        u0454(.A(i_11_), .B(i_1_), .Y(men_men_n477_));
  OR2        u0455(.A(i_11_), .B(i_8_), .Y(men_men_n478_));
  NOi21      u0456(.An(i_2_), .B(i_7_), .Y(men_men_n479_));
  NAi31      u0457(.An(men_men_n478_), .B(men_men_n479_), .C(i_0_), .Y(men_men_n480_));
  NO2        u0458(.A(men_men_n421_), .B(i_6_), .Y(men_men_n481_));
  NA3        u0459(.A(men_men_n481_), .B(men_men_n450_), .C(men_men_n72_), .Y(men_men_n482_));
  NO2        u0460(.A(men_men_n482_), .B(men_men_n480_), .Y(men_men_n483_));
  NO2        u0461(.A(i_3_), .B(men_men_n192_), .Y(men_men_n484_));
  NO2        u0462(.A(i_6_), .B(i_10_), .Y(men_men_n485_));
  NA4        u0463(.A(men_men_n485_), .B(men_men_n316_), .C(men_men_n484_), .D(men_men_n238_), .Y(men_men_n486_));
  NO2        u0464(.A(men_men_n486_), .B(men_men_n155_), .Y(men_men_n487_));
  NA3        u0465(.A(men_men_n246_), .B(men_men_n171_), .C(men_men_n131_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n489_));
  NO2        u0467(.A(men_men_n157_), .B(i_3_), .Y(men_men_n490_));
  NAi31      u0468(.An(men_men_n489_), .B(men_men_n490_), .C(men_men_n227_), .Y(men_men_n491_));
  NA3        u0469(.A(men_men_n397_), .B(men_men_n178_), .C(men_men_n148_), .Y(men_men_n492_));
  NA3        u0470(.A(men_men_n492_), .B(men_men_n491_), .C(men_men_n488_), .Y(men_men_n493_));
  NO4        u0471(.A(men_men_n493_), .B(men_men_n487_), .C(men_men_n483_), .D(men_men_n473_), .Y(men_men_n494_));
  NA2        u0472(.A(men_men_n459_), .B(men_men_n386_), .Y(men_men_n495_));
  NA2        u0473(.A(men_men_n464_), .B(men_men_n393_), .Y(men_men_n496_));
  NO2        u0474(.A(men_men_n496_), .B(men_men_n225_), .Y(men_men_n497_));
  NAi21      u0475(.An(men_men_n216_), .B(men_men_n402_), .Y(men_men_n498_));
  NA2        u0476(.A(men_men_n342_), .B(men_men_n218_), .Y(men_men_n499_));
  NO2        u0477(.A(men_men_n26_), .B(i_5_), .Y(men_men_n500_));
  NO2        u0478(.A(i_0_), .B(men_men_n82_), .Y(men_men_n501_));
  NA3        u0479(.A(men_men_n501_), .B(men_men_n500_), .C(men_men_n141_), .Y(men_men_n502_));
  OAI220     u0480(.A0(men_men_n38_), .A1(men_men_n502_), .B0(men_men_n499_), .B1(men_men_n498_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n316_), .B(men_men_n240_), .Y(men_men_n504_));
  NO2        u0482(.A(men_men_n504_), .B(men_men_n440_), .Y(men_men_n505_));
  NA4        u0483(.A(men_men_n309_), .B(men_men_n224_), .C(men_men_n70_), .D(men_men_n238_), .Y(men_men_n506_));
  NO2        u0484(.A(men_men_n506_), .B(men_men_n476_), .Y(men_men_n507_));
  NO4        u0485(.A(men_men_n507_), .B(men_men_n505_), .C(men_men_n503_), .D(men_men_n497_), .Y(men_men_n508_));
  NA4        u0486(.A(men_men_n508_), .B(men_men_n494_), .C(men_men_n468_), .D(men_men_n466_), .Y(men_men_n509_));
  NA3        u0487(.A(men_men_n309_), .B(men_men_n175_), .C(men_men_n173_), .Y(men_men_n510_));
  OAI210     u0488(.A0(men_men_n304_), .A1(men_men_n179_), .B0(men_men_n510_), .Y(men_men_n511_));
  AN2        u0489(.A(men_men_n290_), .B(men_men_n235_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n512_), .B(men_men_n511_), .Y(men_men_n513_));
  NA2        u0491(.A(men_men_n121_), .B(men_men_n110_), .Y(men_men_n514_));
  AN2        u0492(.A(men_men_n514_), .B(men_men_n459_), .Y(men_men_n515_));
  OAI210     u0493(.A0(i_2_), .A1(men_men_n233_), .B0(men_men_n310_), .Y(men_men_n516_));
  AOI220     u0494(.A0(men_men_n516_), .A1(men_men_n328_), .B0(men_men_n515_), .B1(men_men_n312_), .Y(men_men_n517_));
  NA2        u0495(.A(men_men_n386_), .B(men_men_n226_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n359_), .B(men_men_n70_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n376_), .B(men_men_n369_), .Y(men_men_n520_));
  AO210      u0498(.A0(men_men_n519_), .A1(men_men_n518_), .B0(men_men_n520_), .Y(men_men_n521_));
  NO2        u0499(.A(men_men_n36_), .B(i_8_), .Y(men_men_n522_));
  INV        u0500(.A(men_men_n521_), .Y(men_men_n523_));
  OAI210     u0501(.A0(i_8_), .A1(men_men_n63_), .B0(men_men_n133_), .Y(men_men_n524_));
  AOI210     u0502(.A0(men_men_n193_), .A1(i_9_), .B0(men_men_n269_), .Y(men_men_n525_));
  NO2        u0503(.A(men_men_n525_), .B(men_men_n198_), .Y(men_men_n526_));
  AOI220     u0504(.A0(i_6_), .A1(men_men_n526_), .B0(men_men_n524_), .B1(men_men_n422_), .Y(men_men_n527_));
  NA4        u0505(.A(men_men_n527_), .B(men_men_n521_), .C(men_men_n517_), .D(men_men_n513_), .Y(men_men_n528_));
  NA2        u0506(.A(men_men_n392_), .B(men_men_n298_), .Y(men_men_n529_));
  NA2        u0507(.A(men_men_n169_), .B(men_men_n529_), .Y(men_men_n530_));
  NO2        u0508(.A(i_12_), .B(men_men_n192_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n531_), .B(men_men_n226_), .Y(men_men_n532_));
  NO3        u0510(.A(i_10_), .B(men_men_n532_), .C(men_men_n467_), .Y(men_men_n533_));
  NOi31      u0511(.An(men_men_n319_), .B(men_men_n421_), .C(men_men_n38_), .Y(men_men_n534_));
  OAI210     u0512(.A0(men_men_n534_), .A1(men_men_n533_), .B0(men_men_n530_), .Y(men_men_n535_));
  NO2        u0513(.A(i_8_), .B(i_7_), .Y(men_men_n536_));
  OAI210     u0514(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n537_), .B(men_men_n224_), .Y(men_men_n538_));
  AOI220     u0516(.A0(men_men_n329_), .A1(men_men_n39_), .B0(men_men_n236_), .B1(men_men_n207_), .Y(men_men_n539_));
  OAI220     u0517(.A0(men_men_n539_), .A1(men_men_n181_), .B0(men_men_n538_), .B1(men_men_n244_), .Y(men_men_n540_));
  NA2        u0518(.A(men_men_n44_), .B(i_10_), .Y(men_men_n541_));
  NO2        u0519(.A(men_men_n541_), .B(i_6_), .Y(men_men_n542_));
  NA3        u0520(.A(men_men_n542_), .B(men_men_n540_), .C(men_men_n536_), .Y(men_men_n543_));
  AOI220     u0521(.A0(men_men_n433_), .A1(men_men_n329_), .B0(men_men_n248_), .B1(men_men_n245_), .Y(men_men_n544_));
  OAI220     u0522(.A0(men_men_n544_), .A1(men_men_n266_), .B0(men_men_n469_), .B1(men_men_n132_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n545_), .B(men_men_n269_), .Y(men_men_n546_));
  NOi31      u0524(.An(men_men_n293_), .B(men_men_n304_), .C(men_men_n179_), .Y(men_men_n547_));
  NA3        u0525(.A(men_men_n309_), .B(men_men_n173_), .C(men_men_n94_), .Y(men_men_n548_));
  NO2        u0526(.A(men_men_n157_), .B(i_5_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n549_), .B(men_men_n322_), .Y(men_men_n550_));
  NA2        u0528(.A(men_men_n550_), .B(men_men_n548_), .Y(men_men_n551_));
  OAI210     u0529(.A0(men_men_n551_), .A1(men_men_n547_), .B0(men_men_n464_), .Y(men_men_n552_));
  NA4        u0530(.A(men_men_n552_), .B(men_men_n546_), .C(men_men_n543_), .D(men_men_n535_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n286_), .B(men_men_n81_), .Y(men_men_n554_));
  NO2        u0532(.A(men_men_n350_), .B(men_men_n554_), .Y(men_men_n555_));
  NA2        u0533(.A(men_men_n299_), .B(men_men_n290_), .Y(men_men_n556_));
  NO2        u0534(.A(men_men_n556_), .B(men_men_n172_), .Y(men_men_n557_));
  NA2        u0535(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n558_));
  NA2        u0536(.A(men_men_n452_), .B(men_men_n222_), .Y(men_men_n559_));
  NO2        u0537(.A(men_men_n558_), .B(men_men_n559_), .Y(men_men_n560_));
  NA3        u0538(.A(men_men_n531_), .B(men_men_n278_), .C(i_5_), .Y(men_men_n561_));
  NO2        u0539(.A(i_1_), .B(men_men_n561_), .Y(men_men_n562_));
  NO4        u0540(.A(men_men_n562_), .B(men_men_n560_), .C(men_men_n557_), .D(men_men_n555_), .Y(men_men_n563_));
  NO4        u0541(.A(men_men_n253_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n564_));
  NO3        u0542(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n234_), .B(men_men_n36_), .Y(men_men_n566_));
  AN2        u0544(.A(men_men_n566_), .B(men_men_n565_), .Y(men_men_n567_));
  AN2        u0545(.A(men_men_n567_), .B(men_men_n359_), .Y(men_men_n568_));
  NO2        u0546(.A(men_men_n421_), .B(i_1_), .Y(men_men_n569_));
  NOi31      u0547(.An(men_men_n569_), .B(men_men_n460_), .C(men_men_n70_), .Y(men_men_n570_));
  AN3        u0548(.A(men_men_n570_), .B(men_men_n419_), .C(men_men_n500_), .Y(men_men_n571_));
  NO2        u0549(.A(men_men_n431_), .B(men_men_n176_), .Y(men_men_n572_));
  NO3        u0550(.A(men_men_n572_), .B(men_men_n571_), .C(men_men_n568_), .Y(men_men_n573_));
  NOi21      u0551(.An(i_10_), .B(i_6_), .Y(men_men_n574_));
  NO2        u0552(.A(men_men_n82_), .B(men_men_n25_), .Y(men_men_n575_));
  NO2        u0553(.A(men_men_n113_), .B(men_men_n23_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n319_), .B(men_men_n164_), .Y(men_men_n577_));
  AOI220     u0555(.A0(men_men_n577_), .A1(men_men_n441_), .B0(men_men_n182_), .B1(men_men_n180_), .Y(men_men_n578_));
  NOi21      u0556(.An(men_men_n145_), .B(men_men_n337_), .Y(men_men_n579_));
  NO2        u0557(.A(men_men_n579_), .B(men_men_n578_), .Y(men_men_n580_));
  NO2        u0558(.A(men_men_n519_), .B(men_men_n382_), .Y(men_men_n581_));
  INV        u0559(.A(men_men_n322_), .Y(men_men_n582_));
  NO2        u0560(.A(i_12_), .B(men_men_n82_), .Y(men_men_n583_));
  NA3        u0561(.A(men_men_n583_), .B(men_men_n278_), .C(i_5_), .Y(men_men_n584_));
  NA3        u0562(.A(men_men_n389_), .B(men_men_n286_), .C(men_men_n218_), .Y(men_men_n585_));
  AOI210     u0563(.A0(men_men_n585_), .A1(men_men_n584_), .B0(men_men_n582_), .Y(men_men_n586_));
  NA2        u0564(.A(men_men_n173_), .B(i_0_), .Y(men_men_n587_));
  NO3        u0565(.A(men_men_n587_), .B(men_men_n1042_), .C(men_men_n304_), .Y(men_men_n588_));
  OR2        u0566(.A(i_2_), .B(i_5_), .Y(men_men_n589_));
  OR2        u0567(.A(men_men_n589_), .B(men_men_n414_), .Y(men_men_n590_));
  AOI210     u0568(.A0(men_men_n378_), .A1(men_men_n245_), .B0(men_men_n197_), .Y(men_men_n591_));
  AOI210     u0569(.A0(men_men_n591_), .A1(men_men_n590_), .B0(men_men_n498_), .Y(men_men_n592_));
  NO4        u0570(.A(men_men_n592_), .B(men_men_n588_), .C(men_men_n586_), .D(men_men_n581_), .Y(men_men_n593_));
  NA4        u0571(.A(men_men_n593_), .B(men_men_n580_), .C(men_men_n573_), .D(men_men_n563_), .Y(men_men_n594_));
  NO4        u0572(.A(men_men_n594_), .B(men_men_n553_), .C(men_men_n528_), .D(men_men_n509_), .Y(men_men_n595_));
  NA4        u0573(.A(men_men_n595_), .B(men_men_n449_), .C(men_men_n358_), .D(men_men_n315_), .Y(men7));
  NO2        u0574(.A(men_men_n90_), .B(men_men_n54_), .Y(men_men_n597_));
  NO2        u0575(.A(men_men_n106_), .B(men_men_n87_), .Y(men_men_n598_));
  NA2        u0576(.A(men_men_n387_), .B(men_men_n598_), .Y(men_men_n599_));
  NA2        u0577(.A(men_men_n485_), .B(men_men_n81_), .Y(men_men_n600_));
  NA2        u0578(.A(i_11_), .B(men_men_n192_), .Y(men_men_n601_));
  NA2        u0579(.A(men_men_n143_), .B(men_men_n601_), .Y(men_men_n602_));
  OAI210     u0580(.A0(men_men_n602_), .A1(men_men_n600_), .B0(men_men_n599_), .Y(men_men_n603_));
  NA3        u0581(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n238_), .B(i_4_), .Y(men_men_n605_));
  NA2        u0583(.A(i_2_), .B(men_men_n82_), .Y(men_men_n606_));
  OAI210     u0584(.A0(men_men_n85_), .A1(men_men_n202_), .B0(men_men_n203_), .Y(men_men_n607_));
  NO2        u0585(.A(i_7_), .B(men_men_n37_), .Y(men_men_n608_));
  NA2        u0586(.A(i_4_), .B(i_8_), .Y(men_men_n609_));
  AOI210     u0587(.A0(men_men_n609_), .A1(men_men_n309_), .B0(men_men_n608_), .Y(men_men_n610_));
  OAI220     u0588(.A0(men_men_n610_), .A1(men_men_n606_), .B0(men_men_n607_), .B1(i_13_), .Y(men_men_n611_));
  NO3        u0589(.A(men_men_n611_), .B(men_men_n603_), .C(men_men_n597_), .Y(men_men_n612_));
  INV        u0590(.A(men_men_n161_), .Y(men_men_n613_));
  OR2        u0591(.A(i_6_), .B(i_10_), .Y(men_men_n614_));
  NO2        u0592(.A(men_men_n614_), .B(men_men_n23_), .Y(men_men_n615_));
  OR3        u0593(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n616_));
  NO3        u0594(.A(men_men_n616_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n617_));
  INV        u0595(.A(men_men_n199_), .Y(men_men_n618_));
  NO2        u0596(.A(men_men_n617_), .B(men_men_n615_), .Y(men_men_n619_));
  OA220      u0597(.A0(men_men_n619_), .A1(men_men_n582_), .B0(men_men_n613_), .B1(men_men_n271_), .Y(men_men_n620_));
  AOI210     u0598(.A0(men_men_n620_), .A1(men_men_n612_), .B0(men_men_n63_), .Y(men_men_n621_));
  NOi21      u0599(.An(i_11_), .B(i_7_), .Y(men_men_n622_));
  AO210      u0600(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n623_), .B(men_men_n622_), .Y(men_men_n624_));
  NA3        u0602(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n625_));
  NAi21      u0603(.An(men_men_n625_), .B(i_11_), .Y(men_men_n626_));
  NO2        u0604(.A(men_men_n626_), .B(men_men_n63_), .Y(men_men_n627_));
  NA2        u0605(.A(men_men_n84_), .B(men_men_n63_), .Y(men_men_n628_));
  AO210      u0606(.A0(men_men_n628_), .A1(men_men_n382_), .B0(men_men_n40_), .Y(men_men_n629_));
  NA2        u0607(.A(men_men_n227_), .B(men_men_n63_), .Y(men_men_n630_));
  NA2        u0608(.A(men_men_n415_), .B(men_men_n31_), .Y(men_men_n631_));
  OR2        u0609(.A(men_men_n208_), .B(men_men_n106_), .Y(men_men_n632_));
  NA2        u0610(.A(men_men_n632_), .B(men_men_n631_), .Y(men_men_n633_));
  NO2        u0611(.A(men_men_n63_), .B(i_9_), .Y(men_men_n634_));
  NA2        u0612(.A(men_men_n63_), .B(men_men_n633_), .Y(men_men_n635_));
  NO2        u0613(.A(i_1_), .B(i_12_), .Y(men_men_n636_));
  NA3        u0614(.A(men_men_n635_), .B(men_men_n630_), .C(men_men_n629_), .Y(men_men_n637_));
  OAI210     u0615(.A0(men_men_n637_), .A1(men_men_n627_), .B0(i_6_), .Y(men_men_n638_));
  NO2        u0616(.A(i_6_), .B(i_11_), .Y(men_men_n639_));
  INV        u0617(.A(men_men_n461_), .Y(men_men_n640_));
  NO4        u0618(.A(men_men_n215_), .B(men_men_n127_), .C(i_13_), .D(men_men_n82_), .Y(men_men_n641_));
  NA2        u0619(.A(men_men_n641_), .B(men_men_n634_), .Y(men_men_n642_));
  NO3        u0620(.A(men_men_n614_), .B(men_men_n234_), .C(men_men_n23_), .Y(men_men_n643_));
  AOI210     u0621(.A0(i_1_), .A1(men_men_n261_), .B0(men_men_n643_), .Y(men_men_n644_));
  OAI210     u0622(.A0(men_men_n644_), .A1(men_men_n44_), .B0(men_men_n642_), .Y(men_men_n645_));
  NA3        u0623(.A(men_men_n536_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n646_));
  NA2        u0624(.A(men_men_n137_), .B(i_9_), .Y(men_men_n647_));
  NA3        u0625(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n648_));
  NO2        u0626(.A(men_men_n46_), .B(i_1_), .Y(men_men_n649_));
  NA3        u0627(.A(men_men_n649_), .B(men_men_n270_), .C(men_men_n44_), .Y(men_men_n650_));
  OAI220     u0628(.A0(men_men_n650_), .A1(men_men_n648_), .B0(men_men_n647_), .B1(men_men_n1039_), .Y(men_men_n651_));
  NA3        u0629(.A(men_men_n634_), .B(men_men_n322_), .C(i_6_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n652_), .B(men_men_n23_), .Y(men_men_n653_));
  AOI210     u0631(.A0(men_men_n477_), .A1(men_men_n424_), .B0(men_men_n243_), .Y(men_men_n654_));
  NO2        u0632(.A(men_men_n654_), .B(men_men_n606_), .Y(men_men_n655_));
  NAi21      u0633(.An(men_men_n646_), .B(men_men_n89_), .Y(men_men_n656_));
  NA2        u0634(.A(men_men_n649_), .B(men_men_n270_), .Y(men_men_n657_));
  NO2        u0635(.A(i_11_), .B(men_men_n37_), .Y(men_men_n658_));
  NA2        u0636(.A(men_men_n658_), .B(men_men_n24_), .Y(men_men_n659_));
  OAI210     u0637(.A0(men_men_n659_), .A1(men_men_n657_), .B0(men_men_n656_), .Y(men_men_n660_));
  OR4        u0638(.A(men_men_n660_), .B(men_men_n655_), .C(men_men_n653_), .D(men_men_n651_), .Y(men_men_n661_));
  NO3        u0639(.A(men_men_n661_), .B(men_men_n645_), .C(men_men_n640_), .Y(men_men_n662_));
  NO2        u0640(.A(men_men_n238_), .B(men_men_n99_), .Y(men_men_n663_));
  NO2        u0641(.A(men_men_n663_), .B(men_men_n622_), .Y(men_men_n664_));
  NA2        u0642(.A(men_men_n664_), .B(i_1_), .Y(men_men_n665_));
  NO2        u0643(.A(men_men_n665_), .B(men_men_n616_), .Y(men_men_n666_));
  NA2        u0644(.A(men_men_n666_), .B(men_men_n46_), .Y(men_men_n667_));
  NA2        u0645(.A(i_3_), .B(men_men_n192_), .Y(men_men_n668_));
  NO2        u0646(.A(men_men_n668_), .B(men_men_n113_), .Y(men_men_n669_));
  AN2        u0647(.A(men_men_n669_), .B(men_men_n542_), .Y(men_men_n670_));
  NO2        u0648(.A(men_men_n234_), .B(men_men_n44_), .Y(men_men_n671_));
  NO3        u0649(.A(men_men_n671_), .B(men_men_n312_), .C(men_men_n239_), .Y(men_men_n672_));
  NO2        u0650(.A(men_men_n116_), .B(men_men_n37_), .Y(men_men_n673_));
  NO2        u0651(.A(men_men_n673_), .B(i_6_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n82_), .B(i_9_), .Y(men_men_n675_));
  NO2        u0653(.A(men_men_n675_), .B(men_men_n63_), .Y(men_men_n676_));
  NO2        u0654(.A(men_men_n676_), .B(men_men_n636_), .Y(men_men_n677_));
  NO4        u0655(.A(men_men_n677_), .B(men_men_n674_), .C(men_men_n672_), .D(i_4_), .Y(men_men_n678_));
  NA2        u0656(.A(i_1_), .B(i_3_), .Y(men_men_n679_));
  NO2        u0657(.A(men_men_n462_), .B(men_men_n90_), .Y(men_men_n680_));
  AOI210     u0658(.A0(men_men_n671_), .A1(men_men_n574_), .B0(men_men_n680_), .Y(men_men_n681_));
  NO2        u0659(.A(men_men_n681_), .B(men_men_n679_), .Y(men_men_n682_));
  NO3        u0660(.A(men_men_n682_), .B(men_men_n678_), .C(men_men_n670_), .Y(men_men_n683_));
  NA4        u0661(.A(men_men_n683_), .B(men_men_n667_), .C(men_men_n662_), .D(men_men_n638_), .Y(men_men_n684_));
  NO3        u0662(.A(men_men_n478_), .B(i_3_), .C(i_7_), .Y(men_men_n685_));
  NOi21      u0663(.An(men_men_n685_), .B(i_10_), .Y(men_men_n686_));
  OA210      u0664(.A0(men_men_n686_), .A1(men_men_n246_), .B0(men_men_n82_), .Y(men_men_n687_));
  NA2        u0665(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n688_));
  NA3        u0666(.A(men_men_n485_), .B(men_men_n522_), .C(men_men_n46_), .Y(men_men_n689_));
  NO3        u0667(.A(men_men_n479_), .B(men_men_n609_), .C(men_men_n82_), .Y(men_men_n690_));
  NA2        u0668(.A(men_men_n690_), .B(men_men_n25_), .Y(men_men_n691_));
  NA3        u0669(.A(men_men_n161_), .B(men_men_n81_), .C(men_men_n82_), .Y(men_men_n692_));
  NA4        u0670(.A(men_men_n692_), .B(men_men_n691_), .C(men_men_n689_), .D(men_men_n688_), .Y(men_men_n693_));
  OAI210     u0671(.A0(men_men_n693_), .A1(men_men_n687_), .B0(i_1_), .Y(men_men_n694_));
  AOI210     u0672(.A0(men_men_n270_), .A1(men_men_n95_), .B0(i_1_), .Y(men_men_n695_));
  NO2        u0673(.A(men_men_n374_), .B(i_2_), .Y(men_men_n696_));
  NA2        u0674(.A(men_men_n696_), .B(men_men_n695_), .Y(men_men_n697_));
  OAI210     u0675(.A0(men_men_n652_), .A1(men_men_n453_), .B0(men_men_n697_), .Y(men_men_n698_));
  INV        u0676(.A(men_men_n698_), .Y(men_men_n699_));
  AOI210     u0677(.A0(men_men_n699_), .A1(men_men_n694_), .B0(i_13_), .Y(men_men_n700_));
  OR2        u0678(.A(i_11_), .B(i_7_), .Y(men_men_n701_));
  NA3        u0679(.A(men_men_n701_), .B(men_men_n104_), .C(men_men_n137_), .Y(men_men_n702_));
  AOI220     u0680(.A0(men_men_n471_), .A1(men_men_n161_), .B0(men_men_n455_), .B1(men_men_n137_), .Y(men_men_n703_));
  OAI210     u0681(.A0(men_men_n703_), .A1(men_men_n44_), .B0(men_men_n702_), .Y(men_men_n704_));
  NA2        u0682(.A(men_men_n246_), .B(men_men_n130_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(men_men_n40_), .Y(men_men_n706_));
  AOI210     u0684(.A0(men_men_n704_), .A1(men_men_n339_), .B0(men_men_n706_), .Y(men_men_n707_));
  AOI220     u0685(.A0(i_7_), .A1(men_men_n69_), .B0(men_men_n389_), .B1(men_men_n649_), .Y(men_men_n708_));
  NO2        u0686(.A(men_men_n708_), .B(men_men_n244_), .Y(men_men_n709_));
  AOI210     u0687(.A0(men_men_n453_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n710_));
  NA2        u0688(.A(men_men_n126_), .B(i_13_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n648_), .B(men_men_n113_), .Y(men_men_n712_));
  INV        u0690(.A(men_men_n712_), .Y(men_men_n713_));
  OAI220     u0691(.A0(men_men_n713_), .A1(men_men_n68_), .B0(men_men_n711_), .B1(men_men_n695_), .Y(men_men_n714_));
  NO3        u0692(.A(men_men_n68_), .B(men_men_n32_), .C(men_men_n99_), .Y(men_men_n715_));
  NA2        u0693(.A(men_men_n26_), .B(men_men_n192_), .Y(men_men_n716_));
  NA2        u0694(.A(men_men_n716_), .B(i_7_), .Y(men_men_n717_));
  NO3        u0695(.A(men_men_n479_), .B(men_men_n238_), .C(men_men_n82_), .Y(men_men_n718_));
  AOI210     u0696(.A0(men_men_n718_), .A1(men_men_n717_), .B0(men_men_n715_), .Y(men_men_n719_));
  NO2        u0697(.A(men_men_n719_), .B(men_men_n618_), .Y(men_men_n720_));
  NO3        u0698(.A(men_men_n720_), .B(men_men_n714_), .C(men_men_n709_), .Y(men_men_n721_));
  OR2        u0699(.A(i_11_), .B(i_6_), .Y(men_men_n722_));
  NA3        u0700(.A(men_men_n605_), .B(men_men_n716_), .C(i_7_), .Y(men_men_n723_));
  AOI210     u0701(.A0(men_men_n723_), .A1(men_men_n713_), .B0(men_men_n722_), .Y(men_men_n724_));
  NA2        u0702(.A(men_men_n639_), .B(i_13_), .Y(men_men_n725_));
  NAi21      u0703(.An(i_11_), .B(i_12_), .Y(men_men_n726_));
  NOi41      u0704(.An(men_men_n109_), .B(men_men_n726_), .C(i_13_), .D(men_men_n82_), .Y(men_men_n727_));
  NO3        u0705(.A(men_men_n479_), .B(men_men_n583_), .C(men_men_n609_), .Y(men_men_n728_));
  AOI220     u0706(.A0(men_men_n728_), .A1(men_men_n316_), .B0(men_men_n727_), .B1(men_men_n192_), .Y(men_men_n729_));
  NA2        u0707(.A(men_men_n729_), .B(men_men_n725_), .Y(men_men_n730_));
  OAI210     u0708(.A0(men_men_n730_), .A1(men_men_n724_), .B0(men_men_n63_), .Y(men_men_n731_));
  NA2        u0709(.A(i_8_), .B(men_men_n25_), .Y(men_men_n732_));
  NO3        u0710(.A(men_men_n732_), .B(men_men_n387_), .C(men_men_n605_), .Y(men_men_n733_));
  OAI210     u0711(.A0(men_men_n733_), .A1(men_men_n375_), .B0(men_men_n373_), .Y(men_men_n734_));
  NO2        u0712(.A(men_men_n127_), .B(i_2_), .Y(men_men_n735_));
  NA2        u0713(.A(men_men_n735_), .B(men_men_n636_), .Y(men_men_n736_));
  NA2        u0714(.A(men_men_n736_), .B(men_men_n734_), .Y(men_men_n737_));
  NA3        u0715(.A(men_men_n737_), .B(men_men_n45_), .C(men_men_n226_), .Y(men_men_n738_));
  NA4        u0716(.A(men_men_n738_), .B(men_men_n731_), .C(men_men_n721_), .D(men_men_n707_), .Y(men_men_n739_));
  OR4        u0717(.A(men_men_n739_), .B(men_men_n700_), .C(men_men_n684_), .D(men_men_n621_), .Y(men5));
  AOI210     u0718(.A0(men_men_n664_), .A1(men_men_n273_), .B0(men_men_n422_), .Y(men_men_n741_));
  NO3        u0719(.A(i_11_), .B(men_men_n238_), .C(i_13_), .Y(men_men_n742_));
  NO2        u0720(.A(men_men_n123_), .B(men_men_n23_), .Y(men_men_n743_));
  NA2        u0721(.A(i_12_), .B(i_8_), .Y(men_men_n744_));
  OAI210     u0722(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n744_), .Y(men_men_n745_));
  INV        u0723(.A(men_men_n452_), .Y(men_men_n746_));
  AOI220     u0724(.A0(men_men_n322_), .A1(men_men_n576_), .B0(men_men_n745_), .B1(men_men_n743_), .Y(men_men_n747_));
  INV        u0725(.A(men_men_n747_), .Y(men_men_n748_));
  NO2        u0726(.A(men_men_n748_), .B(men_men_n1041_), .Y(men_men_n749_));
  INV        u0727(.A(men_men_n171_), .Y(men_men_n750_));
  INV        u0728(.A(men_men_n246_), .Y(men_men_n751_));
  OAI210     u0729(.A0(men_men_n696_), .A1(men_men_n454_), .B0(men_men_n109_), .Y(men_men_n752_));
  AOI210     u0730(.A0(men_men_n752_), .A1(men_men_n751_), .B0(men_men_n750_), .Y(men_men_n753_));
  NO2        u0731(.A(men_men_n462_), .B(men_men_n26_), .Y(men_men_n754_));
  NO2        u0732(.A(men_men_n754_), .B(men_men_n424_), .Y(men_men_n755_));
  NA2        u0733(.A(men_men_n755_), .B(i_2_), .Y(men_men_n756_));
  INV        u0734(.A(men_men_n756_), .Y(men_men_n757_));
  AOI210     u0735(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n421_), .Y(men_men_n758_));
  AOI210     u0736(.A0(men_men_n758_), .A1(men_men_n757_), .B0(men_men_n753_), .Y(men_men_n759_));
  NO2        u0737(.A(men_men_n189_), .B(men_men_n124_), .Y(men_men_n760_));
  OAI210     u0738(.A0(men_men_n760_), .A1(men_men_n743_), .B0(i_2_), .Y(men_men_n761_));
  NO2        u0739(.A(men_men_n761_), .B(men_men_n192_), .Y(men_men_n762_));
  OA210      u0740(.A0(men_men_n624_), .A1(men_men_n125_), .B0(i_13_), .Y(men_men_n763_));
  NA2        u0741(.A(men_men_n199_), .B(men_men_n202_), .Y(men_men_n764_));
  NA2        u0742(.A(men_men_n151_), .B(men_men_n601_), .Y(men_men_n765_));
  AOI210     u0743(.A0(men_men_n765_), .A1(men_men_n764_), .B0(men_men_n378_), .Y(men_men_n766_));
  AOI210     u0744(.A0(men_men_n208_), .A1(men_men_n147_), .B0(men_men_n522_), .Y(men_men_n767_));
  NA2        u0745(.A(men_men_n767_), .B(men_men_n424_), .Y(men_men_n768_));
  NO2        u0746(.A(men_men_n100_), .B(men_men_n44_), .Y(men_men_n769_));
  INV        u0747(.A(men_men_n305_), .Y(men_men_n770_));
  NA4        u0748(.A(men_men_n770_), .B(men_men_n309_), .C(men_men_n123_), .D(men_men_n42_), .Y(men_men_n771_));
  OAI210     u0749(.A0(men_men_n771_), .A1(men_men_n769_), .B0(men_men_n768_), .Y(men_men_n772_));
  NO4        u0750(.A(men_men_n772_), .B(men_men_n766_), .C(men_men_n763_), .D(men_men_n762_), .Y(men_men_n773_));
  NA2        u0751(.A(men_men_n576_), .B(men_men_n28_), .Y(men_men_n774_));
  NA2        u0752(.A(men_men_n742_), .B(men_men_n279_), .Y(men_men_n775_));
  NA2        u0753(.A(men_men_n775_), .B(men_men_n774_), .Y(men_men_n776_));
  NO2        u0754(.A(men_men_n62_), .B(i_12_), .Y(men_men_n777_));
  NO2        u0755(.A(men_men_n777_), .B(men_men_n125_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n778_), .B(men_men_n601_), .Y(men_men_n779_));
  AOI220     u0757(.A0(men_men_n779_), .A1(men_men_n36_), .B0(men_men_n776_), .B1(men_men_n46_), .Y(men_men_n780_));
  NA4        u0758(.A(men_men_n780_), .B(men_men_n773_), .C(men_men_n759_), .D(men_men_n749_), .Y(men6));
  NA2        u0759(.A(men_men_n1044_), .B(men_men_n735_), .Y(men_men_n782_));
  NA4        u0760(.A(men_men_n393_), .B(men_men_n484_), .C(men_men_n68_), .D(men_men_n99_), .Y(men_men_n783_));
  INV        u0761(.A(men_men_n783_), .Y(men_men_n784_));
  NO2        u0762(.A(men_men_n221_), .B(men_men_n489_), .Y(men_men_n785_));
  NO2        u0763(.A(i_11_), .B(i_9_), .Y(men_men_n786_));
  NO2        u0764(.A(men_men_n784_), .B(men_men_n334_), .Y(men_men_n787_));
  AO210      u0765(.A0(men_men_n787_), .A1(men_men_n782_), .B0(i_12_), .Y(men_men_n788_));
  NA2        u0766(.A(men_men_n379_), .B(men_men_n342_), .Y(men_men_n789_));
  NA2        u0767(.A(men_men_n583_), .B(men_men_n63_), .Y(men_men_n790_));
  NA2        u0768(.A(men_men_n686_), .B(men_men_n68_), .Y(men_men_n791_));
  NA4        u0769(.A(men_men_n628_), .B(men_men_n791_), .C(men_men_n790_), .D(men_men_n789_), .Y(men_men_n792_));
  INV        u0770(.A(men_men_n196_), .Y(men_men_n793_));
  AOI220     u0771(.A0(men_men_n793_), .A1(men_men_n786_), .B0(men_men_n792_), .B1(men_men_n70_), .Y(men_men_n794_));
  INV        u0772(.A(men_men_n333_), .Y(men_men_n795_));
  NA2        u0773(.A(men_men_n72_), .B(men_men_n130_), .Y(men_men_n796_));
  NO2        u0774(.A(men_men_n796_), .B(men_men_n795_), .Y(men_men_n797_));
  NA2        u0775(.A(men_men_n1040_), .B(men_men_n777_), .Y(men_men_n798_));
  AOI210     u0776(.A0(men_men_n798_), .A1(men_men_n520_), .B0(men_men_n184_), .Y(men_men_n799_));
  INV        u0777(.A(i_11_), .Y(men_men_n800_));
  NA3        u0778(.A(men_men_n800_), .B(men_men_n475_), .C(men_men_n393_), .Y(men_men_n801_));
  NAi32      u0779(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n802_));
  AOI210     u0780(.A0(men_men_n722_), .A1(men_men_n83_), .B0(men_men_n802_), .Y(men_men_n803_));
  OAI210     u0781(.A0(men_men_n685_), .A1(men_men_n566_), .B0(men_men_n565_), .Y(men_men_n804_));
  NAi31      u0782(.An(men_men_n803_), .B(men_men_n804_), .C(men_men_n801_), .Y(men_men_n805_));
  OR3        u0783(.A(men_men_n805_), .B(men_men_n799_), .C(men_men_n797_), .Y(men_men_n806_));
  NA3        u0784(.A(men_men_n354_), .B(men_men_n257_), .C(i_7_), .Y(men_men_n807_));
  NA3        u0785(.A(men_men_n454_), .B(men_men_n146_), .C(men_men_n67_), .Y(men_men_n808_));
  OR2        u0786(.A(men_men_n746_), .B(men_men_n36_), .Y(men_men_n809_));
  NA3        u0787(.A(men_men_n809_), .B(men_men_n808_), .C(men_men_n807_), .Y(men_men_n810_));
  OAI210     u0788(.A0(i_6_), .A1(i_11_), .B0(men_men_n83_), .Y(men_men_n811_));
  AOI220     u0789(.A0(men_men_n811_), .A1(men_men_n565_), .B0(men_men_n785_), .B1(men_men_n717_), .Y(men_men_n812_));
  NA3        u0790(.A(men_men_n378_), .B(men_men_n240_), .C(men_men_n146_), .Y(men_men_n813_));
  NA3        u0791(.A(men_men_n813_), .B(men_men_n812_), .C(men_men_n607_), .Y(men_men_n814_));
  AO210      u0792(.A0(men_men_n522_), .A1(men_men_n46_), .B0(men_men_n84_), .Y(men_men_n815_));
  NA3        u0793(.A(men_men_n815_), .B(men_men_n485_), .C(men_men_n218_), .Y(men_men_n816_));
  INV        u0794(.A(men_men_n564_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n614_), .B(men_men_n100_), .Y(men_men_n818_));
  OAI210     u0796(.A0(men_men_n818_), .A1(men_men_n110_), .B0(men_men_n413_), .Y(men_men_n819_));
  INV        u0797(.A(men_men_n590_), .Y(men_men_n820_));
  NA3        u0798(.A(men_men_n820_), .B(men_men_n333_), .C(i_7_), .Y(men_men_n821_));
  NA4        u0799(.A(men_men_n821_), .B(men_men_n819_), .C(men_men_n817_), .D(men_men_n816_), .Y(men_men_n822_));
  NO4        u0800(.A(men_men_n822_), .B(men_men_n814_), .C(men_men_n810_), .D(men_men_n806_), .Y(men_men_n823_));
  NA4        u0801(.A(men_men_n823_), .B(men_men_n794_), .C(men_men_n788_), .D(men_men_n383_), .Y(men3));
  NA2        u0802(.A(i_12_), .B(i_10_), .Y(men_men_n825_));
  NA2        u0803(.A(i_6_), .B(i_7_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n826_), .B(i_0_), .Y(men_men_n827_));
  NO2        u0805(.A(i_11_), .B(men_men_n238_), .Y(men_men_n828_));
  OAI210     u0806(.A0(men_men_n827_), .A1(men_men_n293_), .B0(men_men_n828_), .Y(men_men_n829_));
  NO2        u0807(.A(men_men_n829_), .B(men_men_n192_), .Y(men_men_n830_));
  NO3        u0808(.A(men_men_n458_), .B(men_men_n87_), .C(men_men_n44_), .Y(men_men_n831_));
  OA210      u0809(.A0(men_men_n831_), .A1(men_men_n830_), .B0(men_men_n173_), .Y(men_men_n832_));
  NA3        u0810(.A(men_men_n813_), .B(men_men_n607_), .C(men_men_n377_), .Y(men_men_n833_));
  NA2        u0811(.A(men_men_n833_), .B(men_men_n39_), .Y(men_men_n834_));
  NO2        u0812(.A(men_men_n632_), .B(men_men_n462_), .Y(men_men_n835_));
  NA2        u0813(.A(men_men_n415_), .B(men_men_n45_), .Y(men_men_n836_));
  AN2        u0814(.A(men_men_n460_), .B(men_men_n55_), .Y(men_men_n837_));
  NO2        u0815(.A(men_men_n837_), .B(men_men_n835_), .Y(men_men_n838_));
  AOI210     u0816(.A0(men_men_n838_), .A1(men_men_n834_), .B0(men_men_n48_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n184_), .B(men_men_n574_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n710_), .B(men_men_n675_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n340_), .B(men_men_n443_), .Y(men_men_n842_));
  OAI220     u0820(.A0(men_men_n842_), .A1(men_men_n841_), .B0(men_men_n840_), .B1(men_men_n63_), .Y(men_men_n843_));
  NOi21      u0821(.An(i_5_), .B(i_9_), .Y(men_men_n844_));
  NA2        u0822(.A(men_men_n844_), .B(men_men_n451_), .Y(men_men_n845_));
  AOI210     u0823(.A0(men_men_n270_), .A1(men_men_n477_), .B0(men_men_n690_), .Y(men_men_n846_));
  NO2        u0824(.A(men_men_n174_), .B(men_men_n147_), .Y(men_men_n847_));
  NA2        u0825(.A(men_men_n847_), .B(men_men_n245_), .Y(men_men_n848_));
  OAI220     u0826(.A0(men_men_n848_), .A1(men_men_n179_), .B0(men_men_n846_), .B1(men_men_n845_), .Y(men_men_n849_));
  NO4        u0827(.A(men_men_n849_), .B(men_men_n843_), .C(men_men_n839_), .D(men_men_n832_), .Y(men_men_n850_));
  NA2        u0828(.A(men_men_n184_), .B(men_men_n24_), .Y(men_men_n851_));
  NO2        u0829(.A(men_men_n673_), .B(men_men_n598_), .Y(men_men_n852_));
  NO2        u0830(.A(men_men_n852_), .B(men_men_n851_), .Y(men_men_n853_));
  NA2        u0831(.A(men_men_n316_), .B(men_men_n128_), .Y(men_men_n854_));
  NAi21      u0832(.An(men_men_n162_), .B(men_men_n443_), .Y(men_men_n855_));
  NO2        u0833(.A(men_men_n854_), .B(men_men_n405_), .Y(men_men_n856_));
  NO2        u0834(.A(men_men_n856_), .B(men_men_n853_), .Y(men_men_n857_));
  NA2        u0835(.A(men_men_n575_), .B(i_0_), .Y(men_men_n858_));
  NO3        u0836(.A(men_men_n858_), .B(men_men_n388_), .C(men_men_n85_), .Y(men_men_n859_));
  NO4        u0837(.A(men_men_n589_), .B(men_men_n215_), .C(men_men_n421_), .D(men_men_n414_), .Y(men_men_n860_));
  AOI210     u0838(.A0(men_men_n860_), .A1(i_11_), .B0(men_men_n859_), .Y(men_men_n861_));
  NA2        u0839(.A(men_men_n742_), .B(men_men_n334_), .Y(men_men_n862_));
  AOI210     u0840(.A0(men_men_n485_), .A1(men_men_n85_), .B0(men_men_n58_), .Y(men_men_n863_));
  OAI220     u0841(.A0(men_men_n863_), .A1(men_men_n862_), .B0(men_men_n659_), .B1(men_men_n538_), .Y(men_men_n864_));
  NA2        u0842(.A(i_0_), .B(i_10_), .Y(men_men_n865_));
  OAI210     u0843(.A0(men_men_n865_), .A1(men_men_n82_), .B0(men_men_n541_), .Y(men_men_n866_));
  NO4        u0844(.A(men_men_n113_), .B(men_men_n58_), .C(men_men_n668_), .D(i_5_), .Y(men_men_n867_));
  AN2        u0845(.A(men_men_n867_), .B(men_men_n866_), .Y(men_men_n868_));
  AOI220     u0846(.A0(men_men_n340_), .A1(men_men_n96_), .B0(men_men_n184_), .B1(men_men_n81_), .Y(men_men_n869_));
  NA2        u0847(.A(men_men_n569_), .B(i_4_), .Y(men_men_n870_));
  NA2        u0848(.A(men_men_n187_), .B(men_men_n202_), .Y(men_men_n871_));
  OAI220     u0849(.A0(men_men_n871_), .A1(men_men_n862_), .B0(men_men_n870_), .B1(men_men_n869_), .Y(men_men_n872_));
  NO3        u0850(.A(men_men_n872_), .B(men_men_n868_), .C(men_men_n864_), .Y(men_men_n873_));
  NA3        u0851(.A(men_men_n873_), .B(men_men_n861_), .C(men_men_n857_), .Y(men_men_n874_));
  NO2        u0852(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n875_));
  NA2        u0853(.A(i_11_), .B(i_9_), .Y(men_men_n876_));
  NO3        u0854(.A(i_12_), .B(men_men_n876_), .C(men_men_n606_), .Y(men_men_n877_));
  AN2        u0855(.A(men_men_n877_), .B(men_men_n875_), .Y(men_men_n878_));
  NA2        u0856(.A(men_men_n397_), .B(men_men_n178_), .Y(men_men_n879_));
  NA2        u0857(.A(men_men_n879_), .B(men_men_n160_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n876_), .B(men_men_n70_), .Y(men_men_n881_));
  NO2        u0859(.A(men_men_n174_), .B(i_0_), .Y(men_men_n882_));
  INV        u0860(.A(men_men_n882_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n475_), .B(men_men_n232_), .Y(men_men_n884_));
  AOI210     u0862(.A0(men_men_n376_), .A1(men_men_n41_), .B0(men_men_n412_), .Y(men_men_n885_));
  OAI220     u0863(.A0(men_men_n885_), .A1(men_men_n845_), .B0(men_men_n884_), .B1(men_men_n883_), .Y(men_men_n886_));
  NO3        u0864(.A(men_men_n886_), .B(men_men_n880_), .C(men_men_n878_), .Y(men_men_n887_));
  NA2        u0865(.A(men_men_n658_), .B(men_men_n120_), .Y(men_men_n888_));
  NO2        u0866(.A(i_6_), .B(men_men_n888_), .Y(men_men_n889_));
  AOI210     u0867(.A0(men_men_n453_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n890_));
  NA2        u0868(.A(men_men_n171_), .B(men_men_n101_), .Y(men_men_n891_));
  NOi32      u0869(.An(men_men_n890_), .Bn(men_men_n187_), .C(men_men_n891_), .Y(men_men_n892_));
  NA2        u0870(.A(men_men_n608_), .B(men_men_n334_), .Y(men_men_n893_));
  NO2        u0871(.A(men_men_n893_), .B(men_men_n836_), .Y(men_men_n894_));
  NO3        u0872(.A(men_men_n894_), .B(men_men_n892_), .C(men_men_n889_), .Y(men_men_n895_));
  NOi21      u0873(.An(i_7_), .B(i_5_), .Y(men_men_n896_));
  NOi31      u0874(.An(men_men_n896_), .B(i_0_), .C(men_men_n726_), .Y(men_men_n897_));
  NA3        u0875(.A(men_men_n897_), .B(men_men_n387_), .C(i_6_), .Y(men_men_n898_));
  OA210      u0876(.A0(men_men_n891_), .A1(men_men_n520_), .B0(men_men_n898_), .Y(men_men_n899_));
  NO3        u0877(.A(men_men_n408_), .B(men_men_n366_), .C(men_men_n362_), .Y(men_men_n900_));
  NO2        u0878(.A(men_men_n264_), .B(men_men_n323_), .Y(men_men_n901_));
  NO2        u0879(.A(men_men_n726_), .B(men_men_n259_), .Y(men_men_n902_));
  AOI210     u0880(.A0(men_men_n902_), .A1(men_men_n901_), .B0(men_men_n900_), .Y(men_men_n903_));
  NA4        u0881(.A(men_men_n903_), .B(men_men_n899_), .C(men_men_n895_), .D(men_men_n887_), .Y(men_men_n904_));
  NO2        u0882(.A(men_men_n851_), .B(men_men_n241_), .Y(men_men_n905_));
  AN2        u0883(.A(men_men_n339_), .B(men_men_n334_), .Y(men_men_n906_));
  NA2        u0884(.A(men_men_n905_), .B(i_10_), .Y(men_men_n907_));
  NO2        u0885(.A(men_men_n825_), .B(men_men_n322_), .Y(men_men_n908_));
  OA210      u0886(.A0(men_men_n475_), .A1(men_men_n224_), .B0(men_men_n474_), .Y(men_men_n909_));
  NA2        u0887(.A(men_men_n908_), .B(men_men_n881_), .Y(men_men_n910_));
  NA3        u0888(.A(men_men_n474_), .B(men_men_n415_), .C(men_men_n45_), .Y(men_men_n911_));
  OAI210     u0889(.A0(men_men_n855_), .A1(i_6_), .B0(men_men_n911_), .Y(men_men_n912_));
  NA2        u0890(.A(men_men_n881_), .B(men_men_n309_), .Y(men_men_n913_));
  NA2        u0891(.A(men_men_n186_), .B(men_men_n913_), .Y(men_men_n914_));
  AOI220     u0892(.A0(men_men_n914_), .A1(men_men_n475_), .B0(men_men_n912_), .B1(men_men_n70_), .Y(men_men_n915_));
  NO2        u0893(.A(men_men_n72_), .B(men_men_n744_), .Y(men_men_n916_));
  AOI210     u0894(.A0(men_men_n173_), .A1(men_men_n598_), .B0(men_men_n916_), .Y(men_men_n917_));
  NO2        u0895(.A(men_men_n917_), .B(men_men_n47_), .Y(men_men_n918_));
  NO3        u0896(.A(men_men_n589_), .B(men_men_n361_), .C(men_men_n24_), .Y(men_men_n919_));
  INV        u0897(.A(men_men_n919_), .Y(men_men_n920_));
  NAi21      u0898(.An(i_9_), .B(i_5_), .Y(men_men_n921_));
  NO2        u0899(.A(men_men_n921_), .B(men_men_n408_), .Y(men_men_n922_));
  NO2        u0900(.A(men_men_n604_), .B(men_men_n103_), .Y(men_men_n923_));
  AOI220     u0901(.A0(men_men_n923_), .A1(i_0_), .B0(men_men_n922_), .B1(men_men_n624_), .Y(men_men_n924_));
  OAI220     u0902(.A0(men_men_n924_), .A1(men_men_n82_), .B0(men_men_n920_), .B1(men_men_n172_), .Y(men_men_n925_));
  NO3        u0903(.A(men_men_n925_), .B(men_men_n918_), .C(men_men_n523_), .Y(men_men_n926_));
  NA4        u0904(.A(men_men_n926_), .B(men_men_n915_), .C(men_men_n910_), .D(men_men_n907_), .Y(men_men_n927_));
  NO3        u0905(.A(men_men_n927_), .B(men_men_n904_), .C(men_men_n874_), .Y(men_men_n928_));
  NO2        u0906(.A(i_0_), .B(men_men_n726_), .Y(men_men_n929_));
  NA2        u0907(.A(men_men_n70_), .B(men_men_n44_), .Y(men_men_n930_));
  NA2        u0908(.A(men_men_n865_), .B(men_men_n930_), .Y(men_men_n931_));
  NO2        u0909(.A(i_5_), .B(men_men_n25_), .Y(men_men_n932_));
  AO220      u0910(.A0(men_men_n932_), .A1(men_men_n931_), .B0(men_men_n929_), .B1(men_men_n173_), .Y(men_men_n933_));
  AOI210     u0911(.A0(men_men_n790_), .A1(men_men_n688_), .B0(men_men_n891_), .Y(men_men_n934_));
  AOI210     u0912(.A0(men_men_n933_), .A1(men_men_n351_), .B0(men_men_n934_), .Y(men_men_n935_));
  NA2        u0913(.A(men_men_n735_), .B(men_men_n145_), .Y(men_men_n936_));
  INV        u0914(.A(men_men_n936_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n937_), .B(men_men_n675_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n804_), .B(men_men_n408_), .Y(men_men_n939_));
  NA3        u0917(.A(men_men_n827_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n828_), .B(i_9_), .Y(men_men_n941_));
  AOI210     u0919(.A0(men_men_n940_), .A1(men_men_n502_), .B0(men_men_n941_), .Y(men_men_n942_));
  OAI210     u0920(.A0(men_men_n245_), .A1(i_9_), .B0(men_men_n231_), .Y(men_men_n943_));
  AOI210     u0921(.A0(men_men_n943_), .A1(men_men_n858_), .B0(men_men_n153_), .Y(men_men_n944_));
  NO3        u0922(.A(men_men_n944_), .B(men_men_n942_), .C(men_men_n939_), .Y(men_men_n945_));
  NA3        u0923(.A(men_men_n945_), .B(men_men_n938_), .C(men_men_n935_), .Y(men_men_n946_));
  NA2        u0924(.A(men_men_n906_), .B(men_men_n378_), .Y(men_men_n947_));
  AOI210     u0925(.A0(men_men_n304_), .A1(men_men_n162_), .B0(men_men_n947_), .Y(men_men_n948_));
  NA3        u0926(.A(men_men_n39_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n949_));
  NA2        u0927(.A(i_5_), .B(men_men_n490_), .Y(men_men_n950_));
  AOI210     u0928(.A0(men_men_n949_), .A1(men_men_n162_), .B0(men_men_n950_), .Y(men_men_n951_));
  NO2        u0929(.A(men_men_n951_), .B(men_men_n948_), .Y(men_men_n952_));
  NO3        u0930(.A(men_men_n865_), .B(men_men_n844_), .C(men_men_n189_), .Y(men_men_n953_));
  AOI220     u0931(.A0(men_men_n953_), .A1(i_11_), .B0(men_men_n570_), .B1(men_men_n72_), .Y(men_men_n954_));
  NO3        u0932(.A(men_men_n209_), .B(men_men_n386_), .C(i_0_), .Y(men_men_n955_));
  OAI210     u0933(.A0(men_men_n955_), .A1(men_men_n73_), .B0(i_13_), .Y(men_men_n956_));
  OAI220     u0934(.A0(men_men_n532_), .A1(men_men_n138_), .B0(i_12_), .B1(men_men_n618_), .Y(men_men_n957_));
  NA3        u0935(.A(men_men_n957_), .B(men_men_n400_), .C(i_0_), .Y(men_men_n958_));
  NA4        u0936(.A(men_men_n958_), .B(men_men_n956_), .C(men_men_n954_), .D(men_men_n952_), .Y(men_men_n959_));
  NO2        u0937(.A(men_men_n244_), .B(men_men_n90_), .Y(men_men_n960_));
  AOI210     u0938(.A0(men_men_n960_), .A1(men_men_n929_), .B0(men_men_n107_), .Y(men_men_n961_));
  AOI220     u0939(.A0(men_men_n896_), .A1(men_men_n490_), .B0(men_men_n827_), .B1(men_men_n163_), .Y(men_men_n962_));
  NA2        u0940(.A(men_men_n354_), .B(men_men_n175_), .Y(men_men_n963_));
  OA220      u0941(.A0(men_men_n963_), .A1(men_men_n962_), .B0(men_men_n961_), .B1(i_5_), .Y(men_men_n964_));
  AOI210     u0942(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n174_), .Y(men_men_n965_));
  NA2        u0943(.A(men_men_n965_), .B(men_men_n909_), .Y(men_men_n966_));
  NA3        u0944(.A(men_men_n495_), .B(men_men_n488_), .C(men_men_n472_), .Y(men_men_n967_));
  INV        u0945(.A(men_men_n967_), .Y(men_men_n968_));
  NA3        u0946(.A(men_men_n393_), .B(men_men_n171_), .C(men_men_n170_), .Y(men_men_n969_));
  NA3        u0947(.A(i_5_), .B(men_men_n293_), .C(men_men_n231_), .Y(men_men_n970_));
  NA2        u0948(.A(men_men_n970_), .B(men_men_n969_), .Y(men_men_n971_));
  NA3        u0949(.A(men_men_n393_), .B(men_men_n341_), .C(men_men_n222_), .Y(men_men_n972_));
  INV        u0950(.A(men_men_n972_), .Y(men_men_n973_));
  NOi31      u0951(.An(men_men_n392_), .B(men_men_n930_), .C(men_men_n241_), .Y(men_men_n974_));
  NO3        u0952(.A(men_men_n974_), .B(men_men_n973_), .C(men_men_n971_), .Y(men_men_n975_));
  NA4        u0953(.A(men_men_n975_), .B(men_men_n968_), .C(men_men_n966_), .D(men_men_n964_), .Y(men_men_n976_));
  NO2        u0954(.A(men_men_n82_), .B(i_5_), .Y(men_men_n977_));
  NA3        u0955(.A(men_men_n828_), .B(men_men_n108_), .C(men_men_n123_), .Y(men_men_n978_));
  INV        u0956(.A(men_men_n978_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n979_), .B(men_men_n977_), .Y(men_men_n980_));
  NA3        u0958(.A(men_men_n309_), .B(i_5_), .C(men_men_n192_), .Y(men_men_n981_));
  NO3        u0959(.A(men_men_n241_), .B(i_0_), .C(i_12_), .Y(men_men_n982_));
  AOI220     u0960(.A0(men_men_n982_), .A1(men_men_n243_), .B0(men_men_n784_), .B1(men_men_n175_), .Y(men_men_n983_));
  AN2        u0961(.A(men_men_n865_), .B(men_men_n153_), .Y(men_men_n984_));
  NO3        u0962(.A(men_men_n984_), .B(i_12_), .C(men_men_n646_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n985_), .B(men_men_n218_), .Y(men_men_n986_));
  NA3        u0964(.A(men_men_n96_), .B(men_men_n574_), .C(i_11_), .Y(men_men_n987_));
  NO2        u0965(.A(men_men_n987_), .B(men_men_n155_), .Y(men_men_n988_));
  NA2        u0966(.A(men_men_n896_), .B(men_men_n471_), .Y(men_men_n989_));
  INV        u0967(.A(men_men_n64_), .Y(men_men_n990_));
  OAI220     u0968(.A0(men_men_n990_), .A1(men_men_n981_), .B0(men_men_n989_), .B1(men_men_n676_), .Y(men_men_n991_));
  AOI210     u0969(.A0(men_men_n991_), .A1(men_men_n882_), .B0(men_men_n988_), .Y(men_men_n992_));
  NA4        u0970(.A(men_men_n992_), .B(men_men_n986_), .C(men_men_n983_), .D(men_men_n980_), .Y(men_men_n993_));
  NO4        u0971(.A(men_men_n993_), .B(men_men_n976_), .C(men_men_n959_), .D(men_men_n946_), .Y(men_men_n994_));
  NA3        u0972(.A(men_men_n890_), .B(men_men_n373_), .C(i_5_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n995_), .B(men_men_n613_), .Y(men_men_n996_));
  NA2        u0974(.A(men_men_n996_), .B(men_men_n207_), .Y(men_men_n997_));
  AN2        u0975(.A(men_men_n701_), .B(men_men_n374_), .Y(men_men_n998_));
  NA2        u0976(.A(men_men_n185_), .B(men_men_n187_), .Y(men_men_n999_));
  AO210      u0977(.A0(men_men_n998_), .A1(men_men_n33_), .B0(men_men_n999_), .Y(men_men_n1000_));
  OAI210     u0978(.A0(men_men_n617_), .A1(men_men_n615_), .B0(men_men_n322_), .Y(men_men_n1001_));
  NA2        u0979(.A(men_men_n1001_), .B(men_men_n1000_), .Y(men_men_n1002_));
  NO2        u0980(.A(men_men_n465_), .B(men_men_n270_), .Y(men_men_n1003_));
  NO4        u0981(.A(men_men_n234_), .B(men_men_n144_), .C(men_men_n679_), .D(men_men_n37_), .Y(men_men_n1004_));
  NO3        u0982(.A(men_men_n1004_), .B(men_men_n1003_), .C(men_men_n860_), .Y(men_men_n1005_));
  OAI210     u0983(.A0(men_men_n987_), .A1(men_men_n147_), .B0(men_men_n1005_), .Y(men_men_n1006_));
  AOI210     u0984(.A0(men_men_n1002_), .A1(men_men_n48_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  AOI210     u0985(.A0(men_men_n1007_), .A1(men_men_n997_), .B0(men_men_n70_), .Y(men_men_n1008_));
  INV        u0986(.A(men_men_n567_), .Y(men_men_n1009_));
  NO2        u0987(.A(men_men_n1009_), .B(men_men_n750_), .Y(men_men_n1010_));
  INV        u0988(.A(men_men_n73_), .Y(men_men_n1011_));
  AOI210     u0989(.A0(men_men_n965_), .A1(i_5_), .B0(men_men_n897_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n1012_), .A1(men_men_n1011_), .B0(men_men_n679_), .Y(men_men_n1013_));
  NA2        u0991(.A(i_8_), .B(men_men_n73_), .Y(men_men_n1014_));
  NO2        u0992(.A(men_men_n1014_), .B(men_men_n238_), .Y(men_men_n1015_));
  NA3        u0993(.A(men_men_n94_), .B(men_men_n311_), .C(men_men_n31_), .Y(men_men_n1016_));
  INV        u0994(.A(men_men_n1016_), .Y(men_men_n1017_));
  NO3        u0995(.A(men_men_n1017_), .B(men_men_n1015_), .C(men_men_n1013_), .Y(men_men_n1018_));
  OAI210     u0996(.A0(men_men_n272_), .A1(men_men_n158_), .B0(men_men_n85_), .Y(men_men_n1019_));
  NA3        u0997(.A(men_men_n754_), .B(men_men_n293_), .C(men_men_n77_), .Y(men_men_n1020_));
  AOI210     u0998(.A0(men_men_n1020_), .A1(men_men_n1019_), .B0(i_11_), .Y(men_men_n1021_));
  NA2        u0999(.A(men_men_n609_), .B(men_men_n215_), .Y(men_men_n1022_));
  OAI210     u1000(.A0(men_men_n1022_), .A1(men_men_n890_), .B0(men_men_n207_), .Y(men_men_n1023_));
  NA2        u1001(.A(men_men_n164_), .B(i_5_), .Y(men_men_n1024_));
  AOI210     u1002(.A0(men_men_n1023_), .A1(men_men_n764_), .B0(men_men_n1024_), .Y(men_men_n1025_));
  NO3        u1003(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1026_));
  OAI210     u1004(.A0(men_men_n901_), .A1(men_men_n311_), .B0(men_men_n1026_), .Y(men_men_n1027_));
  NO2        u1005(.A(men_men_n1027_), .B(men_men_n726_), .Y(men_men_n1028_));
  NO4        u1006(.A(men_men_n921_), .B(men_men_n478_), .C(men_men_n254_), .D(men_men_n253_), .Y(men_men_n1029_));
  NO2        u1007(.A(men_men_n1029_), .B(men_men_n564_), .Y(men_men_n1030_));
  INV        u1008(.A(men_men_n367_), .Y(men_men_n1031_));
  AOI210     u1009(.A0(men_men_n1031_), .A1(men_men_n1030_), .B0(men_men_n40_), .Y(men_men_n1032_));
  NO4        u1010(.A(men_men_n1032_), .B(men_men_n1028_), .C(men_men_n1025_), .D(men_men_n1021_), .Y(men_men_n1033_));
  OAI210     u1011(.A0(men_men_n1018_), .A1(i_4_), .B0(men_men_n1033_), .Y(men_men_n1034_));
  NO3        u1012(.A(men_men_n1034_), .B(men_men_n1010_), .C(men_men_n1008_), .Y(men_men_n1035_));
  NA4        u1013(.A(men_men_n1035_), .B(men_men_n994_), .C(men_men_n928_), .D(men_men_n850_), .Y(men4));
  INV        u1014(.A(i_2_), .Y(men_men_n1039_));
  INV        u1015(.A(i_9_), .Y(men_men_n1040_));
  INV        u1016(.A(men_men_n741_), .Y(men_men_n1041_));
  INV        u1017(.A(i_6_), .Y(men_men_n1042_));
  INV        u1018(.A(i_10_), .Y(men_men_n1043_));
  INV        u1019(.A(i_9_), .Y(men_men_n1044_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule