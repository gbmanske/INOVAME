//Benchmark atmr_max1024_476_0.0625

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n411_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  INV        o012(.A(ori_ori_n24_), .Y(ori_ori_n29_));
  NO2        o013(.A(x4), .B(x3), .Y(ori_ori_n30_));
  INV        o014(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  OA210      o015(.A0(ori_ori_n31_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n32_));
  NOi31      o016(.An(ori_ori_n23_), .B(ori_ori_n32_), .C(ori_ori_n29_), .Y(ori00));
  NO2        o017(.A(x1), .B(x0), .Y(ori_ori_n34_));
  INV        o018(.A(x6), .Y(ori_ori_n35_));
  NO2        o019(.A(ori_ori_n35_), .B(ori_ori_n25_), .Y(ori_ori_n36_));
  AN2        o020(.A(x8), .B(x7), .Y(ori_ori_n37_));
  NA2        o021(.A(x4), .B(x3), .Y(ori_ori_n38_));
  NO2        o022(.A(ori_ori_n23_), .B(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o023(.A(x2), .B(x0), .Y(ori_ori_n40_));
  INV        o024(.A(x3), .Y(ori_ori_n41_));
  NO2        o025(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n42_));
  INV        o026(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n36_), .B(x4), .Y(ori_ori_n44_));
  OAI210     o028(.A0(ori_ori_n44_), .A1(ori_ori_n43_), .B0(ori_ori_n40_), .Y(ori_ori_n45_));
  INV        o029(.A(x4), .Y(ori_ori_n46_));
  NO2        o030(.A(ori_ori_n46_), .B(ori_ori_n17_), .Y(ori_ori_n47_));
  NA2        o031(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n48_));
  OAI210     o032(.A0(ori_ori_n48_), .A1(ori_ori_n20_), .B0(ori_ori_n45_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n50_));
  AOI220     o034(.A0(ori_ori_n50_), .A1(ori_ori_n34_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n51_));
  INV        o035(.A(x2), .Y(ori_ori_n52_));
  NO2        o036(.A(ori_ori_n52_), .B(ori_ori_n17_), .Y(ori_ori_n53_));
  NA2        o037(.A(ori_ori_n41_), .B(ori_ori_n18_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  OAI210     o039(.A0(ori_ori_n51_), .A1(ori_ori_n31_), .B0(ori_ori_n55_), .Y(ori_ori_n56_));
  NO3        o040(.A(ori_ori_n56_), .B(ori_ori_n49_), .C(ori_ori_n39_), .Y(ori01));
  NA2        o041(.A(x8), .B(x7), .Y(ori_ori_n58_));
  NA2        o042(.A(ori_ori_n41_), .B(x1), .Y(ori_ori_n59_));
  INV        o043(.A(x9), .Y(ori_ori_n60_));
  NO2        o044(.A(x7), .B(x6), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n59_), .B(x5), .Y(ori_ori_n62_));
  AN2        o046(.A(ori_ori_n62_), .B(ori_ori_n61_), .Y(ori_ori_n63_));
  OAI210     o047(.A0(ori_ori_n42_), .A1(ori_ori_n25_), .B0(ori_ori_n52_), .Y(ori_ori_n64_));
  OAI210     o048(.A0(ori_ori_n54_), .A1(ori_ori_n20_), .B0(ori_ori_n64_), .Y(ori_ori_n65_));
  NO2        o049(.A(ori_ori_n65_), .B(ori_ori_n63_), .Y(ori_ori_n66_));
  NA2        o050(.A(ori_ori_n66_), .B(x4), .Y(ori_ori_n67_));
  NA2        o051(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n68_));
  OAI210     o052(.A0(ori_ori_n68_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n69_));
  NA2        o053(.A(x5), .B(x3), .Y(ori_ori_n70_));
  NO2        o054(.A(x8), .B(x6), .Y(ori_ori_n71_));
  NO4        o055(.A(ori_ori_n71_), .B(ori_ori_n70_), .C(ori_ori_n61_), .D(ori_ori_n52_), .Y(ori_ori_n72_));
  NAi21      o056(.An(x4), .B(x3), .Y(ori_ori_n73_));
  INV        o057(.A(ori_ori_n73_), .Y(ori_ori_n74_));
  NO2        o058(.A(ori_ori_n74_), .B(ori_ori_n22_), .Y(ori_ori_n75_));
  NO2        o059(.A(x4), .B(x2), .Y(ori_ori_n76_));
  NO2        o060(.A(ori_ori_n76_), .B(x3), .Y(ori_ori_n77_));
  NO3        o061(.A(ori_ori_n77_), .B(ori_ori_n75_), .C(ori_ori_n18_), .Y(ori_ori_n78_));
  NO3        o062(.A(ori_ori_n78_), .B(ori_ori_n72_), .C(ori_ori_n69_), .Y(ori_ori_n79_));
  NA2        o063(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n80_));
  NO2        o064(.A(ori_ori_n80_), .B(ori_ori_n25_), .Y(ori_ori_n81_));
  INV        o065(.A(x8), .Y(ori_ori_n82_));
  NA2        o066(.A(x2), .B(x1), .Y(ori_ori_n83_));
  INV        o067(.A(ori_ori_n81_), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n84_), .B(ori_ori_n26_), .Y(ori_ori_n85_));
  AOI210     o069(.A0(ori_ori_n54_), .A1(ori_ori_n25_), .B0(ori_ori_n52_), .Y(ori_ori_n86_));
  OAI210     o070(.A0(ori_ori_n43_), .A1(ori_ori_n36_), .B0(ori_ori_n46_), .Y(ori_ori_n87_));
  NO3        o071(.A(ori_ori_n87_), .B(ori_ori_n86_), .C(ori_ori_n85_), .Y(ori_ori_n88_));
  NA2        o072(.A(x4), .B(ori_ori_n41_), .Y(ori_ori_n89_));
  NO2        o073(.A(ori_ori_n46_), .B(ori_ori_n52_), .Y(ori_ori_n90_));
  OAI210     o074(.A0(ori_ori_n90_), .A1(ori_ori_n41_), .B0(ori_ori_n18_), .Y(ori_ori_n91_));
  AOI210     o075(.A0(ori_ori_n89_), .A1(ori_ori_n50_), .B0(ori_ori_n91_), .Y(ori_ori_n92_));
  NO2        o076(.A(x3), .B(x2), .Y(ori_ori_n93_));
  NA3        o077(.A(ori_ori_n93_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n94_));
  AOI210     o078(.A0(x8), .A1(x6), .B0(ori_ori_n94_), .Y(ori_ori_n95_));
  NA2        o079(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n96_));
  OAI210     o080(.A0(ori_ori_n96_), .A1(ori_ori_n38_), .B0(ori_ori_n17_), .Y(ori_ori_n97_));
  NO4        o081(.A(ori_ori_n97_), .B(ori_ori_n95_), .C(ori_ori_n92_), .D(ori_ori_n88_), .Y(ori_ori_n98_));
  AO210      o082(.A0(ori_ori_n79_), .A1(ori_ori_n67_), .B0(ori_ori_n98_), .Y(ori02));
  NO2        o083(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n100_));
  NO2        o084(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n101_));
  NA2        o085(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n102_));
  INV        o086(.A(ori_ori_n102_), .Y(ori_ori_n103_));
  AOI220     o087(.A0(ori_ori_n103_), .A1(ori_ori_n101_), .B0(ori_ori_n100_), .B1(x4), .Y(ori_ori_n104_));
  NO3        o088(.A(ori_ori_n104_), .B(x7), .C(x5), .Y(ori_ori_n105_));
  OR2        o089(.A(x8), .B(x0), .Y(ori_ori_n106_));
  INV        o090(.A(ori_ori_n106_), .Y(ori_ori_n107_));
  NO2        o091(.A(x4), .B(x1), .Y(ori_ori_n108_));
  NA3        o092(.A(ori_ori_n108_), .B(x2), .C(ori_ori_n58_), .Y(ori_ori_n109_));
  NOi21      o093(.An(x0), .B(x1), .Y(ori_ori_n110_));
  NOi21      o094(.An(x0), .B(x4), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n109_), .B(ori_ori_n70_), .Y(ori_ori_n112_));
  NO2        o096(.A(x5), .B(ori_ori_n46_), .Y(ori_ori_n113_));
  NA2        o097(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n114_));
  AOI210     o098(.A0(ori_ori_n114_), .A1(ori_ori_n96_), .B0(ori_ori_n102_), .Y(ori_ori_n115_));
  OAI210     o099(.A0(ori_ori_n115_), .A1(ori_ori_n34_), .B0(ori_ori_n113_), .Y(ori_ori_n116_));
  NAi21      o100(.An(x0), .B(x4), .Y(ori_ori_n117_));
  NO2        o101(.A(ori_ori_n117_), .B(x1), .Y(ori_ori_n118_));
  NO2        o102(.A(x7), .B(x0), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n76_), .B(ori_ori_n90_), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n120_), .B(x3), .Y(ori_ori_n121_));
  OAI210     o105(.A0(ori_ori_n119_), .A1(ori_ori_n118_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n21_), .B(ori_ori_n41_), .Y(ori_ori_n123_));
  NA2        o107(.A(x5), .B(x0), .Y(ori_ori_n124_));
  NO2        o108(.A(ori_ori_n46_), .B(x2), .Y(ori_ori_n125_));
  NA3        o109(.A(ori_ori_n125_), .B(ori_ori_n124_), .C(ori_ori_n123_), .Y(ori_ori_n126_));
  NA4        o110(.A(ori_ori_n126_), .B(ori_ori_n122_), .C(ori_ori_n116_), .D(ori_ori_n35_), .Y(ori_ori_n127_));
  NO3        o111(.A(ori_ori_n127_), .B(ori_ori_n112_), .C(ori_ori_n105_), .Y(ori_ori_n128_));
  NO3        o112(.A(ori_ori_n70_), .B(ori_ori_n68_), .C(ori_ori_n24_), .Y(ori_ori_n129_));
  NO2        o113(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n130_));
  NA2        o114(.A(x7), .B(x3), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n89_), .B(x5), .Y(ori_ori_n132_));
  NO2        o116(.A(x9), .B(x7), .Y(ori_ori_n133_));
  NOi21      o117(.An(x8), .B(x0), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n41_), .B(x2), .Y(ori_ori_n135_));
  INV        o119(.A(x7), .Y(ori_ori_n136_));
  NA2        o120(.A(ori_ori_n136_), .B(ori_ori_n18_), .Y(ori_ori_n137_));
  AOI220     o121(.A0(ori_ori_n137_), .A1(ori_ori_n135_), .B0(ori_ori_n100_), .B1(ori_ori_n37_), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n139_), .B(ori_ori_n111_), .Y(ori_ori_n140_));
  NO2        o124(.A(ori_ori_n140_), .B(ori_ori_n138_), .Y(ori_ori_n141_));
  INV        o125(.A(ori_ori_n141_), .Y(ori_ori_n142_));
  OAI210     o126(.A0(ori_ori_n131_), .A1(ori_ori_n48_), .B0(ori_ori_n142_), .Y(ori_ori_n143_));
  NA2        o127(.A(x5), .B(x1), .Y(ori_ori_n144_));
  INV        o128(.A(ori_ori_n144_), .Y(ori_ori_n145_));
  AOI210     o129(.A0(ori_ori_n145_), .A1(ori_ori_n111_), .B0(ori_ori_n35_), .Y(ori_ori_n146_));
  NAi21      o130(.An(x2), .B(x7), .Y(ori_ori_n147_));
  NO2        o131(.A(ori_ori_n147_), .B(ori_ori_n46_), .Y(ori_ori_n148_));
  NA2        o132(.A(ori_ori_n148_), .B(ori_ori_n62_), .Y(ori_ori_n149_));
  NA2        o133(.A(ori_ori_n149_), .B(ori_ori_n146_), .Y(ori_ori_n150_));
  NO3        o134(.A(ori_ori_n150_), .B(ori_ori_n143_), .C(ori_ori_n129_), .Y(ori_ori_n151_));
  NO2        o135(.A(ori_ori_n151_), .B(ori_ori_n128_), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n124_), .B(ori_ori_n120_), .Y(ori_ori_n153_));
  NA2        o137(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n154_));
  NA2        o138(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n155_));
  NA3        o139(.A(ori_ori_n155_), .B(ori_ori_n154_), .C(ori_ori_n24_), .Y(ori_ori_n156_));
  AN2        o140(.A(ori_ori_n156_), .B(ori_ori_n125_), .Y(ori_ori_n157_));
  NA2        o141(.A(x8), .B(x0), .Y(ori_ori_n158_));
  NO2        o142(.A(ori_ori_n136_), .B(ori_ori_n25_), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n110_), .B(x4), .Y(ori_ori_n160_));
  NA2        o144(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  AOI210     o145(.A0(ori_ori_n158_), .A1(ori_ori_n114_), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  NA2        o146(.A(x2), .B(x0), .Y(ori_ori_n163_));
  NA2        o147(.A(x4), .B(x1), .Y(ori_ori_n164_));
  NAi21      o148(.An(ori_ori_n108_), .B(ori_ori_n164_), .Y(ori_ori_n165_));
  NOi31      o149(.An(ori_ori_n165_), .B(ori_ori_n139_), .C(ori_ori_n163_), .Y(ori_ori_n166_));
  NO4        o150(.A(ori_ori_n166_), .B(ori_ori_n162_), .C(ori_ori_n157_), .D(ori_ori_n153_), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n167_), .B(ori_ori_n41_), .Y(ori_ori_n168_));
  NO2        o152(.A(ori_ori_n156_), .B(ori_ori_n68_), .Y(ori_ori_n169_));
  INV        o153(.A(ori_ori_n113_), .Y(ori_ori_n170_));
  NO2        o154(.A(ori_ori_n96_), .B(ori_ori_n17_), .Y(ori_ori_n171_));
  AOI210     o155(.A0(ori_ori_n34_), .A1(ori_ori_n82_), .B0(ori_ori_n171_), .Y(ori_ori_n172_));
  NO3        o156(.A(ori_ori_n172_), .B(ori_ori_n170_), .C(x7), .Y(ori_ori_n173_));
  NA3        o157(.A(ori_ori_n165_), .B(ori_ori_n170_), .C(ori_ori_n40_), .Y(ori_ori_n174_));
  OAI210     o158(.A0(ori_ori_n155_), .A1(ori_ori_n120_), .B0(ori_ori_n174_), .Y(ori_ori_n175_));
  NO3        o159(.A(ori_ori_n175_), .B(ori_ori_n173_), .C(ori_ori_n169_), .Y(ori_ori_n176_));
  NO2        o160(.A(ori_ori_n176_), .B(x3), .Y(ori_ori_n177_));
  NO3        o161(.A(ori_ori_n177_), .B(ori_ori_n168_), .C(ori_ori_n152_), .Y(ori03));
  NO2        o162(.A(ori_ori_n46_), .B(x3), .Y(ori_ori_n179_));
  NO2        o163(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n180_));
  NO2        o164(.A(ori_ori_n52_), .B(x1), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n70_), .B(x6), .Y(ori_ori_n182_));
  NA2        o166(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n183_), .B(x4), .Y(ori_ori_n184_));
  NO2        o168(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n185_));
  AO220      o169(.A0(ori_ori_n185_), .A1(ori_ori_n184_), .B0(ori_ori_n182_), .B1(ori_ori_n53_), .Y(ori_ori_n186_));
  INV        o170(.A(ori_ori_n186_), .Y(ori_ori_n187_));
  NA2        o171(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n188_));
  NA2        o172(.A(x9), .B(ori_ori_n52_), .Y(ori_ori_n189_));
  NA2        o173(.A(ori_ori_n183_), .B(ori_ori_n73_), .Y(ori_ori_n190_));
  AOI210     o174(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n163_), .Y(ori_ori_n191_));
  NA2        o175(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n192_));
  NO3        o176(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n193_));
  NO2        o177(.A(x5), .B(x1), .Y(ori_ori_n194_));
  NO2        o178(.A(ori_ori_n188_), .B(ori_ori_n154_), .Y(ori_ori_n195_));
  NO3        o179(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n196_));
  NO2        o180(.A(ori_ori_n196_), .B(ori_ori_n195_), .Y(ori_ori_n197_));
  INV        o181(.A(ori_ori_n197_), .Y(ori_ori_n198_));
  NA2        o182(.A(ori_ori_n198_), .B(ori_ori_n46_), .Y(ori_ori_n199_));
  NA3        o183(.A(ori_ori_n199_), .B(ori_ori_n192_), .C(ori_ori_n187_), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n46_), .B(ori_ori_n41_), .Y(ori_ori_n201_));
  NA2        o185(.A(ori_ori_n201_), .B(ori_ori_n19_), .Y(ori_ori_n202_));
  NO2        o186(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n203_), .B(x6), .Y(ori_ori_n204_));
  NOi21      o188(.An(ori_ori_n76_), .B(ori_ori_n204_), .Y(ori_ori_n205_));
  NA2        o189(.A(ori_ori_n60_), .B(ori_ori_n82_), .Y(ori_ori_n206_));
  NA3        o190(.A(ori_ori_n206_), .B(ori_ori_n203_), .C(x6), .Y(ori_ori_n207_));
  AOI210     o191(.A0(ori_ori_n207_), .A1(ori_ori_n205_), .B0(ori_ori_n136_), .Y(ori_ori_n208_));
  AO210      o192(.A0(ori_ori_n208_), .A1(ori_ori_n202_), .B0(ori_ori_n159_), .Y(ori_ori_n209_));
  NA2        o193(.A(ori_ori_n41_), .B(ori_ori_n52_), .Y(ori_ori_n210_));
  OAI210     o194(.A0(ori_ori_n210_), .A1(ori_ori_n25_), .B0(ori_ori_n155_), .Y(ori_ori_n211_));
  NO2        o195(.A(ori_ori_n164_), .B(x6), .Y(ori_ori_n212_));
  AOI220     o196(.A0(ori_ori_n212_), .A1(ori_ori_n211_), .B0(ori_ori_n125_), .B1(ori_ori_n81_), .Y(ori_ori_n213_));
  NA2        o197(.A(x6), .B(ori_ori_n46_), .Y(ori_ori_n214_));
  OAI210     o198(.A0(ori_ori_n107_), .A1(ori_ori_n71_), .B0(x4), .Y(ori_ori_n215_));
  AOI210     o199(.A0(ori_ori_n215_), .A1(ori_ori_n214_), .B0(ori_ori_n70_), .Y(ori_ori_n216_));
  NA2        o200(.A(ori_ori_n180_), .B(ori_ori_n118_), .Y(ori_ori_n217_));
  NA3        o201(.A(ori_ori_n188_), .B(ori_ori_n113_), .C(x6), .Y(ori_ori_n218_));
  OAI210     o202(.A0(ori_ori_n82_), .A1(ori_ori_n35_), .B0(ori_ori_n62_), .Y(ori_ori_n219_));
  NA3        o203(.A(ori_ori_n219_), .B(ori_ori_n218_), .C(ori_ori_n217_), .Y(ori_ori_n220_));
  OAI210     o204(.A0(ori_ori_n220_), .A1(ori_ori_n216_), .B0(x2), .Y(ori_ori_n221_));
  NA3        o205(.A(ori_ori_n221_), .B(ori_ori_n213_), .C(ori_ori_n209_), .Y(ori_ori_n222_));
  AOI210     o206(.A0(ori_ori_n200_), .A1(x8), .B0(ori_ori_n222_), .Y(ori_ori_n223_));
  NO2        o207(.A(ori_ori_n82_), .B(x3), .Y(ori_ori_n224_));
  NA2        o208(.A(ori_ori_n224_), .B(ori_ori_n184_), .Y(ori_ori_n225_));
  NO2        o209(.A(ori_ori_n80_), .B(ori_ori_n25_), .Y(ori_ori_n226_));
  AOI210     o210(.A0(ori_ori_n204_), .A1(ori_ori_n139_), .B0(ori_ori_n226_), .Y(ori_ori_n227_));
  AOI210     o211(.A0(ori_ori_n227_), .A1(ori_ori_n225_), .B0(x2), .Y(ori_ori_n228_));
  NO2        o212(.A(x4), .B(ori_ori_n52_), .Y(ori_ori_n229_));
  AOI220     o213(.A0(ori_ori_n184_), .A1(ori_ori_n171_), .B0(ori_ori_n229_), .B1(ori_ori_n62_), .Y(ori_ori_n230_));
  NA2        o214(.A(ori_ori_n41_), .B(ori_ori_n17_), .Y(ori_ori_n231_));
  NO2        o215(.A(ori_ori_n231_), .B(ori_ori_n25_), .Y(ori_ori_n232_));
  NA2        o216(.A(ori_ori_n232_), .B(ori_ori_n108_), .Y(ori_ori_n233_));
  NA2        o217(.A(ori_ori_n188_), .B(x6), .Y(ori_ori_n234_));
  NO2        o218(.A(ori_ori_n188_), .B(x6), .Y(ori_ori_n235_));
  INV        o219(.A(ori_ori_n235_), .Y(ori_ori_n236_));
  NA3        o220(.A(ori_ori_n236_), .B(ori_ori_n234_), .C(ori_ori_n130_), .Y(ori_ori_n237_));
  NA4        o221(.A(ori_ori_n237_), .B(ori_ori_n233_), .C(ori_ori_n230_), .D(ori_ori_n136_), .Y(ori_ori_n238_));
  NA2        o222(.A(ori_ori_n180_), .B(ori_ori_n203_), .Y(ori_ori_n239_));
  NAi21      o223(.An(x1), .B(x4), .Y(ori_ori_n240_));
  AOI210     o224(.A0(x3), .A1(x2), .B0(ori_ori_n46_), .Y(ori_ori_n241_));
  OAI210     o225(.A0(ori_ori_n124_), .A1(x3), .B0(ori_ori_n241_), .Y(ori_ori_n242_));
  NA2        o226(.A(ori_ori_n242_), .B(ori_ori_n240_), .Y(ori_ori_n243_));
  NA2        o227(.A(ori_ori_n243_), .B(ori_ori_n239_), .Y(ori_ori_n244_));
  NA2        o228(.A(ori_ori_n60_), .B(x2), .Y(ori_ori_n245_));
  NA2        o229(.A(x6), .B(x2), .Y(ori_ori_n246_));
  NO2        o230(.A(ori_ori_n160_), .B(ori_ori_n44_), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n247_), .B(ori_ori_n244_), .Y(ori_ori_n248_));
  OR2        o232(.A(ori_ori_n182_), .B(ori_ori_n132_), .Y(ori_ori_n249_));
  NA2        o233(.A(x4), .B(x0), .Y(ori_ori_n250_));
  NA2        o234(.A(ori_ori_n249_), .B(ori_ori_n40_), .Y(ori_ori_n251_));
  AOI210     o235(.A0(ori_ori_n251_), .A1(ori_ori_n248_), .B0(x8), .Y(ori_ori_n252_));
  INV        o236(.A(ori_ori_n158_), .Y(ori_ori_n253_));
  OAI210     o237(.A0(ori_ori_n253_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n254_));
  NO2        o238(.A(ori_ori_n254_), .B(ori_ori_n210_), .Y(ori_ori_n255_));
  NO4        o239(.A(ori_ori_n255_), .B(ori_ori_n252_), .C(ori_ori_n238_), .D(ori_ori_n228_), .Y(ori_ori_n256_));
  INV        o240(.A(x1), .Y(ori_ori_n257_));
  NO3        o241(.A(ori_ori_n257_), .B(x3), .C(ori_ori_n35_), .Y(ori_ori_n258_));
  OAI210     o242(.A0(ori_ori_n258_), .A1(ori_ori_n235_), .B0(x2), .Y(ori_ori_n259_));
  OAI210     o243(.A0(ori_ori_n253_), .A1(x6), .B0(ori_ori_n42_), .Y(ori_ori_n260_));
  AOI210     o244(.A0(ori_ori_n260_), .A1(ori_ori_n259_), .B0(ori_ori_n170_), .Y(ori_ori_n261_));
  NOi21      o245(.An(ori_ori_n246_), .B(ori_ori_n17_), .Y(ori_ori_n262_));
  NA3        o246(.A(ori_ori_n262_), .B(ori_ori_n194_), .C(ori_ori_n38_), .Y(ori_ori_n263_));
  AOI210     o247(.A0(ori_ori_n35_), .A1(ori_ori_n52_), .B0(x0), .Y(ori_ori_n264_));
  NA3        o248(.A(ori_ori_n264_), .B(ori_ori_n145_), .C(ori_ori_n31_), .Y(ori_ori_n265_));
  NA2        o249(.A(x3), .B(x2), .Y(ori_ori_n266_));
  AOI220     o250(.A0(ori_ori_n266_), .A1(ori_ori_n210_), .B0(ori_ori_n265_), .B1(ori_ori_n263_), .Y(ori_ori_n267_));
  NAi21      o251(.An(x4), .B(x0), .Y(ori_ori_n268_));
  NO3        o252(.A(ori_ori_n268_), .B(ori_ori_n42_), .C(x2), .Y(ori_ori_n269_));
  OAI210     o253(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n269_), .Y(ori_ori_n270_));
  OAI220     o254(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n271_));
  NO2        o255(.A(ori_ori_n264_), .B(ori_ori_n262_), .Y(ori_ori_n272_));
  AOI220     o256(.A0(ori_ori_n272_), .A1(ori_ori_n74_), .B0(ori_ori_n271_), .B1(ori_ori_n30_), .Y(ori_ori_n273_));
  AOI210     o257(.A0(ori_ori_n273_), .A1(ori_ori_n270_), .B0(ori_ori_n25_), .Y(ori_ori_n274_));
  NA3        o258(.A(ori_ori_n35_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n275_));
  OAI210     o259(.A0(ori_ori_n264_), .A1(ori_ori_n262_), .B0(ori_ori_n275_), .Y(ori_ori_n276_));
  INV        o260(.A(ori_ori_n195_), .Y(ori_ori_n277_));
  NA2        o261(.A(ori_ori_n35_), .B(ori_ori_n41_), .Y(ori_ori_n278_));
  OR2        o262(.A(ori_ori_n278_), .B(ori_ori_n250_), .Y(ori_ori_n279_));
  OAI220     o263(.A0(ori_ori_n279_), .A1(ori_ori_n144_), .B0(ori_ori_n214_), .B1(ori_ori_n277_), .Y(ori_ori_n280_));
  AO210      o264(.A0(ori_ori_n276_), .A1(ori_ori_n132_), .B0(ori_ori_n280_), .Y(ori_ori_n281_));
  NO4        o265(.A(ori_ori_n281_), .B(ori_ori_n274_), .C(ori_ori_n267_), .D(ori_ori_n261_), .Y(ori_ori_n282_));
  OAI210     o266(.A0(ori_ori_n256_), .A1(ori_ori_n223_), .B0(ori_ori_n282_), .Y(ori04));
  NO2        o267(.A(x2), .B(x1), .Y(ori_ori_n284_));
  OAI210     o268(.A0(ori_ori_n231_), .A1(ori_ori_n284_), .B0(ori_ori_n35_), .Y(ori_ori_n285_));
  NO2        o269(.A(ori_ori_n284_), .B(ori_ori_n268_), .Y(ori_ori_n286_));
  OAI210     o270(.A0(ori_ori_n52_), .A1(ori_ori_n286_), .B0(ori_ori_n224_), .Y(ori_ori_n287_));
  NO2        o271(.A(ori_ori_n245_), .B(ori_ori_n80_), .Y(ori_ori_n288_));
  NO2        o272(.A(ori_ori_n288_), .B(ori_ori_n35_), .Y(ori_ori_n289_));
  NO2        o273(.A(ori_ori_n266_), .B(ori_ori_n185_), .Y(ori_ori_n290_));
  NA2        o274(.A(ori_ori_n290_), .B(ori_ori_n82_), .Y(ori_ori_n291_));
  NA3        o275(.A(ori_ori_n291_), .B(ori_ori_n289_), .C(ori_ori_n287_), .Y(ori_ori_n292_));
  NA2        o276(.A(ori_ori_n292_), .B(ori_ori_n285_), .Y(ori_ori_n293_));
  OAI210     o277(.A0(ori_ori_n106_), .A1(ori_ori_n96_), .B0(ori_ori_n158_), .Y(ori_ori_n294_));
  NA3        o278(.A(ori_ori_n294_), .B(x6), .C(x3), .Y(ori_ori_n295_));
  AOI210     o279(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n296_));
  OAI220     o280(.A0(ori_ori_n296_), .A1(ori_ori_n278_), .B0(ori_ori_n245_), .B1(ori_ori_n275_), .Y(ori_ori_n297_));
  INV        o281(.A(ori_ori_n297_), .Y(ori_ori_n298_));
  NA2        o282(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n299_));
  OAI210     o283(.A0(ori_ori_n96_), .A1(ori_ori_n17_), .B0(ori_ori_n299_), .Y(ori_ori_n300_));
  NA2        o284(.A(ori_ori_n300_), .B(ori_ori_n71_), .Y(ori_ori_n301_));
  NA3        o285(.A(ori_ori_n301_), .B(ori_ori_n298_), .C(ori_ori_n295_), .Y(ori_ori_n302_));
  OAI210     o286(.A0(ori_ori_n101_), .A1(x3), .B0(ori_ori_n269_), .Y(ori_ori_n303_));
  NA2        o287(.A(ori_ori_n193_), .B(ori_ori_n76_), .Y(ori_ori_n304_));
  NA3        o288(.A(ori_ori_n304_), .B(ori_ori_n303_), .C(ori_ori_n136_), .Y(ori_ori_n305_));
  AOI210     o289(.A0(ori_ori_n302_), .A1(x4), .B0(ori_ori_n305_), .Y(ori_ori_n306_));
  NA3        o290(.A(ori_ori_n286_), .B(ori_ori_n189_), .C(ori_ori_n82_), .Y(ori_ori_n307_));
  NOi21      o291(.An(x4), .B(x0), .Y(ori_ori_n308_));
  XO2        o292(.A(x4), .B(x0), .Y(ori_ori_n309_));
  INV        o293(.A(ori_ori_n240_), .Y(ori_ori_n310_));
  AOI220     o294(.A0(ori_ori_n310_), .A1(x8), .B0(ori_ori_n308_), .B1(ori_ori_n83_), .Y(ori_ori_n311_));
  AOI210     o295(.A0(ori_ori_n311_), .A1(ori_ori_n307_), .B0(x3), .Y(ori_ori_n312_));
  INV        o296(.A(ori_ori_n83_), .Y(ori_ori_n313_));
  NO2        o297(.A(ori_ori_n82_), .B(x4), .Y(ori_ori_n314_));
  AOI220     o298(.A0(ori_ori_n314_), .A1(ori_ori_n42_), .B0(ori_ori_n111_), .B1(ori_ori_n313_), .Y(ori_ori_n315_));
  NO2        o299(.A(ori_ori_n309_), .B(x2), .Y(ori_ori_n316_));
  INV        o300(.A(ori_ori_n316_), .Y(ori_ori_n317_));
  NA4        o301(.A(ori_ori_n317_), .B(ori_ori_n315_), .C(ori_ori_n202_), .D(x6), .Y(ori_ori_n318_));
  OAI220     o302(.A0(ori_ori_n268_), .A1(ori_ori_n80_), .B0(ori_ori_n163_), .B1(ori_ori_n82_), .Y(ori_ori_n319_));
  NO2        o303(.A(ori_ori_n41_), .B(x0), .Y(ori_ori_n320_));
  NA2        o304(.A(ori_ori_n319_), .B(ori_ori_n59_), .Y(ori_ori_n321_));
  NO2        o305(.A(ori_ori_n134_), .B(ori_ori_n73_), .Y(ori_ori_n322_));
  NO2        o306(.A(ori_ori_n34_), .B(x2), .Y(ori_ori_n323_));
  NOi21      o307(.An(ori_ori_n108_), .B(ori_ori_n27_), .Y(ori_ori_n324_));
  AOI210     o308(.A0(ori_ori_n323_), .A1(ori_ori_n322_), .B0(ori_ori_n324_), .Y(ori_ori_n325_));
  OAI210     o309(.A0(ori_ori_n321_), .A1(ori_ori_n60_), .B0(ori_ori_n325_), .Y(ori_ori_n326_));
  OAI220     o310(.A0(ori_ori_n326_), .A1(x6), .B0(ori_ori_n318_), .B1(ori_ori_n312_), .Y(ori_ori_n327_));
  NA2        o311(.A(ori_ori_n46_), .B(ori_ori_n40_), .Y(ori_ori_n328_));
  OAI210     o312(.A0(ori_ori_n328_), .A1(ori_ori_n82_), .B0(ori_ori_n279_), .Y(ori_ori_n329_));
  AOI210     o313(.A0(ori_ori_n329_), .A1(ori_ori_n18_), .B0(ori_ori_n136_), .Y(ori_ori_n330_));
  AO220      o314(.A0(ori_ori_n330_), .A1(ori_ori_n327_), .B0(ori_ori_n306_), .B1(ori_ori_n293_), .Y(ori_ori_n331_));
  NA2        o315(.A(ori_ori_n323_), .B(x6), .Y(ori_ori_n332_));
  AOI210     o316(.A0(x6), .A1(x1), .B0(ori_ori_n135_), .Y(ori_ori_n333_));
  NA2        o317(.A(ori_ori_n314_), .B(x0), .Y(ori_ori_n334_));
  NA2        o318(.A(ori_ori_n76_), .B(x6), .Y(ori_ori_n335_));
  OAI210     o319(.A0(ori_ori_n334_), .A1(ori_ori_n333_), .B0(ori_ori_n335_), .Y(ori_ori_n336_));
  AOI220     o320(.A0(ori_ori_n336_), .A1(ori_ori_n332_), .B0(ori_ori_n196_), .B1(ori_ori_n47_), .Y(ori_ori_n337_));
  NA2        o321(.A(ori_ori_n337_), .B(ori_ori_n331_), .Y(ori_ori_n338_));
  AOI210     o322(.A0(ori_ori_n181_), .A1(x8), .B0(ori_ori_n101_), .Y(ori_ori_n339_));
  NA2        o323(.A(ori_ori_n339_), .B(ori_ori_n299_), .Y(ori_ori_n340_));
  NA3        o324(.A(ori_ori_n340_), .B(ori_ori_n179_), .C(ori_ori_n136_), .Y(ori_ori_n341_));
  OAI210     o325(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n210_), .Y(ori_ori_n342_));
  AO220      o326(.A0(ori_ori_n342_), .A1(ori_ori_n133_), .B0(ori_ori_n100_), .B1(x4), .Y(ori_ori_n343_));
  NA3        o327(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n344_));
  NA2        o328(.A(ori_ori_n201_), .B(x0), .Y(ori_ori_n345_));
  OAI220     o329(.A0(ori_ori_n345_), .A1(ori_ori_n189_), .B0(ori_ori_n344_), .B1(ori_ori_n313_), .Y(ori_ori_n346_));
  AOI210     o330(.A0(ori_ori_n343_), .A1(ori_ori_n107_), .B0(ori_ori_n346_), .Y(ori_ori_n347_));
  AOI210     o331(.A0(ori_ori_n347_), .A1(ori_ori_n341_), .B0(ori_ori_n25_), .Y(ori_ori_n348_));
  NAi31      o332(.An(ori_ori_n48_), .B(ori_ori_n257_), .C(ori_ori_n159_), .Y(ori_ori_n349_));
  INV        o333(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  OAI210     o334(.A0(ori_ori_n350_), .A1(ori_ori_n348_), .B0(x6), .Y(ori_ori_n351_));
  NA2        o335(.A(ori_ori_n46_), .B(ori_ori_n119_), .Y(ori_ori_n352_));
  NA3        o336(.A(ori_ori_n53_), .B(ori_ori_n37_), .C(ori_ori_n30_), .Y(ori_ori_n353_));
  AOI220     o337(.A0(ori_ori_n353_), .A1(ori_ori_n352_), .B0(ori_ori_n38_), .B1(ori_ori_n31_), .Y(ori_ori_n354_));
  NO2        o338(.A(ori_ori_n136_), .B(x0), .Y(ori_ori_n355_));
  AOI220     o339(.A0(ori_ori_n355_), .A1(ori_ori_n201_), .B0(ori_ori_n179_), .B1(ori_ori_n136_), .Y(ori_ori_n356_));
  OAI210     o340(.A0(ori_ori_n356_), .A1(x8), .B0(ori_ori_n411_), .Y(ori_ori_n357_));
  NAi31      o341(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n358_));
  OAI210     o342(.A0(ori_ori_n358_), .A1(x4), .B0(ori_ori_n147_), .Y(ori_ori_n359_));
  NA3        o343(.A(ori_ori_n359_), .B(ori_ori_n131_), .C(x9), .Y(ori_ori_n360_));
  NO3        o344(.A(x9), .B(ori_ori_n136_), .C(x0), .Y(ori_ori_n361_));
  AOI220     o345(.A0(ori_ori_n361_), .A1(ori_ori_n224_), .B0(ori_ori_n322_), .B1(ori_ori_n136_), .Y(ori_ori_n362_));
  NA4        o346(.A(ori_ori_n362_), .B(x1), .C(ori_ori_n360_), .D(ori_ori_n48_), .Y(ori_ori_n363_));
  OAI210     o347(.A0(ori_ori_n357_), .A1(ori_ori_n354_), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  NOi31      o348(.An(ori_ori_n355_), .B(ori_ori_n31_), .C(x8), .Y(ori_ori_n365_));
  AOI210     o349(.A0(ori_ori_n37_), .A1(x9), .B0(ori_ori_n117_), .Y(ori_ori_n366_));
  NO2        o350(.A(ori_ori_n366_), .B(ori_ori_n41_), .Y(ori_ori_n367_));
  NOi31      o351(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n368_));
  INV        o352(.A(ori_ori_n368_), .Y(ori_ori_n369_));
  AOI210     o353(.A0(ori_ori_n240_), .A1(ori_ori_n58_), .B0(ori_ori_n110_), .Y(ori_ori_n370_));
  OAI210     o354(.A0(ori_ori_n370_), .A1(x3), .B0(ori_ori_n369_), .Y(ori_ori_n371_));
  NO3        o355(.A(ori_ori_n371_), .B(ori_ori_n367_), .C(x2), .Y(ori_ori_n372_));
  OAI210     o356(.A0(ori_ori_n268_), .A1(ori_ori_n41_), .B0(ori_ori_n309_), .Y(ori_ori_n373_));
  INV        o357(.A(ori_ori_n344_), .Y(ori_ori_n374_));
  AOI220     o358(.A0(ori_ori_n374_), .A1(ori_ori_n82_), .B0(ori_ori_n373_), .B1(ori_ori_n136_), .Y(ori_ori_n375_));
  NO2        o359(.A(ori_ori_n375_), .B(ori_ori_n52_), .Y(ori_ori_n376_));
  NO3        o360(.A(ori_ori_n376_), .B(ori_ori_n372_), .C(ori_ori_n365_), .Y(ori_ori_n377_));
  AOI210     o361(.A0(ori_ori_n377_), .A1(ori_ori_n364_), .B0(ori_ori_n25_), .Y(ori_ori_n378_));
  NA4        o362(.A(ori_ori_n30_), .B(ori_ori_n82_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n379_));
  NO2        o363(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n380_));
  NA2        o364(.A(ori_ori_n380_), .B(ori_ori_n241_), .Y(ori_ori_n381_));
  NO2        o365(.A(ori_ori_n381_), .B(ori_ori_n93_), .Y(ori_ori_n382_));
  NO3        o366(.A(ori_ori_n245_), .B(ori_ori_n158_), .C(ori_ori_n38_), .Y(ori_ori_n383_));
  OAI210     o367(.A0(ori_ori_n383_), .A1(ori_ori_n382_), .B0(x7), .Y(ori_ori_n384_));
  NA2        o368(.A(ori_ori_n206_), .B(x7), .Y(ori_ori_n385_));
  NA3        o369(.A(ori_ori_n385_), .B(ori_ori_n135_), .C(ori_ori_n118_), .Y(ori_ori_n386_));
  NA3        o370(.A(ori_ori_n386_), .B(ori_ori_n384_), .C(ori_ori_n379_), .Y(ori_ori_n387_));
  OAI210     o371(.A0(ori_ori_n387_), .A1(ori_ori_n378_), .B0(ori_ori_n35_), .Y(ori_ori_n388_));
  NO2        o372(.A(ori_ori_n361_), .B(ori_ori_n185_), .Y(ori_ori_n389_));
  NO4        o373(.A(ori_ori_n389_), .B(ori_ori_n70_), .C(x4), .D(ori_ori_n52_), .Y(ori_ori_n390_));
  NA2        o374(.A(ori_ori_n231_), .B(ori_ori_n21_), .Y(ori_ori_n391_));
  NO2        o375(.A(ori_ori_n144_), .B(ori_ori_n119_), .Y(ori_ori_n392_));
  NA2        o376(.A(ori_ori_n392_), .B(ori_ori_n391_), .Y(ori_ori_n393_));
  NO2        o377(.A(ori_ori_n393_), .B(ori_ori_n28_), .Y(ori_ori_n394_));
  AOI220     o378(.A0(ori_ori_n320_), .A1(ori_ori_n82_), .B0(ori_ori_n134_), .B1(ori_ori_n181_), .Y(ori_ori_n395_));
  NA3        o379(.A(ori_ori_n395_), .B(ori_ori_n358_), .C(ori_ori_n80_), .Y(ori_ori_n396_));
  NA2        o380(.A(ori_ori_n396_), .B(ori_ori_n159_), .Y(ori_ori_n397_));
  NO2        o381(.A(ori_ori_n144_), .B(ori_ori_n41_), .Y(ori_ori_n398_));
  NA2        o382(.A(x3), .B(ori_ori_n52_), .Y(ori_ori_n399_));
  OAI210     o383(.A0(ori_ori_n133_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n400_));
  NO3        o384(.A(ori_ori_n368_), .B(x3), .C(ori_ori_n52_), .Y(ori_ori_n401_));
  NA2        o385(.A(ori_ori_n401_), .B(ori_ori_n400_), .Y(ori_ori_n402_));
  OAI210     o386(.A0(ori_ori_n137_), .A1(ori_ori_n399_), .B0(ori_ori_n402_), .Y(ori_ori_n403_));
  AOI220     o387(.A0(ori_ori_n403_), .A1(x0), .B0(ori_ori_n398_), .B1(ori_ori_n119_), .Y(ori_ori_n404_));
  AOI210     o388(.A0(ori_ori_n404_), .A1(ori_ori_n397_), .B0(ori_ori_n214_), .Y(ori_ori_n405_));
  NO3        o389(.A(ori_ori_n405_), .B(ori_ori_n394_), .C(ori_ori_n390_), .Y(ori_ori_n406_));
  NA3        o390(.A(ori_ori_n406_), .B(ori_ori_n388_), .C(ori_ori_n351_), .Y(ori_ori_n407_));
  AOI210     o391(.A0(ori_ori_n338_), .A1(ori_ori_n25_), .B0(ori_ori_n407_), .Y(ori05));
  INV        o392(.A(x1), .Y(ori_ori_n411_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  INV        m005(.A(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x7), .B(x6), .Y(mai_mai_n25_));
  NA2        m009(.A(x8), .B(x3), .Y(mai_mai_n26_));
  NA2        m010(.A(x4), .B(x2), .Y(mai_mai_n27_));
  NO4        m011(.A(mai_mai_n27_), .B(mai_mai_n26_), .C(mai_mai_n25_), .D(mai_mai_n24_), .Y(mai_mai_n28_));
  NO2        m012(.A(mai_mai_n28_), .B(mai_mai_n23_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  NOi21      m015(.An(mai_mai_n22_), .B(mai_mai_n29_), .Y(mai00));
  NO2        m016(.A(x1), .B(x0), .Y(mai_mai_n33_));
  INV        m017(.A(x6), .Y(mai_mai_n34_));
  NO2        m018(.A(mai_mai_n34_), .B(mai_mai_n24_), .Y(mai_mai_n35_));
  AN2        m019(.A(x8), .B(x7), .Y(mai_mai_n36_));
  NA3        m020(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(mai_mai_n33_), .Y(mai_mai_n37_));
  NA2        m021(.A(x4), .B(x3), .Y(mai_mai_n38_));
  AOI210     m022(.A0(mai_mai_n37_), .A1(mai_mai_n22_), .B0(mai_mai_n38_), .Y(mai_mai_n39_));
  NO2        m023(.A(x2), .B(x0), .Y(mai_mai_n40_));
  INV        m024(.A(x3), .Y(mai_mai_n41_));
  NO2        m025(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n42_));
  INV        m026(.A(mai_mai_n42_), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n35_), .B(x4), .Y(mai_mai_n44_));
  OAI210     m028(.A0(mai_mai_n44_), .A1(mai_mai_n43_), .B0(mai_mai_n40_), .Y(mai_mai_n45_));
  INV        m029(.A(x4), .Y(mai_mai_n46_));
  NO2        m030(.A(mai_mai_n46_), .B(mai_mai_n17_), .Y(mai_mai_n47_));
  NA2        m031(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n48_));
  OAI210     m032(.A0(mai_mai_n48_), .A1(mai_mai_n20_), .B0(mai_mai_n45_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n50_), .B(mai_mai_n33_), .Y(mai_mai_n51_));
  INV        m035(.A(x2), .Y(mai_mai_n52_));
  NO2        m036(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n55_));
  OAI210     m039(.A0(mai_mai_n51_), .A1(mai_mai_n31_), .B0(mai_mai_n55_), .Y(mai_mai_n56_));
  NO3        m040(.A(mai_mai_n56_), .B(mai_mai_n49_), .C(mai_mai_n39_), .Y(mai01));
  NA2        m041(.A(x8), .B(x7), .Y(mai_mai_n58_));
  NA2        m042(.A(mai_mai_n41_), .B(x1), .Y(mai_mai_n59_));
  INV        m043(.A(x9), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n60_), .B(mai_mai_n34_), .Y(mai_mai_n61_));
  INV        m045(.A(mai_mai_n61_), .Y(mai_mai_n62_));
  NO3        m046(.A(mai_mai_n62_), .B(mai_mai_n59_), .C(mai_mai_n58_), .Y(mai_mai_n63_));
  NO2        m047(.A(x7), .B(x6), .Y(mai_mai_n64_));
  NO2        m048(.A(mai_mai_n59_), .B(x5), .Y(mai_mai_n65_));
  NO2        m049(.A(x8), .B(x2), .Y(mai_mai_n66_));
  INV        m050(.A(mai_mai_n66_), .Y(mai_mai_n67_));
  NO2        m051(.A(mai_mai_n67_), .B(x1), .Y(mai_mai_n68_));
  OA210      m052(.A0(mai_mai_n68_), .A1(mai_mai_n65_), .B0(mai_mai_n64_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n42_), .A1(mai_mai_n24_), .B0(mai_mai_n52_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n54_), .A1(mai_mai_n20_), .B0(mai_mai_n70_), .Y(mai_mai_n71_));
  NAi31      m055(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n72_));
  NO2        m056(.A(mai_mai_n71_), .B(mai_mai_n69_), .Y(mai_mai_n73_));
  OAI210     m057(.A0(mai_mai_n73_), .A1(mai_mai_n63_), .B0(x4), .Y(mai_mai_n74_));
  NA2        m058(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n75_));
  OAI210     m059(.A0(mai_mai_n75_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n76_));
  NA2        m060(.A(x5), .B(x3), .Y(mai_mai_n77_));
  NO2        m061(.A(x8), .B(x6), .Y(mai_mai_n78_));
  NO4        m062(.A(mai_mai_n78_), .B(mai_mai_n77_), .C(mai_mai_n64_), .D(mai_mai_n52_), .Y(mai_mai_n79_));
  NAi21      m063(.An(x4), .B(x3), .Y(mai_mai_n80_));
  INV        m064(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m065(.A(x4), .B(x2), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(x3), .Y(mai_mai_n83_));
  NO2        m067(.A(mai_mai_n80_), .B(mai_mai_n18_), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n79_), .C(mai_mai_n76_), .Y(mai_mai_n85_));
  NO4        m069(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n41_), .D(x1), .Y(mai_mai_n86_));
  NA2        m070(.A(mai_mai_n60_), .B(mai_mai_n46_), .Y(mai_mai_n87_));
  INV        m071(.A(mai_mai_n87_), .Y(mai_mai_n88_));
  OAI210     m072(.A0(mai_mai_n86_), .A1(mai_mai_n65_), .B0(mai_mai_n88_), .Y(mai_mai_n89_));
  NA2        m073(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n24_), .Y(mai_mai_n91_));
  INV        m075(.A(x8), .Y(mai_mai_n92_));
  NA2        m076(.A(x2), .B(x1), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n92_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n91_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n25_), .Y(mai_mai_n96_));
  AOI210     m080(.A0(mai_mai_n54_), .A1(mai_mai_n24_), .B0(mai_mai_n52_), .Y(mai_mai_n97_));
  OAI210     m081(.A0(mai_mai_n43_), .A1(mai_mai_n35_), .B0(mai_mai_n46_), .Y(mai_mai_n98_));
  NO3        m082(.A(mai_mai_n98_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n99_));
  NA2        m083(.A(x4), .B(mai_mai_n41_), .Y(mai_mai_n100_));
  NO2        m084(.A(mai_mai_n46_), .B(mai_mai_n52_), .Y(mai_mai_n101_));
  OAI210     m085(.A0(mai_mai_n101_), .A1(mai_mai_n41_), .B0(mai_mai_n18_), .Y(mai_mai_n102_));
  AOI210     m086(.A0(mai_mai_n100_), .A1(mai_mai_n50_), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m087(.A(x3), .B(x2), .Y(mai_mai_n104_));
  NA3        m088(.A(mai_mai_n104_), .B(mai_mai_n25_), .C(mai_mai_n24_), .Y(mai_mai_n105_));
  AOI210     m089(.A0(x8), .A1(x6), .B0(mai_mai_n105_), .Y(mai_mai_n106_));
  NA2        m090(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n107_));
  OAI210     m091(.A0(mai_mai_n107_), .A1(mai_mai_n38_), .B0(mai_mai_n17_), .Y(mai_mai_n108_));
  NO4        m092(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n103_), .D(mai_mai_n99_), .Y(mai_mai_n109_));
  AO220      m093(.A0(mai_mai_n109_), .A1(mai_mai_n89_), .B0(mai_mai_n85_), .B1(mai_mai_n74_), .Y(mai02));
  NO2        m094(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n111_));
  NO2        m095(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n112_));
  NA2        m096(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n113_));
  NA2        m097(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n114_));
  OAI210     m098(.A0(mai_mai_n87_), .A1(mai_mai_n113_), .B0(mai_mai_n114_), .Y(mai_mai_n115_));
  AOI220     m099(.A0(mai_mai_n115_), .A1(mai_mai_n112_), .B0(mai_mai_n111_), .B1(x4), .Y(mai_mai_n116_));
  NO3        m100(.A(mai_mai_n116_), .B(x7), .C(x5), .Y(mai_mai_n117_));
  NA2        m101(.A(x9), .B(x2), .Y(mai_mai_n118_));
  OR2        m102(.A(x8), .B(x0), .Y(mai_mai_n119_));
  INV        m103(.A(mai_mai_n119_), .Y(mai_mai_n120_));
  NAi21      m104(.An(x2), .B(x8), .Y(mai_mai_n121_));
  INV        m105(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  OAI220     m106(.A0(mai_mai_n122_), .A1(mai_mai_n120_), .B0(mai_mai_n118_), .B1(x7), .Y(mai_mai_n123_));
  NO2        m107(.A(x4), .B(x1), .Y(mai_mai_n124_));
  NA3        m108(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n58_), .Y(mai_mai_n125_));
  NOi21      m109(.An(x0), .B(x1), .Y(mai_mai_n126_));
  NO3        m110(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n127_));
  NOi21      m111(.An(x0), .B(x4), .Y(mai_mai_n128_));
  NAi21      m112(.An(x8), .B(x7), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n129_), .B(mai_mai_n60_), .Y(mai_mai_n130_));
  AOI220     m114(.A0(mai_mai_n130_), .A1(mai_mai_n128_), .B0(mai_mai_n127_), .B1(mai_mai_n126_), .Y(mai_mai_n131_));
  AOI210     m115(.A0(mai_mai_n131_), .A1(mai_mai_n125_), .B0(mai_mai_n77_), .Y(mai_mai_n132_));
  NO2        m116(.A(x5), .B(mai_mai_n46_), .Y(mai_mai_n133_));
  NA2        m117(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n134_));
  AOI210     m118(.A0(mai_mai_n134_), .A1(mai_mai_n107_), .B0(mai_mai_n114_), .Y(mai_mai_n135_));
  OAI210     m119(.A0(mai_mai_n135_), .A1(mai_mai_n33_), .B0(mai_mai_n133_), .Y(mai_mai_n136_));
  NAi21      m120(.An(x0), .B(x4), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n137_), .B(x1), .Y(mai_mai_n138_));
  NO2        m122(.A(x7), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n82_), .B(mai_mai_n101_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n140_), .B(x3), .Y(mai_mai_n141_));
  OAI210     m125(.A0(mai_mai_n139_), .A1(mai_mai_n138_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NA2        m126(.A(x5), .B(x0), .Y(mai_mai_n143_));
  NO2        m127(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n144_));
  NA3        m128(.A(mai_mai_n142_), .B(mai_mai_n136_), .C(mai_mai_n34_), .Y(mai_mai_n145_));
  NO3        m129(.A(mai_mai_n145_), .B(mai_mai_n132_), .C(mai_mai_n117_), .Y(mai_mai_n146_));
  NO3        m130(.A(mai_mai_n77_), .B(mai_mai_n75_), .C(mai_mai_n23_), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n27_), .B(mai_mai_n24_), .Y(mai_mai_n148_));
  AOI220     m132(.A0(mai_mai_n126_), .A1(mai_mai_n148_), .B0(mai_mai_n65_), .B1(mai_mai_n17_), .Y(mai_mai_n149_));
  NO3        m133(.A(mai_mai_n149_), .B(mai_mai_n58_), .C(mai_mai_n60_), .Y(mai_mai_n150_));
  NA2        m134(.A(x7), .B(x3), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n100_), .B(x5), .Y(mai_mai_n152_));
  NO2        m136(.A(x9), .B(x7), .Y(mai_mai_n153_));
  NOi21      m137(.An(x8), .B(x0), .Y(mai_mai_n154_));
  OA210      m138(.A0(mai_mai_n153_), .A1(x1), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n41_), .B(x2), .Y(mai_mai_n156_));
  INV        m140(.A(x7), .Y(mai_mai_n157_));
  NA2        m141(.A(mai_mai_n157_), .B(mai_mai_n18_), .Y(mai_mai_n158_));
  AOI220     m142(.A0(mai_mai_n158_), .A1(mai_mai_n156_), .B0(mai_mai_n111_), .B1(mai_mai_n36_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n24_), .B(x4), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n128_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n161_), .B(mai_mai_n159_), .Y(mai_mai_n162_));
  AOI210     m146(.A0(mai_mai_n155_), .A1(mai_mai_n152_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  OAI210     m147(.A0(mai_mai_n151_), .A1(mai_mai_n48_), .B0(mai_mai_n163_), .Y(mai_mai_n164_));
  NA2        m148(.A(x5), .B(x1), .Y(mai_mai_n165_));
  INV        m149(.A(mai_mai_n165_), .Y(mai_mai_n166_));
  AOI210     m150(.A0(mai_mai_n166_), .A1(mai_mai_n128_), .B0(mai_mai_n34_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n60_), .B(mai_mai_n92_), .Y(mai_mai_n168_));
  NAi21      m152(.An(x2), .B(x7), .Y(mai_mai_n169_));
  NO3        m153(.A(mai_mai_n169_), .B(mai_mai_n168_), .C(mai_mai_n46_), .Y(mai_mai_n170_));
  NA2        m154(.A(mai_mai_n170_), .B(mai_mai_n65_), .Y(mai_mai_n171_));
  NAi31      m155(.An(mai_mai_n77_), .B(mai_mai_n36_), .C(mai_mai_n33_), .Y(mai_mai_n172_));
  NA3        m156(.A(mai_mai_n172_), .B(mai_mai_n171_), .C(mai_mai_n167_), .Y(mai_mai_n173_));
  NO4        m157(.A(mai_mai_n173_), .B(mai_mai_n164_), .C(mai_mai_n150_), .D(mai_mai_n147_), .Y(mai_mai_n174_));
  NO2        m158(.A(mai_mai_n174_), .B(mai_mai_n146_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n143_), .B(mai_mai_n140_), .Y(mai_mai_n176_));
  NA2        m160(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n177_));
  NA2        m161(.A(mai_mai_n24_), .B(mai_mai_n17_), .Y(mai_mai_n178_));
  NA3        m162(.A(mai_mai_n178_), .B(mai_mai_n177_), .C(mai_mai_n23_), .Y(mai_mai_n179_));
  AN2        m163(.A(mai_mai_n179_), .B(mai_mai_n144_), .Y(mai_mai_n180_));
  NA2        m164(.A(x8), .B(x0), .Y(mai_mai_n181_));
  NO2        m165(.A(mai_mai_n157_), .B(mai_mai_n24_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n126_), .B(x4), .Y(mai_mai_n183_));
  NA2        m167(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  AOI210     m168(.A0(mai_mai_n181_), .A1(mai_mai_n134_), .B0(mai_mai_n184_), .Y(mai_mai_n185_));
  NA2        m169(.A(x2), .B(x0), .Y(mai_mai_n186_));
  NA2        m170(.A(x4), .B(x1), .Y(mai_mai_n187_));
  NAi21      m171(.An(mai_mai_n124_), .B(mai_mai_n187_), .Y(mai_mai_n188_));
  NOi31      m172(.An(mai_mai_n188_), .B(mai_mai_n160_), .C(mai_mai_n186_), .Y(mai_mai_n189_));
  NO4        m173(.A(mai_mai_n189_), .B(mai_mai_n185_), .C(mai_mai_n180_), .D(mai_mai_n176_), .Y(mai_mai_n190_));
  NO2        m174(.A(mai_mai_n190_), .B(mai_mai_n41_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n179_), .B(mai_mai_n75_), .Y(mai_mai_n192_));
  INV        m176(.A(mai_mai_n133_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n107_), .B(mai_mai_n17_), .Y(mai_mai_n194_));
  AOI210     m178(.A0(mai_mai_n33_), .A1(mai_mai_n92_), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  NO3        m179(.A(mai_mai_n195_), .B(mai_mai_n193_), .C(x7), .Y(mai_mai_n196_));
  NA3        m180(.A(mai_mai_n188_), .B(mai_mai_n193_), .C(mai_mai_n40_), .Y(mai_mai_n197_));
  OAI210     m181(.A0(mai_mai_n178_), .A1(mai_mai_n140_), .B0(mai_mai_n197_), .Y(mai_mai_n198_));
  NO3        m182(.A(mai_mai_n198_), .B(mai_mai_n196_), .C(mai_mai_n192_), .Y(mai_mai_n199_));
  NO2        m183(.A(mai_mai_n199_), .B(x3), .Y(mai_mai_n200_));
  NO3        m184(.A(mai_mai_n200_), .B(mai_mai_n191_), .C(mai_mai_n175_), .Y(mai03));
  NO2        m185(.A(mai_mai_n46_), .B(x3), .Y(mai_mai_n202_));
  NO2        m186(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n204_));
  OAI210     m188(.A0(mai_mai_n204_), .A1(mai_mai_n24_), .B0(mai_mai_n61_), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n205_), .B(mai_mai_n17_), .Y(mai_mai_n206_));
  NA2        m190(.A(mai_mai_n206_), .B(mai_mai_n202_), .Y(mai_mai_n207_));
  NA2        m191(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n208_));
  NO2        m192(.A(mai_mai_n208_), .B(x4), .Y(mai_mai_n209_));
  NO2        m193(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n210_));
  NA2        m194(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n211_));
  NO2        m195(.A(mai_mai_n211_), .B(mai_mai_n208_), .Y(mai_mai_n212_));
  NA2        m196(.A(x9), .B(mai_mai_n52_), .Y(mai_mai_n213_));
  NA2        m197(.A(mai_mai_n213_), .B(x4), .Y(mai_mai_n214_));
  NA2        m198(.A(mai_mai_n208_), .B(mai_mai_n80_), .Y(mai_mai_n215_));
  AOI210     m199(.A0(mai_mai_n24_), .A1(x3), .B0(mai_mai_n186_), .Y(mai_mai_n216_));
  AOI220     m200(.A0(mai_mai_n216_), .A1(mai_mai_n215_), .B0(mai_mai_n214_), .B1(mai_mai_n212_), .Y(mai_mai_n217_));
  NO2        m201(.A(x5), .B(x1), .Y(mai_mai_n218_));
  AOI220     m202(.A0(mai_mai_n218_), .A1(mai_mai_n17_), .B0(mai_mai_n104_), .B1(x5), .Y(mai_mai_n219_));
  NO2        m203(.A(mai_mai_n211_), .B(mai_mai_n177_), .Y(mai_mai_n220_));
  NO3        m204(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  OAI210     m206(.A0(mai_mai_n219_), .A1(mai_mai_n62_), .B0(mai_mai_n222_), .Y(mai_mai_n223_));
  NA2        m207(.A(mai_mai_n223_), .B(mai_mai_n46_), .Y(mai_mai_n224_));
  NA3        m208(.A(mai_mai_n224_), .B(mai_mai_n217_), .C(mai_mai_n207_), .Y(mai_mai_n225_));
  NO2        m209(.A(mai_mai_n46_), .B(mai_mai_n41_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n226_), .B(mai_mai_n19_), .Y(mai_mai_n227_));
  NO2        m211(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n228_));
  NO2        m212(.A(mai_mai_n228_), .B(x6), .Y(mai_mai_n229_));
  NOi21      m213(.An(mai_mai_n82_), .B(mai_mai_n229_), .Y(mai_mai_n230_));
  NA2        m214(.A(mai_mai_n60_), .B(mai_mai_n92_), .Y(mai_mai_n231_));
  NA3        m215(.A(mai_mai_n231_), .B(mai_mai_n228_), .C(x6), .Y(mai_mai_n232_));
  AOI210     m216(.A0(mai_mai_n232_), .A1(mai_mai_n230_), .B0(mai_mai_n157_), .Y(mai_mai_n233_));
  AO210      m217(.A0(mai_mai_n233_), .A1(mai_mai_n227_), .B0(mai_mai_n182_), .Y(mai_mai_n234_));
  NA2        m218(.A(mai_mai_n41_), .B(mai_mai_n52_), .Y(mai_mai_n235_));
  NA2        m219(.A(mai_mai_n144_), .B(mai_mai_n91_), .Y(mai_mai_n236_));
  NA2        m220(.A(x6), .B(mai_mai_n46_), .Y(mai_mai_n237_));
  OAI210     m221(.A0(mai_mai_n120_), .A1(mai_mai_n78_), .B0(x4), .Y(mai_mai_n238_));
  AOI210     m222(.A0(mai_mai_n238_), .A1(mai_mai_n237_), .B0(mai_mai_n77_), .Y(mai_mai_n239_));
  NO2        m223(.A(mai_mai_n60_), .B(x6), .Y(mai_mai_n240_));
  NO2        m224(.A(mai_mai_n165_), .B(mai_mai_n41_), .Y(mai_mai_n241_));
  OAI210     m225(.A0(mai_mai_n241_), .A1(mai_mai_n220_), .B0(mai_mai_n240_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n203_), .B(mai_mai_n138_), .Y(mai_mai_n243_));
  NA3        m227(.A(mai_mai_n211_), .B(mai_mai_n133_), .C(x6), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n92_), .A1(mai_mai_n34_), .B0(mai_mai_n65_), .Y(mai_mai_n245_));
  NA4        m229(.A(mai_mai_n245_), .B(mai_mai_n244_), .C(mai_mai_n243_), .D(mai_mai_n242_), .Y(mai_mai_n246_));
  OAI210     m230(.A0(mai_mai_n246_), .A1(mai_mai_n239_), .B0(x2), .Y(mai_mai_n247_));
  NA3        m231(.A(mai_mai_n247_), .B(mai_mai_n236_), .C(mai_mai_n234_), .Y(mai_mai_n248_));
  AOI210     m232(.A0(mai_mai_n225_), .A1(x8), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  NO2        m233(.A(mai_mai_n92_), .B(x3), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n250_), .B(mai_mai_n209_), .Y(mai_mai_n251_));
  NO3        m235(.A(mai_mai_n90_), .B(mai_mai_n78_), .C(mai_mai_n24_), .Y(mai_mai_n252_));
  AOI210     m236(.A0(mai_mai_n229_), .A1(mai_mai_n160_), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  AOI210     m237(.A0(mai_mai_n253_), .A1(mai_mai_n251_), .B0(x2), .Y(mai_mai_n254_));
  NO2        m238(.A(x4), .B(mai_mai_n52_), .Y(mai_mai_n255_));
  AOI220     m239(.A0(mai_mai_n209_), .A1(mai_mai_n194_), .B0(mai_mai_n255_), .B1(mai_mai_n65_), .Y(mai_mai_n256_));
  NA2        m240(.A(mai_mai_n60_), .B(x6), .Y(mai_mai_n257_));
  NA3        m241(.A(mai_mai_n24_), .B(x3), .C(x2), .Y(mai_mai_n258_));
  AOI210     m242(.A0(mai_mai_n258_), .A1(mai_mai_n143_), .B0(mai_mai_n257_), .Y(mai_mai_n259_));
  NA2        m243(.A(mai_mai_n41_), .B(mai_mai_n17_), .Y(mai_mai_n260_));
  NO2        m244(.A(mai_mai_n260_), .B(mai_mai_n24_), .Y(mai_mai_n261_));
  OAI210     m245(.A0(mai_mai_n261_), .A1(mai_mai_n259_), .B0(mai_mai_n124_), .Y(mai_mai_n262_));
  NA2        m246(.A(mai_mai_n211_), .B(x6), .Y(mai_mai_n263_));
  NO2        m247(.A(mai_mai_n211_), .B(x6), .Y(mai_mai_n264_));
  NAi21      m248(.An(mai_mai_n168_), .B(mai_mai_n264_), .Y(mai_mai_n265_));
  NA3        m249(.A(mai_mai_n265_), .B(mai_mai_n263_), .C(mai_mai_n148_), .Y(mai_mai_n266_));
  NA4        m250(.A(mai_mai_n266_), .B(mai_mai_n262_), .C(mai_mai_n256_), .D(mai_mai_n157_), .Y(mai_mai_n267_));
  NA2        m251(.A(mai_mai_n203_), .B(mai_mai_n228_), .Y(mai_mai_n268_));
  NO2        m252(.A(x9), .B(x6), .Y(mai_mai_n269_));
  NO2        m253(.A(mai_mai_n143_), .B(mai_mai_n18_), .Y(mai_mai_n270_));
  NAi21      m254(.An(mai_mai_n270_), .B(mai_mai_n258_), .Y(mai_mai_n271_));
  NAi21      m255(.An(x1), .B(x4), .Y(mai_mai_n272_));
  AOI210     m256(.A0(x3), .A1(x2), .B0(mai_mai_n46_), .Y(mai_mai_n273_));
  OAI210     m257(.A0(mai_mai_n143_), .A1(x3), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  AOI220     m258(.A0(mai_mai_n274_), .A1(mai_mai_n272_), .B0(mai_mai_n271_), .B1(mai_mai_n269_), .Y(mai_mai_n275_));
  NA2        m259(.A(mai_mai_n275_), .B(mai_mai_n268_), .Y(mai_mai_n276_));
  NA2        m260(.A(mai_mai_n60_), .B(x2), .Y(mai_mai_n277_));
  NO2        m261(.A(mai_mai_n277_), .B(mai_mai_n268_), .Y(mai_mai_n278_));
  NO3        m262(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n279_));
  NA2        m263(.A(mai_mai_n107_), .B(mai_mai_n24_), .Y(mai_mai_n280_));
  NA2        m264(.A(x6), .B(x2), .Y(mai_mai_n281_));
  NO2        m265(.A(mai_mai_n281_), .B(mai_mai_n177_), .Y(mai_mai_n282_));
  AOI210     m266(.A0(mai_mai_n280_), .A1(mai_mai_n279_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  OAI220     m267(.A0(mai_mai_n283_), .A1(mai_mai_n41_), .B0(mai_mai_n183_), .B1(mai_mai_n44_), .Y(mai_mai_n284_));
  OAI210     m268(.A0(mai_mai_n284_), .A1(mai_mai_n278_), .B0(mai_mai_n276_), .Y(mai_mai_n285_));
  NO2        m269(.A(x3), .B(mai_mai_n208_), .Y(mai_mai_n286_));
  NA2        m270(.A(x4), .B(x0), .Y(mai_mai_n287_));
  NA2        m271(.A(mai_mai_n286_), .B(mai_mai_n40_), .Y(mai_mai_n288_));
  AOI210     m272(.A0(mai_mai_n288_), .A1(mai_mai_n285_), .B0(x8), .Y(mai_mai_n289_));
  INV        m273(.A(mai_mai_n257_), .Y(mai_mai_n290_));
  OAI210     m274(.A0(mai_mai_n270_), .A1(mai_mai_n218_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  OAI210     m275(.A0(x0), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n292_));
  AOI210     m276(.A0(mai_mai_n292_), .A1(mai_mai_n291_), .B0(mai_mai_n235_), .Y(mai_mai_n293_));
  NO4        m277(.A(mai_mai_n293_), .B(mai_mai_n289_), .C(mai_mai_n267_), .D(mai_mai_n254_), .Y(mai_mai_n294_));
  NO2        m278(.A(mai_mai_n168_), .B(x1), .Y(mai_mai_n295_));
  NO3        m279(.A(mai_mai_n295_), .B(x3), .C(mai_mai_n34_), .Y(mai_mai_n296_));
  OAI210     m280(.A0(mai_mai_n296_), .A1(mai_mai_n264_), .B0(x2), .Y(mai_mai_n297_));
  OAI210     m281(.A0(x0), .A1(x6), .B0(mai_mai_n42_), .Y(mai_mai_n298_));
  AOI210     m282(.A0(mai_mai_n298_), .A1(mai_mai_n297_), .B0(mai_mai_n193_), .Y(mai_mai_n299_));
  NOi21      m283(.An(mai_mai_n281_), .B(mai_mai_n17_), .Y(mai_mai_n300_));
  NA3        m284(.A(mai_mai_n300_), .B(mai_mai_n218_), .C(mai_mai_n38_), .Y(mai_mai_n301_));
  AOI210     m285(.A0(mai_mai_n34_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n302_));
  NA3        m286(.A(mai_mai_n302_), .B(mai_mai_n166_), .C(mai_mai_n31_), .Y(mai_mai_n303_));
  NA2        m287(.A(x3), .B(x2), .Y(mai_mai_n304_));
  AOI220     m288(.A0(mai_mai_n304_), .A1(mai_mai_n235_), .B0(mai_mai_n303_), .B1(mai_mai_n301_), .Y(mai_mai_n305_));
  NAi21      m289(.An(x4), .B(x0), .Y(mai_mai_n306_));
  NO3        m290(.A(mai_mai_n306_), .B(mai_mai_n42_), .C(x2), .Y(mai_mai_n307_));
  OAI210     m291(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n307_), .Y(mai_mai_n308_));
  OAI220     m292(.A0(mai_mai_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n309_));
  NO2        m293(.A(x9), .B(x8), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n34_), .C(mai_mai_n52_), .Y(mai_mai_n311_));
  OAI210     m295(.A0(mai_mai_n302_), .A1(mai_mai_n300_), .B0(mai_mai_n311_), .Y(mai_mai_n312_));
  AOI220     m296(.A0(mai_mai_n312_), .A1(mai_mai_n81_), .B0(mai_mai_n309_), .B1(mai_mai_n30_), .Y(mai_mai_n313_));
  AOI210     m297(.A0(mai_mai_n313_), .A1(mai_mai_n308_), .B0(mai_mai_n24_), .Y(mai_mai_n314_));
  NA3        m298(.A(mai_mai_n34_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n315_));
  OAI210     m299(.A0(mai_mai_n302_), .A1(mai_mai_n300_), .B0(mai_mai_n315_), .Y(mai_mai_n316_));
  INV        m300(.A(mai_mai_n220_), .Y(mai_mai_n317_));
  NA2        m301(.A(mai_mai_n34_), .B(mai_mai_n41_), .Y(mai_mai_n318_));
  OR2        m302(.A(mai_mai_n318_), .B(mai_mai_n287_), .Y(mai_mai_n319_));
  OAI220     m303(.A0(mai_mai_n319_), .A1(mai_mai_n165_), .B0(mai_mai_n237_), .B1(mai_mai_n317_), .Y(mai_mai_n320_));
  AO210      m304(.A0(mai_mai_n316_), .A1(mai_mai_n152_), .B0(mai_mai_n320_), .Y(mai_mai_n321_));
  NO4        m305(.A(mai_mai_n321_), .B(mai_mai_n314_), .C(mai_mai_n305_), .D(mai_mai_n299_), .Y(mai_mai_n322_));
  OAI210     m306(.A0(mai_mai_n294_), .A1(mai_mai_n249_), .B0(mai_mai_n322_), .Y(mai04));
  OAI210     m307(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n324_));
  NA3        m308(.A(mai_mai_n324_), .B(mai_mai_n279_), .C(mai_mai_n83_), .Y(mai_mai_n325_));
  NO2        m309(.A(x2), .B(x1), .Y(mai_mai_n326_));
  OAI210     m310(.A0(mai_mai_n260_), .A1(mai_mai_n326_), .B0(mai_mai_n34_), .Y(mai_mai_n327_));
  NO2        m311(.A(mai_mai_n326_), .B(mai_mai_n306_), .Y(mai_mai_n328_));
  AOI210     m312(.A0(mai_mai_n60_), .A1(x4), .B0(mai_mai_n113_), .Y(mai_mai_n329_));
  OAI210     m313(.A0(mai_mai_n329_), .A1(mai_mai_n328_), .B0(mai_mai_n250_), .Y(mai_mai_n330_));
  NO2        m314(.A(mai_mai_n277_), .B(mai_mai_n90_), .Y(mai_mai_n331_));
  NO2        m315(.A(mai_mai_n331_), .B(mai_mai_n34_), .Y(mai_mai_n332_));
  NO2        m316(.A(mai_mai_n304_), .B(mai_mai_n210_), .Y(mai_mai_n333_));
  NA2        m317(.A(x9), .B(x0), .Y(mai_mai_n334_));
  AOI210     m318(.A0(mai_mai_n90_), .A1(mai_mai_n75_), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  OAI210     m319(.A0(mai_mai_n335_), .A1(mai_mai_n333_), .B0(mai_mai_n92_), .Y(mai_mai_n336_));
  NA3        m320(.A(mai_mai_n336_), .B(mai_mai_n332_), .C(mai_mai_n330_), .Y(mai_mai_n337_));
  NA2        m321(.A(mai_mai_n337_), .B(mai_mai_n327_), .Y(mai_mai_n338_));
  NO2        m322(.A(mai_mai_n213_), .B(mai_mai_n114_), .Y(mai_mai_n339_));
  NO3        m323(.A(mai_mai_n257_), .B(mai_mai_n121_), .C(mai_mai_n18_), .Y(mai_mai_n340_));
  NO2        m324(.A(mai_mai_n340_), .B(mai_mai_n339_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n119_), .A1(mai_mai_n107_), .B0(mai_mai_n181_), .Y(mai_mai_n342_));
  NA3        m326(.A(mai_mai_n342_), .B(x6), .C(x3), .Y(mai_mai_n343_));
  NOi21      m327(.An(mai_mai_n154_), .B(mai_mai_n134_), .Y(mai_mai_n344_));
  AOI210     m328(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n345_));
  OAI220     m329(.A0(mai_mai_n345_), .A1(mai_mai_n318_), .B0(mai_mai_n277_), .B1(mai_mai_n315_), .Y(mai_mai_n346_));
  AOI210     m330(.A0(mai_mai_n344_), .A1(mai_mai_n61_), .B0(mai_mai_n346_), .Y(mai_mai_n347_));
  NA2        m331(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n348_));
  NA2        m332(.A(mai_mai_n331_), .B(mai_mai_n92_), .Y(mai_mai_n349_));
  NA4        m333(.A(mai_mai_n349_), .B(mai_mai_n347_), .C(mai_mai_n343_), .D(mai_mai_n341_), .Y(mai_mai_n350_));
  OAI210     m334(.A0(mai_mai_n112_), .A1(x3), .B0(mai_mai_n307_), .Y(mai_mai_n351_));
  NA2        m335(.A(mai_mai_n351_), .B(mai_mai_n157_), .Y(mai_mai_n352_));
  AOI210     m336(.A0(mai_mai_n350_), .A1(x4), .B0(mai_mai_n352_), .Y(mai_mai_n353_));
  NA3        m337(.A(mai_mai_n328_), .B(mai_mai_n213_), .C(mai_mai_n92_), .Y(mai_mai_n354_));
  NOi21      m338(.An(x4), .B(x0), .Y(mai_mai_n355_));
  XO2        m339(.A(x4), .B(x0), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n356_), .A1(mai_mai_n118_), .B0(mai_mai_n272_), .Y(mai_mai_n357_));
  AOI220     m341(.A0(mai_mai_n357_), .A1(x8), .B0(mai_mai_n355_), .B1(mai_mai_n93_), .Y(mai_mai_n358_));
  AOI210     m342(.A0(mai_mai_n358_), .A1(mai_mai_n354_), .B0(x3), .Y(mai_mai_n359_));
  INV        m343(.A(mai_mai_n93_), .Y(mai_mai_n360_));
  NO2        m344(.A(mai_mai_n92_), .B(x4), .Y(mai_mai_n361_));
  AOI220     m345(.A0(mai_mai_n361_), .A1(mai_mai_n42_), .B0(mai_mai_n128_), .B1(mai_mai_n360_), .Y(mai_mai_n362_));
  NO3        m346(.A(mai_mai_n356_), .B(mai_mai_n168_), .C(x2), .Y(mai_mai_n363_));
  NO3        m347(.A(mai_mai_n231_), .B(mai_mai_n27_), .C(mai_mai_n23_), .Y(mai_mai_n364_));
  NO2        m348(.A(mai_mai_n364_), .B(mai_mai_n363_), .Y(mai_mai_n365_));
  NA4        m349(.A(mai_mai_n365_), .B(mai_mai_n362_), .C(mai_mai_n227_), .D(x6), .Y(mai_mai_n366_));
  NO2        m350(.A(mai_mai_n186_), .B(mai_mai_n92_), .Y(mai_mai_n367_));
  NO2        m351(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n368_));
  BUFFER     m352(.A(mai_mai_n361_), .Y(mai_mai_n369_));
  NO2        m353(.A(mai_mai_n154_), .B(mai_mai_n107_), .Y(mai_mai_n370_));
  AOI220     m354(.A0(mai_mai_n370_), .A1(mai_mai_n369_), .B0(mai_mai_n367_), .B1(mai_mai_n59_), .Y(mai_mai_n371_));
  NO2        m355(.A(mai_mai_n154_), .B(mai_mai_n80_), .Y(mai_mai_n372_));
  NO2        m356(.A(mai_mai_n33_), .B(x2), .Y(mai_mai_n373_));
  NOi21      m357(.An(mai_mai_n124_), .B(mai_mai_n26_), .Y(mai_mai_n374_));
  AOI210     m358(.A0(mai_mai_n373_), .A1(mai_mai_n372_), .B0(mai_mai_n374_), .Y(mai_mai_n375_));
  OAI210     m359(.A0(mai_mai_n371_), .A1(mai_mai_n60_), .B0(mai_mai_n375_), .Y(mai_mai_n376_));
  OAI220     m360(.A0(mai_mai_n376_), .A1(x6), .B0(mai_mai_n366_), .B1(mai_mai_n359_), .Y(mai_mai_n377_));
  OAI210     m361(.A0(mai_mai_n61_), .A1(mai_mai_n46_), .B0(mai_mai_n40_), .Y(mai_mai_n378_));
  OAI210     m362(.A0(mai_mai_n378_), .A1(mai_mai_n92_), .B0(mai_mai_n319_), .Y(mai_mai_n379_));
  AOI210     m363(.A0(mai_mai_n379_), .A1(mai_mai_n18_), .B0(mai_mai_n157_), .Y(mai_mai_n380_));
  AO220      m364(.A0(mai_mai_n380_), .A1(mai_mai_n377_), .B0(mai_mai_n353_), .B1(mai_mai_n338_), .Y(mai_mai_n381_));
  NA2        m365(.A(mai_mai_n221_), .B(mai_mai_n47_), .Y(mai_mai_n382_));
  NA3        m366(.A(mai_mai_n382_), .B(mai_mai_n381_), .C(mai_mai_n325_), .Y(mai_mai_n383_));
  AOI210     m367(.A0(mai_mai_n204_), .A1(x8), .B0(mai_mai_n112_), .Y(mai_mai_n384_));
  NA2        m368(.A(mai_mai_n384_), .B(mai_mai_n348_), .Y(mai_mai_n385_));
  NA3        m369(.A(mai_mai_n385_), .B(mai_mai_n202_), .C(mai_mai_n157_), .Y(mai_mai_n386_));
  NA3        m370(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n387_));
  NO2        m371(.A(mai_mai_n387_), .B(mai_mai_n360_), .Y(mai_mai_n388_));
  INV        m372(.A(mai_mai_n388_), .Y(mai_mai_n389_));
  AOI210     m373(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n24_), .Y(mai_mai_n390_));
  NA3        m374(.A(mai_mai_n122_), .B(mai_mai_n226_), .C(x0), .Y(mai_mai_n391_));
  OAI210     m375(.A0(mai_mai_n202_), .A1(mai_mai_n66_), .B0(mai_mai_n210_), .Y(mai_mai_n392_));
  NA3        m376(.A(mai_mai_n204_), .B(mai_mai_n228_), .C(x8), .Y(mai_mai_n393_));
  AOI210     m377(.A0(mai_mai_n393_), .A1(mai_mai_n392_), .B0(mai_mai_n24_), .Y(mai_mai_n394_));
  AOI210     m378(.A0(mai_mai_n121_), .A1(mai_mai_n119_), .B0(mai_mai_n40_), .Y(mai_mai_n395_));
  NOi31      m379(.An(mai_mai_n395_), .B(mai_mai_n368_), .C(mai_mai_n187_), .Y(mai_mai_n396_));
  OAI210     m380(.A0(mai_mai_n396_), .A1(mai_mai_n394_), .B0(mai_mai_n153_), .Y(mai_mai_n397_));
  NA2        m381(.A(mai_mai_n397_), .B(mai_mai_n391_), .Y(mai_mai_n398_));
  OAI210     m382(.A0(mai_mai_n398_), .A1(mai_mai_n390_), .B0(x6), .Y(mai_mai_n399_));
  OAI210     m383(.A0(mai_mai_n168_), .A1(mai_mai_n46_), .B0(mai_mai_n139_), .Y(mai_mai_n400_));
  AOI210     m384(.A0(mai_mai_n38_), .A1(mai_mai_n31_), .B0(mai_mai_n400_), .Y(mai_mai_n401_));
  NO2        m385(.A(mai_mai_n157_), .B(x0), .Y(mai_mai_n402_));
  AOI220     m386(.A0(mai_mai_n402_), .A1(mai_mai_n226_), .B0(mai_mai_n202_), .B1(mai_mai_n157_), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n130_), .A1(mai_mai_n255_), .B0(x1), .Y(mai_mai_n404_));
  OAI210     m388(.A0(mai_mai_n403_), .A1(x8), .B0(mai_mai_n404_), .Y(mai_mai_n405_));
  NO4        m389(.A(mai_mai_n129_), .B(mai_mai_n306_), .C(x9), .D(x2), .Y(mai_mai_n406_));
  NOi21      m390(.An(mai_mai_n127_), .B(mai_mai_n186_), .Y(mai_mai_n407_));
  NO3        m391(.A(mai_mai_n407_), .B(mai_mai_n406_), .C(mai_mai_n18_), .Y(mai_mai_n408_));
  NA2        m392(.A(mai_mai_n372_), .B(mai_mai_n157_), .Y(mai_mai_n409_));
  NA3        m393(.A(mai_mai_n409_), .B(mai_mai_n408_), .C(mai_mai_n48_), .Y(mai_mai_n410_));
  OAI210     m394(.A0(mai_mai_n405_), .A1(mai_mai_n401_), .B0(mai_mai_n410_), .Y(mai_mai_n411_));
  NOi31      m395(.An(mai_mai_n402_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n412_));
  INV        m396(.A(mai_mai_n137_), .Y(mai_mai_n413_));
  NO3        m397(.A(mai_mai_n413_), .B(mai_mai_n127_), .C(mai_mai_n41_), .Y(mai_mai_n414_));
  AOI210     m398(.A0(mai_mai_n272_), .A1(mai_mai_n58_), .B0(mai_mai_n126_), .Y(mai_mai_n415_));
  NO2        m399(.A(mai_mai_n415_), .B(x3), .Y(mai_mai_n416_));
  NO3        m400(.A(mai_mai_n416_), .B(mai_mai_n414_), .C(x2), .Y(mai_mai_n417_));
  OAI220     m401(.A0(mai_mai_n356_), .A1(mai_mai_n310_), .B0(mai_mai_n306_), .B1(mai_mai_n41_), .Y(mai_mai_n418_));
  AOI210     m402(.A0(x9), .A1(mai_mai_n46_), .B0(mai_mai_n387_), .Y(mai_mai_n419_));
  AOI220     m403(.A0(mai_mai_n419_), .A1(mai_mai_n92_), .B0(mai_mai_n418_), .B1(mai_mai_n157_), .Y(mai_mai_n420_));
  NO2        m404(.A(mai_mai_n420_), .B(mai_mai_n52_), .Y(mai_mai_n421_));
  NO3        m405(.A(mai_mai_n421_), .B(mai_mai_n417_), .C(mai_mai_n412_), .Y(mai_mai_n422_));
  AOI210     m406(.A0(mai_mai_n422_), .A1(mai_mai_n411_), .B0(mai_mai_n24_), .Y(mai_mai_n423_));
  NO3        m407(.A(mai_mai_n60_), .B(x4), .C(x1), .Y(mai_mai_n424_));
  NA2        m408(.A(mai_mai_n424_), .B(mai_mai_n395_), .Y(mai_mai_n425_));
  NO2        m409(.A(mai_mai_n425_), .B(mai_mai_n104_), .Y(mai_mai_n426_));
  NA2        m410(.A(mai_mai_n426_), .B(x7), .Y(mai_mai_n427_));
  NA2        m411(.A(mai_mai_n231_), .B(x7), .Y(mai_mai_n428_));
  NA3        m412(.A(mai_mai_n428_), .B(mai_mai_n156_), .C(mai_mai_n138_), .Y(mai_mai_n429_));
  NA2        m413(.A(mai_mai_n429_), .B(mai_mai_n427_), .Y(mai_mai_n430_));
  OAI210     m414(.A0(mai_mai_n430_), .A1(mai_mai_n423_), .B0(mai_mai_n34_), .Y(mai_mai_n431_));
  INV        m415(.A(mai_mai_n210_), .Y(mai_mai_n432_));
  NO4        m416(.A(mai_mai_n432_), .B(mai_mai_n77_), .C(x4), .D(mai_mai_n52_), .Y(mai_mai_n433_));
  NA2        m417(.A(mai_mai_n260_), .B(mai_mai_n21_), .Y(mai_mai_n434_));
  NO2        m418(.A(mai_mai_n165_), .B(mai_mai_n139_), .Y(mai_mai_n435_));
  NA2        m419(.A(mai_mai_n435_), .B(mai_mai_n434_), .Y(mai_mai_n436_));
  AOI210     m420(.A0(mai_mai_n436_), .A1(mai_mai_n172_), .B0(mai_mai_n27_), .Y(mai_mai_n437_));
  AOI220     m421(.A0(mai_mai_n368_), .A1(mai_mai_n92_), .B0(mai_mai_n154_), .B1(mai_mai_n204_), .Y(mai_mai_n438_));
  NA2        m422(.A(mai_mai_n438_), .B(mai_mai_n90_), .Y(mai_mai_n439_));
  NA2        m423(.A(mai_mai_n439_), .B(mai_mai_n182_), .Y(mai_mai_n440_));
  OAI220     m424(.A0(x3), .A1(mai_mai_n67_), .B0(mai_mai_n165_), .B1(mai_mai_n41_), .Y(mai_mai_n441_));
  NA2        m425(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n442_));
  AOI210     m426(.A0(mai_mai_n169_), .A1(mai_mai_n26_), .B0(mai_mai_n72_), .Y(mai_mai_n443_));
  OAI210     m427(.A0(mai_mai_n153_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n444_));
  NO2        m428(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n445_));
  AOI210     m429(.A0(mai_mai_n445_), .A1(mai_mai_n444_), .B0(mai_mai_n443_), .Y(mai_mai_n446_));
  OAI210     m430(.A0(mai_mai_n158_), .A1(mai_mai_n442_), .B0(mai_mai_n446_), .Y(mai_mai_n447_));
  AOI220     m431(.A0(mai_mai_n447_), .A1(x0), .B0(mai_mai_n441_), .B1(mai_mai_n139_), .Y(mai_mai_n448_));
  AOI210     m432(.A0(mai_mai_n448_), .A1(mai_mai_n440_), .B0(mai_mai_n237_), .Y(mai_mai_n449_));
  NA2        m433(.A(x9), .B(x5), .Y(mai_mai_n450_));
  NO4        m434(.A(mai_mai_n107_), .B(mai_mai_n450_), .C(mai_mai_n58_), .D(mai_mai_n31_), .Y(mai_mai_n451_));
  NO4        m435(.A(mai_mai_n451_), .B(mai_mai_n449_), .C(mai_mai_n437_), .D(mai_mai_n433_), .Y(mai_mai_n452_));
  NA3        m436(.A(mai_mai_n452_), .B(mai_mai_n431_), .C(mai_mai_n399_), .Y(mai_mai_n453_));
  AOI210     m437(.A0(mai_mai_n383_), .A1(mai_mai_n24_), .B0(mai_mai_n453_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  AOI210     u035(.A0(men_men_n22_), .A1(men_men_n19_), .B0(men_men_n35_), .Y(men_men_n52_));
  INV        u036(.A(x2), .Y(men_men_n53_));
  NO2        u037(.A(men_men_n53_), .B(men_men_n17_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  OAI210     u040(.A0(men_men_n52_), .A1(men_men_n32_), .B0(men_men_n56_), .Y(men_men_n57_));
  NO3        u041(.A(men_men_n57_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u042(.A(x8), .B(x7), .Y(men_men_n59_));
  NA2        u043(.A(men_men_n43_), .B(x1), .Y(men_men_n60_));
  INV        u044(.A(x9), .Y(men_men_n61_));
  NO2        u045(.A(men_men_n61_), .B(men_men_n36_), .Y(men_men_n62_));
  INV        u046(.A(men_men_n62_), .Y(men_men_n63_));
  NO3        u047(.A(men_men_n63_), .B(men_men_n60_), .C(men_men_n59_), .Y(men_men_n64_));
  NO2        u048(.A(x7), .B(x6), .Y(men_men_n65_));
  NO2        u049(.A(men_men_n60_), .B(x5), .Y(men_men_n66_));
  NO2        u050(.A(x8), .B(x2), .Y(men_men_n67_));
  INV        u051(.A(men_men_n67_), .Y(men_men_n68_));
  NO2        u052(.A(men_men_n68_), .B(x1), .Y(men_men_n69_));
  OA210      u053(.A0(men_men_n69_), .A1(men_men_n66_), .B0(men_men_n65_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n53_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n55_), .A1(men_men_n20_), .B0(men_men_n71_), .Y(men_men_n72_));
  NAi31      u056(.An(x1), .B(x9), .C(x5), .Y(men_men_n73_));
  OAI220     u057(.A0(men_men_n73_), .A1(men_men_n43_), .B0(men_men_n72_), .B1(men_men_n70_), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n64_), .B0(x4), .Y(men_men_n75_));
  NA2        u059(.A(men_men_n48_), .B(x2), .Y(men_men_n76_));
  OAI210     u060(.A0(men_men_n76_), .A1(men_men_n55_), .B0(x0), .Y(men_men_n77_));
  NA2        u061(.A(x5), .B(x3), .Y(men_men_n78_));
  NO2        u062(.A(x8), .B(x6), .Y(men_men_n79_));
  NO4        u063(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n65_), .D(men_men_n53_), .Y(men_men_n80_));
  NAi21      u064(.An(x4), .B(x3), .Y(men_men_n81_));
  INV        u065(.A(men_men_n81_), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(men_men_n22_), .Y(men_men_n83_));
  NO2        u067(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u068(.A(men_men_n84_), .B(x3), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n83_), .C(men_men_n18_), .Y(men_men_n86_));
  NO3        u070(.A(men_men_n86_), .B(men_men_n80_), .C(men_men_n77_), .Y(men_men_n87_));
  NO4        u071(.A(men_men_n21_), .B(x6), .C(men_men_n43_), .D(x1), .Y(men_men_n88_));
  NA2        u072(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n89_));
  INV        u073(.A(men_men_n89_), .Y(men_men_n90_));
  OAI210     u074(.A0(men_men_n88_), .A1(men_men_n66_), .B0(men_men_n90_), .Y(men_men_n91_));
  NA2        u075(.A(x3), .B(men_men_n18_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n25_), .Y(men_men_n93_));
  INV        u077(.A(x8), .Y(men_men_n94_));
  NA2        u078(.A(x2), .B(x1), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n94_), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n93_), .Y(men_men_n97_));
  NO2        u081(.A(men_men_n97_), .B(men_men_n26_), .Y(men_men_n98_));
  AOI210     u082(.A0(men_men_n55_), .A1(men_men_n25_), .B0(men_men_n53_), .Y(men_men_n99_));
  OAI210     u083(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n100_));
  NO3        u084(.A(men_men_n100_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n101_));
  NA2        u085(.A(x4), .B(men_men_n43_), .Y(men_men_n102_));
  NO2        u086(.A(men_men_n48_), .B(men_men_n53_), .Y(men_men_n103_));
  NO2        u087(.A(men_men_n102_), .B(x1), .Y(men_men_n104_));
  NO2        u088(.A(x3), .B(x2), .Y(men_men_n105_));
  NA3        u089(.A(men_men_n105_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n106_));
  AOI210     u090(.A0(x8), .A1(x6), .B0(men_men_n106_), .Y(men_men_n107_));
  NA2        u091(.A(men_men_n53_), .B(x1), .Y(men_men_n108_));
  OAI210     u092(.A0(men_men_n108_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n109_));
  NO4        u093(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n104_), .D(men_men_n101_), .Y(men_men_n110_));
  AO220      u094(.A0(men_men_n110_), .A1(men_men_n91_), .B0(men_men_n87_), .B1(men_men_n75_), .Y(men02));
  NO2        u095(.A(x3), .B(men_men_n53_), .Y(men_men_n112_));
  NO2        u096(.A(x8), .B(men_men_n18_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n53_), .B(men_men_n17_), .Y(men_men_n114_));
  NA2        u098(.A(men_men_n43_), .B(x0), .Y(men_men_n115_));
  OAI210     u099(.A0(men_men_n89_), .A1(men_men_n114_), .B0(men_men_n115_), .Y(men_men_n116_));
  AOI220     u100(.A0(men_men_n116_), .A1(men_men_n113_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n117_));
  NO3        u101(.A(men_men_n117_), .B(x7), .C(x5), .Y(men_men_n118_));
  NA2        u102(.A(x9), .B(x2), .Y(men_men_n119_));
  OR2        u103(.A(x8), .B(x0), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  NAi21      u105(.An(x2), .B(x8), .Y(men_men_n122_));
  INV        u106(.A(men_men_n122_), .Y(men_men_n123_));
  NO2        u107(.A(x4), .B(x1), .Y(men_men_n124_));
  NA3        u108(.A(men_men_n124_), .B(x0), .C(men_men_n59_), .Y(men_men_n125_));
  NOi21      u109(.An(x0), .B(x1), .Y(men_men_n126_));
  NO3        u110(.A(x9), .B(x8), .C(x7), .Y(men_men_n127_));
  NOi21      u111(.An(x0), .B(x4), .Y(men_men_n128_));
  NAi21      u112(.An(x8), .B(x7), .Y(men_men_n129_));
  NO2        u113(.A(men_men_n129_), .B(men_men_n61_), .Y(men_men_n130_));
  AOI220     u114(.A0(men_men_n130_), .A1(men_men_n128_), .B0(men_men_n127_), .B1(men_men_n126_), .Y(men_men_n131_));
  AOI210     u115(.A0(men_men_n131_), .A1(men_men_n125_), .B0(men_men_n78_), .Y(men_men_n132_));
  NO2        u116(.A(x5), .B(men_men_n48_), .Y(men_men_n133_));
  NA2        u117(.A(x2), .B(men_men_n18_), .Y(men_men_n134_));
  AOI210     u118(.A0(men_men_n134_), .A1(men_men_n108_), .B0(men_men_n115_), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n135_), .A1(men_men_n35_), .B0(men_men_n133_), .Y(men_men_n136_));
  NAi21      u120(.An(x0), .B(x4), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x1), .Y(men_men_n138_));
  NO2        u122(.A(x7), .B(x0), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n84_), .B(men_men_n103_), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n140_), .B(x3), .Y(men_men_n141_));
  OAI210     u125(.A0(men_men_n139_), .A1(men_men_n138_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n21_), .B(men_men_n43_), .Y(men_men_n143_));
  NA2        u127(.A(x5), .B(x0), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n48_), .B(x2), .Y(men_men_n145_));
  NA3        u129(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .Y(men_men_n146_));
  NA4        u130(.A(men_men_n146_), .B(men_men_n142_), .C(men_men_n136_), .D(men_men_n36_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n147_), .B(men_men_n132_), .C(men_men_n118_), .Y(men_men_n148_));
  NO3        u132(.A(men_men_n78_), .B(men_men_n76_), .C(men_men_n24_), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n150_));
  AOI220     u134(.A0(men_men_n126_), .A1(men_men_n150_), .B0(men_men_n66_), .B1(men_men_n17_), .Y(men_men_n151_));
  NO3        u135(.A(men_men_n151_), .B(men_men_n59_), .C(men_men_n61_), .Y(men_men_n152_));
  NA2        u136(.A(x7), .B(x3), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n102_), .B(x5), .Y(men_men_n154_));
  NO2        u138(.A(x9), .B(x7), .Y(men_men_n155_));
  NOi21      u139(.An(x8), .B(x0), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n43_), .B(x2), .Y(men_men_n157_));
  INV        u141(.A(x7), .Y(men_men_n158_));
  NA2        u142(.A(men_men_n158_), .B(men_men_n18_), .Y(men_men_n159_));
  AOI220     u143(.A0(men_men_n159_), .A1(men_men_n157_), .B0(men_men_n112_), .B1(men_men_n38_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n25_), .B(x4), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n161_), .B(men_men_n128_), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n160_), .Y(men_men_n163_));
  AOI210     u147(.A0(men_men_n156_), .A1(men_men_n154_), .B0(men_men_n163_), .Y(men_men_n164_));
  OAI210     u148(.A0(men_men_n153_), .A1(men_men_n50_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA2        u149(.A(x5), .B(x1), .Y(men_men_n166_));
  INV        u150(.A(men_men_n166_), .Y(men_men_n167_));
  AOI210     u151(.A0(men_men_n167_), .A1(men_men_n128_), .B0(men_men_n36_), .Y(men_men_n168_));
  NO2        u152(.A(men_men_n61_), .B(men_men_n94_), .Y(men_men_n169_));
  NAi21      u153(.An(x2), .B(x7), .Y(men_men_n170_));
  NO3        u154(.A(men_men_n170_), .B(men_men_n169_), .C(men_men_n48_), .Y(men_men_n171_));
  NA2        u155(.A(men_men_n171_), .B(men_men_n66_), .Y(men_men_n172_));
  NAi31      u156(.An(men_men_n78_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n173_));
  NA3        u157(.A(men_men_n173_), .B(men_men_n172_), .C(men_men_n168_), .Y(men_men_n174_));
  NO4        u158(.A(men_men_n174_), .B(men_men_n165_), .C(men_men_n152_), .D(men_men_n149_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n175_), .B(men_men_n148_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n144_), .B(men_men_n140_), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n178_));
  NA2        u162(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n179_));
  NA3        u163(.A(men_men_n179_), .B(men_men_n178_), .C(men_men_n24_), .Y(men_men_n180_));
  AN2        u164(.A(men_men_n180_), .B(men_men_n145_), .Y(men_men_n181_));
  NA2        u165(.A(x8), .B(x0), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n158_), .B(men_men_n25_), .Y(men_men_n183_));
  NO2        u167(.A(men_men_n126_), .B(x4), .Y(men_men_n184_));
  NA2        u168(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  AOI210     u169(.A0(men_men_n182_), .A1(men_men_n134_), .B0(men_men_n185_), .Y(men_men_n186_));
  NA2        u170(.A(x2), .B(x0), .Y(men_men_n187_));
  NA2        u171(.A(x4), .B(x1), .Y(men_men_n188_));
  NAi21      u172(.An(men_men_n124_), .B(men_men_n188_), .Y(men_men_n189_));
  NOi31      u173(.An(men_men_n189_), .B(men_men_n161_), .C(men_men_n187_), .Y(men_men_n190_));
  NO4        u174(.A(men_men_n190_), .B(men_men_n186_), .C(men_men_n181_), .D(men_men_n177_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n191_), .B(men_men_n43_), .Y(men_men_n192_));
  NO2        u176(.A(men_men_n180_), .B(men_men_n76_), .Y(men_men_n193_));
  INV        u177(.A(men_men_n133_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n108_), .B(men_men_n17_), .Y(men_men_n195_));
  AOI210     u179(.A0(men_men_n35_), .A1(men_men_n94_), .B0(men_men_n195_), .Y(men_men_n196_));
  NO3        u180(.A(men_men_n196_), .B(men_men_n194_), .C(x7), .Y(men_men_n197_));
  NA3        u181(.A(men_men_n189_), .B(men_men_n194_), .C(men_men_n42_), .Y(men_men_n198_));
  OAI210     u182(.A0(men_men_n179_), .A1(men_men_n140_), .B0(men_men_n198_), .Y(men_men_n199_));
  NO3        u183(.A(men_men_n199_), .B(men_men_n197_), .C(men_men_n193_), .Y(men_men_n200_));
  NO2        u184(.A(men_men_n200_), .B(x3), .Y(men_men_n201_));
  NO3        u185(.A(men_men_n201_), .B(men_men_n192_), .C(men_men_n176_), .Y(men03));
  NO2        u186(.A(men_men_n48_), .B(x3), .Y(men_men_n203_));
  NO2        u187(.A(x6), .B(men_men_n25_), .Y(men_men_n204_));
  INV        u188(.A(men_men_n204_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n53_), .B(x1), .Y(men_men_n206_));
  OAI210     u190(.A0(men_men_n206_), .A1(men_men_n25_), .B0(men_men_n62_), .Y(men_men_n207_));
  OAI220     u191(.A0(men_men_n207_), .A1(men_men_n17_), .B0(men_men_n205_), .B1(men_men_n108_), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n208_), .B(men_men_n203_), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n78_), .B(x6), .Y(men_men_n210_));
  NA2        u194(.A(x6), .B(men_men_n25_), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n211_), .B(x4), .Y(men_men_n212_));
  NO2        u196(.A(men_men_n18_), .B(x0), .Y(men_men_n213_));
  AO220      u197(.A0(men_men_n213_), .A1(men_men_n212_), .B0(men_men_n210_), .B1(men_men_n54_), .Y(men_men_n214_));
  NA2        u198(.A(men_men_n214_), .B(men_men_n61_), .Y(men_men_n215_));
  NA2        u199(.A(x3), .B(men_men_n17_), .Y(men_men_n216_));
  NO2        u200(.A(men_men_n216_), .B(men_men_n211_), .Y(men_men_n217_));
  NA2        u201(.A(x9), .B(men_men_n53_), .Y(men_men_n218_));
  NA2        u202(.A(x9), .B(men_men_n217_), .Y(men_men_n219_));
  NO3        u203(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n220_));
  NO2        u204(.A(x5), .B(x1), .Y(men_men_n221_));
  AOI220     u205(.A0(men_men_n221_), .A1(men_men_n17_), .B0(men_men_n105_), .B1(x5), .Y(men_men_n222_));
  NO2        u206(.A(men_men_n216_), .B(men_men_n178_), .Y(men_men_n223_));
  NO3        u207(.A(x3), .B(x2), .C(x1), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n225_));
  OAI210     u209(.A0(men_men_n222_), .A1(men_men_n63_), .B0(men_men_n225_), .Y(men_men_n226_));
  AOI220     u210(.A0(men_men_n226_), .A1(men_men_n48_), .B0(men_men_n220_), .B1(men_men_n133_), .Y(men_men_n227_));
  NA4        u211(.A(men_men_n227_), .B(men_men_n219_), .C(men_men_n215_), .D(men_men_n209_), .Y(men_men_n228_));
  NO2        u212(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n229_));
  NA2        u213(.A(men_men_n229_), .B(men_men_n19_), .Y(men_men_n230_));
  NO2        u214(.A(x3), .B(men_men_n17_), .Y(men_men_n231_));
  NO2        u215(.A(men_men_n231_), .B(x6), .Y(men_men_n232_));
  NOi21      u216(.An(men_men_n84_), .B(men_men_n232_), .Y(men_men_n233_));
  NA2        u217(.A(men_men_n61_), .B(men_men_n94_), .Y(men_men_n234_));
  NO2        u218(.A(men_men_n233_), .B(men_men_n158_), .Y(men_men_n235_));
  AO210      u219(.A0(men_men_n235_), .A1(men_men_n230_), .B0(men_men_n183_), .Y(men_men_n236_));
  NA2        u220(.A(men_men_n43_), .B(men_men_n53_), .Y(men_men_n237_));
  OAI210     u221(.A0(men_men_n237_), .A1(men_men_n25_), .B0(men_men_n179_), .Y(men_men_n238_));
  NO3        u222(.A(men_men_n188_), .B(men_men_n61_), .C(x6), .Y(men_men_n239_));
  AOI220     u223(.A0(men_men_n239_), .A1(men_men_n238_), .B0(men_men_n145_), .B1(men_men_n93_), .Y(men_men_n240_));
  NA2        u224(.A(x6), .B(men_men_n48_), .Y(men_men_n241_));
  OAI210     u225(.A0(men_men_n121_), .A1(men_men_n79_), .B0(x4), .Y(men_men_n242_));
  AOI210     u226(.A0(men_men_n242_), .A1(men_men_n241_), .B0(men_men_n78_), .Y(men_men_n243_));
  NO2        u227(.A(men_men_n61_), .B(x6), .Y(men_men_n244_));
  NO2        u228(.A(men_men_n166_), .B(men_men_n43_), .Y(men_men_n245_));
  OAI210     u229(.A0(men_men_n245_), .A1(men_men_n223_), .B0(men_men_n244_), .Y(men_men_n246_));
  NA2        u230(.A(men_men_n204_), .B(men_men_n138_), .Y(men_men_n247_));
  NA3        u231(.A(men_men_n216_), .B(men_men_n133_), .C(x6), .Y(men_men_n248_));
  OAI210     u232(.A0(men_men_n94_), .A1(men_men_n36_), .B0(men_men_n66_), .Y(men_men_n249_));
  NA4        u233(.A(men_men_n249_), .B(men_men_n248_), .C(men_men_n247_), .D(men_men_n246_), .Y(men_men_n250_));
  OAI210     u234(.A0(men_men_n250_), .A1(men_men_n243_), .B0(x2), .Y(men_men_n251_));
  NA3        u235(.A(men_men_n251_), .B(men_men_n240_), .C(men_men_n236_), .Y(men_men_n252_));
  AOI210     u236(.A0(men_men_n228_), .A1(x8), .B0(men_men_n252_), .Y(men_men_n253_));
  NO2        u237(.A(men_men_n94_), .B(x3), .Y(men_men_n254_));
  NO3        u238(.A(men_men_n92_), .B(men_men_n79_), .C(men_men_n25_), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n232_), .A1(men_men_n161_), .B0(men_men_n255_), .Y(men_men_n256_));
  NO2        u240(.A(men_men_n256_), .B(x2), .Y(men_men_n257_));
  NO2        u241(.A(x4), .B(men_men_n53_), .Y(men_men_n258_));
  AOI220     u242(.A0(men_men_n212_), .A1(men_men_n195_), .B0(men_men_n258_), .B1(men_men_n66_), .Y(men_men_n259_));
  NA2        u243(.A(men_men_n61_), .B(x6), .Y(men_men_n260_));
  NA3        u244(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n261_));
  AOI210     u245(.A0(men_men_n261_), .A1(men_men_n144_), .B0(men_men_n260_), .Y(men_men_n262_));
  NA2        u246(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n263_), .B(men_men_n25_), .Y(men_men_n264_));
  OAI210     u248(.A0(men_men_n264_), .A1(men_men_n262_), .B0(men_men_n124_), .Y(men_men_n265_));
  NA2        u249(.A(men_men_n216_), .B(x6), .Y(men_men_n266_));
  NO2        u250(.A(men_men_n216_), .B(x6), .Y(men_men_n267_));
  NA2        u251(.A(men_men_n266_), .B(men_men_n150_), .Y(men_men_n268_));
  NA4        u252(.A(men_men_n268_), .B(men_men_n265_), .C(men_men_n259_), .D(men_men_n158_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n204_), .B(men_men_n231_), .Y(men_men_n270_));
  NO2        u254(.A(x9), .B(x6), .Y(men_men_n271_));
  NO2        u255(.A(men_men_n144_), .B(men_men_n18_), .Y(men_men_n272_));
  NAi21      u256(.An(men_men_n272_), .B(men_men_n261_), .Y(men_men_n273_));
  NAi21      u257(.An(x1), .B(x4), .Y(men_men_n274_));
  AOI210     u258(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n275_));
  OAI210     u259(.A0(men_men_n144_), .A1(x3), .B0(men_men_n275_), .Y(men_men_n276_));
  AOI220     u260(.A0(men_men_n276_), .A1(men_men_n274_), .B0(men_men_n273_), .B1(men_men_n271_), .Y(men_men_n277_));
  NA2        u261(.A(men_men_n277_), .B(men_men_n270_), .Y(men_men_n278_));
  NA2        u262(.A(men_men_n61_), .B(x2), .Y(men_men_n279_));
  NO2        u263(.A(men_men_n279_), .B(men_men_n270_), .Y(men_men_n280_));
  NO3        u264(.A(x9), .B(x6), .C(x0), .Y(men_men_n281_));
  NA2        u265(.A(men_men_n108_), .B(men_men_n25_), .Y(men_men_n282_));
  NA2        u266(.A(x6), .B(x2), .Y(men_men_n283_));
  NO2        u267(.A(men_men_n283_), .B(men_men_n178_), .Y(men_men_n284_));
  AOI210     u268(.A0(men_men_n282_), .A1(men_men_n281_), .B0(men_men_n284_), .Y(men_men_n285_));
  OAI220     u269(.A0(men_men_n285_), .A1(men_men_n43_), .B0(men_men_n184_), .B1(men_men_n46_), .Y(men_men_n286_));
  OAI210     u270(.A0(men_men_n286_), .A1(men_men_n280_), .B0(men_men_n278_), .Y(men_men_n287_));
  NA2        u271(.A(x9), .B(men_men_n43_), .Y(men_men_n288_));
  NO2        u272(.A(men_men_n288_), .B(men_men_n211_), .Y(men_men_n289_));
  OR3        u273(.A(men_men_n289_), .B(men_men_n210_), .C(men_men_n154_), .Y(men_men_n290_));
  NA2        u274(.A(x4), .B(x0), .Y(men_men_n291_));
  NO3        u275(.A(men_men_n73_), .B(men_men_n291_), .C(x6), .Y(men_men_n292_));
  AOI210     u276(.A0(men_men_n290_), .A1(men_men_n42_), .B0(men_men_n292_), .Y(men_men_n293_));
  AOI210     u277(.A0(men_men_n293_), .A1(men_men_n287_), .B0(x8), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n272_), .A1(men_men_n221_), .B0(x6), .Y(men_men_n295_));
  INV        u279(.A(men_men_n182_), .Y(men_men_n296_));
  OAI210     u280(.A0(men_men_n296_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n297_));
  AOI210     u281(.A0(men_men_n297_), .A1(men_men_n295_), .B0(men_men_n237_), .Y(men_men_n298_));
  NO4        u282(.A(men_men_n298_), .B(men_men_n294_), .C(men_men_n269_), .D(men_men_n257_), .Y(men_men_n299_));
  NO2        u283(.A(men_men_n169_), .B(x1), .Y(men_men_n300_));
  NO3        u284(.A(men_men_n300_), .B(x3), .C(men_men_n36_), .Y(men_men_n301_));
  OAI210     u285(.A0(men_men_n301_), .A1(men_men_n267_), .B0(x2), .Y(men_men_n302_));
  OAI210     u286(.A0(men_men_n296_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n303_));
  AOI210     u287(.A0(men_men_n303_), .A1(men_men_n302_), .B0(men_men_n194_), .Y(men_men_n304_));
  NOi21      u288(.An(men_men_n283_), .B(men_men_n17_), .Y(men_men_n305_));
  NA3        u289(.A(men_men_n305_), .B(men_men_n221_), .C(men_men_n40_), .Y(men_men_n306_));
  AOI210     u290(.A0(men_men_n36_), .A1(men_men_n53_), .B0(x0), .Y(men_men_n307_));
  NA3        u291(.A(men_men_n307_), .B(men_men_n167_), .C(men_men_n32_), .Y(men_men_n308_));
  NA2        u292(.A(x3), .B(x2), .Y(men_men_n309_));
  AOI220     u293(.A0(men_men_n309_), .A1(men_men_n237_), .B0(men_men_n308_), .B1(men_men_n306_), .Y(men_men_n310_));
  NAi21      u294(.An(x4), .B(x0), .Y(men_men_n311_));
  NO3        u295(.A(men_men_n311_), .B(men_men_n44_), .C(x2), .Y(men_men_n312_));
  OAI210     u296(.A0(x6), .A1(men_men_n18_), .B0(men_men_n312_), .Y(men_men_n313_));
  OAI220     u297(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n314_));
  NO2        u298(.A(x9), .B(x8), .Y(men_men_n315_));
  NA3        u299(.A(men_men_n315_), .B(men_men_n36_), .C(men_men_n53_), .Y(men_men_n316_));
  OAI210     u300(.A0(men_men_n307_), .A1(men_men_n305_), .B0(men_men_n316_), .Y(men_men_n317_));
  AOI220     u301(.A0(men_men_n317_), .A1(men_men_n82_), .B0(men_men_n314_), .B1(men_men_n31_), .Y(men_men_n318_));
  AOI210     u302(.A0(men_men_n318_), .A1(men_men_n313_), .B0(men_men_n25_), .Y(men_men_n319_));
  NA3        u303(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n320_));
  OAI210     u304(.A0(men_men_n307_), .A1(men_men_n305_), .B0(men_men_n320_), .Y(men_men_n321_));
  INV        u305(.A(men_men_n223_), .Y(men_men_n322_));
  NA2        u306(.A(men_men_n36_), .B(men_men_n43_), .Y(men_men_n323_));
  OR2        u307(.A(men_men_n323_), .B(men_men_n291_), .Y(men_men_n324_));
  OAI220     u308(.A0(men_men_n324_), .A1(men_men_n166_), .B0(men_men_n241_), .B1(men_men_n322_), .Y(men_men_n325_));
  AO210      u309(.A0(men_men_n321_), .A1(men_men_n154_), .B0(men_men_n325_), .Y(men_men_n326_));
  NO4        u310(.A(men_men_n326_), .B(men_men_n319_), .C(men_men_n310_), .D(men_men_n304_), .Y(men_men_n327_));
  OAI210     u311(.A0(men_men_n299_), .A1(men_men_n253_), .B0(men_men_n327_), .Y(men04));
  OAI210     u312(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n329_));
  NA3        u313(.A(men_men_n329_), .B(men_men_n281_), .C(men_men_n85_), .Y(men_men_n330_));
  NO2        u314(.A(x2), .B(x1), .Y(men_men_n331_));
  OAI210     u315(.A0(men_men_n263_), .A1(men_men_n331_), .B0(men_men_n36_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n331_), .B(men_men_n311_), .Y(men_men_n333_));
  NA2        u317(.A(men_men_n333_), .B(men_men_n254_), .Y(men_men_n334_));
  NO2        u318(.A(men_men_n279_), .B(men_men_n92_), .Y(men_men_n335_));
  NO2        u319(.A(men_men_n335_), .B(men_men_n36_), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n309_), .B(men_men_n213_), .Y(men_men_n337_));
  NA2        u321(.A(x9), .B(x0), .Y(men_men_n338_));
  AOI210     u322(.A0(men_men_n92_), .A1(men_men_n76_), .B0(men_men_n338_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n339_), .A1(men_men_n337_), .B0(men_men_n94_), .Y(men_men_n340_));
  NA3        u324(.A(men_men_n340_), .B(men_men_n336_), .C(men_men_n334_), .Y(men_men_n341_));
  NA2        u325(.A(men_men_n341_), .B(men_men_n332_), .Y(men_men_n342_));
  NO2        u326(.A(men_men_n218_), .B(men_men_n115_), .Y(men_men_n343_));
  NO3        u327(.A(men_men_n260_), .B(men_men_n122_), .C(men_men_n18_), .Y(men_men_n344_));
  NO2        u328(.A(men_men_n344_), .B(men_men_n343_), .Y(men_men_n345_));
  NOi21      u329(.An(men_men_n156_), .B(men_men_n134_), .Y(men_men_n346_));
  AOI210     u330(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n347_));
  NO2        u331(.A(men_men_n347_), .B(men_men_n323_), .Y(men_men_n348_));
  AOI210     u332(.A0(men_men_n346_), .A1(men_men_n62_), .B0(men_men_n348_), .Y(men_men_n349_));
  NA2        u333(.A(x2), .B(men_men_n17_), .Y(men_men_n350_));
  OAI210     u334(.A0(men_men_n108_), .A1(men_men_n17_), .B0(men_men_n350_), .Y(men_men_n351_));
  AOI220     u335(.A0(men_men_n351_), .A1(men_men_n79_), .B0(men_men_n335_), .B1(men_men_n94_), .Y(men_men_n352_));
  NA3        u336(.A(men_men_n352_), .B(men_men_n349_), .C(men_men_n345_), .Y(men_men_n353_));
  OAI210     u337(.A0(men_men_n113_), .A1(x3), .B0(men_men_n312_), .Y(men_men_n354_));
  NA3        u338(.A(men_men_n234_), .B(men_men_n220_), .C(men_men_n84_), .Y(men_men_n355_));
  NA3        u339(.A(men_men_n355_), .B(men_men_n354_), .C(men_men_n158_), .Y(men_men_n356_));
  AOI210     u340(.A0(men_men_n353_), .A1(x4), .B0(men_men_n356_), .Y(men_men_n357_));
  NOi21      u341(.An(x4), .B(x0), .Y(men_men_n358_));
  XO2        u342(.A(x4), .B(x0), .Y(men_men_n359_));
  OAI210     u343(.A0(men_men_n359_), .A1(men_men_n119_), .B0(men_men_n274_), .Y(men_men_n360_));
  AOI220     u344(.A0(men_men_n360_), .A1(x8), .B0(men_men_n358_), .B1(men_men_n95_), .Y(men_men_n361_));
  NO2        u345(.A(men_men_n361_), .B(x3), .Y(men_men_n362_));
  INV        u346(.A(men_men_n95_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n94_), .B(x4), .Y(men_men_n364_));
  AOI220     u348(.A0(men_men_n364_), .A1(men_men_n44_), .B0(men_men_n128_), .B1(men_men_n363_), .Y(men_men_n365_));
  NO3        u349(.A(men_men_n359_), .B(men_men_n169_), .C(x2), .Y(men_men_n366_));
  NO3        u350(.A(men_men_n234_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n367_));
  NO2        u351(.A(men_men_n367_), .B(men_men_n366_), .Y(men_men_n368_));
  NA4        u352(.A(men_men_n368_), .B(men_men_n365_), .C(men_men_n230_), .D(x6), .Y(men_men_n369_));
  OAI220     u353(.A0(men_men_n311_), .A1(men_men_n92_), .B0(men_men_n187_), .B1(men_men_n94_), .Y(men_men_n370_));
  NO2        u354(.A(men_men_n43_), .B(x0), .Y(men_men_n371_));
  OR2        u355(.A(men_men_n364_), .B(men_men_n371_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n156_), .B(men_men_n108_), .Y(men_men_n373_));
  AOI220     u357(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n370_), .B1(men_men_n60_), .Y(men_men_n374_));
  NO2        u358(.A(men_men_n156_), .B(men_men_n81_), .Y(men_men_n375_));
  NO2        u359(.A(men_men_n35_), .B(x2), .Y(men_men_n376_));
  NA2        u360(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n374_), .A1(men_men_n61_), .B0(men_men_n377_), .Y(men_men_n378_));
  OAI220     u362(.A0(men_men_n378_), .A1(x6), .B0(men_men_n369_), .B1(men_men_n362_), .Y(men_men_n379_));
  OAI210     u363(.A0(men_men_n62_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n380_));
  OAI210     u364(.A0(men_men_n380_), .A1(men_men_n94_), .B0(men_men_n324_), .Y(men_men_n381_));
  AOI210     u365(.A0(men_men_n381_), .A1(men_men_n18_), .B0(men_men_n158_), .Y(men_men_n382_));
  AO220      u366(.A0(men_men_n382_), .A1(men_men_n379_), .B0(men_men_n357_), .B1(men_men_n342_), .Y(men_men_n383_));
  NA2        u367(.A(men_men_n376_), .B(x6), .Y(men_men_n384_));
  AOI210     u368(.A0(x6), .A1(x1), .B0(men_men_n157_), .Y(men_men_n385_));
  NA2        u369(.A(men_men_n364_), .B(x0), .Y(men_men_n386_));
  NA2        u370(.A(men_men_n84_), .B(x6), .Y(men_men_n387_));
  OAI210     u371(.A0(men_men_n386_), .A1(men_men_n385_), .B0(men_men_n387_), .Y(men_men_n388_));
  AOI220     u372(.A0(men_men_n388_), .A1(men_men_n384_), .B0(men_men_n224_), .B1(men_men_n49_), .Y(men_men_n389_));
  NA3        u373(.A(men_men_n389_), .B(men_men_n383_), .C(men_men_n330_), .Y(men_men_n390_));
  NA3        u374(.A(men_men_n113_), .B(men_men_n203_), .C(men_men_n158_), .Y(men_men_n391_));
  OAI210     u375(.A0(men_men_n28_), .A1(x1), .B0(men_men_n237_), .Y(men_men_n392_));
  AO220      u376(.A0(men_men_n392_), .A1(men_men_n155_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n393_));
  NA3        u377(.A(x7), .B(x3), .C(x0), .Y(men_men_n394_));
  NA2        u378(.A(men_men_n229_), .B(x0), .Y(men_men_n395_));
  OAI220     u379(.A0(men_men_n395_), .A1(men_men_n218_), .B0(men_men_n394_), .B1(men_men_n363_), .Y(men_men_n396_));
  AOI210     u380(.A0(men_men_n393_), .A1(men_men_n121_), .B0(men_men_n396_), .Y(men_men_n397_));
  AOI210     u381(.A0(men_men_n397_), .A1(men_men_n391_), .B0(men_men_n25_), .Y(men_men_n398_));
  NA3        u382(.A(men_men_n123_), .B(men_men_n229_), .C(x0), .Y(men_men_n399_));
  OAI210     u383(.A0(men_men_n203_), .A1(men_men_n67_), .B0(men_men_n213_), .Y(men_men_n400_));
  NA3        u384(.A(men_men_n206_), .B(men_men_n231_), .C(x8), .Y(men_men_n401_));
  AOI210     u385(.A0(men_men_n401_), .A1(men_men_n400_), .B0(men_men_n25_), .Y(men_men_n402_));
  AOI210     u386(.A0(men_men_n122_), .A1(men_men_n120_), .B0(men_men_n42_), .Y(men_men_n403_));
  NOi31      u387(.An(men_men_n403_), .B(men_men_n371_), .C(men_men_n188_), .Y(men_men_n404_));
  OAI210     u388(.A0(men_men_n404_), .A1(men_men_n402_), .B0(men_men_n155_), .Y(men_men_n405_));
  NAi31      u389(.An(men_men_n50_), .B(men_men_n300_), .C(men_men_n183_), .Y(men_men_n406_));
  NA3        u390(.A(men_men_n406_), .B(men_men_n405_), .C(men_men_n399_), .Y(men_men_n407_));
  OAI210     u391(.A0(men_men_n407_), .A1(men_men_n398_), .B0(x6), .Y(men_men_n408_));
  INV        u392(.A(men_men_n139_), .Y(men_men_n409_));
  NA3        u393(.A(men_men_n54_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n410_));
  AOI220     u394(.A0(men_men_n410_), .A1(men_men_n409_), .B0(men_men_n40_), .B1(men_men_n32_), .Y(men_men_n411_));
  NA2        u395(.A(men_men_n203_), .B(men_men_n158_), .Y(men_men_n412_));
  AOI210     u396(.A0(men_men_n130_), .A1(men_men_n258_), .B0(x1), .Y(men_men_n413_));
  OAI210     u397(.A0(men_men_n412_), .A1(x8), .B0(men_men_n413_), .Y(men_men_n414_));
  NAi31      u398(.An(x2), .B(x8), .C(x0), .Y(men_men_n415_));
  OAI210     u399(.A0(men_men_n415_), .A1(x4), .B0(men_men_n170_), .Y(men_men_n416_));
  NA3        u400(.A(men_men_n416_), .B(men_men_n153_), .C(x9), .Y(men_men_n417_));
  NO4        u401(.A(men_men_n129_), .B(men_men_n311_), .C(x9), .D(x2), .Y(men_men_n418_));
  NOi21      u402(.An(men_men_n127_), .B(men_men_n187_), .Y(men_men_n419_));
  NO3        u403(.A(men_men_n419_), .B(men_men_n418_), .C(men_men_n18_), .Y(men_men_n420_));
  NO3        u404(.A(x9), .B(men_men_n158_), .C(x0), .Y(men_men_n421_));
  AOI220     u405(.A0(men_men_n421_), .A1(men_men_n254_), .B0(men_men_n375_), .B1(men_men_n158_), .Y(men_men_n422_));
  NA4        u406(.A(men_men_n422_), .B(men_men_n420_), .C(men_men_n417_), .D(men_men_n50_), .Y(men_men_n423_));
  OAI210     u407(.A0(men_men_n414_), .A1(men_men_n411_), .B0(men_men_n423_), .Y(men_men_n424_));
  AOI210     u408(.A0(men_men_n38_), .A1(x9), .B0(men_men_n137_), .Y(men_men_n425_));
  NO3        u409(.A(men_men_n425_), .B(men_men_n127_), .C(men_men_n43_), .Y(men_men_n426_));
  NOi31      u410(.An(x1), .B(x8), .C(x7), .Y(men_men_n427_));
  AOI220     u411(.A0(men_men_n427_), .A1(men_men_n358_), .B0(men_men_n128_), .B1(x3), .Y(men_men_n428_));
  AOI210     u412(.A0(men_men_n274_), .A1(men_men_n59_), .B0(men_men_n126_), .Y(men_men_n429_));
  OAI210     u413(.A0(men_men_n429_), .A1(x3), .B0(men_men_n428_), .Y(men_men_n430_));
  NO3        u414(.A(men_men_n430_), .B(men_men_n426_), .C(x2), .Y(men_men_n431_));
  OAI220     u415(.A0(men_men_n359_), .A1(men_men_n315_), .B0(men_men_n311_), .B1(men_men_n43_), .Y(men_men_n432_));
  AOI210     u416(.A0(x9), .A1(men_men_n48_), .B0(men_men_n394_), .Y(men_men_n433_));
  AOI220     u417(.A0(men_men_n433_), .A1(men_men_n94_), .B0(men_men_n432_), .B1(men_men_n158_), .Y(men_men_n434_));
  NO2        u418(.A(men_men_n434_), .B(men_men_n53_), .Y(men_men_n435_));
  NO2        u419(.A(men_men_n435_), .B(men_men_n431_), .Y(men_men_n436_));
  AOI210     u420(.A0(men_men_n436_), .A1(men_men_n424_), .B0(men_men_n25_), .Y(men_men_n437_));
  NA4        u421(.A(men_men_n31_), .B(men_men_n94_), .C(x2), .D(men_men_n17_), .Y(men_men_n438_));
  NO3        u422(.A(men_men_n61_), .B(x4), .C(x1), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n67_), .B(men_men_n18_), .C(x0), .Y(men_men_n440_));
  AOI220     u424(.A0(men_men_n440_), .A1(men_men_n275_), .B0(men_men_n439_), .B1(men_men_n403_), .Y(men_men_n441_));
  NO2        u425(.A(men_men_n441_), .B(men_men_n105_), .Y(men_men_n442_));
  NO3        u426(.A(men_men_n279_), .B(men_men_n182_), .C(men_men_n40_), .Y(men_men_n443_));
  OAI210     u427(.A0(men_men_n443_), .A1(men_men_n442_), .B0(x7), .Y(men_men_n444_));
  NA2        u428(.A(men_men_n234_), .B(x7), .Y(men_men_n445_));
  NA3        u429(.A(men_men_n445_), .B(men_men_n157_), .C(men_men_n138_), .Y(men_men_n446_));
  NA3        u430(.A(men_men_n446_), .B(men_men_n444_), .C(men_men_n438_), .Y(men_men_n447_));
  OAI210     u431(.A0(men_men_n447_), .A1(men_men_n437_), .B0(men_men_n36_), .Y(men_men_n448_));
  NO2        u432(.A(men_men_n421_), .B(men_men_n213_), .Y(men_men_n449_));
  NO4        u433(.A(men_men_n449_), .B(men_men_n78_), .C(x4), .D(men_men_n53_), .Y(men_men_n450_));
  NO2        u434(.A(men_men_n173_), .B(men_men_n28_), .Y(men_men_n451_));
  NA2        u435(.A(men_men_n415_), .B(men_men_n92_), .Y(men_men_n452_));
  NA2        u436(.A(men_men_n452_), .B(men_men_n183_), .Y(men_men_n453_));
  OAI220     u437(.A0(men_men_n288_), .A1(men_men_n68_), .B0(men_men_n166_), .B1(men_men_n43_), .Y(men_men_n454_));
  AOI210     u438(.A0(men_men_n170_), .A1(men_men_n27_), .B0(men_men_n73_), .Y(men_men_n455_));
  AOI220     u439(.A0(men_men_n455_), .A1(x0), .B0(men_men_n454_), .B1(men_men_n139_), .Y(men_men_n456_));
  AOI210     u440(.A0(men_men_n456_), .A1(men_men_n453_), .B0(men_men_n241_), .Y(men_men_n457_));
  NA2        u441(.A(x9), .B(x5), .Y(men_men_n458_));
  NO4        u442(.A(men_men_n108_), .B(men_men_n458_), .C(men_men_n59_), .D(men_men_n32_), .Y(men_men_n459_));
  NO4        u443(.A(men_men_n459_), .B(men_men_n457_), .C(men_men_n451_), .D(men_men_n450_), .Y(men_men_n460_));
  NA3        u444(.A(men_men_n460_), .B(men_men_n448_), .C(men_men_n408_), .Y(men_men_n461_));
  AOI210     u445(.A0(men_men_n390_), .A1(men_men_n25_), .B0(men_men_n461_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule