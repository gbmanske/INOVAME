//Benchmark atmr_misex3_1774_0.5

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  NOi32      o000(.An(i), .Bn(g), .C(h), .Y(ori_ori_n29_));
  NOi32      o001(.An(j), .Bn(g), .C(k), .Y(ori_ori_n30_));
  NA2        o002(.A(ori_ori_n30_), .B(m), .Y(ori_ori_n31_));
  INV        o003(.A(h), .Y(ori_ori_n32_));
  INV        o004(.A(i), .Y(ori_ori_n33_));
  AN2        o005(.A(h), .B(g), .Y(ori_ori_n34_));
  NAi21      o006(.An(n), .B(m), .Y(ori_ori_n35_));
  NOi32      o007(.An(k), .Bn(h), .C(g), .Y(ori_ori_n36_));
  INV        o008(.A(c), .Y(ori_ori_n37_));
  INV        o009(.A(d), .Y(ori_ori_n38_));
  NAi21      o010(.An(i), .B(h), .Y(ori_ori_n39_));
  INV        o011(.A(n), .Y(ori_ori_n40_));
  NOi32      o012(.An(m), .Bn(j), .C(k), .Y(ori_ori_n41_));
  NAi41      o013(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n42_));
  AN2        o014(.A(e), .B(b), .Y(ori_ori_n43_));
  INV        o015(.A(a), .Y(ori_ori_n44_));
  NOi21      o016(.An(m), .B(n), .Y(ori_ori_n45_));
  INV        o017(.A(b), .Y(ori_ori_n46_));
  NOi31      o018(.An(k), .B(m), .C(j), .Y(ori_ori_n47_));
  NA3        o019(.A(ori_ori_n47_), .B(h), .C(n), .Y(ori_ori_n48_));
  NOi31      o020(.An(k), .B(m), .C(i), .Y(ori_ori_n49_));
  INV        o021(.A(ori_ori_n48_), .Y(ori_ori_n50_));
  NOi32      o022(.An(f), .Bn(b), .C(e), .Y(ori_ori_n51_));
  NAi21      o023(.An(m), .B(n), .Y(ori_ori_n52_));
  NAi31      o024(.An(j), .B(k), .C(h), .Y(ori_ori_n53_));
  NA2        o025(.A(d), .B(b), .Y(ori_ori_n54_));
  NAi21      o026(.An(e), .B(g), .Y(ori_ori_n55_));
  NAi21      o027(.An(c), .B(d), .Y(ori_ori_n56_));
  NAi31      o028(.An(l), .B(k), .C(h), .Y(ori_ori_n57_));
  NO2        o029(.A(ori_ori_n52_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NAi31      o030(.An(e), .B(f), .C(b), .Y(ori_ori_n59_));
  NOi21      o031(.An(k), .B(m), .Y(ori_ori_n60_));
  NOi21      o032(.An(h), .B(g), .Y(ori_ori_n61_));
  NAi31      o033(.An(d), .B(f), .C(c), .Y(ori_ori_n62_));
  NAi31      o034(.An(e), .B(f), .C(c), .Y(ori_ori_n63_));
  NA2        o035(.A(j), .B(h), .Y(ori_ori_n64_));
  OR3        o036(.A(n), .B(m), .C(k), .Y(ori_ori_n65_));
  NO2        o037(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  NO2        o038(.A(n), .B(m), .Y(ori_ori_n67_));
  NA2        o039(.A(ori_ori_n67_), .B(k), .Y(ori_ori_n68_));
  NAi21      o040(.An(f), .B(e), .Y(ori_ori_n69_));
  NA2        o041(.A(d), .B(c), .Y(ori_ori_n70_));
  NO2        o042(.A(ori_ori_n70_), .B(ori_ori_n69_), .Y(ori_ori_n71_));
  NOi21      o043(.An(ori_ori_n71_), .B(ori_ori_n68_), .Y(ori_ori_n72_));
  NAi31      o044(.An(m), .B(n), .C(b), .Y(ori_ori_n73_));
  NAi21      o045(.An(h), .B(f), .Y(ori_ori_n74_));
  NO2        o046(.A(ori_ori_n73_), .B(ori_ori_n56_), .Y(ori_ori_n75_));
  NA2        o047(.A(ori_ori_n75_), .B(k), .Y(ori_ori_n76_));
  NOi32      o048(.An(f), .Bn(c), .C(d), .Y(ori_ori_n77_));
  NOi32      o049(.An(f), .Bn(c), .C(e), .Y(ori_ori_n78_));
  NO2        o050(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  NAi21      o051(.An(ori_ori_n72_), .B(ori_ori_n76_), .Y(ori_ori_n80_));
  OR2        o052(.A(ori_ori_n80_), .B(ori_ori_n50_), .Y(ori_ori_n81_));
  INV        o053(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  NA2        o054(.A(m), .B(j), .Y(ori_ori_n83_));
  NAi31      o055(.An(n), .B(h), .C(g), .Y(ori_ori_n84_));
  NAi41      o056(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n85_));
  INV        o057(.A(f), .Y(ori_ori_n86_));
  INV        o058(.A(g), .Y(ori_ori_n87_));
  NOi31      o059(.An(i), .B(j), .C(h), .Y(ori_ori_n88_));
  NOi21      o060(.An(n), .B(m), .Y(ori_ori_n89_));
  NAi21      o061(.An(j), .B(h), .Y(ori_ori_n90_));
  XN2        o062(.A(i), .B(h), .Y(ori_ori_n91_));
  NOi31      o063(.An(k), .B(n), .C(m), .Y(ori_ori_n92_));
  NAi31      o064(.An(f), .B(e), .C(c), .Y(ori_ori_n93_));
  NO3        o065(.A(ori_ori_n93_), .B(ori_ori_n65_), .C(ori_ori_n64_), .Y(ori_ori_n94_));
  NA3        o066(.A(e), .B(c), .C(b), .Y(ori_ori_n95_));
  NAi32      o067(.An(m), .Bn(i), .C(k), .Y(ori_ori_n96_));
  INV        o068(.A(k), .Y(ori_ori_n97_));
  INV        o069(.A(ori_ori_n94_), .Y(ori_ori_n98_));
  BUFFER     o070(.A(n), .Y(ori_ori_n99_));
  NAi41      o071(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n100_));
  NO2        o072(.A(ori_ori_n100_), .B(e), .Y(ori_ori_n101_));
  BUFFER     o073(.A(g), .Y(ori_ori_n102_));
  NO2        o074(.A(ori_ori_n102_), .B(ori_ori_n42_), .Y(ori_ori_n103_));
  NA2        o075(.A(ori_ori_n103_), .B(ori_ori_n51_), .Y(ori_ori_n104_));
  NO2        o076(.A(n), .B(a), .Y(ori_ori_n105_));
  NAi31      o077(.An(ori_ori_n100_), .B(ori_ori_n105_), .C(ori_ori_n43_), .Y(ori_ori_n106_));
  NAi21      o078(.An(h), .B(i), .Y(ori_ori_n107_));
  NA2        o079(.A(ori_ori_n67_), .B(k), .Y(ori_ori_n108_));
  NO2        o080(.A(ori_ori_n108_), .B(ori_ori_n107_), .Y(ori_ori_n109_));
  NA2        o081(.A(ori_ori_n109_), .B(ori_ori_n77_), .Y(ori_ori_n110_));
  NA3        o082(.A(ori_ori_n110_), .B(ori_ori_n106_), .C(ori_ori_n104_), .Y(ori_ori_n111_));
  NOi21      o083(.An(ori_ori_n98_), .B(ori_ori_n111_), .Y(ori_ori_n112_));
  NA3        o084(.A(ori_ori_n38_), .B(c), .C(b), .Y(ori_ori_n113_));
  NA2        o085(.A(k), .B(h), .Y(ori_ori_n114_));
  NA3        o086(.A(ori_ori_n60_), .B(h), .C(ori_ori_n40_), .Y(ori_ori_n115_));
  NO2        o087(.A(ori_ori_n115_), .B(ori_ori_n79_), .Y(ori_ori_n116_));
  INV        o088(.A(e), .Y(ori_ori_n117_));
  NAi32      o089(.An(j), .Bn(h), .C(i), .Y(ori_ori_n118_));
  NAi21      o090(.An(m), .B(l), .Y(ori_ori_n119_));
  NO3        o091(.A(ori_ori_n119_), .B(ori_ori_n118_), .C(ori_ori_n40_), .Y(ori_ori_n120_));
  NA2        o092(.A(h), .B(g), .Y(ori_ori_n121_));
  NAi32      o093(.An(n), .Bn(m), .C(l), .Y(ori_ori_n122_));
  NO2        o094(.A(ori_ori_n122_), .B(ori_ori_n118_), .Y(ori_ori_n123_));
  NA2        o095(.A(ori_ori_n123_), .B(ori_ori_n71_), .Y(ori_ori_n124_));
  NO2        o096(.A(ori_ori_n463_), .B(ori_ori_n116_), .Y(ori_ori_n125_));
  NA2        o097(.A(ori_ori_n109_), .B(ori_ori_n78_), .Y(ori_ori_n126_));
  NAi21      o098(.An(m), .B(k), .Y(ori_ori_n127_));
  NO2        o099(.A(ori_ori_n91_), .B(ori_ori_n127_), .Y(ori_ori_n128_));
  NAi41      o100(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n129_));
  NA2        o101(.A(n), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  NA2        o102(.A(e), .B(c), .Y(ori_ori_n131_));
  NO3        o103(.A(ori_ori_n131_), .B(n), .C(d), .Y(ori_ori_n132_));
  NOi21      o104(.An(f), .B(h), .Y(ori_ori_n133_));
  NAi31      o105(.An(d), .B(e), .C(b), .Y(ori_ori_n134_));
  NA2        o106(.A(ori_ori_n130_), .B(ori_ori_n126_), .Y(ori_ori_n135_));
  NA2        o107(.A(ori_ori_n105_), .B(ori_ori_n43_), .Y(ori_ori_n136_));
  NOi31      o108(.An(l), .B(n), .C(m), .Y(ori_ori_n137_));
  NA2        o109(.A(ori_ori_n137_), .B(ori_ori_n88_), .Y(ori_ori_n138_));
  NO2        o110(.A(ori_ori_n138_), .B(ori_ori_n79_), .Y(ori_ori_n139_));
  NAi32      o111(.An(m), .Bn(j), .C(k), .Y(ori_ori_n140_));
  NAi41      o112(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n141_));
  INV        o113(.A(ori_ori_n141_), .Y(ori_ori_n142_));
  NOi31      o114(.An(j), .B(m), .C(k), .Y(ori_ori_n143_));
  NO2        o115(.A(ori_ori_n47_), .B(ori_ori_n143_), .Y(ori_ori_n144_));
  NAi21      o116(.An(ori_ori_n144_), .B(ori_ori_n142_), .Y(ori_ori_n145_));
  NO2        o117(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n146_));
  INV        o118(.A(ori_ori_n145_), .Y(ori_ori_n147_));
  NA2        o119(.A(h), .B(g), .Y(ori_ori_n148_));
  NOi32      o120(.An(e), .Bn(b), .C(a), .Y(ori_ori_n149_));
  NA2        o121(.A(ori_ori_n36_), .B(ori_ori_n45_), .Y(ori_ori_n150_));
  NO3        o122(.A(ori_ori_n147_), .B(ori_ori_n139_), .C(ori_ori_n135_), .Y(ori_ori_n151_));
  NA4        o123(.A(ori_ori_n151_), .B(ori_ori_n125_), .C(ori_ori_n112_), .D(ori_ori_n82_), .Y(ori10));
  NO3        o124(.A(ori_ori_n56_), .B(n), .C(ori_ori_n44_), .Y(ori_ori_n153_));
  NAi31      o125(.An(b), .B(f), .C(c), .Y(ori_ori_n154_));
  INV        o126(.A(ori_ori_n154_), .Y(ori_ori_n155_));
  AN2        o127(.A(k), .B(h), .Y(ori_ori_n156_));
  NA2        o128(.A(ori_ori_n156_), .B(ori_ori_n89_), .Y(ori_ori_n157_));
  AN2        o129(.A(j), .B(h), .Y(ori_ori_n158_));
  NO3        o130(.A(n), .B(m), .C(k), .Y(ori_ori_n159_));
  INV        o131(.A(ori_ori_n159_), .Y(ori_ori_n160_));
  NO3        o132(.A(ori_ori_n160_), .B(ori_ori_n56_), .C(ori_ori_n86_), .Y(ori_ori_n161_));
  OR2        o133(.A(m), .B(k), .Y(ori_ori_n162_));
  NO2        o134(.A(ori_ori_n64_), .B(ori_ori_n162_), .Y(ori_ori_n163_));
  NA4        o135(.A(n), .B(f), .C(c), .D(ori_ori_n46_), .Y(ori_ori_n164_));
  INV        o136(.A(ori_ori_n161_), .Y(ori_ori_n165_));
  NO2        o137(.A(ori_ori_n164_), .B(ori_ori_n119_), .Y(ori_ori_n166_));
  NOi32      o138(.An(f), .Bn(d), .C(c), .Y(ori_ori_n167_));
  AOI220     o139(.A0(ori_ori_n167_), .A1(ori_ori_n123_), .B0(ori_ori_n166_), .B1(ori_ori_n88_), .Y(ori_ori_n168_));
  NA2        o140(.A(ori_ori_n168_), .B(ori_ori_n165_), .Y(ori_ori_n169_));
  INV        o141(.A(e), .Y(ori_ori_n170_));
  NA2        o142(.A(ori_ori_n34_), .B(e), .Y(ori_ori_n171_));
  NO2        o143(.A(ori_ori_n171_), .B(ori_ori_n83_), .Y(ori_ori_n172_));
  INV        o144(.A(ori_ori_n172_), .Y(ori_ori_n173_));
  NO2        o145(.A(ori_ori_n173_), .B(a), .Y(ori_ori_n174_));
  NO2        o146(.A(ori_ori_n174_), .B(ori_ori_n169_), .Y(ori_ori_n175_));
  NOi21      o147(.An(d), .B(c), .Y(ori_ori_n176_));
  OR2        o148(.A(n), .B(m), .Y(ori_ori_n177_));
  NO2        o149(.A(ori_ori_n177_), .B(ori_ori_n57_), .Y(ori_ori_n178_));
  INV        o150(.A(ori_ori_n150_), .Y(ori_ori_n179_));
  NA2        o151(.A(ori_ori_n179_), .B(ori_ori_n149_), .Y(ori_ori_n180_));
  NAi21      o152(.An(k), .B(j), .Y(ori_ori_n181_));
  NAi21      o153(.An(e), .B(d), .Y(ori_ori_n182_));
  INV        o154(.A(ori_ori_n182_), .Y(ori_ori_n183_));
  NO2        o155(.A(ori_ori_n108_), .B(ori_ori_n86_), .Y(ori_ori_n184_));
  NA2        o156(.A(ori_ori_n184_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NA2        o157(.A(ori_ori_n185_), .B(ori_ori_n180_), .Y(ori_ori_n186_));
  NO2        o158(.A(ori_ori_n138_), .B(ori_ori_n86_), .Y(ori_ori_n187_));
  NA2        o159(.A(ori_ori_n187_), .B(ori_ori_n183_), .Y(ori_ori_n188_));
  NOi31      o160(.An(n), .B(m), .C(k), .Y(ori_ori_n189_));
  AOI220     o161(.A0(ori_ori_n189_), .A1(ori_ori_n158_), .B0(ori_ori_n89_), .B1(k), .Y(ori_ori_n190_));
  NAi31      o162(.An(g), .B(f), .C(c), .Y(ori_ori_n191_));
  NA2        o163(.A(ori_ori_n188_), .B(ori_ori_n124_), .Y(ori_ori_n192_));
  NO2        o164(.A(ori_ori_n192_), .B(ori_ori_n186_), .Y(ori_ori_n193_));
  AN2        o165(.A(e), .B(d), .Y(ori_ori_n194_));
  NO4        o166(.A(ori_ori_n74_), .B(ori_ori_n42_), .C(ori_ori_n37_), .D(b), .Y(ori_ori_n195_));
  INV        o167(.A(ori_ori_n58_), .Y(ori_ori_n196_));
  AOI210     o168(.A0(ori_ori_n96_), .A1(ori_ori_n140_), .B0(ori_ori_n40_), .Y(ori_ori_n197_));
  INV        o169(.A(ori_ori_n48_), .Y(ori_ori_n198_));
  NA2        o170(.A(ori_ori_n48_), .B(ori_ori_n196_), .Y(ori_ori_n199_));
  NO2        o171(.A(ori_ori_n199_), .B(ori_ori_n195_), .Y(ori_ori_n200_));
  INV        o172(.A(ori_ori_n72_), .Y(ori_ori_n201_));
  NA2        o173(.A(ori_ori_n201_), .B(ori_ori_n98_), .Y(ori_ori_n202_));
  OAI210     o174(.A0(ori_ori_n49_), .A1(ori_ori_n47_), .B0(n), .Y(ori_ori_n203_));
  XO2        o175(.A(i), .B(h), .Y(ori_ori_n204_));
  NA2        o176(.A(ori_ori_n60_), .B(n), .Y(ori_ori_n205_));
  NAi41      o177(.An(ori_ori_n120_), .B(ori_ori_n205_), .C(ori_ori_n190_), .D(ori_ori_n157_), .Y(ori_ori_n206_));
  NOi21      o178(.An(ori_ori_n206_), .B(ori_ori_n113_), .Y(ori_ori_n207_));
  NAi31      o179(.An(c), .B(f), .C(d), .Y(ori_ori_n208_));
  NO2        o180(.A(ori_ori_n115_), .B(ori_ori_n208_), .Y(ori_ori_n209_));
  NO3        o181(.A(ori_ori_n209_), .B(ori_ori_n207_), .C(ori_ori_n202_), .Y(ori_ori_n210_));
  NA4        o182(.A(ori_ori_n210_), .B(ori_ori_n200_), .C(ori_ori_n193_), .D(ori_ori_n175_), .Y(ori11));
  INV        o183(.A(k), .Y(ori_ori_n212_));
  INV        o184(.A(j), .Y(ori_ori_n213_));
  NO2        o185(.A(ori_ori_n114_), .B(ori_ori_n35_), .Y(ori_ori_n214_));
  NOi41      o186(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n215_));
  NAi32      o187(.An(e), .Bn(b), .C(c), .Y(ori_ori_n216_));
  OR2        o188(.A(ori_ori_n216_), .B(ori_ori_n40_), .Y(ori_ori_n217_));
  AN2        o189(.A(ori_ori_n141_), .B(ori_ori_n129_), .Y(ori_ori_n218_));
  NA2        o190(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  OA210      o191(.A0(ori_ori_n219_), .A1(ori_ori_n215_), .B0(ori_ori_n469_), .Y(ori_ori_n220_));
  NO2        o192(.A(ori_ori_n54_), .B(c), .Y(ori_ori_n221_));
  NA3        o193(.A(ori_ori_n221_), .B(j), .C(ori_ori_n189_), .Y(ori_ori_n222_));
  NA3        o194(.A(f), .B(d), .C(b), .Y(ori_ori_n223_));
  NO4        o195(.A(ori_ori_n223_), .B(m), .C(ori_ori_n64_), .D(g), .Y(ori_ori_n224_));
  INV        o196(.A(ori_ori_n222_), .Y(ori_ori_n225_));
  NO2        o197(.A(ori_ori_n225_), .B(ori_ori_n220_), .Y(ori_ori_n226_));
  NO3        o198(.A(ori_ori_n127_), .B(ori_ori_n39_), .C(n), .Y(ori_ori_n227_));
  NA3        o199(.A(ori_ori_n208_), .B(ori_ori_n63_), .C(ori_ori_n62_), .Y(ori_ori_n228_));
  NA2        o200(.A(ori_ori_n191_), .B(ori_ori_n93_), .Y(ori_ori_n229_));
  OR2        o201(.A(ori_ori_n229_), .B(ori_ori_n228_), .Y(ori_ori_n230_));
  NA2        o202(.A(ori_ori_n230_), .B(ori_ori_n227_), .Y(ori_ori_n231_));
  INV        o203(.A(ori_ori_n231_), .Y(ori_ori_n232_));
  NOi32      o204(.An(e), .Bn(c), .C(f), .Y(ori_ori_n233_));
  INV        o205(.A(ori_ori_n85_), .Y(ori_ori_n234_));
  NA2        o206(.A(ori_ori_n204_), .B(ori_ori_n60_), .Y(ori_ori_n235_));
  AN3        o207(.A(f), .B(d), .C(b), .Y(ori_ori_n236_));
  OAI210     o208(.A0(ori_ori_n236_), .A1(ori_ori_n51_), .B0(n), .Y(ori_ori_n237_));
  NA2        o209(.A(ori_ori_n60_), .B(ori_ori_n87_), .Y(ori_ori_n238_));
  AOI210     o210(.A0(ori_ori_n237_), .A1(ori_ori_n95_), .B0(ori_ori_n238_), .Y(ori_ori_n239_));
  NAi31      o211(.An(m), .B(n), .C(k), .Y(ori_ori_n240_));
  INV        o212(.A(ori_ori_n106_), .Y(ori_ori_n241_));
  NO2        o213(.A(ori_ori_n241_), .B(ori_ori_n239_), .Y(ori_ori_n242_));
  INV        o214(.A(ori_ori_n242_), .Y(ori_ori_n243_));
  NO2        o215(.A(ori_ori_n243_), .B(ori_ori_n232_), .Y(ori_ori_n244_));
  NA2        o216(.A(ori_ori_n153_), .B(ori_ori_n61_), .Y(ori_ori_n245_));
  NO2        o217(.A(ori_ori_n245_), .B(ori_ori_n212_), .Y(ori_ori_n246_));
  NO3        o218(.A(g), .B(ori_ori_n86_), .C(ori_ori_n37_), .Y(ori_ori_n247_));
  OAI210     o219(.A0(ori_ori_n92_), .A1(ori_ori_n163_), .B0(ori_ori_n247_), .Y(ori_ori_n248_));
  NA2        o220(.A(h), .B(ori_ori_n30_), .Y(ori_ori_n249_));
  NA2        o221(.A(ori_ori_n41_), .B(ori_ori_n34_), .Y(ori_ori_n250_));
  NO2        o222(.A(ori_ori_n250_), .B(ori_ori_n136_), .Y(ori_ori_n251_));
  INV        o223(.A(ori_ori_n251_), .Y(ori_ori_n252_));
  NA2        o224(.A(ori_ori_n252_), .B(ori_ori_n248_), .Y(ori_ori_n253_));
  NO3        o225(.A(ori_ori_n167_), .B(ori_ori_n78_), .C(ori_ori_n77_), .Y(ori_ori_n254_));
  NA2        o226(.A(ori_ori_n254_), .B(ori_ori_n93_), .Y(ori_ori_n255_));
  NA2        o227(.A(ori_ori_n255_), .B(ori_ori_n109_), .Y(ori_ori_n256_));
  NO2        o228(.A(ori_ori_n191_), .B(ori_ori_n64_), .Y(ori_ori_n257_));
  NA2        o229(.A(ori_ori_n256_), .B(ori_ori_n165_), .Y(ori_ori_n258_));
  NO3        o230(.A(ori_ori_n258_), .B(ori_ori_n253_), .C(ori_ori_n246_), .Y(ori_ori_n259_));
  NA3        o231(.A(ori_ori_n259_), .B(ori_ori_n244_), .C(ori_ori_n226_), .Y(ori08));
  NO2        o232(.A(k), .B(h), .Y(ori_ori_n261_));
  AO210      o233(.A0(ori_ori_n107_), .A1(ori_ori_n181_), .B0(ori_ori_n261_), .Y(ori_ori_n262_));
  NO2        o234(.A(ori_ori_n262_), .B(ori_ori_n119_), .Y(ori_ori_n263_));
  NA2        o235(.A(ori_ori_n233_), .B(ori_ori_n40_), .Y(ori_ori_n264_));
  NA2        o236(.A(ori_ori_n264_), .B(ori_ori_n191_), .Y(ori_ori_n265_));
  NA2        o237(.A(ori_ori_n265_), .B(ori_ori_n263_), .Y(ori_ori_n266_));
  AOI210     o238(.A0(ori_ori_n223_), .A1(ori_ori_n59_), .B0(ori_ori_n40_), .Y(ori_ori_n267_));
  INV        o239(.A(ori_ori_n266_), .Y(ori_ori_n268_));
  NO2        o240(.A(ori_ori_n127_), .B(g), .Y(ori_ori_n269_));
  NA3        o241(.A(ori_ori_n255_), .B(ori_ori_n137_), .C(ori_ori_n156_), .Y(ori_ori_n270_));
  INV        o242(.A(ori_ori_n270_), .Y(ori_ori_n271_));
  NO3        o243(.A(ori_ori_n271_), .B(ori_ori_n166_), .C(ori_ori_n268_), .Y(ori_ori_n272_));
  NA2        o244(.A(ori_ori_n234_), .B(ori_ori_n163_), .Y(ori_ori_n273_));
  NA3        o245(.A(ori_ori_n150_), .B(ori_ori_n273_), .C(ori_ori_n106_), .Y(ori_ori_n274_));
  NO2        o246(.A(ori_ori_n274_), .B(ori_ori_n257_), .Y(ori_ori_n275_));
  NA2        o247(.A(ori_ori_n229_), .B(ori_ori_n123_), .Y(ori_ori_n276_));
  INV        o248(.A(ori_ori_n276_), .Y(ori_ori_n277_));
  NO2        o249(.A(ori_ori_n119_), .B(ori_ori_n53_), .Y(ori_ori_n278_));
  AOI220     o250(.A0(ori_ori_n278_), .A1(ori_ori_n234_), .B0(ori_ori_n269_), .B1(ori_ori_n267_), .Y(ori_ori_n279_));
  INV        o251(.A(ori_ori_n279_), .Y(ori_ori_n280_));
  OR2        o252(.A(ori_ori_n280_), .B(ori_ori_n277_), .Y(ori_ori_n281_));
  INV        o253(.A(ori_ori_n217_), .Y(ori_ori_n282_));
  NA2        o254(.A(ori_ori_n282_), .B(ori_ori_n29_), .Y(ori_ori_n283_));
  NO2        o255(.A(ori_ori_n136_), .B(ori_ori_n31_), .Y(ori_ori_n284_));
  INV        o256(.A(ori_ori_n284_), .Y(ori_ori_n285_));
  NA2        o257(.A(ori_ori_n285_), .B(ori_ori_n283_), .Y(ori_ori_n286_));
  NO3        o258(.A(ori_ori_n139_), .B(ori_ori_n286_), .C(ori_ori_n281_), .Y(ori_ori_n287_));
  INV        o259(.A(ori_ori_n144_), .Y(ori_ori_n288_));
  INV        o260(.A(ori_ori_n168_), .Y(ori_ori_n289_));
  NO2        o261(.A(ori_ori_n216_), .B(ori_ori_n40_), .Y(ori_ori_n290_));
  NA2        o262(.A(ori_ori_n288_), .B(ori_ori_n290_), .Y(ori_ori_n291_));
  INV        o263(.A(ori_ori_n291_), .Y(ori_ori_n292_));
  NO2        o264(.A(ori_ori_n254_), .B(n), .Y(ori_ori_n293_));
  BUFFER     o265(.A(ori_ori_n278_), .Y(ori_ori_n294_));
  AOI220     o266(.A0(ori_ori_n294_), .A1(ori_ori_n247_), .B0(ori_ori_n293_), .B1(ori_ori_n263_), .Y(ori_ori_n295_));
  INV        o267(.A(ori_ori_n295_), .Y(ori_ori_n296_));
  NO3        o268(.A(ori_ori_n296_), .B(ori_ori_n292_), .C(ori_ori_n289_), .Y(ori_ori_n297_));
  NA4        o269(.A(ori_ori_n297_), .B(ori_ori_n287_), .C(ori_ori_n275_), .D(ori_ori_n272_), .Y(ori09));
  NO2        o270(.A(ori_ori_n49_), .B(ori_ori_n47_), .Y(ori_ori_n299_));
  NO2        o271(.A(ori_ori_n299_), .B(f), .Y(ori_ori_n300_));
  NA2        o272(.A(ori_ori_n300_), .B(n), .Y(ori_ori_n301_));
  NA2        o273(.A(ori_ori_n262_), .B(ori_ori_n53_), .Y(ori_ori_n302_));
  NA2        o274(.A(ori_ori_n302_), .B(ori_ori_n75_), .Y(ori_ori_n303_));
  NA2        o275(.A(ori_ori_n303_), .B(ori_ori_n301_), .Y(ori_ori_n304_));
  NO2        o276(.A(ori_ori_n240_), .B(ori_ori_n134_), .Y(ori_ori_n305_));
  NO3        o277(.A(ori_ori_n120_), .B(ori_ori_n198_), .C(ori_ori_n304_), .Y(ori_ori_n306_));
  NO2        o278(.A(ori_ori_n93_), .B(ori_ori_n90_), .Y(ori_ori_n307_));
  NA2        o279(.A(ori_ori_n307_), .B(ori_ori_n92_), .Y(ori_ori_n308_));
  NA2        o280(.A(e), .B(d), .Y(ori_ori_n309_));
  OAI220     o281(.A0(ori_ori_n309_), .A1(c), .B0(ori_ori_n131_), .B1(d), .Y(ori_ori_n310_));
  NA3        o282(.A(ori_ori_n310_), .B(ori_ori_n184_), .C(ori_ori_n204_), .Y(ori_ori_n311_));
  AOI220     o283(.A0(h), .A1(ori_ori_n305_), .B0(ori_ori_n227_), .B1(ori_ori_n233_), .Y(ori_ori_n312_));
  AO210      o284(.A0(ori_ori_n184_), .A1(h), .B0(ori_ori_n66_), .Y(ori_ori_n313_));
  OAI210     o285(.A0(ori_ori_n313_), .A1(ori_ori_n187_), .B0(ori_ori_n310_), .Y(ori_ori_n314_));
  AN3        o286(.A(ori_ori_n314_), .B(ori_ori_n312_), .C(ori_ori_n264_), .Y(ori_ori_n315_));
  NA3        o287(.A(ori_ori_n315_), .B(ori_ori_n311_), .C(ori_ori_n306_), .Y(ori12));
  NO2        o288(.A(ori_ori_n182_), .B(c), .Y(ori_ori_n317_));
  NO3        o289(.A(ori_ori_n177_), .B(ori_ori_n107_), .C(ori_ori_n87_), .Y(ori_ori_n318_));
  NA2        o290(.A(ori_ori_n318_), .B(ori_ori_n317_), .Y(ori_ori_n319_));
  INV        o291(.A(ori_ori_n182_), .Y(ori_ori_n320_));
  NO2        o292(.A(ori_ori_n299_), .B(ori_ori_n148_), .Y(ori_ori_n321_));
  NA2        o293(.A(ori_ori_n321_), .B(ori_ori_n320_), .Y(ori_ori_n322_));
  NA2        o294(.A(ori_ori_n322_), .B(ori_ori_n319_), .Y(ori_ori_n323_));
  AOI210     o295(.A0(ori_ori_n96_), .A1(ori_ori_n140_), .B0(ori_ori_n84_), .Y(ori_ori_n324_));
  OR2        o296(.A(ori_ori_n324_), .B(ori_ori_n318_), .Y(ori_ori_n325_));
  OAI210     o297(.A0(ori_ori_n159_), .A1(ori_ori_n325_), .B0(ori_ori_n167_), .Y(ori_ori_n326_));
  NO2        o298(.A(ori_ori_n56_), .B(ori_ori_n99_), .Y(ori_ori_n327_));
  NA2        o299(.A(ori_ori_n327_), .B(ori_ori_n101_), .Y(ori_ori_n328_));
  NA2        o300(.A(ori_ori_n328_), .B(ori_ori_n326_), .Y(ori_ori_n329_));
  NA2        o301(.A(ori_ori_n178_), .B(ori_ori_n176_), .Y(ori_ori_n330_));
  INV        o302(.A(ori_ori_n330_), .Y(ori_ori_n331_));
  NO3        o303(.A(ori_ori_n331_), .B(ori_ori_n329_), .C(ori_ori_n323_), .Y(ori_ori_n332_));
  NOi21      o304(.An(ori_ori_n29_), .B(ori_ori_n240_), .Y(ori_ori_n333_));
  INV        o305(.A(ori_ori_n106_), .Y(ori_ori_n334_));
  INV        o306(.A(ori_ori_n130_), .Y(ori_ori_n335_));
  INV        o307(.A(ori_ori_n203_), .Y(ori_ori_n336_));
  NO2        o308(.A(ori_ori_n335_), .B(ori_ori_n334_), .Y(ori_ori_n337_));
  INV        o309(.A(ori_ori_n146_), .Y(ori_ori_n338_));
  NA2        o310(.A(ori_ori_n61_), .B(i), .Y(ori_ori_n339_));
  NA2        o311(.A(ori_ori_n34_), .B(i), .Y(ori_ori_n340_));
  NO2        o312(.A(ori_ori_n340_), .B(ori_ori_n83_), .Y(ori_ori_n341_));
  INV        o313(.A(ori_ori_n341_), .Y(ori_ori_n342_));
  NO2        o314(.A(n), .B(ori_ori_n215_), .Y(ori_ori_n343_));
  OAI220     o315(.A0(ori_ori_n343_), .A1(ori_ori_n338_), .B0(ori_ori_n342_), .B1(ori_ori_n136_), .Y(ori_ori_n344_));
  NA3        o316(.A(ori_ori_n133_), .B(i), .C(g), .Y(ori_ori_n345_));
  AOI210     o317(.A0(ori_ori_n249_), .A1(ori_ori_n345_), .B0(m), .Y(ori_ori_n346_));
  OAI210     o318(.A0(ori_ori_n346_), .A1(ori_ori_n321_), .B0(ori_ori_n132_), .Y(ori_ori_n347_));
  INV        o319(.A(ori_ori_n347_), .Y(ori_ori_n348_));
  NO2        o320(.A(ori_ori_n190_), .B(ori_ori_n87_), .Y(ori_ori_n349_));
  NA2        o321(.A(ori_ori_n349_), .B(ori_ori_n155_), .Y(ori_ori_n350_));
  INV        o322(.A(ori_ori_n350_), .Y(ori_ori_n351_));
  NA2        o323(.A(ori_ori_n346_), .B(ori_ori_n320_), .Y(ori_ori_n352_));
  INV        o324(.A(ori_ori_n352_), .Y(ori_ori_n353_));
  NO4        o325(.A(ori_ori_n353_), .B(ori_ori_n351_), .C(ori_ori_n348_), .D(ori_ori_n344_), .Y(ori_ori_n354_));
  NA2        o326(.A(h), .B(n), .Y(ori_ori_n355_));
  NO2        o327(.A(ori_ori_n47_), .B(ori_ori_n143_), .Y(ori_ori_n356_));
  NO2        o328(.A(ori_ori_n356_), .B(ori_ori_n355_), .Y(ori_ori_n357_));
  NA2        o329(.A(ori_ori_n93_), .B(ori_ori_n63_), .Y(ori_ori_n358_));
  NO2        o330(.A(ori_ori_n178_), .B(ori_ori_n66_), .Y(ori_ori_n359_));
  NOi31      o331(.An(ori_ori_n358_), .B(ori_ori_n359_), .C(ori_ori_n87_), .Y(ori_ori_n360_));
  NAi21      o332(.An(ori_ori_n216_), .B(ori_ori_n349_), .Y(ori_ori_n361_));
  INV        o333(.A(ori_ori_n195_), .Y(ori_ori_n362_));
  NA2        o334(.A(ori_ori_n362_), .B(ori_ori_n361_), .Y(ori_ori_n363_));
  NA2        o335(.A(ori_ori_n324_), .B(ori_ori_n317_), .Y(ori_ori_n364_));
  OAI210     o336(.A0(ori_ori_n324_), .A1(ori_ori_n318_), .B0(ori_ori_n358_), .Y(ori_ori_n365_));
  NA2        o337(.A(ori_ori_n197_), .B(ori_ori_n34_), .Y(ori_ori_n366_));
  NA2        o338(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n367_));
  NO4        o339(.A(ori_ori_n367_), .B(ori_ori_n363_), .C(ori_ori_n360_), .D(ori_ori_n357_), .Y(ori_ori_n368_));
  NA4        o340(.A(ori_ori_n368_), .B(ori_ori_n354_), .C(ori_ori_n337_), .D(ori_ori_n332_), .Y(ori13));
  NA3        o341(.A(k), .B(j), .C(i), .Y(ori_ori_n370_));
  NO2        o342(.A(f), .B(c), .Y(ori_ori_n371_));
  OR2        o343(.A(m), .B(i), .Y(ori_ori_n372_));
  AN3        o344(.A(g), .B(f), .C(c), .Y(ori_ori_n373_));
  NA2        o345(.A(i), .B(h), .Y(ori_ori_n374_));
  NO2        o346(.A(n), .B(f), .Y(ori_ori_n375_));
  NO2        o347(.A(ori_ori_n117_), .B(a), .Y(ori_ori_n376_));
  NA2        o348(.A(ori_ori_n172_), .B(ori_ori_n468_), .Y(ori_ori_n377_));
  NA2        o349(.A(ori_ori_n214_), .B(ori_ori_n376_), .Y(ori_ori_n378_));
  NA2        o350(.A(ori_ori_n378_), .B(ori_ori_n377_), .Y(ori00));
  OAI210     o351(.A0(ori_ori_n356_), .A1(ori_ori_n32_), .B0(ori_ori_n235_), .Y(ori_ori_n380_));
  NA2        o352(.A(ori_ori_n380_), .B(n), .Y(ori_ori_n381_));
  AOI210     o353(.A0(ori_ori_n381_), .A1(ori_ori_n465_), .B0(b), .Y(ori_ori_n382_));
  INV        o354(.A(ori_ori_n382_), .Y(ori_ori_n383_));
  NA3        o355(.A(d), .B(ori_ori_n37_), .C(b), .Y(ori_ori_n384_));
  NA2        o356(.A(ori_ori_n156_), .B(ori_ori_n89_), .Y(ori_ori_n385_));
  OR2        o357(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n386_));
  INV        o358(.A(ori_ori_n224_), .Y(ori_ori_n387_));
  AN3        o359(.A(ori_ori_n387_), .B(ori_ori_n386_), .C(ori_ori_n222_), .Y(ori_ori_n388_));
  NA3        o360(.A(ori_ori_n236_), .B(ori_ori_n89_), .C(ori_ori_n61_), .Y(ori_ori_n389_));
  INV        o361(.A(ori_ori_n389_), .Y(ori_ori_n390_));
  AOI220     o362(.A0(ori_ori_n333_), .A1(ori_ori_n221_), .B0(ori_ori_n236_), .B1(ori_ori_n103_), .Y(ori_ori_n391_));
  INV        o363(.A(ori_ori_n391_), .Y(ori_ori_n392_));
  NO2        o364(.A(ori_ori_n392_), .B(ori_ori_n390_), .Y(ori_ori_n393_));
  NA3        o365(.A(ori_ori_n393_), .B(ori_ori_n388_), .C(ori_ori_n383_), .Y(ori01));
  INV        o366(.A(ori_ori_n116_), .Y(ori_ori_n395_));
  NA3        o367(.A(ori_ori_n164_), .B(ori_ori_n395_), .C(ori_ori_n364_), .Y(ori_ori_n396_));
  NA2        o368(.A(ori_ori_n216_), .B(ori_ori_n113_), .Y(ori_ori_n397_));
  NA2        o369(.A(ori_ori_n336_), .B(ori_ori_n397_), .Y(ori_ori_n398_));
  NA2        o370(.A(ori_ori_n398_), .B(ori_ori_n312_), .Y(ori_ori_n399_));
  NA2        o371(.A(ori_ori_n389_), .B(ori_ori_n308_), .Y(ori_ori_n400_));
  NO2        o372(.A(ori_ori_n251_), .B(ori_ori_n209_), .Y(ori_ori_n401_));
  INV        o373(.A(ori_ori_n401_), .Y(ori_ori_n402_));
  NO4        o374(.A(ori_ori_n402_), .B(ori_ori_n400_), .C(ori_ori_n399_), .D(ori_ori_n396_), .Y(ori_ori_n403_));
  INV        o375(.A(ori_ori_n115_), .Y(ori_ori_n404_));
  NA2        o376(.A(ori_ori_n404_), .B(ori_ori_n247_), .Y(ori_ori_n405_));
  NO2        o377(.A(ori_ori_n339_), .B(ori_ori_n95_), .Y(ori_ori_n406_));
  NO2        o378(.A(ori_ori_n340_), .B(ori_ori_n218_), .Y(ori_ori_n407_));
  OAI210     o379(.A0(ori_ori_n407_), .A1(ori_ori_n406_), .B0(ori_ori_n143_), .Y(ori_ori_n408_));
  OR2        o380(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n409_));
  INV        o381(.A(ori_ori_n409_), .Y(ori_ori_n410_));
  NOi21      o382(.An(ori_ori_n408_), .B(ori_ori_n410_), .Y(ori_ori_n411_));
  NO2        o383(.A(ori_ori_n374_), .B(m), .Y(ori_ori_n412_));
  NO2        o384(.A(ori_ori_n229_), .B(ori_ori_n228_), .Y(ori_ori_n413_));
  NO3        o385(.A(ori_ori_n374_), .B(ori_ori_n413_), .C(ori_ori_n65_), .Y(ori_ori_n414_));
  INV        o386(.A(ori_ori_n414_), .Y(ori_ori_n415_));
  NA4        o387(.A(ori_ori_n415_), .B(ori_ori_n411_), .C(ori_ori_n405_), .D(ori_ori_n403_), .Y(ori06));
  OAI210     o388(.A0(n), .A1(ori_ori_n412_), .B0(ori_ori_n155_), .Y(ori_ori_n417_));
  NA2        o389(.A(ori_ori_n417_), .B(ori_ori_n408_), .Y(ori_ori_n418_));
  NO2        o390(.A(ori_ori_n418_), .B(ori_ori_n111_), .Y(ori_ori_n419_));
  NO2        o391(.A(ori_ori_n121_), .B(ori_ori_n33_), .Y(ori_ori_n420_));
  AOI210     o392(.A0(ori_ori_n420_), .A1(ori_ori_n215_), .B0(ori_ori_n406_), .Y(ori_ori_n421_));
  AOI210     o393(.A0(ori_ori_n420_), .A1(ori_ori_n219_), .B0(ori_ori_n234_), .Y(ori_ori_n422_));
  AOI210     o394(.A0(ori_ori_n422_), .A1(ori_ori_n421_), .B0(ori_ori_n140_), .Y(ori_ori_n423_));
  INV        o395(.A(ori_ori_n250_), .Y(ori_ori_n424_));
  NA2        o396(.A(ori_ori_n424_), .B(ori_ori_n149_), .Y(ori_ori_n425_));
  INV        o397(.A(ori_ori_n425_), .Y(ori_ori_n426_));
  NO2        o398(.A(ori_ori_n426_), .B(ori_ori_n423_), .Y(ori_ori_n427_));
  AN2        o399(.A(ori_ori_n318_), .B(ori_ori_n317_), .Y(ori_ori_n428_));
  NO2        o400(.A(ori_ori_n428_), .B(ori_ori_n195_), .Y(ori_ori_n429_));
  INV        o401(.A(ori_ori_n429_), .Y(ori_ori_n430_));
  INV        o402(.A(i), .Y(ori_ori_n431_));
  NO4        o403(.A(ori_ori_n413_), .B(ori_ori_n431_), .C(ori_ori_n177_), .D(ori_ori_n97_), .Y(ori_ori_n432_));
  NO3        o404(.A(ori_ori_n432_), .B(ori_ori_n430_), .C(ori_ori_n467_), .Y(ori_ori_n433_));
  NA4        o405(.A(ori_ori_n433_), .B(ori_ori_n427_), .C(ori_ori_n419_), .D(ori_ori_n415_), .Y(ori07));
  NO2        o406(.A(m), .B(h), .Y(ori_ori_n435_));
  NO2        o407(.A(ori_ori_n370_), .B(ori_ori_n122_), .Y(ori_ori_n436_));
  NO2        o408(.A(l), .B(k), .Y(ori_ori_n437_));
  NO3        o409(.A(ori_ori_n177_), .B(d), .C(c), .Y(ori_ori_n438_));
  NA2        o410(.A(ori_ori_n373_), .B(ori_ori_n194_), .Y(ori_ori_n439_));
  NA2        o411(.A(ori_ori_n435_), .B(ori_ori_n437_), .Y(ori_ori_n440_));
  INV        o412(.A(ori_ori_n440_), .Y(ori_ori_n441_));
  NA2        o413(.A(ori_ori_n375_), .B(ori_ori_n170_), .Y(ori_ori_n442_));
  NO2        o414(.A(ori_ori_n442_), .B(ori_ori_n176_), .Y(ori_ori_n443_));
  OR2        o415(.A(ori_ori_n443_), .B(ori_ori_n441_), .Y(ori_ori_n444_));
  NO2        o416(.A(ori_ori_n444_), .B(ori_ori_n464_), .Y(ori_ori_n445_));
  NA3        o417(.A(ori_ori_n445_), .B(ori_ori_n439_), .C(ori_ori_n35_), .Y(ori_ori_n446_));
  NO2        o418(.A(ori_ori_n162_), .B(j), .Y(ori_ori_n447_));
  NA2        o419(.A(ori_ori_n371_), .B(ori_ori_n55_), .Y(ori_ori_n448_));
  INV        o420(.A(ori_ori_n448_), .Y(ori_ori_n449_));
  NA2        o421(.A(ori_ori_n447_), .B(h), .Y(ori_ori_n450_));
  INV        o422(.A(ori_ori_n450_), .Y(ori_ori_n451_));
  NO2        o423(.A(ori_ori_n451_), .B(ori_ori_n449_), .Y(ori_ori_n452_));
  NO2        o424(.A(ori_ori_n372_), .B(h), .Y(ori_ori_n453_));
  NA2        o425(.A(ori_ori_n466_), .B(ori_ori_n452_), .Y(ori_ori_n454_));
  NA2        o426(.A(h), .B(ori_ori_n436_), .Y(ori_ori_n455_));
  OR2        o427(.A(h), .B(ori_ori_n213_), .Y(ori_ori_n456_));
  NO2        o428(.A(ori_ori_n456_), .B(ori_ori_n65_), .Y(ori_ori_n457_));
  NO2        o429(.A(ori_ori_n457_), .B(ori_ori_n438_), .Y(ori_ori_n458_));
  NA2        o430(.A(ori_ori_n458_), .B(ori_ori_n455_), .Y(ori_ori_n459_));
  OR3        o431(.A(ori_ori_n459_), .B(ori_ori_n454_), .C(ori_ori_n446_), .Y(ori04));
  INV        o432(.A(ori_ori_n124_), .Y(ori_ori_n463_));
  INV        o433(.A(ori_ori_n52_), .Y(ori_ori_n464_));
  INV        o434(.A(ori_ori_n120_), .Y(ori_ori_n465_));
  INV        o435(.A(ori_ori_n453_), .Y(ori_ori_n466_));
  INV        o436(.A(ori_ori_n391_), .Y(ori_ori_n467_));
  INV        o437(.A(a), .Y(ori_ori_n468_));
  INV        o438(.A(m), .Y(ori_ori_n469_));
  ZERO       o439(.Y(ori02));
  ZERO       o440(.Y(ori03));
  ZERO       o441(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(i), .Bn(g), .C(h), .Y(mai_mai_n33_));
  NA2        m0005(.A(mai_mai_n33_), .B(m), .Y(mai_mai_n34_));
  AN2        m0006(.A(m), .B(l), .Y(mai_mai_n35_));
  NOi32      m0007(.An(j), .Bn(g), .C(k), .Y(mai_mai_n36_));
  NA2        m0008(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n37_));
  NO2        m0009(.A(mai_mai_n37_), .B(n), .Y(mai_mai_n38_));
  INV        m0010(.A(h), .Y(mai_mai_n39_));
  NAi21      m0011(.An(j), .B(l), .Y(mai_mai_n40_));
  INV        m0012(.A(i), .Y(mai_mai_n41_));
  AN2        m0013(.A(h), .B(g), .Y(mai_mai_n42_));
  NAi21      m0014(.An(n), .B(m), .Y(mai_mai_n43_));
  NOi32      m0015(.An(k), .Bn(h), .C(l), .Y(mai_mai_n44_));
  NOi32      m0016(.An(k), .Bn(h), .C(g), .Y(mai_mai_n45_));
  INV        m0017(.A(mai_mai_n45_), .Y(mai_mai_n46_));
  NO2        m0018(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n43_), .B(mai_mai_n32_), .Y(mai_mai_n48_));
  INV        m0020(.A(c), .Y(mai_mai_n49_));
  NA2        m0021(.A(e), .B(b), .Y(mai_mai_n50_));
  NO2        m0022(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n51_));
  INV        m0023(.A(d), .Y(mai_mai_n52_));
  NAi21      m0024(.An(i), .B(h), .Y(mai_mai_n53_));
  NAi21      m0025(.An(i), .B(j), .Y(mai_mai_n54_));
  NAi32      m0026(.An(n), .Bn(k), .C(m), .Y(mai_mai_n55_));
  NAi31      m0027(.An(l), .B(m), .C(k), .Y(mai_mai_n56_));
  NAi21      m0028(.An(e), .B(h), .Y(mai_mai_n57_));
  NAi41      m0029(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n58_));
  INV        m0030(.A(m), .Y(mai_mai_n59_));
  NOi21      m0031(.An(k), .B(l), .Y(mai_mai_n60_));
  AN4        m0032(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n61_));
  NOi31      m0033(.An(h), .B(g), .C(f), .Y(mai_mai_n62_));
  NA2        m0034(.A(mai_mai_n62_), .B(mai_mai_n61_), .Y(mai_mai_n63_));
  NAi32      m0035(.An(m), .Bn(k), .C(j), .Y(mai_mai_n64_));
  NOi32      m0036(.An(h), .Bn(g), .C(f), .Y(mai_mai_n65_));
  NA2        m0037(.A(mai_mai_n65_), .B(mai_mai_n61_), .Y(mai_mai_n66_));
  OA220      m0038(.A0(mai_mai_n66_), .A1(mai_mai_n64_), .B0(mai_mai_n63_), .B1(l), .Y(mai_mai_n67_));
  INV        m0039(.A(mai_mai_n67_), .Y(mai_mai_n68_));
  INV        m0040(.A(n), .Y(mai_mai_n69_));
  NOi32      m0041(.An(e), .Bn(b), .C(d), .Y(mai_mai_n70_));
  INV        m0042(.A(j), .Y(mai_mai_n71_));
  AN3        m0043(.A(m), .B(k), .C(i), .Y(mai_mai_n72_));
  NAi32      m0044(.An(g), .Bn(f), .C(h), .Y(mai_mai_n73_));
  NAi31      m0045(.An(j), .B(m), .C(l), .Y(mai_mai_n74_));
  NO2        m0046(.A(mai_mai_n74_), .B(mai_mai_n73_), .Y(mai_mai_n75_));
  NA2        m0047(.A(m), .B(l), .Y(mai_mai_n76_));
  NO2        m0048(.A(mai_mai_n76_), .B(f), .Y(mai_mai_n77_));
  NOi32      m0049(.An(m), .Bn(l), .C(i), .Y(mai_mai_n78_));
  NOi21      m0050(.An(g), .B(i), .Y(mai_mai_n79_));
  NAi41      m0051(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n80_));
  AN2        m0052(.A(e), .B(b), .Y(mai_mai_n81_));
  NOi31      m0053(.An(c), .B(h), .C(f), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n83_));
  NOi21      m0055(.An(i), .B(h), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(g), .C(mai_mai_n35_), .Y(mai_mai_n85_));
  INV        m0057(.A(a), .Y(mai_mai_n86_));
  INV        m0058(.A(mai_mai_n81_), .Y(mai_mai_n87_));
  INV        m0059(.A(l), .Y(mai_mai_n88_));
  NOi21      m0060(.An(m), .B(n), .Y(mai_mai_n89_));
  AN2        m0061(.A(k), .B(h), .Y(mai_mai_n90_));
  INV        m0062(.A(mai_mai_n85_), .Y(mai_mai_n91_));
  INV        m0063(.A(b), .Y(mai_mai_n92_));
  NA2        m0064(.A(l), .B(j), .Y(mai_mai_n93_));
  NOi32      m0065(.An(c), .Bn(a), .C(d), .Y(mai_mai_n94_));
  NOi31      m0066(.An(k), .B(m), .C(j), .Y(mai_mai_n95_));
  NOi31      m0067(.An(k), .B(m), .C(i), .Y(mai_mai_n96_));
  NA3        m0068(.A(mai_mai_n96_), .B(mai_mai_n65_), .C(mai_mai_n61_), .Y(mai_mai_n97_));
  INV        m0069(.A(mai_mai_n97_), .Y(mai_mai_n98_));
  NOi32      m0070(.An(f), .Bn(b), .C(e), .Y(mai_mai_n99_));
  NAi21      m0071(.An(g), .B(h), .Y(mai_mai_n100_));
  NAi21      m0072(.An(m), .B(n), .Y(mai_mai_n101_));
  NAi21      m0073(.An(j), .B(k), .Y(mai_mai_n102_));
  NO3        m0074(.A(mai_mai_n102_), .B(mai_mai_n101_), .C(mai_mai_n100_), .Y(mai_mai_n103_));
  NAi41      m0075(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n104_));
  NAi31      m0076(.An(j), .B(k), .C(h), .Y(mai_mai_n105_));
  NO3        m0077(.A(mai_mai_n105_), .B(mai_mai_n104_), .C(mai_mai_n101_), .Y(mai_mai_n106_));
  AOI210     m0078(.A0(mai_mai_n103_), .A1(mai_mai_n99_), .B0(mai_mai_n106_), .Y(mai_mai_n107_));
  NO2        m0079(.A(k), .B(j), .Y(mai_mai_n108_));
  NO2        m0080(.A(mai_mai_n108_), .B(mai_mai_n101_), .Y(mai_mai_n109_));
  AN2        m0081(.A(k), .B(j), .Y(mai_mai_n110_));
  NAi21      m0082(.An(c), .B(b), .Y(mai_mai_n111_));
  NA2        m0083(.A(f), .B(d), .Y(mai_mai_n112_));
  NO4        m0084(.A(mai_mai_n112_), .B(mai_mai_n111_), .C(mai_mai_n110_), .D(mai_mai_n100_), .Y(mai_mai_n113_));
  NA2        m0085(.A(h), .B(c), .Y(mai_mai_n114_));
  NAi31      m0086(.An(f), .B(e), .C(b), .Y(mai_mai_n115_));
  NA2        m0087(.A(mai_mai_n113_), .B(mai_mai_n109_), .Y(mai_mai_n116_));
  NA2        m0088(.A(d), .B(b), .Y(mai_mai_n117_));
  NAi21      m0089(.An(e), .B(f), .Y(mai_mai_n118_));
  NO2        m0090(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n119_));
  NA2        m0091(.A(b), .B(a), .Y(mai_mai_n120_));
  NAi21      m0092(.An(c), .B(d), .Y(mai_mai_n121_));
  NAi31      m0093(.An(l), .B(k), .C(h), .Y(mai_mai_n122_));
  NO2        m0094(.A(mai_mai_n101_), .B(mai_mai_n122_), .Y(mai_mai_n123_));
  NA2        m0095(.A(mai_mai_n123_), .B(mai_mai_n119_), .Y(mai_mai_n124_));
  NAi41      m0096(.An(mai_mai_n98_), .B(mai_mai_n124_), .C(mai_mai_n116_), .D(mai_mai_n107_), .Y(mai_mai_n125_));
  NAi31      m0097(.An(e), .B(f), .C(b), .Y(mai_mai_n126_));
  NOi21      m0098(.An(g), .B(d), .Y(mai_mai_n127_));
  NO2        m0099(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n128_));
  NOi21      m0100(.An(h), .B(i), .Y(mai_mai_n129_));
  NOi21      m0101(.An(k), .B(m), .Y(mai_mai_n130_));
  NA3        m0102(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(n), .Y(mai_mai_n131_));
  NOi21      m0103(.An(mai_mai_n128_), .B(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m0104(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n133_));
  NA2        m0105(.A(mai_mai_n133_), .B(h), .Y(mai_mai_n134_));
  NOi32      m0106(.An(n), .Bn(k), .C(m), .Y(mai_mai_n135_));
  NA2        m0107(.A(l), .B(i), .Y(mai_mai_n136_));
  NA2        m0108(.A(mai_mai_n136_), .B(mai_mai_n135_), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n137_), .B(mai_mai_n134_), .Y(mai_mai_n138_));
  NAi31      m0110(.An(d), .B(f), .C(c), .Y(mai_mai_n139_));
  NAi31      m0111(.An(e), .B(f), .C(c), .Y(mai_mai_n140_));
  NA2        m0112(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n141_));
  NA2        m0113(.A(j), .B(h), .Y(mai_mai_n142_));
  OR3        m0114(.A(n), .B(m), .C(k), .Y(mai_mai_n143_));
  NO2        m0115(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NAi32      m0116(.An(m), .Bn(k), .C(n), .Y(mai_mai_n145_));
  NO2        m0117(.A(mai_mai_n145_), .B(mai_mai_n142_), .Y(mai_mai_n146_));
  AOI220     m0118(.A0(mai_mai_n146_), .A1(mai_mai_n128_), .B0(mai_mai_n144_), .B1(mai_mai_n141_), .Y(mai_mai_n147_));
  NO2        m0119(.A(n), .B(m), .Y(mai_mai_n148_));
  NA2        m0120(.A(mai_mai_n148_), .B(mai_mai_n44_), .Y(mai_mai_n149_));
  NAi21      m0121(.An(f), .B(e), .Y(mai_mai_n150_));
  NA2        m0122(.A(d), .B(c), .Y(mai_mai_n151_));
  NAi31      m0123(.An(m), .B(n), .C(b), .Y(mai_mai_n152_));
  NA2        m0124(.A(k), .B(i), .Y(mai_mai_n153_));
  NAi21      m0125(.An(h), .B(f), .Y(mai_mai_n154_));
  NO2        m0126(.A(mai_mai_n152_), .B(mai_mai_n121_), .Y(mai_mai_n155_));
  NOi32      m0127(.An(f), .Bn(c), .C(d), .Y(mai_mai_n156_));
  NOi32      m0128(.An(f), .Bn(c), .C(e), .Y(mai_mai_n157_));
  NO2        m0129(.A(mai_mai_n157_), .B(mai_mai_n156_), .Y(mai_mai_n158_));
  NO3        m0130(.A(n), .B(m), .C(j), .Y(mai_mai_n159_));
  NA2        m0131(.A(mai_mai_n159_), .B(mai_mai_n90_), .Y(mai_mai_n160_));
  AO210      m0132(.A0(mai_mai_n160_), .A1(mai_mai_n149_), .B0(mai_mai_n158_), .Y(mai_mai_n161_));
  NA2        m0133(.A(mai_mai_n161_), .B(mai_mai_n147_), .Y(mai_mai_n162_));
  OR4        m0134(.A(mai_mai_n162_), .B(mai_mai_n138_), .C(mai_mai_n132_), .D(mai_mai_n125_), .Y(mai_mai_n163_));
  NO4        m0135(.A(mai_mai_n163_), .B(mai_mai_n91_), .C(mai_mai_n68_), .D(mai_mai_n48_), .Y(mai_mai_n164_));
  NA3        m0136(.A(m), .B(mai_mai_n88_), .C(j), .Y(mai_mai_n165_));
  NAi31      m0137(.An(n), .B(h), .C(g), .Y(mai_mai_n166_));
  NO2        m0138(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  NOi32      m0139(.An(m), .Bn(k), .C(l), .Y(mai_mai_n168_));
  NA3        m0140(.A(mai_mai_n168_), .B(mai_mai_n71_), .C(g), .Y(mai_mai_n169_));
  AN2        m0141(.A(i), .B(g), .Y(mai_mai_n170_));
  NA3        m0142(.A(mai_mai_n60_), .B(mai_mai_n170_), .C(mai_mai_n89_), .Y(mai_mai_n171_));
  NAi41      m0143(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n172_));
  INV        m0144(.A(mai_mai_n172_), .Y(mai_mai_n173_));
  INV        m0145(.A(f), .Y(mai_mai_n174_));
  INV        m0146(.A(g), .Y(mai_mai_n175_));
  NOi31      m0147(.An(i), .B(j), .C(h), .Y(mai_mai_n176_));
  NOi21      m0148(.An(l), .B(m), .Y(mai_mai_n177_));
  NA2        m0149(.A(mai_mai_n177_), .B(mai_mai_n176_), .Y(mai_mai_n178_));
  NO3        m0150(.A(mai_mai_n178_), .B(mai_mai_n175_), .C(mai_mai_n174_), .Y(mai_mai_n179_));
  NA2        m0151(.A(mai_mai_n179_), .B(mai_mai_n173_), .Y(mai_mai_n180_));
  INV        m0152(.A(mai_mai_n180_), .Y(mai_mai_n181_));
  NOi21      m0153(.An(n), .B(m), .Y(mai_mai_n182_));
  NOi32      m0154(.An(l), .Bn(i), .C(j), .Y(mai_mai_n183_));
  NA2        m0155(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  OA220      m0156(.A0(mai_mai_n184_), .A1(mai_mai_n83_), .B0(mai_mai_n64_), .B1(mai_mai_n63_), .Y(mai_mai_n185_));
  NAi21      m0157(.An(j), .B(h), .Y(mai_mai_n186_));
  XN2        m0158(.A(i), .B(h), .Y(mai_mai_n187_));
  NA2        m0159(.A(mai_mai_n187_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  NOi31      m0160(.An(k), .B(n), .C(m), .Y(mai_mai_n189_));
  NOi31      m0161(.An(mai_mai_n189_), .B(mai_mai_n151_), .C(mai_mai_n150_), .Y(mai_mai_n190_));
  NA2        m0162(.A(mai_mai_n190_), .B(mai_mai_n188_), .Y(mai_mai_n191_));
  NAi31      m0163(.An(f), .B(e), .C(c), .Y(mai_mai_n192_));
  NO4        m0164(.A(mai_mai_n192_), .B(mai_mai_n143_), .C(mai_mai_n142_), .D(mai_mai_n52_), .Y(mai_mai_n193_));
  NA4        m0165(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n194_));
  NAi32      m0166(.An(m), .Bn(i), .C(k), .Y(mai_mai_n195_));
  NO3        m0167(.A(mai_mai_n195_), .B(mai_mai_n73_), .C(mai_mai_n194_), .Y(mai_mai_n196_));
  INV        m0168(.A(k), .Y(mai_mai_n197_));
  NO2        m0169(.A(mai_mai_n196_), .B(mai_mai_n193_), .Y(mai_mai_n198_));
  NAi21      m0170(.An(n), .B(a), .Y(mai_mai_n199_));
  NO2        m0171(.A(mai_mai_n199_), .B(mai_mai_n117_), .Y(mai_mai_n200_));
  NAi41      m0172(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n201_));
  NO2        m0173(.A(mai_mai_n201_), .B(e), .Y(mai_mai_n202_));
  NA2        m0174(.A(mai_mai_n202_), .B(mai_mai_n200_), .Y(mai_mai_n203_));
  AN4        m0175(.A(mai_mai_n203_), .B(mai_mai_n198_), .C(mai_mai_n191_), .D(mai_mai_n185_), .Y(mai_mai_n204_));
  NAi41      m0176(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n205_));
  NO2        m0177(.A(mai_mai_n205_), .B(mai_mai_n174_), .Y(mai_mai_n206_));
  NA2        m0178(.A(mai_mai_n130_), .B(mai_mai_n84_), .Y(mai_mai_n207_));
  NAi21      m0179(.An(mai_mai_n207_), .B(mai_mai_n206_), .Y(mai_mai_n208_));
  NO2        m0180(.A(n), .B(a), .Y(mai_mai_n209_));
  NAi21      m0181(.An(h), .B(i), .Y(mai_mai_n210_));
  NA2        m0182(.A(mai_mai_n148_), .B(k), .Y(mai_mai_n211_));
  NO2        m0183(.A(mai_mai_n211_), .B(mai_mai_n210_), .Y(mai_mai_n212_));
  NA2        m0184(.A(mai_mai_n212_), .B(mai_mai_n156_), .Y(mai_mai_n213_));
  NA2        m0185(.A(mai_mai_n213_), .B(mai_mai_n208_), .Y(mai_mai_n214_));
  NOi21      m0186(.An(g), .B(e), .Y(mai_mai_n215_));
  NO2        m0187(.A(mai_mai_n58_), .B(mai_mai_n59_), .Y(mai_mai_n216_));
  NA2        m0188(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  INV        m0189(.A(mai_mai_n55_), .Y(mai_mai_n218_));
  INV        m0190(.A(mai_mai_n217_), .Y(mai_mai_n219_));
  NOi41      m0191(.An(mai_mai_n204_), .B(mai_mai_n219_), .C(mai_mai_n214_), .D(mai_mai_n181_), .Y(mai_mai_n220_));
  NO2        m0192(.A(mai_mai_n167_), .B(mai_mai_n38_), .Y(mai_mai_n221_));
  NO2        m0193(.A(mai_mai_n221_), .B(mai_mai_n87_), .Y(mai_mai_n222_));
  NA3        m0194(.A(mai_mai_n52_), .B(c), .C(b), .Y(mai_mai_n223_));
  NAi21      m0195(.An(h), .B(g), .Y(mai_mai_n224_));
  OR4        m0196(.A(mai_mai_n224_), .B(mai_mai_n223_), .C(mai_mai_n184_), .D(e), .Y(mai_mai_n225_));
  NO2        m0197(.A(mai_mai_n207_), .B(f), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n226_), .B(mai_mai_n61_), .Y(mai_mai_n227_));
  NAi31      m0199(.An(e), .B(d), .C(a), .Y(mai_mai_n228_));
  NA2        m0200(.A(mai_mai_n227_), .B(mai_mai_n225_), .Y(mai_mai_n229_));
  NA4        m0201(.A(mai_mai_n130_), .B(mai_mai_n65_), .C(mai_mai_n61_), .D(mai_mai_n93_), .Y(mai_mai_n230_));
  NA3        m0202(.A(mai_mai_n130_), .B(mai_mai_n129_), .C(mai_mai_n69_), .Y(mai_mai_n231_));
  NO2        m0203(.A(mai_mai_n231_), .B(mai_mai_n158_), .Y(mai_mai_n232_));
  NOi21      m0204(.An(mai_mai_n230_), .B(mai_mai_n232_), .Y(mai_mai_n233_));
  NA3        m0205(.A(e), .B(c), .C(b), .Y(mai_mai_n234_));
  INV        m0206(.A(mai_mai_n43_), .Y(mai_mai_n235_));
  NOi21      m0207(.An(l), .B(j), .Y(mai_mai_n236_));
  OR3        m0208(.A(mai_mai_n58_), .B(mai_mai_n59_), .C(e), .Y(mai_mai_n237_));
  NO2        m0209(.A(j), .B(mai_mai_n237_), .Y(mai_mai_n238_));
  INV        m0210(.A(mai_mai_n238_), .Y(mai_mai_n239_));
  NAi32      m0211(.An(j), .Bn(h), .C(i), .Y(mai_mai_n240_));
  NAi21      m0212(.An(m), .B(l), .Y(mai_mai_n241_));
  NO2        m0213(.A(mai_mai_n240_), .B(mai_mai_n69_), .Y(mai_mai_n242_));
  NA2        m0214(.A(h), .B(g), .Y(mai_mai_n243_));
  NA2        m0215(.A(mai_mai_n135_), .B(mai_mai_n41_), .Y(mai_mai_n244_));
  NA2        m0216(.A(mai_mai_n242_), .B(mai_mai_n133_), .Y(mai_mai_n245_));
  NA3        m0217(.A(mai_mai_n245_), .B(mai_mai_n239_), .C(mai_mai_n233_), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n115_), .B(d), .Y(mai_mai_n247_));
  NO2        m0219(.A(mai_mai_n83_), .B(mai_mai_n80_), .Y(mai_mai_n248_));
  NAi32      m0220(.An(n), .Bn(m), .C(l), .Y(mai_mai_n249_));
  NO4        m0221(.A(mai_mai_n47_), .B(mai_mai_n246_), .C(mai_mai_n229_), .D(mai_mai_n222_), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n212_), .B(mai_mai_n157_), .Y(mai_mai_n251_));
  NAi21      m0223(.An(m), .B(k), .Y(mai_mai_n252_));
  NO2        m0224(.A(mai_mai_n187_), .B(mai_mai_n252_), .Y(mai_mai_n253_));
  NAi41      m0225(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n254_));
  NA2        m0226(.A(e), .B(c), .Y(mai_mai_n255_));
  NO3        m0227(.A(mai_mai_n255_), .B(n), .C(d), .Y(mai_mai_n256_));
  NA2        m0228(.A(f), .B(k), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n175_), .Y(mai_mai_n258_));
  NAi31      m0230(.An(d), .B(e), .C(b), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n101_), .B(mai_mai_n259_), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n260_), .B(mai_mai_n258_), .Y(mai_mai_n261_));
  NA2        m0233(.A(mai_mai_n261_), .B(mai_mai_n251_), .Y(mai_mai_n262_));
  NO4        m0234(.A(mai_mai_n254_), .B(mai_mai_n64_), .C(mai_mai_n57_), .D(mai_mai_n175_), .Y(mai_mai_n263_));
  NA2        m0235(.A(mai_mai_n209_), .B(mai_mai_n81_), .Y(mai_mai_n264_));
  OR2        m0236(.A(mai_mai_n264_), .B(mai_mai_n169_), .Y(mai_mai_n265_));
  NOi31      m0237(.An(l), .B(n), .C(m), .Y(mai_mai_n266_));
  BUFFER     m0238(.A(mai_mai_n263_), .Y(mai_mai_n267_));
  NAi32      m0239(.An(m), .Bn(j), .C(k), .Y(mai_mai_n268_));
  NAi41      m0240(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n269_));
  NOi31      m0241(.An(j), .B(m), .C(k), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n95_), .B(mai_mai_n270_), .Y(mai_mai_n271_));
  AN3        m0243(.A(h), .B(g), .C(f), .Y(mai_mai_n272_));
  NOi32      m0244(.An(m), .Bn(j), .C(l), .Y(mai_mai_n273_));
  INV        m0245(.A(mai_mai_n273_), .Y(mai_mai_n274_));
  NO2        m0246(.A(mai_mai_n241_), .B(mai_mai_n240_), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n178_), .B(g), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n126_), .B(mai_mai_n69_), .Y(mai_mai_n277_));
  AOI220     m0249(.A0(mai_mai_n277_), .A1(mai_mai_n276_), .B0(mai_mai_n206_), .B1(mai_mai_n275_), .Y(mai_mai_n278_));
  NA2        m0250(.A(mai_mai_n272_), .B(mai_mai_n173_), .Y(mai_mai_n279_));
  NA2        m0251(.A(mai_mai_n279_), .B(mai_mai_n278_), .Y(mai_mai_n280_));
  NA3        m0252(.A(h), .B(g), .C(f), .Y(mai_mai_n281_));
  NA2        m0253(.A(h), .B(e), .Y(mai_mai_n282_));
  NO2        m0254(.A(mai_mai_n282_), .B(mai_mai_n40_), .Y(mai_mai_n283_));
  NA2        m0255(.A(mai_mai_n283_), .B(mai_mai_n89_), .Y(mai_mai_n284_));
  NOi32      m0256(.An(j), .Bn(g), .C(i), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n285_), .B(mai_mai_n89_), .Y(mai_mai_n286_));
  BUFFER     m0258(.A(mai_mai_n286_), .Y(mai_mai_n287_));
  NOi32      m0259(.An(e), .Bn(b), .C(a), .Y(mai_mai_n288_));
  NO3        m0260(.A(mai_mai_n254_), .B(mai_mai_n57_), .C(mai_mai_n175_), .Y(mai_mai_n289_));
  NA2        m0261(.A(mai_mai_n171_), .B(mai_mai_n34_), .Y(mai_mai_n290_));
  AOI220     m0262(.A0(mai_mai_n290_), .A1(mai_mai_n288_), .B0(mai_mai_n289_), .B1(k), .Y(mai_mai_n291_));
  INV        m0263(.A(n), .Y(mai_mai_n292_));
  NA2        m0264(.A(mai_mai_n170_), .B(k), .Y(mai_mai_n293_));
  NA3        m0265(.A(m), .B(mai_mai_n88_), .C(mai_mai_n174_), .Y(mai_mai_n294_));
  NA4        m0266(.A(mai_mai_n168_), .B(mai_mai_n71_), .C(g), .D(mai_mai_n174_), .Y(mai_mai_n295_));
  NAi41      m0267(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n45_), .B(mai_mai_n89_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  AOI220     m0270(.A0(mai_mai_n298_), .A1(b), .B0(mai_mai_n168_), .B1(mai_mai_n292_), .Y(mai_mai_n299_));
  NA4        m0271(.A(mai_mai_n299_), .B(mai_mai_n291_), .C(mai_mai_n287_), .D(mai_mai_n284_), .Y(mai_mai_n300_));
  NO4        m0272(.A(mai_mai_n300_), .B(mai_mai_n280_), .C(mai_mai_n267_), .D(mai_mai_n262_), .Y(mai_mai_n301_));
  NA4        m0273(.A(mai_mai_n301_), .B(mai_mai_n250_), .C(mai_mai_n220_), .D(mai_mai_n164_), .Y(mai10));
  NA3        m0274(.A(m), .B(k), .C(i), .Y(mai_mai_n303_));
  NO3        m0275(.A(mai_mai_n303_), .B(j), .C(mai_mai_n175_), .Y(mai_mai_n304_));
  NOi21      m0276(.An(e), .B(f), .Y(mai_mai_n305_));
  NO3        m0277(.A(mai_mai_n121_), .B(n), .C(mai_mai_n86_), .Y(mai_mai_n306_));
  NAi31      m0278(.An(b), .B(f), .C(c), .Y(mai_mai_n307_));
  INV        m0279(.A(mai_mai_n307_), .Y(mai_mai_n308_));
  NOi32      m0280(.An(k), .Bn(h), .C(j), .Y(mai_mai_n309_));
  NA2        m0281(.A(mai_mai_n309_), .B(mai_mai_n182_), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n131_), .B(mai_mai_n310_), .Y(mai_mai_n311_));
  AOI220     m0283(.A0(mai_mai_n311_), .A1(mai_mai_n308_), .B0(mai_mai_n306_), .B1(mai_mai_n304_), .Y(mai_mai_n312_));
  AN2        m0284(.A(j), .B(h), .Y(mai_mai_n313_));
  NO3        m0285(.A(n), .B(m), .C(k), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n314_), .B(mai_mai_n313_), .Y(mai_mai_n315_));
  NO3        m0287(.A(mai_mai_n315_), .B(mai_mai_n121_), .C(mai_mai_n174_), .Y(mai_mai_n316_));
  OR2        m0288(.A(m), .B(k), .Y(mai_mai_n317_));
  NO2        m0289(.A(mai_mai_n142_), .B(mai_mai_n317_), .Y(mai_mai_n318_));
  NA4        m0290(.A(n), .B(f), .C(c), .D(mai_mai_n92_), .Y(mai_mai_n319_));
  NOi21      m0291(.An(mai_mai_n318_), .B(mai_mai_n319_), .Y(mai_mai_n320_));
  NOi32      m0292(.An(d), .Bn(a), .C(c), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n321_), .B(mai_mai_n150_), .Y(mai_mai_n322_));
  NAi31      m0294(.An(k), .B(m), .C(j), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n320_), .B(mai_mai_n316_), .Y(mai_mai_n324_));
  NO2        m0296(.A(mai_mai_n319_), .B(mai_mai_n241_), .Y(mai_mai_n325_));
  NOi32      m0297(.An(f), .Bn(d), .C(c), .Y(mai_mai_n326_));
  NA2        m0298(.A(mai_mai_n324_), .B(mai_mai_n312_), .Y(mai_mai_n327_));
  NA2        m0299(.A(mai_mai_n209_), .B(d), .Y(mai_mai_n328_));
  INV        m0300(.A(e), .Y(mai_mai_n329_));
  OAI220     m0301(.A0(mai_mai_n1093_), .A1(mai_mai_n165_), .B0(mai_mai_n169_), .B1(mai_mai_n329_), .Y(mai_mai_n330_));
  NA3        m0302(.A(e), .B(mai_mai_n236_), .C(m), .Y(mai_mai_n331_));
  NOi21      m0303(.An(g), .B(h), .Y(mai_mai_n332_));
  NA3        m0304(.A(m), .B(mai_mai_n332_), .C(e), .Y(mai_mai_n333_));
  AN3        m0305(.A(h), .B(g), .C(e), .Y(mai_mai_n334_));
  AN2        m0306(.A(mai_mai_n333_), .B(mai_mai_n331_), .Y(mai_mai_n335_));
  NO2        m0307(.A(mai_mai_n335_), .B(mai_mai_n328_), .Y(mai_mai_n336_));
  NA3        m0308(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(e), .Y(mai_mai_n337_));
  NA3        m0309(.A(mai_mai_n321_), .B(mai_mai_n150_), .C(mai_mai_n69_), .Y(mai_mai_n338_));
  NAi31      m0310(.An(b), .B(c), .C(a), .Y(mai_mai_n339_));
  NO2        m0311(.A(mai_mai_n339_), .B(n), .Y(mai_mai_n340_));
  NA2        m0312(.A(mai_mai_n44_), .B(m), .Y(mai_mai_n341_));
  NO2        m0313(.A(mai_mai_n336_), .B(mai_mai_n327_), .Y(mai_mai_n342_));
  NA2        m0314(.A(i), .B(g), .Y(mai_mai_n343_));
  NO3        m0315(.A(mai_mai_n228_), .B(mai_mai_n343_), .C(c), .Y(mai_mai_n344_));
  NOi21      m0316(.An(a), .B(n), .Y(mai_mai_n345_));
  NA2        m0317(.A(d), .B(mai_mai_n345_), .Y(mai_mai_n346_));
  NA3        m0318(.A(i), .B(g), .C(f), .Y(mai_mai_n347_));
  OR2        m0319(.A(mai_mai_n347_), .B(mai_mai_n56_), .Y(mai_mai_n348_));
  NA3        m0320(.A(m), .B(mai_mai_n332_), .C(mai_mai_n150_), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n349_), .B(mai_mai_n346_), .Y(mai_mai_n350_));
  AOI210     m0322(.A0(mai_mai_n344_), .A1(mai_mai_n235_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  OR2        m0323(.A(n), .B(m), .Y(mai_mai_n352_));
  NO2        m0324(.A(mai_mai_n352_), .B(mai_mai_n122_), .Y(mai_mai_n353_));
  NO2        m0325(.A(mai_mai_n151_), .B(mai_mai_n118_), .Y(mai_mai_n354_));
  OAI210     m0326(.A0(mai_mai_n353_), .A1(mai_mai_n144_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NAi21      m0327(.An(k), .B(j), .Y(mai_mai_n356_));
  NAi21      m0328(.An(e), .B(d), .Y(mai_mai_n357_));
  INV        m0329(.A(mai_mai_n357_), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n211_), .B(mai_mai_n174_), .Y(mai_mai_n359_));
  NA3        m0331(.A(mai_mai_n359_), .B(mai_mai_n358_), .C(mai_mai_n188_), .Y(mai_mai_n360_));
  NA2        m0332(.A(mai_mai_n360_), .B(mai_mai_n355_), .Y(mai_mai_n361_));
  NOi31      m0333(.An(n), .B(m), .C(k), .Y(mai_mai_n362_));
  AOI220     m0334(.A0(mai_mai_n362_), .A1(mai_mai_n313_), .B0(mai_mai_n182_), .B1(mai_mai_n44_), .Y(mai_mai_n363_));
  NOi31      m0335(.An(mai_mai_n351_), .B(mai_mai_n361_), .C(mai_mai_n219_), .Y(mai_mai_n364_));
  NOi32      m0336(.An(c), .Bn(a), .C(b), .Y(mai_mai_n365_));
  NA2        m0337(.A(mai_mai_n365_), .B(mai_mai_n89_), .Y(mai_mai_n366_));
  AN2        m0338(.A(e), .B(d), .Y(mai_mai_n367_));
  NO2        m0339(.A(mai_mai_n118_), .B(mai_mai_n366_), .Y(mai_mai_n368_));
  NA3        m0340(.A(e), .B(d), .C(c), .Y(mai_mai_n369_));
  NAi21      m0341(.An(mai_mai_n369_), .B(a), .Y(mai_mai_n370_));
  INV        m0342(.A(mai_mai_n169_), .Y(mai_mai_n371_));
  NOi21      m0343(.An(mai_mai_n370_), .B(mai_mai_n371_), .Y(mai_mai_n372_));
  NO2        m0344(.A(mai_mai_n1092_), .B(mai_mai_n372_), .Y(mai_mai_n373_));
  NO4        m0345(.A(mai_mai_n154_), .B(mai_mai_n80_), .C(mai_mai_n49_), .D(b), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n308_), .B(mai_mai_n123_), .Y(mai_mai_n375_));
  NA2        m0347(.A(l), .B(k), .Y(mai_mai_n376_));
  NA3        m0348(.A(mai_mai_n376_), .B(j), .C(mai_mai_n182_), .Y(mai_mai_n377_));
  AOI210     m0349(.A0(mai_mai_n195_), .A1(mai_mai_n268_), .B0(mai_mai_n69_), .Y(mai_mai_n378_));
  NOi21      m0350(.An(mai_mai_n377_), .B(mai_mai_n378_), .Y(mai_mai_n379_));
  OR3        m0351(.A(mai_mai_n379_), .B(mai_mai_n114_), .C(mai_mai_n104_), .Y(mai_mai_n380_));
  NA2        m0352(.A(mai_mai_n230_), .B(mai_mai_n97_), .Y(mai_mai_n381_));
  NA2        m0353(.A(mai_mai_n321_), .B(mai_mai_n89_), .Y(mai_mai_n382_));
  NO3        m0354(.A(mai_mai_n338_), .B(mai_mai_n74_), .C(mai_mai_n100_), .Y(mai_mai_n383_));
  NO2        m0355(.A(mai_mai_n383_), .B(mai_mai_n381_), .Y(mai_mai_n384_));
  NA3        m0356(.A(mai_mai_n384_), .B(mai_mai_n380_), .C(mai_mai_n375_), .Y(mai_mai_n385_));
  NO4        m0357(.A(mai_mai_n385_), .B(mai_mai_n374_), .C(mai_mai_n373_), .D(mai_mai_n368_), .Y(mai_mai_n386_));
  NOi21      m0358(.An(d), .B(e), .Y(mai_mai_n387_));
  NO2        m0359(.A(mai_mai_n154_), .B(mai_mai_n49_), .Y(mai_mai_n388_));
  NAi31      m0360(.An(j), .B(l), .C(i), .Y(mai_mai_n389_));
  OAI210     m0361(.A0(mai_mai_n389_), .A1(mai_mai_n101_), .B0(mai_mai_n80_), .Y(mai_mai_n390_));
  NA3        m0362(.A(mai_mai_n390_), .B(mai_mai_n388_), .C(mai_mai_n387_), .Y(mai_mai_n391_));
  NO3        m0363(.A(mai_mai_n322_), .B(mai_mai_n274_), .C(mai_mai_n166_), .Y(mai_mai_n392_));
  NO2        m0364(.A(mai_mai_n322_), .B(mai_mai_n297_), .Y(mai_mai_n393_));
  NO3        m0365(.A(mai_mai_n393_), .B(mai_mai_n392_), .C(mai_mai_n248_), .Y(mai_mai_n394_));
  NA3        m0366(.A(mai_mai_n394_), .B(mai_mai_n391_), .C(mai_mai_n204_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n96_), .B(mai_mai_n95_), .Y(mai_mai_n396_));
  NO2        m0368(.A(mai_mai_n396_), .B(mai_mai_n100_), .Y(mai_mai_n397_));
  XO2        m0369(.A(i), .B(h), .Y(mai_mai_n398_));
  NA3        m0370(.A(mai_mai_n398_), .B(mai_mai_n130_), .C(n), .Y(mai_mai_n399_));
  NA3        m0371(.A(mai_mai_n399_), .B(mai_mai_n363_), .C(mai_mai_n310_), .Y(mai_mai_n400_));
  NAi31      m0372(.An(c), .B(f), .C(d), .Y(mai_mai_n401_));
  AOI210     m0373(.A0(mai_mai_n231_), .A1(mai_mai_n160_), .B0(mai_mai_n401_), .Y(mai_mai_n402_));
  NOi21      m0374(.An(mai_mai_n67_), .B(mai_mai_n402_), .Y(mai_mai_n403_));
  NA3        m0375(.A(mai_mai_n306_), .B(mai_mai_n78_), .C(g), .Y(mai_mai_n404_));
  NA2        m0376(.A(mai_mai_n189_), .B(mai_mai_n84_), .Y(mai_mai_n405_));
  AOI210     m0377(.A0(mai_mai_n405_), .A1(mai_mai_n149_), .B0(mai_mai_n401_), .Y(mai_mai_n406_));
  NOi21      m0378(.An(mai_mai_n404_), .B(mai_mai_n406_), .Y(mai_mai_n407_));
  NA3        m0379(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(f), .Y(mai_mai_n408_));
  NO2        m0380(.A(mai_mai_n408_), .B(mai_mai_n346_), .Y(mai_mai_n409_));
  NO2        m0381(.A(mai_mai_n409_), .B(mai_mai_n238_), .Y(mai_mai_n410_));
  NA3        m0382(.A(mai_mai_n410_), .B(mai_mai_n407_), .C(mai_mai_n403_), .Y(mai_mai_n411_));
  NO2        m0383(.A(mai_mai_n411_), .B(mai_mai_n395_), .Y(mai_mai_n412_));
  NA4        m0384(.A(mai_mai_n412_), .B(mai_mai_n386_), .C(mai_mai_n364_), .D(mai_mai_n342_), .Y(mai11));
  INV        m0385(.A(mai_mai_n58_), .Y(mai_mai_n414_));
  NA2        m0386(.A(j), .B(g), .Y(mai_mai_n415_));
  NAi31      m0387(.An(i), .B(m), .C(l), .Y(mai_mai_n416_));
  NA3        m0388(.A(m), .B(k), .C(j), .Y(mai_mai_n417_));
  OAI220     m0389(.A0(mai_mai_n417_), .A1(mai_mai_n100_), .B0(mai_mai_n416_), .B1(mai_mai_n415_), .Y(mai_mai_n418_));
  NA2        m0390(.A(mai_mai_n418_), .B(mai_mai_n414_), .Y(mai_mai_n419_));
  NOi32      m0391(.An(e), .Bn(b), .C(f), .Y(mai_mai_n420_));
  NA2        m0392(.A(mai_mai_n42_), .B(j), .Y(mai_mai_n421_));
  NO2        m0393(.A(mai_mai_n421_), .B(mai_mai_n244_), .Y(mai_mai_n422_));
  NAi31      m0394(.An(d), .B(e), .C(a), .Y(mai_mai_n423_));
  NO2        m0395(.A(mai_mai_n423_), .B(n), .Y(mai_mai_n424_));
  INV        m0396(.A(mai_mai_n422_), .Y(mai_mai_n425_));
  NAi41      m0397(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n426_));
  AN2        m0398(.A(mai_mai_n426_), .B(mai_mai_n296_), .Y(mai_mai_n427_));
  NAi31      m0399(.An(n), .B(m), .C(k), .Y(mai_mai_n428_));
  NO2        m0400(.A(n), .B(d), .Y(mai_mai_n429_));
  NO2        m0401(.A(n), .B(mai_mai_n120_), .Y(mai_mai_n430_));
  NA2        m0402(.A(mai_mai_n418_), .B(f), .Y(mai_mai_n431_));
  NO2        m0403(.A(mai_mai_n431_), .B(n), .Y(mai_mai_n432_));
  INV        m0404(.A(mai_mai_n432_), .Y(mai_mai_n433_));
  NA2        m0405(.A(mai_mai_n110_), .B(mai_mai_n33_), .Y(mai_mai_n434_));
  NOi41      m0406(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n435_));
  NAi32      m0407(.An(e), .Bn(b), .C(c), .Y(mai_mai_n436_));
  AN2        m0408(.A(mai_mai_n269_), .B(mai_mai_n254_), .Y(mai_mai_n437_));
  OAI220     m0409(.A0(mai_mai_n323_), .A1(i), .B0(mai_mai_n416_), .B1(mai_mai_n415_), .Y(mai_mai_n438_));
  NAi31      m0410(.An(d), .B(c), .C(a), .Y(mai_mai_n439_));
  NO2        m0411(.A(mai_mai_n439_), .B(n), .Y(mai_mai_n440_));
  NA3        m0412(.A(mai_mai_n440_), .B(mai_mai_n438_), .C(e), .Y(mai_mai_n441_));
  NO3        m0413(.A(i), .B(mai_mai_n43_), .C(mai_mai_n175_), .Y(mai_mai_n442_));
  INV        m0414(.A(mai_mai_n441_), .Y(mai_mai_n443_));
  NA2        m0415(.A(mai_mai_n438_), .B(f), .Y(mai_mai_n444_));
  NO3        m0416(.A(mai_mai_n145_), .B(mai_mai_n142_), .C(g), .Y(mai_mai_n445_));
  NA2        m0417(.A(mai_mai_n445_), .B(mai_mai_n51_), .Y(mai_mai_n446_));
  INV        m0418(.A(mai_mai_n446_), .Y(mai_mai_n447_));
  NA3        m0419(.A(f), .B(d), .C(b), .Y(mai_mai_n448_));
  NO3        m0420(.A(mai_mai_n448_), .B(mai_mai_n145_), .C(mai_mai_n142_), .Y(mai_mai_n449_));
  NO2        m0421(.A(mai_mai_n449_), .B(mai_mai_n447_), .Y(mai_mai_n450_));
  AN4        m0422(.A(mai_mai_n450_), .B(mai_mai_n433_), .C(mai_mai_n425_), .D(mai_mai_n419_), .Y(mai_mai_n451_));
  INV        m0423(.A(k), .Y(mai_mai_n452_));
  NA4        m0424(.A(mai_mai_n321_), .B(mai_mai_n332_), .C(mai_mai_n150_), .D(mai_mai_n89_), .Y(mai_mai_n453_));
  NAi32      m0425(.An(h), .Bn(f), .C(g), .Y(mai_mai_n454_));
  NAi41      m0426(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n455_));
  OAI210     m0427(.A0(mai_mai_n423_), .A1(n), .B0(mai_mai_n455_), .Y(mai_mai_n456_));
  NA2        m0428(.A(mai_mai_n456_), .B(m), .Y(mai_mai_n457_));
  NAi31      m0429(.An(h), .B(g), .C(f), .Y(mai_mai_n458_));
  NO3        m0430(.A(mai_mai_n454_), .B(mai_mai_n58_), .C(mai_mai_n59_), .Y(mai_mai_n459_));
  NO4        m0431(.A(mai_mai_n458_), .B(n), .C(mai_mai_n120_), .D(mai_mai_n59_), .Y(mai_mai_n460_));
  OR2        m0432(.A(mai_mai_n460_), .B(mai_mai_n459_), .Y(mai_mai_n461_));
  NAi31      m0433(.An(mai_mai_n461_), .B(mai_mai_n457_), .C(mai_mai_n453_), .Y(mai_mai_n462_));
  NAi31      m0434(.An(f), .B(h), .C(g), .Y(mai_mai_n463_));
  NOi31      m0435(.An(b), .B(mai_mai_n281_), .C(mai_mai_n55_), .Y(mai_mai_n464_));
  NOi32      m0436(.An(d), .Bn(a), .C(e), .Y(mai_mai_n465_));
  INV        m0437(.A(mai_mai_n89_), .Y(mai_mai_n466_));
  NO2        m0438(.A(n), .B(c), .Y(mai_mai_n467_));
  NOi32      m0439(.An(e), .Bn(a), .C(d), .Y(mai_mai_n468_));
  AOI210     m0440(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n468_), .Y(mai_mai_n469_));
  NO2        m0441(.A(mai_mai_n174_), .B(mai_mai_n434_), .Y(mai_mai_n470_));
  AOI210     m0442(.A0(mai_mai_n470_), .A1(mai_mai_n89_), .B0(mai_mai_n464_), .Y(mai_mai_n471_));
  OAI210     m0443(.A0(mai_mai_n208_), .A1(mai_mai_n71_), .B0(mai_mai_n471_), .Y(mai_mai_n472_));
  NO2        m0444(.A(mai_mai_n462_), .B(mai_mai_n472_), .Y(mai_mai_n473_));
  NO2        m0445(.A(mai_mai_n252_), .B(mai_mai_n53_), .Y(mai_mai_n474_));
  NA3        m0446(.A(mai_mai_n401_), .B(mai_mai_n140_), .C(mai_mai_n139_), .Y(mai_mai_n475_));
  INV        m0447(.A(mai_mai_n192_), .Y(mai_mai_n476_));
  NA2        m0448(.A(mai_mai_n475_), .B(mai_mai_n474_), .Y(mai_mai_n477_));
  NO2        m0449(.A(mai_mai_n477_), .B(mai_mai_n71_), .Y(mai_mai_n478_));
  NOi32      m0450(.An(e), .Bn(c), .C(f), .Y(mai_mai_n479_));
  NOi21      m0451(.An(f), .B(g), .Y(mai_mai_n480_));
  NO2        m0452(.A(mai_mai_n480_), .B(mai_mai_n172_), .Y(mai_mai_n481_));
  AOI220     m0453(.A0(mai_mai_n481_), .A1(mai_mai_n318_), .B0(mai_mai_n479_), .B1(mai_mai_n144_), .Y(mai_mai_n482_));
  NA2        m0454(.A(mai_mai_n482_), .B(mai_mai_n147_), .Y(mai_mai_n483_));
  AOI210     m0455(.A0(mai_mai_n427_), .A1(mai_mai_n322_), .B0(mai_mai_n243_), .Y(mai_mai_n484_));
  NA2        m0456(.A(mai_mai_n484_), .B(mai_mai_n218_), .Y(mai_mai_n485_));
  NAi21      m0457(.An(k), .B(h), .Y(mai_mai_n486_));
  NO2        m0458(.A(mai_mai_n486_), .B(f), .Y(mai_mai_n487_));
  OR2        m0459(.A(mai_mai_n486_), .B(mai_mai_n457_), .Y(mai_mai_n488_));
  NOi31      m0460(.An(m), .B(n), .C(k), .Y(mai_mai_n489_));
  INV        m0461(.A(mai_mai_n43_), .Y(mai_mai_n490_));
  NA2        m0462(.A(mai_mai_n488_), .B(mai_mai_n485_), .Y(mai_mai_n491_));
  NA2        m0463(.A(mai_mai_n84_), .B(mai_mai_n35_), .Y(mai_mai_n492_));
  NO2        m0464(.A(mai_mai_n420_), .B(mai_mai_n288_), .Y(mai_mai_n493_));
  NO2        m0465(.A(mai_mai_n493_), .B(n), .Y(mai_mai_n494_));
  NAi21      m0466(.An(mai_mai_n492_), .B(mai_mai_n494_), .Y(mai_mai_n495_));
  NO2        m0467(.A(mai_mai_n421_), .B(mai_mai_n145_), .Y(mai_mai_n496_));
  NA2        m0468(.A(mai_mai_n398_), .B(mai_mai_n130_), .Y(mai_mai_n497_));
  NO3        m0469(.A(mai_mai_n319_), .B(mai_mai_n497_), .C(mai_mai_n71_), .Y(mai_mai_n498_));
  AOI210     m0470(.A0(c), .A1(mai_mai_n496_), .B0(mai_mai_n498_), .Y(mai_mai_n499_));
  NAi31      m0471(.An(m), .B(n), .C(k), .Y(mai_mai_n500_));
  OR2        m0472(.A(mai_mai_n104_), .B(mai_mai_n53_), .Y(mai_mai_n501_));
  NO2        m0473(.A(mai_mai_n501_), .B(mai_mai_n500_), .Y(mai_mai_n502_));
  NA2        m0474(.A(mai_mai_n502_), .B(j), .Y(mai_mai_n503_));
  NA3        m0475(.A(mai_mai_n503_), .B(mai_mai_n499_), .C(mai_mai_n495_), .Y(mai_mai_n504_));
  NO4        m0476(.A(mai_mai_n504_), .B(mai_mai_n491_), .C(mai_mai_n483_), .D(mai_mai_n478_), .Y(mai_mai_n505_));
  NAi31      m0477(.An(g), .B(h), .C(f), .Y(mai_mai_n506_));
  OR3        m0478(.A(mai_mai_n506_), .B(mai_mai_n228_), .C(n), .Y(mai_mai_n507_));
  BUFFER     m0479(.A(mai_mai_n455_), .Y(mai_mai_n508_));
  NA3        m0480(.A(e), .B(mai_mai_n94_), .C(mai_mai_n69_), .Y(mai_mai_n509_));
  OR2        m0481(.A(mai_mai_n58_), .B(mai_mai_n59_), .Y(mai_mai_n510_));
  OR2        m0482(.A(mai_mai_n486_), .B(mai_mai_n510_), .Y(mai_mai_n511_));
  AN2        m0483(.A(h), .B(f), .Y(mai_mai_n512_));
  NA2        m0484(.A(mai_mai_n512_), .B(mai_mai_n36_), .Y(mai_mai_n513_));
  NO2        m0485(.A(mai_mai_n513_), .B(mai_mai_n366_), .Y(mai_mai_n514_));
  AOI210     m0486(.A0(d), .A1(mai_mai_n339_), .B0(mai_mai_n43_), .Y(mai_mai_n515_));
  NO2        m0487(.A(mai_mai_n458_), .B(k), .Y(mai_mai_n516_));
  AOI210     m0488(.A0(mai_mai_n516_), .A1(mai_mai_n515_), .B0(mai_mai_n514_), .Y(mai_mai_n517_));
  NA2        m0489(.A(mai_mai_n517_), .B(mai_mai_n511_), .Y(mai_mai_n518_));
  NO2        m0490(.A(mai_mai_n210_), .B(f), .Y(mai_mai_n519_));
  INV        m0491(.A(mai_mai_n53_), .Y(mai_mai_n520_));
  NO3        m0492(.A(mai_mai_n520_), .B(mai_mai_n519_), .C(mai_mai_n33_), .Y(mai_mai_n521_));
  NA2        m0493(.A(mai_mai_n260_), .B(mai_mai_n110_), .Y(mai_mai_n522_));
  OA220      m0494(.A0(mai_mai_n1091_), .A1(mai_mai_n434_), .B0(mai_mai_n286_), .B1(mai_mai_n87_), .Y(mai_mai_n523_));
  OAI210     m0495(.A0(mai_mai_n522_), .A1(mai_mai_n521_), .B0(mai_mai_n523_), .Y(mai_mai_n524_));
  NO3        m0496(.A(mai_mai_n326_), .B(mai_mai_n157_), .C(mai_mai_n156_), .Y(mai_mai_n525_));
  NA2        m0497(.A(mai_mai_n525_), .B(mai_mai_n192_), .Y(mai_mai_n526_));
  NA3        m0498(.A(mai_mai_n526_), .B(mai_mai_n212_), .C(j), .Y(mai_mai_n527_));
  NA2        m0499(.A(mai_mai_n365_), .B(mai_mai_n69_), .Y(mai_mai_n528_));
  NA3        m0500(.A(mai_mai_n527_), .B(mai_mai_n404_), .C(mai_mai_n324_), .Y(mai_mai_n529_));
  NO3        m0501(.A(mai_mai_n529_), .B(mai_mai_n524_), .C(mai_mai_n518_), .Y(mai_mai_n530_));
  NA4        m0502(.A(mai_mai_n530_), .B(mai_mai_n505_), .C(mai_mai_n473_), .D(mai_mai_n451_), .Y(mai08));
  NO2        m0503(.A(k), .B(h), .Y(mai_mai_n532_));
  AO210      m0504(.A0(mai_mai_n210_), .A1(mai_mai_n356_), .B0(mai_mai_n532_), .Y(mai_mai_n533_));
  NO2        m0505(.A(mai_mai_n533_), .B(mai_mai_n241_), .Y(mai_mai_n534_));
  NA2        m0506(.A(mai_mai_n479_), .B(mai_mai_n69_), .Y(mai_mai_n535_));
  AOI210     m0507(.A0(mai_mai_n479_), .A1(mai_mai_n534_), .B0(mai_mai_n383_), .Y(mai_mai_n536_));
  NA2        m0508(.A(mai_mai_n69_), .B(mai_mai_n86_), .Y(mai_mai_n537_));
  NO2        m0509(.A(mai_mai_n537_), .B(mai_mai_n50_), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n303_), .B(mai_mai_n88_), .Y(mai_mai_n539_));
  NA2        m0511(.A(mai_mai_n448_), .B(mai_mai_n194_), .Y(mai_mai_n540_));
  AOI220     m0512(.A0(mai_mai_n540_), .A1(mai_mai_n276_), .B0(mai_mai_n539_), .B1(mai_mai_n538_), .Y(mai_mai_n541_));
  NA4        m0513(.A(mai_mai_n177_), .B(mai_mai_n110_), .C(mai_mai_n41_), .D(h), .Y(mai_mai_n542_));
  AN2        m0514(.A(l), .B(k), .Y(mai_mai_n543_));
  NA4        m0515(.A(mai_mai_n543_), .B(mai_mai_n84_), .C(mai_mai_n59_), .D(mai_mai_n175_), .Y(mai_mai_n544_));
  NA3        m0516(.A(mai_mai_n541_), .B(mai_mai_n536_), .C(mai_mai_n278_), .Y(mai_mai_n545_));
  NO4        m0517(.A(mai_mai_n142_), .B(mai_mai_n317_), .C(mai_mai_n88_), .D(g), .Y(mai_mai_n546_));
  AOI210     m0518(.A0(mai_mai_n546_), .A1(mai_mai_n540_), .B0(mai_mai_n409_), .Y(mai_mai_n547_));
  NA2        m0519(.A(mai_mai_n481_), .B(mai_mai_n275_), .Y(mai_mai_n548_));
  NA2        m0520(.A(mai_mai_n548_), .B(mai_mai_n547_), .Y(mai_mai_n549_));
  NO2        m0521(.A(mai_mai_n376_), .B(mai_mai_n101_), .Y(mai_mai_n550_));
  NA2        m0522(.A(mai_mai_n550_), .B(mai_mai_n1096_), .Y(mai_mai_n551_));
  NO3        m0523(.A(mai_mai_n252_), .B(mai_mai_n100_), .C(mai_mai_n40_), .Y(mai_mai_n552_));
  NAi21      m0524(.An(mai_mai_n552_), .B(mai_mai_n544_), .Y(mai_mai_n553_));
  NA2        m0525(.A(mai_mai_n533_), .B(mai_mai_n105_), .Y(mai_mai_n554_));
  AOI220     m0526(.A0(mai_mai_n554_), .A1(mai_mai_n325_), .B0(mai_mai_n553_), .B1(mai_mai_n61_), .Y(mai_mai_n555_));
  OAI210     m0527(.A0(mai_mai_n551_), .A1(mai_mai_n71_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  NA3        m0528(.A(mai_mai_n526_), .B(mai_mai_n266_), .C(mai_mai_n309_), .Y(mai_mai_n557_));
  NA2        m0529(.A(mai_mai_n543_), .B(mai_mai_n182_), .Y(mai_mai_n558_));
  NO2        m0530(.A(mai_mai_n558_), .B(mai_mai_n259_), .Y(mai_mai_n559_));
  NA2        m0531(.A(mai_mai_n559_), .B(mai_mai_n519_), .Y(mai_mai_n560_));
  NA3        m0532(.A(m), .B(l), .C(k), .Y(mai_mai_n561_));
  AOI210     m0533(.A0(mai_mai_n509_), .A1(mai_mai_n507_), .B0(mai_mai_n561_), .Y(mai_mai_n562_));
  INV        m0534(.A(mai_mai_n562_), .Y(mai_mai_n563_));
  NA3        m0535(.A(mai_mai_n563_), .B(mai_mai_n560_), .C(mai_mai_n557_), .Y(mai_mai_n564_));
  NO4        m0536(.A(mai_mai_n564_), .B(mai_mai_n556_), .C(mai_mai_n549_), .D(mai_mai_n545_), .Y(mai_mai_n565_));
  NA2        m0537(.A(g), .B(mai_mai_n89_), .Y(mai_mai_n566_));
  NA2        m0538(.A(mai_mai_n566_), .B(mai_mai_n208_), .Y(mai_mai_n567_));
  NA2        m0539(.A(mai_mai_n543_), .B(mai_mai_n59_), .Y(mai_mai_n568_));
  NO3        m0540(.A(mai_mai_n525_), .B(mai_mai_n142_), .C(i), .Y(mai_mai_n569_));
  NOi21      m0541(.An(h), .B(j), .Y(mai_mai_n570_));
  NA2        m0542(.A(mai_mai_n570_), .B(f), .Y(mai_mai_n571_));
  NO2        m0543(.A(mai_mai_n571_), .B(mai_mai_n205_), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n572_), .B(mai_mai_n569_), .Y(mai_mai_n573_));
  NO2        m0545(.A(mai_mai_n573_), .B(mai_mai_n568_), .Y(mai_mai_n574_));
  AOI210     m0546(.A0(mai_mai_n567_), .A1(l), .B0(mai_mai_n574_), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n65_), .B(l), .Y(mai_mai_n576_));
  OR2        m0548(.A(mai_mai_n576_), .B(mai_mai_n457_), .Y(mai_mai_n577_));
  NO2        m0549(.A(mai_mai_n43_), .B(mai_mai_n86_), .Y(mai_mai_n578_));
  NO3        m0550(.A(n), .B(mai_mai_n120_), .C(mai_mai_n59_), .Y(mai_mai_n579_));
  NA2        m0551(.A(k), .B(j), .Y(mai_mai_n580_));
  NO2        m0552(.A(mai_mai_n580_), .B(mai_mai_n39_), .Y(mai_mai_n581_));
  AOI210     m0553(.A0(mai_mai_n420_), .A1(n), .B0(mai_mai_n435_), .Y(mai_mai_n582_));
  NA2        m0554(.A(mai_mai_n582_), .B(mai_mai_n437_), .Y(mai_mai_n583_));
  AN3        m0555(.A(mai_mai_n583_), .B(mai_mai_n581_), .C(mai_mai_n79_), .Y(mai_mai_n584_));
  NO3        m0556(.A(mai_mai_n142_), .B(mai_mai_n317_), .C(mai_mai_n88_), .Y(mai_mai_n585_));
  NA2        m0557(.A(mai_mai_n585_), .B(mai_mai_n206_), .Y(mai_mai_n586_));
  NAi31      m0558(.An(mai_mai_n469_), .B(mai_mai_n75_), .C(mai_mai_n69_), .Y(mai_mai_n587_));
  NA2        m0559(.A(mai_mai_n587_), .B(mai_mai_n586_), .Y(mai_mai_n588_));
  NO2        m0560(.A(mai_mai_n561_), .B(mai_mai_n73_), .Y(mai_mai_n589_));
  NA2        m0561(.A(mai_mai_n589_), .B(mai_mai_n456_), .Y(mai_mai_n590_));
  INV        m0562(.A(mai_mai_n590_), .Y(mai_mai_n591_));
  OR3        m0563(.A(mai_mai_n591_), .B(mai_mai_n588_), .C(mai_mai_n584_), .Y(mai_mai_n592_));
  NA2        m0564(.A(mai_mai_n582_), .B(mai_mai_n437_), .Y(mai_mai_n593_));
  NA4        m0565(.A(mai_mai_n593_), .B(mai_mai_n177_), .C(mai_mai_n356_), .D(mai_mai_n33_), .Y(mai_mai_n594_));
  NA3        m0566(.A(g), .B(mai_mai_n236_), .C(h), .Y(mai_mai_n595_));
  NOi21      m0567(.An(mai_mai_n515_), .B(mai_mai_n595_), .Y(mai_mai_n596_));
  INV        m0568(.A(mai_mai_n74_), .Y(mai_mai_n597_));
  NO2        m0569(.A(mai_mai_n576_), .B(mai_mai_n510_), .Y(mai_mai_n598_));
  AOI210     m0570(.A0(mai_mai_n597_), .A1(mai_mai_n494_), .B0(mai_mai_n598_), .Y(mai_mai_n599_));
  NAi31      m0571(.An(mai_mai_n596_), .B(mai_mai_n599_), .C(mai_mai_n594_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n589_), .B(mai_mai_n200_), .Y(mai_mai_n601_));
  OAI210     m0573(.A0(mai_mai_n561_), .A1(mai_mai_n506_), .B0(mai_mai_n408_), .Y(mai_mai_n602_));
  NA3        m0574(.A(mai_mai_n209_), .B(mai_mai_n52_), .C(b), .Y(mai_mai_n603_));
  AOI220     m0575(.A0(mai_mai_n467_), .A1(mai_mai_n29_), .B0(mai_mai_n365_), .B1(mai_mai_n69_), .Y(mai_mai_n604_));
  NA2        m0576(.A(mai_mai_n604_), .B(mai_mai_n603_), .Y(mai_mai_n605_));
  NO2        m0577(.A(mai_mai_n595_), .B(mai_mai_n382_), .Y(mai_mai_n606_));
  AOI210     m0578(.A0(mai_mai_n605_), .A1(mai_mai_n602_), .B0(mai_mai_n606_), .Y(mai_mai_n607_));
  NA2        m0579(.A(mai_mai_n607_), .B(mai_mai_n601_), .Y(mai_mai_n608_));
  NOi41      m0580(.An(mai_mai_n577_), .B(mai_mai_n608_), .C(mai_mai_n600_), .D(mai_mai_n592_), .Y(mai_mai_n609_));
  OR2        m0581(.A(mai_mai_n542_), .B(mai_mai_n194_), .Y(mai_mai_n610_));
  NO3        m0582(.A(mai_mai_n271_), .B(mai_mai_n243_), .C(mai_mai_n88_), .Y(mai_mai_n611_));
  NA2        m0583(.A(mai_mai_n611_), .B(mai_mai_n583_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n610_), .Y(mai_mai_n613_));
  OR2        m0585(.A(mai_mai_n506_), .B(mai_mai_n74_), .Y(mai_mai_n614_));
  NOi31      m0586(.An(b), .B(d), .C(a), .Y(mai_mai_n615_));
  NO2        m0587(.A(mai_mai_n615_), .B(mai_mai_n465_), .Y(mai_mai_n616_));
  NO2        m0588(.A(mai_mai_n616_), .B(n), .Y(mai_mai_n617_));
  NOi21      m0589(.An(mai_mai_n604_), .B(mai_mai_n617_), .Y(mai_mai_n618_));
  OAI220     m0590(.A0(mai_mai_n618_), .A1(mai_mai_n614_), .B0(mai_mai_n595_), .B1(mai_mai_n466_), .Y(mai_mai_n619_));
  NO2        m0591(.A(mai_mai_n525_), .B(n), .Y(mai_mai_n620_));
  NA2        m0592(.A(mai_mai_n620_), .B(mai_mai_n534_), .Y(mai_mai_n621_));
  NO2        m0593(.A(mai_mai_n255_), .B(mai_mai_n199_), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n77_), .B(mai_mai_n622_), .Y(mai_mai_n623_));
  NA2        m0595(.A(mai_mai_n94_), .B(mai_mai_n69_), .Y(mai_mai_n624_));
  AOI210     m0596(.A0(mai_mai_n337_), .A1(mai_mai_n331_), .B0(mai_mai_n624_), .Y(mai_mai_n625_));
  NAi21      m0597(.An(mai_mai_n625_), .B(mai_mai_n623_), .Y(mai_mai_n626_));
  NA2        m0598(.A(mai_mai_n559_), .B(mai_mai_n33_), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n224_), .B(i), .Y(mai_mai_n628_));
  NA2        m0600(.A(mai_mai_n546_), .B(mai_mai_n277_), .Y(mai_mai_n629_));
  NAi41      m0601(.An(mai_mai_n626_), .B(mai_mai_n629_), .C(mai_mai_n627_), .D(mai_mai_n621_), .Y(mai_mai_n630_));
  NO3        m0602(.A(mai_mai_n630_), .B(mai_mai_n619_), .C(mai_mai_n613_), .Y(mai_mai_n631_));
  NA4        m0603(.A(mai_mai_n631_), .B(mai_mai_n609_), .C(mai_mai_n575_), .D(mai_mai_n565_), .Y(mai09));
  NA4        m0604(.A(k), .B(l), .C(i), .D(j), .Y(mai_mai_n633_));
  NA2        m0605(.A(mai_mai_n353_), .B(e), .Y(mai_mai_n634_));
  NO2        m0606(.A(mai_mai_n169_), .B(mai_mai_n174_), .Y(mai_mai_n635_));
  NA3        m0607(.A(m), .B(l), .C(i), .Y(mai_mai_n636_));
  OAI220     m0608(.A0(mai_mai_n458_), .A1(mai_mai_n636_), .B0(mai_mai_n281_), .B1(mai_mai_n416_), .Y(mai_mai_n637_));
  NA4        m0609(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(g), .D(f), .Y(mai_mai_n638_));
  NAi31      m0610(.An(mai_mai_n637_), .B(mai_mai_n638_), .C(mai_mai_n348_), .Y(mai_mai_n639_));
  OR2        m0611(.A(mai_mai_n639_), .B(mai_mai_n635_), .Y(mai_mai_n640_));
  NA3        m0612(.A(mai_mai_n614_), .B(mai_mai_n444_), .C(mai_mai_n408_), .Y(mai_mai_n641_));
  OA210      m0613(.A0(mai_mai_n641_), .A1(mai_mai_n640_), .B0(mai_mai_n617_), .Y(mai_mai_n642_));
  INV        m0614(.A(mai_mai_n269_), .Y(mai_mai_n643_));
  NOi31      m0615(.An(k), .B(m), .C(l), .Y(mai_mai_n644_));
  NO2        m0616(.A(m), .B(mai_mai_n463_), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n272_), .B(mai_mai_n273_), .Y(mai_mai_n646_));
  OAI210     m0618(.A0(mai_mai_n169_), .A1(mai_mai_n174_), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  AOI220     m0619(.A0(mai_mai_n647_), .A1(mai_mai_n209_), .B0(mai_mai_n645_), .B1(mai_mai_n643_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n90_), .B(mai_mai_n155_), .C(mai_mai_n31_), .Y(mai_mai_n649_));
  NA4        m0621(.A(mai_mai_n649_), .B(mai_mai_n648_), .C(mai_mai_n482_), .D(mai_mai_n67_), .Y(mai_mai_n650_));
  NO2        m0622(.A(mai_mai_n454_), .B(mai_mai_n389_), .Y(mai_mai_n651_));
  NA2        m0623(.A(mai_mai_n651_), .B(mai_mai_n155_), .Y(mai_mai_n652_));
  NA2        m0624(.A(f), .B(m), .Y(mai_mai_n653_));
  NO2        m0625(.A(mai_mai_n653_), .B(mai_mai_n46_), .Y(mai_mai_n654_));
  NA4        m0626(.A(g), .B(mai_mai_n467_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n655_));
  INV        m0627(.A(mai_mai_n655_), .Y(mai_mai_n656_));
  AOI210     m0628(.A0(mai_mai_n654_), .A1(mai_mai_n430_), .B0(mai_mai_n656_), .Y(mai_mai_n657_));
  NA3        m0629(.A(k), .B(i), .C(j), .Y(mai_mai_n658_));
  NA3        m0630(.A(a), .B(f), .C(mai_mai_n69_), .Y(mai_mai_n659_));
  NO2        m0631(.A(mai_mai_n659_), .B(mai_mai_n59_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n658_), .B(mai_mai_n660_), .Y(mai_mai_n661_));
  NAi31      m0633(.An(mai_mai_n381_), .B(mai_mai_n661_), .C(mai_mai_n652_), .Y(mai_mai_n662_));
  NO4        m0634(.A(mai_mai_n480_), .B(mai_mai_n101_), .C(mai_mai_n259_), .D(mai_mai_n122_), .Y(mai_mai_n663_));
  NO2        m0635(.A(mai_mai_n500_), .B(mai_mai_n259_), .Y(mai_mai_n664_));
  AN2        m0636(.A(mai_mai_n664_), .B(mai_mai_n519_), .Y(mai_mai_n665_));
  NO3        m0637(.A(mai_mai_n665_), .B(mai_mai_n663_), .C(mai_mai_n196_), .Y(mai_mai_n666_));
  NO2        m0638(.A(mai_mai_n659_), .B(mai_mai_n341_), .Y(mai_mai_n667_));
  NOi31      m0639(.An(mai_mai_n185_), .B(mai_mai_n667_), .C(mai_mai_n248_), .Y(mai_mai_n668_));
  NA2        m0640(.A(c), .B(mai_mai_n92_), .Y(mai_mai_n669_));
  NO2        m0641(.A(mai_mai_n669_), .B(mai_mai_n329_), .Y(mai_mai_n670_));
  NA3        m0642(.A(mai_mai_n670_), .B(mai_mai_n400_), .C(f), .Y(mai_mai_n671_));
  OR2        m0643(.A(mai_mai_n506_), .B(mai_mai_n428_), .Y(mai_mai_n672_));
  NA4        m0644(.A(mai_mai_n672_), .B(mai_mai_n671_), .C(mai_mai_n668_), .D(mai_mai_n666_), .Y(mai_mai_n673_));
  NO4        m0645(.A(mai_mai_n673_), .B(mai_mai_n662_), .C(mai_mai_n650_), .D(mai_mai_n642_), .Y(mai_mai_n674_));
  OR2        m0646(.A(mai_mai_n659_), .B(mai_mai_n59_), .Y(mai_mai_n675_));
  NO2        m0647(.A(h), .B(mai_mai_n675_), .Y(mai_mai_n676_));
  NO2        m0648(.A(mai_mai_n264_), .B(mai_mai_n638_), .Y(mai_mai_n677_));
  NO2        m0649(.A(mai_mai_n105_), .B(mai_mai_n101_), .Y(mai_mai_n678_));
  NO2        m0650(.A(mai_mai_n192_), .B(mai_mai_n186_), .Y(mai_mai_n679_));
  AOI220     m0651(.A0(mai_mai_n679_), .A1(mai_mai_n189_), .B0(mai_mai_n247_), .B1(mai_mai_n678_), .Y(mai_mai_n680_));
  INV        m0652(.A(mai_mai_n680_), .Y(mai_mai_n681_));
  NA2        m0653(.A(e), .B(d), .Y(mai_mai_n682_));
  OAI220     m0654(.A0(mai_mai_n682_), .A1(c), .B0(mai_mai_n255_), .B1(d), .Y(mai_mai_n683_));
  NA3        m0655(.A(mai_mai_n683_), .B(mai_mai_n359_), .C(mai_mai_n398_), .Y(mai_mai_n684_));
  AOI210     m0656(.A0(mai_mai_n405_), .A1(mai_mai_n149_), .B0(mai_mai_n192_), .Y(mai_mai_n685_));
  AOI210     m0657(.A0(mai_mai_n481_), .A1(mai_mai_n275_), .B0(mai_mai_n685_), .Y(mai_mai_n686_));
  NA3        m0658(.A(mai_mai_n135_), .B(mai_mai_n70_), .C(mai_mai_n33_), .Y(mai_mai_n687_));
  NA3        m0659(.A(mai_mai_n687_), .B(mai_mai_n686_), .C(mai_mai_n684_), .Y(mai_mai_n688_));
  NO4        m0660(.A(mai_mai_n688_), .B(mai_mai_n681_), .C(mai_mai_n677_), .D(mai_mai_n676_), .Y(mai_mai_n689_));
  NA2        m0661(.A(mai_mai_n643_), .B(mai_mai_n31_), .Y(mai_mai_n690_));
  OR2        m0662(.A(mai_mai_n690_), .B(mai_mai_n178_), .Y(mai_mai_n691_));
  NO2        m0663(.A(mai_mai_n480_), .B(mai_mai_n53_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n692_), .B(mai_mai_n664_), .Y(mai_mai_n693_));
  OAI210     m0665(.A0(mai_mai_n634_), .A1(mai_mai_n139_), .B0(mai_mai_n693_), .Y(mai_mai_n694_));
  AN2        m0666(.A(mai_mai_n209_), .B(mai_mai_n637_), .Y(mai_mai_n695_));
  NOi31      m0667(.An(mai_mai_n430_), .B(mai_mai_n653_), .C(j), .Y(mai_mai_n696_));
  NO2        m0668(.A(mai_mai_n695_), .B(mai_mai_n694_), .Y(mai_mai_n697_));
  AO220      m0669(.A0(mai_mai_n359_), .A1(mai_mai_n570_), .B0(mai_mai_n144_), .B1(f), .Y(mai_mai_n698_));
  NA2        m0670(.A(mai_mai_n698_), .B(mai_mai_n683_), .Y(mai_mai_n699_));
  NO2        m0671(.A(mai_mai_n347_), .B(mai_mai_n56_), .Y(mai_mai_n700_));
  OAI210     m0672(.A0(mai_mai_n641_), .A1(mai_mai_n700_), .B0(mai_mai_n538_), .Y(mai_mai_n701_));
  AN4        m0673(.A(mai_mai_n701_), .B(mai_mai_n699_), .C(mai_mai_n697_), .D(mai_mai_n691_), .Y(mai_mai_n702_));
  NA3        m0674(.A(mai_mai_n702_), .B(mai_mai_n689_), .C(mai_mai_n674_), .Y(mai12));
  NO4        m0675(.A(mai_mai_n352_), .B(mai_mai_n210_), .C(mai_mai_n452_), .D(mai_mai_n175_), .Y(mai_mai_n704_));
  NO2        m0676(.A(mai_mai_n357_), .B(mai_mai_n92_), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n506_), .B(mai_mai_n303_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n706_), .B(mai_mai_n429_), .Y(mai_mai_n707_));
  NA2        m0679(.A(mai_mai_n707_), .B(mai_mai_n351_), .Y(mai_mai_n708_));
  AOI210     m0680(.A0(mai_mai_n195_), .A1(mai_mai_n268_), .B0(mai_mai_n166_), .Y(mai_mai_n709_));
  OR2        m0681(.A(mai_mai_n709_), .B(mai_mai_n704_), .Y(mai_mai_n710_));
  NO2        m0682(.A(mai_mai_n315_), .B(mai_mai_n175_), .Y(mai_mai_n711_));
  OAI210     m0683(.A0(mai_mai_n711_), .A1(mai_mai_n710_), .B0(mai_mai_n326_), .Y(mai_mai_n712_));
  INV        m0684(.A(mai_mai_n492_), .Y(mai_mai_n713_));
  NO2        m0685(.A(mai_mai_n458_), .B(mai_mai_n636_), .Y(mai_mai_n714_));
  NA2        m0686(.A(mai_mai_n622_), .B(mai_mai_n713_), .Y(mai_mai_n715_));
  NO2        m0687(.A(mai_mai_n121_), .B(mai_mai_n199_), .Y(mai_mai_n716_));
  NA2        m0688(.A(mai_mai_n715_), .B(mai_mai_n712_), .Y(mai_mai_n717_));
  OR2        m0689(.A(mai_mai_n256_), .B(mai_mai_n705_), .Y(mai_mai_n718_));
  NO3        m0690(.A(mai_mai_n101_), .B(mai_mai_n122_), .C(mai_mai_n175_), .Y(mai_mai_n719_));
  NA2        m0691(.A(mai_mai_n719_), .B(mai_mai_n420_), .Y(mai_mai_n720_));
  INV        m0692(.A(mai_mai_n720_), .Y(mai_mai_n721_));
  NO2        m0693(.A(mai_mai_n508_), .B(mai_mai_n74_), .Y(mai_mai_n722_));
  NO4        m0694(.A(mai_mai_n722_), .B(mai_mai_n721_), .C(mai_mai_n717_), .D(mai_mai_n708_), .Y(mai_mai_n723_));
  NA2        m0695(.A(mai_mai_n436_), .B(mai_mai_n115_), .Y(mai_mai_n724_));
  NOi21      m0696(.An(mai_mai_n33_), .B(mai_mai_n500_), .Y(mai_mai_n725_));
  NA2        m0697(.A(mai_mai_n725_), .B(mai_mai_n724_), .Y(mai_mai_n726_));
  INV        m0698(.A(mai_mai_n726_), .Y(mai_mai_n727_));
  INV        m0699(.A(mai_mai_n291_), .Y(mai_mai_n728_));
  NO2        m0700(.A(mai_mai_n728_), .B(mai_mai_n727_), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n275_), .B(g), .Y(mai_mai_n730_));
  NA2        m0702(.A(h), .B(i), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n731_), .B(mai_mai_n74_), .Y(mai_mai_n732_));
  INV        m0704(.A(mai_mai_n732_), .Y(mai_mai_n733_));
  OAI220     m0705(.A0(mai_mai_n115_), .A1(mai_mai_n730_), .B0(mai_mai_n733_), .B1(mai_mai_n264_), .Y(mai_mai_n734_));
  INV        m0706(.A(mai_mai_n389_), .Y(mai_mai_n735_));
  NO2        m0707(.A(mai_mai_n347_), .B(k), .Y(mai_mai_n736_));
  OAI220     m0708(.A0(mai_mai_n736_), .A1(mai_mai_n735_), .B0(mai_mai_n515_), .B1(mai_mai_n579_), .Y(mai_mai_n737_));
  NA3        m0709(.A(f), .B(k), .C(g), .Y(mai_mai_n738_));
  AOI210     m0710(.A0(mai_mai_n513_), .A1(mai_mai_n738_), .B0(m), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n739_), .B(mai_mai_n256_), .Y(mai_mai_n740_));
  INV        m0712(.A(mai_mai_n348_), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n183_), .B(mai_mai_n62_), .Y(mai_mai_n742_));
  NA2        m0714(.A(mai_mai_n742_), .B(mai_mai_n1098_), .Y(mai_mai_n743_));
  AOI220     m0715(.A0(mai_mai_n743_), .A1(mai_mai_n216_), .B0(mai_mai_n741_), .B1(mai_mai_n69_), .Y(mai_mai_n744_));
  NA3        m0716(.A(mai_mai_n744_), .B(mai_mai_n740_), .C(mai_mai_n737_), .Y(mai_mai_n745_));
  NO2        m0717(.A(mai_mai_n303_), .B(mai_mai_n73_), .Y(mai_mai_n746_));
  NA2        m0718(.A(mai_mai_n746_), .B(mai_mai_n200_), .Y(mai_mai_n747_));
  NA2        m0719(.A(mai_mai_n1097_), .B(mai_mai_n72_), .Y(mai_mai_n748_));
  NO2        m0720(.A(mai_mai_n363_), .B(mai_mai_n175_), .Y(mai_mai_n749_));
  AOI220     m0721(.A0(mai_mai_n749_), .A1(mai_mai_n308_), .B0(mai_mai_n718_), .B1(mai_mai_n179_), .Y(mai_mai_n750_));
  NA2        m0722(.A(mai_mai_n706_), .B(mai_mai_n716_), .Y(mai_mai_n751_));
  NA4        m0723(.A(mai_mai_n751_), .B(mai_mai_n750_), .C(mai_mai_n748_), .D(mai_mai_n747_), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n714_), .B(mai_mai_n429_), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n333_), .B(mai_mai_n624_), .Y(mai_mai_n754_));
  AOI210     m0726(.A0(m), .A1(mai_mai_n424_), .B0(mai_mai_n754_), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n739_), .B(mai_mai_n705_), .Y(mai_mai_n756_));
  INV        m0728(.A(mai_mai_n43_), .Y(mai_mai_n757_));
  AOI220     m0729(.A0(mai_mai_n757_), .A1(mai_mai_n484_), .B0(mai_mai_n496_), .B1(mai_mai_n420_), .Y(mai_mai_n758_));
  NA4        m0730(.A(mai_mai_n758_), .B(mai_mai_n756_), .C(mai_mai_n755_), .D(mai_mai_n753_), .Y(mai_mai_n759_));
  NO4        m0731(.A(mai_mai_n759_), .B(mai_mai_n752_), .C(mai_mai_n745_), .D(mai_mai_n734_), .Y(mai_mai_n760_));
  NAi31      m0732(.An(mai_mai_n111_), .B(mai_mai_n334_), .C(n), .Y(mai_mai_n761_));
  NO2        m0733(.A(mai_mai_n270_), .B(mai_mai_n644_), .Y(mai_mai_n762_));
  NO2        m0734(.A(mai_mai_n762_), .B(mai_mai_n761_), .Y(mai_mai_n763_));
  NO3        m0735(.A(mai_mai_n224_), .B(mai_mai_n111_), .C(mai_mai_n329_), .Y(mai_mai_n764_));
  AOI210     m0736(.A0(mai_mai_n764_), .A1(mai_mai_n390_), .B0(mai_mai_n763_), .Y(mai_mai_n765_));
  NA2        m0737(.A(mai_mai_n383_), .B(i), .Y(mai_mai_n766_));
  NA2        m0738(.A(mai_mai_n766_), .B(mai_mai_n765_), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n192_), .B(mai_mai_n140_), .Y(mai_mai_n768_));
  NA2        m0740(.A(mai_mai_n374_), .B(g), .Y(mai_mai_n769_));
  INV        m0741(.A(mai_mai_n769_), .Y(mai_mai_n770_));
  NO2        m0742(.A(mai_mai_n761_), .B(mai_mai_n195_), .Y(mai_mai_n771_));
  OAI220     m0743(.A0(mai_mai_n706_), .A1(mai_mai_n714_), .B0(mai_mai_n430_), .B1(mai_mai_n340_), .Y(mai_mai_n772_));
  INV        m0744(.A(mai_mai_n772_), .Y(mai_mai_n773_));
  OAI210     m0745(.A0(mai_mai_n709_), .A1(mai_mai_n704_), .B0(mai_mai_n768_), .Y(mai_mai_n774_));
  INV        m0746(.A(mai_mai_n263_), .Y(mai_mai_n775_));
  NA3        m0747(.A(mai_mai_n775_), .B(mai_mai_n774_), .C(mai_mai_n225_), .Y(mai_mai_n776_));
  OR3        m0748(.A(mai_mai_n776_), .B(mai_mai_n773_), .C(mai_mai_n771_), .Y(mai_mai_n777_));
  NO3        m0749(.A(mai_mai_n777_), .B(mai_mai_n770_), .C(mai_mai_n767_), .Y(mai_mai_n778_));
  NA4        m0750(.A(mai_mai_n778_), .B(mai_mai_n760_), .C(mai_mai_n729_), .D(mai_mai_n723_), .Y(mai13));
  NA3        m0751(.A(mai_mai_n209_), .B(b), .C(m), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n387_), .B(f), .Y(mai_mai_n781_));
  NO3        m0753(.A(mai_mai_n781_), .B(mai_mai_n780_), .C(k), .Y(mai_mai_n782_));
  NAi32      m0754(.An(d), .Bn(c), .C(e), .Y(mai_mai_n783_));
  NO4        m0755(.A(i), .B(mai_mai_n783_), .C(mai_mai_n458_), .D(mai_mai_n249_), .Y(mai_mai_n784_));
  AN2        m0756(.A(d), .B(c), .Y(mai_mai_n785_));
  NA2        m0757(.A(mai_mai_n785_), .B(mai_mai_n92_), .Y(mai_mai_n786_));
  NO4        m0758(.A(mai_mai_n786_), .B(mai_mai_n1094_), .C(mai_mai_n145_), .D(mai_mai_n136_), .Y(mai_mai_n787_));
  NA2        m0759(.A(mai_mai_n387_), .B(c), .Y(mai_mai_n788_));
  NO4        m0760(.A(i), .B(mai_mai_n454_), .C(mai_mai_n788_), .D(mai_mai_n249_), .Y(mai_mai_n789_));
  OR2        m0761(.A(mai_mai_n787_), .B(mai_mai_n789_), .Y(mai_mai_n790_));
  OR3        m0762(.A(mai_mai_n790_), .B(mai_mai_n784_), .C(mai_mai_n782_), .Y(mai_mai_n791_));
  NO2        m0763(.A(f), .B(mai_mai_n117_), .Y(mai_mai_n792_));
  NA2        m0764(.A(mai_mai_n792_), .B(g), .Y(mai_mai_n793_));
  OR3        m0765(.A(mai_mai_n186_), .B(mai_mai_n145_), .C(mai_mai_n136_), .Y(mai_mai_n794_));
  NO2        m0766(.A(mai_mai_n794_), .B(mai_mai_n793_), .Y(mai_mai_n795_));
  NO2        m0767(.A(mai_mai_n788_), .B(mai_mai_n249_), .Y(mai_mai_n796_));
  NO2        m0768(.A(j), .B(mai_mai_n41_), .Y(mai_mai_n797_));
  NA2        m0769(.A(mai_mai_n487_), .B(mai_mai_n797_), .Y(mai_mai_n798_));
  NOi21      m0770(.An(mai_mai_n796_), .B(mai_mai_n798_), .Y(mai_mai_n799_));
  NO2        m0771(.A(mai_mai_n580_), .B(mai_mai_n88_), .Y(mai_mai_n800_));
  NOi41      m0772(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n801_), .B(mai_mai_n800_), .Y(mai_mai_n802_));
  NO2        m0774(.A(mai_mai_n802_), .B(mai_mai_n793_), .Y(mai_mai_n803_));
  OR3        m0775(.A(e), .B(d), .C(c), .Y(mai_mai_n804_));
  NA3        m0776(.A(k), .B(j), .C(i), .Y(mai_mai_n805_));
  NO3        m0777(.A(mai_mai_n805_), .B(mai_mai_n249_), .C(mai_mai_n73_), .Y(mai_mai_n806_));
  NOi21      m0778(.An(mai_mai_n806_), .B(mai_mai_n804_), .Y(mai_mai_n807_));
  OR4        m0779(.A(mai_mai_n807_), .B(mai_mai_n803_), .C(mai_mai_n799_), .D(mai_mai_n795_), .Y(mai_mai_n808_));
  NA3        m0780(.A(mai_mai_n367_), .B(mai_mai_n266_), .C(mai_mai_n49_), .Y(mai_mai_n809_));
  NO2        m0781(.A(mai_mai_n809_), .B(mai_mai_n798_), .Y(mai_mai_n810_));
  NO3        m0782(.A(mai_mai_n809_), .B(mai_mai_n454_), .C(mai_mai_n356_), .Y(mai_mai_n811_));
  NO2        m0783(.A(f), .B(c), .Y(mai_mai_n812_));
  NOi21      m0784(.An(mai_mai_n812_), .B(mai_mai_n352_), .Y(mai_mai_n813_));
  NA2        m0785(.A(mai_mai_n813_), .B(mai_mai_n52_), .Y(mai_mai_n814_));
  NO3        m0786(.A(i), .B(h), .C(l), .Y(mai_mai_n815_));
  NOi31      m0787(.An(mai_mai_n815_), .B(mai_mai_n814_), .C(j), .Y(mai_mai_n816_));
  OR3        m0788(.A(mai_mai_n816_), .B(mai_mai_n811_), .C(mai_mai_n810_), .Y(mai_mai_n817_));
  OR3        m0789(.A(mai_mai_n817_), .B(mai_mai_n808_), .C(mai_mai_n791_), .Y(mai02));
  OR3        m0790(.A(n), .B(m), .C(i), .Y(mai_mai_n819_));
  NO4        m0791(.A(mai_mai_n819_), .B(h), .C(l), .D(mai_mai_n804_), .Y(mai_mai_n820_));
  NOi31      m0792(.An(e), .B(d), .C(c), .Y(mai_mai_n821_));
  AOI210     m0793(.A0(mai_mai_n806_), .A1(mai_mai_n821_), .B0(mai_mai_n784_), .Y(mai_mai_n822_));
  AN3        m0794(.A(g), .B(f), .C(c), .Y(mai_mai_n823_));
  INV        m0795(.A(mai_mai_n823_), .Y(mai_mai_n824_));
  OR2        m0796(.A(mai_mai_n805_), .B(mai_mai_n249_), .Y(mai_mai_n825_));
  OR2        m0797(.A(mai_mai_n825_), .B(mai_mai_n824_), .Y(mai_mai_n826_));
  NO3        m0798(.A(mai_mai_n809_), .B(i), .C(mai_mai_n454_), .Y(mai_mai_n827_));
  NO2        m0799(.A(mai_mai_n827_), .B(mai_mai_n795_), .Y(mai_mai_n828_));
  NA3        m0800(.A(l), .B(k), .C(j), .Y(mai_mai_n829_));
  NA2        m0801(.A(i), .B(h), .Y(mai_mai_n830_));
  NO3        m0802(.A(mai_mai_n830_), .B(mai_mai_n829_), .C(mai_mai_n101_), .Y(mai_mai_n831_));
  NO3        m0803(.A(mai_mai_n112_), .B(mai_mai_n234_), .C(mai_mai_n175_), .Y(mai_mai_n832_));
  AOI210     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n831_), .B0(mai_mai_n799_), .Y(mai_mai_n833_));
  NA3        m0805(.A(c), .B(b), .C(a), .Y(mai_mai_n834_));
  INV        m0806(.A(mai_mai_n834_), .Y(mai_mai_n835_));
  NO2        m0807(.A(mai_mai_n805_), .B(mai_mai_n43_), .Y(mai_mai_n836_));
  AOI210     m0808(.A0(mai_mai_n836_), .A1(mai_mai_n835_), .B0(mai_mai_n810_), .Y(mai_mai_n837_));
  AN4        m0809(.A(mai_mai_n837_), .B(mai_mai_n833_), .C(mai_mai_n828_), .D(mai_mai_n826_), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n802_), .B(mai_mai_n794_), .Y(mai_mai_n839_));
  AOI210     m0811(.A0(mai_mai_n839_), .A1(e), .B0(mai_mai_n782_), .Y(mai_mai_n840_));
  NAi41      m0812(.An(mai_mai_n820_), .B(mai_mai_n840_), .C(mai_mai_n838_), .D(mai_mai_n822_), .Y(mai03));
  NOi41      m0813(.An(mai_mai_n614_), .B(mai_mai_n647_), .C(mai_mai_n639_), .D(mai_mai_n36_), .Y(mai_mai_n842_));
  OAI220     m0814(.A0(mai_mai_n842_), .A1(mai_mai_n528_), .B0(mai_mai_n294_), .B1(mai_mai_n455_), .Y(mai_mai_n843_));
  NA4        m0815(.A(i), .B(mai_mai_n821_), .C(mai_mai_n272_), .D(mai_mai_n266_), .Y(mai_mai_n844_));
  INV        m0816(.A(mai_mai_n844_), .Y(mai_mai_n845_));
  NOi31      m0817(.An(m), .B(n), .C(f), .Y(mai_mai_n846_));
  NA2        m0818(.A(mai_mai_n846_), .B(mai_mai_n45_), .Y(mai_mai_n847_));
  AN2        m0819(.A(e), .B(c), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n848_), .B(a), .Y(mai_mai_n849_));
  OAI220     m0821(.A0(mai_mai_n849_), .A1(mai_mai_n847_), .B0(mai_mai_n672_), .B1(mai_mai_n339_), .Y(mai_mai_n850_));
  NOi31      m0822(.An(g), .B(mai_mai_n780_), .C(h), .Y(mai_mai_n851_));
  NO4        m0823(.A(mai_mai_n851_), .B(mai_mai_n850_), .C(mai_mai_n845_), .D(mai_mai_n754_), .Y(mai_mai_n852_));
  INV        m0824(.A(mai_mai_n784_), .Y(mai_mai_n853_));
  NO2        m0825(.A(mai_mai_n830_), .B(mai_mai_n376_), .Y(mai_mai_n854_));
  NO2        m0826(.A(mai_mai_n71_), .B(g), .Y(mai_mai_n855_));
  NO2        m0827(.A(mai_mai_n854_), .B(mai_mai_n815_), .Y(mai_mai_n856_));
  OR2        m0828(.A(mai_mai_n856_), .B(mai_mai_n814_), .Y(mai_mai_n857_));
  NA3        m0829(.A(mai_mai_n857_), .B(mai_mai_n853_), .C(mai_mai_n852_), .Y(mai_mai_n858_));
  NO4        m0830(.A(mai_mai_n858_), .B(mai_mai_n843_), .C(mai_mai_n626_), .D(mai_mai_n443_), .Y(mai_mai_n859_));
  NA2        m0831(.A(c), .B(b), .Y(mai_mai_n860_));
  NO2        m0832(.A(mai_mai_n537_), .B(mai_mai_n860_), .Y(mai_mai_n861_));
  NO2        m0833(.A(mai_mai_n653_), .B(mai_mai_n1095_), .Y(mai_mai_n862_));
  OAI210     m0834(.A0(mai_mai_n862_), .A1(mai_mai_n654_), .B0(mai_mai_n861_), .Y(mai_mai_n863_));
  NAi21      m0835(.An(mai_mai_n335_), .B(mai_mai_n861_), .Y(mai_mai_n864_));
  NA3        m0836(.A(mai_mai_n340_), .B(mai_mai_n438_), .C(f), .Y(mai_mai_n865_));
  NA2        m0837(.A(mai_mai_n865_), .B(mai_mai_n864_), .Y(mai_mai_n866_));
  NAi21      m0838(.An(f), .B(d), .Y(mai_mai_n867_));
  NO2        m0839(.A(mai_mai_n867_), .B(mai_mai_n834_), .Y(mai_mai_n868_));
  AOI210     m0840(.A0(mai_mai_n868_), .A1(mai_mai_n89_), .B0(mai_mai_n866_), .Y(mai_mai_n869_));
  INV        m0841(.A(mai_mai_n199_), .Y(mai_mai_n870_));
  NA2        m0842(.A(mai_mai_n870_), .B(m), .Y(mai_mai_n871_));
  NO2        m0843(.A(mai_mai_n118_), .B(mai_mai_n871_), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n440_), .B(mai_mai_n330_), .Y(mai_mai_n873_));
  NO2        m0845(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n874_));
  NAi21      m0846(.An(mai_mai_n874_), .B(mai_mai_n873_), .Y(mai_mai_n875_));
  NO2        m0847(.A(mai_mai_n875_), .B(mai_mai_n872_), .Y(mai_mai_n876_));
  NA4        m0848(.A(mai_mai_n876_), .B(mai_mai_n869_), .C(mai_mai_n863_), .D(mai_mai_n859_), .Y(mai00));
  INV        m0849(.A(mai_mai_n827_), .Y(mai_mai_n878_));
  NA3        m0850(.A(mai_mai_n878_), .B(mai_mai_n844_), .C(mai_mai_n755_), .Y(mai_mai_n879_));
  NA2        m0851(.A(mai_mai_n400_), .B(f), .Y(mai_mai_n880_));
  NA3        m0852(.A(mai_mai_n644_), .B(mai_mai_n215_), .C(n), .Y(mai_mai_n881_));
  AOI210     m0853(.A0(mai_mai_n881_), .A1(mai_mai_n880_), .B0(mai_mai_n786_), .Y(mai_mai_n882_));
  NO3        m0854(.A(mai_mai_n882_), .B(mai_mai_n879_), .C(mai_mai_n808_), .Y(mai_mai_n883_));
  NA3        m0855(.A(mai_mai_n135_), .B(mai_mai_n42_), .C(mai_mai_n41_), .Y(mai_mai_n884_));
  NA2        m0856(.A(d), .B(b), .Y(mai_mai_n885_));
  NO2        m0857(.A(mai_mai_n885_), .B(mai_mai_n884_), .Y(mai_mai_n886_));
  NO3        m0858(.A(mai_mai_n886_), .B(mai_mai_n874_), .C(mai_mai_n696_), .Y(mai_mai_n887_));
  NO4        m0859(.A(mai_mai_n379_), .B(mai_mai_n282_), .C(mai_mai_n860_), .D(mai_mai_n52_), .Y(mai_mai_n888_));
  NA3        m0860(.A(mai_mai_n309_), .B(mai_mai_n182_), .C(g), .Y(mai_mai_n889_));
  OR2        m0861(.A(mai_mai_n310_), .B(mai_mai_n104_), .Y(mai_mai_n890_));
  NO2        m0862(.A(h), .B(g), .Y(mai_mai_n891_));
  NA4        m0863(.A(mai_mai_n390_), .B(mai_mai_n367_), .C(mai_mai_n891_), .D(b), .Y(mai_mai_n892_));
  NA2        m0864(.A(mai_mai_n719_), .B(b), .Y(mai_mai_n893_));
  AOI220     m0865(.A0(mai_mai_n253_), .A1(mai_mai_n206_), .B0(mai_mai_n146_), .B1(mai_mai_n119_), .Y(mai_mai_n894_));
  NA4        m0866(.A(mai_mai_n894_), .B(mai_mai_n893_), .C(mai_mai_n892_), .D(mai_mai_n890_), .Y(mai_mai_n895_));
  NO3        m0867(.A(mai_mai_n895_), .B(mai_mai_n888_), .C(mai_mai_n219_), .Y(mai_mai_n896_));
  NA2        m0868(.A(mai_mai_n206_), .B(mai_mai_n275_), .Y(mai_mai_n897_));
  NA2        m0869(.A(mai_mai_n897_), .B(mai_mai_n124_), .Y(mai_mai_n898_));
  NA3        m0870(.A(mai_mai_n148_), .B(mai_mai_n88_), .C(g), .Y(mai_mai_n899_));
  NOi31      m0871(.An(c), .B(mai_mai_n1099_), .C(mai_mai_n899_), .Y(mai_mai_n900_));
  NAi21      m0872(.An(mai_mai_n152_), .B(mai_mai_n651_), .Y(mai_mai_n901_));
  NAi21      m0873(.An(mai_mai_n900_), .B(mai_mai_n901_), .Y(mai_mai_n902_));
  INV        m0874(.A(mai_mai_n820_), .Y(mai_mai_n903_));
  NAi21      m0875(.An(mai_mai_n789_), .B(mai_mai_n903_), .Y(mai_mai_n904_));
  NO3        m0876(.A(mai_mai_n904_), .B(mai_mai_n902_), .C(mai_mai_n898_), .Y(mai_mai_n905_));
  AN3        m0877(.A(mai_mai_n905_), .B(mai_mai_n896_), .C(mai_mai_n887_), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n424_), .B(m), .Y(mai_mai_n907_));
  NA3        m0879(.A(mai_mai_n441_), .B(mai_mai_n907_), .C(mai_mai_n203_), .Y(mai_mai_n908_));
  OR4        m0880(.A(mai_mai_n786_), .B(mai_mai_n224_), .C(mai_mai_n184_), .D(e), .Y(mai_mai_n909_));
  AOI220     m0881(.A0(b), .A1(mai_mai_n226_), .B0(mai_mai_n643_), .B1(mai_mai_n176_), .Y(mai_mai_n910_));
  NA2        m0882(.A(mai_mai_n910_), .B(mai_mai_n909_), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n54_), .B(h), .Y(mai_mai_n912_));
  NO3        m0884(.A(mai_mai_n786_), .B(mai_mai_n1094_), .C(mai_mai_n558_), .Y(mai_mai_n913_));
  OAI210     m0885(.A0(mai_mai_n832_), .A1(mai_mai_n913_), .B0(mai_mai_n912_), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n914_), .B(mai_mai_n657_), .Y(mai_mai_n915_));
  NO4        m0887(.A(mai_mai_n915_), .B(mai_mai_n911_), .C(mai_mai_n238_), .D(mai_mai_n908_), .Y(mai_mai_n916_));
  NA2        m0888(.A(e), .B(mai_mai_n578_), .Y(mai_mai_n917_));
  NA4        m0889(.A(mai_mai_n917_), .B(mai_mai_n916_), .C(mai_mai_n906_), .D(mai_mai_n883_), .Y(mai01));
  NO2        m0890(.A(mai_mai_n606_), .B(mai_mai_n232_), .Y(mai_mai_n919_));
  INV        m0891(.A(mai_mai_n919_), .Y(mai_mai_n920_));
  NA2        m0892(.A(mai_mai_n693_), .B(mai_mai_n265_), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n1100_), .B(mai_mai_n1090_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n922_), .B(mai_mai_n490_), .Y(mai_mai_n923_));
  INV        m0895(.A(k), .Y(mai_mai_n924_));
  OR2        m0896(.A(mai_mai_n924_), .B(mai_mai_n453_), .Y(mai_mai_n925_));
  NAi41      m0897(.An(mai_mai_n132_), .B(mai_mai_n925_), .C(mai_mai_n923_), .D(mai_mai_n680_), .Y(mai_mai_n926_));
  NO3        m0898(.A(mai_mai_n596_), .B(mai_mai_n514_), .C(mai_mai_n402_), .Y(mai_mai_n927_));
  OR2        m0899(.A(mai_mai_n160_), .B(mai_mai_n158_), .Y(mai_mai_n928_));
  NA3        m0900(.A(mai_mai_n928_), .B(mai_mai_n927_), .C(mai_mai_n107_), .Y(mai_mai_n929_));
  NO4        m0901(.A(mai_mai_n929_), .B(mai_mai_n926_), .C(mai_mai_n921_), .D(mai_mai_n920_), .Y(mai_mai_n930_));
  NA2        m0902(.A(mai_mai_n427_), .B(mai_mai_n322_), .Y(mai_mai_n931_));
  NOi21      m0903(.An(mai_mai_n442_), .B(mai_mai_n452_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n932_), .B(mai_mai_n931_), .Y(mai_mai_n933_));
  NA2        m0905(.A(mai_mai_n617_), .B(mai_mai_n168_), .Y(mai_mai_n934_));
  OAI210     m0906(.A0(mai_mai_n285_), .A1(mai_mai_n33_), .B0(k), .Y(mai_mai_n935_));
  OR2        m0907(.A(mai_mai_n935_), .B(mai_mai_n264_), .Y(mai_mai_n936_));
  NA4        m0908(.A(mai_mai_n936_), .B(mai_mai_n934_), .C(mai_mai_n933_), .D(mai_mai_n889_), .Y(mai_mai_n937_));
  AOI210     m0909(.A0(mai_mai_n461_), .A1(k), .B0(mai_mai_n464_), .Y(mai_mai_n938_));
  OAI210     m0910(.A0(mai_mai_n924_), .A1(mai_mai_n457_), .B0(mai_mai_n938_), .Y(mai_mai_n939_));
  NA2        m0911(.A(mai_mai_n258_), .B(mai_mai_n515_), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n940_), .B(mai_mai_n599_), .Y(mai_mai_n941_));
  NO3        m0913(.A(mai_mai_n941_), .B(mai_mai_n939_), .C(mai_mai_n937_), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n397_), .B(mai_mai_n51_), .Y(mai_mai_n943_));
  NA3        m0915(.A(mai_mai_n884_), .B(mai_mai_n943_), .C(mai_mai_n577_), .Y(mai_mai_n944_));
  NO2        m0916(.A(mai_mai_n731_), .B(mai_mai_n194_), .Y(mai_mai_n945_));
  NO3        m0917(.A(mai_mai_n64_), .B(mai_mai_n243_), .C(mai_mai_n41_), .Y(mai_mai_n946_));
  NA2        m0918(.A(mai_mai_n946_), .B(mai_mai_n435_), .Y(mai_mai_n947_));
  NA2        m0919(.A(mai_mai_n947_), .B(mai_mai_n511_), .Y(mai_mai_n948_));
  NO2        m0920(.A(mai_mai_n295_), .B(mai_mai_n58_), .Y(mai_mai_n949_));
  INV        m0921(.A(mai_mai_n949_), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n946_), .B(n), .Y(mai_mai_n951_));
  NA3        m0923(.A(mai_mai_n951_), .B(mai_mai_n950_), .C(mai_mai_n312_), .Y(mai_mai_n952_));
  NO3        m0924(.A(mai_mai_n952_), .B(mai_mai_n948_), .C(mai_mai_n944_), .Y(mai_mai_n953_));
  NO3        m0925(.A(mai_mai_n830_), .B(mai_mai_n145_), .C(mai_mai_n71_), .Y(mai_mai_n954_));
  NO2        m0926(.A(mai_mai_n476_), .B(mai_mai_n475_), .Y(mai_mai_n955_));
  NO4        m0927(.A(mai_mai_n830_), .B(mai_mai_n955_), .C(mai_mai_n143_), .D(mai_mai_n71_), .Y(mai_mai_n956_));
  NO3        m0928(.A(mai_mai_n956_), .B(mai_mai_n954_), .C(mai_mai_n491_), .Y(mai_mai_n957_));
  NA4        m0929(.A(mai_mai_n957_), .B(mai_mai_n953_), .C(mai_mai_n942_), .D(mai_mai_n930_), .Y(mai06));
  NO2        m0930(.A(mai_mai_n186_), .B(mai_mai_n80_), .Y(mai_mai_n959_));
  OAI210     m0931(.A0(mai_mai_n959_), .A1(mai_mai_n954_), .B0(mai_mai_n308_), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n672_), .B(mai_mai_n960_), .Y(mai_mai_n961_));
  NO3        m0933(.A(mai_mai_n961_), .B(mai_mai_n948_), .C(mai_mai_n214_), .Y(mai_mai_n962_));
  INV        m0934(.A(mai_mai_n945_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n963_), .B(mai_mai_n268_), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n405_), .B(mai_mai_n140_), .Y(mai_mai_n965_));
  NOi21      m0937(.An(mai_mai_n106_), .B(mai_mai_n41_), .Y(mai_mai_n966_));
  NO2        m0938(.A(mai_mai_n469_), .B(mai_mai_n847_), .Y(mai_mai_n967_));
  NO3        m0939(.A(mai_mai_n967_), .B(mai_mai_n966_), .C(mai_mai_n965_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n55_), .B(mai_mai_n968_), .Y(mai_mai_n969_));
  BUFFER     m0941(.A(mai_mai_n725_), .Y(mai_mai_n970_));
  NO3        m0942(.A(mai_mai_n970_), .B(mai_mai_n969_), .C(mai_mai_n964_), .Y(mai_mai_n971_));
  NO3        m0943(.A(h), .B(mai_mai_n80_), .C(mai_mai_n234_), .Y(mai_mai_n972_));
  OAI220     m0944(.A0(mai_mai_n535_), .A1(mai_mai_n207_), .B0(mai_mai_n401_), .B1(mai_mai_n405_), .Y(mai_mai_n973_));
  NO2        m0945(.A(mai_mai_n463_), .B(j), .Y(mai_mai_n974_));
  NO3        m0946(.A(mai_mai_n973_), .B(mai_mai_n972_), .C(mai_mai_n850_), .Y(mai_mai_n975_));
  NAi31      m0947(.An(mai_mai_n571_), .B(mai_mai_n69_), .C(mai_mai_n168_), .Y(mai_mai_n976_));
  NA2        m0948(.A(mai_mai_n976_), .B(mai_mai_n975_), .Y(mai_mai_n977_));
  OR2        m0949(.A(mai_mai_n595_), .B(mai_mai_n428_), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n974_), .B(m), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n979_), .B(mai_mai_n978_), .Y(mai_mai_n980_));
  NO3        m0952(.A(mai_mai_n665_), .B(mai_mai_n393_), .C(mai_mai_n374_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n981_), .B(mai_mai_n951_), .Y(mai_mai_n982_));
  NAi21      m0954(.An(j), .B(i), .Y(mai_mai_n983_));
  NO4        m0955(.A(mai_mai_n955_), .B(mai_mai_n983_), .C(mai_mai_n352_), .D(mai_mai_n197_), .Y(mai_mai_n984_));
  NO4        m0956(.A(mai_mai_n984_), .B(mai_mai_n982_), .C(mai_mai_n980_), .D(mai_mai_n977_), .Y(mai_mai_n985_));
  NA4        m0957(.A(mai_mai_n985_), .B(mai_mai_n971_), .C(mai_mai_n962_), .D(mai_mai_n957_), .Y(mai07));
  NAi21      m0958(.An(f), .B(c), .Y(mai_mai_n987_));
  OR2        m0959(.A(e), .B(d), .Y(mai_mai_n988_));
  NO2        m0960(.A(mai_mai_n486_), .B(mai_mai_n255_), .Y(mai_mai_n989_));
  NA3        m0961(.A(mai_mai_n989_), .B(mai_mai_n797_), .C(mai_mai_n148_), .Y(mai_mai_n990_));
  NOi31      m0962(.An(n), .B(m), .C(b), .Y(mai_mai_n991_));
  NO3        m0963(.A(mai_mai_n101_), .B(mai_mai_n356_), .C(h), .Y(mai_mai_n992_));
  INV        m0964(.A(mai_mai_n990_), .Y(mai_mai_n993_));
  NO2        m0965(.A(k), .B(i), .Y(mai_mai_n994_));
  NA3        m0966(.A(mai_mai_n994_), .B(mai_mai_n679_), .C(mai_mai_n148_), .Y(mai_mai_n995_));
  NA2        m0967(.A(mai_mai_n71_), .B(mai_mai_n41_), .Y(mai_mai_n996_));
  NO2        m0968(.A(mai_mai_n805_), .B(mai_mai_n249_), .Y(mai_mai_n997_));
  INV        m0969(.A(mai_mai_n995_), .Y(mai_mai_n998_));
  NO2        m0970(.A(mai_mai_n998_), .B(mai_mai_n993_), .Y(mai_mai_n999_));
  NO2        m0971(.A(g), .B(c), .Y(mai_mai_n1000_));
  NA2        m0972(.A(mai_mai_n1000_), .B(mai_mai_n153_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(mai_mai_n1001_), .B(mai_mai_n1089_), .Y(mai_mai_n1002_));
  NA2        m0974(.A(mai_mai_n1002_), .B(mai_mai_n148_), .Y(mai_mai_n1003_));
  NO2        m0975(.A(mai_mai_n357_), .B(a), .Y(mai_mai_n1004_));
  NA3        m0976(.A(mai_mai_n1004_), .B(k), .C(mai_mai_n89_), .Y(mai_mai_n1005_));
  NO2        m0977(.A(i), .B(h), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n867_), .B(h), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n108_), .B(mai_mai_n182_), .Y(mai_mai_n1008_));
  NO2        m0980(.A(mai_mai_n1008_), .B(mai_mai_n1007_), .Y(mai_mai_n1009_));
  NOi31      m0981(.An(m), .B(n), .C(b), .Y(mai_mai_n1010_));
  INV        m0982(.A(mai_mai_n1009_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n823_), .B(mai_mai_n367_), .Y(mai_mai_n1012_));
  NO4        m0984(.A(mai_mai_n1012_), .B(mai_mai_n800_), .C(mai_mai_n352_), .D(mai_mai_n41_), .Y(mai_mai_n1013_));
  OAI210     m0985(.A0(mai_mai_n151_), .A1(mai_mai_n415_), .B0(mai_mai_n801_), .Y(mai_mai_n1014_));
  INV        m0986(.A(mai_mai_n1014_), .Y(mai_mai_n1015_));
  NO2        m0987(.A(mai_mai_n1015_), .B(mai_mai_n1013_), .Y(mai_mai_n1016_));
  AN4        m0988(.A(mai_mai_n1016_), .B(mai_mai_n1011_), .C(mai_mai_n1005_), .D(mai_mai_n1003_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n991_), .B(mai_mai_n305_), .Y(mai_mai_n1018_));
  NA2        m0990(.A(mai_mai_n831_), .B(mai_mai_n1012_), .Y(mai_mai_n1019_));
  INV        m0991(.A(mai_mai_n1019_), .Y(mai_mai_n1020_));
  NO4        m0992(.A(mai_mai_n101_), .B(g), .C(f), .D(e), .Y(mai_mai_n1021_));
  NA3        m0993(.A(mai_mai_n994_), .B(mai_mai_n236_), .C(h), .Y(mai_mai_n1022_));
  OR2        m0994(.A(e), .B(a), .Y(mai_mai_n1023_));
  NO2        m0995(.A(mai_mai_n988_), .B(mai_mai_n987_), .Y(mai_mai_n1024_));
  AOI210     m0996(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1024_), .Y(mai_mai_n1025_));
  NO2        m0997(.A(mai_mai_n1025_), .B(mai_mai_n819_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n846_), .B(mai_mai_n329_), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n1026_), .B(mai_mai_n1020_), .Y(mai_mai_n1028_));
  NA3        m1000(.A(mai_mai_n1028_), .B(mai_mai_n1017_), .C(mai_mai_n999_), .Y(mai_mai_n1029_));
  NO2        m1001(.A(mai_mai_n317_), .B(j), .Y(mai_mai_n1030_));
  NAi31      m1002(.An(mai_mai_n1006_), .B(mai_mai_n813_), .C(mai_mai_n136_), .Y(mai_mai_n1031_));
  INV        m1003(.A(mai_mai_n1031_), .Y(mai_mai_n1032_));
  NA3        m1004(.A(g), .B(mai_mai_n1030_), .C(mai_mai_n129_), .Y(mai_mai_n1033_));
  INV        m1005(.A(mai_mai_n1033_), .Y(mai_mai_n1034_));
  NO2        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1032_), .Y(mai_mai_n1035_));
  NA2        m1007(.A(mai_mai_n628_), .B(mai_mai_n159_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n148_), .B(mai_mai_n88_), .Y(mai_mai_n1037_));
  NOi21      m1009(.An(d), .B(f), .Y(mai_mai_n1038_));
  NO2        m1010(.A(mai_mai_n988_), .B(f), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n1036_), .B(mai_mai_n1035_), .Y(mai_mai_n1040_));
  NO3        m1012(.A(mai_mai_n823_), .B(mai_mai_n812_), .C(mai_mai_n39_), .Y(mai_mai_n1041_));
  NA2        m1013(.A(mai_mai_n1041_), .B(mai_mai_n997_), .Y(mai_mai_n1042_));
  OAI210     m1014(.A0(mai_mai_n1021_), .A1(mai_mai_n991_), .B0(mai_mai_n669_), .Y(mai_mai_n1043_));
  OAI220     m1015(.A0(mai_mai_n783_), .A1(mai_mai_n101_), .B0(h), .B1(mai_mai_n143_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n1044_), .B(mai_mai_n480_), .Y(mai_mai_n1045_));
  NA3        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1043_), .C(mai_mai_n1042_), .Y(mai_mai_n1046_));
  NA2        m1018(.A(mai_mai_n1000_), .B(mai_mai_n1038_), .Y(mai_mai_n1047_));
  NO2        m1019(.A(mai_mai_n1047_), .B(m), .Y(mai_mai_n1048_));
  NO2        m1020(.A(mai_mai_n121_), .B(mai_mai_n150_), .Y(mai_mai_n1049_));
  OAI210     m1021(.A0(mai_mai_n1049_), .A1(mai_mai_n86_), .B0(mai_mai_n1010_), .Y(mai_mai_n1050_));
  INV        m1022(.A(mai_mai_n1050_), .Y(mai_mai_n1051_));
  NO3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1048_), .C(mai_mai_n1046_), .Y(mai_mai_n1052_));
  NO2        m1024(.A(mai_mai_n987_), .B(e), .Y(mai_mai_n1053_));
  NA2        m1025(.A(mai_mai_n855_), .B(mai_mai_n489_), .Y(mai_mai_n1054_));
  NO2        m1026(.A(mai_mai_n1054_), .B(mai_mai_n354_), .Y(mai_mai_n1055_));
  INV        m1027(.A(mai_mai_n1055_), .Y(mai_mai_n1056_));
  NO2        m1028(.A(mai_mai_n150_), .B(c), .Y(mai_mai_n1057_));
  OAI210     m1029(.A0(mai_mai_n1057_), .A1(mai_mai_n1053_), .B0(mai_mai_n148_), .Y(mai_mai_n1058_));
  AOI220     m1030(.A0(mai_mai_n1058_), .A1(mai_mai_n814_), .B0(mai_mai_n421_), .B1(mai_mai_n293_), .Y(mai_mai_n1059_));
  NO2        m1031(.A(mai_mai_n1023_), .B(f), .Y(mai_mai_n1060_));
  AOI210     m1032(.A0(mai_mai_n682_), .A1(mai_mai_n332_), .B0(mai_mai_n82_), .Y(mai_mai_n1061_));
  NA2        m1033(.A(mai_mai_n1060_), .B(mai_mai_n996_), .Y(mai_mai_n1062_));
  OAI220     m1034(.A0(mai_mai_n1062_), .A1(mai_mai_n43_), .B0(mai_mai_n1061_), .B1(mai_mai_n143_), .Y(mai_mai_n1063_));
  NA2        m1035(.A(mai_mai_n992_), .B(mai_mai_n151_), .Y(mai_mai_n1064_));
  INV        m1036(.A(mai_mai_n1064_), .Y(mai_mai_n1065_));
  NO3        m1037(.A(mai_mai_n1065_), .B(mai_mai_n1063_), .C(mai_mai_n1059_), .Y(mai_mai_n1066_));
  NA3        m1038(.A(mai_mai_n1066_), .B(mai_mai_n1056_), .C(mai_mai_n1052_), .Y(mai_mai_n1067_));
  AO210      m1039(.A0(mai_mai_n102_), .A1(l), .B0(mai_mai_n1018_), .Y(mai_mai_n1068_));
  NO2        m1040(.A(mai_mai_n127_), .B(mai_mai_n1053_), .Y(mai_mai_n1069_));
  NO2        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1037_), .Y(mai_mai_n1070_));
  NOi21      m1042(.An(mai_mai_n992_), .B(e), .Y(mai_mai_n1071_));
  NO2        m1043(.A(mai_mai_n1071_), .B(mai_mai_n1070_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n52_), .B(a), .Y(mai_mai_n1073_));
  NO2        m1045(.A(mai_mai_n1027_), .B(mai_mai_n1073_), .Y(mai_mai_n1074_));
  INV        m1046(.A(mai_mai_n1074_), .Y(mai_mai_n1075_));
  NA3        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1072_), .C(mai_mai_n1068_), .Y(mai_mai_n1076_));
  OR4        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1067_), .C(mai_mai_n1040_), .D(mai_mai_n1029_), .Y(mai04));
  NOi31      m1049(.An(mai_mai_n1021_), .B(mai_mai_n1022_), .C(mai_mai_n786_), .Y(mai_mai_n1078_));
  NA2        m1050(.A(mai_mai_n1039_), .B(mai_mai_n628_), .Y(mai_mai_n1079_));
  NO2        m1051(.A(mai_mai_n1079_), .B(j), .Y(mai_mai_n1080_));
  OR3        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1078_), .C(mai_mai_n803_), .Y(mai_mai_n1081_));
  INV        m1053(.A(mai_mai_n73_), .Y(mai_mai_n1082_));
  AOI210     m1054(.A0(mai_mai_n1082_), .A1(mai_mai_n796_), .B0(mai_mai_n900_), .Y(mai_mai_n1083_));
  NA2        m1055(.A(mai_mai_n1083_), .B(mai_mai_n914_), .Y(mai_mai_n1084_));
  NO4        m1056(.A(mai_mai_n1084_), .B(mai_mai_n1081_), .C(mai_mai_n811_), .D(mai_mai_n791_), .Y(mai_mai_n1085_));
  NA4        m1057(.A(mai_mai_n1085_), .B(mai_mai_n857_), .C(mai_mai_n844_), .D(mai_mai_n838_), .Y(mai05));
  INV        m1058(.A(l), .Y(mai_mai_n1089_));
  INV        m1059(.A(f), .Y(mai_mai_n1090_));
  INV        m1060(.A(mai_mai_n420_), .Y(mai_mai_n1091_));
  INV        m1061(.A(mai_mai_n89_), .Y(mai_mai_n1092_));
  INV        m1062(.A(e), .Y(mai_mai_n1093_));
  INV        m1063(.A(e), .Y(mai_mai_n1094_));
  INV        m1064(.A(mai_mai_n633_), .Y(mai_mai_n1095_));
  INV        m1065(.A(mai_mai_n53_), .Y(mai_mai_n1096_));
  INV        m1066(.A(mai_mai_n455_), .Y(mai_mai_n1097_));
  INV        m1067(.A(g), .Y(mai_mai_n1098_));
  INV        m1068(.A(e), .Y(mai_mai_n1099_));
  INV        m1069(.A(k), .Y(mai_mai_n1100_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NAi21      u0031(.An(i), .B(h), .Y(men_men_n60_));
  NAi31      u0032(.An(i), .B(l), .C(j), .Y(men_men_n61_));
  OAI220     u0033(.A0(men_men_n61_), .A1(men_men_n49_), .B0(men_men_n60_), .B1(men_men_n44_), .Y(men_men_n62_));
  NAi31      u0034(.An(d), .B(men_men_n62_), .C(men_men_n58_), .Y(men_men_n63_));
  NAi41      u0035(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n64_));
  NA2        u0036(.A(g), .B(f), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi21      u0038(.An(i), .B(j), .Y(men_men_n67_));
  NAi32      u0039(.An(n), .Bn(k), .C(m), .Y(men_men_n68_));
  NO2        u0040(.A(men_men_n68_), .B(men_men_n67_), .Y(men_men_n69_));
  NAi31      u0041(.An(l), .B(m), .C(k), .Y(men_men_n70_));
  NAi21      u0042(.An(e), .B(h), .Y(men_men_n71_));
  NAi41      u0043(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n73_));
  INV        u0045(.A(m), .Y(men_men_n74_));
  NOi21      u0046(.An(k), .B(l), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  AN4        u0048(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n77_));
  NOi31      u0049(.An(h), .B(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n77_), .Y(men_men_n79_));
  NAi32      u0051(.An(m), .Bn(k), .C(j), .Y(men_men_n80_));
  NOi32      u0052(.An(h), .Bn(g), .C(f), .Y(men_men_n81_));
  NA2        u0053(.A(men_men_n81_), .B(men_men_n77_), .Y(men_men_n82_));
  OA220      u0054(.A0(men_men_n82_), .A1(men_men_n80_), .B0(men_men_n79_), .B1(men_men_n76_), .Y(men_men_n83_));
  NA3        u0055(.A(men_men_n83_), .B(men_men_n73_), .C(men_men_n63_), .Y(men_men_n84_));
  INV        u0056(.A(n), .Y(men_men_n85_));
  NOi32      u0057(.An(e), .Bn(b), .C(d), .Y(men_men_n86_));
  NA2        u0058(.A(men_men_n86_), .B(men_men_n85_), .Y(men_men_n87_));
  INV        u0059(.A(j), .Y(men_men_n88_));
  AN3        u0060(.A(m), .B(k), .C(i), .Y(men_men_n89_));
  NA3        u0061(.A(men_men_n89_), .B(men_men_n88_), .C(g), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(f), .Y(men_men_n91_));
  NAi32      u0063(.An(g), .Bn(f), .C(h), .Y(men_men_n92_));
  NAi31      u0064(.An(j), .B(m), .C(l), .Y(men_men_n93_));
  NO2        u0065(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  NA2        u0066(.A(m), .B(l), .Y(men_men_n95_));
  NAi31      u0067(.An(k), .B(j), .C(g), .Y(men_men_n96_));
  NO3        u0068(.A(men_men_n96_), .B(men_men_n95_), .C(f), .Y(men_men_n97_));
  AN2        u0069(.A(j), .B(g), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(l), .C(i), .Y(men_men_n99_));
  NOi21      u0071(.An(g), .B(i), .Y(men_men_n100_));
  NOi32      u0072(.An(m), .Bn(j), .C(k), .Y(men_men_n101_));
  AOI220     u0073(.A0(men_men_n101_), .A1(men_men_n100_), .B0(men_men_n99_), .B1(men_men_n98_), .Y(men_men_n102_));
  NO2        u0074(.A(men_men_n102_), .B(f), .Y(men_men_n103_));
  NO4        u0075(.A(men_men_n103_), .B(men_men_n97_), .C(men_men_n94_), .D(men_men_n91_), .Y(men_men_n104_));
  NAi41      u0076(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n105_));
  AN2        u0077(.A(e), .B(b), .Y(men_men_n106_));
  NOi31      u0078(.An(c), .B(h), .C(f), .Y(men_men_n107_));
  NA2        u0079(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NOi21      u0080(.An(g), .B(f), .Y(men_men_n109_));
  NOi21      u0081(.An(i), .B(h), .Y(men_men_n110_));
  NA3        u0082(.A(men_men_n110_), .B(men_men_n109_), .C(men_men_n36_), .Y(men_men_n111_));
  INV        u0083(.A(a), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n106_), .B(men_men_n112_), .Y(men_men_n113_));
  INV        u0085(.A(l), .Y(men_men_n114_));
  NOi21      u0086(.An(m), .B(n), .Y(men_men_n115_));
  NO2        u0087(.A(men_men_n111_), .B(men_men_n87_), .Y(men_men_n116_));
  INV        u0088(.A(b), .Y(men_men_n117_));
  NA2        u0089(.A(l), .B(j), .Y(men_men_n118_));
  AN2        u0090(.A(k), .B(i), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u0092(.A(g), .B(e), .Y(men_men_n121_));
  NOi32      u0093(.An(c), .Bn(a), .C(d), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n115_), .Y(men_men_n123_));
  NO4        u0095(.A(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n124_));
  NO2        u0096(.A(men_men_n124_), .B(men_men_n116_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n104_), .A1(men_men_n87_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n78_), .C(men_men_n77_), .Y(men_men_n128_));
  NOi31      u0100(.An(k), .B(m), .C(i), .Y(men_men_n129_));
  NA3        u0101(.A(men_men_n129_), .B(men_men_n81_), .C(men_men_n77_), .Y(men_men_n130_));
  NA2        u0102(.A(men_men_n130_), .B(men_men_n128_), .Y(men_men_n131_));
  NOi32      u0103(.An(f), .Bn(b), .C(e), .Y(men_men_n132_));
  NAi21      u0104(.An(g), .B(h), .Y(men_men_n133_));
  NAi21      u0105(.An(m), .B(n), .Y(men_men_n134_));
  NAi21      u0106(.An(j), .B(k), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n133_), .Y(men_men_n136_));
  NAi41      u0108(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n137_));
  NAi31      u0109(.An(j), .B(k), .C(h), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n134_), .Y(men_men_n139_));
  AOI210     u0111(.A0(men_men_n136_), .A1(men_men_n132_), .B0(men_men_n139_), .Y(men_men_n140_));
  NO2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  AN2        u0113(.A(k), .B(j), .Y(men_men_n142_));
  NAi21      u0114(.An(c), .B(b), .Y(men_men_n143_));
  NA2        u0115(.A(f), .B(d), .Y(men_men_n144_));
  NO4        u0116(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n142_), .D(men_men_n133_), .Y(men_men_n145_));
  NA2        u0117(.A(h), .B(c), .Y(men_men_n146_));
  NAi31      u0118(.An(f), .B(e), .C(b), .Y(men_men_n147_));
  NA2        u0119(.A(men_men_n145_), .B(n), .Y(men_men_n148_));
  NA2        u0120(.A(d), .B(b), .Y(men_men_n149_));
  NAi21      u0121(.An(e), .B(f), .Y(men_men_n150_));
  NO2        u0122(.A(men_men_n150_), .B(men_men_n149_), .Y(men_men_n151_));
  NA2        u0123(.A(b), .B(a), .Y(men_men_n152_));
  NAi21      u0124(.An(c), .B(d), .Y(men_men_n153_));
  NAi31      u0125(.An(l), .B(k), .C(h), .Y(men_men_n154_));
  NO2        u0126(.A(men_men_n134_), .B(men_men_n154_), .Y(men_men_n155_));
  NA2        u0127(.A(men_men_n155_), .B(men_men_n151_), .Y(men_men_n156_));
  NAi41      u0128(.An(men_men_n131_), .B(men_men_n156_), .C(men_men_n148_), .D(men_men_n140_), .Y(men_men_n157_));
  NAi31      u0129(.An(e), .B(f), .C(b), .Y(men_men_n158_));
  NOi21      u0130(.An(g), .B(d), .Y(men_men_n159_));
  NO2        u0131(.A(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  NOi21      u0132(.An(h), .B(i), .Y(men_men_n161_));
  NOi21      u0133(.An(k), .B(m), .Y(men_men_n162_));
  NA3        u0134(.A(men_men_n162_), .B(men_men_n161_), .C(n), .Y(men_men_n163_));
  NOi21      u0135(.An(men_men_n160_), .B(men_men_n163_), .Y(men_men_n164_));
  NOi21      u0136(.An(h), .B(g), .Y(men_men_n165_));
  NO2        u0137(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n166_));
  NA2        u0138(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  NAi31      u0139(.An(l), .B(j), .C(h), .Y(men_men_n168_));
  NO2        u0140(.A(men_men_n168_), .B(men_men_n49_), .Y(men_men_n169_));
  NA2        u0141(.A(men_men_n169_), .B(men_men_n66_), .Y(men_men_n170_));
  NA2        u0142(.A(l), .B(i), .Y(men_men_n171_));
  NA2        u0143(.A(men_men_n171_), .B(n), .Y(men_men_n172_));
  OAI210     u0144(.A0(men_men_n172_), .A1(men_men_n167_), .B0(men_men_n170_), .Y(men_men_n173_));
  NAi31      u0145(.An(e), .B(f), .C(c), .Y(men_men_n174_));
  NA2        u0146(.A(j), .B(h), .Y(men_men_n175_));
  OR3        u0147(.A(n), .B(m), .C(k), .Y(men_men_n176_));
  NO2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  NAi32      u0149(.An(m), .Bn(k), .C(n), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n175_), .Y(men_men_n179_));
  AOI220     u0151(.A0(men_men_n179_), .A1(men_men_n160_), .B0(men_men_n177_), .B1(f), .Y(men_men_n180_));
  NO2        u0152(.A(n), .B(m), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n50_), .Y(men_men_n182_));
  NAi21      u0154(.An(f), .B(e), .Y(men_men_n183_));
  NA2        u0155(.A(d), .B(c), .Y(men_men_n184_));
  NOi21      u0156(.An(c), .B(men_men_n182_), .Y(men_men_n185_));
  NAi21      u0157(.An(d), .B(c), .Y(men_men_n186_));
  NAi31      u0158(.An(m), .B(n), .C(b), .Y(men_men_n187_));
  NA2        u0159(.A(k), .B(i), .Y(men_men_n188_));
  NAi21      u0160(.An(h), .B(f), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NO2        u0162(.A(men_men_n187_), .B(men_men_n153_), .Y(men_men_n191_));
  NA2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi32      u0164(.An(f), .Bn(c), .C(e), .Y(men_men_n193_));
  NO3        u0165(.A(n), .B(m), .C(j), .Y(men_men_n194_));
  NA2        u0166(.A(men_men_n194_), .B(k), .Y(men_men_n195_));
  NAi31      u0167(.An(men_men_n185_), .B(men_men_n192_), .C(men_men_n180_), .Y(men_men_n196_));
  OR4        u0168(.A(men_men_n196_), .B(men_men_n173_), .C(men_men_n164_), .D(men_men_n157_), .Y(men_men_n197_));
  NO4        u0169(.A(men_men_n197_), .B(men_men_n126_), .C(men_men_n84_), .D(men_men_n55_), .Y(men_men_n198_));
  NA3        u0170(.A(m), .B(men_men_n114_), .C(j), .Y(men_men_n199_));
  NAi31      u0171(.An(n), .B(h), .C(g), .Y(men_men_n200_));
  NO2        u0172(.A(men_men_n200_), .B(men_men_n199_), .Y(men_men_n201_));
  NOi32      u0173(.An(m), .Bn(k), .C(l), .Y(men_men_n202_));
  NA3        u0174(.A(men_men_n202_), .B(men_men_n88_), .C(g), .Y(men_men_n203_));
  NO2        u0175(.A(men_men_n203_), .B(n), .Y(men_men_n204_));
  NOi21      u0176(.An(k), .B(j), .Y(men_men_n205_));
  NA4        u0177(.A(men_men_n205_), .B(men_men_n115_), .C(i), .D(g), .Y(men_men_n206_));
  AN2        u0178(.A(i), .B(g), .Y(men_men_n207_));
  NA3        u0179(.A(men_men_n75_), .B(men_men_n207_), .C(men_men_n115_), .Y(men_men_n208_));
  NA2        u0180(.A(men_men_n208_), .B(men_men_n206_), .Y(men_men_n209_));
  NO3        u0181(.A(men_men_n209_), .B(men_men_n204_), .C(men_men_n201_), .Y(men_men_n210_));
  NAi41      u0182(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n211_));
  INV        u0183(.A(men_men_n211_), .Y(men_men_n212_));
  INV        u0184(.A(f), .Y(men_men_n213_));
  INV        u0185(.A(g), .Y(men_men_n214_));
  NOi31      u0186(.An(i), .B(j), .C(h), .Y(men_men_n215_));
  NOi21      u0187(.An(l), .B(m), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NO3        u0189(.A(men_men_n217_), .B(men_men_n214_), .C(men_men_n213_), .Y(men_men_n218_));
  NA2        u0190(.A(men_men_n218_), .B(men_men_n212_), .Y(men_men_n219_));
  OAI210     u0191(.A0(men_men_n210_), .A1(men_men_n32_), .B0(men_men_n219_), .Y(men_men_n220_));
  NOi21      u0192(.An(n), .B(m), .Y(men_men_n221_));
  NA2        u0193(.A(i), .B(men_men_n221_), .Y(men_men_n222_));
  OA220      u0194(.A0(men_men_n222_), .A1(men_men_n108_), .B0(men_men_n80_), .B1(men_men_n79_), .Y(men_men_n223_));
  NAi21      u0195(.An(j), .B(h), .Y(men_men_n224_));
  XN2        u0196(.A(i), .B(h), .Y(men_men_n225_));
  NOi31      u0197(.An(k), .B(n), .C(m), .Y(men_men_n226_));
  NAi31      u0198(.An(f), .B(e), .C(c), .Y(men_men_n227_));
  NA4        u0199(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n228_));
  NAi32      u0200(.An(m), .Bn(i), .C(k), .Y(men_men_n229_));
  NO3        u0201(.A(men_men_n229_), .B(men_men_n92_), .C(men_men_n228_), .Y(men_men_n230_));
  INV        u0202(.A(k), .Y(men_men_n231_));
  INV        u0203(.A(men_men_n230_), .Y(men_men_n232_));
  NAi21      u0204(.An(n), .B(a), .Y(men_men_n233_));
  NO2        u0205(.A(men_men_n233_), .B(men_men_n149_), .Y(men_men_n234_));
  NAi41      u0206(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n235_));
  NO2        u0207(.A(men_men_n235_), .B(e), .Y(men_men_n236_));
  NO3        u0208(.A(men_men_n150_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n237_));
  OAI210     u0209(.A0(men_men_n237_), .A1(men_men_n236_), .B0(men_men_n234_), .Y(men_men_n238_));
  AN3        u0210(.A(men_men_n238_), .B(men_men_n232_), .C(men_men_n223_), .Y(men_men_n239_));
  OR2        u0211(.A(h), .B(g), .Y(men_men_n240_));
  NO2        u0212(.A(men_men_n240_), .B(men_men_n105_), .Y(men_men_n241_));
  NA2        u0213(.A(men_men_n241_), .B(men_men_n132_), .Y(men_men_n242_));
  NAi41      u0214(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n243_), .B(men_men_n213_), .Y(men_men_n244_));
  NA2        u0216(.A(men_men_n162_), .B(men_men_n110_), .Y(men_men_n245_));
  NAi21      u0217(.An(men_men_n245_), .B(men_men_n244_), .Y(men_men_n246_));
  NO2        u0218(.A(n), .B(a), .Y(men_men_n247_));
  NAi31      u0219(.An(men_men_n235_), .B(men_men_n247_), .C(men_men_n106_), .Y(men_men_n248_));
  AN2        u0220(.A(men_men_n248_), .B(men_men_n246_), .Y(men_men_n249_));
  NAi21      u0221(.An(h), .B(i), .Y(men_men_n250_));
  NA2        u0222(.A(men_men_n249_), .B(men_men_n242_), .Y(men_men_n251_));
  NOi21      u0223(.An(g), .B(e), .Y(men_men_n252_));
  NO2        u0224(.A(men_men_n72_), .B(men_men_n74_), .Y(men_men_n253_));
  NA2        u0225(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NOi32      u0226(.An(l), .Bn(j), .C(i), .Y(men_men_n255_));
  AOI210     u0227(.A0(men_men_n75_), .A1(men_men_n88_), .B0(men_men_n255_), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n250_), .B(men_men_n44_), .Y(men_men_n257_));
  NAi21      u0229(.An(f), .B(g), .Y(men_men_n258_));
  NO2        u0230(.A(men_men_n258_), .B(men_men_n64_), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n68_), .B(men_men_n118_), .Y(men_men_n260_));
  AOI220     u0232(.A0(men_men_n260_), .A1(men_men_n259_), .B0(men_men_n257_), .B1(men_men_n66_), .Y(men_men_n261_));
  OAI210     u0233(.A0(men_men_n256_), .A1(men_men_n254_), .B0(men_men_n261_), .Y(men_men_n262_));
  NO3        u0234(.A(men_men_n135_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n263_));
  NOi41      u0235(.An(men_men_n239_), .B(men_men_n262_), .C(men_men_n251_), .D(men_men_n220_), .Y(men_men_n264_));
  NO4        u0236(.A(men_men_n201_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n265_), .B(men_men_n113_), .Y(men_men_n266_));
  NA3        u0238(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n267_));
  NAi21      u0239(.An(h), .B(g), .Y(men_men_n268_));
  OR4        u0240(.A(men_men_n268_), .B(men_men_n267_), .C(men_men_n222_), .D(e), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n245_), .B(men_men_n258_), .Y(men_men_n270_));
  NAi31      u0242(.An(g), .B(k), .C(h), .Y(men_men_n271_));
  NO3        u0243(.A(men_men_n134_), .B(men_men_n271_), .C(l), .Y(men_men_n272_));
  NAi31      u0244(.An(e), .B(d), .C(a), .Y(men_men_n273_));
  NA2        u0245(.A(men_men_n272_), .B(men_men_n132_), .Y(men_men_n274_));
  NA2        u0246(.A(men_men_n274_), .B(men_men_n269_), .Y(men_men_n275_));
  NA4        u0247(.A(men_men_n162_), .B(men_men_n81_), .C(men_men_n77_), .D(men_men_n118_), .Y(men_men_n276_));
  NA2        u0248(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n277_));
  NA3        u0249(.A(e), .B(c), .C(b), .Y(men_men_n278_));
  NO2        u0250(.A(d), .B(men_men_n278_), .Y(men_men_n279_));
  NAi32      u0251(.An(k), .Bn(i), .C(j), .Y(men_men_n280_));
  NAi31      u0252(.An(h), .B(l), .C(i), .Y(men_men_n281_));
  NA3        u0253(.A(men_men_n281_), .B(men_men_n280_), .C(men_men_n168_), .Y(men_men_n282_));
  NOi21      u0254(.An(men_men_n282_), .B(men_men_n49_), .Y(men_men_n283_));
  OAI210     u0255(.A0(men_men_n259_), .A1(men_men_n279_), .B0(men_men_n283_), .Y(men_men_n284_));
  NAi21      u0256(.An(l), .B(k), .Y(men_men_n285_));
  NO2        u0257(.A(men_men_n285_), .B(men_men_n49_), .Y(men_men_n286_));
  NOi21      u0258(.An(l), .B(j), .Y(men_men_n287_));
  NA2        u0259(.A(men_men_n165_), .B(men_men_n287_), .Y(men_men_n288_));
  NA3        u0260(.A(men_men_n119_), .B(men_men_n118_), .C(g), .Y(men_men_n289_));
  OR3        u0261(.A(men_men_n72_), .B(men_men_n74_), .C(e), .Y(men_men_n290_));
  AOI210     u0262(.A0(men_men_n289_), .A1(men_men_n288_), .B0(men_men_n290_), .Y(men_men_n291_));
  INV        u0263(.A(men_men_n291_), .Y(men_men_n292_));
  NAi32      u0264(.An(j), .Bn(h), .C(i), .Y(men_men_n293_));
  NAi21      u0265(.An(m), .B(l), .Y(men_men_n294_));
  NO2        u0266(.A(men_men_n294_), .B(men_men_n293_), .Y(men_men_n295_));
  NA2        u0267(.A(h), .B(g), .Y(men_men_n296_));
  NA2        u0268(.A(n), .B(men_men_n45_), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n297_), .B(men_men_n296_), .Y(men_men_n298_));
  OAI210     u0270(.A0(men_men_n298_), .A1(men_men_n295_), .B0(men_men_n166_), .Y(men_men_n299_));
  NA4        u0271(.A(men_men_n299_), .B(men_men_n292_), .C(men_men_n284_), .D(men_men_n276_), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n147_), .B(d), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n301_), .B(men_men_n53_), .Y(men_men_n302_));
  NAi32      u0274(.An(n), .Bn(m), .C(l), .Y(men_men_n303_));
  NO2        u0275(.A(men_men_n303_), .B(men_men_n293_), .Y(men_men_n304_));
  INV        u0276(.A(men_men_n304_), .Y(men_men_n305_));
  NO2        u0277(.A(men_men_n123_), .B(men_men_n117_), .Y(men_men_n306_));
  NAi31      u0278(.An(k), .B(l), .C(j), .Y(men_men_n307_));
  OAI210     u0279(.A0(men_men_n285_), .A1(j), .B0(men_men_n307_), .Y(men_men_n308_));
  NOi21      u0280(.An(men_men_n308_), .B(men_men_n121_), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n309_), .B(men_men_n306_), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n310_), .B(men_men_n302_), .Y(men_men_n311_));
  NO4        u0283(.A(men_men_n311_), .B(men_men_n300_), .C(men_men_n275_), .D(men_men_n266_), .Y(men_men_n312_));
  NAi21      u0284(.An(m), .B(k), .Y(men_men_n313_));
  NO2        u0285(.A(men_men_n225_), .B(men_men_n313_), .Y(men_men_n314_));
  NAi41      u0286(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n315_));
  NAi31      u0287(.An(i), .B(l), .C(h), .Y(men_men_n316_));
  NO4        u0288(.A(men_men_n316_), .B(e), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n317_));
  NA2        u0289(.A(e), .B(c), .Y(men_men_n318_));
  NOi21      u0290(.An(f), .B(h), .Y(men_men_n319_));
  NA2        u0291(.A(men_men_n319_), .B(men_men_n119_), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n214_), .Y(men_men_n321_));
  NAi31      u0293(.An(d), .B(e), .C(b), .Y(men_men_n322_));
  NO2        u0294(.A(men_men_n134_), .B(men_men_n322_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n321_), .Y(men_men_n324_));
  NAi21      u0296(.An(men_men_n317_), .B(men_men_n324_), .Y(men_men_n325_));
  NO4        u0297(.A(men_men_n315_), .B(men_men_n80_), .C(men_men_n71_), .D(men_men_n214_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n247_), .B(men_men_n106_), .Y(men_men_n327_));
  OR2        u0299(.A(men_men_n327_), .B(men_men_n203_), .Y(men_men_n328_));
  NOi31      u0300(.An(l), .B(n), .C(m), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n329_), .B(men_men_n215_), .Y(men_men_n330_));
  INV        u0302(.A(men_men_n330_), .Y(men_men_n331_));
  NAi32      u0303(.An(men_men_n331_), .Bn(men_men_n326_), .C(men_men_n328_), .Y(men_men_n332_));
  NAi32      u0304(.An(m), .Bn(j), .C(k), .Y(men_men_n333_));
  NAi41      u0305(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n334_));
  OAI210     u0306(.A0(men_men_n211_), .A1(men_men_n333_), .B0(men_men_n334_), .Y(men_men_n335_));
  NOi31      u0307(.An(j), .B(m), .C(k), .Y(men_men_n336_));
  NO2        u0308(.A(men_men_n127_), .B(men_men_n336_), .Y(men_men_n337_));
  AN3        u0309(.A(h), .B(g), .C(f), .Y(men_men_n338_));
  NAi31      u0310(.An(men_men_n337_), .B(men_men_n338_), .C(men_men_n335_), .Y(men_men_n339_));
  NOi32      u0311(.An(m), .Bn(j), .C(l), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n340_), .B(men_men_n99_), .Y(men_men_n341_));
  NAi32      u0313(.An(men_men_n341_), .Bn(men_men_n200_), .C(men_men_n301_), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n294_), .B(men_men_n293_), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n217_), .B(g), .Y(men_men_n344_));
  INV        u0316(.A(men_men_n158_), .Y(men_men_n345_));
  AOI220     u0317(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n244_), .B1(men_men_n343_), .Y(men_men_n346_));
  NA2        u0318(.A(men_men_n229_), .B(men_men_n80_), .Y(men_men_n347_));
  NA3        u0319(.A(men_men_n347_), .B(men_men_n338_), .C(men_men_n212_), .Y(men_men_n348_));
  NA4        u0320(.A(men_men_n348_), .B(men_men_n346_), .C(men_men_n342_), .D(men_men_n339_), .Y(men_men_n349_));
  NA3        u0321(.A(h), .B(g), .C(f), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n350_), .B(men_men_n76_), .Y(men_men_n351_));
  NA2        u0323(.A(men_men_n334_), .B(men_men_n211_), .Y(men_men_n352_));
  NA2        u0324(.A(men_men_n165_), .B(e), .Y(men_men_n353_));
  NO2        u0325(.A(men_men_n353_), .B(men_men_n41_), .Y(men_men_n354_));
  AOI220     u0326(.A0(men_men_n354_), .A1(men_men_n306_), .B0(men_men_n352_), .B1(men_men_n351_), .Y(men_men_n355_));
  NOi32      u0327(.An(j), .Bn(g), .C(i), .Y(men_men_n356_));
  NA3        u0328(.A(men_men_n356_), .B(men_men_n285_), .C(men_men_n115_), .Y(men_men_n357_));
  AO210      u0329(.A0(men_men_n113_), .A1(men_men_n32_), .B0(men_men_n357_), .Y(men_men_n358_));
  NOi32      u0330(.An(e), .Bn(b), .C(a), .Y(men_men_n359_));
  AN2        u0331(.A(l), .B(j), .Y(men_men_n360_));
  NO2        u0332(.A(men_men_n313_), .B(men_men_n360_), .Y(men_men_n361_));
  NO3        u0333(.A(men_men_n315_), .B(men_men_n71_), .C(men_men_n214_), .Y(men_men_n362_));
  NA3        u0334(.A(men_men_n208_), .B(men_men_n206_), .C(men_men_n35_), .Y(men_men_n363_));
  AOI220     u0335(.A0(men_men_n363_), .A1(men_men_n359_), .B0(men_men_n362_), .B1(men_men_n361_), .Y(men_men_n364_));
  NO2        u0336(.A(men_men_n322_), .B(n), .Y(men_men_n365_));
  NA2        u0337(.A(men_men_n207_), .B(k), .Y(men_men_n366_));
  NA3        u0338(.A(m), .B(men_men_n114_), .C(men_men_n213_), .Y(men_men_n367_));
  NA4        u0339(.A(men_men_n202_), .B(men_men_n88_), .C(g), .D(men_men_n213_), .Y(men_men_n368_));
  OAI210     u0340(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n368_), .Y(men_men_n369_));
  NAi41      u0341(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n370_));
  NA2        u0342(.A(men_men_n51_), .B(men_men_n115_), .Y(men_men_n371_));
  NO2        u0343(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  AOI220     u0344(.A0(men_men_n372_), .A1(b), .B0(men_men_n369_), .B1(men_men_n365_), .Y(men_men_n373_));
  NA4        u0345(.A(men_men_n373_), .B(men_men_n364_), .C(men_men_n358_), .D(men_men_n355_), .Y(men_men_n374_));
  NO4        u0346(.A(men_men_n374_), .B(men_men_n349_), .C(men_men_n332_), .D(men_men_n325_), .Y(men_men_n375_));
  NA4        u0347(.A(men_men_n375_), .B(men_men_n312_), .C(men_men_n264_), .D(men_men_n198_), .Y(men10));
  NA3        u0348(.A(m), .B(k), .C(i), .Y(men_men_n377_));
  NO3        u0349(.A(men_men_n377_), .B(j), .C(men_men_n214_), .Y(men_men_n378_));
  NOi21      u0350(.An(e), .B(f), .Y(men_men_n379_));
  NO4        u0351(.A(men_men_n153_), .B(men_men_n379_), .C(n), .D(men_men_n112_), .Y(men_men_n380_));
  NAi31      u0352(.An(b), .B(f), .C(c), .Y(men_men_n381_));
  INV        u0353(.A(men_men_n381_), .Y(men_men_n382_));
  NOi32      u0354(.An(k), .Bn(h), .C(j), .Y(men_men_n383_));
  NA2        u0355(.A(men_men_n383_), .B(men_men_n221_), .Y(men_men_n384_));
  NA2        u0356(.A(men_men_n163_), .B(men_men_n384_), .Y(men_men_n385_));
  AOI220     u0357(.A0(men_men_n385_), .A1(men_men_n382_), .B0(men_men_n380_), .B1(men_men_n378_), .Y(men_men_n386_));
  OR2        u0358(.A(m), .B(k), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n175_), .B(men_men_n387_), .Y(men_men_n388_));
  NA4        u0360(.A(n), .B(f), .C(c), .D(men_men_n117_), .Y(men_men_n389_));
  NOi21      u0361(.An(men_men_n388_), .B(men_men_n389_), .Y(men_men_n390_));
  NOi32      u0362(.An(d), .Bn(a), .C(c), .Y(men_men_n391_));
  NA2        u0363(.A(men_men_n391_), .B(men_men_n183_), .Y(men_men_n392_));
  NAi21      u0364(.An(i), .B(g), .Y(men_men_n393_));
  NAi31      u0365(.An(k), .B(m), .C(j), .Y(men_men_n394_));
  NO3        u0366(.A(men_men_n394_), .B(men_men_n393_), .C(n), .Y(men_men_n395_));
  NOi21      u0367(.An(men_men_n395_), .B(men_men_n392_), .Y(men_men_n396_));
  NO2        u0368(.A(men_men_n396_), .B(men_men_n390_), .Y(men_men_n397_));
  NO2        u0369(.A(men_men_n389_), .B(men_men_n294_), .Y(men_men_n398_));
  AOI220     u0370(.A0(f), .A1(men_men_n304_), .B0(men_men_n398_), .B1(men_men_n215_), .Y(men_men_n399_));
  NA3        u0371(.A(men_men_n399_), .B(men_men_n397_), .C(men_men_n386_), .Y(men_men_n400_));
  NO2        u0372(.A(men_men_n59_), .B(men_men_n117_), .Y(men_men_n401_));
  NA2        u0373(.A(men_men_n247_), .B(men_men_n401_), .Y(men_men_n402_));
  INV        u0374(.A(e), .Y(men_men_n403_));
  NA2        u0375(.A(men_men_n46_), .B(e), .Y(men_men_n404_));
  OAI220     u0376(.A0(men_men_n404_), .A1(men_men_n199_), .B0(men_men_n203_), .B1(men_men_n403_), .Y(men_men_n405_));
  AN2        u0377(.A(g), .B(e), .Y(men_men_n406_));
  NA3        u0378(.A(men_men_n406_), .B(men_men_n202_), .C(i), .Y(men_men_n407_));
  OAI210     u0379(.A0(men_men_n90_), .A1(men_men_n403_), .B0(men_men_n407_), .Y(men_men_n408_));
  NO2        u0380(.A(men_men_n102_), .B(men_men_n403_), .Y(men_men_n409_));
  NO3        u0381(.A(men_men_n409_), .B(men_men_n408_), .C(men_men_n405_), .Y(men_men_n410_));
  NOi32      u0382(.An(h), .Bn(e), .C(g), .Y(men_men_n411_));
  NA3        u0383(.A(men_men_n411_), .B(men_men_n287_), .C(m), .Y(men_men_n412_));
  NOi21      u0384(.An(g), .B(h), .Y(men_men_n413_));
  AN3        u0385(.A(m), .B(l), .C(i), .Y(men_men_n414_));
  NA3        u0386(.A(men_men_n414_), .B(men_men_n413_), .C(e), .Y(men_men_n415_));
  AN3        u0387(.A(h), .B(g), .C(e), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n416_), .B(men_men_n99_), .Y(men_men_n417_));
  AN3        u0389(.A(men_men_n417_), .B(men_men_n415_), .C(men_men_n412_), .Y(men_men_n418_));
  AOI210     u0390(.A0(men_men_n418_), .A1(men_men_n410_), .B0(men_men_n402_), .Y(men_men_n419_));
  NA3        u0391(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n420_));
  NO2        u0392(.A(men_men_n420_), .B(men_men_n402_), .Y(men_men_n421_));
  NA3        u0393(.A(men_men_n391_), .B(men_men_n183_), .C(men_men_n85_), .Y(men_men_n422_));
  NAi31      u0394(.An(b), .B(c), .C(a), .Y(men_men_n423_));
  NO2        u0395(.A(men_men_n423_), .B(n), .Y(men_men_n424_));
  OAI210     u0396(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n425_));
  NO3        u0397(.A(men_men_n421_), .B(men_men_n419_), .C(men_men_n400_), .Y(men_men_n426_));
  NA2        u0398(.A(i), .B(g), .Y(men_men_n427_));
  NO3        u0399(.A(men_men_n273_), .B(men_men_n427_), .C(c), .Y(men_men_n428_));
  NOi21      u0400(.An(d), .B(c), .Y(men_men_n429_));
  NA2        u0401(.A(men_men_n429_), .B(a), .Y(men_men_n430_));
  NA3        u0402(.A(i), .B(g), .C(f), .Y(men_men_n431_));
  OR2        u0403(.A(men_men_n431_), .B(men_men_n70_), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n414_), .B(men_men_n413_), .C(men_men_n183_), .Y(men_men_n433_));
  AOI210     u0405(.A0(men_men_n433_), .A1(men_men_n432_), .B0(men_men_n430_), .Y(men_men_n434_));
  AOI210     u0406(.A0(men_men_n428_), .A1(men_men_n286_), .B0(men_men_n434_), .Y(men_men_n435_));
  OR2        u0407(.A(n), .B(m), .Y(men_men_n436_));
  NO2        u0408(.A(men_men_n436_), .B(men_men_n154_), .Y(men_men_n437_));
  OAI210     u0409(.A0(men_men_n437_), .A1(men_men_n177_), .B0(f), .Y(men_men_n438_));
  INV        u0410(.A(men_men_n371_), .Y(men_men_n439_));
  NA3        u0411(.A(men_men_n439_), .B(men_men_n359_), .C(d), .Y(men_men_n440_));
  NO2        u0412(.A(men_men_n423_), .B(men_men_n49_), .Y(men_men_n441_));
  NO3        u0413(.A(men_men_n65_), .B(men_men_n114_), .C(e), .Y(men_men_n442_));
  NAi21      u0414(.An(k), .B(j), .Y(men_men_n443_));
  NA2        u0415(.A(men_men_n250_), .B(men_men_n443_), .Y(men_men_n444_));
  NA3        u0416(.A(men_men_n444_), .B(men_men_n442_), .C(men_men_n441_), .Y(men_men_n445_));
  NAi21      u0417(.An(e), .B(d), .Y(men_men_n446_));
  NA3        u0418(.A(men_men_n445_), .B(men_men_n440_), .C(men_men_n438_), .Y(men_men_n447_));
  NOi31      u0419(.An(n), .B(m), .C(k), .Y(men_men_n448_));
  AOI220     u0420(.A0(men_men_n448_), .A1(h), .B0(men_men_n221_), .B1(men_men_n50_), .Y(men_men_n449_));
  NAi31      u0421(.An(g), .B(f), .C(c), .Y(men_men_n450_));
  OR3        u0422(.A(men_men_n450_), .B(men_men_n449_), .C(e), .Y(men_men_n451_));
  NA2        u0423(.A(men_men_n451_), .B(men_men_n305_), .Y(men_men_n452_));
  NOi41      u0424(.An(men_men_n435_), .B(men_men_n452_), .C(men_men_n447_), .D(men_men_n262_), .Y(men_men_n453_));
  NOi32      u0425(.An(c), .Bn(a), .C(b), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n115_), .Y(men_men_n455_));
  INV        u0427(.A(men_men_n271_), .Y(men_men_n456_));
  AN2        u0428(.A(e), .B(d), .Y(men_men_n457_));
  NO2        u0429(.A(men_men_n133_), .B(men_men_n41_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n65_), .B(e), .Y(men_men_n459_));
  NOi31      u0431(.An(j), .B(k), .C(i), .Y(men_men_n460_));
  NOi21      u0432(.An(men_men_n168_), .B(men_men_n460_), .Y(men_men_n461_));
  NA4        u0433(.A(men_men_n316_), .B(men_men_n461_), .C(men_men_n256_), .D(men_men_n120_), .Y(men_men_n462_));
  AOI210     u0434(.A0(men_men_n462_), .A1(men_men_n459_), .B0(men_men_n458_), .Y(men_men_n463_));
  AOI210     u0435(.A0(men_men_n463_), .A1(men_men_n271_), .B0(men_men_n455_), .Y(men_men_n464_));
  NO2        u0436(.A(men_men_n209_), .B(men_men_n204_), .Y(men_men_n465_));
  NOi21      u0437(.An(a), .B(b), .Y(men_men_n466_));
  NA3        u0438(.A(e), .B(d), .C(c), .Y(men_men_n467_));
  NAi21      u0439(.An(men_men_n467_), .B(men_men_n466_), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n422_), .B(men_men_n203_), .Y(men_men_n469_));
  NOi21      u0441(.An(men_men_n468_), .B(men_men_n469_), .Y(men_men_n470_));
  AOI210     u0442(.A0(men_men_n265_), .A1(men_men_n465_), .B0(men_men_n470_), .Y(men_men_n471_));
  OR2        u0443(.A(k), .B(j), .Y(men_men_n472_));
  NA2        u0444(.A(l), .B(k), .Y(men_men_n473_));
  NA3        u0445(.A(men_men_n473_), .B(men_men_n472_), .C(men_men_n221_), .Y(men_men_n474_));
  AOI210     u0446(.A0(men_men_n229_), .A1(men_men_n333_), .B0(men_men_n85_), .Y(men_men_n475_));
  NOi21      u0447(.An(men_men_n474_), .B(men_men_n475_), .Y(men_men_n476_));
  OR3        u0448(.A(men_men_n476_), .B(men_men_n146_), .C(men_men_n137_), .Y(men_men_n477_));
  NA3        u0449(.A(men_men_n276_), .B(men_men_n130_), .C(men_men_n128_), .Y(men_men_n478_));
  NA2        u0450(.A(men_men_n391_), .B(men_men_n115_), .Y(men_men_n479_));
  NO4        u0451(.A(men_men_n479_), .B(men_men_n96_), .C(men_men_n114_), .D(e), .Y(men_men_n480_));
  NO3        u0452(.A(men_men_n422_), .B(men_men_n93_), .C(men_men_n133_), .Y(men_men_n481_));
  NO4        u0453(.A(men_men_n481_), .B(men_men_n480_), .C(men_men_n478_), .D(men_men_n317_), .Y(men_men_n482_));
  NA2        u0454(.A(men_men_n482_), .B(men_men_n477_), .Y(men_men_n483_));
  NO3        u0455(.A(men_men_n483_), .B(men_men_n471_), .C(men_men_n464_), .Y(men_men_n484_));
  NA2        u0456(.A(men_men_n69_), .B(men_men_n66_), .Y(men_men_n485_));
  INV        u0457(.A(men_men_n189_), .Y(men_men_n486_));
  NAi31      u0458(.An(j), .B(l), .C(i), .Y(men_men_n487_));
  OAI210     u0459(.A0(men_men_n487_), .A1(men_men_n134_), .B0(men_men_n105_), .Y(men_men_n488_));
  NA3        u0460(.A(men_men_n488_), .B(men_men_n486_), .C(d), .Y(men_men_n489_));
  NO3        u0461(.A(men_men_n392_), .B(men_men_n341_), .C(men_men_n200_), .Y(men_men_n490_));
  NO2        u0462(.A(men_men_n392_), .B(men_men_n371_), .Y(men_men_n491_));
  NO3        u0463(.A(men_men_n491_), .B(men_men_n490_), .C(men_men_n185_), .Y(men_men_n492_));
  NA4        u0464(.A(men_men_n492_), .B(men_men_n489_), .C(men_men_n485_), .D(men_men_n239_), .Y(men_men_n493_));
  OAI210     u0465(.A0(men_men_n129_), .A1(men_men_n127_), .B0(n), .Y(men_men_n494_));
  NO2        u0466(.A(men_men_n494_), .B(men_men_n133_), .Y(men_men_n495_));
  OR2        u0467(.A(men_men_n295_), .B(men_men_n241_), .Y(men_men_n496_));
  OA210      u0468(.A0(men_men_n496_), .A1(men_men_n495_), .B0(men_men_n193_), .Y(men_men_n497_));
  XO2        u0469(.A(i), .B(h), .Y(men_men_n498_));
  NA3        u0470(.A(men_men_n498_), .B(men_men_n162_), .C(n), .Y(men_men_n499_));
  NAi41      u0471(.An(men_men_n295_), .B(men_men_n499_), .C(men_men_n449_), .D(men_men_n384_), .Y(men_men_n500_));
  NOi32      u0472(.An(men_men_n500_), .Bn(men_men_n459_), .C(men_men_n267_), .Y(men_men_n501_));
  BUFFER     u0473(.A(men_men_n83_), .Y(men_men_n502_));
  NA3        u0474(.A(men_men_n380_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n503_));
  NA2        u0475(.A(men_men_n226_), .B(men_men_n110_), .Y(men_men_n504_));
  NA2        u0476(.A(men_men_n504_), .B(men_men_n182_), .Y(men_men_n505_));
  AOI210     u0477(.A0(men_men_n357_), .A1(men_men_n35_), .B0(men_men_n468_), .Y(men_men_n506_));
  NOi31      u0478(.An(men_men_n503_), .B(men_men_n506_), .C(men_men_n505_), .Y(men_men_n507_));
  AO220      u0479(.A0(men_men_n283_), .A1(men_men_n259_), .B0(men_men_n169_), .B1(men_men_n66_), .Y(men_men_n508_));
  NA3        u0480(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n509_));
  NO2        u0481(.A(men_men_n509_), .B(men_men_n430_), .Y(men_men_n510_));
  NO2        u0482(.A(men_men_n510_), .B(men_men_n291_), .Y(men_men_n511_));
  NAi41      u0483(.An(men_men_n508_), .B(men_men_n511_), .C(men_men_n507_), .D(men_men_n502_), .Y(men_men_n512_));
  NO4        u0484(.A(men_men_n512_), .B(men_men_n501_), .C(men_men_n497_), .D(men_men_n493_), .Y(men_men_n513_));
  NA4        u0485(.A(men_men_n513_), .B(men_men_n484_), .C(men_men_n453_), .D(men_men_n426_), .Y(men11));
  NO2        u0486(.A(men_men_n72_), .B(f), .Y(men_men_n515_));
  NA2        u0487(.A(j), .B(g), .Y(men_men_n516_));
  NAi31      u0488(.An(i), .B(m), .C(l), .Y(men_men_n517_));
  NA3        u0489(.A(m), .B(k), .C(j), .Y(men_men_n518_));
  OAI220     u0490(.A0(men_men_n518_), .A1(men_men_n133_), .B0(men_men_n517_), .B1(men_men_n516_), .Y(men_men_n519_));
  NA2        u0491(.A(men_men_n519_), .B(men_men_n515_), .Y(men_men_n520_));
  NOi32      u0492(.An(e), .Bn(b), .C(f), .Y(men_men_n521_));
  NA2        u0493(.A(men_men_n255_), .B(men_men_n115_), .Y(men_men_n522_));
  NA2        u0494(.A(men_men_n46_), .B(j), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n523_), .B(men_men_n297_), .Y(men_men_n524_));
  NAi31      u0496(.An(d), .B(e), .C(a), .Y(men_men_n525_));
  NO2        u0497(.A(men_men_n525_), .B(n), .Y(men_men_n526_));
  AOI220     u0498(.A0(men_men_n526_), .A1(men_men_n103_), .B0(men_men_n524_), .B1(men_men_n521_), .Y(men_men_n527_));
  NAi41      u0499(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n528_));
  AN2        u0500(.A(men_men_n528_), .B(men_men_n370_), .Y(men_men_n529_));
  AOI210     u0501(.A0(men_men_n529_), .A1(men_men_n392_), .B0(men_men_n268_), .Y(men_men_n530_));
  NA2        u0502(.A(j), .B(i), .Y(men_men_n531_));
  NAi31      u0503(.An(n), .B(m), .C(k), .Y(men_men_n532_));
  NO3        u0504(.A(men_men_n532_), .B(men_men_n531_), .C(men_men_n114_), .Y(men_men_n533_));
  NO4        u0505(.A(n), .B(d), .C(men_men_n117_), .D(a), .Y(men_men_n534_));
  NO2        u0506(.A(c), .B(men_men_n152_), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n535_), .B(men_men_n534_), .Y(men_men_n536_));
  NOi32      u0508(.An(g), .Bn(f), .C(i), .Y(men_men_n537_));
  AOI220     u0509(.A0(men_men_n537_), .A1(men_men_n101_), .B0(men_men_n519_), .B1(f), .Y(men_men_n538_));
  NO2        u0510(.A(men_men_n271_), .B(men_men_n49_), .Y(men_men_n539_));
  NO2        u0511(.A(men_men_n538_), .B(men_men_n536_), .Y(men_men_n540_));
  AOI210     u0512(.A0(men_men_n533_), .A1(men_men_n530_), .B0(men_men_n540_), .Y(men_men_n541_));
  NA2        u0513(.A(men_men_n142_), .B(men_men_n34_), .Y(men_men_n542_));
  OAI220     u0514(.A0(men_men_n542_), .A1(m), .B0(men_men_n523_), .B1(men_men_n229_), .Y(men_men_n543_));
  NOi41      u0515(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n544_));
  NAi32      u0516(.An(e), .Bn(b), .C(c), .Y(men_men_n545_));
  AN2        u0517(.A(men_men_n334_), .B(men_men_n315_), .Y(men_men_n546_));
  NA2        u0518(.A(men_men_n546_), .B(men_men_n545_), .Y(men_men_n547_));
  OA210      u0519(.A0(men_men_n547_), .A1(men_men_n544_), .B0(men_men_n543_), .Y(men_men_n548_));
  OAI220     u0520(.A0(men_men_n394_), .A1(men_men_n393_), .B0(men_men_n517_), .B1(men_men_n516_), .Y(men_men_n549_));
  NAi31      u0521(.An(d), .B(c), .C(a), .Y(men_men_n550_));
  NO2        u0522(.A(men_men_n550_), .B(n), .Y(men_men_n551_));
  NA3        u0523(.A(men_men_n551_), .B(men_men_n549_), .C(e), .Y(men_men_n552_));
  NO3        u0524(.A(men_men_n61_), .B(men_men_n49_), .C(men_men_n214_), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n227_), .B(men_men_n112_), .Y(men_men_n554_));
  OAI210     u0526(.A0(men_men_n553_), .A1(men_men_n395_), .B0(men_men_n554_), .Y(men_men_n555_));
  NA2        u0527(.A(men_men_n555_), .B(men_men_n552_), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n273_), .B(n), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n424_), .B(men_men_n557_), .Y(men_men_n558_));
  NA2        u0530(.A(men_men_n549_), .B(f), .Y(men_men_n559_));
  NAi32      u0531(.An(d), .Bn(a), .C(b), .Y(men_men_n560_));
  NO2        u0532(.A(men_men_n560_), .B(men_men_n49_), .Y(men_men_n561_));
  NA2        u0533(.A(h), .B(f), .Y(men_men_n562_));
  NO2        u0534(.A(men_men_n562_), .B(men_men_n96_), .Y(men_men_n563_));
  NO3        u0535(.A(men_men_n178_), .B(men_men_n175_), .C(g), .Y(men_men_n564_));
  AOI220     u0536(.A0(men_men_n564_), .A1(men_men_n58_), .B0(men_men_n563_), .B1(men_men_n561_), .Y(men_men_n565_));
  OAI210     u0537(.A0(men_men_n559_), .A1(men_men_n558_), .B0(men_men_n565_), .Y(men_men_n566_));
  AN3        u0538(.A(j), .B(h), .C(g), .Y(men_men_n567_));
  NO2        u0539(.A(men_men_n149_), .B(c), .Y(men_men_n568_));
  NA3        u0540(.A(men_men_n568_), .B(men_men_n567_), .C(men_men_n448_), .Y(men_men_n569_));
  NA3        u0541(.A(f), .B(d), .C(b), .Y(men_men_n570_));
  NO4        u0542(.A(men_men_n570_), .B(men_men_n178_), .C(men_men_n175_), .D(g), .Y(men_men_n571_));
  NAi21      u0543(.An(men_men_n571_), .B(men_men_n569_), .Y(men_men_n572_));
  NO4        u0544(.A(men_men_n572_), .B(men_men_n566_), .C(men_men_n556_), .D(men_men_n548_), .Y(men_men_n573_));
  AN4        u0545(.A(men_men_n573_), .B(men_men_n541_), .C(men_men_n527_), .D(men_men_n520_), .Y(men_men_n574_));
  INV        u0546(.A(k), .Y(men_men_n575_));
  NA3        u0547(.A(l), .B(men_men_n575_), .C(i), .Y(men_men_n576_));
  INV        u0548(.A(men_men_n576_), .Y(men_men_n577_));
  NA4        u0549(.A(men_men_n391_), .B(men_men_n413_), .C(men_men_n183_), .D(men_men_n115_), .Y(men_men_n578_));
  NAi32      u0550(.An(h), .Bn(f), .C(g), .Y(men_men_n579_));
  NAi41      u0551(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n580_));
  OAI210     u0552(.A0(men_men_n525_), .A1(n), .B0(men_men_n580_), .Y(men_men_n581_));
  NA2        u0553(.A(men_men_n581_), .B(m), .Y(men_men_n582_));
  NAi31      u0554(.An(h), .B(g), .C(f), .Y(men_men_n583_));
  OR3        u0555(.A(men_men_n583_), .B(men_men_n273_), .C(men_men_n49_), .Y(men_men_n584_));
  NA4        u0556(.A(men_men_n413_), .B(men_men_n122_), .C(men_men_n115_), .D(e), .Y(men_men_n585_));
  AN2        u0557(.A(men_men_n585_), .B(men_men_n584_), .Y(men_men_n586_));
  OA210      u0558(.A0(men_men_n582_), .A1(men_men_n579_), .B0(men_men_n586_), .Y(men_men_n587_));
  NO3        u0559(.A(men_men_n579_), .B(men_men_n72_), .C(men_men_n74_), .Y(men_men_n588_));
  NO4        u0560(.A(men_men_n583_), .B(c), .C(men_men_n152_), .D(men_men_n74_), .Y(men_men_n589_));
  OR2        u0561(.A(men_men_n589_), .B(men_men_n588_), .Y(men_men_n590_));
  NAi31      u0562(.An(men_men_n590_), .B(men_men_n587_), .C(men_men_n578_), .Y(men_men_n591_));
  NAi31      u0563(.An(f), .B(h), .C(g), .Y(men_men_n592_));
  NO4        u0564(.A(men_men_n307_), .B(men_men_n592_), .C(men_men_n72_), .D(men_men_n74_), .Y(men_men_n593_));
  NOi32      u0565(.An(b), .Bn(a), .C(c), .Y(men_men_n594_));
  NOi41      u0566(.An(men_men_n594_), .B(men_men_n350_), .C(men_men_n68_), .D(men_men_n118_), .Y(men_men_n595_));
  OR2        u0567(.A(men_men_n595_), .B(men_men_n593_), .Y(men_men_n596_));
  NOi32      u0568(.An(d), .Bn(a), .C(e), .Y(men_men_n597_));
  NA2        u0569(.A(men_men_n597_), .B(men_men_n115_), .Y(men_men_n598_));
  NO2        u0570(.A(n), .B(c), .Y(men_men_n599_));
  NA3        u0571(.A(men_men_n599_), .B(men_men_n29_), .C(m), .Y(men_men_n600_));
  NAi32      u0572(.An(n), .Bn(f), .C(m), .Y(men_men_n601_));
  NA3        u0573(.A(men_men_n601_), .B(men_men_n600_), .C(men_men_n598_), .Y(men_men_n602_));
  NOi32      u0574(.An(e), .Bn(a), .C(d), .Y(men_men_n603_));
  AOI210     u0575(.A0(men_men_n29_), .A1(d), .B0(men_men_n603_), .Y(men_men_n604_));
  INV        u0576(.A(men_men_n542_), .Y(men_men_n605_));
  AOI210     u0577(.A0(men_men_n605_), .A1(men_men_n602_), .B0(men_men_n596_), .Y(men_men_n606_));
  OAI210     u0578(.A0(men_men_n246_), .A1(men_men_n88_), .B0(men_men_n606_), .Y(men_men_n607_));
  AOI210     u0579(.A0(men_men_n591_), .A1(men_men_n577_), .B0(men_men_n607_), .Y(men_men_n608_));
  NO3        u0580(.A(men_men_n313_), .B(men_men_n60_), .C(n), .Y(men_men_n609_));
  NA2        u0581(.A(men_men_n75_), .B(men_men_n115_), .Y(men_men_n610_));
  NO2        u0582(.A(men_men_n610_), .B(men_men_n45_), .Y(men_men_n611_));
  AOI220     u0583(.A0(men_men_n611_), .A1(men_men_n530_), .B0(c), .B1(men_men_n609_), .Y(men_men_n612_));
  NO2        u0584(.A(men_men_n612_), .B(men_men_n88_), .Y(men_men_n613_));
  NA3        u0585(.A(men_men_n544_), .B(men_men_n336_), .C(men_men_n46_), .Y(men_men_n614_));
  NOi32      u0586(.An(e), .Bn(c), .C(f), .Y(men_men_n615_));
  NOi21      u0587(.An(f), .B(g), .Y(men_men_n616_));
  NO2        u0588(.A(men_men_n616_), .B(men_men_n211_), .Y(men_men_n617_));
  AOI220     u0589(.A0(men_men_n617_), .A1(men_men_n388_), .B0(men_men_n615_), .B1(men_men_n177_), .Y(men_men_n618_));
  NA3        u0590(.A(men_men_n618_), .B(men_men_n614_), .C(men_men_n180_), .Y(men_men_n619_));
  AOI210     u0591(.A0(men_men_n529_), .A1(men_men_n392_), .B0(men_men_n296_), .Y(men_men_n620_));
  NA2        u0592(.A(men_men_n620_), .B(men_men_n260_), .Y(men_men_n621_));
  NOi21      u0593(.An(j), .B(l), .Y(men_men_n622_));
  NAi21      u0594(.An(k), .B(h), .Y(men_men_n623_));
  NO2        u0595(.A(men_men_n623_), .B(men_men_n258_), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n624_), .B(men_men_n622_), .Y(men_men_n625_));
  OR2        u0597(.A(men_men_n625_), .B(men_men_n582_), .Y(men_men_n626_));
  NOi31      u0598(.An(m), .B(n), .C(k), .Y(men_men_n627_));
  NA2        u0599(.A(men_men_n622_), .B(men_men_n627_), .Y(men_men_n628_));
  AOI210     u0600(.A0(men_men_n392_), .A1(men_men_n370_), .B0(men_men_n296_), .Y(men_men_n629_));
  NAi21      u0601(.An(men_men_n628_), .B(men_men_n629_), .Y(men_men_n630_));
  NO2        u0602(.A(men_men_n273_), .B(men_men_n49_), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n307_), .B(men_men_n592_), .Y(men_men_n632_));
  NO2        u0604(.A(men_men_n525_), .B(men_men_n49_), .Y(men_men_n633_));
  AOI220     u0605(.A0(men_men_n633_), .A1(men_men_n632_), .B0(men_men_n631_), .B1(men_men_n563_), .Y(men_men_n634_));
  NA4        u0606(.A(men_men_n634_), .B(men_men_n630_), .C(men_men_n626_), .D(men_men_n621_), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n110_), .B(men_men_n36_), .Y(men_men_n636_));
  NO2        u0608(.A(k), .B(men_men_n214_), .Y(men_men_n637_));
  NO2        u0609(.A(men_men_n521_), .B(men_men_n359_), .Y(men_men_n638_));
  NO2        u0610(.A(men_men_n638_), .B(n), .Y(men_men_n639_));
  NAi31      u0611(.An(men_men_n636_), .B(men_men_n639_), .C(men_men_n637_), .Y(men_men_n640_));
  NO2        u0612(.A(men_men_n523_), .B(men_men_n178_), .Y(men_men_n641_));
  NA3        u0613(.A(men_men_n545_), .B(men_men_n267_), .C(men_men_n147_), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n498_), .B(men_men_n162_), .Y(men_men_n643_));
  NO3        u0615(.A(men_men_n389_), .B(men_men_n643_), .C(men_men_n88_), .Y(men_men_n644_));
  AOI210     u0616(.A0(men_men_n642_), .A1(men_men_n641_), .B0(men_men_n644_), .Y(men_men_n645_));
  AN3        u0617(.A(f), .B(d), .C(b), .Y(men_men_n646_));
  NO2        u0618(.A(men_men_n646_), .B(men_men_n132_), .Y(men_men_n647_));
  NA3        u0619(.A(men_men_n498_), .B(men_men_n162_), .C(men_men_n214_), .Y(men_men_n648_));
  AOI210     u0620(.A0(men_men_n647_), .A1(men_men_n228_), .B0(men_men_n648_), .Y(men_men_n649_));
  NAi31      u0621(.An(m), .B(n), .C(k), .Y(men_men_n650_));
  OR2        u0622(.A(men_men_n137_), .B(men_men_n60_), .Y(men_men_n651_));
  OAI210     u0623(.A0(men_men_n651_), .A1(men_men_n650_), .B0(men_men_n248_), .Y(men_men_n652_));
  OAI210     u0624(.A0(men_men_n652_), .A1(men_men_n649_), .B0(j), .Y(men_men_n653_));
  NA3        u0625(.A(men_men_n653_), .B(men_men_n645_), .C(men_men_n640_), .Y(men_men_n654_));
  NO4        u0626(.A(men_men_n654_), .B(men_men_n635_), .C(men_men_n619_), .D(men_men_n613_), .Y(men_men_n655_));
  NA2        u0627(.A(men_men_n380_), .B(men_men_n165_), .Y(men_men_n656_));
  NAi31      u0628(.An(g), .B(h), .C(f), .Y(men_men_n657_));
  OR3        u0629(.A(men_men_n657_), .B(men_men_n273_), .C(n), .Y(men_men_n658_));
  OA210      u0630(.A0(men_men_n525_), .A1(n), .B0(men_men_n580_), .Y(men_men_n659_));
  NA3        u0631(.A(men_men_n411_), .B(men_men_n122_), .C(men_men_n85_), .Y(men_men_n660_));
  OAI210     u0632(.A0(men_men_n659_), .A1(men_men_n92_), .B0(men_men_n660_), .Y(men_men_n661_));
  NOi21      u0633(.An(men_men_n658_), .B(men_men_n661_), .Y(men_men_n662_));
  AOI210     u0634(.A0(men_men_n662_), .A1(men_men_n656_), .B0(men_men_n518_), .Y(men_men_n663_));
  NO3        u0635(.A(g), .B(men_men_n213_), .C(men_men_n56_), .Y(men_men_n664_));
  NAi21      u0636(.An(h), .B(j), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n504_), .B(men_men_n88_), .Y(men_men_n666_));
  OAI210     u0638(.A0(men_men_n666_), .A1(men_men_n388_), .B0(men_men_n664_), .Y(men_men_n667_));
  NA2        u0639(.A(men_men_n594_), .B(men_men_n338_), .Y(men_men_n668_));
  OA220      u0640(.A0(men_men_n628_), .A1(men_men_n668_), .B0(men_men_n625_), .B1(men_men_n72_), .Y(men_men_n669_));
  NA3        u0641(.A(men_men_n515_), .B(men_men_n101_), .C(men_men_n100_), .Y(men_men_n670_));
  NA2        u0642(.A(h), .B(men_men_n37_), .Y(men_men_n671_));
  NA2        u0643(.A(men_men_n101_), .B(men_men_n46_), .Y(men_men_n672_));
  OAI220     u0644(.A0(men_men_n672_), .A1(men_men_n327_), .B0(men_men_n671_), .B1(men_men_n455_), .Y(men_men_n673_));
  AOI210     u0645(.A0(men_men_n560_), .A1(men_men_n423_), .B0(men_men_n49_), .Y(men_men_n674_));
  OAI220     u0646(.A0(men_men_n583_), .A1(men_men_n576_), .B0(men_men_n320_), .B1(men_men_n516_), .Y(men_men_n675_));
  AOI210     u0647(.A0(men_men_n675_), .A1(men_men_n674_), .B0(men_men_n673_), .Y(men_men_n676_));
  NA4        u0648(.A(men_men_n676_), .B(men_men_n670_), .C(men_men_n669_), .D(men_men_n667_), .Y(men_men_n677_));
  NO2        u0649(.A(men_men_n250_), .B(f), .Y(men_men_n678_));
  NO2        u0650(.A(men_men_n616_), .B(men_men_n60_), .Y(men_men_n679_));
  NO3        u0651(.A(men_men_n679_), .B(men_men_n678_), .C(men_men_n34_), .Y(men_men_n680_));
  NA2        u0652(.A(men_men_n323_), .B(men_men_n142_), .Y(men_men_n681_));
  NA2        u0653(.A(men_men_n134_), .B(men_men_n49_), .Y(men_men_n682_));
  AOI220     u0654(.A0(men_men_n682_), .A1(men_men_n521_), .B0(men_men_n359_), .B1(men_men_n115_), .Y(men_men_n683_));
  OA220      u0655(.A0(men_men_n683_), .A1(men_men_n542_), .B0(men_men_n357_), .B1(men_men_n113_), .Y(men_men_n684_));
  OAI210     u0656(.A0(men_men_n681_), .A1(men_men_n680_), .B0(men_men_n684_), .Y(men_men_n685_));
  NA2        u0657(.A(men_men_n454_), .B(men_men_n85_), .Y(men_men_n686_));
  NO4        u0658(.A(men_men_n518_), .B(men_men_n686_), .C(men_men_n133_), .D(men_men_n213_), .Y(men_men_n687_));
  INV        u0659(.A(men_men_n687_), .Y(men_men_n688_));
  NA3        u0660(.A(men_men_n688_), .B(men_men_n503_), .C(men_men_n397_), .Y(men_men_n689_));
  NO4        u0661(.A(men_men_n689_), .B(men_men_n685_), .C(men_men_n677_), .D(men_men_n663_), .Y(men_men_n690_));
  NA4        u0662(.A(men_men_n690_), .B(men_men_n655_), .C(men_men_n608_), .D(men_men_n574_), .Y(men08));
  NO2        u0663(.A(k), .B(h), .Y(men_men_n692_));
  AO210      u0664(.A0(men_men_n250_), .A1(men_men_n443_), .B0(men_men_n692_), .Y(men_men_n693_));
  NO2        u0665(.A(men_men_n693_), .B(men_men_n294_), .Y(men_men_n694_));
  AOI210     u0666(.A0(men_men_n1513_), .A1(men_men_n694_), .B0(men_men_n481_), .Y(men_men_n695_));
  NA2        u0667(.A(men_men_n85_), .B(men_men_n112_), .Y(men_men_n696_));
  NO2        u0668(.A(men_men_n696_), .B(men_men_n57_), .Y(men_men_n697_));
  NO4        u0669(.A(men_men_n377_), .B(men_men_n114_), .C(j), .D(men_men_n214_), .Y(men_men_n698_));
  NA2        u0670(.A(men_men_n570_), .B(men_men_n228_), .Y(men_men_n699_));
  AOI220     u0671(.A0(men_men_n699_), .A1(men_men_n344_), .B0(men_men_n698_), .B1(men_men_n697_), .Y(men_men_n700_));
  AOI210     u0672(.A0(men_men_n570_), .A1(men_men_n158_), .B0(men_men_n85_), .Y(men_men_n701_));
  NA4        u0673(.A(men_men_n216_), .B(men_men_n142_), .C(men_men_n45_), .D(h), .Y(men_men_n702_));
  AN2        u0674(.A(l), .B(k), .Y(men_men_n703_));
  NA3        u0675(.A(men_men_n703_), .B(men_men_n110_), .C(men_men_n214_), .Y(men_men_n704_));
  OAI210     u0676(.A0(men_men_n702_), .A1(g), .B0(men_men_n704_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n705_), .B(men_men_n701_), .Y(men_men_n706_));
  NA4        u0678(.A(men_men_n706_), .B(men_men_n700_), .C(men_men_n695_), .D(men_men_n346_), .Y(men_men_n707_));
  AN2        u0679(.A(men_men_n526_), .B(men_men_n97_), .Y(men_men_n708_));
  NO4        u0680(.A(men_men_n175_), .B(men_men_n387_), .C(men_men_n114_), .D(g), .Y(men_men_n709_));
  AOI210     u0681(.A0(men_men_n709_), .A1(men_men_n699_), .B0(men_men_n510_), .Y(men_men_n710_));
  NO2        u0682(.A(men_men_n38_), .B(men_men_n213_), .Y(men_men_n711_));
  NA2        u0683(.A(men_men_n711_), .B(men_men_n557_), .Y(men_men_n712_));
  NAi31      u0684(.An(men_men_n708_), .B(men_men_n712_), .C(men_men_n710_), .Y(men_men_n713_));
  NO2        u0685(.A(men_men_n529_), .B(men_men_n35_), .Y(men_men_n714_));
  OAI210     u0686(.A0(men_men_n545_), .A1(men_men_n47_), .B0(men_men_n651_), .Y(men_men_n715_));
  NO2        u0687(.A(men_men_n473_), .B(men_men_n134_), .Y(men_men_n716_));
  AOI210     u0688(.A0(men_men_n716_), .A1(men_men_n715_), .B0(men_men_n714_), .Y(men_men_n717_));
  NO3        u0689(.A(men_men_n313_), .B(men_men_n133_), .C(men_men_n41_), .Y(men_men_n718_));
  NAi21      u0690(.An(men_men_n718_), .B(men_men_n704_), .Y(men_men_n719_));
  NA2        u0691(.A(men_men_n719_), .B(men_men_n77_), .Y(men_men_n720_));
  OAI210     u0692(.A0(men_men_n717_), .A1(men_men_n88_), .B0(men_men_n720_), .Y(men_men_n721_));
  NA2        u0693(.A(men_men_n359_), .B(men_men_n43_), .Y(men_men_n722_));
  NO2        u0694(.A(men_men_n1515_), .B(men_men_n322_), .Y(men_men_n723_));
  AOI210     u0695(.A0(men_men_n723_), .A1(men_men_n678_), .B0(men_men_n480_), .Y(men_men_n724_));
  NA3        u0696(.A(m), .B(l), .C(k), .Y(men_men_n725_));
  AOI210     u0697(.A0(men_men_n660_), .A1(men_men_n658_), .B0(men_men_n725_), .Y(men_men_n726_));
  NO2        u0698(.A(men_men_n528_), .B(men_men_n268_), .Y(men_men_n727_));
  NOi21      u0699(.An(men_men_n727_), .B(men_men_n522_), .Y(men_men_n728_));
  NA4        u0700(.A(men_men_n115_), .B(l), .C(k), .D(men_men_n88_), .Y(men_men_n729_));
  NA3        u0701(.A(men_men_n122_), .B(men_men_n406_), .C(i), .Y(men_men_n730_));
  NO2        u0702(.A(men_men_n730_), .B(men_men_n729_), .Y(men_men_n731_));
  NO3        u0703(.A(men_men_n731_), .B(men_men_n728_), .C(men_men_n726_), .Y(men_men_n732_));
  NA3        u0704(.A(men_men_n732_), .B(men_men_n724_), .C(men_men_n722_), .Y(men_men_n733_));
  NO4        u0705(.A(men_men_n733_), .B(men_men_n721_), .C(men_men_n713_), .D(men_men_n707_), .Y(men_men_n734_));
  NA2        u0706(.A(men_men_n617_), .B(men_men_n388_), .Y(men_men_n735_));
  NOi31      u0707(.An(g), .B(h), .C(f), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n633_), .B(men_men_n736_), .Y(men_men_n737_));
  AO210      u0709(.A0(men_men_n737_), .A1(men_men_n584_), .B0(men_men_n531_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n392_), .B(men_men_n516_), .C(h), .Y(men_men_n739_));
  NO2        u0711(.A(men_men_n739_), .B(men_men_n491_), .Y(men_men_n740_));
  NA4        u0712(.A(men_men_n740_), .B(men_men_n738_), .C(men_men_n735_), .D(men_men_n249_), .Y(men_men_n741_));
  INV        u0713(.A(men_men_n703_), .Y(men_men_n742_));
  NOi21      u0714(.An(h), .B(j), .Y(men_men_n743_));
  NA2        u0715(.A(men_men_n743_), .B(f), .Y(men_men_n744_));
  NO2        u0716(.A(men_men_n744_), .B(men_men_n243_), .Y(men_men_n745_));
  INV        u0717(.A(men_men_n745_), .Y(men_men_n746_));
  OAI220     u0718(.A0(men_men_n746_), .A1(men_men_n742_), .B0(men_men_n586_), .B1(men_men_n61_), .Y(men_men_n747_));
  AOI210     u0719(.A0(men_men_n741_), .A1(l), .B0(men_men_n747_), .Y(men_men_n748_));
  NO2        u0720(.A(j), .B(i), .Y(men_men_n749_));
  NA3        u0721(.A(men_men_n749_), .B(men_men_n81_), .C(l), .Y(men_men_n750_));
  NA2        u0722(.A(men_men_n749_), .B(men_men_n33_), .Y(men_men_n751_));
  NA2        u0723(.A(men_men_n416_), .B(men_men_n122_), .Y(men_men_n752_));
  OA220      u0724(.A0(men_men_n752_), .A1(men_men_n751_), .B0(men_men_n750_), .B1(men_men_n582_), .Y(men_men_n753_));
  NO3        u0725(.A(men_men_n153_), .B(men_men_n49_), .C(men_men_n112_), .Y(men_men_n754_));
  NO3        u0726(.A(c), .B(men_men_n152_), .C(men_men_n74_), .Y(men_men_n755_));
  NO3        u0727(.A(men_men_n473_), .B(men_men_n431_), .C(j), .Y(men_men_n756_));
  OAI210     u0728(.A0(men_men_n755_), .A1(men_men_n754_), .B0(men_men_n756_), .Y(men_men_n757_));
  OAI210     u0729(.A0(men_men_n737_), .A1(men_men_n61_), .B0(men_men_n757_), .Y(men_men_n758_));
  NA2        u0730(.A(k), .B(j), .Y(men_men_n759_));
  NO2        u0731(.A(men_men_n294_), .B(men_men_n40_), .Y(men_men_n760_));
  AOI210     u0732(.A0(men_men_n521_), .A1(n), .B0(men_men_n544_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n761_), .B(men_men_n546_), .Y(men_men_n762_));
  AN3        u0734(.A(men_men_n762_), .B(men_men_n760_), .C(men_men_n100_), .Y(men_men_n763_));
  NO3        u0735(.A(men_men_n175_), .B(men_men_n387_), .C(men_men_n114_), .Y(men_men_n764_));
  AOI210     u0736(.A0(men_men_n764_), .A1(men_men_n244_), .B0(men_men_n304_), .Y(men_men_n765_));
  NAi21      u0737(.An(men_men_n604_), .B(men_men_n94_), .Y(men_men_n766_));
  NA2        u0738(.A(men_men_n766_), .B(men_men_n765_), .Y(men_men_n767_));
  NO2        u0739(.A(men_men_n294_), .B(men_men_n138_), .Y(men_men_n768_));
  AOI220     u0740(.A0(men_men_n768_), .A1(men_men_n617_), .B0(men_men_n718_), .B1(men_men_n701_), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n725_), .B(men_men_n92_), .Y(men_men_n770_));
  NA2        u0742(.A(men_men_n770_), .B(men_men_n581_), .Y(men_men_n771_));
  NO2        u0743(.A(men_men_n583_), .B(men_men_n118_), .Y(men_men_n772_));
  OAI210     u0744(.A0(men_men_n772_), .A1(men_men_n756_), .B0(men_men_n674_), .Y(men_men_n773_));
  NA3        u0745(.A(men_men_n773_), .B(men_men_n771_), .C(men_men_n769_), .Y(men_men_n774_));
  OR4        u0746(.A(men_men_n774_), .B(men_men_n767_), .C(men_men_n763_), .D(men_men_n758_), .Y(men_men_n775_));
  NA3        u0747(.A(men_men_n761_), .B(men_men_n546_), .C(men_men_n545_), .Y(men_men_n776_));
  NA4        u0748(.A(men_men_n776_), .B(men_men_n216_), .C(men_men_n443_), .D(men_men_n34_), .Y(men_men_n777_));
  NO4        u0749(.A(men_men_n473_), .B(men_men_n427_), .C(j), .D(f), .Y(men_men_n778_));
  OAI220     u0750(.A0(men_men_n702_), .A1(n), .B0(men_men_n327_), .B1(men_men_n38_), .Y(men_men_n779_));
  AOI210     u0751(.A0(men_men_n778_), .A1(men_men_n253_), .B0(men_men_n779_), .Y(men_men_n780_));
  NA3        u0752(.A(men_men_n537_), .B(men_men_n287_), .C(h), .Y(men_men_n781_));
  NOi21      u0753(.An(men_men_n674_), .B(men_men_n781_), .Y(men_men_n782_));
  NO2        u0754(.A(men_men_n93_), .B(men_men_n47_), .Y(men_men_n783_));
  OAI220     u0755(.A0(men_men_n781_), .A1(men_men_n600_), .B0(men_men_n750_), .B1(men_men_n72_), .Y(men_men_n784_));
  AOI210     u0756(.A0(men_men_n783_), .A1(men_men_n639_), .B0(men_men_n784_), .Y(men_men_n785_));
  NAi41      u0757(.An(men_men_n782_), .B(men_men_n785_), .C(men_men_n780_), .D(men_men_n777_), .Y(men_men_n786_));
  OR2        u0758(.A(men_men_n770_), .B(men_men_n97_), .Y(men_men_n787_));
  AOI220     u0759(.A0(men_men_n787_), .A1(men_men_n234_), .B0(men_men_n756_), .B1(men_men_n631_), .Y(men_men_n788_));
  NO2        u0760(.A(men_men_n659_), .B(men_men_n74_), .Y(men_men_n789_));
  AOI210     u0761(.A0(men_men_n778_), .A1(men_men_n789_), .B0(men_men_n331_), .Y(men_men_n790_));
  OAI210     u0762(.A0(men_men_n725_), .A1(men_men_n657_), .B0(men_men_n509_), .Y(men_men_n791_));
  NA3        u0763(.A(men_men_n247_), .B(men_men_n59_), .C(b), .Y(men_men_n792_));
  AOI220     u0764(.A0(men_men_n599_), .A1(men_men_n29_), .B0(men_men_n454_), .B1(men_men_n85_), .Y(men_men_n793_));
  NA2        u0765(.A(men_men_n793_), .B(men_men_n792_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n781_), .B(men_men_n479_), .Y(men_men_n795_));
  AOI210     u0767(.A0(men_men_n794_), .A1(men_men_n791_), .B0(men_men_n795_), .Y(men_men_n796_));
  NA3        u0768(.A(men_men_n796_), .B(men_men_n790_), .C(men_men_n788_), .Y(men_men_n797_));
  NOi41      u0769(.An(men_men_n753_), .B(men_men_n797_), .C(men_men_n786_), .D(men_men_n775_), .Y(men_men_n798_));
  OR3        u0770(.A(men_men_n702_), .B(men_men_n228_), .C(g), .Y(men_men_n799_));
  NO3        u0771(.A(men_men_n337_), .B(men_men_n296_), .C(men_men_n114_), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n800_), .B(men_men_n762_), .Y(men_men_n801_));
  NA2        u0773(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n802_));
  NO3        u0774(.A(men_men_n802_), .B(men_men_n751_), .C(men_men_n273_), .Y(men_men_n803_));
  NO3        u0775(.A(men_men_n516_), .B(men_men_n95_), .C(h), .Y(men_men_n804_));
  AOI210     u0776(.A0(men_men_n804_), .A1(men_men_n697_), .B0(men_men_n803_), .Y(men_men_n805_));
  NA4        u0777(.A(men_men_n805_), .B(men_men_n801_), .C(men_men_n799_), .D(men_men_n399_), .Y(men_men_n806_));
  OR2        u0778(.A(men_men_n657_), .B(men_men_n93_), .Y(men_men_n807_));
  NOi31      u0779(.An(b), .B(d), .C(a), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n808_), .B(men_men_n597_), .Y(men_men_n809_));
  NO2        u0781(.A(men_men_n809_), .B(n), .Y(men_men_n810_));
  NOi21      u0782(.An(men_men_n793_), .B(men_men_n810_), .Y(men_men_n811_));
  OAI220     u0783(.A0(men_men_n811_), .A1(men_men_n807_), .B0(men_men_n781_), .B1(men_men_n598_), .Y(men_men_n812_));
  INV        u0784(.A(men_men_n545_), .Y(men_men_n813_));
  NO3        u0785(.A(men_men_n616_), .B(men_men_n322_), .C(men_men_n118_), .Y(men_men_n814_));
  NOi21      u0786(.An(men_men_n814_), .B(men_men_n163_), .Y(men_men_n815_));
  AOI210     u0787(.A0(men_men_n800_), .A1(men_men_n813_), .B0(men_men_n815_), .Y(men_men_n816_));
  OAI210     u0788(.A0(men_men_n702_), .A1(men_men_n389_), .B0(men_men_n816_), .Y(men_men_n817_));
  NA2        u0789(.A(men_men_n768_), .B(men_men_n664_), .Y(men_men_n818_));
  NO2        u0790(.A(men_men_n318_), .B(men_men_n233_), .Y(men_men_n819_));
  OAI210     u0791(.A0(men_men_n97_), .A1(men_men_n94_), .B0(men_men_n819_), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n122_), .B(men_men_n85_), .Y(men_men_n821_));
  AOI210     u0793(.A0(men_men_n420_), .A1(men_men_n412_), .B0(men_men_n821_), .Y(men_men_n822_));
  NAi21      u0794(.An(men_men_n822_), .B(men_men_n820_), .Y(men_men_n823_));
  NA2        u0795(.A(men_men_n723_), .B(men_men_n34_), .Y(men_men_n824_));
  NAi21      u0796(.An(men_men_n729_), .B(men_men_n428_), .Y(men_men_n825_));
  NA2        u0797(.A(men_men_n709_), .B(men_men_n345_), .Y(men_men_n826_));
  OAI210     u0798(.A0(men_men_n589_), .A1(men_men_n588_), .B0(men_men_n360_), .Y(men_men_n827_));
  AN3        u0799(.A(men_men_n827_), .B(men_men_n826_), .C(men_men_n825_), .Y(men_men_n828_));
  NAi41      u0800(.An(men_men_n823_), .B(men_men_n828_), .C(men_men_n824_), .D(men_men_n818_), .Y(men_men_n829_));
  NO4        u0801(.A(men_men_n829_), .B(men_men_n817_), .C(men_men_n812_), .D(men_men_n806_), .Y(men_men_n830_));
  NA4        u0802(.A(men_men_n830_), .B(men_men_n798_), .C(men_men_n748_), .D(men_men_n734_), .Y(men09));
  INV        u0803(.A(men_men_n123_), .Y(men_men_n832_));
  NA2        u0804(.A(f), .B(e), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n225_), .B(men_men_n114_), .Y(men_men_n834_));
  NA2        u0806(.A(men_men_n834_), .B(g), .Y(men_men_n835_));
  NA4        u0807(.A(men_men_n307_), .B(men_men_n461_), .C(men_men_n256_), .D(men_men_n120_), .Y(men_men_n836_));
  AOI210     u0808(.A0(men_men_n836_), .A1(g), .B0(men_men_n458_), .Y(men_men_n837_));
  AOI210     u0809(.A0(men_men_n837_), .A1(men_men_n835_), .B0(men_men_n833_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n437_), .B(e), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n838_), .B(men_men_n832_), .Y(men_men_n840_));
  NO2        u0812(.A(men_men_n203_), .B(men_men_n213_), .Y(men_men_n841_));
  NA3        u0813(.A(m), .B(l), .C(i), .Y(men_men_n842_));
  OAI220     u0814(.A0(men_men_n583_), .A1(men_men_n842_), .B0(men_men_n350_), .B1(men_men_n517_), .Y(men_men_n843_));
  NA4        u0815(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(f), .Y(men_men_n844_));
  NAi31      u0816(.An(men_men_n843_), .B(men_men_n844_), .C(men_men_n432_), .Y(men_men_n845_));
  OA210      u0817(.A0(men_men_n845_), .A1(men_men_n841_), .B0(men_men_n557_), .Y(men_men_n846_));
  NA3        u0818(.A(men_men_n807_), .B(men_men_n559_), .C(men_men_n509_), .Y(men_men_n847_));
  OA210      u0819(.A0(men_men_n847_), .A1(men_men_n846_), .B0(men_men_n810_), .Y(men_men_n848_));
  INV        u0820(.A(men_men_n334_), .Y(men_men_n849_));
  NO2        u0821(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n850_));
  NOi31      u0822(.An(k), .B(m), .C(l), .Y(men_men_n851_));
  NO2        u0823(.A(men_men_n336_), .B(men_men_n851_), .Y(men_men_n852_));
  AOI210     u0824(.A0(men_men_n852_), .A1(men_men_n850_), .B0(men_men_n592_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n792_), .B(men_men_n327_), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n338_), .B(men_men_n340_), .Y(men_men_n855_));
  OAI210     u0827(.A0(men_men_n203_), .A1(men_men_n213_), .B0(men_men_n855_), .Y(men_men_n856_));
  AOI220     u0828(.A0(men_men_n856_), .A1(men_men_n854_), .B0(men_men_n853_), .B1(men_men_n849_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n171_), .B(k), .Y(men_men_n858_));
  NA2        u0830(.A(men_men_n858_), .B(men_men_n693_), .Y(men_men_n859_));
  NA3        u0831(.A(men_men_n859_), .B(men_men_n191_), .C(men_men_n31_), .Y(men_men_n860_));
  NA4        u0832(.A(men_men_n860_), .B(men_men_n857_), .C(men_men_n618_), .D(men_men_n83_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n579_), .B(men_men_n487_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n862_), .B(men_men_n191_), .Y(men_men_n863_));
  NOi21      u0835(.An(f), .B(d), .Y(men_men_n864_));
  NA2        u0836(.A(men_men_n864_), .B(m), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n865_), .B(men_men_n52_), .Y(men_men_n866_));
  NOi32      u0838(.An(g), .Bn(f), .C(d), .Y(men_men_n867_));
  NA4        u0839(.A(men_men_n867_), .B(men_men_n599_), .C(men_men_n29_), .D(m), .Y(men_men_n868_));
  NOi21      u0840(.An(men_men_n308_), .B(men_men_n868_), .Y(men_men_n869_));
  AOI210     u0841(.A0(men_men_n866_), .A1(men_men_n535_), .B0(men_men_n869_), .Y(men_men_n870_));
  NA3        u0842(.A(men_men_n307_), .B(men_men_n256_), .C(men_men_n120_), .Y(men_men_n871_));
  AN2        u0843(.A(f), .B(d), .Y(men_men_n872_));
  NA3        u0844(.A(men_men_n466_), .B(men_men_n872_), .C(men_men_n85_), .Y(men_men_n873_));
  NO3        u0845(.A(men_men_n873_), .B(men_men_n74_), .C(men_men_n214_), .Y(men_men_n874_));
  INV        u0846(.A(men_men_n280_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n871_), .B(men_men_n874_), .Y(men_men_n876_));
  NAi41      u0848(.An(men_men_n478_), .B(men_men_n876_), .C(men_men_n870_), .D(men_men_n863_), .Y(men_men_n877_));
  NO4        u0849(.A(men_men_n616_), .B(men_men_n134_), .C(men_men_n322_), .D(men_men_n154_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n650_), .B(men_men_n322_), .Y(men_men_n879_));
  AN2        u0851(.A(men_men_n879_), .B(men_men_n678_), .Y(men_men_n880_));
  NO3        u0852(.A(men_men_n880_), .B(men_men_n878_), .C(men_men_n230_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n597_), .B(men_men_n85_), .Y(men_men_n882_));
  OAI220     u0854(.A0(men_men_n855_), .A1(men_men_n882_), .B0(men_men_n792_), .B1(men_men_n432_), .Y(men_men_n883_));
  NA3        u0855(.A(men_men_n162_), .B(men_men_n110_), .C(men_men_n109_), .Y(men_men_n884_));
  OAI220     u0856(.A0(men_men_n873_), .A1(men_men_n425_), .B0(men_men_n334_), .B1(men_men_n884_), .Y(men_men_n885_));
  NOi31      u0857(.An(men_men_n223_), .B(men_men_n885_), .C(men_men_n883_), .Y(men_men_n886_));
  NA2        u0858(.A(c), .B(men_men_n117_), .Y(men_men_n887_));
  NO2        u0859(.A(men_men_n887_), .B(men_men_n403_), .Y(men_men_n888_));
  NA3        u0860(.A(men_men_n888_), .B(men_men_n500_), .C(f), .Y(men_men_n889_));
  OR2        u0861(.A(men_men_n657_), .B(men_men_n532_), .Y(men_men_n890_));
  INV        u0862(.A(men_men_n890_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n809_), .B(men_men_n113_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n892_), .B(men_men_n891_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n889_), .C(men_men_n886_), .D(men_men_n881_), .Y(men_men_n894_));
  NO4        u0866(.A(men_men_n894_), .B(men_men_n877_), .C(men_men_n861_), .D(men_men_n848_), .Y(men_men_n895_));
  BUFFER     u0867(.A(men_men_n873_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n114_), .B(j), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n834_), .B(g), .Y(men_men_n898_));
  AOI210     u0870(.A0(men_men_n898_), .A1(men_men_n288_), .B0(men_men_n896_), .Y(men_men_n899_));
  AOI210     u0871(.A0(men_men_n792_), .A1(men_men_n327_), .B0(men_men_n844_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n138_), .B(men_men_n134_), .Y(men_men_n901_));
  NA2        u0873(.A(men_men_n301_), .B(men_men_n901_), .Y(men_men_n902_));
  NO2        u0874(.A(men_men_n425_), .B(men_men_n833_), .Y(men_men_n903_));
  NA2        u0875(.A(men_men_n903_), .B(men_men_n551_), .Y(men_men_n904_));
  NA2        u0876(.A(men_men_n904_), .B(men_men_n902_), .Y(men_men_n905_));
  NA2        u0877(.A(e), .B(d), .Y(men_men_n906_));
  NA2        u0878(.A(men_men_n617_), .B(men_men_n343_), .Y(men_men_n907_));
  NA2        u0879(.A(men_men_n280_), .B(men_men_n168_), .Y(men_men_n908_));
  NA2        u0880(.A(men_men_n874_), .B(men_men_n908_), .Y(men_men_n909_));
  NA3        u0881(.A(n), .B(men_men_n86_), .C(men_men_n34_), .Y(men_men_n910_));
  NA3        u0882(.A(men_men_n910_), .B(men_men_n909_), .C(men_men_n907_), .Y(men_men_n911_));
  NO4        u0883(.A(men_men_n911_), .B(men_men_n905_), .C(men_men_n900_), .D(men_men_n899_), .Y(men_men_n912_));
  NA2        u0884(.A(men_men_n849_), .B(men_men_n31_), .Y(men_men_n913_));
  OR2        u0885(.A(men_men_n913_), .B(men_men_n217_), .Y(men_men_n914_));
  NO2        u0886(.A(men_men_n296_), .B(j), .Y(men_men_n915_));
  AOI220     u0887(.A0(men_men_n915_), .A1(men_men_n879_), .B0(men_men_n609_), .B1(men_men_n615_), .Y(men_men_n916_));
  NA2        u0888(.A(men_men_n839_), .B(men_men_n916_), .Y(men_men_n917_));
  OAI210     u0889(.A0(men_men_n834_), .A1(men_men_n908_), .B0(men_men_n867_), .Y(men_men_n918_));
  NO2        u0890(.A(men_men_n918_), .B(men_men_n600_), .Y(men_men_n919_));
  AOI210     u0891(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n255_), .Y(men_men_n920_));
  NO2        u0892(.A(men_men_n920_), .B(men_men_n868_), .Y(men_men_n921_));
  AO210      u0893(.A0(men_men_n854_), .A1(men_men_n843_), .B0(men_men_n921_), .Y(men_men_n922_));
  NOi31      u0894(.An(men_men_n535_), .B(men_men_n865_), .C(men_men_n288_), .Y(men_men_n923_));
  NO4        u0895(.A(men_men_n923_), .B(men_men_n922_), .C(men_men_n919_), .D(men_men_n917_), .Y(men_men_n924_));
  NO2        u0896(.A(men_men_n431_), .B(men_men_n70_), .Y(men_men_n925_));
  OAI210     u0897(.A0(men_men_n847_), .A1(men_men_n925_), .B0(men_men_n697_), .Y(men_men_n926_));
  AN4        u0898(.A(men_men_n926_), .B(men_men_n330_), .C(men_men_n924_), .D(men_men_n914_), .Y(men_men_n927_));
  NA4        u0899(.A(men_men_n927_), .B(men_men_n912_), .C(men_men_n895_), .D(men_men_n840_), .Y(men12));
  NO2        u0900(.A(men_men_n446_), .B(c), .Y(men_men_n929_));
  NO4        u0901(.A(men_men_n436_), .B(men_men_n250_), .C(men_men_n575_), .D(men_men_n214_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n930_), .B(men_men_n929_), .Y(men_men_n931_));
  NA2        u0903(.A(men_men_n535_), .B(men_men_n925_), .Y(men_men_n932_));
  NO2        u0904(.A(men_men_n446_), .B(men_men_n117_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n850_), .B(men_men_n350_), .Y(men_men_n934_));
  NO2        u0906(.A(men_men_n657_), .B(men_men_n377_), .Y(men_men_n935_));
  AOI220     u0907(.A0(men_men_n935_), .A1(men_men_n534_), .B0(men_men_n934_), .B1(men_men_n933_), .Y(men_men_n936_));
  NA4        u0908(.A(men_men_n936_), .B(men_men_n932_), .C(men_men_n931_), .D(men_men_n435_), .Y(men_men_n937_));
  AOI210     u0909(.A0(men_men_n229_), .A1(men_men_n333_), .B0(men_men_n200_), .Y(men_men_n938_));
  NO2        u0910(.A(men_men_n330_), .B(men_men_n214_), .Y(men_men_n939_));
  NA2        u0911(.A(men_men_n939_), .B(f), .Y(men_men_n940_));
  NO2        u0912(.A(men_men_n636_), .B(men_men_n258_), .Y(men_men_n941_));
  NO2        u0913(.A(men_men_n583_), .B(men_men_n842_), .Y(men_men_n942_));
  AOI220     u0914(.A0(men_men_n942_), .A1(men_men_n557_), .B0(men_men_n819_), .B1(men_men_n941_), .Y(men_men_n943_));
  NO2        u0915(.A(men_men_n153_), .B(men_men_n233_), .Y(men_men_n944_));
  NA3        u0916(.A(men_men_n944_), .B(men_men_n236_), .C(i), .Y(men_men_n945_));
  NA3        u0917(.A(men_men_n945_), .B(men_men_n943_), .C(men_men_n940_), .Y(men_men_n946_));
  OR2        u0918(.A(men_men_n1514_), .B(men_men_n933_), .Y(men_men_n947_));
  NA2        u0919(.A(men_men_n947_), .B(men_men_n351_), .Y(men_men_n948_));
  NO3        u0920(.A(men_men_n134_), .B(men_men_n154_), .C(men_men_n214_), .Y(men_men_n949_));
  NA2        u0921(.A(men_men_n949_), .B(men_men_n521_), .Y(men_men_n950_));
  NA4        u0922(.A(men_men_n437_), .B(men_men_n429_), .C(men_men_n183_), .D(g), .Y(men_men_n951_));
  NA3        u0923(.A(men_men_n951_), .B(men_men_n950_), .C(men_men_n948_), .Y(men_men_n952_));
  NO3        u0924(.A(men_men_n662_), .B(men_men_n93_), .C(men_men_n45_), .Y(men_men_n953_));
  NO4        u0925(.A(men_men_n953_), .B(men_men_n952_), .C(men_men_n946_), .D(men_men_n937_), .Y(men_men_n954_));
  NO2        u0926(.A(men_men_n367_), .B(men_men_n366_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n580_), .B(men_men_n72_), .Y(men_men_n956_));
  NA2        u0928(.A(men_men_n545_), .B(men_men_n147_), .Y(men_men_n957_));
  NOi21      u0929(.An(men_men_n34_), .B(men_men_n650_), .Y(men_men_n958_));
  AOI220     u0930(.A0(men_men_n958_), .A1(men_men_n957_), .B0(men_men_n956_), .B1(men_men_n955_), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n248_), .A1(men_men_n45_), .B0(men_men_n959_), .Y(men_men_n960_));
  NA2        u0932(.A(men_men_n428_), .B(men_men_n260_), .Y(men_men_n961_));
  NO3        u0933(.A(men_men_n821_), .B(men_men_n90_), .C(men_men_n403_), .Y(men_men_n962_));
  NAi21      u0934(.An(men_men_n962_), .B(men_men_n961_), .Y(men_men_n963_));
  NO2        u0935(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n494_), .B(men_men_n296_), .Y(men_men_n965_));
  NO2        u0937(.A(men_men_n965_), .B(men_men_n363_), .Y(men_men_n966_));
  NO2        u0938(.A(men_men_n966_), .B(men_men_n147_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n627_), .B(men_men_n360_), .Y(men_men_n968_));
  OAI210     u0940(.A0(men_men_n730_), .A1(men_men_n968_), .B0(men_men_n364_), .Y(men_men_n969_));
  NO4        u0941(.A(men_men_n969_), .B(men_men_n967_), .C(men_men_n963_), .D(men_men_n960_), .Y(men_men_n970_));
  NA2        u0942(.A(men_men_n343_), .B(g), .Y(men_men_n971_));
  NA2        u0943(.A(men_men_n165_), .B(i), .Y(men_men_n972_));
  NA2        u0944(.A(men_men_n46_), .B(i), .Y(men_men_n973_));
  OAI220     u0945(.A0(men_men_n973_), .A1(men_men_n199_), .B0(men_men_n972_), .B1(men_men_n93_), .Y(men_men_n974_));
  AOI210     u0946(.A0(men_men_n414_), .A1(men_men_n37_), .B0(men_men_n974_), .Y(men_men_n975_));
  NO2        u0947(.A(men_men_n147_), .B(men_men_n85_), .Y(men_men_n976_));
  OR2        u0948(.A(men_men_n976_), .B(men_men_n544_), .Y(men_men_n977_));
  NA2        u0949(.A(men_men_n545_), .B(men_men_n381_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n978_), .B(men_men_n977_), .Y(men_men_n979_));
  OAI220     u0951(.A0(men_men_n979_), .A1(men_men_n971_), .B0(men_men_n975_), .B1(men_men_n327_), .Y(men_men_n980_));
  NO2        u0952(.A(men_men_n657_), .B(men_men_n487_), .Y(men_men_n981_));
  NA3        u0953(.A(men_men_n338_), .B(men_men_n622_), .C(i), .Y(men_men_n982_));
  OAI210     u0954(.A0(men_men_n431_), .A1(men_men_n307_), .B0(men_men_n982_), .Y(men_men_n983_));
  OAI220     u0955(.A0(men_men_n983_), .A1(men_men_n981_), .B0(men_men_n674_), .B1(men_men_n755_), .Y(men_men_n984_));
  NA2        u0956(.A(men_men_n603_), .B(men_men_n115_), .Y(men_men_n985_));
  OR3        u0957(.A(men_men_n307_), .B(men_men_n427_), .C(f), .Y(men_men_n986_));
  NA3        u0958(.A(men_men_n622_), .B(men_men_n81_), .C(i), .Y(men_men_n987_));
  OA220      u0959(.A0(men_men_n987_), .A1(men_men_n985_), .B0(men_men_n986_), .B1(men_men_n582_), .Y(men_men_n988_));
  NA2        u0960(.A(men_men_n934_), .B(men_men_n1514_), .Y(men_men_n989_));
  NA2        u0961(.A(men_men_n686_), .B(men_men_n882_), .Y(men_men_n990_));
  NA2        u0962(.A(men_men_n844_), .B(men_men_n432_), .Y(men_men_n991_));
  NA2        u0963(.A(i), .B(men_men_n78_), .Y(men_men_n992_));
  NA3        u0964(.A(men_men_n992_), .B(men_men_n987_), .C(men_men_n986_), .Y(men_men_n993_));
  AOI220     u0965(.A0(men_men_n993_), .A1(men_men_n253_), .B0(men_men_n991_), .B1(men_men_n990_), .Y(men_men_n994_));
  NA4        u0966(.A(men_men_n994_), .B(men_men_n989_), .C(men_men_n988_), .D(men_men_n984_), .Y(men_men_n995_));
  NA2        u0967(.A(men_men_n941_), .B(men_men_n234_), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n661_), .B(men_men_n89_), .Y(men_men_n997_));
  NO2        u0969(.A(men_men_n449_), .B(men_men_n214_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n947_), .B(men_men_n218_), .Y(men_men_n999_));
  AOI220     u0971(.A0(men_men_n935_), .A1(men_men_n944_), .B0(men_men_n581_), .B1(men_men_n91_), .Y(men_men_n1000_));
  NA4        u0972(.A(men_men_n1000_), .B(men_men_n999_), .C(men_men_n997_), .D(men_men_n996_), .Y(men_men_n1001_));
  OAI210     u0973(.A0(men_men_n991_), .A1(men_men_n942_), .B0(men_men_n534_), .Y(men_men_n1002_));
  AOI210     u0974(.A0(men_men_n415_), .A1(men_men_n407_), .B0(men_men_n821_), .Y(men_men_n1003_));
  OAI210     u0975(.A0(men_men_n367_), .A1(men_men_n366_), .B0(men_men_n111_), .Y(men_men_n1004_));
  AOI210     u0976(.A0(men_men_n1004_), .A1(men_men_n526_), .B0(men_men_n1003_), .Y(men_men_n1005_));
  NO3        u0977(.A(men_men_n897_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1006_));
  AOI220     u0978(.A0(men_men_n1006_), .A1(men_men_n620_), .B0(men_men_n641_), .B1(men_men_n521_), .Y(men_men_n1007_));
  NA3        u0979(.A(men_men_n1007_), .B(men_men_n1005_), .C(men_men_n1002_), .Y(men_men_n1008_));
  NO4        u0980(.A(men_men_n1008_), .B(men_men_n1001_), .C(men_men_n995_), .D(men_men_n980_), .Y(men_men_n1009_));
  NAi31      u0981(.An(men_men_n143_), .B(men_men_n416_), .C(n), .Y(men_men_n1010_));
  NO2        u0982(.A(m), .B(men_men_n1010_), .Y(men_men_n1011_));
  NO3        u0983(.A(men_men_n268_), .B(men_men_n143_), .C(men_men_n403_), .Y(men_men_n1012_));
  AOI210     u0984(.A0(men_men_n1012_), .A1(men_men_n488_), .B0(men_men_n1011_), .Y(men_men_n1013_));
  NA2        u0985(.A(men_men_n481_), .B(i), .Y(men_men_n1014_));
  NA2        u0986(.A(men_men_n1014_), .B(men_men_n1013_), .Y(men_men_n1015_));
  NA2        u0987(.A(men_men_n227_), .B(men_men_n174_), .Y(men_men_n1016_));
  NO3        u0988(.A(men_men_n304_), .B(men_men_n437_), .C(men_men_n177_), .Y(men_men_n1017_));
  NOi21      u0989(.An(men_men_n1016_), .B(men_men_n1017_), .Y(men_men_n1018_));
  NAi21      u0990(.An(men_men_n545_), .B(men_men_n998_), .Y(men_men_n1019_));
  NA2        u0991(.A(men_men_n430_), .B(men_men_n882_), .Y(men_men_n1020_));
  NO3        u0992(.A(men_men_n431_), .B(men_men_n307_), .C(men_men_n74_), .Y(men_men_n1021_));
  NA2        u0993(.A(men_men_n1021_), .B(men_men_n1020_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n1022_), .B(men_men_n1019_), .Y(men_men_n1023_));
  NO2        u0995(.A(men_men_n982_), .B(men_men_n598_), .Y(men_men_n1024_));
  NO2        u0996(.A(men_men_n658_), .B(men_men_n377_), .Y(men_men_n1025_));
  NA2        u0997(.A(men_men_n938_), .B(men_men_n929_), .Y(men_men_n1026_));
  NO3        u0998(.A(c), .B(men_men_n152_), .C(men_men_n213_), .Y(men_men_n1027_));
  OAI210     u0999(.A0(men_men_n1027_), .A1(men_men_n515_), .B0(men_men_n378_), .Y(men_men_n1028_));
  OAI220     u1000(.A0(men_men_n935_), .A1(men_men_n942_), .B0(men_men_n535_), .B1(men_men_n424_), .Y(men_men_n1029_));
  NA4        u1001(.A(men_men_n1029_), .B(men_men_n1028_), .C(men_men_n1026_), .D(men_men_n614_), .Y(men_men_n1030_));
  NA3        u1002(.A(men_men_n978_), .B(men_men_n475_), .C(men_men_n46_), .Y(men_men_n1031_));
  AOI210     u1003(.A0(men_men_n380_), .A1(men_men_n378_), .B0(men_men_n326_), .Y(men_men_n1032_));
  NA3        u1004(.A(men_men_n1032_), .B(men_men_n1031_), .C(men_men_n269_), .Y(men_men_n1033_));
  OR4        u1005(.A(men_men_n1033_), .B(men_men_n1030_), .C(men_men_n1025_), .D(men_men_n1024_), .Y(men_men_n1034_));
  NO4        u1006(.A(men_men_n1034_), .B(men_men_n1023_), .C(men_men_n1018_), .D(men_men_n1015_), .Y(men_men_n1035_));
  NA4        u1007(.A(men_men_n1035_), .B(men_men_n1009_), .C(men_men_n970_), .D(men_men_n954_), .Y(men13));
  NA2        u1008(.A(men_men_n46_), .B(men_men_n88_), .Y(men_men_n1037_));
  AN2        u1009(.A(c), .B(b), .Y(men_men_n1038_));
  NA3        u1010(.A(men_men_n247_), .B(men_men_n1038_), .C(m), .Y(men_men_n1039_));
  NO4        u1011(.A(e), .B(men_men_n1039_), .C(men_men_n1037_), .D(men_men_n576_), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n260_), .B(men_men_n1038_), .Y(men_men_n1041_));
  NO4        u1013(.A(men_men_n1041_), .B(e), .C(men_men_n972_), .D(a), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1043_));
  NO4        u1015(.A(men_men_n1043_), .B(d), .C(men_men_n583_), .D(men_men_n303_), .Y(men_men_n1044_));
  NA2        u1016(.A(men_men_n665_), .B(men_men_n224_), .Y(men_men_n1045_));
  NA2        u1017(.A(men_men_n406_), .B(men_men_n213_), .Y(men_men_n1046_));
  AN2        u1018(.A(d), .B(c), .Y(men_men_n1047_));
  NA2        u1019(.A(men_men_n1047_), .B(men_men_n117_), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n1048_), .B(men_men_n1046_), .C(men_men_n178_), .Y(men_men_n1049_));
  NO3        u1021(.A(men_men_n1043_), .B(men_men_n579_), .C(men_men_n303_), .Y(men_men_n1050_));
  AO210      u1022(.A0(men_men_n1049_), .A1(men_men_n1045_), .B0(men_men_n1050_), .Y(men_men_n1051_));
  OR4        u1023(.A(men_men_n1051_), .B(men_men_n1044_), .C(men_men_n1042_), .D(men_men_n1040_), .Y(men_men_n1052_));
  NAi32      u1024(.An(f), .Bn(e), .C(c), .Y(men_men_n1053_));
  OR2        u1025(.A(men_men_n224_), .B(men_men_n178_), .Y(men_men_n1054_));
  NO2        u1026(.A(men_men_n1054_), .B(men_men_n1053_), .Y(men_men_n1055_));
  INV        u1027(.A(men_men_n303_), .Y(men_men_n1056_));
  NA2        u1028(.A(men_men_n624_), .B(men_men_n1512_), .Y(men_men_n1057_));
  NOi21      u1029(.An(men_men_n1056_), .B(men_men_n1057_), .Y(men_men_n1058_));
  NO2        u1030(.A(men_men_n759_), .B(men_men_n114_), .Y(men_men_n1059_));
  NOi41      u1031(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n1060_), .B(men_men_n1059_), .Y(men_men_n1061_));
  NO2        u1033(.A(men_men_n1061_), .B(men_men_n1053_), .Y(men_men_n1062_));
  NA3        u1034(.A(k), .B(j), .C(i), .Y(men_men_n1063_));
  NO3        u1035(.A(men_men_n1063_), .B(men_men_n303_), .C(men_men_n92_), .Y(men_men_n1064_));
  OR4        u1036(.A(men_men_n1064_), .B(men_men_n1062_), .C(men_men_n1058_), .D(men_men_n1055_), .Y(men_men_n1065_));
  NA3        u1037(.A(men_men_n457_), .B(men_men_n329_), .C(men_men_n56_), .Y(men_men_n1066_));
  NO3        u1038(.A(men_men_n1066_), .B(men_men_n579_), .C(men_men_n45_), .Y(men_men_n1067_));
  NO2        u1039(.A(f), .B(c), .Y(men_men_n1068_));
  NOi21      u1040(.An(men_men_n1068_), .B(men_men_n436_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n1069_), .B(men_men_n59_), .Y(men_men_n1070_));
  NO3        u1042(.A(k), .B(men_men_n240_), .C(l), .Y(men_men_n1071_));
  NOi21      u1043(.An(men_men_n1071_), .B(men_men_n1070_), .Y(men_men_n1072_));
  OR2        u1044(.A(men_men_n1072_), .B(men_men_n1067_), .Y(men_men_n1073_));
  OR3        u1045(.A(men_men_n1073_), .B(men_men_n1065_), .C(men_men_n1052_), .Y(men02));
  OR2        u1046(.A(l), .B(k), .Y(men_men_n1075_));
  OR3        u1047(.A(h), .B(g), .C(f), .Y(men_men_n1076_));
  OR3        u1048(.A(n), .B(m), .C(i), .Y(men_men_n1077_));
  NO4        u1049(.A(men_men_n1077_), .B(men_men_n1076_), .C(men_men_n1075_), .D(e), .Y(men_men_n1078_));
  NO2        u1050(.A(men_men_n1064_), .B(men_men_n1044_), .Y(men_men_n1079_));
  NA3        u1051(.A(g), .B(men_men_n457_), .C(h), .Y(men_men_n1080_));
  OR2        u1052(.A(men_men_n303_), .B(men_men_n1080_), .Y(men_men_n1081_));
  NO3        u1053(.A(men_men_n1066_), .B(men_men_n1043_), .C(men_men_n579_), .Y(men_men_n1082_));
  NO2        u1054(.A(men_men_n1082_), .B(men_men_n1055_), .Y(men_men_n1083_));
  NA3        u1055(.A(l), .B(k), .C(j), .Y(men_men_n1084_));
  NA2        u1056(.A(i), .B(h), .Y(men_men_n1085_));
  NO2        u1057(.A(men_men_n1085_), .B(men_men_n1084_), .Y(men_men_n1086_));
  NO3        u1058(.A(men_men_n144_), .B(men_men_n278_), .C(men_men_n214_), .Y(men_men_n1087_));
  AOI210     u1059(.A0(men_men_n1087_), .A1(men_men_n1086_), .B0(men_men_n1058_), .Y(men_men_n1088_));
  NA3        u1060(.A(c), .B(b), .C(a), .Y(men_men_n1089_));
  NO3        u1061(.A(men_men_n1089_), .B(men_men_n906_), .C(men_men_n213_), .Y(men_men_n1090_));
  AN3        u1062(.A(men_men_n1088_), .B(men_men_n1083_), .C(men_men_n1081_), .Y(men_men_n1091_));
  NO2        u1063(.A(men_men_n1048_), .B(men_men_n1046_), .Y(men_men_n1092_));
  AOI210     u1064(.A0(l), .A1(men_men_n1092_), .B0(men_men_n1040_), .Y(men_men_n1093_));
  NAi41      u1065(.An(men_men_n1078_), .B(men_men_n1093_), .C(men_men_n1091_), .D(men_men_n1079_), .Y(men03));
  NO2        u1066(.A(men_men_n517_), .B(men_men_n592_), .Y(men_men_n1095_));
  NA4        u1067(.A(men_men_n89_), .B(men_men_n88_), .C(g), .D(men_men_n213_), .Y(men_men_n1096_));
  NA4        u1068(.A(men_men_n567_), .B(m), .C(men_men_n114_), .D(men_men_n213_), .Y(men_men_n1097_));
  NA3        u1069(.A(men_men_n1097_), .B(men_men_n368_), .C(men_men_n1096_), .Y(men_men_n1098_));
  NO3        u1070(.A(men_men_n1098_), .B(men_men_n1095_), .C(men_men_n1004_), .Y(men_men_n1099_));
  NOi41      u1071(.An(men_men_n807_), .B(men_men_n856_), .C(men_men_n845_), .D(men_men_n711_), .Y(men_men_n1100_));
  OAI220     u1072(.A0(men_men_n1100_), .A1(men_men_n686_), .B0(men_men_n1099_), .B1(men_men_n580_), .Y(men_men_n1101_));
  NOi31      u1073(.An(i), .B(k), .C(j), .Y(men_men_n1102_));
  NA4        u1074(.A(men_men_n1102_), .B(e), .C(men_men_n338_), .D(men_men_n329_), .Y(men_men_n1103_));
  OAI210     u1075(.A0(men_men_n821_), .A1(men_men_n417_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  NOi31      u1076(.An(m), .B(n), .C(f), .Y(men_men_n1105_));
  NA2        u1077(.A(men_men_n1105_), .B(men_men_n51_), .Y(men_men_n1106_));
  AN2        u1078(.A(e), .B(c), .Y(men_men_n1107_));
  NA2        u1079(.A(men_men_n1107_), .B(a), .Y(men_men_n1108_));
  OAI220     u1080(.A0(men_men_n1108_), .A1(men_men_n1106_), .B0(men_men_n890_), .B1(men_men_n423_), .Y(men_men_n1109_));
  NA2        u1081(.A(men_men_n498_), .B(l), .Y(men_men_n1110_));
  NOi31      u1082(.An(men_men_n867_), .B(men_men_n1039_), .C(men_men_n1110_), .Y(men_men_n1111_));
  NO4        u1083(.A(men_men_n1111_), .B(men_men_n1109_), .C(men_men_n1104_), .D(men_men_n1003_), .Y(men_men_n1112_));
  NO2        u1084(.A(men_men_n278_), .B(a), .Y(men_men_n1113_));
  INV        u1085(.A(men_men_n1044_), .Y(men_men_n1114_));
  NO2        u1086(.A(men_men_n88_), .B(g), .Y(men_men_n1115_));
  AOI210     u1087(.A0(men_men_n1115_), .A1(i), .B0(men_men_n1071_), .Y(men_men_n1116_));
  OR2        u1088(.A(men_men_n1116_), .B(men_men_n1070_), .Y(men_men_n1117_));
  NA3        u1089(.A(men_men_n1117_), .B(men_men_n1114_), .C(men_men_n1112_), .Y(men_men_n1118_));
  NO4        u1090(.A(men_men_n1118_), .B(men_men_n1101_), .C(men_men_n823_), .D(men_men_n556_), .Y(men_men_n1119_));
  NA2        u1091(.A(c), .B(b), .Y(men_men_n1120_));
  NO2        u1092(.A(men_men_n696_), .B(men_men_n1120_), .Y(men_men_n1121_));
  OAI210     u1093(.A0(men_men_n865_), .A1(men_men_n837_), .B0(men_men_n410_), .Y(men_men_n1122_));
  OAI210     u1094(.A0(men_men_n1122_), .A1(men_men_n866_), .B0(men_men_n1121_), .Y(men_men_n1123_));
  NAi21      u1095(.An(men_men_n418_), .B(men_men_n1121_), .Y(men_men_n1124_));
  NA3        u1096(.A(men_men_n424_), .B(men_men_n549_), .C(f), .Y(men_men_n1125_));
  OAI210     u1097(.A0(men_men_n539_), .A1(men_men_n39_), .B0(men_men_n1113_), .Y(men_men_n1126_));
  NA3        u1098(.A(men_men_n1126_), .B(men_men_n1125_), .C(men_men_n1124_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n256_), .B(men_men_n120_), .Y(men_men_n1128_));
  OAI210     u1100(.A0(men_men_n1128_), .A1(men_men_n282_), .B0(g), .Y(men_men_n1129_));
  NO2        u1101(.A(f), .B(men_men_n1089_), .Y(men_men_n1130_));
  INV        u1102(.A(men_men_n1130_), .Y(men_men_n1131_));
  AOI210     u1103(.A0(men_men_n1129_), .A1(men_men_n288_), .B0(men_men_n1131_), .Y(men_men_n1132_));
  NO2        u1104(.A(men_men_n1132_), .B(men_men_n1127_), .Y(men_men_n1133_));
  INV        u1105(.A(men_men_n458_), .Y(men_men_n1134_));
  NO2        u1106(.A(men_men_n184_), .B(men_men_n233_), .Y(men_men_n1135_));
  NA2        u1107(.A(men_men_n1135_), .B(m), .Y(men_men_n1136_));
  NA3        u1108(.A(men_men_n920_), .B(men_men_n1110_), .C(men_men_n461_), .Y(men_men_n1137_));
  OAI210     u1109(.A0(men_men_n1137_), .A1(men_men_n308_), .B0(men_men_n459_), .Y(men_men_n1138_));
  AOI210     u1110(.A0(men_men_n1138_), .A1(men_men_n1134_), .B0(men_men_n1136_), .Y(men_men_n1139_));
  NA2        u1111(.A(men_men_n551_), .B(men_men_n405_), .Y(men_men_n1140_));
  NA2        u1112(.A(men_men_n161_), .B(men_men_n33_), .Y(men_men_n1141_));
  AOI210     u1113(.A0(men_men_n968_), .A1(men_men_n1141_), .B0(men_men_n214_), .Y(men_men_n1142_));
  NA2        u1114(.A(men_men_n1142_), .B(men_men_n1130_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n1144_));
  AOI210     u1116(.A0(men_men_n1135_), .A1(men_men_n51_), .B0(men_men_n962_), .Y(men_men_n1145_));
  NAi41      u1117(.An(men_men_n1144_), .B(men_men_n1145_), .C(men_men_n1143_), .D(men_men_n1140_), .Y(men_men_n1146_));
  NO2        u1118(.A(men_men_n1146_), .B(men_men_n1139_), .Y(men_men_n1147_));
  NA4        u1119(.A(men_men_n1147_), .B(men_men_n1133_), .C(men_men_n1123_), .D(men_men_n1119_), .Y(men00));
  NO2        u1120(.A(men_men_n295_), .B(men_men_n272_), .Y(men_men_n1149_));
  NO2        u1121(.A(men_men_n1149_), .B(men_men_n570_), .Y(men_men_n1150_));
  AOI210     u1122(.A0(men_men_n903_), .A1(men_men_n944_), .B0(men_men_n1104_), .Y(men_men_n1151_));
  NO2        u1123(.A(men_men_n962_), .B(men_men_n708_), .Y(men_men_n1152_));
  NA3        u1124(.A(men_men_n1152_), .B(men_men_n1151_), .C(men_men_n1005_), .Y(men_men_n1153_));
  NA2        u1125(.A(men_men_n500_), .B(f), .Y(men_men_n1154_));
  NA2        u1126(.A(h), .B(men_men_n252_), .Y(men_men_n1155_));
  AOI210     u1127(.A0(men_men_n1155_), .A1(men_men_n1154_), .B0(men_men_n1048_), .Y(men_men_n1156_));
  NO4        u1128(.A(men_men_n1156_), .B(men_men_n1153_), .C(men_men_n1150_), .D(men_men_n1065_), .Y(men_men_n1157_));
  NA3        u1129(.A(n), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1158_));
  NA3        u1130(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1159_));
  NOi31      u1131(.An(n), .B(m), .C(i), .Y(men_men_n1160_));
  NA3        u1132(.A(men_men_n1160_), .B(men_men_n646_), .C(men_men_n51_), .Y(men_men_n1161_));
  OAI210     u1133(.A0(men_men_n1159_), .A1(men_men_n1158_), .B0(men_men_n1161_), .Y(men_men_n1162_));
  INV        u1134(.A(men_men_n569_), .Y(men_men_n1163_));
  NO4        u1135(.A(men_men_n1163_), .B(men_men_n1162_), .C(men_men_n1144_), .D(men_men_n923_), .Y(men_men_n1164_));
  NO3        u1136(.A(men_men_n476_), .B(men_men_n353_), .C(men_men_n1120_), .Y(men_men_n1165_));
  NA3        u1137(.A(men_men_n383_), .B(men_men_n221_), .C(g), .Y(men_men_n1166_));
  OA220      u1138(.A0(men_men_n1166_), .A1(men_men_n1159_), .B0(men_men_n384_), .B1(men_men_n137_), .Y(men_men_n1167_));
  NO2        u1139(.A(h), .B(g), .Y(men_men_n1168_));
  NA4        u1140(.A(men_men_n488_), .B(men_men_n457_), .C(men_men_n1168_), .D(men_men_n1038_), .Y(men_men_n1169_));
  OAI220     u1141(.A0(men_men_n517_), .A1(men_men_n592_), .B0(men_men_n93_), .B1(men_men_n92_), .Y(men_men_n1170_));
  AOI220     u1142(.A0(men_men_n1170_), .A1(men_men_n526_), .B0(men_men_n949_), .B1(men_men_n568_), .Y(men_men_n1171_));
  AOI220     u1143(.A0(men_men_n314_), .A1(men_men_n244_), .B0(men_men_n179_), .B1(men_men_n151_), .Y(men_men_n1172_));
  NA4        u1144(.A(men_men_n1172_), .B(men_men_n1171_), .C(men_men_n1169_), .D(men_men_n1167_), .Y(men_men_n1173_));
  NO3        u1145(.A(men_men_n1173_), .B(men_men_n1165_), .C(men_men_n262_), .Y(men_men_n1174_));
  INV        u1146(.A(men_men_n317_), .Y(men_men_n1175_));
  AOI210     u1147(.A0(men_men_n244_), .A1(men_men_n343_), .B0(men_men_n571_), .Y(men_men_n1176_));
  NA3        u1148(.A(men_men_n1176_), .B(men_men_n1175_), .C(men_men_n156_), .Y(men_men_n1177_));
  NO2        u1149(.A(men_men_n235_), .B(men_men_n183_), .Y(men_men_n1178_));
  NA2        u1150(.A(men_men_n1178_), .B(men_men_n424_), .Y(men_men_n1179_));
  NA3        u1151(.A(men_men_n181_), .B(men_men_n114_), .C(g), .Y(men_men_n1180_));
  NA3        u1152(.A(men_men_n457_), .B(men_men_n40_), .C(f), .Y(men_men_n1181_));
  NOi31      u1153(.An(men_men_n875_), .B(men_men_n1181_), .C(men_men_n1180_), .Y(men_men_n1182_));
  NAi31      u1154(.An(men_men_n187_), .B(men_men_n862_), .C(men_men_n457_), .Y(men_men_n1183_));
  NAi31      u1155(.An(men_men_n1182_), .B(men_men_n1183_), .C(men_men_n1179_), .Y(men_men_n1184_));
  NO2        u1156(.A(men_men_n271_), .B(men_men_n74_), .Y(men_men_n1185_));
  NO3        u1157(.A(men_men_n423_), .B(men_men_n833_), .C(n), .Y(men_men_n1186_));
  AOI210     u1158(.A0(men_men_n1186_), .A1(men_men_n1185_), .B0(men_men_n1078_), .Y(men_men_n1187_));
  NAi31      u1159(.An(men_men_n1050_), .B(men_men_n1187_), .C(men_men_n73_), .Y(men_men_n1188_));
  NO4        u1160(.A(men_men_n1188_), .B(men_men_n1184_), .C(men_men_n1177_), .D(men_men_n508_), .Y(men_men_n1189_));
  AN3        u1161(.A(men_men_n1189_), .B(men_men_n1174_), .C(men_men_n1164_), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n526_), .B(men_men_n103_), .Y(men_men_n1191_));
  NA3        u1163(.A(men_men_n1105_), .B(men_men_n603_), .C(men_men_n456_), .Y(men_men_n1192_));
  NA4        u1164(.A(men_men_n1192_), .B(men_men_n552_), .C(men_men_n1191_), .D(men_men_n238_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n1098_), .B(men_men_n526_), .Y(men_men_n1194_));
  NA4        u1166(.A(men_men_n646_), .B(men_men_n205_), .C(men_men_n221_), .D(men_men_n165_), .Y(men_men_n1195_));
  NA3        u1167(.A(men_men_n1195_), .B(men_men_n1194_), .C(men_men_n292_), .Y(men_men_n1196_));
  OAI210     u1168(.A0(men_men_n455_), .A1(men_men_n121_), .B0(men_men_n868_), .Y(men_men_n1197_));
  AOI220     u1169(.A0(men_men_n1197_), .A1(men_men_n1137_), .B0(men_men_n551_), .B1(men_men_n405_), .Y(men_men_n1198_));
  OR4        u1170(.A(men_men_n1048_), .B(men_men_n268_), .C(men_men_n222_), .D(e), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n217_), .B(men_men_n214_), .Y(men_men_n1200_));
  NA2        u1172(.A(n), .B(e), .Y(men_men_n1201_));
  NO2        u1173(.A(men_men_n1201_), .B(men_men_n149_), .Y(men_men_n1202_));
  AOI220     u1174(.A0(men_men_n1202_), .A1(men_men_n270_), .B0(men_men_n849_), .B1(men_men_n1200_), .Y(men_men_n1203_));
  OAI210     u1175(.A0(men_men_n354_), .A1(men_men_n309_), .B0(men_men_n441_), .Y(men_men_n1204_));
  NA4        u1176(.A(men_men_n1204_), .B(men_men_n1203_), .C(men_men_n1199_), .D(men_men_n1198_), .Y(men_men_n1205_));
  AOI210     u1177(.A0(men_men_n1202_), .A1(men_men_n853_), .B0(men_men_n822_), .Y(men_men_n1206_));
  AOI220     u1178(.A0(men_men_n958_), .A1(men_men_n568_), .B0(men_men_n646_), .B1(men_men_n241_), .Y(men_men_n1207_));
  NO2        u1179(.A(men_men_n67_), .B(h), .Y(men_men_n1208_));
  NO3        u1180(.A(men_men_n1048_), .B(men_men_n1046_), .C(men_men_n1515_), .Y(men_men_n1209_));
  NO2        u1181(.A(men_men_n1075_), .B(men_men_n134_), .Y(men_men_n1210_));
  AN2        u1182(.A(men_men_n1210_), .B(men_men_n1087_), .Y(men_men_n1211_));
  OAI210     u1183(.A0(men_men_n1211_), .A1(men_men_n1209_), .B0(men_men_n1208_), .Y(men_men_n1212_));
  NA4        u1184(.A(men_men_n1212_), .B(men_men_n1207_), .C(men_men_n1206_), .D(men_men_n870_), .Y(men_men_n1213_));
  NO4        u1185(.A(men_men_n1213_), .B(men_men_n1205_), .C(men_men_n1196_), .D(men_men_n1193_), .Y(men_men_n1214_));
  NA2        u1186(.A(men_men_n838_), .B(men_men_n754_), .Y(men_men_n1215_));
  NA4        u1187(.A(men_men_n1215_), .B(men_men_n1214_), .C(men_men_n1190_), .D(men_men_n1157_), .Y(men01));
  AN2        u1188(.A(men_men_n1028_), .B(men_men_n1026_), .Y(men_men_n1217_));
  NO3        u1189(.A(men_men_n803_), .B(men_men_n795_), .C(men_men_n469_), .Y(men_men_n1218_));
  NO2        u1190(.A(men_men_n585_), .B(men_men_n285_), .Y(men_men_n1219_));
  NA2        u1191(.A(men_men_n1219_), .B(i), .Y(men_men_n1220_));
  NA3        u1192(.A(men_men_n1220_), .B(men_men_n1218_), .C(men_men_n1217_), .Y(men_men_n1221_));
  NA2        u1193(.A(men_men_n581_), .B(men_men_n91_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n545_), .B(men_men_n267_), .Y(men_men_n1223_));
  NA2        u1195(.A(men_men_n965_), .B(men_men_n1223_), .Y(men_men_n1224_));
  NA4        u1196(.A(men_men_n1224_), .B(men_men_n1222_), .C(men_men_n916_), .D(men_men_n328_), .Y(men_men_n1225_));
  NA2        u1197(.A(men_men_n703_), .B(men_men_n98_), .Y(men_men_n1226_));
  NO2        u1198(.A(men_men_n1226_), .B(i), .Y(men_men_n1227_));
  OAI210     u1199(.A0(men_men_n781_), .A1(men_men_n598_), .B0(men_men_n1195_), .Y(men_men_n1228_));
  AOI210     u1200(.A0(men_men_n1227_), .A1(men_men_n631_), .B0(men_men_n1228_), .Y(men_men_n1229_));
  NA2        u1201(.A(men_men_n119_), .B(l), .Y(men_men_n1230_));
  OA220      u1202(.A0(men_men_n1230_), .A1(men_men_n578_), .B0(men_men_n659_), .B1(men_men_n368_), .Y(men_men_n1231_));
  NAi41      u1203(.An(men_men_n164_), .B(men_men_n1231_), .C(men_men_n1229_), .D(men_men_n902_), .Y(men_men_n1232_));
  NO2        u1204(.A(men_men_n782_), .B(men_men_n673_), .Y(men_men_n1233_));
  NA4        u1205(.A(men_men_n703_), .B(men_men_n98_), .C(men_men_n45_), .D(men_men_n213_), .Y(men_men_n1234_));
  NA2        u1206(.A(men_men_n1233_), .B(men_men_n140_), .Y(men_men_n1235_));
  NO4        u1207(.A(men_men_n1235_), .B(men_men_n1232_), .C(men_men_n1225_), .D(men_men_n1221_), .Y(men_men_n1236_));
  NA2        u1208(.A(men_men_n1166_), .B(men_men_n206_), .Y(men_men_n1237_));
  OAI210     u1209(.A0(men_men_n1237_), .A1(men_men_n298_), .B0(men_men_n521_), .Y(men_men_n1238_));
  NA2        u1210(.A(men_men_n529_), .B(men_men_n392_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n75_), .B(i), .Y(men_men_n1240_));
  AOI210     u1212(.A0(men_men_n584_), .A1(men_men_n578_), .B0(men_men_n1240_), .Y(men_men_n1241_));
  AOI210     u1213(.A0(men_men_n553_), .A1(men_men_n1239_), .B0(men_men_n1241_), .Y(men_men_n1242_));
  AOI210     u1214(.A0(men_men_n203_), .A1(men_men_n90_), .B0(men_men_n213_), .Y(men_men_n1243_));
  OAI210     u1215(.A0(men_men_n810_), .A1(men_men_n424_), .B0(men_men_n1243_), .Y(men_men_n1244_));
  AN3        u1216(.A(m), .B(l), .C(k), .Y(men_men_n1245_));
  OAI210     u1217(.A0(men_men_n356_), .A1(men_men_n34_), .B0(men_men_n1245_), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n202_), .B(men_men_n34_), .Y(men_men_n1247_));
  AO210      u1219(.A0(men_men_n1247_), .A1(men_men_n1246_), .B0(men_men_n327_), .Y(men_men_n1248_));
  NA4        u1220(.A(men_men_n1248_), .B(men_men_n1244_), .C(men_men_n1242_), .D(men_men_n1238_), .Y(men_men_n1249_));
  AOI210     u1221(.A0(men_men_n590_), .A1(men_men_n119_), .B0(men_men_n596_), .Y(men_men_n1250_));
  OAI210     u1222(.A0(men_men_n1230_), .A1(men_men_n587_), .B0(men_men_n1250_), .Y(men_men_n1251_));
  NA2        u1223(.A(men_men_n277_), .B(men_men_n195_), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n1252_), .B(men_men_n664_), .Y(men_men_n1253_));
  NO3        u1225(.A(men_men_n821_), .B(men_men_n203_), .C(men_men_n403_), .Y(men_men_n1254_));
  NO2        u1226(.A(men_men_n1254_), .B(men_men_n962_), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n1227_), .A1(men_men_n321_), .B0(men_men_n674_), .Y(men_men_n1256_));
  NA4        u1228(.A(men_men_n1256_), .B(men_men_n1255_), .C(men_men_n1253_), .D(men_men_n785_), .Y(men_men_n1257_));
  NO3        u1229(.A(men_men_n1257_), .B(men_men_n1251_), .C(men_men_n1249_), .Y(men_men_n1258_));
  NA3        u1230(.A(men_men_n599_), .B(men_men_n29_), .C(f), .Y(men_men_n1259_));
  NO2        u1231(.A(men_men_n1259_), .B(men_men_n203_), .Y(men_men_n1260_));
  AOI210     u1232(.A0(men_men_n495_), .A1(men_men_n58_), .B0(men_men_n1260_), .Y(men_men_n1261_));
  OR3        u1233(.A(men_men_n1226_), .B(men_men_n600_), .C(i), .Y(men_men_n1262_));
  NA3        u1234(.A(men_men_n736_), .B(men_men_n75_), .C(i), .Y(men_men_n1263_));
  AOI210     u1235(.A0(men_men_n1263_), .A1(men_men_n1234_), .B0(men_men_n985_), .Y(men_men_n1264_));
  NO2        u1236(.A(men_men_n206_), .B(men_men_n113_), .Y(men_men_n1265_));
  NO3        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .C(men_men_n1162_), .Y(men_men_n1266_));
  NA4        u1238(.A(men_men_n1266_), .B(men_men_n1262_), .C(men_men_n1261_), .D(men_men_n753_), .Y(men_men_n1267_));
  NA2        u1239(.A(men_men_n563_), .B(men_men_n561_), .Y(men_men_n1268_));
  NO3        u1240(.A(men_men_n80_), .B(men_men_n296_), .C(men_men_n45_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n544_), .Y(men_men_n1270_));
  NA3        u1242(.A(men_men_n1270_), .B(men_men_n1268_), .C(men_men_n669_), .Y(men_men_n1271_));
  OR2        u1243(.A(men_men_n1166_), .B(men_men_n1159_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n368_), .B(men_men_n72_), .Y(men_men_n1273_));
  AOI210     u1245(.A0(men_men_n727_), .A1(men_men_n611_), .B0(men_men_n1273_), .Y(men_men_n1274_));
  NA2        u1246(.A(men_men_n1269_), .B(men_men_n813_), .Y(men_men_n1275_));
  NA4        u1247(.A(men_men_n1275_), .B(men_men_n1274_), .C(men_men_n1272_), .D(men_men_n386_), .Y(men_men_n1276_));
  NO3        u1248(.A(men_men_n1276_), .B(men_men_n1271_), .C(men_men_n1267_), .Y(men_men_n1277_));
  NO2        u1249(.A(men_men_n133_), .B(men_men_n45_), .Y(men_men_n1278_));
  AO220      u1250(.A0(i), .A1(men_men_n617_), .B0(men_men_n1278_), .B1(men_men_n701_), .Y(men_men_n1279_));
  NA2        u1251(.A(men_men_n1279_), .B(men_men_n336_), .Y(men_men_n1280_));
  NA2        u1252(.A(men_men_n450_), .B(men_men_n137_), .Y(men_men_n1281_));
  NO3        u1253(.A(men_men_n1085_), .B(men_men_n178_), .C(men_men_n88_), .Y(men_men_n1282_));
  AOI220     u1254(.A0(men_men_n1282_), .A1(men_men_n1281_), .B0(men_men_n1269_), .B1(men_men_n976_), .Y(men_men_n1283_));
  NA2        u1255(.A(men_men_n1283_), .B(men_men_n1280_), .Y(men_men_n1284_));
  NO3        u1256(.A(men_men_n450_), .B(men_men_n176_), .C(men_men_n88_), .Y(men_men_n1285_));
  NO3        u1257(.A(men_men_n1285_), .B(men_men_n1284_), .C(men_men_n635_), .Y(men_men_n1286_));
  NA4        u1258(.A(men_men_n1286_), .B(men_men_n1277_), .C(men_men_n1258_), .D(men_men_n1236_), .Y(men06));
  NO2        u1259(.A(men_men_n404_), .B(men_men_n550_), .Y(men_men_n1288_));
  NO2        u1260(.A(men_men_n729_), .B(i), .Y(men_men_n1289_));
  OAI210     u1261(.A0(men_men_n1289_), .A1(men_men_n263_), .B0(men_men_n1288_), .Y(men_men_n1290_));
  NO3        u1262(.A(men_men_n594_), .B(men_men_n808_), .C(men_men_n597_), .Y(men_men_n1291_));
  OR2        u1263(.A(men_men_n1291_), .B(men_men_n890_), .Y(men_men_n1292_));
  NA2        u1264(.A(men_men_n1292_), .B(men_men_n1290_), .Y(men_men_n1293_));
  NO3        u1265(.A(men_men_n1293_), .B(men_men_n1271_), .C(men_men_n251_), .Y(men_men_n1294_));
  NA2        u1266(.A(i), .B(men_men_n977_), .Y(men_men_n1295_));
  AOI210     u1267(.A0(i), .A1(men_men_n547_), .B0(men_men_n1279_), .Y(men_men_n1296_));
  AOI210     u1268(.A0(men_men_n1296_), .A1(men_men_n1295_), .B0(men_men_n333_), .Y(men_men_n1297_));
  OAI210     u1269(.A0(men_men_n90_), .A1(men_men_n40_), .B0(men_men_n672_), .Y(men_men_n1298_));
  NA2        u1270(.A(men_men_n1298_), .B(men_men_n639_), .Y(men_men_n1299_));
  NO2        u1271(.A(men_men_n604_), .B(men_men_n1106_), .Y(men_men_n1300_));
  OAI210     u1272(.A0(men_men_n450_), .A1(men_men_n245_), .B0(men_men_n910_), .Y(men_men_n1301_));
  NO3        u1273(.A(men_men_n1301_), .B(men_men_n1300_), .C(men_men_n139_), .Y(men_men_n1302_));
  OR2        u1274(.A(men_men_n595_), .B(men_men_n593_), .Y(men_men_n1303_));
  NO2        u1275(.A(men_men_n367_), .B(men_men_n138_), .Y(men_men_n1304_));
  AOI210     u1276(.A0(men_men_n1304_), .A1(men_men_n581_), .B0(men_men_n1303_), .Y(men_men_n1305_));
  NA3        u1277(.A(men_men_n1305_), .B(men_men_n1302_), .C(men_men_n1299_), .Y(men_men_n1306_));
  NO2        u1278(.A(men_men_n744_), .B(men_men_n366_), .Y(men_men_n1307_));
  NO3        u1279(.A(men_men_n674_), .B(men_men_n755_), .C(men_men_n631_), .Y(men_men_n1308_));
  NOi21      u1280(.An(men_men_n1307_), .B(men_men_n1308_), .Y(men_men_n1309_));
  AN2        u1281(.A(men_men_n958_), .B(men_men_n642_), .Y(men_men_n1310_));
  NO4        u1282(.A(men_men_n1310_), .B(men_men_n1309_), .C(men_men_n1306_), .D(men_men_n1297_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n802_), .B(men_men_n273_), .Y(men_men_n1312_));
  OAI220     u1284(.A0(men_men_n729_), .A1(men_men_n47_), .B0(men_men_n224_), .B1(men_men_n610_), .Y(men_men_n1313_));
  OAI210     u1285(.A0(men_men_n273_), .A1(c), .B0(men_men_n638_), .Y(men_men_n1314_));
  AOI220     u1286(.A0(men_men_n1314_), .A1(men_men_n1313_), .B0(men_men_n1312_), .B1(men_men_n263_), .Y(men_men_n1315_));
  NO3        u1287(.A(men_men_n240_), .B(men_men_n105_), .C(men_men_n278_), .Y(men_men_n1316_));
  OAI210     u1288(.A0(l), .A1(i), .B0(k), .Y(men_men_n1317_));
  NO3        u1289(.A(men_men_n1317_), .B(men_men_n592_), .C(j), .Y(men_men_n1318_));
  NOi21      u1290(.An(men_men_n1318_), .B(men_men_n72_), .Y(men_men_n1319_));
  NO3        u1291(.A(men_men_n1319_), .B(men_men_n1316_), .C(men_men_n1109_), .Y(men_men_n1320_));
  NA4        u1292(.A(men_men_n793_), .B(men_men_n792_), .C(men_men_n430_), .D(men_men_n882_), .Y(men_men_n1321_));
  NAi31      u1293(.An(men_men_n744_), .B(men_men_n1321_), .C(men_men_n202_), .Y(men_men_n1322_));
  NA4        u1294(.A(men_men_n1322_), .B(men_men_n1320_), .C(men_men_n1315_), .D(men_men_n1207_), .Y(men_men_n1323_));
  NOi31      u1295(.An(men_men_n1291_), .B(men_men_n454_), .C(men_men_n391_), .Y(men_men_n1324_));
  OR3        u1296(.A(men_men_n1324_), .B(men_men_n781_), .C(men_men_n532_), .Y(men_men_n1325_));
  OR2        u1297(.A(men_men_n370_), .B(men_men_n610_), .Y(men_men_n1326_));
  AOI210     u1298(.A0(men_men_n563_), .A1(men_men_n441_), .B0(men_men_n372_), .Y(men_men_n1327_));
  NA2        u1299(.A(men_men_n1318_), .B(men_men_n789_), .Y(men_men_n1328_));
  NA4        u1300(.A(men_men_n1328_), .B(men_men_n1327_), .C(men_men_n1326_), .D(men_men_n1325_), .Y(men_men_n1329_));
  AOI220     u1301(.A0(men_men_n1307_), .A1(men_men_n754_), .B0(men_men_n1304_), .B1(men_men_n234_), .Y(men_men_n1330_));
  NO3        u1302(.A(men_men_n930_), .B(men_men_n880_), .C(men_men_n491_), .Y(men_men_n1331_));
  NA3        u1303(.A(men_men_n1331_), .B(men_men_n1330_), .C(men_men_n1275_), .Y(men_men_n1332_));
  NO4        u1304(.A(men_men_n450_), .B(j), .C(men_men_n436_), .D(men_men_n231_), .Y(men_men_n1333_));
  NO4        u1305(.A(men_men_n1333_), .B(men_men_n1332_), .C(men_men_n1329_), .D(men_men_n1323_), .Y(men_men_n1334_));
  NA4        u1306(.A(men_men_n1334_), .B(men_men_n1311_), .C(men_men_n1294_), .D(men_men_n1286_), .Y(men07));
  NOi21      u1307(.An(j), .B(k), .Y(men_men_n1336_));
  NAi32      u1308(.An(m), .Bn(b), .C(n), .Y(men_men_n1337_));
  NO3        u1309(.A(men_men_n1337_), .B(g), .C(f), .Y(men_men_n1338_));
  OAI210     u1310(.A0(men_men_n316_), .A1(men_men_n472_), .B0(men_men_n1338_), .Y(men_men_n1339_));
  NAi21      u1311(.An(f), .B(c), .Y(men_men_n1340_));
  OR2        u1312(.A(e), .B(d), .Y(men_men_n1341_));
  NOi31      u1313(.An(n), .B(m), .C(b), .Y(men_men_n1342_));
  INV        u1314(.A(men_men_n1339_), .Y(men_men_n1343_));
  NOi41      u1315(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1344_));
  NA3        u1316(.A(men_men_n1344_), .B(men_men_n872_), .C(men_men_n406_), .Y(men_men_n1345_));
  INV        u1317(.A(men_men_n1345_), .Y(men_men_n1346_));
  NA2        u1318(.A(men_men_n1087_), .B(men_men_n221_), .Y(men_men_n1347_));
  NO2        u1319(.A(men_men_n1347_), .B(men_men_n60_), .Y(men_men_n1348_));
  NO2        u1320(.A(k), .B(i), .Y(men_men_n1349_));
  NA2        u1321(.A(men_men_n88_), .B(men_men_n45_), .Y(men_men_n1350_));
  NO2        u1322(.A(men_men_n1053_), .B(men_men_n436_), .Y(men_men_n1351_));
  NA3        u1323(.A(men_men_n1351_), .B(men_men_n1350_), .C(men_men_n214_), .Y(men_men_n1352_));
  NO2        u1324(.A(men_men_n1063_), .B(men_men_n303_), .Y(men_men_n1353_));
  NA2        u1325(.A(men_men_n533_), .B(men_men_n81_), .Y(men_men_n1354_));
  NA2        u1326(.A(men_men_n1208_), .B(men_men_n286_), .Y(men_men_n1355_));
  NA3        u1327(.A(men_men_n1355_), .B(men_men_n1354_), .C(men_men_n1352_), .Y(men_men_n1356_));
  NO4        u1328(.A(men_men_n1356_), .B(men_men_n1348_), .C(men_men_n1346_), .D(men_men_n1343_), .Y(men_men_n1357_));
  NO3        u1329(.A(e), .B(d), .C(c), .Y(men_men_n1358_));
  OAI210     u1330(.A0(men_men_n134_), .A1(men_men_n214_), .B0(men_men_n601_), .Y(men_men_n1359_));
  NA2        u1331(.A(men_men_n1359_), .B(men_men_n1358_), .Y(men_men_n1360_));
  INV        u1332(.A(men_men_n1360_), .Y(men_men_n1361_));
  OR2        u1333(.A(h), .B(f), .Y(men_men_n1362_));
  NO3        u1334(.A(n), .B(m), .C(i), .Y(men_men_n1363_));
  OAI210     u1335(.A0(men_men_n1107_), .A1(men_men_n159_), .B0(men_men_n1363_), .Y(men_men_n1364_));
  NO2        u1336(.A(i), .B(g), .Y(men_men_n1365_));
  OR3        u1337(.A(men_men_n1365_), .B(men_men_n1337_), .C(men_men_n71_), .Y(men_men_n1366_));
  OAI220     u1338(.A0(men_men_n1366_), .A1(men_men_n472_), .B0(men_men_n1364_), .B1(men_men_n1362_), .Y(men_men_n1367_));
  NA3        u1339(.A(men_men_n692_), .B(men_men_n682_), .C(men_men_n114_), .Y(men_men_n1368_));
  NA3        u1340(.A(men_men_n1342_), .B(men_men_n1059_), .C(h), .Y(men_men_n1369_));
  AOI210     u1341(.A0(men_men_n1369_), .A1(men_men_n1368_), .B0(men_men_n45_), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n1363_), .B(men_men_n637_), .Y(men_men_n1371_));
  NO2        u1343(.A(l), .B(k), .Y(men_men_n1372_));
  NOi41      u1344(.An(men_men_n537_), .B(men_men_n1372_), .C(men_men_n467_), .D(men_men_n436_), .Y(men_men_n1373_));
  NO3        u1345(.A(men_men_n436_), .B(d), .C(c), .Y(men_men_n1374_));
  NO4        u1346(.A(men_men_n1373_), .B(men_men_n1370_), .C(men_men_n1367_), .D(men_men_n1361_), .Y(men_men_n1375_));
  NO2        u1347(.A(men_men_n150_), .B(h), .Y(men_men_n1376_));
  NO2        u1348(.A(men_men_n446_), .B(a), .Y(men_men_n1377_));
  NA3        u1349(.A(men_men_n1377_), .B(men_men_n1511_), .C(men_men_n115_), .Y(men_men_n1378_));
  NO2        u1350(.A(i), .B(h), .Y(men_men_n1379_));
  NA2        u1351(.A(men_men_n1379_), .B(men_men_n221_), .Y(men_men_n1380_));
  AOI210     u1352(.A0(men_men_n252_), .A1(men_men_n117_), .B0(men_men_n521_), .Y(men_men_n1381_));
  NO2        u1353(.A(men_men_n1381_), .B(men_men_n1380_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n751_), .B(men_men_n189_), .Y(men_men_n1383_));
  NOi31      u1355(.An(m), .B(n), .C(b), .Y(men_men_n1384_));
  NOi31      u1356(.An(f), .B(d), .C(c), .Y(men_men_n1385_));
  NA2        u1357(.A(men_men_n1385_), .B(men_men_n1384_), .Y(men_men_n1386_));
  INV        u1358(.A(men_men_n1386_), .Y(men_men_n1387_));
  NO3        u1359(.A(men_men_n1387_), .B(men_men_n1383_), .C(men_men_n1382_), .Y(men_men_n1388_));
  NO3        u1360(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1389_));
  AN2        u1361(.A(men_men_n1388_), .B(men_men_n1378_), .Y(men_men_n1390_));
  NA2        u1362(.A(men_men_n1342_), .B(men_men_n379_), .Y(men_men_n1391_));
  NO2        u1363(.A(men_men_n1391_), .B(men_men_n1045_), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n189_), .B(b), .Y(men_men_n1393_));
  NA2        u1365(.A(men_men_n1160_), .B(men_men_n1393_), .Y(men_men_n1394_));
  NO2        u1366(.A(i), .B(men_men_n213_), .Y(men_men_n1395_));
  NA4        u1367(.A(men_men_n1135_), .B(men_men_n1395_), .C(men_men_n106_), .D(m), .Y(men_men_n1396_));
  NAi31      u1368(.An(men_men_n1392_), .B(men_men_n1396_), .C(men_men_n1394_), .Y(men_men_n1397_));
  NA2        u1369(.A(men_men_n194_), .B(men_men_n100_), .Y(men_men_n1398_));
  OR2        u1370(.A(e), .B(a), .Y(men_men_n1399_));
  NOi41      u1371(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n1400_), .B(men_men_n115_), .Y(men_men_n1401_));
  INV        u1373(.A(men_men_n1401_), .Y(men_men_n1402_));
  OR3        u1374(.A(men_men_n532_), .B(men_men_n531_), .C(men_men_n114_), .Y(men_men_n1403_));
  NA2        u1375(.A(men_men_n1105_), .B(men_men_n403_), .Y(men_men_n1404_));
  OAI220     u1376(.A0(men_men_n1404_), .A1(men_men_n429_), .B0(men_men_n1403_), .B1(men_men_n296_), .Y(men_men_n1405_));
  AO210      u1377(.A0(men_men_n1405_), .A1(men_men_n117_), .B0(men_men_n1402_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1406_), .B(men_men_n1397_), .Y(men_men_n1407_));
  NA4        u1379(.A(men_men_n1407_), .B(men_men_n1390_), .C(men_men_n1375_), .D(men_men_n1357_), .Y(men_men_n1408_));
  NO2        u1380(.A(men_men_n1120_), .B(men_men_n112_), .Y(men_men_n1409_));
  NA2        u1381(.A(men_men_n379_), .B(men_men_n56_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1410_), .B(men_men_n1371_), .Y(men_men_n1411_));
  NA2        u1383(.A(men_men_n215_), .B(men_men_n181_), .Y(men_men_n1412_));
  AOI210     u1384(.A0(men_men_n1412_), .A1(men_men_n1180_), .B0(men_men_n1410_), .Y(men_men_n1413_));
  NO2        u1385(.A(men_men_n1080_), .B(men_men_n1077_), .Y(men_men_n1414_));
  NO3        u1386(.A(men_men_n1414_), .B(men_men_n1413_), .C(men_men_n1411_), .Y(men_men_n1415_));
  NA3        u1387(.A(men_men_n1389_), .B(men_men_n1341_), .C(men_men_n1105_), .Y(men_men_n1416_));
  NO3        u1388(.A(men_men_n1077_), .B(men_men_n575_), .C(g), .Y(men_men_n1417_));
  INV        u1389(.A(men_men_n1417_), .Y(men_men_n1418_));
  AOI210     u1390(.A0(men_men_n1418_), .A1(men_men_n1398_), .B0(men_men_n1053_), .Y(men_men_n1419_));
  INV        u1391(.A(men_men_n49_), .Y(men_men_n1420_));
  NA2        u1392(.A(men_men_n1420_), .B(men_men_n1168_), .Y(men_men_n1421_));
  INV        u1393(.A(men_men_n1421_), .Y(men_men_n1422_));
  OAI220     u1394(.A0(men_men_n665_), .A1(g), .B0(men_men_n224_), .B1(c), .Y(men_men_n1423_));
  AOI210     u1395(.A0(men_men_n1393_), .A1(men_men_n41_), .B0(men_men_n1423_), .Y(men_men_n1424_));
  NO2        u1396(.A(men_men_n134_), .B(l), .Y(men_men_n1425_));
  NO2        u1397(.A(men_men_n224_), .B(k), .Y(men_men_n1426_));
  OAI210     u1398(.A0(men_men_n1426_), .A1(men_men_n1379_), .B0(men_men_n1425_), .Y(men_men_n1427_));
  OAI220     u1399(.A0(men_men_n1427_), .A1(men_men_n31_), .B0(men_men_n1424_), .B1(men_men_n178_), .Y(men_men_n1428_));
  NO3        u1400(.A(men_men_n1403_), .B(men_men_n457_), .C(men_men_n350_), .Y(men_men_n1429_));
  NO4        u1401(.A(men_men_n1429_), .B(men_men_n1428_), .C(men_men_n1422_), .D(men_men_n1419_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n49_), .B(men_men_n575_), .Y(men_men_n1431_));
  NO3        u1403(.A(men_men_n1089_), .B(men_men_n1341_), .C(men_men_n49_), .Y(men_men_n1432_));
  NA2        u1404(.A(men_men_n1090_), .B(men_men_n1431_), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n1077_), .B(h), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1434_), .B(d), .C(men_men_n1046_), .Y(men_men_n1435_));
  OAI220     u1407(.A0(men_men_n1435_), .A1(c), .B0(men_men_n1433_), .B1(j), .Y(men_men_n1436_));
  NA3        u1408(.A(men_men_n1409_), .B(men_men_n457_), .C(f), .Y(men_men_n1437_));
  NO2        u1409(.A(men_men_n1336_), .B(men_men_n42_), .Y(men_men_n1438_));
  AOI210     u1410(.A0(men_men_n115_), .A1(men_men_n40_), .B0(men_men_n1438_), .Y(men_men_n1439_));
  NO2        u1411(.A(men_men_n1439_), .B(men_men_n1437_), .Y(men_men_n1440_));
  AOI210     u1412(.A0(men_men_n516_), .A1(h), .B0(men_men_n68_), .Y(men_men_n1441_));
  NA2        u1413(.A(men_men_n1441_), .B(men_men_n1377_), .Y(men_men_n1442_));
  NO2        u1414(.A(j), .B(men_men_n176_), .Y(men_men_n1443_));
  NOi21      u1415(.An(d), .B(f), .Y(men_men_n1444_));
  NO3        u1416(.A(men_men_n1385_), .B(men_men_n1444_), .C(men_men_n40_), .Y(men_men_n1445_));
  NA2        u1417(.A(men_men_n1445_), .B(men_men_n1443_), .Y(men_men_n1446_));
  NA2        u1418(.A(men_men_n1377_), .B(men_men_n1438_), .Y(men_men_n1447_));
  NO2        u1419(.A(men_men_n296_), .B(c), .Y(men_men_n1448_));
  NA2        u1420(.A(men_men_n1448_), .B(men_men_n533_), .Y(men_men_n1449_));
  NA4        u1421(.A(men_men_n1449_), .B(men_men_n1447_), .C(men_men_n1446_), .D(men_men_n1442_), .Y(men_men_n1450_));
  NO3        u1422(.A(men_men_n1450_), .B(men_men_n1440_), .C(men_men_n1436_), .Y(men_men_n1451_));
  NA4        u1423(.A(men_men_n1451_), .B(men_men_n1430_), .C(men_men_n1416_), .D(men_men_n1415_), .Y(men_men_n1452_));
  OAI220     u1424(.A0(men_men_n457_), .A1(men_men_n296_), .B0(men_men_n133_), .B1(men_men_n59_), .Y(men_men_n1453_));
  NA2        u1425(.A(men_men_n1453_), .B(men_men_n1353_), .Y(men_men_n1454_));
  INV        u1426(.A(men_men_n1454_), .Y(men_men_n1455_));
  NA3        u1427(.A(men_men_n1087_), .B(men_men_n110_), .C(men_men_n221_), .Y(men_men_n1456_));
  INV        u1428(.A(men_men_n1456_), .Y(men_men_n1457_));
  NO2        u1429(.A(men_men_n1457_), .B(men_men_n1455_), .Y(men_men_n1458_));
  NO2        u1430(.A(men_men_n1340_), .B(e), .Y(men_men_n1459_));
  NA2        u1431(.A(men_men_n1459_), .B(men_men_n401_), .Y(men_men_n1460_));
  OR3        u1432(.A(men_men_n1426_), .B(men_men_n1208_), .C(men_men_n134_), .Y(men_men_n1461_));
  NO2        u1433(.A(men_men_n1461_), .B(men_men_n1460_), .Y(men_men_n1462_));
  NO3        u1434(.A(men_men_n1403_), .B(men_men_n350_), .C(a), .Y(men_men_n1463_));
  NO2        u1435(.A(men_men_n1463_), .B(men_men_n1462_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n531_), .B(g), .Y(men_men_n1465_));
  AOI210     u1437(.A0(men_men_n1465_), .A1(men_men_n1374_), .B0(men_men_n1432_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n1399_), .B(f), .Y(men_men_n1467_));
  AOI210     u1439(.A0(men_men_n1115_), .A1(a), .B0(men_men_n1467_), .Y(men_men_n1468_));
  OAI220     u1440(.A0(men_men_n1468_), .A1(men_men_n68_), .B0(men_men_n1466_), .B1(men_men_n213_), .Y(men_men_n1469_));
  NA4        u1441(.A(men_men_n1087_), .B(men_men_n1084_), .C(men_men_n221_), .D(men_men_n67_), .Y(men_men_n1470_));
  NO2        u1442(.A(men_men_n49_), .B(l), .Y(men_men_n1471_));
  OAI210     u1443(.A0(men_men_n1399_), .A1(men_men_n864_), .B0(men_men_n472_), .Y(men_men_n1472_));
  OAI210     u1444(.A0(men_men_n1472_), .A1(men_men_n1090_), .B0(men_men_n1471_), .Y(men_men_n1473_));
  NO2        u1445(.A(men_men_n250_), .B(g), .Y(men_men_n1474_));
  NO2        u1446(.A(m), .B(i), .Y(men_men_n1475_));
  AOI220     u1447(.A0(men_men_n1475_), .A1(men_men_n1376_), .B0(men_men_n1069_), .B1(men_men_n1474_), .Y(men_men_n1476_));
  NA3        u1448(.A(men_men_n1476_), .B(men_men_n1473_), .C(men_men_n1470_), .Y(men_men_n1477_));
  NO2        u1449(.A(men_men_n1477_), .B(men_men_n1469_), .Y(men_men_n1478_));
  NA3        u1450(.A(men_men_n1478_), .B(men_men_n1464_), .C(men_men_n1458_), .Y(men_men_n1479_));
  NA3        u1451(.A(men_men_n964_), .B(men_men_n141_), .C(men_men_n46_), .Y(men_men_n1480_));
  AOI210     u1452(.A0(men_men_n151_), .A1(c), .B0(men_men_n1480_), .Y(men_men_n1481_));
  OAI210     u1453(.A0(men_men_n575_), .A1(g), .B0(men_men_n186_), .Y(men_men_n1482_));
  NA2        u1454(.A(men_men_n1482_), .B(men_men_n1434_), .Y(men_men_n1483_));
  NO2        u1455(.A(men_men_n71_), .B(c), .Y(men_men_n1484_));
  NO4        u1456(.A(men_men_n1362_), .B(men_men_n187_), .C(men_men_n443_), .D(men_men_n45_), .Y(men_men_n1485_));
  AOI210     u1457(.A0(men_men_n1443_), .A1(men_men_n1484_), .B0(men_men_n1485_), .Y(men_men_n1486_));
  NA2        u1458(.A(men_men_n1486_), .B(men_men_n1483_), .Y(men_men_n1487_));
  NO2        u1459(.A(men_men_n1487_), .B(men_men_n1481_), .Y(men_men_n1488_));
  NO4        u1460(.A(men_men_n224_), .B(men_men_n187_), .C(men_men_n252_), .D(k), .Y(men_men_n1489_));
  NO2        u1461(.A(men_men_n1480_), .B(men_men_n112_), .Y(men_men_n1490_));
  NO2        u1462(.A(men_men_n1490_), .B(men_men_n1489_), .Y(men_men_n1491_));
  AN2        u1463(.A(men_men_n1087_), .B(men_men_n1075_), .Y(men_men_n1492_));
  NA2        u1464(.A(men_men_n1512_), .B(men_men_n162_), .Y(men_men_n1493_));
  NOi31      u1465(.An(men_men_n30_), .B(men_men_n1493_), .C(n), .Y(men_men_n1494_));
  AOI210     u1466(.A0(men_men_n1492_), .A1(men_men_n1160_), .B0(men_men_n1494_), .Y(men_men_n1495_));
  NO2        u1467(.A(men_men_n1437_), .B(men_men_n68_), .Y(men_men_n1496_));
  NO2        u1468(.A(men_men_n1349_), .B(men_men_n119_), .Y(men_men_n1497_));
  NO2        u1469(.A(men_men_n1497_), .B(men_men_n1391_), .Y(men_men_n1498_));
  NO2        u1470(.A(men_men_n1498_), .B(men_men_n1496_), .Y(men_men_n1499_));
  NA4        u1471(.A(men_men_n1499_), .B(men_men_n1495_), .C(men_men_n1491_), .D(men_men_n1488_), .Y(men_men_n1500_));
  OR4        u1472(.A(men_men_n1500_), .B(men_men_n1479_), .C(men_men_n1452_), .D(men_men_n1408_), .Y(men04));
  NO4        u1473(.A(men_men_n268_), .B(men_men_n1039_), .C(men_men_n473_), .D(j), .Y(men_men_n1502_));
  OR2        u1474(.A(men_men_n1502_), .B(men_men_n1062_), .Y(men_men_n1503_));
  NO3        u1475(.A(men_men_n1350_), .B(men_men_n92_), .C(k), .Y(men_men_n1504_));
  NO2        u1476(.A(men_men_n1504_), .B(men_men_n1182_), .Y(men_men_n1505_));
  NA2        u1477(.A(men_men_n1505_), .B(men_men_n1212_), .Y(men_men_n1506_));
  NO4        u1478(.A(men_men_n1506_), .B(men_men_n1503_), .C(men_men_n1067_), .D(men_men_n1052_), .Y(men_men_n1507_));
  NA4        u1479(.A(men_men_n1507_), .B(men_men_n1117_), .C(men_men_n1103_), .D(men_men_n1091_), .Y(men05));
  INV        u1480(.A(i), .Y(men_men_n1511_));
  INV        u1481(.A(j), .Y(men_men_n1512_));
  INV        u1482(.A(men_men_n450_), .Y(men_men_n1513_));
  INV        u1483(.A(n), .Y(men_men_n1514_));
  INV        u1484(.A(n), .Y(men_men_n1515_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule