// Código templatep ara função duplica.
// Autor: Caio Vieira

module swap;
  // Substitua "?" pelos valores adequados
  parameter WIDTH = 3;

  reg [WIDTH-1:0] data_1;
  reg [WIDTH-1:0] data_2;
  
  // Escreva uma função duplica que recebe como entrada um vetor de tamanho
  // INP_WIDTH e retorna um outro vetor de tamanho OUT_WIDTH. O valor retornado
  //deve ser a entrada duplicada.
  task swap (input [WIDTH-1:0] d1, d2, output [WIDTH-1:0] s1, s2);
    begin
      	s1 = d2;
      	s2 = d1;
    end
  endtask
  
  initial begin
    integer i,j;
    for ( i = 0; i < 4'b1000; i = i+1) begin
      for ( j = 0; j < 4'b1000; j = j+1) begin
        $display("Before: data1: %0d | data2: %0d", i, j);
        swap(i,j,data_1,data_2);
        #1
        $display("After : data1: %0d | data2: %0d", data_1, data_2);
      end
    end
  end
  
endmodule

  
  