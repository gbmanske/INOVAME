library verilog;
use verilog.vl_types.all;
entity tb_sad is
end tb_sad;
