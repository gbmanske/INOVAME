// Benchmark "top" written by ABC on Thu Jun 20 14:59:19 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n142_, new_new_n143_,
    new_new_n144_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1012_, new_new_n1013_, new_new_n1014_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g040(.A(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g063(.A(i_6_), .Y(new_new_n86_));
  OR4        g064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n88_), .B(new_new_n89_), .Y(new_new_n90_));
  OAI210     g068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g073(.A(new_new_n95_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n98_));
  AN3        g076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g080(.A0(new_new_n102_), .A1(new_new_n62_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g081(.A(i_7_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n46_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(new_new_n86_), .Y(new_new_n107_));
  NA2        g085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  NO3        g089(.A(new_new_n111_), .B(new_new_n92_), .C(new_new_n53_), .Y(new_new_n112_));
  AN2        g090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g092(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n115_));
  NO2        g093(.A(i_8_), .B(new_new_n104_), .Y(new_new_n116_));
  NO3        g094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_0_), .Y(new_new_n120_));
  NA2        g098(.A(i_11_), .B(i_12_), .Y(new_new_n121_));
  OAI210     g099(.A0(new_new_n120_), .A1(new_new_n118_), .B0(new_new_n121_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n122_), .B(new_new_n117_), .Y(new_new_n123_));
  NAi41      g101(.An(new_new_n112_), .B(new_new_n123_), .C(new_new_n110_), .D(new_new_n103_), .Y(new_new_n124_));
  NOi21      g102(.An(i_1_), .B(i_5_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(i_11_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g105(.A(i_7_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NO2        g107(.A(new_new_n129_), .B(new_new_n46_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n131_));
  NAi21      g109(.An(i_3_), .B(i_8_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n132_), .B(new_new_n62_), .Y(new_new_n133_));
  NOi31      g111(.An(new_new_n133_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n134_));
  NO2        g112(.A(i_1_), .B(new_new_n86_), .Y(new_new_n135_));
  NO2        g113(.A(i_6_), .B(i_5_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_3_), .Y(new_new_n137_));
  AO210      g115(.A0(new_new_n137_), .A1(new_new_n47_), .B0(new_new_n135_), .Y(new_new_n138_));
  OAI220     g116(.A0(new_new_n138_), .A1(new_new_n111_), .B0(new_new_n134_), .B1(new_new_n126_), .Y(new_new_n139_));
  NO3        g117(.A(new_new_n139_), .B(new_new_n124_), .C(new_new_n98_), .Y(new_new_n140_));
  NA3        g118(.A(new_new_n140_), .B(new_new_n79_), .C(new_new_n56_), .Y(ori2));
  NO2        g119(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n142_));
  NA2        g120(.A(i_6_), .B(new_new_n25_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NA4        g122(.A(new_new_n144_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(ori0));
  AN2        g123(.A(i_8_), .B(i_7_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(i_6_), .Y(new_new_n147_));
  NO2        g125(.A(i_12_), .B(i_13_), .Y(new_new_n148_));
  NAi21      g126(.An(i_5_), .B(i_11_), .Y(new_new_n149_));
  NOi21      g127(.An(new_new_n148_), .B(new_new_n149_), .Y(new_new_n150_));
  NO2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NA2        g129(.A(i_2_), .B(i_3_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n152_), .B(i_4_), .Y(new_new_n153_));
  NA3        g131(.A(new_new_n153_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n154_));
  OR2        g132(.A(new_new_n154_), .B(new_new_n25_), .Y(new_new_n155_));
  AN2        g133(.A(new_new_n148_), .B(new_new_n83_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n156_), .B(new_new_n27_), .Y(new_new_n157_));
  NA2        g135(.A(i_1_), .B(i_5_), .Y(new_new_n158_));
  NO2        g136(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n159_), .B(new_new_n36_), .Y(new_new_n160_));
  NO3        g138(.A(new_new_n160_), .B(new_new_n158_), .C(new_new_n157_), .Y(new_new_n161_));
  OR2        g139(.A(i_0_), .B(i_1_), .Y(new_new_n162_));
  NO3        g140(.A(new_new_n162_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n163_));
  NAi32      g141(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n164_));
  NAi21      g142(.An(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  NOi21      g143(.An(i_4_), .B(i_10_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(new_new_n40_), .Y(new_new_n167_));
  NO2        g145(.A(i_3_), .B(i_5_), .Y(new_new_n168_));
  NO3        g146(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n169_));
  NA2        g147(.A(new_new_n169_), .B(new_new_n168_), .Y(new_new_n170_));
  OAI210     g148(.A0(new_new_n170_), .A1(new_new_n167_), .B0(new_new_n165_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n171_), .B(new_new_n161_), .Y(new_new_n172_));
  AOI210     g150(.A0(new_new_n172_), .A1(new_new_n155_), .B0(new_new_n147_), .Y(new_new_n173_));
  NA2        g151(.A(i_3_), .B(new_new_n48_), .Y(new_new_n174_));
  NOi21      g152(.An(i_4_), .B(i_9_), .Y(new_new_n175_));
  NOi21      g153(.An(i_11_), .B(i_13_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n176_), .B(new_new_n175_), .Y(new_new_n177_));
  NO2        g155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n83_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(new_new_n46_), .Y(new_new_n183_));
  NA2        g161(.A(new_new_n36_), .B(i_5_), .Y(new_new_n184_));
  NAi31      g162(.An(new_new_n184_), .B(new_new_n156_), .C(i_11_), .Y(new_new_n185_));
  NA2        g163(.A(i_3_), .B(i_5_), .Y(new_new_n186_));
  OR2        g164(.A(new_new_n186_), .B(new_new_n177_), .Y(new_new_n187_));
  AOI210     g165(.A0(new_new_n187_), .A1(new_new_n185_), .B0(new_new_n183_), .Y(new_new_n188_));
  NO2        g166(.A(new_new_n73_), .B(i_5_), .Y(new_new_n189_));
  NO2        g167(.A(i_13_), .B(i_10_), .Y(new_new_n190_));
  NO2        g168(.A(i_2_), .B(i_1_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(i_3_), .Y(new_new_n192_));
  NAi21      g170(.An(i_4_), .B(i_12_), .Y(new_new_n193_));
  INV        g171(.A(new_new_n188_), .Y(new_new_n194_));
  INV        g172(.A(i_8_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n195_), .B(i_7_), .Y(new_new_n196_));
  NA2        g174(.A(new_new_n196_), .B(i_6_), .Y(new_new_n197_));
  NO3        g175(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n198_));
  NA2        g176(.A(new_new_n198_), .B(new_new_n116_), .Y(new_new_n199_));
  NO3        g177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n200_));
  NA3        g178(.A(new_new_n200_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n201_));
  NO3        g179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n202_));
  OAI210     g180(.A0(new_new_n99_), .A1(i_12_), .B0(new_new_n202_), .Y(new_new_n203_));
  AOI210     g181(.A0(new_new_n203_), .A1(new_new_n201_), .B0(new_new_n199_), .Y(new_new_n204_));
  NO2        g182(.A(i_3_), .B(i_8_), .Y(new_new_n205_));
  NO3        g183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n206_));
  NA3        g184(.A(new_new_n206_), .B(new_new_n205_), .C(new_new_n40_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n106_), .B(new_new_n58_), .Y(new_new_n208_));
  INV        g186(.A(new_new_n208_), .Y(new_new_n209_));
  NO2        g187(.A(i_13_), .B(i_9_), .Y(new_new_n210_));
  NAi21      g188(.An(i_12_), .B(i_3_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n44_), .B(i_5_), .Y(new_new_n212_));
  NO3        g190(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n209_), .B(new_new_n207_), .Y(new_new_n214_));
  AOI210     g192(.A0(new_new_n214_), .A1(i_7_), .B0(new_new_n204_), .Y(new_new_n215_));
  OAI220     g193(.A0(new_new_n215_), .A1(i_4_), .B0(new_new_n197_), .B1(new_new_n194_), .Y(new_new_n216_));
  NAi21      g194(.An(i_12_), .B(i_7_), .Y(new_new_n217_));
  NA3        g195(.A(i_13_), .B(new_new_n195_), .C(i_10_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  NA2        g197(.A(i_0_), .B(i_5_), .Y(new_new_n220_));
  NA2        g198(.A(new_new_n220_), .B(new_new_n107_), .Y(new_new_n221_));
  OAI220     g199(.A0(new_new_n221_), .A1(new_new_n192_), .B0(new_new_n183_), .B1(new_new_n137_), .Y(new_new_n222_));
  NAi31      g200(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n36_), .B(i_13_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n226_));
  NA3        g204(.A(new_new_n226_), .B(new_new_n225_), .C(new_new_n224_), .Y(new_new_n227_));
  INV        g205(.A(i_13_), .Y(new_new_n228_));
  NO2        g206(.A(i_12_), .B(new_new_n228_), .Y(new_new_n229_));
  NA3        g207(.A(new_new_n229_), .B(new_new_n200_), .C(new_new_n198_), .Y(new_new_n230_));
  OAI210     g208(.A0(new_new_n227_), .A1(new_new_n223_), .B0(new_new_n230_), .Y(new_new_n231_));
  AOI220     g209(.A0(new_new_n231_), .A1(new_new_n146_), .B0(new_new_n222_), .B1(new_new_n219_), .Y(new_new_n232_));
  NO2        g210(.A(i_12_), .B(new_new_n37_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n186_), .B(i_4_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n234_), .B(new_new_n233_), .Y(new_new_n235_));
  OR2        g213(.A(i_8_), .B(i_7_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n236_), .B(new_new_n86_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n53_), .B(i_1_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n237_), .Y(new_new_n239_));
  INV        g217(.A(i_12_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n44_), .B(new_new_n240_), .Y(new_new_n241_));
  NO3        g219(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n242_));
  NA2        g220(.A(i_2_), .B(i_1_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n239_), .B(new_new_n235_), .Y(new_new_n244_));
  NO3        g222(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n245_));
  NAi21      g223(.An(i_4_), .B(i_3_), .Y(new_new_n246_));
  NO2        g224(.A(new_new_n246_), .B(new_new_n75_), .Y(new_new_n247_));
  NO2        g225(.A(i_0_), .B(i_6_), .Y(new_new_n248_));
  NOi41      g226(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n249_), .B(new_new_n248_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n243_), .B(new_new_n186_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n244_), .B(new_new_n210_), .Y(new_new_n252_));
  NO2        g230(.A(i_11_), .B(new_new_n228_), .Y(new_new_n253_));
  NOi21      g231(.An(i_1_), .B(i_6_), .Y(new_new_n254_));
  NAi21      g232(.An(i_3_), .B(i_7_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n240_), .B(i_9_), .Y(new_new_n256_));
  OR4        g234(.A(new_new_n256_), .B(new_new_n255_), .C(new_new_n254_), .D(new_new_n189_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n258_));
  NO2        g236(.A(i_12_), .B(i_3_), .Y(new_new_n259_));
  NA2        g237(.A(new_new_n73_), .B(i_5_), .Y(new_new_n260_));
  NA2        g238(.A(i_3_), .B(i_9_), .Y(new_new_n261_));
  NAi21      g239(.An(i_7_), .B(i_10_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n262_), .B(new_new_n261_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n263_), .B(new_new_n260_), .C(new_new_n64_), .Y(new_new_n264_));
  NA2        g242(.A(new_new_n264_), .B(new_new_n257_), .Y(new_new_n265_));
  NA3        g243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n266_));
  INV        g244(.A(new_new_n147_), .Y(new_new_n267_));
  NA2        g245(.A(new_new_n240_), .B(i_13_), .Y(new_new_n268_));
  NO2        g246(.A(new_new_n268_), .B(new_new_n75_), .Y(new_new_n269_));
  AOI220     g247(.A0(new_new_n269_), .A1(new_new_n267_), .B0(new_new_n265_), .B1(new_new_n253_), .Y(new_new_n270_));
  NO2        g248(.A(new_new_n236_), .B(new_new_n37_), .Y(new_new_n271_));
  NA2        g249(.A(i_12_), .B(i_6_), .Y(new_new_n272_));
  OR2        g250(.A(i_13_), .B(i_9_), .Y(new_new_n273_));
  NO3        g251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n48_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n246_), .B(i_2_), .Y(new_new_n275_));
  NA3        g253(.A(new_new_n275_), .B(new_new_n274_), .C(new_new_n44_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n253_), .B(i_9_), .Y(new_new_n277_));
  NA2        g255(.A(new_new_n260_), .B(new_new_n64_), .Y(new_new_n278_));
  OAI210     g256(.A0(new_new_n278_), .A1(new_new_n277_), .B0(new_new_n276_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n159_), .B(new_new_n63_), .Y(new_new_n280_));
  NO3        g258(.A(i_11_), .B(new_new_n228_), .C(new_new_n25_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n255_), .B(i_8_), .Y(new_new_n282_));
  NO2        g260(.A(i_6_), .B(new_new_n48_), .Y(new_new_n283_));
  NA3        g261(.A(new_new_n283_), .B(new_new_n282_), .C(new_new_n281_), .Y(new_new_n284_));
  NO3        g262(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n285_));
  NA3        g263(.A(new_new_n285_), .B(new_new_n271_), .C(new_new_n229_), .Y(new_new_n286_));
  AOI210     g264(.A0(new_new_n286_), .A1(new_new_n284_), .B0(new_new_n280_), .Y(new_new_n287_));
  AOI210     g265(.A0(new_new_n279_), .A1(new_new_n271_), .B0(new_new_n287_), .Y(new_new_n288_));
  NA4        g266(.A(new_new_n288_), .B(new_new_n270_), .C(new_new_n252_), .D(new_new_n232_), .Y(new_new_n289_));
  NO3        g267(.A(i_12_), .B(new_new_n228_), .C(new_new_n37_), .Y(new_new_n290_));
  INV        g268(.A(new_new_n290_), .Y(new_new_n291_));
  NA2        g269(.A(i_8_), .B(new_new_n104_), .Y(new_new_n292_));
  NOi21      g270(.An(new_new_n168_), .B(new_new_n86_), .Y(new_new_n293_));
  NO3        g271(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n294_));
  AOI220     g272(.A0(new_new_n294_), .A1(new_new_n198_), .B0(new_new_n293_), .B1(new_new_n238_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n295_), .B(new_new_n292_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n243_), .B(i_0_), .Y(new_new_n297_));
  NA2        g275(.A(i_0_), .B(i_1_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n298_), .B(i_2_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n59_), .B(i_6_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n170_), .B(new_new_n147_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(new_new_n296_), .Y(new_new_n302_));
  NO2        g280(.A(i_3_), .B(i_10_), .Y(new_new_n303_));
  NA3        g281(.A(new_new_n303_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n304_));
  NO2        g282(.A(i_2_), .B(new_new_n104_), .Y(new_new_n305_));
  NA2        g283(.A(i_1_), .B(new_new_n36_), .Y(new_new_n306_));
  AN2        g284(.A(i_3_), .B(i_10_), .Y(new_new_n307_));
  NA4        g285(.A(new_new_n307_), .B(new_new_n200_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n308_));
  NO2        g286(.A(i_5_), .B(new_new_n37_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n302_), .B(new_new_n291_), .Y(new_new_n311_));
  NO4        g289(.A(new_new_n311_), .B(new_new_n289_), .C(new_new_n216_), .D(new_new_n173_), .Y(new_new_n312_));
  NO3        g290(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n314_));
  NO3        g292(.A(i_6_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n315_));
  NO2        g293(.A(i_2_), .B(i_3_), .Y(new_new_n316_));
  OR2        g294(.A(i_0_), .B(i_5_), .Y(new_new_n317_));
  NA2        g295(.A(new_new_n220_), .B(new_new_n317_), .Y(new_new_n318_));
  NA4        g296(.A(new_new_n318_), .B(new_new_n237_), .C(new_new_n316_), .D(i_1_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n297_), .B(new_new_n293_), .C(new_new_n116_), .Y(new_new_n320_));
  NAi21      g298(.An(i_8_), .B(i_7_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n321_), .B(i_6_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n162_), .B(new_new_n46_), .Y(new_new_n323_));
  NA3        g301(.A(new_new_n323_), .B(new_new_n322_), .C(new_new_n168_), .Y(new_new_n324_));
  NA3        g302(.A(new_new_n324_), .B(new_new_n320_), .C(new_new_n319_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n325_), .B(i_4_), .Y(new_new_n326_));
  NO2        g304(.A(i_12_), .B(i_10_), .Y(new_new_n327_));
  NOi21      g305(.An(i_5_), .B(i_0_), .Y(new_new_n328_));
  NA4        g306(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n329_));
  NO2        g307(.A(i_6_), .B(i_8_), .Y(new_new_n330_));
  NOi21      g308(.An(i_0_), .B(i_2_), .Y(new_new_n331_));
  AN2        g309(.A(new_new_n331_), .B(new_new_n330_), .Y(new_new_n332_));
  NO2        g310(.A(i_1_), .B(i_7_), .Y(new_new_n333_));
  INV        g311(.A(new_new_n326_), .Y(new_new_n334_));
  NO3        g312(.A(new_new_n236_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n335_));
  NO3        g313(.A(new_new_n321_), .B(i_2_), .C(i_1_), .Y(new_new_n336_));
  OAI210     g314(.A0(new_new_n336_), .A1(new_new_n335_), .B0(i_6_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n254_), .B(new_new_n305_), .C(new_new_n195_), .Y(new_new_n338_));
  AOI210     g316(.A0(new_new_n338_), .A1(new_new_n337_), .B0(new_new_n318_), .Y(new_new_n339_));
  NOi21      g317(.An(new_new_n158_), .B(new_new_n107_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n340_), .B(new_new_n128_), .Y(new_new_n341_));
  OAI210     g319(.A0(new_new_n341_), .A1(new_new_n339_), .B0(i_3_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n298_), .B(new_new_n81_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n343_), .B(new_new_n136_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n344_), .B(i_3_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n195_), .B(i_9_), .Y(new_new_n346_));
  NA2        g324(.A(new_new_n346_), .B(new_new_n208_), .Y(new_new_n347_));
  NO2        g325(.A(new_new_n347_), .B(new_new_n46_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n345_), .Y(new_new_n349_));
  AOI210     g327(.A0(new_new_n349_), .A1(new_new_n342_), .B0(new_new_n167_), .Y(new_new_n350_));
  AOI210     g328(.A0(new_new_n334_), .A1(new_new_n313_), .B0(new_new_n350_), .Y(new_new_n351_));
  NOi32      g329(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n352_));
  INV        g330(.A(new_new_n352_), .Y(new_new_n353_));
  NAi21      g331(.An(i_0_), .B(i_6_), .Y(new_new_n354_));
  NAi21      g332(.An(i_1_), .B(i_5_), .Y(new_new_n355_));
  NA2        g333(.A(new_new_n355_), .B(new_new_n354_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n356_), .B(new_new_n25_), .Y(new_new_n357_));
  OAI210     g335(.A0(new_new_n357_), .A1(new_new_n164_), .B0(new_new_n250_), .Y(new_new_n358_));
  NAi41      g336(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n359_));
  OAI220     g337(.A0(new_new_n359_), .A1(new_new_n355_), .B0(new_new_n223_), .B1(new_new_n164_), .Y(new_new_n360_));
  AOI210     g338(.A0(new_new_n359_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n361_));
  NOi32      g339(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n362_));
  NAi21      g340(.An(i_6_), .B(i_1_), .Y(new_new_n363_));
  OR2        g341(.A(new_new_n361_), .B(new_new_n360_), .Y(new_new_n364_));
  NO2        g342(.A(i_1_), .B(new_new_n104_), .Y(new_new_n365_));
  NAi21      g343(.An(i_3_), .B(i_4_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n366_), .B(i_9_), .Y(new_new_n367_));
  AN2        g345(.A(i_6_), .B(i_7_), .Y(new_new_n368_));
  OAI210     g346(.A0(new_new_n368_), .A1(new_new_n365_), .B0(new_new_n367_), .Y(new_new_n369_));
  NA2        g347(.A(i_2_), .B(i_7_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n366_), .B(i_10_), .Y(new_new_n371_));
  NA3        g349(.A(new_new_n371_), .B(new_new_n370_), .C(new_new_n248_), .Y(new_new_n372_));
  AOI210     g350(.A0(new_new_n372_), .A1(new_new_n369_), .B0(new_new_n189_), .Y(new_new_n373_));
  AOI210     g351(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n374_));
  OAI210     g352(.A0(new_new_n374_), .A1(new_new_n191_), .B0(new_new_n371_), .Y(new_new_n375_));
  AOI220     g353(.A0(new_new_n371_), .A1(new_new_n333_), .B0(new_new_n242_), .B1(new_new_n191_), .Y(new_new_n376_));
  AOI210     g354(.A0(new_new_n376_), .A1(new_new_n375_), .B0(i_5_), .Y(new_new_n377_));
  NO4        g355(.A(new_new_n377_), .B(new_new_n373_), .C(new_new_n364_), .D(new_new_n358_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(new_new_n353_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n380_));
  AN2        g358(.A(i_12_), .B(i_5_), .Y(new_new_n381_));
  NO2        g359(.A(i_4_), .B(new_new_n26_), .Y(new_new_n382_));
  NO2        g360(.A(i_11_), .B(i_6_), .Y(new_new_n383_));
  NO2        g361(.A(i_5_), .B(i_10_), .Y(new_new_n384_));
  NO2        g362(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n154_), .B(new_new_n86_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  NO3        g365(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n388_));
  NO2        g366(.A(i_3_), .B(new_new_n104_), .Y(new_new_n389_));
  NO2        g367(.A(i_11_), .B(i_12_), .Y(new_new_n390_));
  NAi21      g368(.An(i_13_), .B(i_0_), .Y(new_new_n391_));
  INV        g369(.A(new_new_n387_), .Y(new_new_n392_));
  NO3        g370(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n393_));
  NO2        g371(.A(i_0_), .B(i_11_), .Y(new_new_n394_));
  INV        g372(.A(i_5_), .Y(new_new_n395_));
  AN2        g373(.A(i_1_), .B(i_6_), .Y(new_new_n396_));
  NOi21      g374(.An(i_2_), .B(i_12_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n397_), .B(new_new_n396_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n395_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n146_), .B(i_9_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n400_), .B(i_4_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n399_), .B(new_new_n401_), .Y(new_new_n402_));
  NAi21      g380(.An(i_9_), .B(i_4_), .Y(new_new_n403_));
  OR2        g381(.A(i_13_), .B(i_10_), .Y(new_new_n404_));
  NO3        g382(.A(new_new_n404_), .B(new_new_n121_), .C(new_new_n403_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n177_), .B(new_new_n127_), .Y(new_new_n406_));
  OR2        g384(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n290_), .B(new_new_n408_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n283_), .B(new_new_n213_), .Y(new_new_n410_));
  OAI220     g388(.A0(new_new_n410_), .A1(new_new_n407_), .B0(new_new_n409_), .B1(new_new_n340_), .Y(new_new_n411_));
  INV        g389(.A(new_new_n411_), .Y(new_new_n412_));
  AOI210     g390(.A0(new_new_n412_), .A1(new_new_n402_), .B0(new_new_n26_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n320_), .B(new_new_n319_), .Y(new_new_n414_));
  AOI220     g392(.A0(new_new_n300_), .A1(new_new_n294_), .B0(new_new_n297_), .B1(new_new_n314_), .Y(new_new_n415_));
  NO2        g393(.A(new_new_n415_), .B(new_new_n174_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n186_), .B(new_new_n86_), .Y(new_new_n417_));
  AOI220     g395(.A0(new_new_n417_), .A1(new_new_n299_), .B0(new_new_n285_), .B1(new_new_n213_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n418_), .B(new_new_n292_), .Y(new_new_n419_));
  NO3        g397(.A(new_new_n419_), .B(new_new_n416_), .C(new_new_n414_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n198_), .B(new_new_n99_), .Y(new_new_n421_));
  NA3        g399(.A(new_new_n323_), .B(new_new_n168_), .C(new_new_n86_), .Y(new_new_n422_));
  AOI210     g400(.A0(new_new_n422_), .A1(new_new_n421_), .B0(new_new_n321_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n195_), .B(i_10_), .Y(new_new_n424_));
  NA3        g402(.A(new_new_n260_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n425_));
  NA2        g403(.A(new_new_n300_), .B(new_new_n238_), .Y(new_new_n426_));
  OAI220     g404(.A0(new_new_n426_), .A1(new_new_n186_), .B0(new_new_n425_), .B1(new_new_n424_), .Y(new_new_n427_));
  NO2        g405(.A(new_new_n427_), .B(new_new_n423_), .Y(new_new_n428_));
  AOI210     g406(.A0(new_new_n428_), .A1(new_new_n420_), .B0(new_new_n277_), .Y(new_new_n429_));
  NO4        g407(.A(new_new_n429_), .B(new_new_n413_), .C(new_new_n392_), .D(new_new_n379_), .Y(new_new_n430_));
  NO2        g408(.A(new_new_n63_), .B(i_4_), .Y(new_new_n431_));
  NO2        g409(.A(new_new_n73_), .B(i_13_), .Y(new_new_n432_));
  NA3        g410(.A(new_new_n432_), .B(new_new_n431_), .C(i_2_), .Y(new_new_n433_));
  NO2        g411(.A(i_10_), .B(i_9_), .Y(new_new_n434_));
  NAi21      g412(.An(i_12_), .B(i_8_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n435_), .B(i_3_), .Y(new_new_n436_));
  NA2        g414(.A(new_new_n436_), .B(new_new_n434_), .Y(new_new_n437_));
  NO2        g415(.A(new_new_n46_), .B(i_4_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(new_new_n107_), .Y(new_new_n439_));
  OAI220     g417(.A0(new_new_n439_), .A1(new_new_n207_), .B0(new_new_n437_), .B1(new_new_n433_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n310_), .B(i_0_), .Y(new_new_n441_));
  NO3        g419(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n272_), .B(new_new_n100_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n443_), .B(new_new_n442_), .Y(new_new_n444_));
  NA2        g422(.A(i_8_), .B(i_9_), .Y(new_new_n445_));
  AOI210     g423(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n446_));
  OR2        g424(.A(new_new_n446_), .B(new_new_n445_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n290_), .B(new_new_n208_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n448_), .B(new_new_n447_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n253_), .B(new_new_n309_), .Y(new_new_n450_));
  NO3        g428(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n451_));
  INV        g429(.A(new_new_n451_), .Y(new_new_n452_));
  NA3        g430(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n453_));
  NA4        g431(.A(new_new_n149_), .B(new_new_n119_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n454_));
  OAI220     g432(.A0(new_new_n454_), .A1(new_new_n453_), .B0(new_new_n452_), .B1(new_new_n450_), .Y(new_new_n455_));
  NO3        g433(.A(new_new_n455_), .B(new_new_n449_), .C(new_new_n440_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n99_), .B(i_13_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n417_), .B(new_new_n380_), .Y(new_new_n458_));
  NO2        g436(.A(i_2_), .B(i_13_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n458_), .B(new_new_n457_), .Y(new_new_n460_));
  NO3        g438(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n461_));
  NO2        g439(.A(i_6_), .B(i_7_), .Y(new_new_n462_));
  NO2        g440(.A(i_11_), .B(i_1_), .Y(new_new_n463_));
  NOi21      g441(.An(i_2_), .B(i_7_), .Y(new_new_n464_));
  NO2        g442(.A(i_3_), .B(new_new_n195_), .Y(new_new_n465_));
  NO2        g443(.A(i_6_), .B(i_10_), .Y(new_new_n466_));
  NA4        g444(.A(new_new_n466_), .B(new_new_n313_), .C(new_new_n465_), .D(new_new_n240_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n467_), .B(new_new_n160_), .Y(new_new_n468_));
  NA3        g446(.A(new_new_n249_), .B(new_new_n176_), .C(new_new_n136_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n162_), .B(i_3_), .Y(new_new_n471_));
  NAi31      g449(.An(new_new_n470_), .B(new_new_n471_), .C(new_new_n229_), .Y(new_new_n472_));
  NA3        g450(.A(new_new_n385_), .B(new_new_n182_), .C(new_new_n153_), .Y(new_new_n473_));
  NA3        g451(.A(new_new_n473_), .B(new_new_n472_), .C(new_new_n469_), .Y(new_new_n474_));
  NO3        g452(.A(new_new_n474_), .B(new_new_n468_), .C(new_new_n460_), .Y(new_new_n475_));
  NA2        g453(.A(new_new_n442_), .B(new_new_n381_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n451_), .B(new_new_n384_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n477_), .B(new_new_n227_), .Y(new_new_n478_));
  NAi21      g456(.An(new_new_n218_), .B(new_new_n390_), .Y(new_new_n479_));
  NA2        g457(.A(new_new_n333_), .B(new_new_n220_), .Y(new_new_n480_));
  NO2        g458(.A(new_new_n26_), .B(i_5_), .Y(new_new_n481_));
  NO2        g459(.A(i_0_), .B(new_new_n86_), .Y(new_new_n482_));
  NA3        g460(.A(new_new_n482_), .B(new_new_n481_), .C(new_new_n146_), .Y(new_new_n483_));
  OR3        g461(.A(new_new_n306_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n484_));
  OAI220     g462(.A0(new_new_n484_), .A1(new_new_n483_), .B0(new_new_n480_), .B1(new_new_n479_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n27_), .B(i_10_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n313_), .B(new_new_n242_), .Y(new_new_n487_));
  OAI220     g465(.A0(new_new_n487_), .A1(new_new_n425_), .B0(new_new_n486_), .B1(new_new_n457_), .Y(new_new_n488_));
  NO3        g466(.A(new_new_n488_), .B(new_new_n485_), .C(new_new_n478_), .Y(new_new_n489_));
  NA3        g467(.A(new_new_n489_), .B(new_new_n475_), .C(new_new_n456_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n126_), .B(new_new_n115_), .Y(new_new_n491_));
  AN2        g469(.A(new_new_n491_), .B(new_new_n442_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n313_), .B(new_new_n169_), .Y(new_new_n493_));
  OAI210     g471(.A0(new_new_n493_), .A1(new_new_n235_), .B0(new_new_n308_), .Y(new_new_n494_));
  AOI220     g472(.A0(new_new_n494_), .A1(new_new_n322_), .B0(new_new_n492_), .B1(new_new_n310_), .Y(new_new_n495_));
  NA4        g473(.A(new_new_n432_), .B(new_new_n431_), .C(new_new_n205_), .D(i_2_), .Y(new_new_n496_));
  INV        g474(.A(new_new_n496_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n381_), .B(new_new_n228_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n368_), .B(new_new_n362_), .Y(new_new_n499_));
  OR2        g477(.A(new_new_n498_), .B(new_new_n499_), .Y(new_new_n500_));
  NO2        g478(.A(new_new_n36_), .B(i_8_), .Y(new_new_n501_));
  AOI210     g479(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n405_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n502_), .B(new_new_n500_), .Y(new_new_n503_));
  AOI210     g481(.A0(new_new_n497_), .A1(new_new_n206_), .B0(new_new_n503_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n260_), .B(new_new_n64_), .Y(new_new_n505_));
  OAI210     g483(.A0(i_8_), .A1(new_new_n505_), .B0(new_new_n138_), .Y(new_new_n506_));
  AOI210     g484(.A0(new_new_n196_), .A1(i_9_), .B0(new_new_n271_), .Y(new_new_n507_));
  NO2        g485(.A(new_new_n507_), .B(new_new_n201_), .Y(new_new_n508_));
  OR2        g486(.A(new_new_n186_), .B(i_4_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n509_), .B(new_new_n86_), .Y(new_new_n510_));
  AOI220     g488(.A0(new_new_n510_), .A1(new_new_n508_), .B0(new_new_n506_), .B1(new_new_n406_), .Y(new_new_n511_));
  NA3        g489(.A(new_new_n511_), .B(new_new_n504_), .C(new_new_n495_), .Y(new_new_n512_));
  NO2        g490(.A(i_12_), .B(new_new_n195_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n513_), .B(new_new_n228_), .Y(new_new_n514_));
  NO2        g492(.A(i_8_), .B(i_7_), .Y(new_new_n515_));
  OAI210     g493(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n516_), .B(new_new_n226_), .Y(new_new_n517_));
  AOI220     g495(.A0(new_new_n323_), .A1(new_new_n40_), .B0(new_new_n238_), .B1(new_new_n210_), .Y(new_new_n518_));
  OAI220     g496(.A0(new_new_n518_), .A1(new_new_n509_), .B0(new_new_n517_), .B1(new_new_n246_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n44_), .B(i_10_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n520_), .B(i_6_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n521_), .B(new_new_n519_), .C(new_new_n515_), .Y(new_new_n522_));
  AOI220     g500(.A0(new_new_n417_), .A1(new_new_n323_), .B0(new_new_n251_), .B1(new_new_n248_), .Y(new_new_n523_));
  OAI220     g501(.A0(new_new_n523_), .A1(new_new_n268_), .B0(new_new_n457_), .B1(new_new_n137_), .Y(new_new_n524_));
  NA2        g502(.A(new_new_n524_), .B(new_new_n271_), .Y(new_new_n525_));
  NOi31      g503(.An(new_new_n297_), .B(new_new_n304_), .C(new_new_n184_), .Y(new_new_n526_));
  NA3        g504(.A(new_new_n307_), .B(new_new_n178_), .C(new_new_n99_), .Y(new_new_n527_));
  OAI210     g505(.A0(new_new_n1013_), .A1(new_new_n526_), .B0(new_new_n451_), .Y(new_new_n528_));
  NA3        g506(.A(new_new_n528_), .B(new_new_n525_), .C(new_new_n522_), .Y(new_new_n529_));
  NA3        g507(.A(new_new_n220_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n530_));
  NA2        g508(.A(new_new_n290_), .B(new_new_n84_), .Y(new_new_n531_));
  AOI210     g509(.A0(new_new_n530_), .A1(new_new_n344_), .B0(new_new_n531_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n226_), .B(new_new_n225_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n434_), .B(new_new_n224_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n533_), .B(new_new_n534_), .Y(new_new_n535_));
  AOI210     g513(.A0(new_new_n363_), .A1(new_new_n46_), .B0(new_new_n365_), .Y(new_new_n536_));
  NA2        g514(.A(i_0_), .B(new_new_n48_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n513_), .B(new_new_n281_), .C(new_new_n537_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n536_), .B(new_new_n538_), .Y(new_new_n539_));
  NO3        g517(.A(new_new_n539_), .B(new_new_n535_), .C(new_new_n532_), .Y(new_new_n540_));
  NO4        g518(.A(new_new_n254_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n541_));
  NO3        g519(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n236_), .B(new_new_n36_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n404_), .B(i_1_), .Y(new_new_n544_));
  NOi31      g522(.An(new_new_n544_), .B(new_new_n443_), .C(new_new_n73_), .Y(new_new_n545_));
  AN4        g523(.A(new_new_n545_), .B(new_new_n401_), .C(new_new_n481_), .D(i_2_), .Y(new_new_n546_));
  NO2        g524(.A(new_new_n415_), .B(new_new_n181_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n547_), .B(new_new_n546_), .Y(new_new_n548_));
  NOi21      g526(.An(i_10_), .B(i_6_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n551_));
  NA2        g529(.A(new_new_n315_), .B(new_new_n169_), .Y(new_new_n552_));
  AOI220     g530(.A0(new_new_n552_), .A1(new_new_n426_), .B0(new_new_n187_), .B1(new_new_n185_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n200_), .B(new_new_n37_), .Y(new_new_n554_));
  NOi31      g532(.An(new_new_n150_), .B(new_new_n554_), .C(new_new_n329_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n555_), .B(new_new_n553_), .Y(new_new_n556_));
  INV        g534(.A(new_new_n316_), .Y(new_new_n557_));
  NO2        g535(.A(i_12_), .B(new_new_n86_), .Y(new_new_n558_));
  NA3        g536(.A(new_new_n558_), .B(new_new_n281_), .C(new_new_n537_), .Y(new_new_n559_));
  NA3        g537(.A(new_new_n383_), .B(new_new_n290_), .C(new_new_n220_), .Y(new_new_n560_));
  AOI210     g538(.A0(new_new_n560_), .A1(new_new_n559_), .B0(new_new_n557_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n178_), .B(i_0_), .Y(new_new_n562_));
  NO3        g540(.A(new_new_n562_), .B(new_new_n337_), .C(new_new_n304_), .Y(new_new_n563_));
  OR2        g541(.A(i_2_), .B(i_5_), .Y(new_new_n564_));
  OR2        g542(.A(new_new_n564_), .B(new_new_n396_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n565_), .B(new_new_n479_), .Y(new_new_n566_));
  NO3        g544(.A(new_new_n566_), .B(new_new_n563_), .C(new_new_n561_), .Y(new_new_n567_));
  NA4        g545(.A(new_new_n567_), .B(new_new_n556_), .C(new_new_n548_), .D(new_new_n540_), .Y(new_new_n568_));
  NO4        g546(.A(new_new_n568_), .B(new_new_n529_), .C(new_new_n512_), .D(new_new_n490_), .Y(new_new_n569_));
  NA4        g547(.A(new_new_n569_), .B(new_new_n430_), .C(new_new_n351_), .D(new_new_n312_), .Y(ori7));
  NO2        g548(.A(new_new_n95_), .B(new_new_n54_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n111_), .B(new_new_n92_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n382_), .B(new_new_n572_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n466_), .B(new_new_n84_), .Y(new_new_n574_));
  NA2        g552(.A(i_11_), .B(new_new_n195_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n148_), .B(new_new_n575_), .Y(new_new_n576_));
  OAI210     g554(.A0(new_new_n576_), .A1(new_new_n574_), .B0(new_new_n573_), .Y(new_new_n577_));
  NA3        g555(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n240_), .B(i_4_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n579_), .B(i_8_), .Y(new_new_n580_));
  NO2        g558(.A(new_new_n108_), .B(new_new_n578_), .Y(new_new_n581_));
  NA2        g559(.A(i_2_), .B(new_new_n86_), .Y(new_new_n582_));
  OAI210     g560(.A0(new_new_n89_), .A1(new_new_n205_), .B0(new_new_n206_), .Y(new_new_n583_));
  NO2        g561(.A(i_7_), .B(new_new_n37_), .Y(new_new_n584_));
  NA2        g562(.A(i_4_), .B(i_8_), .Y(new_new_n585_));
  AOI210     g563(.A0(new_new_n585_), .A1(new_new_n307_), .B0(new_new_n584_), .Y(new_new_n586_));
  OAI220     g564(.A0(new_new_n586_), .A1(new_new_n582_), .B0(new_new_n583_), .B1(i_13_), .Y(new_new_n587_));
  NO4        g565(.A(new_new_n587_), .B(new_new_n581_), .C(new_new_n577_), .D(new_new_n571_), .Y(new_new_n588_));
  AOI210     g566(.A0(new_new_n132_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n589_));
  AOI210     g567(.A0(new_new_n589_), .A1(new_new_n240_), .B0(new_new_n166_), .Y(new_new_n590_));
  OR2        g568(.A(i_6_), .B(i_10_), .Y(new_new_n591_));
  NO2        g569(.A(new_new_n591_), .B(new_new_n23_), .Y(new_new_n592_));
  OR3        g570(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n593_));
  INV        g571(.A(new_new_n202_), .Y(new_new_n594_));
  INV        g572(.A(new_new_n592_), .Y(new_new_n595_));
  OA220      g573(.A0(new_new_n595_), .A1(new_new_n557_), .B0(new_new_n590_), .B1(new_new_n273_), .Y(new_new_n596_));
  AOI210     g574(.A0(new_new_n596_), .A1(new_new_n588_), .B0(new_new_n63_), .Y(new_new_n597_));
  NOi21      g575(.An(i_11_), .B(i_7_), .Y(new_new_n598_));
  AO210      g576(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n599_), .B(new_new_n598_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n600_), .B(new_new_n210_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n601_), .B(new_new_n63_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n603_));
  AO210      g581(.A0(new_new_n603_), .A1(new_new_n376_), .B0(new_new_n41_), .Y(new_new_n604_));
  NO3        g582(.A(new_new_n262_), .B(new_new_n211_), .C(new_new_n575_), .Y(new_new_n605_));
  OAI210     g583(.A0(new_new_n605_), .A1(new_new_n229_), .B0(new_new_n63_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n397_), .B(new_new_n31_), .Y(new_new_n607_));
  OR2        g585(.A(new_new_n211_), .B(new_new_n111_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n608_), .B(new_new_n607_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n63_), .B(i_9_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n610_), .B(i_4_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n611_), .B(new_new_n609_), .Y(new_new_n612_));
  NO2        g590(.A(i_1_), .B(i_12_), .Y(new_new_n613_));
  NA3        g591(.A(new_new_n612_), .B(new_new_n606_), .C(new_new_n604_), .Y(new_new_n614_));
  OAI210     g592(.A0(new_new_n614_), .A1(new_new_n602_), .B0(i_6_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n240_), .B(new_new_n86_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n616_), .B(i_11_), .Y(new_new_n617_));
  INV        g595(.A(new_new_n444_), .Y(new_new_n618_));
  NO4        g596(.A(new_new_n217_), .B(new_new_n132_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n619_));
  NA2        g597(.A(new_new_n619_), .B(new_new_n610_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n240_), .B(i_6_), .Y(new_new_n621_));
  NO3        g599(.A(new_new_n591_), .B(new_new_n236_), .C(new_new_n23_), .Y(new_new_n622_));
  AOI210     g600(.A0(i_1_), .A1(new_new_n263_), .B0(new_new_n622_), .Y(new_new_n623_));
  OAI210     g601(.A0(new_new_n623_), .A1(new_new_n44_), .B0(new_new_n620_), .Y(new_new_n624_));
  NA3        g602(.A(new_new_n515_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n625_));
  INV        g603(.A(i_2_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n142_), .B(i_9_), .Y(new_new_n627_));
  NA3        g605(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n46_), .B(i_1_), .Y(new_new_n629_));
  NA3        g607(.A(new_new_n629_), .B(new_new_n272_), .C(new_new_n44_), .Y(new_new_n630_));
  OAI220     g608(.A0(new_new_n630_), .A1(new_new_n628_), .B0(new_new_n627_), .B1(new_new_n626_), .Y(new_new_n631_));
  NA3        g609(.A(new_new_n610_), .B(new_new_n316_), .C(i_6_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n23_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n463_), .A1(new_new_n408_), .B0(new_new_n245_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n582_), .Y(new_new_n635_));
  NAi21      g613(.An(new_new_n625_), .B(new_new_n94_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n629_), .B(new_new_n272_), .Y(new_new_n637_));
  NO2        g615(.A(i_11_), .B(new_new_n37_), .Y(new_new_n638_));
  NA2        g616(.A(new_new_n638_), .B(new_new_n24_), .Y(new_new_n639_));
  OAI210     g617(.A0(new_new_n639_), .A1(new_new_n637_), .B0(new_new_n636_), .Y(new_new_n640_));
  OR4        g618(.A(new_new_n640_), .B(new_new_n635_), .C(new_new_n633_), .D(new_new_n631_), .Y(new_new_n641_));
  NO3        g619(.A(new_new_n641_), .B(new_new_n624_), .C(new_new_n618_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n240_), .B(new_new_n104_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(new_new_n598_), .Y(new_new_n644_));
  NA2        g622(.A(new_new_n644_), .B(i_1_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n593_), .Y(new_new_n646_));
  NO2        g624(.A(new_new_n403_), .B(new_new_n86_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n646_), .B(new_new_n46_), .Y(new_new_n648_));
  NA2        g626(.A(i_3_), .B(new_new_n195_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n649_), .B(new_new_n118_), .Y(new_new_n650_));
  AN2        g628(.A(new_new_n650_), .B(new_new_n521_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n236_), .B(new_new_n44_), .Y(new_new_n652_));
  NO3        g630(.A(new_new_n652_), .B(new_new_n310_), .C(new_new_n241_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n121_), .B(new_new_n37_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n654_), .B(i_6_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n86_), .B(i_9_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n656_), .B(new_new_n63_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n657_), .B(new_new_n613_), .Y(new_new_n658_));
  NO4        g636(.A(new_new_n658_), .B(new_new_n655_), .C(new_new_n653_), .D(i_4_), .Y(new_new_n659_));
  NA2        g637(.A(i_1_), .B(i_3_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n445_), .B(new_new_n95_), .Y(new_new_n661_));
  AOI210     g639(.A0(new_new_n652_), .A1(new_new_n549_), .B0(new_new_n661_), .Y(new_new_n662_));
  NO2        g640(.A(new_new_n662_), .B(new_new_n660_), .Y(new_new_n663_));
  NO3        g641(.A(new_new_n663_), .B(new_new_n659_), .C(new_new_n651_), .Y(new_new_n664_));
  NA4        g642(.A(new_new_n664_), .B(new_new_n648_), .C(new_new_n642_), .D(new_new_n615_), .Y(new_new_n665_));
  NO3        g643(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n666_));
  AN2        g644(.A(new_new_n249_), .B(new_new_n86_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n368_), .B(new_new_n367_), .Y(new_new_n668_));
  NA3        g646(.A(new_new_n466_), .B(new_new_n501_), .C(new_new_n46_), .Y(new_new_n669_));
  NO3        g647(.A(new_new_n464_), .B(new_new_n585_), .C(new_new_n86_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n670_), .B(new_new_n25_), .Y(new_new_n671_));
  NA3        g649(.A(new_new_n671_), .B(new_new_n669_), .C(new_new_n668_), .Y(new_new_n672_));
  OAI210     g650(.A0(new_new_n672_), .A1(new_new_n667_), .B0(i_1_), .Y(new_new_n673_));
  AOI210     g651(.A0(new_new_n272_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n674_));
  NO2        g652(.A(new_new_n366_), .B(i_2_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n675_), .B(new_new_n674_), .Y(new_new_n676_));
  OAI210     g654(.A0(new_new_n632_), .A1(new_new_n435_), .B0(new_new_n676_), .Y(new_new_n677_));
  INV        g655(.A(new_new_n677_), .Y(new_new_n678_));
  AOI210     g656(.A0(new_new_n678_), .A1(new_new_n673_), .B0(i_13_), .Y(new_new_n679_));
  OR2        g657(.A(i_11_), .B(i_7_), .Y(new_new_n680_));
  AOI210     g658(.A0(new_new_n628_), .A1(new_new_n54_), .B0(i_12_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n464_), .B(new_new_n24_), .Y(new_new_n682_));
  AOI220     g660(.A0(new_new_n682_), .A1(new_new_n647_), .B0(new_new_n249_), .B1(new_new_n135_), .Y(new_new_n683_));
  OAI220     g661(.A0(new_new_n683_), .A1(new_new_n41_), .B0(new_new_n1012_), .B1(new_new_n95_), .Y(new_new_n684_));
  INV        g662(.A(new_new_n684_), .Y(new_new_n685_));
  INV        g663(.A(new_new_n118_), .Y(new_new_n686_));
  AOI220     g664(.A0(new_new_n686_), .A1(new_new_n72_), .B0(new_new_n383_), .B1(new_new_n629_), .Y(new_new_n687_));
  NO2        g665(.A(new_new_n687_), .B(new_new_n246_), .Y(new_new_n688_));
  AOI210     g666(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n689_));
  NOi31      g667(.An(new_new_n689_), .B(new_new_n574_), .C(new_new_n44_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n131_), .B(i_13_), .Y(new_new_n691_));
  NO2        g669(.A(new_new_n628_), .B(new_new_n118_), .Y(new_new_n692_));
  INV        g670(.A(new_new_n692_), .Y(new_new_n693_));
  OAI220     g671(.A0(new_new_n693_), .A1(new_new_n71_), .B0(new_new_n691_), .B1(new_new_n674_), .Y(new_new_n694_));
  NO3        g672(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n26_), .B(new_new_n195_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n696_), .B(i_7_), .Y(new_new_n697_));
  AOI220     g675(.A0(new_new_n383_), .A1(new_new_n629_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n698_));
  OAI220     g676(.A0(new_new_n698_), .A1(new_new_n580_), .B0(new_new_n1014_), .B1(new_new_n594_), .Y(new_new_n699_));
  NO4        g677(.A(new_new_n699_), .B(new_new_n694_), .C(new_new_n690_), .D(new_new_n688_), .Y(new_new_n700_));
  OR2        g678(.A(i_11_), .B(i_6_), .Y(new_new_n701_));
  NA3        g679(.A(new_new_n579_), .B(new_new_n696_), .C(i_7_), .Y(new_new_n702_));
  AOI210     g680(.A0(new_new_n702_), .A1(new_new_n693_), .B0(new_new_n701_), .Y(new_new_n703_));
  NA3        g681(.A(new_new_n397_), .B(new_new_n584_), .C(new_new_n100_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n617_), .B(i_13_), .Y(new_new_n705_));
  NA2        g683(.A(new_new_n105_), .B(new_new_n696_), .Y(new_new_n706_));
  NAi21      g684(.An(i_11_), .B(i_12_), .Y(new_new_n707_));
  NOi41      g685(.An(new_new_n114_), .B(new_new_n707_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n708_), .B(new_new_n706_), .Y(new_new_n709_));
  NA3        g687(.A(new_new_n709_), .B(new_new_n705_), .C(new_new_n704_), .Y(new_new_n710_));
  OAI210     g688(.A0(new_new_n710_), .A1(new_new_n703_), .B0(new_new_n63_), .Y(new_new_n711_));
  NO2        g689(.A(i_2_), .B(i_12_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n365_), .B(new_new_n712_), .Y(new_new_n713_));
  NA2        g691(.A(i_8_), .B(new_new_n25_), .Y(new_new_n714_));
  NO3        g692(.A(new_new_n714_), .B(new_new_n382_), .C(new_new_n579_), .Y(new_new_n715_));
  OAI210     g693(.A0(new_new_n715_), .A1(new_new_n367_), .B0(new_new_n365_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n132_), .B(i_2_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n717_), .B(new_new_n613_), .Y(new_new_n718_));
  NA3        g696(.A(new_new_n718_), .B(new_new_n716_), .C(new_new_n713_), .Y(new_new_n719_));
  NA3        g697(.A(new_new_n719_), .B(new_new_n45_), .C(new_new_n228_), .Y(new_new_n720_));
  NA4        g698(.A(new_new_n720_), .B(new_new_n711_), .C(new_new_n700_), .D(new_new_n685_), .Y(new_new_n721_));
  OR4        g699(.A(new_new_n721_), .B(new_new_n679_), .C(new_new_n665_), .D(new_new_n597_), .Y(ori5));
  NA2        g700(.A(new_new_n644_), .B(new_new_n275_), .Y(new_new_n723_));
  AN2        g701(.A(new_new_n24_), .B(i_10_), .Y(new_new_n724_));
  NA3        g702(.A(new_new_n724_), .B(new_new_n712_), .C(new_new_n111_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n580_), .B(i_11_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n89_), .B(new_new_n726_), .Y(new_new_n727_));
  NA3        g705(.A(new_new_n727_), .B(new_new_n725_), .C(new_new_n723_), .Y(new_new_n728_));
  NO3        g706(.A(i_11_), .B(new_new_n240_), .C(i_13_), .Y(new_new_n729_));
  NO2        g707(.A(new_new_n128_), .B(new_new_n23_), .Y(new_new_n730_));
  NA2        g708(.A(i_12_), .B(i_8_), .Y(new_new_n731_));
  OAI210     g709(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n731_), .Y(new_new_n732_));
  INV        g710(.A(new_new_n434_), .Y(new_new_n733_));
  AOI220     g711(.A0(new_new_n316_), .A1(new_new_n551_), .B0(new_new_n732_), .B1(new_new_n730_), .Y(new_new_n734_));
  INV        g712(.A(new_new_n734_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n735_), .B(new_new_n728_), .Y(new_new_n736_));
  INV        g714(.A(new_new_n176_), .Y(new_new_n737_));
  INV        g715(.A(new_new_n249_), .Y(new_new_n738_));
  OAI210     g716(.A0(new_new_n675_), .A1(new_new_n436_), .B0(new_new_n114_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n739_), .A1(new_new_n738_), .B0(new_new_n737_), .Y(new_new_n740_));
  NO2        g718(.A(new_new_n445_), .B(new_new_n26_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n741_), .B(new_new_n408_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n742_), .B(i_2_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n743_), .Y(new_new_n744_));
  AOI210     g722(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n404_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n745_), .A1(new_new_n744_), .B0(new_new_n740_), .Y(new_new_n746_));
  NO2        g724(.A(new_new_n193_), .B(new_new_n129_), .Y(new_new_n747_));
  OAI210     g725(.A0(new_new_n747_), .A1(new_new_n730_), .B0(i_2_), .Y(new_new_n748_));
  INV        g726(.A(new_new_n177_), .Y(new_new_n749_));
  NO3        g727(.A(new_new_n599_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n750_));
  AOI210     g728(.A0(new_new_n749_), .A1(new_new_n89_), .B0(new_new_n750_), .Y(new_new_n751_));
  AOI210     g729(.A0(new_new_n751_), .A1(new_new_n748_), .B0(new_new_n195_), .Y(new_new_n752_));
  OA210      g730(.A0(new_new_n600_), .A1(new_new_n130_), .B0(i_13_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n202_), .B(new_new_n205_), .Y(new_new_n754_));
  NA2        g732(.A(new_new_n156_), .B(new_new_n575_), .Y(new_new_n755_));
  AOI210     g733(.A0(new_new_n755_), .A1(new_new_n754_), .B0(new_new_n370_), .Y(new_new_n756_));
  AOI210     g734(.A0(new_new_n211_), .A1(new_new_n152_), .B0(new_new_n501_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n757_), .B(new_new_n408_), .Y(new_new_n758_));
  NO2        g736(.A(new_new_n105_), .B(new_new_n44_), .Y(new_new_n759_));
  INV        g737(.A(new_new_n305_), .Y(new_new_n760_));
  NA4        g738(.A(new_new_n760_), .B(new_new_n307_), .C(new_new_n128_), .D(new_new_n42_), .Y(new_new_n761_));
  OAI210     g739(.A0(new_new_n761_), .A1(new_new_n759_), .B0(new_new_n758_), .Y(new_new_n762_));
  NO4        g740(.A(new_new_n762_), .B(new_new_n756_), .C(new_new_n753_), .D(new_new_n752_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n551_), .B(new_new_n28_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n729_), .B(new_new_n282_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n765_), .B(new_new_n764_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n62_), .B(i_12_), .Y(new_new_n767_));
  NO2        g745(.A(new_new_n767_), .B(new_new_n130_), .Y(new_new_n768_));
  NO2        g746(.A(new_new_n768_), .B(new_new_n575_), .Y(new_new_n769_));
  AOI220     g747(.A0(new_new_n769_), .A1(new_new_n36_), .B0(new_new_n766_), .B1(new_new_n46_), .Y(new_new_n770_));
  NA4        g748(.A(new_new_n770_), .B(new_new_n763_), .C(new_new_n746_), .D(new_new_n736_), .Y(ori6));
  NO3        g749(.A(new_new_n258_), .B(new_new_n309_), .C(i_1_), .Y(new_new_n772_));
  NO2        g750(.A(new_new_n189_), .B(new_new_n143_), .Y(new_new_n773_));
  OAI210     g751(.A0(new_new_n773_), .A1(new_new_n772_), .B0(new_new_n717_), .Y(new_new_n774_));
  NA4        g752(.A(new_new_n384_), .B(new_new_n465_), .C(new_new_n71_), .D(new_new_n104_), .Y(new_new_n775_));
  INV        g753(.A(new_new_n775_), .Y(new_new_n776_));
  NO2        g754(.A(new_new_n223_), .B(new_new_n470_), .Y(new_new_n777_));
  NO2        g755(.A(new_new_n776_), .B(new_new_n328_), .Y(new_new_n778_));
  AO210      g756(.A0(new_new_n778_), .A1(new_new_n774_), .B0(i_12_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n558_), .B(new_new_n63_), .Y(new_new_n780_));
  BUFFER     g758(.A(new_new_n603_), .Y(new_new_n781_));
  NA2        g759(.A(new_new_n781_), .B(new_new_n780_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n782_), .B(new_new_n73_), .Y(new_new_n783_));
  INV        g761(.A(new_new_n327_), .Y(new_new_n784_));
  NA2        g762(.A(new_new_n75_), .B(new_new_n135_), .Y(new_new_n785_));
  INV        g763(.A(new_new_n128_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n786_), .B(new_new_n46_), .Y(new_new_n787_));
  AOI210     g765(.A0(new_new_n787_), .A1(new_new_n785_), .B0(new_new_n784_), .Y(new_new_n788_));
  NO3        g766(.A(new_new_n254_), .B(new_new_n136_), .C(i_9_), .Y(new_new_n789_));
  NA2        g767(.A(new_new_n789_), .B(new_new_n767_), .Y(new_new_n790_));
  AOI210     g768(.A0(new_new_n790_), .A1(new_new_n499_), .B0(new_new_n189_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n32_), .B(i_11_), .Y(new_new_n792_));
  NAi32      g770(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n793_));
  NO2        g771(.A(new_new_n701_), .B(new_new_n793_), .Y(new_new_n794_));
  OAI210     g772(.A0(new_new_n666_), .A1(new_new_n543_), .B0(new_new_n542_), .Y(new_new_n795_));
  NAi21      g773(.An(new_new_n794_), .B(new_new_n795_), .Y(new_new_n796_));
  OR3        g774(.A(new_new_n796_), .B(new_new_n791_), .C(new_new_n788_), .Y(new_new_n797_));
  NO2        g775(.A(new_new_n680_), .B(i_2_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n799_));
  NO2        g777(.A(new_new_n799_), .B(new_new_n396_), .Y(new_new_n800_));
  NA2        g778(.A(new_new_n800_), .B(new_new_n798_), .Y(new_new_n801_));
  AO220      g779(.A0(new_new_n356_), .A1(new_new_n346_), .B0(new_new_n388_), .B1(new_new_n575_), .Y(new_new_n802_));
  NA3        g780(.A(new_new_n802_), .B(new_new_n259_), .C(i_7_), .Y(new_new_n803_));
  OR2        g781(.A(new_new_n600_), .B(new_new_n436_), .Y(new_new_n804_));
  NA3        g782(.A(new_new_n804_), .B(new_new_n151_), .C(new_new_n69_), .Y(new_new_n805_));
  AO210      g783(.A0(new_new_n477_), .A1(new_new_n733_), .B0(new_new_n36_), .Y(new_new_n806_));
  NA4        g784(.A(new_new_n806_), .B(new_new_n805_), .C(new_new_n803_), .D(new_new_n801_), .Y(new_new_n807_));
  OAI210     g785(.A0(new_new_n616_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n808_));
  AOI220     g786(.A0(new_new_n808_), .A1(new_new_n542_), .B0(new_new_n777_), .B1(new_new_n697_), .Y(new_new_n809_));
  NA3        g787(.A(new_new_n370_), .B(new_new_n242_), .C(new_new_n151_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n388_), .B(new_new_n70_), .Y(new_new_n811_));
  NA4        g789(.A(new_new_n811_), .B(new_new_n810_), .C(new_new_n809_), .D(new_new_n583_), .Y(new_new_n812_));
  AO210      g790(.A0(new_new_n501_), .A1(new_new_n46_), .B0(new_new_n88_), .Y(new_new_n813_));
  NA3        g791(.A(new_new_n813_), .B(new_new_n466_), .C(new_new_n220_), .Y(new_new_n814_));
  AOI210     g792(.A0(new_new_n436_), .A1(new_new_n434_), .B0(new_new_n541_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n591_), .B(new_new_n105_), .Y(new_new_n816_));
  OAI210     g794(.A0(new_new_n816_), .A1(new_new_n115_), .B0(new_new_n394_), .Y(new_new_n817_));
  INV        g795(.A(new_new_n565_), .Y(new_new_n818_));
  NA3        g796(.A(new_new_n818_), .B(new_new_n327_), .C(i_7_), .Y(new_new_n819_));
  NA4        g797(.A(new_new_n819_), .B(new_new_n817_), .C(new_new_n815_), .D(new_new_n814_), .Y(new_new_n820_));
  NO4        g798(.A(new_new_n820_), .B(new_new_n812_), .C(new_new_n807_), .D(new_new_n797_), .Y(new_new_n821_));
  NA4        g799(.A(new_new_n821_), .B(new_new_n783_), .C(new_new_n779_), .D(new_new_n378_), .Y(ori3));
  NA2        g800(.A(i_6_), .B(i_7_), .Y(new_new_n823_));
  NO2        g801(.A(new_new_n823_), .B(i_0_), .Y(new_new_n824_));
  NO2        g802(.A(i_11_), .B(new_new_n240_), .Y(new_new_n825_));
  OAI210     g803(.A0(new_new_n824_), .A1(new_new_n297_), .B0(new_new_n825_), .Y(new_new_n826_));
  NO2        g804(.A(new_new_n826_), .B(new_new_n195_), .Y(new_new_n827_));
  NO3        g805(.A(new_new_n441_), .B(new_new_n92_), .C(new_new_n44_), .Y(new_new_n828_));
  OA210      g806(.A0(new_new_n828_), .A1(new_new_n827_), .B0(new_new_n178_), .Y(new_new_n829_));
  NA3        g807(.A(new_new_n810_), .B(new_new_n583_), .C(new_new_n369_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n830_), .B(new_new_n40_), .Y(new_new_n831_));
  NOi21      g809(.An(new_new_n99_), .B(new_new_n742_), .Y(new_new_n832_));
  NO3        g810(.A(new_new_n608_), .B(new_new_n445_), .C(new_new_n135_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n397_), .B(new_new_n45_), .Y(new_new_n834_));
  AN2        g812(.A(new_new_n443_), .B(new_new_n55_), .Y(new_new_n835_));
  NO3        g813(.A(new_new_n835_), .B(new_new_n833_), .C(new_new_n832_), .Y(new_new_n836_));
  AOI210     g814(.A0(new_new_n836_), .A1(new_new_n831_), .B0(new_new_n48_), .Y(new_new_n837_));
  NO4        g815(.A(new_new_n374_), .B(new_new_n381_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n189_), .B(new_new_n549_), .Y(new_new_n839_));
  NOi21      g817(.An(new_new_n839_), .B(new_new_n838_), .Y(new_new_n840_));
  NA2        g818(.A(new_new_n689_), .B(new_new_n656_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n331_), .B(i_5_), .Y(new_new_n842_));
  OAI220     g820(.A0(new_new_n842_), .A1(new_new_n841_), .B0(new_new_n840_), .B1(new_new_n63_), .Y(new_new_n843_));
  NOi21      g821(.An(i_5_), .B(i_9_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n844_), .B(new_new_n432_), .Y(new_new_n845_));
  BUFFER     g823(.A(new_new_n272_), .Y(new_new_n846_));
  AOI210     g824(.A0(new_new_n846_), .A1(new_new_n463_), .B0(new_new_n670_), .Y(new_new_n847_));
  NO3        g825(.A(new_new_n400_), .B(new_new_n272_), .C(new_new_n73_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n179_), .B(new_new_n152_), .Y(new_new_n849_));
  AOI210     g827(.A0(new_new_n849_), .A1(new_new_n248_), .B0(new_new_n848_), .Y(new_new_n850_));
  OAI220     g828(.A0(new_new_n850_), .A1(new_new_n184_), .B0(new_new_n847_), .B1(new_new_n845_), .Y(new_new_n851_));
  NO4        g829(.A(new_new_n851_), .B(new_new_n843_), .C(new_new_n837_), .D(new_new_n829_), .Y(new_new_n852_));
  NA2        g830(.A(new_new_n189_), .B(new_new_n24_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n654_), .B(new_new_n572_), .Y(new_new_n854_));
  NO2        g832(.A(new_new_n854_), .B(new_new_n853_), .Y(new_new_n855_));
  INV        g833(.A(new_new_n855_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n550_), .B(i_0_), .Y(new_new_n857_));
  NO4        g835(.A(new_new_n564_), .B(new_new_n217_), .C(new_new_n404_), .D(new_new_n396_), .Y(new_new_n858_));
  NA2        g836(.A(new_new_n858_), .B(i_11_), .Y(new_new_n859_));
  AN2        g837(.A(new_new_n99_), .B(new_new_n247_), .Y(new_new_n860_));
  NA2        g838(.A(new_new_n729_), .B(new_new_n328_), .Y(new_new_n861_));
  AOI210     g839(.A0(new_new_n466_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n862_));
  OAI220     g840(.A0(new_new_n862_), .A1(new_new_n861_), .B0(new_new_n639_), .B1(new_new_n517_), .Y(new_new_n863_));
  NO2        g841(.A(new_new_n256_), .B(new_new_n158_), .Y(new_new_n864_));
  NA2        g842(.A(i_0_), .B(i_10_), .Y(new_new_n865_));
  INV        g843(.A(new_new_n520_), .Y(new_new_n866_));
  NO4        g844(.A(new_new_n118_), .B(new_new_n58_), .C(new_new_n649_), .D(i_5_), .Y(new_new_n867_));
  AO220      g845(.A0(new_new_n867_), .A1(new_new_n866_), .B0(new_new_n864_), .B1(i_6_), .Y(new_new_n868_));
  AOI220     g846(.A0(new_new_n331_), .A1(new_new_n101_), .B0(new_new_n189_), .B1(new_new_n84_), .Y(new_new_n869_));
  NA2        g847(.A(new_new_n544_), .B(i_4_), .Y(new_new_n870_));
  NA2        g848(.A(new_new_n191_), .B(new_new_n205_), .Y(new_new_n871_));
  OAI220     g849(.A0(new_new_n871_), .A1(new_new_n861_), .B0(new_new_n870_), .B1(new_new_n869_), .Y(new_new_n872_));
  NO4        g850(.A(new_new_n872_), .B(new_new_n868_), .C(new_new_n863_), .D(new_new_n860_), .Y(new_new_n873_));
  NA3        g851(.A(new_new_n873_), .B(new_new_n859_), .C(new_new_n856_), .Y(new_new_n874_));
  NA2        g852(.A(i_11_), .B(i_9_), .Y(new_new_n875_));
  NO2        g853(.A(new_new_n48_), .B(i_7_), .Y(new_new_n876_));
  NA2        g854(.A(new_new_n385_), .B(new_new_n182_), .Y(new_new_n877_));
  NA2        g855(.A(new_new_n877_), .B(new_new_n165_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n179_), .B(i_0_), .Y(new_new_n879_));
  INV        g857(.A(new_new_n879_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n462_), .B(new_new_n234_), .Y(new_new_n881_));
  INV        g859(.A(new_new_n393_), .Y(new_new_n882_));
  OAI220     g860(.A0(new_new_n882_), .A1(new_new_n845_), .B0(new_new_n881_), .B1(new_new_n880_), .Y(new_new_n883_));
  NO2        g861(.A(new_new_n883_), .B(new_new_n878_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n638_), .B(new_new_n125_), .Y(new_new_n885_));
  NO2        g863(.A(i_6_), .B(new_new_n885_), .Y(new_new_n886_));
  AOI210     g864(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n887_));
  NA2        g865(.A(new_new_n176_), .B(new_new_n106_), .Y(new_new_n888_));
  NOi32      g866(.An(new_new_n887_), .Bn(new_new_n191_), .C(new_new_n888_), .Y(new_new_n889_));
  NA2        g867(.A(new_new_n584_), .B(new_new_n328_), .Y(new_new_n890_));
  NO2        g868(.A(new_new_n890_), .B(new_new_n834_), .Y(new_new_n891_));
  NO3        g869(.A(new_new_n891_), .B(new_new_n889_), .C(new_new_n886_), .Y(new_new_n892_));
  NOi21      g870(.An(i_7_), .B(i_5_), .Y(new_new_n893_));
  NOi31      g871(.An(new_new_n893_), .B(i_0_), .C(new_new_n707_), .Y(new_new_n894_));
  NA2        g872(.A(new_new_n892_), .B(new_new_n884_), .Y(new_new_n895_));
  AN2        g873(.A(new_new_n330_), .B(new_new_n328_), .Y(new_new_n896_));
  OA210      g874(.A0(new_new_n462_), .A1(new_new_n226_), .B0(new_new_n461_), .Y(new_new_n897_));
  NA3        g875(.A(new_new_n799_), .B(new_new_n380_), .C(new_new_n616_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n95_), .B(new_new_n44_), .Y(new_new_n899_));
  NO2        g877(.A(new_new_n75_), .B(new_new_n731_), .Y(new_new_n900_));
  AOI220     g878(.A0(new_new_n900_), .A1(new_new_n899_), .B0(new_new_n178_), .B1(new_new_n572_), .Y(new_new_n901_));
  AOI210     g879(.A0(new_new_n901_), .A1(new_new_n898_), .B0(new_new_n47_), .Y(new_new_n902_));
  NO3        g880(.A(new_new_n564_), .B(new_new_n354_), .C(new_new_n24_), .Y(new_new_n903_));
  INV        g881(.A(new_new_n903_), .Y(new_new_n904_));
  NO2        g882(.A(new_new_n578_), .B(new_new_n108_), .Y(new_new_n905_));
  NA2        g883(.A(new_new_n905_), .B(i_0_), .Y(new_new_n906_));
  OAI220     g884(.A0(new_new_n906_), .A1(new_new_n86_), .B0(new_new_n904_), .B1(new_new_n177_), .Y(new_new_n907_));
  NO3        g885(.A(new_new_n907_), .B(new_new_n902_), .C(new_new_n503_), .Y(new_new_n908_));
  INV        g886(.A(new_new_n908_), .Y(new_new_n909_));
  NO3        g887(.A(new_new_n909_), .B(new_new_n895_), .C(new_new_n874_), .Y(new_new_n910_));
  NO2        g888(.A(i_0_), .B(new_new_n707_), .Y(new_new_n911_));
  AOI210     g889(.A0(new_new_n780_), .A1(new_new_n668_), .B0(new_new_n888_), .Y(new_new_n912_));
  INV        g890(.A(new_new_n912_), .Y(new_new_n913_));
  NO2        g891(.A(new_new_n795_), .B(new_new_n391_), .Y(new_new_n914_));
  NA3        g892(.A(new_new_n824_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n915_));
  NA2        g893(.A(new_new_n825_), .B(i_9_), .Y(new_new_n916_));
  AOI210     g894(.A0(new_new_n915_), .A1(new_new_n483_), .B0(new_new_n916_), .Y(new_new_n917_));
  OAI210     g895(.A0(new_new_n248_), .A1(i_9_), .B0(new_new_n233_), .Y(new_new_n918_));
  AOI210     g896(.A0(new_new_n918_), .A1(new_new_n857_), .B0(new_new_n158_), .Y(new_new_n919_));
  NO3        g897(.A(new_new_n919_), .B(new_new_n917_), .C(new_new_n914_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n920_), .B(new_new_n913_), .Y(new_new_n921_));
  NA2        g899(.A(new_new_n896_), .B(new_new_n370_), .Y(new_new_n922_));
  AOI210     g900(.A0(new_new_n304_), .A1(new_new_n167_), .B0(new_new_n922_), .Y(new_new_n923_));
  INV        g901(.A(new_new_n923_), .Y(new_new_n924_));
  NO3        g902(.A(new_new_n865_), .B(new_new_n844_), .C(new_new_n193_), .Y(new_new_n925_));
  AOI220     g903(.A0(new_new_n925_), .A1(i_11_), .B0(new_new_n545_), .B1(new_new_n75_), .Y(new_new_n926_));
  NO3        g904(.A(new_new_n212_), .B(new_new_n381_), .C(i_0_), .Y(new_new_n927_));
  OAI210     g905(.A0(new_new_n927_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n928_));
  INV        g906(.A(new_new_n220_), .Y(new_new_n929_));
  OAI220     g907(.A0(new_new_n514_), .A1(new_new_n143_), .B0(new_new_n621_), .B1(new_new_n594_), .Y(new_new_n930_));
  NA3        g908(.A(new_new_n930_), .B(new_new_n389_), .C(new_new_n929_), .Y(new_new_n931_));
  NA4        g909(.A(new_new_n931_), .B(new_new_n928_), .C(new_new_n926_), .D(new_new_n924_), .Y(new_new_n932_));
  NO2        g910(.A(new_new_n246_), .B(new_new_n95_), .Y(new_new_n933_));
  AOI210     g911(.A0(new_new_n933_), .A1(new_new_n911_), .B0(new_new_n112_), .Y(new_new_n934_));
  AOI220     g912(.A0(new_new_n893_), .A1(new_new_n471_), .B0(new_new_n824_), .B1(new_new_n168_), .Y(new_new_n935_));
  NA2        g913(.A(new_new_n346_), .B(new_new_n180_), .Y(new_new_n936_));
  OA220      g914(.A0(new_new_n936_), .A1(new_new_n935_), .B0(new_new_n934_), .B1(i_5_), .Y(new_new_n937_));
  AOI210     g915(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n938_));
  NA2        g916(.A(new_new_n938_), .B(new_new_n897_), .Y(new_new_n939_));
  NA3        g917(.A(new_new_n592_), .B(new_new_n189_), .C(new_new_n84_), .Y(new_new_n940_));
  NA2        g918(.A(new_new_n940_), .B(new_new_n527_), .Y(new_new_n941_));
  NO3        g919(.A(new_new_n834_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n942_));
  NA2        g920(.A(new_new_n476_), .B(new_new_n469_), .Y(new_new_n943_));
  NO3        g921(.A(new_new_n943_), .B(new_new_n942_), .C(new_new_n941_), .Y(new_new_n944_));
  NA3        g922(.A(new_new_n384_), .B(new_new_n176_), .C(new_new_n175_), .Y(new_new_n945_));
  NA3        g923(.A(new_new_n876_), .B(new_new_n297_), .C(new_new_n233_), .Y(new_new_n946_));
  NA2        g924(.A(new_new_n946_), .B(new_new_n945_), .Y(new_new_n947_));
  NA3        g925(.A(new_new_n384_), .B(new_new_n332_), .C(new_new_n224_), .Y(new_new_n948_));
  INV        g926(.A(new_new_n948_), .Y(new_new_n949_));
  NO3        g927(.A(new_new_n875_), .B(new_new_n220_), .C(new_new_n193_), .Y(new_new_n950_));
  NO3        g928(.A(new_new_n950_), .B(new_new_n949_), .C(new_new_n947_), .Y(new_new_n951_));
  NA4        g929(.A(new_new_n951_), .B(new_new_n944_), .C(new_new_n939_), .D(new_new_n937_), .Y(new_new_n952_));
  NO2        g930(.A(new_new_n86_), .B(i_5_), .Y(new_new_n953_));
  NA3        g931(.A(new_new_n825_), .B(new_new_n113_), .C(new_new_n128_), .Y(new_new_n954_));
  INV        g932(.A(new_new_n954_), .Y(new_new_n955_));
  NA2        g933(.A(new_new_n955_), .B(new_new_n953_), .Y(new_new_n956_));
  NA3        g934(.A(new_new_n307_), .B(i_5_), .C(new_new_n195_), .Y(new_new_n957_));
  NAi31      g935(.An(new_new_n245_), .B(new_new_n957_), .C(new_new_n246_), .Y(new_new_n958_));
  NO4        g936(.A(new_new_n243_), .B(new_new_n212_), .C(i_0_), .D(i_12_), .Y(new_new_n959_));
  AOI220     g937(.A0(new_new_n959_), .A1(new_new_n958_), .B0(new_new_n776_), .B1(new_new_n180_), .Y(new_new_n960_));
  AN2        g938(.A(new_new_n865_), .B(new_new_n158_), .Y(new_new_n961_));
  NO4        g939(.A(new_new_n961_), .B(i_12_), .C(new_new_n625_), .D(new_new_n135_), .Y(new_new_n962_));
  NA2        g940(.A(new_new_n962_), .B(new_new_n220_), .Y(new_new_n963_));
  NA3        g941(.A(new_new_n101_), .B(new_new_n549_), .C(i_11_), .Y(new_new_n964_));
  NO2        g942(.A(new_new_n964_), .B(new_new_n160_), .Y(new_new_n965_));
  NA2        g943(.A(new_new_n893_), .B(new_new_n459_), .Y(new_new_n966_));
  NA2        g944(.A(new_new_n64_), .B(new_new_n104_), .Y(new_new_n967_));
  OAI220     g945(.A0(new_new_n967_), .A1(new_new_n957_), .B0(new_new_n966_), .B1(new_new_n657_), .Y(new_new_n968_));
  AOI210     g946(.A0(new_new_n968_), .A1(new_new_n879_), .B0(new_new_n965_), .Y(new_new_n969_));
  NA4        g947(.A(new_new_n969_), .B(new_new_n963_), .C(new_new_n960_), .D(new_new_n956_), .Y(new_new_n970_));
  NO4        g948(.A(new_new_n970_), .B(new_new_n952_), .C(new_new_n932_), .D(new_new_n921_), .Y(new_new_n971_));
  OAI210     g949(.A0(new_new_n798_), .A1(new_new_n792_), .B0(new_new_n37_), .Y(new_new_n972_));
  NA3        g950(.A(new_new_n887_), .B(new_new_n365_), .C(i_5_), .Y(new_new_n973_));
  NA3        g951(.A(new_new_n973_), .B(new_new_n972_), .C(new_new_n590_), .Y(new_new_n974_));
  NA2        g952(.A(new_new_n974_), .B(new_new_n210_), .Y(new_new_n975_));
  BUFFER     g953(.A(new_new_n366_), .Y(new_new_n976_));
  NA2        g954(.A(new_new_n190_), .B(new_new_n191_), .Y(new_new_n977_));
  AO210      g955(.A0(new_new_n976_), .A1(new_new_n33_), .B0(new_new_n977_), .Y(new_new_n978_));
  NAi31      g956(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n979_));
  AOI210     g957(.A0(new_new_n121_), .A1(new_new_n70_), .B0(new_new_n979_), .Y(new_new_n980_));
  NO2        g958(.A(new_new_n980_), .B(new_new_n622_), .Y(new_new_n981_));
  NA2        g959(.A(new_new_n981_), .B(new_new_n978_), .Y(new_new_n982_));
  NO2        g960(.A(new_new_n453_), .B(new_new_n272_), .Y(new_new_n983_));
  NO2        g961(.A(new_new_n983_), .B(new_new_n858_), .Y(new_new_n984_));
  OAI210     g962(.A0(new_new_n964_), .A1(new_new_n152_), .B0(new_new_n984_), .Y(new_new_n985_));
  AOI210     g963(.A0(new_new_n982_), .A1(new_new_n48_), .B0(new_new_n985_), .Y(new_new_n986_));
  AOI210     g964(.A0(new_new_n986_), .A1(new_new_n975_), .B0(new_new_n73_), .Y(new_new_n987_));
  INV        g965(.A(new_new_n377_), .Y(new_new_n988_));
  NO2        g966(.A(new_new_n988_), .B(new_new_n737_), .Y(new_new_n989_));
  OAI210     g967(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n111_), .Y(new_new_n990_));
  NA2        g968(.A(new_new_n990_), .B(new_new_n76_), .Y(new_new_n991_));
  AOI210     g969(.A0(new_new_n938_), .A1(new_new_n876_), .B0(new_new_n894_), .Y(new_new_n992_));
  AOI210     g970(.A0(new_new_n992_), .A1(new_new_n991_), .B0(new_new_n660_), .Y(new_new_n993_));
  NA2        g971(.A(new_new_n266_), .B(new_new_n57_), .Y(new_new_n994_));
  AOI220     g972(.A0(new_new_n994_), .A1(new_new_n76_), .B0(new_new_n343_), .B1(new_new_n258_), .Y(new_new_n995_));
  NO2        g973(.A(new_new_n995_), .B(new_new_n240_), .Y(new_new_n996_));
  NO2        g974(.A(new_new_n996_), .B(new_new_n993_), .Y(new_new_n997_));
  OAI210     g975(.A0(new_new_n274_), .A1(new_new_n163_), .B0(new_new_n89_), .Y(new_new_n998_));
  NO2        g976(.A(new_new_n998_), .B(i_11_), .Y(new_new_n999_));
  NA2        g977(.A(new_new_n585_), .B(new_new_n217_), .Y(new_new_n1000_));
  OAI210     g978(.A0(new_new_n1000_), .A1(new_new_n887_), .B0(new_new_n210_), .Y(new_new_n1001_));
  NA2        g979(.A(new_new_n169_), .B(i_5_), .Y(new_new_n1002_));
  NO2        g980(.A(new_new_n1001_), .B(new_new_n1002_), .Y(new_new_n1003_));
  INV        g981(.A(new_new_n360_), .Y(new_new_n1004_));
  NO2        g982(.A(new_new_n1004_), .B(new_new_n41_), .Y(new_new_n1005_));
  NO3        g983(.A(new_new_n1005_), .B(new_new_n1003_), .C(new_new_n999_), .Y(new_new_n1006_));
  OAI210     g984(.A0(new_new_n997_), .A1(i_4_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  NO3        g985(.A(new_new_n1007_), .B(new_new_n989_), .C(new_new_n987_), .Y(new_new_n1008_));
  NA4        g986(.A(new_new_n1008_), .B(new_new_n971_), .C(new_new_n910_), .D(new_new_n852_), .Y(ori4));
  INV        g987(.A(new_new_n681_), .Y(new_new_n1012_));
  INV        g988(.A(new_new_n527_), .Y(new_new_n1013_));
  INV        g989(.A(new_new_n695_), .Y(new_new_n1014_));
endmodule


