//Benchmark atmr_intb_466_0.25

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n274_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n314_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n315_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  AOI220     o035(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n60_));
  OAI210     o038(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n60_), .Y(ori_ori_n61_));
  AOI220     o039(.A0(ori_ori_n61_), .A1(ori_ori_n55_), .B0(ori_ori_n59_), .B1(ori_ori_n31_), .Y(ori_ori_n62_));
  NO2        o040(.A(ori_ori_n62_), .B(x05), .Y(ori_ori_n63_));
  NA2        o041(.A(x09), .B(x05), .Y(ori_ori_n64_));
  NA2        o042(.A(x10), .B(x06), .Y(ori_ori_n65_));
  NA3        o043(.A(ori_ori_n65_), .B(ori_ori_n64_), .C(ori_ori_n28_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n66_), .B(x03), .Y(ori_ori_n67_));
  NOi31      o045(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n68_));
  INV        o046(.A(x07), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n24_), .Y(ori_ori_n70_));
  NA2        o048(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n48_), .B(ori_ori_n71_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n73_));
  NO2        o051(.A(x08), .B(x01), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n73_), .B0(ori_ori_n35_), .Y(ori_ori_n75_));
  NO3        o053(.A(ori_ori_n75_), .B(ori_ori_n72_), .C(ori_ori_n70_), .Y(ori_ori_n76_));
  AN2        o054(.A(ori_ori_n76_), .B(ori_ori_n67_), .Y(ori_ori_n77_));
  INV        o055(.A(ori_ori_n75_), .Y(ori_ori_n78_));
  NA2        o056(.A(x11), .B(x00), .Y(ori_ori_n79_));
  NO2        o057(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n80_));
  NOi21      o058(.An(ori_ori_n79_), .B(ori_ori_n80_), .Y(ori_ori_n81_));
  INV        o059(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  NOi21      o060(.An(x01), .B(x10), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n84_));
  NO3        o062(.A(ori_ori_n84_), .B(ori_ori_n83_), .C(x06), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n85_), .B(ori_ori_n27_), .Y(ori_ori_n86_));
  OAI210     o064(.A0(ori_ori_n82_), .A1(x07), .B0(ori_ori_n86_), .Y(ori_ori_n87_));
  NO3        o065(.A(ori_ori_n87_), .B(ori_ori_n77_), .C(ori_ori_n63_), .Y(ori01));
  INV        o066(.A(x12), .Y(ori_ori_n89_));
  INV        o067(.A(x13), .Y(ori_ori_n90_));
  NO2        o068(.A(x10), .B(x01), .Y(ori_ori_n91_));
  NO2        o069(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n92_));
  NO2        o070(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n94_));
  NOi21      o072(.An(ori_ori_n94_), .B(ori_ori_n54_), .Y(ori_ori_n95_));
  NA2        o073(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n96_));
  NO2        o074(.A(ori_ori_n96_), .B(x05), .Y(ori_ori_n97_));
  INV        o075(.A(ori_ori_n95_), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n98_), .B(ori_ori_n65_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n100_));
  NA2        o078(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n104_));
  NA3        o082(.A(ori_ori_n104_), .B(ori_ori_n103_), .C(x13), .Y(ori_ori_n105_));
  NO2        o083(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n106_));
  NOi31      o084(.An(ori_ori_n105_), .B(ori_ori_n106_), .C(ori_ori_n102_), .Y(ori_ori_n107_));
  NO3        o085(.A(ori_ori_n107_), .B(x06), .C(x03), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n108_), .B(ori_ori_n99_), .Y(ori_ori_n109_));
  NA2        o087(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n110_));
  OAI210     o088(.A0(ori_ori_n74_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n111_), .B(ori_ori_n110_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n114_));
  AOI210     o092(.A0(ori_ori_n114_), .A1(ori_ori_n49_), .B0(ori_ori_n113_), .Y(ori_ori_n115_));
  AN2        o093(.A(ori_ori_n115_), .B(ori_ori_n112_), .Y(ori_ori_n116_));
  NO2        o094(.A(x09), .B(x05), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n117_), .B(ori_ori_n47_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n93_), .B(ori_ori_n49_), .Y(ori_ori_n119_));
  NA2        o097(.A(x09), .B(x00), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n119_), .B(ori_ori_n116_), .Y(ori_ori_n121_));
  NO2        o099(.A(x03), .B(x02), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n75_), .B(ori_ori_n90_), .Y(ori_ori_n123_));
  OAI210     o101(.A0(ori_ori_n123_), .A1(ori_ori_n95_), .B0(ori_ori_n122_), .Y(ori_ori_n124_));
  OA210      o102(.A0(ori_ori_n121_), .A1(x11), .B0(ori_ori_n124_), .Y(ori_ori_n125_));
  OAI210     o103(.A0(ori_ori_n109_), .A1(ori_ori_n23_), .B0(ori_ori_n125_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n93_), .B(ori_ori_n40_), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n127_), .B(ori_ori_n41_), .Y(ori_ori_n128_));
  NO2        o106(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n90_), .B(x01), .Y(ori_ori_n130_));
  AOI210     o108(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n128_), .B(ori_ori_n131_), .Y(ori_ori_n132_));
  NA2        o110(.A(x10), .B(x05), .Y(ori_ori_n133_));
  NO2        o111(.A(x09), .B(x01), .Y(ori_ori_n134_));
  INV        o112(.A(ori_ori_n25_), .Y(ori_ori_n135_));
  NAi21      o113(.An(x13), .B(x00), .Y(ori_ori_n136_));
  AN2        o114(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n84_), .B(x06), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n136_), .B(ori_ori_n36_), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n138_), .B(ori_ori_n137_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n140_), .B(ori_ori_n135_), .Y(ori_ori_n141_));
  NOi21      o119(.An(x09), .B(x00), .Y(ori_ori_n142_));
  NO3        o120(.A(ori_ori_n73_), .B(ori_ori_n142_), .C(ori_ori_n47_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(ori_ori_n101_), .Y(ori_ori_n144_));
  NA2        o122(.A(x06), .B(x05), .Y(ori_ori_n145_));
  OAI210     o123(.A0(ori_ori_n145_), .A1(ori_ori_n35_), .B0(ori_ori_n89_), .Y(ori_ori_n146_));
  AOI210     o124(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n146_), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n147_), .B(ori_ori_n144_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n90_), .B(x12), .Y(ori_ori_n149_));
  AOI210     o127(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o128(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n151_));
  NA2        o129(.A(ori_ori_n151_), .B(x02), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n150_), .B(ori_ori_n148_), .Y(ori_ori_n153_));
  NA3        o131(.A(ori_ori_n153_), .B(ori_ori_n141_), .C(ori_ori_n132_), .Y(ori_ori_n154_));
  AOI210     o132(.A0(ori_ori_n126_), .A1(ori_ori_n89_), .B0(ori_ori_n154_), .Y(ori_ori_n155_));
  INV        o133(.A(ori_ori_n66_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n156_), .B(ori_ori_n112_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n100_), .B(x06), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n158_), .Y(ori_ori_n159_));
  AOI210     o137(.A0(ori_ori_n159_), .A1(ori_ori_n157_), .B0(x12), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n83_), .B(x06), .Y(ori_ori_n161_));
  AOI210     o139(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n162_));
  NO3        o140(.A(ori_ori_n162_), .B(ori_ori_n161_), .C(ori_ori_n41_), .Y(ori_ori_n163_));
  INV        o141(.A(ori_ori_n114_), .Y(ori_ori_n164_));
  OAI210     o142(.A0(ori_ori_n164_), .A1(ori_ori_n163_), .B0(x02), .Y(ori_ori_n165_));
  AOI210     o143(.A0(ori_ori_n165_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n166_));
  OAI210     o144(.A0(ori_ori_n160_), .A1(ori_ori_n53_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  INV        o145(.A(ori_ori_n114_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n90_), .B(x03), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n68_), .B(ori_ori_n169_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n172_));
  NOi21      o150(.An(x13), .B(x04), .Y(ori_ori_n173_));
  NO3        o151(.A(ori_ori_n173_), .B(ori_ori_n68_), .C(ori_ori_n142_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n174_), .B(x05), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n172_), .Y(ori_ori_n176_));
  OAI210     o154(.A0(ori_ori_n171_), .A1(ori_ori_n168_), .B0(ori_ori_n176_), .Y(ori_ori_n177_));
  INV        o155(.A(ori_ori_n80_), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n179_));
  NO2        o157(.A(x06), .B(x00), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n181_));
  NA2        o159(.A(x13), .B(ori_ori_n89_), .Y(ori_ori_n182_));
  NA3        o160(.A(ori_ori_n182_), .B(ori_ori_n146_), .C(ori_ori_n81_), .Y(ori_ori_n183_));
  OAI210     o161(.A0(ori_ori_n317_), .A1(ori_ori_n179_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  AOI210     o162(.A0(ori_ori_n80_), .A1(ori_ori_n177_), .B0(ori_ori_n184_), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n185_), .A1(ori_ori_n167_), .B0(x07), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n64_), .B(ori_ori_n29_), .Y(ori_ori_n187_));
  NOi31      o165(.An(ori_ori_n110_), .B(ori_ori_n173_), .C(ori_ori_n142_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n188_), .B(ori_ori_n187_), .Y(ori_ori_n189_));
  OAI210     o167(.A0(ori_ori_n68_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n190_));
  INV        o168(.A(ori_ori_n190_), .Y(ori_ori_n191_));
  NO2        o169(.A(x12), .B(x02), .Y(ori_ori_n192_));
  INV        o170(.A(ori_ori_n192_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n193_), .B(ori_ori_n178_), .Y(ori_ori_n194_));
  OA210      o172(.A0(ori_ori_n191_), .A1(ori_ori_n189_), .B0(ori_ori_n194_), .Y(ori_ori_n195_));
  NA2        o173(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n196_), .B(x01), .Y(ori_ori_n197_));
  INV        o175(.A(ori_ori_n197_), .Y(ori_ori_n198_));
  AOI210     o176(.A0(ori_ori_n198_), .A1(ori_ori_n105_), .B0(ori_ori_n29_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n90_), .B(x04), .Y(ori_ori_n200_));
  NO3        o178(.A(ori_ori_n79_), .B(x12), .C(x03), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n199_), .B(ori_ori_n201_), .Y(ori_ori_n202_));
  NOi21      o180(.An(ori_ori_n187_), .B(ori_ori_n161_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n204_));
  NA2        o182(.A(ori_ori_n203_), .B(ori_ori_n204_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(ori_ori_n138_), .Y(ori_ori_n207_));
  NO2        o185(.A(ori_ori_n179_), .B(ori_ori_n28_), .Y(ori_ori_n208_));
  NA2        o186(.A(ori_ori_n207_), .B(ori_ori_n208_), .Y(ori_ori_n209_));
  NA3        o187(.A(ori_ori_n209_), .B(ori_ori_n205_), .C(ori_ori_n202_), .Y(ori_ori_n210_));
  NO3        o188(.A(ori_ori_n210_), .B(ori_ori_n195_), .C(ori_ori_n186_), .Y(ori_ori_n211_));
  OAI210     o189(.A0(ori_ori_n155_), .A1(ori_ori_n57_), .B0(ori_ori_n211_), .Y(ori02));
  AOI210     o190(.A0(ori_ori_n110_), .A1(ori_ori_n75_), .B0(ori_ori_n103_), .Y(ori_ori_n213_));
  NOi21      o191(.An(ori_ori_n174_), .B(ori_ori_n134_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n214_), .B(ori_ori_n32_), .Y(ori_ori_n215_));
  OAI210     o193(.A0(ori_ori_n215_), .A1(ori_ori_n213_), .B0(ori_ori_n133_), .Y(ori_ori_n216_));
  INV        o194(.A(ori_ori_n133_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n315_), .B(ori_ori_n162_), .Y(ori_ori_n218_));
  OAI220     o196(.A0(ori_ori_n218_), .A1(ori_ori_n90_), .B0(ori_ori_n75_), .B1(ori_ori_n50_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n219_), .B(ori_ori_n217_), .Y(ori_ori_n220_));
  AOI210     o198(.A0(ori_ori_n220_), .A1(ori_ori_n216_), .B0(ori_ori_n48_), .Y(ori_ori_n221_));
  NAi21      o199(.An(ori_ori_n175_), .B(ori_ori_n171_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n181_), .B(ori_ori_n47_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  OAI210     o202(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n313_), .B(ori_ori_n225_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n226_), .B(ori_ori_n84_), .Y(ori_ori_n227_));
  INV        o205(.A(ori_ori_n122_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n228_), .B(ori_ori_n102_), .Y(ori_ori_n229_));
  NA2        o207(.A(ori_ori_n229_), .B(x13), .Y(ori_ori_n230_));
  NA3        o208(.A(ori_ori_n230_), .B(ori_ori_n227_), .C(ori_ori_n224_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n231_), .B(ori_ori_n221_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n113_), .B(x03), .Y(ori_ori_n233_));
  INV        o211(.A(ori_ori_n136_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n35_), .B(ori_ori_n36_), .Y(ori_ori_n235_));
  AOI220     o213(.A0(ori_ori_n235_), .A1(ori_ori_n234_), .B0(ori_ori_n151_), .B1(x08), .Y(ori_ori_n236_));
  OAI210     o214(.A0(ori_ori_n236_), .A1(ori_ori_n206_), .B0(ori_ori_n233_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n237_), .B(ori_ori_n91_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n200_), .B(ori_ori_n89_), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n89_), .B(ori_ori_n41_), .Y(ori_ori_n240_));
  NA3        o218(.A(ori_ori_n240_), .B(ori_ori_n239_), .C(ori_ori_n102_), .Y(ori_ori_n241_));
  NA3        o219(.A(ori_ori_n241_), .B(ori_ori_n238_), .C(ori_ori_n48_), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n151_), .Y(ori_ori_n243_));
  OAI220     o221(.A0(ori_ori_n314_), .A1(ori_ori_n31_), .B0(ori_ori_n243_), .B1(ori_ori_n55_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n244_), .B(x02), .Y(ori_ori_n245_));
  NO3        o223(.A(ori_ori_n149_), .B(ori_ori_n129_), .C(ori_ori_n51_), .Y(ori_ori_n246_));
  OAI210     o224(.A0(ori_ori_n120_), .A1(ori_ori_n36_), .B0(ori_ori_n89_), .Y(ori_ori_n247_));
  OAI210     o225(.A0(ori_ori_n247_), .A1(ori_ori_n143_), .B0(ori_ori_n246_), .Y(ori_ori_n248_));
  NA3        o226(.A(ori_ori_n248_), .B(ori_ori_n245_), .C(x06), .Y(ori_ori_n249_));
  NO3        o227(.A(ori_ori_n206_), .B(ori_ori_n100_), .C(x08), .Y(ori_ori_n250_));
  INV        o228(.A(ori_ori_n250_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n252_));
  NO3        o230(.A(ori_ori_n94_), .B(ori_ori_n101_), .C(ori_ori_n38_), .Y(ori_ori_n253_));
  AOI210     o231(.A0(ori_ori_n246_), .A1(ori_ori_n252_), .B0(ori_ori_n253_), .Y(ori_ori_n254_));
  OAI210     o232(.A0(ori_ori_n251_), .A1(ori_ori_n28_), .B0(ori_ori_n254_), .Y(ori_ori_n255_));
  AN2        o233(.A(ori_ori_n255_), .B(x04), .Y(ori_ori_n256_));
  AOI210     o234(.A0(ori_ori_n249_), .A1(ori_ori_n242_), .B0(ori_ori_n256_), .Y(ori_ori_n257_));
  OAI210     o235(.A0(ori_ori_n232_), .A1(x12), .B0(ori_ori_n257_), .Y(ori03));
  OR2        o236(.A(ori_ori_n42_), .B(ori_ori_n169_), .Y(ori_ori_n259_));
  AOI210     o237(.A0(ori_ori_n123_), .A1(ori_ori_n89_), .B0(ori_ori_n259_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n149_), .B(ori_ori_n122_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n261_), .B(ori_ori_n152_), .Y(ori_ori_n262_));
  OAI210     o240(.A0(ori_ori_n262_), .A1(ori_ori_n260_), .B0(x05), .Y(ori_ori_n263_));
  AOI210     o241(.A0(ori_ori_n170_), .A1(ori_ori_n41_), .B0(ori_ori_n97_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n264_), .B(ori_ori_n55_), .Y(ori_ori_n265_));
  NA2        o243(.A(ori_ori_n265_), .B(ori_ori_n89_), .Y(ori_ori_n266_));
  AOI210     o244(.A0(ori_ori_n118_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n316_), .B(ori_ori_n37_), .Y(ori_ori_n268_));
  OAI210     o246(.A0(ori_ori_n268_), .A1(ori_ori_n267_), .B0(x04), .Y(ori_ori_n269_));
  NO3        o247(.A(ori_ori_n240_), .B(ori_ori_n75_), .C(ori_ori_n55_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n89_), .B(ori_ori_n118_), .Y(ori_ori_n271_));
  NO3        o249(.A(ori_ori_n106_), .B(ori_ori_n271_), .C(ori_ori_n270_), .Y(ori_ori_n272_));
  NA4        o250(.A(ori_ori_n272_), .B(ori_ori_n269_), .C(ori_ori_n266_), .D(ori_ori_n263_), .Y(ori04));
  NO2        o251(.A(ori_ori_n78_), .B(ori_ori_n39_), .Y(ori_ori_n274_));
  XO2        o252(.A(ori_ori_n274_), .B(ori_ori_n182_), .Y(ori05));
  INV        o253(.A(ori_ori_n25_), .Y(ori_ori_n276_));
  AOI210     o254(.A0(x06), .A1(ori_ori_n29_), .B0(ori_ori_n24_), .Y(ori_ori_n277_));
  OAI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n276_), .B0(ori_ori_n89_), .Y(ori_ori_n278_));
  OAI210     o256(.A0(ori_ori_n26_), .A1(ori_ori_n89_), .B0(x07), .Y(ori_ori_n279_));
  INV        o257(.A(ori_ori_n279_), .Y(ori_ori_n280_));
  AOI210     o258(.A0(ori_ori_n71_), .A1(ori_ori_n31_), .B0(ori_ori_n51_), .Y(ori_ori_n281_));
  NO3        o259(.A(ori_ori_n281_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n282_));
  BUFFER     o260(.A(ori_ori_n179_), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n180_), .B(ori_ori_n178_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n284_), .B(ori_ori_n283_), .Y(ori_ori_n285_));
  OAI210     o263(.A0(ori_ori_n285_), .A1(ori_ori_n282_), .B0(ori_ori_n89_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n33_), .B(ori_ori_n89_), .Y(ori_ori_n287_));
  AOI210     o265(.A0(ori_ori_n287_), .A1(ori_ori_n80_), .B0(x07), .Y(ori_ori_n288_));
  AOI220     o266(.A0(ori_ori_n288_), .A1(ori_ori_n286_), .B0(ori_ori_n280_), .B1(ori_ori_n278_), .Y(ori_ori_n289_));
  NOi21      o267(.An(ori_ori_n233_), .B(ori_ori_n106_), .Y(ori_ori_n290_));
  NO2        o268(.A(ori_ori_n290_), .B(ori_ori_n193_), .Y(ori_ori_n291_));
  OAI210     o269(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n292_));
  AOI210     o270(.A0(ori_ori_n182_), .A1(ori_ori_n47_), .B0(ori_ori_n292_), .Y(ori_ori_n293_));
  NO3        o271(.A(ori_ori_n293_), .B(ori_ori_n291_), .C(x08), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n103_), .B(ori_ori_n28_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n295_), .B(ori_ori_n197_), .Y(ori_ori_n296_));
  OR3        o274(.A(ori_ori_n296_), .B(x12), .C(x03), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n297_), .B(x08), .Y(ori_ori_n298_));
  INV        o276(.A(ori_ori_n298_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n294_), .B(ori_ori_n299_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n117_), .B(ori_ori_n43_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n301_), .B(ori_ori_n139_), .Y(ori_ori_n302_));
  NA3        o280(.A(ori_ori_n296_), .B(ori_ori_n290_), .C(ori_ori_n239_), .Y(ori_ori_n303_));
  INV        o281(.A(x14), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n130_), .B(ori_ori_n53_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n305_), .B(ori_ori_n304_), .Y(ori_ori_n306_));
  NA3        o284(.A(ori_ori_n306_), .B(ori_ori_n303_), .C(ori_ori_n302_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n287_), .B(ori_ori_n57_), .Y(ori_ori_n308_));
  NO2        o286(.A(ori_ori_n308_), .B(ori_ori_n79_), .Y(ori_ori_n309_));
  NO4        o287(.A(ori_ori_n309_), .B(ori_ori_n307_), .C(ori_ori_n300_), .D(ori_ori_n289_), .Y(ori06));
  INV        o288(.A(x13), .Y(ori_ori_n313_));
  INV        o289(.A(x05), .Y(ori_ori_n314_));
  INV        o290(.A(x02), .Y(ori_ori_n315_));
  INV        o291(.A(ori_ori_n134_), .Y(ori_ori_n316_));
  INV        o292(.A(ori_ori_n181_), .Y(ori_ori_n317_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NO3        m026(.A(x06), .B(x11), .C(x09), .Y(mai_mai_n49_));
  INV        m027(.A(x09), .Y(mai_mai_n50_));
  NO2        m028(.A(x10), .B(x02), .Y(mai_mai_n51_));
  NO2        m029(.A(x09), .B(x07), .Y(mai_mai_n52_));
  OAI210     m030(.A0(mai_mai_n52_), .A1(mai_mai_n49_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NOi21      m031(.An(x01), .B(x09), .Y(mai_mai_n54_));
  INV        m032(.A(x00), .Y(mai_mai_n55_));
  NO2        m033(.A(mai_mai_n50_), .B(mai_mai_n55_), .Y(mai_mai_n56_));
  NO2        m034(.A(mai_mai_n56_), .B(mai_mai_n54_), .Y(mai_mai_n57_));
  NA2        m035(.A(x09), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  INV        m036(.A(x07), .Y(mai_mai_n59_));
  INV        m037(.A(mai_mai_n57_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n61_), .B(mai_mai_n24_), .Y(mai_mai_n62_));
  NO2        m040(.A(mai_mai_n62_), .B(mai_mai_n60_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n63_), .B(mai_mai_n31_), .Y(mai_mai_n64_));
  AOI210     m042(.A0(mai_mai_n64_), .A1(mai_mai_n53_), .B0(x05), .Y(mai_mai_n65_));
  NA2        m043(.A(x09), .B(x05), .Y(mai_mai_n66_));
  NA2        m044(.A(x10), .B(x06), .Y(mai_mai_n67_));
  NA2        m045(.A(x07), .B(x03), .Y(mai_mai_n68_));
  NOi31      m046(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n69_));
  NO2        m047(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n70_), .B(mai_mai_n36_), .Y(mai_mai_n71_));
  OAI210     m049(.A0(mai_mai_n70_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n72_));
  AOI210     m050(.A0(mai_mai_n71_), .A1(mai_mai_n48_), .B0(mai_mai_n72_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n74_));
  NO2        m052(.A(x08), .B(x01), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n35_), .Y(mai_mai_n76_));
  NA2        m054(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n76_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  AN2        m056(.A(mai_mai_n78_), .B(mai_mai_n68_), .Y(mai_mai_n79_));
  INV        m057(.A(mai_mai_n76_), .Y(mai_mai_n80_));
  NO2        m058(.A(x06), .B(x05), .Y(mai_mai_n81_));
  NA2        m059(.A(x11), .B(x00), .Y(mai_mai_n82_));
  NO2        m060(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n83_));
  NOi21      m061(.An(mai_mai_n82_), .B(mai_mai_n83_), .Y(mai_mai_n84_));
  NOi21      m062(.An(x01), .B(x10), .Y(mai_mai_n85_));
  NO2        m063(.A(mai_mai_n29_), .B(mai_mai_n55_), .Y(mai_mai_n86_));
  NO3        m064(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(x06), .Y(mai_mai_n87_));
  NA2        m065(.A(mai_mai_n87_), .B(mai_mai_n27_), .Y(mai_mai_n88_));
  OAI210     m066(.A0(mai_mai_n364_), .A1(x07), .B0(mai_mai_n88_), .Y(mai_mai_n89_));
  NO3        m067(.A(mai_mai_n89_), .B(mai_mai_n79_), .C(mai_mai_n65_), .Y(mai01));
  INV        m068(.A(x12), .Y(mai_mai_n91_));
  INV        m069(.A(x13), .Y(mai_mai_n92_));
  NA2        m070(.A(x08), .B(x04), .Y(mai_mai_n93_));
  NA2        m071(.A(x08), .B(mai_mai_n81_), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n85_), .B(mai_mai_n28_), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n95_), .B(mai_mai_n66_), .Y(mai_mai_n96_));
  NO2        m074(.A(x10), .B(x01), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n98_));
  NO2        m076(.A(mai_mai_n98_), .B(mai_mai_n97_), .Y(mai_mai_n99_));
  NO3        m077(.A(x02), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n100_));
  AOI210     m078(.A0(mai_mai_n100_), .A1(mai_mai_n99_), .B0(mai_mai_n96_), .Y(mai_mai_n101_));
  AOI210     m079(.A0(mai_mai_n101_), .A1(mai_mai_n94_), .B0(mai_mai_n92_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n54_), .B(x05), .Y(mai_mai_n103_));
  NOi21      m081(.An(mai_mai_n103_), .B(mai_mai_n56_), .Y(mai_mai_n104_));
  INV        m082(.A(x02), .Y(mai_mai_n105_));
  NA3        m083(.A(x13), .B(mai_mai_n105_), .C(x06), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(mai_mai_n104_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n75_), .B(x13), .Y(mai_mai_n108_));
  NA2        m086(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NA2        m088(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n111_), .B(x05), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(mai_mai_n110_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n35_), .B(mai_mai_n55_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n114_), .B(mai_mai_n92_), .Y(mai_mai_n115_));
  AOI210     m093(.A0(mai_mai_n115_), .A1(mai_mai_n71_), .B0(mai_mai_n104_), .Y(mai_mai_n116_));
  AOI210     m094(.A0(mai_mai_n116_), .A1(mai_mai_n113_), .B0(mai_mai_n67_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n118_));
  NA2        m096(.A(x10), .B(mai_mai_n55_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n50_), .B(x05), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n122_));
  NO3        m100(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n123_));
  NO4        m101(.A(mai_mai_n123_), .B(mai_mai_n117_), .C(mai_mai_n107_), .D(mai_mai_n102_), .Y(mai_mai_n124_));
  OAI210     m102(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n125_));
  NO2        m103(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n127_));
  NO2        m105(.A(x09), .B(x05), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n47_), .Y(mai_mai_n129_));
  AOI210     m107(.A0(mai_mai_n129_), .A1(mai_mai_n99_), .B0(x06), .Y(mai_mai_n130_));
  NA2        m108(.A(x09), .B(x00), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n103_), .B(mai_mai_n131_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n69_), .B(mai_mai_n50_), .Y(mai_mai_n133_));
  AOI210     m111(.A0(mai_mai_n133_), .A1(mai_mai_n132_), .B0(mai_mai_n127_), .Y(mai_mai_n134_));
  NO2        m112(.A(mai_mai_n134_), .B(mai_mai_n130_), .Y(mai_mai_n135_));
  NO2        m113(.A(x03), .B(x02), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n76_), .B(mai_mai_n92_), .Y(mai_mai_n137_));
  OAI210     m115(.A0(mai_mai_n137_), .A1(mai_mai_n104_), .B0(mai_mai_n136_), .Y(mai_mai_n138_));
  OA210      m116(.A0(mai_mai_n135_), .A1(x11), .B0(mai_mai_n138_), .Y(mai_mai_n139_));
  OAI210     m117(.A0(mai_mai_n124_), .A1(mai_mai_n23_), .B0(mai_mai_n139_), .Y(mai_mai_n140_));
  NAi21      m118(.An(x06), .B(x10), .Y(mai_mai_n141_));
  INV        m119(.A(x01), .Y(mai_mai_n142_));
  BUFFER     m120(.A(mai_mai_n142_), .Y(mai_mai_n143_));
  AOI210     m121(.A0(mai_mai_n143_), .A1(mai_mai_n368_), .B0(mai_mai_n41_), .Y(mai_mai_n144_));
  NO2        m122(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n92_), .B(x01), .Y(mai_mai_n146_));
  NO2        m124(.A(mai_mai_n146_), .B(x08), .Y(mai_mai_n147_));
  AOI210     m125(.A0(x09), .A1(mai_mai_n145_), .B0(mai_mai_n48_), .Y(mai_mai_n148_));
  AOI210     m126(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n148_), .A1(mai_mai_n144_), .B0(mai_mai_n149_), .Y(mai_mai_n150_));
  NA2        m128(.A(x04), .B(x02), .Y(mai_mai_n151_));
  NA2        m129(.A(x10), .B(x05), .Y(mai_mai_n152_));
  INV        m130(.A(x03), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n103_), .B(x08), .Y(mai_mai_n154_));
  OAI210     m132(.A0(mai_mai_n363_), .A1(x11), .B0(mai_mai_n153_), .Y(mai_mai_n155_));
  NAi21      m133(.An(mai_mai_n151_), .B(mai_mai_n155_), .Y(mai_mai_n156_));
  INV        m134(.A(mai_mai_n25_), .Y(mai_mai_n157_));
  NAi21      m135(.An(x13), .B(x00), .Y(mai_mai_n158_));
  AOI210     m136(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n158_), .Y(mai_mai_n159_));
  AOI220     m137(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n160_));
  OAI210     m138(.A0(mai_mai_n152_), .A1(mai_mai_n35_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  AN2        m139(.A(mai_mai_n161_), .B(mai_mai_n159_), .Y(mai_mai_n162_));
  NO2        m140(.A(mai_mai_n158_), .B(mai_mai_n36_), .Y(mai_mai_n163_));
  OAI210     m141(.A0(mai_mai_n163_), .A1(mai_mai_n162_), .B0(mai_mai_n157_), .Y(mai_mai_n164_));
  NOi21      m142(.An(x09), .B(x00), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n92_), .B(x12), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n85_), .B(mai_mai_n50_), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n369_), .B(x12), .Y(mai_mai_n169_));
  NA4        m147(.A(mai_mai_n169_), .B(mai_mai_n164_), .C(mai_mai_n156_), .D(mai_mai_n150_), .Y(mai_mai_n170_));
  AOI210     m148(.A0(mai_mai_n140_), .A1(mai_mai_n91_), .B0(mai_mai_n170_), .Y(mai_mai_n171_));
  NA2        m149(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n172_));
  NA2        m150(.A(mai_mai_n172_), .B(mai_mai_n125_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n365_), .B(mai_mai_n173_), .Y(mai_mai_n174_));
  NO2        m152(.A(mai_mai_n174_), .B(x12), .Y(mai_mai_n175_));
  INV        m153(.A(mai_mai_n69_), .Y(mai_mai_n176_));
  NO2        m154(.A(x05), .B(mai_mai_n50_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n177_), .B(mai_mai_n55_), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n178_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n179_), .B(mai_mai_n23_), .Y(mai_mai_n180_));
  OAI210     m158(.A0(mai_mai_n175_), .A1(mai_mai_n55_), .B0(mai_mai_n180_), .Y(mai_mai_n181_));
  INV        m159(.A(mai_mai_n127_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n50_), .B(x03), .Y(mai_mai_n183_));
  OAI210     m161(.A0(mai_mai_n70_), .A1(mai_mai_n36_), .B0(mai_mai_n109_), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n92_), .B(x03), .Y(mai_mai_n185_));
  NA2        m163(.A(mai_mai_n185_), .B(mai_mai_n184_), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n141_), .Y(mai_mai_n187_));
  NOi21      m165(.An(x13), .B(x04), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n188_), .B(mai_mai_n165_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n187_), .B(mai_mai_n55_), .Y(mai_mai_n190_));
  OAI210     m168(.A0(mai_mai_n186_), .A1(mai_mai_n182_), .B0(mai_mai_n190_), .Y(mai_mai_n191_));
  INV        m169(.A(mai_mai_n83_), .Y(mai_mai_n192_));
  NO2        m170(.A(mai_mai_n192_), .B(x12), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n194_));
  NO2        m172(.A(mai_mai_n50_), .B(mai_mai_n36_), .Y(mai_mai_n195_));
  OAI210     m173(.A0(mai_mai_n195_), .A1(mai_mai_n161_), .B0(mai_mai_n159_), .Y(mai_mai_n196_));
  AOI210     m174(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n197_));
  NO2        m175(.A(x06), .B(x00), .Y(mai_mai_n198_));
  NO3        m176(.A(mai_mai_n198_), .B(mai_mai_n197_), .C(mai_mai_n41_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n93_), .B(mai_mai_n131_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n200_), .B(mai_mai_n199_), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n202_));
  NA2        m180(.A(mai_mai_n202_), .B(x03), .Y(mai_mai_n203_));
  OA210      m181(.A0(mai_mai_n203_), .A1(mai_mai_n201_), .B0(mai_mai_n196_), .Y(mai_mai_n204_));
  NA2        m182(.A(x13), .B(mai_mai_n91_), .Y(mai_mai_n205_));
  NA3        m183(.A(mai_mai_n205_), .B(x12), .C(mai_mai_n84_), .Y(mai_mai_n206_));
  OAI210     m184(.A0(mai_mai_n204_), .A1(mai_mai_n194_), .B0(mai_mai_n206_), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n193_), .A1(mai_mai_n191_), .B0(mai_mai_n207_), .Y(mai_mai_n208_));
  AOI210     m186(.A0(mai_mai_n208_), .A1(mai_mai_n181_), .B0(x07), .Y(mai_mai_n209_));
  NA2        m187(.A(mai_mai_n66_), .B(mai_mai_n29_), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n188_), .B(mai_mai_n165_), .Y(mai_mai_n211_));
  AOI210     m189(.A0(mai_mai_n211_), .A1(mai_mai_n133_), .B0(mai_mai_n210_), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n92_), .B(x06), .Y(mai_mai_n213_));
  INV        m191(.A(mai_mai_n213_), .Y(mai_mai_n214_));
  NO2        m192(.A(x08), .B(x05), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n215_), .B(mai_mai_n197_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n216_), .B(mai_mai_n214_), .Y(mai_mai_n217_));
  NO2        m195(.A(x12), .B(x02), .Y(mai_mai_n218_));
  INV        m196(.A(mai_mai_n218_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n219_), .B(mai_mai_n192_), .Y(mai_mai_n220_));
  OA210      m198(.A0(mai_mai_n217_), .A1(mai_mai_n212_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  NA2        m199(.A(mai_mai_n50_), .B(mai_mai_n41_), .Y(mai_mai_n222_));
  NOi21      m200(.An(mai_mai_n75_), .B(mai_mai_n109_), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n213_), .B(mai_mai_n184_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n92_), .B(x04), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n225_), .B(mai_mai_n28_), .Y(mai_mai_n226_));
  OAI210     m204(.A0(mai_mai_n226_), .A1(mai_mai_n108_), .B0(mai_mai_n224_), .Y(mai_mai_n227_));
  NO3        m205(.A(mai_mai_n82_), .B(x12), .C(x03), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n227_), .A1(mai_mai_n223_), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  INV        m207(.A(mai_mai_n167_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n231_));
  NA2        m209(.A(mai_mai_n230_), .B(mai_mai_n231_), .Y(mai_mai_n232_));
  NA2        m210(.A(mai_mai_n232_), .B(mai_mai_n229_), .Y(mai_mai_n233_));
  NO3        m211(.A(mai_mai_n233_), .B(mai_mai_n221_), .C(mai_mai_n209_), .Y(mai_mai_n234_));
  OAI210     m212(.A0(mai_mai_n171_), .A1(mai_mai_n59_), .B0(mai_mai_n234_), .Y(mai02));
  BUFFER     m213(.A(mai_mai_n189_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n92_), .B(mai_mai_n35_), .Y(mai_mai_n237_));
  NA3        m215(.A(mai_mai_n237_), .B(x10), .C(mai_mai_n54_), .Y(mai_mai_n238_));
  OAI210     m216(.A0(mai_mai_n236_), .A1(mai_mai_n32_), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NA2        m217(.A(mai_mai_n239_), .B(mai_mai_n152_), .Y(mai_mai_n240_));
  NO2        m218(.A(mai_mai_n76_), .B(mai_mai_n50_), .Y(mai_mai_n241_));
  AOI220     m219(.A0(mai_mai_n241_), .A1(x10), .B0(mai_mai_n137_), .B1(mai_mai_n136_), .Y(mai_mai_n242_));
  AOI210     m220(.A0(mai_mai_n242_), .A1(mai_mai_n240_), .B0(mai_mai_n48_), .Y(mai_mai_n243_));
  NO2        m221(.A(x05), .B(x02), .Y(mai_mai_n244_));
  OAI210     m222(.A0(mai_mai_n173_), .A1(mai_mai_n165_), .B0(mai_mai_n244_), .Y(mai_mai_n245_));
  AOI220     m223(.A0(mai_mai_n215_), .A1(mai_mai_n56_), .B0(mai_mai_n54_), .B1(mai_mai_n36_), .Y(mai_mai_n246_));
  NOi21      m224(.An(mai_mai_n237_), .B(mai_mai_n246_), .Y(mai_mai_n247_));
  AOI210     m225(.A0(mai_mai_n188_), .A1(mai_mai_n70_), .B0(mai_mai_n247_), .Y(mai_mai_n248_));
  AOI210     m226(.A0(mai_mai_n248_), .A1(mai_mai_n245_), .B0(mai_mai_n127_), .Y(mai_mai_n249_));
  INV        m227(.A(mai_mai_n186_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n202_), .B(mai_mai_n47_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  AN2        m230(.A(mai_mai_n185_), .B(mai_mai_n184_), .Y(mai_mai_n253_));
  OAI210     m231(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n254_));
  NA2        m232(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n255_));
  OA210      m233(.A0(mai_mai_n255_), .A1(x08), .B0(mai_mai_n129_), .Y(mai_mai_n256_));
  AOI210     m234(.A0(mai_mai_n256_), .A1(mai_mai_n125_), .B0(mai_mai_n254_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n257_), .A1(mai_mai_n253_), .B0(mai_mai_n86_), .Y(mai_mai_n258_));
  NA3        m236(.A(mai_mai_n86_), .B(mai_mai_n75_), .C(mai_mai_n183_), .Y(mai_mai_n259_));
  NA3        m237(.A(mai_mai_n85_), .B(mai_mai_n74_), .C(mai_mai_n42_), .Y(mai_mai_n260_));
  AOI210     m238(.A0(mai_mai_n260_), .A1(mai_mai_n259_), .B0(x04), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n216_), .B(mai_mai_n95_), .Y(mai_mai_n262_));
  AOI210     m240(.A0(mai_mai_n262_), .A1(x13), .B0(mai_mai_n261_), .Y(mai_mai_n263_));
  NA3        m241(.A(mai_mai_n263_), .B(mai_mai_n258_), .C(mai_mai_n252_), .Y(mai_mai_n264_));
  NO3        m242(.A(mai_mai_n264_), .B(mai_mai_n249_), .C(mai_mai_n243_), .Y(mai_mai_n265_));
  NA2        m243(.A(mai_mai_n126_), .B(x03), .Y(mai_mai_n266_));
  NA2        m244(.A(mai_mai_n168_), .B(mai_mai_n97_), .Y(mai_mai_n267_));
  INV        m245(.A(mai_mai_n54_), .Y(mai_mai_n268_));
  OAI220     m246(.A0(mai_mai_n225_), .A1(mai_mai_n268_), .B0(mai_mai_n121_), .B1(mai_mai_n28_), .Y(mai_mai_n269_));
  OAI210     m247(.A0(mai_mai_n269_), .A1(mai_mai_n154_), .B0(mai_mai_n98_), .Y(mai_mai_n270_));
  NA3        m248(.A(x12), .B(x12), .C(mai_mai_n120_), .Y(mai_mai_n271_));
  NA4        m249(.A(mai_mai_n271_), .B(mai_mai_n270_), .C(mai_mai_n267_), .D(mai_mai_n48_), .Y(mai_mai_n272_));
  INV        m250(.A(mai_mai_n168_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n147_), .B(mai_mai_n40_), .Y(mai_mai_n274_));
  NA2        m252(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n275_));
  OAI220     m253(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n273_), .B1(mai_mai_n57_), .Y(mai_mai_n276_));
  NA2        m254(.A(mai_mai_n276_), .B(x02), .Y(mai_mai_n277_));
  INV        m255(.A(mai_mai_n195_), .Y(mai_mai_n278_));
  NA2        m256(.A(mai_mai_n166_), .B(x04), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n279_), .B(mai_mai_n278_), .Y(mai_mai_n280_));
  NO2        m258(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n281_));
  OAI210     m259(.A0(mai_mai_n281_), .A1(mai_mai_n280_), .B0(mai_mai_n86_), .Y(mai_mai_n282_));
  NO3        m260(.A(mai_mai_n166_), .B(mai_mai_n145_), .C(mai_mai_n51_), .Y(mai_mai_n283_));
  OAI210     m261(.A0(mai_mai_n131_), .A1(mai_mai_n36_), .B0(mai_mai_n91_), .Y(mai_mai_n284_));
  NA2        m262(.A(mai_mai_n284_), .B(mai_mai_n283_), .Y(mai_mai_n285_));
  NA4        m263(.A(mai_mai_n285_), .B(mai_mai_n282_), .C(mai_mai_n277_), .D(x06), .Y(mai_mai_n286_));
  NA2        m264(.A(x09), .B(x03), .Y(mai_mai_n287_));
  OAI220     m265(.A0(mai_mai_n287_), .A1(mai_mai_n119_), .B0(mai_mai_n172_), .B1(mai_mai_n61_), .Y(mai_mai_n288_));
  OAI220     m266(.A0(mai_mai_n146_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n118_), .B(x08), .Y(mai_mai_n290_));
  AOI210     m268(.A0(mai_mai_n289_), .A1(mai_mai_n182_), .B0(mai_mai_n290_), .Y(mai_mai_n291_));
  NO3        m269(.A(mai_mai_n103_), .B(mai_mai_n119_), .C(mai_mai_n38_), .Y(mai_mai_n292_));
  INV        m270(.A(mai_mai_n292_), .Y(mai_mai_n293_));
  OAI210     m271(.A0(mai_mai_n291_), .A1(mai_mai_n28_), .B0(mai_mai_n293_), .Y(mai_mai_n294_));
  AO220      m272(.A0(mai_mai_n294_), .A1(x04), .B0(mai_mai_n288_), .B1(x05), .Y(mai_mai_n295_));
  AOI210     m273(.A0(mai_mai_n286_), .A1(mai_mai_n272_), .B0(mai_mai_n295_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n265_), .A1(x12), .B0(mai_mai_n296_), .Y(mai03));
  OR2        m275(.A(mai_mai_n42_), .B(mai_mai_n183_), .Y(mai_mai_n298_));
  AOI210     m276(.A0(mai_mai_n137_), .A1(mai_mai_n91_), .B0(mai_mai_n298_), .Y(mai_mai_n299_));
  AO210      m277(.A0(mai_mai_n278_), .A1(mai_mai_n77_), .B0(mai_mai_n279_), .Y(mai_mai_n300_));
  INV        m278(.A(mai_mai_n300_), .Y(mai_mai_n301_));
  OAI210     m279(.A0(mai_mai_n301_), .A1(mai_mai_n299_), .B0(x05), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n298_), .B(x05), .Y(mai_mai_n303_));
  AOI210     m281(.A0(mai_mai_n125_), .A1(mai_mai_n176_), .B0(mai_mai_n303_), .Y(mai_mai_n304_));
  AOI210     m282(.A0(mai_mai_n185_), .A1(mai_mai_n71_), .B0(mai_mai_n112_), .Y(mai_mai_n305_));
  OAI220     m283(.A0(mai_mai_n305_), .A1(mai_mai_n57_), .B0(mai_mai_n255_), .B1(mai_mai_n246_), .Y(mai_mai_n306_));
  OAI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n304_), .B0(mai_mai_n91_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n132_), .B(x13), .Y(mai_mai_n308_));
  NA2        m286(.A(mai_mai_n308_), .B(x04), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n158_), .A1(mai_mai_n91_), .B0(mai_mai_n129_), .Y(mai_mai_n310_));
  OA210      m288(.A0(mai_mai_n147_), .A1(x12), .B0(mai_mai_n122_), .Y(mai_mai_n311_));
  NO2        m289(.A(mai_mai_n311_), .B(mai_mai_n310_), .Y(mai_mai_n312_));
  NA4        m290(.A(mai_mai_n312_), .B(mai_mai_n309_), .C(mai_mai_n307_), .D(mai_mai_n302_), .Y(mai04));
  NO2        m291(.A(mai_mai_n80_), .B(mai_mai_n39_), .Y(mai_mai_n314_));
  XO2        m292(.A(mai_mai_n314_), .B(mai_mai_n205_), .Y(mai05));
  NA2        m293(.A(mai_mai_n121_), .B(mai_mai_n31_), .Y(mai_mai_n316_));
  NA2        m294(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n317_));
  NA2        m295(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n317_), .A1(mai_mai_n72_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  AOI210     m297(.A0(mai_mai_n319_), .A1(x06), .B0(mai_mai_n367_), .Y(mai_mai_n320_));
  NA2        m298(.A(x01), .B(x05), .Y(mai_mai_n321_));
  NA2        m299(.A(mai_mai_n321_), .B(mai_mai_n198_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n322_), .B(mai_mai_n366_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n323_), .B(mai_mai_n91_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n83_), .B(x07), .Y(mai_mai_n325_));
  AOI220     m303(.A0(mai_mai_n325_), .A1(mai_mai_n324_), .B0(mai_mai_n320_), .B1(mai_mai_n316_), .Y(mai_mai_n326_));
  OR2        m304(.A(mai_mai_n222_), .B(mai_mai_n219_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(x11), .A1(x07), .B0(mai_mai_n126_), .Y(mai_mai_n328_));
  OR2        m306(.A(mai_mai_n328_), .B(x03), .Y(mai_mai_n329_));
  NO2        m307(.A(mai_mai_n128_), .B(mai_mai_n28_), .Y(mai_mai_n330_));
  AOI220     m308(.A0(mai_mai_n330_), .A1(mai_mai_n329_), .B0(mai_mai_n327_), .B1(mai_mai_n47_), .Y(mai_mai_n331_));
  NA2        m309(.A(mai_mai_n331_), .B(mai_mai_n92_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n279_), .A1(x02), .B0(mai_mai_n218_), .Y(mai_mai_n333_));
  NOi21      m311(.An(mai_mai_n266_), .B(mai_mai_n122_), .Y(mai_mai_n334_));
  NO2        m312(.A(mai_mai_n334_), .B(mai_mai_n219_), .Y(mai_mai_n335_));
  OAI210     m313(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n205_), .A1(mai_mai_n47_), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  NO4        m315(.A(mai_mai_n337_), .B(mai_mai_n335_), .C(mai_mai_n333_), .D(x08), .Y(mai_mai_n338_));
  NO2        m316(.A(x05), .B(x03), .Y(mai_mai_n339_));
  NO2        m317(.A(x13), .B(x12), .Y(mai_mai_n340_));
  OR3        m318(.A(x09), .B(x12), .C(x03), .Y(mai_mai_n341_));
  NA3        m319(.A(mai_mai_n273_), .B(mai_mai_n114_), .C(x12), .Y(mai_mai_n342_));
  AO210      m320(.A0(mai_mai_n273_), .A1(mai_mai_n114_), .B0(mai_mai_n205_), .Y(mai_mai_n343_));
  NA4        m321(.A(mai_mai_n343_), .B(mai_mai_n342_), .C(mai_mai_n341_), .D(x08), .Y(mai_mai_n344_));
  AOI210     m322(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(mai_mai_n344_), .Y(mai_mai_n345_));
  AOI210     m323(.A0(mai_mai_n338_), .A1(mai_mai_n332_), .B0(mai_mai_n345_), .Y(mai_mai_n346_));
  INV        m324(.A(x07), .Y(mai_mai_n347_));
  OAI220     m325(.A0(mai_mai_n347_), .A1(mai_mai_n318_), .B0(mai_mai_n128_), .B1(mai_mai_n43_), .Y(mai_mai_n348_));
  NA2        m326(.A(mai_mai_n348_), .B(mai_mai_n163_), .Y(mai_mai_n349_));
  INV        m327(.A(x14), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n95_), .B(x11), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n351_), .B(mai_mai_n350_), .Y(mai_mai_n352_));
  NA2        m330(.A(mai_mai_n352_), .B(mai_mai_n349_), .Y(mai_mai_n353_));
  NO2        m331(.A(mai_mai_n145_), .B(mai_mai_n59_), .Y(mai_mai_n354_));
  NOi21      m332(.An(mai_mai_n225_), .B(mai_mai_n132_), .Y(mai_mai_n355_));
  NA2        m333(.A(mai_mai_n231_), .B(mai_mai_n187_), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  OAI210     m335(.A0(mai_mai_n357_), .A1(mai_mai_n355_), .B0(mai_mai_n91_), .Y(mai_mai_n358_));
  OAI210     m336(.A0(mai_mai_n354_), .A1(mai_mai_n82_), .B0(mai_mai_n358_), .Y(mai_mai_n359_));
  NO4        m337(.A(mai_mai_n359_), .B(mai_mai_n353_), .C(mai_mai_n346_), .D(mai_mai_n326_), .Y(mai06));
  INV        m338(.A(x01), .Y(mai_mai_n363_));
  INV        m339(.A(mai_mai_n84_), .Y(mai_mai_n364_));
  INV        m340(.A(x05), .Y(mai_mai_n365_));
  INV        m341(.A(mai_mai_n213_), .Y(mai_mai_n366_));
  INV        m342(.A(x07), .Y(mai_mai_n367_));
  INV        m343(.A(mai_mai_n40_), .Y(mai_mai_n368_));
  INV        m344(.A(mai_mai_n25_), .Y(mai_mai_n369_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NO2        u026(.A(x02), .B(x11), .Y(men_men_n49_));
  INV        u027(.A(x09), .Y(men_men_n50_));
  NO2        u028(.A(x10), .B(x02), .Y(men_men_n51_));
  INV        u029(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u030(.A(men_men_n52_), .B(x07), .Y(men_men_n53_));
  OAI210     u031(.A0(men_men_n53_), .A1(men_men_n49_), .B0(men_men_n47_), .Y(men_men_n54_));
  NOi21      u032(.An(x01), .B(x09), .Y(men_men_n55_));
  INV        u033(.A(x00), .Y(men_men_n56_));
  NO2        u034(.A(men_men_n50_), .B(men_men_n56_), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n57_), .B(men_men_n55_), .Y(men_men_n58_));
  NA2        u036(.A(x09), .B(men_men_n56_), .Y(men_men_n59_));
  INV        u037(.A(x07), .Y(men_men_n60_));
  AOI210     u038(.A0(x11), .A1(men_men_n48_), .B0(men_men_n60_), .Y(men_men_n61_));
  INV        u039(.A(men_men_n58_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n29_), .B(x02), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n24_), .Y(men_men_n64_));
  OAI220     u042(.A0(men_men_n64_), .A1(men_men_n62_), .B0(men_men_n61_), .B1(men_men_n59_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n60_), .B(men_men_n48_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n30_), .A1(x11), .B0(men_men_n66_), .Y(men_men_n67_));
  AOI220     u045(.A0(men_men_n67_), .A1(men_men_n58_), .B0(men_men_n65_), .B1(men_men_n31_), .Y(men_men_n68_));
  AOI210     u046(.A0(men_men_n68_), .A1(men_men_n54_), .B0(x05), .Y(men_men_n69_));
  NA2        u047(.A(x10), .B(x09), .Y(men_men_n70_));
  NA2        u048(.A(x09), .B(x05), .Y(men_men_n71_));
  NA2        u049(.A(x10), .B(x06), .Y(men_men_n72_));
  NA3        u050(.A(men_men_n72_), .B(men_men_n71_), .C(men_men_n28_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n60_), .B(men_men_n41_), .Y(men_men_n74_));
  OAI210     u052(.A0(men_men_n73_), .A1(x11), .B0(x03), .Y(men_men_n75_));
  NOi31      u053(.An(x08), .B(x04), .C(x00), .Y(men_men_n76_));
  NO2        u054(.A(x10), .B(x09), .Y(men_men_n77_));
  NO2        u055(.A(x09), .B(men_men_n41_), .Y(men_men_n78_));
  OAI210     u056(.A0(men_men_n78_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n36_), .B(x00), .Y(men_men_n80_));
  NO2        u058(.A(x08), .B(x01), .Y(men_men_n81_));
  OAI210     u059(.A0(men_men_n81_), .A1(men_men_n80_), .B0(men_men_n35_), .Y(men_men_n82_));
  NA2        u060(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n83_));
  NO2        u061(.A(men_men_n82_), .B(x02), .Y(men_men_n84_));
  AN2        u062(.A(men_men_n84_), .B(men_men_n75_), .Y(men_men_n85_));
  INV        u063(.A(men_men_n82_), .Y(men_men_n86_));
  NO2        u064(.A(x06), .B(x05), .Y(men_men_n87_));
  NA2        u065(.A(x11), .B(x00), .Y(men_men_n88_));
  NO2        u066(.A(x11), .B(men_men_n47_), .Y(men_men_n89_));
  NOi21      u067(.An(men_men_n88_), .B(men_men_n89_), .Y(men_men_n90_));
  AOI210     u068(.A0(men_men_n87_), .A1(men_men_n86_), .B0(men_men_n90_), .Y(men_men_n91_));
  NOi21      u069(.An(x01), .B(x10), .Y(men_men_n92_));
  NO2        u070(.A(men_men_n29_), .B(men_men_n56_), .Y(men_men_n93_));
  NO3        u071(.A(men_men_n93_), .B(men_men_n92_), .C(x06), .Y(men_men_n94_));
  NA2        u072(.A(men_men_n94_), .B(men_men_n27_), .Y(men_men_n95_));
  OAI210     u073(.A0(men_men_n91_), .A1(x07), .B0(men_men_n95_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n85_), .C(men_men_n69_), .Y(men01));
  INV        u075(.A(x12), .Y(men_men_n98_));
  INV        u076(.A(x13), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n384_), .B(men_men_n70_), .Y(men_men_n100_));
  NA2        u078(.A(x08), .B(x04), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n101_), .B(men_men_n56_), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n102_), .B(men_men_n100_), .Y(men_men_n103_));
  NA2        u081(.A(men_men_n92_), .B(men_men_n28_), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n71_), .Y(men_men_n105_));
  NO2        u083(.A(x10), .B(x01), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n29_), .B(x00), .Y(men_men_n107_));
  NA2        u085(.A(x04), .B(men_men_n28_), .Y(men_men_n108_));
  NO3        u086(.A(men_men_n108_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n105_), .Y(men_men_n110_));
  AOI210     u088(.A0(men_men_n110_), .A1(men_men_n103_), .B0(men_men_n99_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n55_), .B(x05), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n35_), .B(x02), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n99_), .B(men_men_n36_), .Y(men_men_n114_));
  NA3        u092(.A(men_men_n114_), .B(men_men_n113_), .C(x06), .Y(men_men_n115_));
  INV        u093(.A(men_men_n115_), .Y(men_men_n116_));
  NA2        u094(.A(men_men_n35_), .B(men_men_n56_), .Y(men_men_n117_));
  INV        u095(.A(men_men_n72_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n119_));
  NA2        u097(.A(x10), .B(men_men_n56_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NA2        u099(.A(men_men_n50_), .B(x05), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n36_), .B(x04), .Y(men_men_n123_));
  NA3        u101(.A(men_men_n123_), .B(men_men_n122_), .C(x13), .Y(men_men_n124_));
  NO3        u102(.A(men_men_n117_), .B(men_men_n78_), .C(men_men_n36_), .Y(men_men_n125_));
  NO2        u103(.A(men_men_n59_), .B(x05), .Y(men_men_n126_));
  NOi41      u104(.An(men_men_n124_), .B(men_men_n126_), .C(men_men_n125_), .D(men_men_n121_), .Y(men_men_n127_));
  NO3        u105(.A(men_men_n127_), .B(x06), .C(x03), .Y(men_men_n128_));
  NO4        u106(.A(men_men_n128_), .B(men_men_n118_), .C(men_men_n116_), .D(men_men_n111_), .Y(men_men_n129_));
  NO2        u107(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n130_));
  OA210      u108(.A0(x00), .A1(men_men_n77_), .B0(men_men_n130_), .Y(men_men_n131_));
  NO2        u109(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n29_), .B(x06), .Y(men_men_n133_));
  OA210      u111(.A0(men_men_n28_), .A1(men_men_n131_), .B0(men_men_n386_), .Y(men_men_n134_));
  NO2        u112(.A(x09), .B(x05), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(men_men_n47_), .Y(men_men_n136_));
  NA2        u114(.A(x09), .B(x00), .Y(men_men_n137_));
  NA2        u115(.A(men_men_n112_), .B(men_men_n137_), .Y(men_men_n138_));
  NO2        u116(.A(men_men_n28_), .B(men_men_n134_), .Y(men_men_n139_));
  NO2        u117(.A(x03), .B(x02), .Y(men_men_n140_));
  OR2        u118(.A(men_men_n139_), .B(x11), .Y(men_men_n141_));
  OAI210     u119(.A0(men_men_n129_), .A1(men_men_n23_), .B0(men_men_n141_), .Y(men_men_n142_));
  NAi21      u120(.An(x06), .B(x10), .Y(men_men_n143_));
  NOi21      u121(.An(x01), .B(x13), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n144_), .B(men_men_n143_), .Y(men_men_n145_));
  OR2        u123(.A(men_men_n145_), .B(x08), .Y(men_men_n146_));
  NO2        u124(.A(men_men_n146_), .B(men_men_n41_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n29_), .B(x03), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n99_), .B(x01), .Y(men_men_n149_));
  NO2        u127(.A(men_men_n149_), .B(x08), .Y(men_men_n150_));
  OAI210     u128(.A0(x05), .A1(men_men_n150_), .B0(men_men_n50_), .Y(men_men_n151_));
  AOI210     u129(.A0(men_men_n151_), .A1(men_men_n148_), .B0(men_men_n48_), .Y(men_men_n152_));
  AOI210     u130(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n153_));
  OAI210     u131(.A0(men_men_n152_), .A1(men_men_n147_), .B0(men_men_n153_), .Y(men_men_n154_));
  NA2        u132(.A(x04), .B(x02), .Y(men_men_n155_));
  NA2        u133(.A(x10), .B(x05), .Y(men_men_n156_));
  NA2        u134(.A(x09), .B(x06), .Y(men_men_n157_));
  NO2        u135(.A(x09), .B(x01), .Y(men_men_n158_));
  NO3        u136(.A(men_men_n158_), .B(men_men_n106_), .C(men_men_n31_), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n159_), .B(x00), .Y(men_men_n160_));
  NO2        u138(.A(men_men_n112_), .B(x08), .Y(men_men_n161_));
  NA3        u139(.A(men_men_n144_), .B(men_men_n143_), .C(men_men_n50_), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n92_), .B(x05), .Y(men_men_n163_));
  OAI210     u141(.A0(men_men_n163_), .A1(men_men_n114_), .B0(men_men_n162_), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n161_), .A1(x06), .B0(men_men_n164_), .Y(men_men_n165_));
  OAI210     u143(.A0(men_men_n165_), .A1(x11), .B0(men_men_n160_), .Y(men_men_n166_));
  NAi21      u144(.An(men_men_n155_), .B(men_men_n166_), .Y(men_men_n167_));
  INV        u145(.A(men_men_n25_), .Y(men_men_n168_));
  NAi21      u146(.An(x13), .B(x00), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n169_), .Y(men_men_n170_));
  AOI220     u148(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n156_), .A1(men_men_n35_), .B0(men_men_n171_), .Y(men_men_n172_));
  AN2        u150(.A(men_men_n172_), .B(men_men_n170_), .Y(men_men_n173_));
  BUFFER     u151(.A(men_men_n71_), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n93_), .B(x06), .Y(men_men_n175_));
  NO2        u153(.A(men_men_n169_), .B(men_men_n36_), .Y(men_men_n176_));
  INV        u154(.A(men_men_n176_), .Y(men_men_n177_));
  OAI220     u155(.A0(men_men_n177_), .A1(men_men_n157_), .B0(men_men_n175_), .B1(men_men_n174_), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n178_), .A1(men_men_n173_), .B0(men_men_n168_), .Y(men_men_n179_));
  NOi21      u157(.An(x09), .B(x00), .Y(men_men_n180_));
  NO3        u158(.A(men_men_n80_), .B(men_men_n180_), .C(men_men_n47_), .Y(men_men_n181_));
  NA2        u159(.A(men_men_n181_), .B(men_men_n120_), .Y(men_men_n182_));
  NA2        u160(.A(x10), .B(x08), .Y(men_men_n183_));
  INV        u161(.A(men_men_n183_), .Y(men_men_n184_));
  NA2        u162(.A(x06), .B(x05), .Y(men_men_n185_));
  OAI210     u163(.A0(men_men_n185_), .A1(men_men_n35_), .B0(men_men_n98_), .Y(men_men_n186_));
  AOI210     u164(.A0(men_men_n184_), .A1(men_men_n57_), .B0(men_men_n186_), .Y(men_men_n187_));
  NA2        u165(.A(men_men_n187_), .B(men_men_n182_), .Y(men_men_n188_));
  NO2        u166(.A(men_men_n99_), .B(x12), .Y(men_men_n189_));
  AOI210     u167(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n189_), .Y(men_men_n190_));
  NA2        u168(.A(men_men_n92_), .B(men_men_n50_), .Y(men_men_n191_));
  NO2        u169(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n192_));
  NA2        u170(.A(men_men_n192_), .B(x02), .Y(men_men_n193_));
  NO2        u171(.A(men_men_n193_), .B(men_men_n191_), .Y(men_men_n194_));
  AOI210     u172(.A0(men_men_n190_), .A1(men_men_n188_), .B0(men_men_n194_), .Y(men_men_n195_));
  NA4        u173(.A(men_men_n195_), .B(men_men_n179_), .C(men_men_n167_), .D(men_men_n154_), .Y(men_men_n196_));
  AOI210     u174(.A0(men_men_n142_), .A1(men_men_n98_), .B0(men_men_n196_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n119_), .B(x06), .Y(men_men_n198_));
  AOI210     u176(.A0(x06), .A1(men_men_n73_), .B0(x12), .Y(men_men_n199_));
  INV        u177(.A(men_men_n76_), .Y(men_men_n200_));
  NA2        u178(.A(men_men_n145_), .B(men_men_n56_), .Y(men_men_n201_));
  NA2        u179(.A(men_men_n201_), .B(men_men_n200_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n92_), .B(x06), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n36_), .A1(x04), .B0(men_men_n50_), .Y(men_men_n204_));
  NO3        u182(.A(men_men_n204_), .B(men_men_n203_), .C(men_men_n41_), .Y(men_men_n205_));
  NA4        u183(.A(men_men_n143_), .B(men_men_n55_), .C(men_men_n36_), .D(x04), .Y(men_men_n206_));
  NA2        u184(.A(men_men_n206_), .B(men_men_n133_), .Y(men_men_n207_));
  OAI210     u185(.A0(men_men_n207_), .A1(men_men_n205_), .B0(x02), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n208_), .A1(men_men_n202_), .B0(men_men_n23_), .Y(men_men_n209_));
  OAI210     u187(.A0(men_men_n199_), .A1(men_men_n56_), .B0(men_men_n209_), .Y(men_men_n210_));
  INV        u188(.A(men_men_n133_), .Y(men_men_n211_));
  NO2        u189(.A(men_men_n50_), .B(x03), .Y(men_men_n212_));
  INV        u190(.A(men_men_n143_), .Y(men_men_n213_));
  INV        u191(.A(men_men_n89_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n214_), .B(x12), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n217_));
  OAI210     u195(.A0(men_men_n217_), .A1(men_men_n172_), .B0(men_men_n170_), .Y(men_men_n218_));
  OAI210     u196(.A0(men_men_n101_), .A1(men_men_n137_), .B0(men_men_n72_), .Y(men_men_n219_));
  INV        u197(.A(men_men_n219_), .Y(men_men_n220_));
  INV        u198(.A(x03), .Y(men_men_n221_));
  OA210      u199(.A0(men_men_n221_), .A1(men_men_n220_), .B0(men_men_n218_), .Y(men_men_n222_));
  NA2        u200(.A(x13), .B(men_men_n98_), .Y(men_men_n223_));
  NA3        u201(.A(men_men_n223_), .B(men_men_n186_), .C(men_men_n90_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n222_), .A1(men_men_n216_), .B0(men_men_n224_), .Y(men_men_n225_));
  NO2        u203(.A(men_men_n215_), .B(men_men_n225_), .Y(men_men_n226_));
  AOI210     u204(.A0(men_men_n226_), .A1(men_men_n210_), .B0(x07), .Y(men_men_n227_));
  NA2        u205(.A(men_men_n71_), .B(men_men_n29_), .Y(men_men_n228_));
  NO2        u206(.A(x12), .B(x02), .Y(men_men_n229_));
  INV        u207(.A(men_men_n229_), .Y(men_men_n230_));
  NA2        u208(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n231_), .B(x01), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n99_), .B(x04), .Y(men_men_n233_));
  NA2        u211(.A(x02), .B(x06), .Y(men_men_n234_));
  NO3        u212(.A(men_men_n88_), .B(x12), .C(x03), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n234_), .A1(x10), .B0(men_men_n235_), .Y(men_men_n236_));
  AOI210     u214(.A0(men_men_n191_), .A1(men_men_n185_), .B0(men_men_n101_), .Y(men_men_n237_));
  NOi21      u215(.An(men_men_n228_), .B(men_men_n203_), .Y(men_men_n238_));
  NO2        u216(.A(men_men_n25_), .B(x00), .Y(men_men_n239_));
  OAI210     u217(.A0(men_men_n238_), .A1(men_men_n237_), .B0(men_men_n239_), .Y(men_men_n240_));
  NO2        u218(.A(men_men_n57_), .B(x05), .Y(men_men_n241_));
  NO3        u219(.A(men_men_n241_), .B(men_men_n204_), .C(men_men_n175_), .Y(men_men_n242_));
  NO2        u220(.A(men_men_n216_), .B(men_men_n28_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n242_), .A1(men_men_n211_), .B0(men_men_n243_), .Y(men_men_n244_));
  NA3        u222(.A(men_men_n244_), .B(men_men_n240_), .C(men_men_n236_), .Y(men_men_n245_));
  NO2        u223(.A(men_men_n245_), .B(men_men_n227_), .Y(men_men_n246_));
  OAI210     u224(.A0(men_men_n197_), .A1(men_men_n60_), .B0(men_men_n246_), .Y(men02));
  NA2        u225(.A(men_men_n184_), .B(men_men_n55_), .Y(men_men_n248_));
  OAI210     u226(.A0(x01), .A1(men_men_n32_), .B0(men_men_n248_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n249_), .B(men_men_n156_), .Y(men_men_n250_));
  INV        u228(.A(men_men_n156_), .Y(men_men_n251_));
  AOI210     u229(.A0(men_men_n113_), .A1(men_men_n83_), .B0(men_men_n204_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(men_men_n99_), .Y(men_men_n253_));
  AOI210     u231(.A0(men_men_n253_), .A1(men_men_n251_), .B0(men_men_n140_), .Y(men_men_n254_));
  AOI210     u232(.A0(men_men_n254_), .A1(men_men_n250_), .B0(men_men_n48_), .Y(men_men_n255_));
  AOI210     u233(.A0(men_men_n55_), .A1(men_men_n36_), .B0(men_men_n57_), .Y(men_men_n256_));
  NO2        u234(.A(x02), .B(men_men_n133_), .Y(men_men_n257_));
  NO2        u235(.A(x10), .B(men_men_n47_), .Y(men_men_n258_));
  INV        u236(.A(men_men_n258_), .Y(men_men_n259_));
  AN2        u237(.A(men_men_n387_), .B(x08), .Y(men_men_n260_));
  OAI210     u238(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n261_));
  BUFFER     u239(.A(men_men_n136_), .Y(men_men_n262_));
  AOI210     u240(.A0(men_men_n262_), .A1(x04), .B0(men_men_n261_), .Y(men_men_n263_));
  OAI210     u241(.A0(men_men_n263_), .A1(men_men_n260_), .B0(men_men_n93_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n93_), .B(men_men_n212_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n265_), .B(x04), .Y(men_men_n266_));
  INV        u244(.A(men_men_n140_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n267_), .B(men_men_n121_), .Y(men_men_n268_));
  AOI210     u246(.A0(men_men_n268_), .A1(x13), .B0(men_men_n266_), .Y(men_men_n269_));
  NA3        u247(.A(men_men_n269_), .B(men_men_n264_), .C(men_men_n259_), .Y(men_men_n270_));
  NO3        u248(.A(men_men_n270_), .B(men_men_n257_), .C(men_men_n255_), .Y(men_men_n271_));
  NA2        u249(.A(men_men_n132_), .B(x03), .Y(men_men_n272_));
  OAI210     u250(.A0(men_men_n169_), .A1(men_men_n241_), .B0(men_men_n272_), .Y(men_men_n273_));
  NA2        u251(.A(men_men_n273_), .B(men_men_n106_), .Y(men_men_n274_));
  NA2        u252(.A(men_men_n155_), .B(men_men_n149_), .Y(men_men_n275_));
  BUFFER     u253(.A(men_men_n275_), .Y(men_men_n276_));
  OAI220     u254(.A0(men_men_n233_), .A1(x09), .B0(men_men_n122_), .B1(men_men_n28_), .Y(men_men_n277_));
  OAI210     u255(.A0(men_men_n277_), .A1(men_men_n276_), .B0(men_men_n107_), .Y(men_men_n278_));
  NA2        u256(.A(men_men_n233_), .B(men_men_n98_), .Y(men_men_n279_));
  NA2        u257(.A(men_men_n98_), .B(men_men_n41_), .Y(men_men_n280_));
  NA3        u258(.A(men_men_n280_), .B(men_men_n279_), .C(men_men_n121_), .Y(men_men_n281_));
  NA4        u259(.A(men_men_n281_), .B(men_men_n278_), .C(men_men_n274_), .D(men_men_n48_), .Y(men_men_n282_));
  INV        u260(.A(men_men_n192_), .Y(men_men_n283_));
  NA2        u261(.A(men_men_n189_), .B(x04), .Y(men_men_n284_));
  NO2        u262(.A(men_men_n284_), .B(men_men_n36_), .Y(men_men_n285_));
  NO3        u263(.A(men_men_n171_), .B(x13), .C(men_men_n31_), .Y(men_men_n286_));
  OAI210     u264(.A0(men_men_n286_), .A1(men_men_n285_), .B0(men_men_n93_), .Y(men_men_n287_));
  NO3        u265(.A(men_men_n189_), .B(men_men_n148_), .C(men_men_n51_), .Y(men_men_n288_));
  OAI210     u266(.A0(x12), .A1(men_men_n181_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA3        u267(.A(men_men_n289_), .B(men_men_n287_), .C(x06), .Y(men_men_n290_));
  NA2        u268(.A(x09), .B(x03), .Y(men_men_n291_));
  OAI220     u269(.A0(men_men_n291_), .A1(men_men_n120_), .B0(x01), .B1(men_men_n63_), .Y(men_men_n292_));
  NO2        u270(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n288_), .B(men_men_n293_), .Y(men_men_n294_));
  INV        u272(.A(men_men_n294_), .Y(men_men_n295_));
  AO220      u273(.A0(men_men_n295_), .A1(x04), .B0(men_men_n292_), .B1(x05), .Y(men_men_n296_));
  AOI210     u274(.A0(men_men_n290_), .A1(men_men_n282_), .B0(men_men_n296_), .Y(men_men_n297_));
  OAI210     u275(.A0(men_men_n271_), .A1(x12), .B0(men_men_n297_), .Y(men03));
  OR2        u276(.A(men_men_n42_), .B(men_men_n212_), .Y(men_men_n299_));
  AOI210     u277(.A0(men_men_n35_), .A1(men_men_n98_), .B0(men_men_n299_), .Y(men_men_n300_));
  OAI210     u278(.A0(men_men_n385_), .A1(men_men_n300_), .B0(x05), .Y(men_men_n301_));
  NA2        u279(.A(men_men_n299_), .B(x05), .Y(men_men_n302_));
  NO2        u280(.A(x04), .B(men_men_n302_), .Y(men_men_n303_));
  NO2        u281(.A(x02), .B(men_men_n256_), .Y(men_men_n304_));
  OAI210     u282(.A0(men_men_n304_), .A1(men_men_n303_), .B0(men_men_n98_), .Y(men_men_n305_));
  AOI210     u283(.A0(men_men_n136_), .A1(men_men_n59_), .B0(men_men_n38_), .Y(men_men_n306_));
  NO2        u284(.A(men_men_n158_), .B(men_men_n126_), .Y(men_men_n307_));
  OAI220     u285(.A0(men_men_n307_), .A1(men_men_n37_), .B0(men_men_n138_), .B1(x13), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n308_), .A1(men_men_n306_), .B0(x04), .Y(men_men_n309_));
  NO3        u287(.A(men_men_n280_), .B(men_men_n82_), .C(men_men_n58_), .Y(men_men_n310_));
  AOI210     u288(.A0(men_men_n177_), .A1(men_men_n98_), .B0(men_men_n136_), .Y(men_men_n311_));
  OA210      u289(.A0(men_men_n150_), .A1(x12), .B0(men_men_n126_), .Y(men_men_n312_));
  NO3        u290(.A(men_men_n312_), .B(men_men_n311_), .C(men_men_n310_), .Y(men_men_n313_));
  NA4        u291(.A(men_men_n313_), .B(men_men_n309_), .C(men_men_n305_), .D(men_men_n301_), .Y(men04));
  NO2        u292(.A(men_men_n86_), .B(men_men_n39_), .Y(men_men_n315_));
  XO2        u293(.A(men_men_n315_), .B(men_men_n223_), .Y(men05));
  AOI210     u294(.A0(men_men_n71_), .A1(men_men_n51_), .B0(men_men_n198_), .Y(men_men_n317_));
  AOI210     u295(.A0(men_men_n317_), .A1(men_men_n261_), .B0(men_men_n25_), .Y(men_men_n318_));
  AOI210     u296(.A0(men_men_n213_), .A1(men_men_n56_), .B0(men_men_n87_), .Y(men_men_n319_));
  NO2        u297(.A(men_men_n319_), .B(men_men_n24_), .Y(men_men_n320_));
  OAI210     u298(.A0(men_men_n320_), .A1(men_men_n318_), .B0(men_men_n98_), .Y(men_men_n321_));
  NA2        u299(.A(x11), .B(men_men_n31_), .Y(men_men_n322_));
  NA2        u300(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n228_), .B(x03), .Y(men_men_n324_));
  OAI220     u302(.A0(men_men_n324_), .A1(men_men_n323_), .B0(men_men_n322_), .B1(men_men_n79_), .Y(men_men_n325_));
  OAI210     u303(.A0(men_men_n26_), .A1(men_men_n98_), .B0(x07), .Y(men_men_n326_));
  AOI210     u304(.A0(men_men_n325_), .A1(x06), .B0(men_men_n326_), .Y(men_men_n327_));
  AOI220     u305(.A0(men_men_n79_), .A1(men_men_n31_), .B0(men_men_n51_), .B1(men_men_n50_), .Y(men_men_n328_));
  NO3        u306(.A(men_men_n328_), .B(men_men_n23_), .C(x00), .Y(men_men_n329_));
  NA2        u307(.A(men_men_n70_), .B(x02), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(men_men_n324_), .Y(men_men_n331_));
  OR2        u309(.A(men_men_n331_), .B(men_men_n216_), .Y(men_men_n332_));
  NO2        u310(.A(men_men_n23_), .B(x10), .Y(men_men_n333_));
  OAI210     u311(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n334_));
  OR3        u312(.A(men_men_n334_), .B(men_men_n333_), .C(men_men_n44_), .Y(men_men_n335_));
  NA2        u313(.A(men_men_n335_), .B(men_men_n332_), .Y(men_men_n336_));
  OAI210     u314(.A0(men_men_n336_), .A1(men_men_n329_), .B0(men_men_n98_), .Y(men_men_n337_));
  AOI220     u315(.A0(men_men_n388_), .A1(men_men_n337_), .B0(men_men_n327_), .B1(men_men_n321_), .Y(men_men_n338_));
  NA3        u316(.A(men_men_n23_), .B(men_men_n60_), .C(men_men_n48_), .Y(men_men_n339_));
  AO210      u317(.A0(men_men_n339_), .A1(men_men_n231_), .B0(men_men_n230_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n333_), .A1(men_men_n74_), .B0(men_men_n132_), .Y(men_men_n341_));
  OR2        u319(.A(men_men_n341_), .B(x03), .Y(men_men_n342_));
  NA2        u320(.A(men_men_n293_), .B(men_men_n60_), .Y(men_men_n343_));
  NO2        u321(.A(men_men_n343_), .B(x11), .Y(men_men_n344_));
  NO3        u322(.A(men_men_n344_), .B(men_men_n135_), .C(men_men_n28_), .Y(men_men_n345_));
  AOI220     u323(.A0(men_men_n345_), .A1(men_men_n342_), .B0(men_men_n340_), .B1(men_men_n47_), .Y(men_men_n346_));
  NO4        u324(.A(men_men_n280_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n347_));
  OAI210     u325(.A0(men_men_n347_), .A1(men_men_n346_), .B0(men_men_n99_), .Y(men_men_n348_));
  AOI210     u326(.A0(men_men_n284_), .A1(men_men_n108_), .B0(men_men_n229_), .Y(men_men_n349_));
  NOi21      u327(.An(men_men_n272_), .B(men_men_n126_), .Y(men_men_n350_));
  NO2        u328(.A(men_men_n349_), .B(x08), .Y(men_men_n351_));
  AOI210     u329(.A0(men_men_n333_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n352_));
  NA2        u330(.A(x09), .B(men_men_n41_), .Y(men_men_n353_));
  OAI220     u331(.A0(men_men_n353_), .A1(men_men_n352_), .B0(men_men_n322_), .B1(men_men_n66_), .Y(men_men_n354_));
  NO2        u332(.A(x13), .B(x12), .Y(men_men_n355_));
  NO2        u333(.A(men_men_n122_), .B(men_men_n28_), .Y(men_men_n356_));
  NO2        u334(.A(men_men_n356_), .B(men_men_n232_), .Y(men_men_n357_));
  NA3        u335(.A(men_men_n283_), .B(men_men_n117_), .C(x12), .Y(men_men_n358_));
  AO210      u336(.A0(men_men_n283_), .A1(men_men_n117_), .B0(men_men_n223_), .Y(men_men_n359_));
  NA3        u337(.A(men_men_n359_), .B(men_men_n358_), .C(x08), .Y(men_men_n360_));
  AOI210     u338(.A0(men_men_n355_), .A1(men_men_n354_), .B0(men_men_n360_), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n351_), .A1(men_men_n348_), .B0(men_men_n361_), .Y(men_men_n362_));
  OAI210     u340(.A0(men_men_n343_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n363_));
  NA2        u341(.A(men_men_n251_), .B(x07), .Y(men_men_n364_));
  NO2        u342(.A(men_men_n364_), .B(men_men_n323_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n363_), .B0(men_men_n176_), .Y(men_men_n366_));
  NA3        u344(.A(men_men_n357_), .B(men_men_n350_), .C(men_men_n279_), .Y(men_men_n367_));
  INV        u345(.A(x14), .Y(men_men_n368_));
  NO3        u346(.A(men_men_n272_), .B(men_men_n104_), .C(x11), .Y(men_men_n369_));
  NO3        u347(.A(men_men_n149_), .B(men_men_n74_), .C(men_men_n56_), .Y(men_men_n370_));
  NO3        u348(.A(men_men_n339_), .B(men_men_n280_), .C(men_men_n169_), .Y(men_men_n371_));
  NO4        u349(.A(men_men_n371_), .B(men_men_n370_), .C(men_men_n369_), .D(men_men_n368_), .Y(men_men_n372_));
  NA3        u350(.A(men_men_n372_), .B(men_men_n367_), .C(men_men_n366_), .Y(men_men_n373_));
  AOI220     u351(.A0(x12), .A1(men_men_n60_), .B0(men_men_n356_), .B1(men_men_n148_), .Y(men_men_n374_));
  NOi21      u352(.An(men_men_n233_), .B(men_men_n138_), .Y(men_men_n375_));
  NO3        u353(.A(men_men_n119_), .B(men_men_n24_), .C(x06), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n239_), .A1(men_men_n213_), .B0(men_men_n376_), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n44_), .A1(x04), .B0(men_men_n377_), .Y(men_men_n378_));
  OAI210     u356(.A0(men_men_n378_), .A1(men_men_n375_), .B0(men_men_n98_), .Y(men_men_n379_));
  OAI210     u357(.A0(men_men_n374_), .A1(men_men_n88_), .B0(men_men_n379_), .Y(men_men_n380_));
  NO4        u358(.A(men_men_n380_), .B(men_men_n373_), .C(men_men_n362_), .D(men_men_n338_), .Y(men06));
  INV        u359(.A(x01), .Y(men_men_n384_));
  INV        u360(.A(men_men_n284_), .Y(men_men_n385_));
  INV        u361(.A(x08), .Y(men_men_n386_));
  INV        u362(.A(x03), .Y(men_men_n387_));
  INV        u363(.A(x07), .Y(men_men_n388_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule