// Benchmark "top" written by ABC on Thu Jun 20 14:59:11 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n42_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n776_, new_new_n777_,
    new_new_n778_, new_new_n779_, new_new_n780_, new_new_n781_,
    new_new_n782_, new_new_n783_, new_new_n784_, new_new_n785_,
    new_new_n786_, new_new_n787_, new_new_n788_, new_new_n789_,
    new_new_n790_, new_new_n791_, new_new_n792_, new_new_n793_,
    new_new_n794_, new_new_n795_, new_new_n796_, new_new_n797_,
    new_new_n798_, new_new_n799_, new_new_n800_, new_new_n801_,
    new_new_n802_, new_new_n803_, new_new_n804_, new_new_n805_,
    new_new_n806_, new_new_n807_, new_new_n808_, new_new_n809_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n825_, new_new_n826_,
    new_new_n827_, new_new_n828_, new_new_n829_, new_new_n830_,
    new_new_n831_, new_new_n832_, new_new_n833_, new_new_n834_,
    new_new_n835_, new_new_n836_, new_new_n837_, new_new_n838_,
    new_new_n839_, new_new_n840_, new_new_n841_, new_new_n842_,
    new_new_n843_, new_new_n844_, new_new_n845_, new_new_n846_,
    new_new_n847_, new_new_n848_, new_new_n849_, new_new_n850_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n875_,
    new_new_n876_, new_new_n877_, new_new_n878_, new_new_n879_,
    new_new_n880_, new_new_n881_, new_new_n882_, new_new_n883_,
    new_new_n884_, new_new_n885_, new_new_n886_, new_new_n887_,
    new_new_n888_, new_new_n889_, new_new_n890_, new_new_n891_,
    new_new_n892_, new_new_n893_, new_new_n894_, new_new_n895_,
    new_new_n896_, new_new_n897_, new_new_n898_, new_new_n899_,
    new_new_n900_, new_new_n901_, new_new_n902_, new_new_n903_,
    new_new_n904_, new_new_n905_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1100_,
    new_new_n1101_, new_new_n1102_, new_new_n1103_, new_new_n1104_,
    new_new_n1105_, new_new_n1106_, new_new_n1107_, new_new_n1108_,
    new_new_n1109_, new_new_n1110_, new_new_n1111_, new_new_n1112_,
    new_new_n1113_, new_new_n1114_, new_new_n1115_, new_new_n1116_,
    new_new_n1117_, new_new_n1118_, new_new_n1119_, new_new_n1120_,
    new_new_n1121_, new_new_n1122_, new_new_n1123_, new_new_n1124_,
    new_new_n1125_, new_new_n1126_, new_new_n1127_, new_new_n1128_,
    new_new_n1129_, new_new_n1130_, new_new_n1131_, new_new_n1132_,
    new_new_n1133_, new_new_n1134_, new_new_n1135_, new_new_n1136_,
    new_new_n1137_, new_new_n1138_, new_new_n1139_, new_new_n1140_,
    new_new_n1141_, new_new_n1142_, new_new_n1146_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  NOi21      g0006(.An(i_11_), .B(i_8_), .Y(new_new_n29_));
  AO210      g0007(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n30_));
  OR2        g0008(.A(new_new_n30_), .B(new_new_n29_), .Y(new_new_n31_));
  NA2        g0009(.A(new_new_n31_), .B(new_new_n26_), .Y(new_new_n32_));
  XO2        g0010(.A(new_new_n32_), .B(new_new_n23_), .Y(new_new_n33_));
  INV        g0011(.A(i_4_), .Y(new_new_n34_));
  INV        g0012(.A(i_10_), .Y(new_new_n35_));
  NAi21      g0013(.An(i_11_), .B(i_9_), .Y(new_new_n36_));
  NOi21      g0014(.An(i_12_), .B(i_13_), .Y(new_new_n37_));
  INV        g0015(.A(new_new_n37_), .Y(new_new_n38_));
  NO2        g0016(.A(new_new_n34_), .B(i_3_), .Y(new_new_n39_));
  NAi31      g0017(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n33_), .Y(men1));
  INV        g0019(.A(i_11_), .Y(new_new_n42_));
  NO2        g0020(.A(new_new_n42_), .B(i_6_), .Y(new_new_n43_));
  INV        g0021(.A(i_2_), .Y(new_new_n44_));
  NA2        g0022(.A(i_0_), .B(i_3_), .Y(new_new_n45_));
  INV        g0023(.A(i_5_), .Y(new_new_n46_));
  NO2        g0024(.A(i_7_), .B(i_10_), .Y(new_new_n47_));
  AOI210     g0025(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n47_), .Y(new_new_n48_));
  OAI210     g0026(.A0(new_new_n48_), .A1(i_3_), .B0(new_new_n46_), .Y(new_new_n49_));
  AOI210     g0027(.A0(new_new_n49_), .A1(new_new_n45_), .B0(new_new_n44_), .Y(new_new_n50_));
  NA2        g0028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g0029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g0030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  OAI210     g0031(.A0(new_new_n53_), .A1(new_new_n50_), .B0(new_new_n43_), .Y(new_new_n54_));
  NA3        g0032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g0033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g0034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  OAI210     g0035(.A0(new_new_n57_), .A1(new_new_n56_), .B0(new_new_n55_), .Y(new_new_n58_));
  NA2        g0036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g0037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g0038(.A(i_1_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g0040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n29_), .Y(new_new_n63_));
  NA2        g0041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi31      g0043(.An(new_new_n65_), .B(new_new_n63_), .C(new_new_n59_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n48_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g0053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(new_new_n79_), .B(new_new_n56_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  NO3        g0060(.A(new_new_n82_), .B(new_new_n81_), .C(new_new_n61_), .Y(new_new_n83_));
  INV        g0061(.A(i_6_), .Y(new_new_n84_));
  OR4        g0062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n85_));
  INV        g0063(.A(new_new_n85_), .Y(new_new_n86_));
  NO2        g0064(.A(i_2_), .B(i_7_), .Y(new_new_n87_));
  AOI210     g0065(.A0(new_new_n86_), .A1(new_new_n84_), .B0(new_new_n87_), .Y(new_new_n88_));
  OAI210     g0066(.A0(new_new_n83_), .A1(new_new_n80_), .B0(new_new_n88_), .Y(new_new_n89_));
  NAi21      g0067(.An(i_6_), .B(i_10_), .Y(new_new_n90_));
  NA2        g0068(.A(i_6_), .B(i_9_), .Y(new_new_n91_));
  AOI210     g0069(.A0(new_new_n91_), .A1(new_new_n90_), .B0(new_new_n61_), .Y(new_new_n92_));
  NA2        g0070(.A(i_2_), .B(i_6_), .Y(new_new_n93_));
  NO3        g0071(.A(new_new_n93_), .B(new_new_n47_), .C(new_new_n25_), .Y(new_new_n94_));
  NO2        g0072(.A(new_new_n94_), .B(new_new_n92_), .Y(new_new_n95_));
  AOI210     g0073(.A0(new_new_n95_), .A1(new_new_n89_), .B0(new_new_n78_), .Y(new_new_n96_));
  AN3        g0074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n97_));
  NAi21      g0075(.An(i_6_), .B(i_11_), .Y(new_new_n98_));
  NO2        g0076(.A(i_5_), .B(i_8_), .Y(new_new_n99_));
  NOi21      g0077(.An(new_new_n99_), .B(new_new_n98_), .Y(new_new_n100_));
  AOI220     g0078(.A0(new_new_n100_), .A1(new_new_n60_), .B0(new_new_n97_), .B1(new_new_n30_), .Y(new_new_n101_));
  INV        g0079(.A(i_7_), .Y(new_new_n102_));
  NA2        g0080(.A(new_new_n44_), .B(new_new_n102_), .Y(new_new_n103_));
  NO2        g0081(.A(i_0_), .B(i_5_), .Y(new_new_n104_));
  NO2        g0082(.A(new_new_n104_), .B(new_new_n84_), .Y(new_new_n105_));
  NA2        g0083(.A(i_12_), .B(i_3_), .Y(new_new_n106_));
  INV        g0084(.A(new_new_n106_), .Y(new_new_n107_));
  NA3        g0085(.A(new_new_n107_), .B(new_new_n105_), .C(new_new_n103_), .Y(new_new_n108_));
  NAi21      g0086(.An(i_7_), .B(i_11_), .Y(new_new_n109_));
  NO3        g0087(.A(new_new_n109_), .B(new_new_n90_), .C(new_new_n51_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g0089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g0090(.A(new_new_n78_), .B(new_new_n56_), .Y(new_new_n113_));
  NO2        g0091(.A(i_8_), .B(new_new_n102_), .Y(new_new_n114_));
  NO3        g0092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g0093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g0094(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g0096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g0097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g0098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NAi41      g0099(.An(new_new_n110_), .B(new_new_n121_), .C(new_new_n108_), .D(new_new_n101_), .Y(new_new_n122_));
  NOi21      g0100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n102_), .B(new_new_n35_), .Y(new_new_n125_));
  NA2        g0103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g0105(.A(new_new_n127_), .B(new_new_n44_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n91_), .B(new_new_n90_), .Y(new_new_n129_));
  NAi21      g0107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n130_), .B(new_new_n60_), .Y(new_new_n131_));
  NOi31      g0109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g0110(.A(i_1_), .B(new_new_n84_), .Y(new_new_n133_));
  NO2        g0111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g0113(.A0(new_new_n135_), .A1(new_new_n45_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g0114(.A0(new_new_n136_), .A1(new_new_n109_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g0115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n96_), .Y(new_new_n138_));
  NA3        g0116(.A(new_new_n138_), .B(new_new_n77_), .C(new_new_n54_), .Y(men2));
  NO2        g0117(.A(new_new_n61_), .B(new_new_n35_), .Y(new_new_n140_));
  NA2        g0118(.A(i_6_), .B(new_new_n25_), .Y(new_new_n141_));
  NA3        g0119(.A(new_new_n75_), .B(new_new_n67_), .C(new_new_n26_), .Y(men0));
  AN2        g0120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g0122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g0123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g0124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g0125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g0126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  OR2        g0129(.A(new_new_n151_), .B(new_new_n25_), .Y(new_new_n152_));
  AN2        g0130(.A(new_new_n145_), .B(new_new_n81_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(new_new_n27_), .Y(new_new_n154_));
  NA2        g0132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n71_), .B(new_new_n44_), .Y(new_new_n156_));
  NA2        g0134(.A(new_new_n156_), .B(new_new_n34_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n158_));
  OR2        g0136(.A(i_0_), .B(i_1_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n160_));
  NAi32      g0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n161_));
  NAi21      g0139(.An(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NOi21      g0140(.An(i_4_), .B(i_10_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n37_), .Y(new_new_n164_));
  NO2        g0142(.A(i_3_), .B(i_5_), .Y(new_new_n165_));
  NO3        g0143(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  OAI210     g0145(.A0(new_new_n167_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n168_));
  NO2        g0146(.A(new_new_n168_), .B(new_new_n158_), .Y(new_new_n169_));
  AOI210     g0147(.A0(new_new_n169_), .A1(new_new_n152_), .B0(new_new_n144_), .Y(new_new_n170_));
  NA3        g0148(.A(new_new_n71_), .B(new_new_n44_), .C(i_1_), .Y(new_new_n171_));
  NA2        g0149(.A(i_3_), .B(new_new_n46_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_4_), .B(i_9_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_11_), .B(i_13_), .Y(new_new_n174_));
  NA2        g0152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  OR2        g0153(.A(new_new_n175_), .B(new_new_n172_), .Y(new_new_n176_));
  NO2        g0154(.A(i_4_), .B(i_5_), .Y(new_new_n177_));
  NAi21      g0155(.An(i_12_), .B(i_11_), .Y(new_new_n178_));
  NO2        g0156(.A(new_new_n178_), .B(i_13_), .Y(new_new_n179_));
  NA3        g0157(.A(new_new_n179_), .B(new_new_n177_), .C(new_new_n81_), .Y(new_new_n180_));
  AOI210     g0158(.A0(new_new_n180_), .A1(new_new_n176_), .B0(new_new_n171_), .Y(new_new_n181_));
  NO2        g0159(.A(new_new_n71_), .B(new_new_n61_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n182_), .B(new_new_n44_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n34_), .B(i_5_), .Y(new_new_n184_));
  NAi31      g0162(.An(new_new_n184_), .B(new_new_n153_), .C(i_11_), .Y(new_new_n185_));
  NA2        g0163(.A(i_3_), .B(i_5_), .Y(new_new_n186_));
  OR2        g0164(.A(new_new_n186_), .B(new_new_n175_), .Y(new_new_n187_));
  AOI210     g0165(.A0(new_new_n187_), .A1(new_new_n185_), .B0(new_new_n183_), .Y(new_new_n188_));
  NO2        g0166(.A(new_new_n71_), .B(i_5_), .Y(new_new_n189_));
  NO2        g0167(.A(i_13_), .B(i_10_), .Y(new_new_n190_));
  NA3        g0168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n42_), .Y(new_new_n191_));
  NO2        g0169(.A(i_2_), .B(i_1_), .Y(new_new_n192_));
  NA2        g0170(.A(new_new_n192_), .B(i_3_), .Y(new_new_n193_));
  NAi21      g0171(.An(i_4_), .B(i_12_), .Y(new_new_n194_));
  NO4        g0172(.A(new_new_n194_), .B(new_new_n193_), .C(new_new_n191_), .D(new_new_n25_), .Y(new_new_n195_));
  NO3        g0173(.A(new_new_n195_), .B(new_new_n188_), .C(new_new_n181_), .Y(new_new_n196_));
  INV        g0174(.A(i_8_), .Y(new_new_n197_));
  NO2        g0175(.A(new_new_n197_), .B(i_7_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(i_6_), .Y(new_new_n199_));
  NO3        g0177(.A(i_3_), .B(new_new_n84_), .C(new_new_n46_), .Y(new_new_n200_));
  NA2        g0178(.A(new_new_n200_), .B(new_new_n114_), .Y(new_new_n201_));
  NO3        g0179(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n202_));
  NA3        g0180(.A(new_new_n202_), .B(new_new_n37_), .C(new_new_n42_), .Y(new_new_n203_));
  NO3        g0181(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n204_));
  OAI210     g0182(.A0(new_new_n97_), .A1(i_12_), .B0(new_new_n204_), .Y(new_new_n205_));
  AOI210     g0183(.A0(new_new_n205_), .A1(new_new_n203_), .B0(new_new_n201_), .Y(new_new_n206_));
  NO2        g0184(.A(i_3_), .B(i_8_), .Y(new_new_n207_));
  NO3        g0185(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(new_new_n207_), .C(new_new_n37_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n104_), .B(new_new_n56_), .Y(new_new_n210_));
  NA2        g0188(.A(new_new_n210_), .B(new_new_n159_), .Y(new_new_n211_));
  NO2        g0189(.A(i_13_), .B(i_9_), .Y(new_new_n212_));
  NA3        g0190(.A(new_new_n212_), .B(i_6_), .C(new_new_n197_), .Y(new_new_n213_));
  NAi21      g0191(.An(i_12_), .B(i_3_), .Y(new_new_n214_));
  OR2        g0192(.A(new_new_n214_), .B(new_new_n213_), .Y(new_new_n215_));
  NO2        g0193(.A(new_new_n42_), .B(i_5_), .Y(new_new_n216_));
  NO3        g0194(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n217_));
  NA3        g0195(.A(new_new_n217_), .B(new_new_n216_), .C(i_10_), .Y(new_new_n218_));
  OAI220     g0196(.A0(new_new_n218_), .A1(new_new_n215_), .B0(new_new_n211_), .B1(new_new_n209_), .Y(new_new_n219_));
  AOI210     g0197(.A0(new_new_n219_), .A1(i_7_), .B0(new_new_n206_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n220_), .A1(i_4_), .B0(new_new_n199_), .B1(new_new_n196_), .Y(new_new_n221_));
  NAi21      g0199(.An(i_12_), .B(i_7_), .Y(new_new_n222_));
  NA3        g0200(.A(i_13_), .B(new_new_n197_), .C(i_10_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  NA2        g0202(.A(i_0_), .B(i_5_), .Y(new_new_n225_));
  NA2        g0203(.A(new_new_n225_), .B(new_new_n105_), .Y(new_new_n226_));
  OAI220     g0204(.A0(new_new_n226_), .A1(new_new_n193_), .B0(new_new_n183_), .B1(new_new_n135_), .Y(new_new_n227_));
  NAi31      g0205(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n34_), .B(i_13_), .Y(new_new_n229_));
  NO2        g0207(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n44_), .B(new_new_n61_), .Y(new_new_n231_));
  NA3        g0209(.A(new_new_n231_), .B(new_new_n230_), .C(new_new_n229_), .Y(new_new_n232_));
  INV        g0210(.A(i_13_), .Y(new_new_n233_));
  NO2        g0211(.A(i_12_), .B(new_new_n233_), .Y(new_new_n234_));
  NA3        g0212(.A(new_new_n234_), .B(new_new_n202_), .C(new_new_n200_), .Y(new_new_n235_));
  OAI210     g0213(.A0(new_new_n232_), .A1(new_new_n228_), .B0(new_new_n235_), .Y(new_new_n236_));
  AOI220     g0214(.A0(new_new_n236_), .A1(new_new_n143_), .B0(new_new_n227_), .B1(new_new_n224_), .Y(new_new_n237_));
  NO2        g0215(.A(i_12_), .B(new_new_n35_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n186_), .B(i_4_), .Y(new_new_n239_));
  NA2        g0217(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n240_));
  OR2        g0218(.A(i_8_), .B(i_7_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n241_), .B(new_new_n84_), .Y(new_new_n242_));
  NO2        g0220(.A(new_new_n51_), .B(i_1_), .Y(new_new_n243_));
  NA2        g0221(.A(new_new_n243_), .B(new_new_n242_), .Y(new_new_n244_));
  INV        g0222(.A(i_12_), .Y(new_new_n245_));
  NO2        g0223(.A(new_new_n42_), .B(new_new_n245_), .Y(new_new_n246_));
  NO3        g0224(.A(new_new_n34_), .B(i_8_), .C(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(i_2_), .B(i_1_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n244_), .B(new_new_n240_), .Y(new_new_n249_));
  NO3        g0227(.A(i_11_), .B(i_7_), .C(new_new_n35_), .Y(new_new_n250_));
  NAi21      g0228(.An(i_4_), .B(i_3_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n251_), .B(new_new_n73_), .Y(new_new_n252_));
  NO2        g0230(.A(i_0_), .B(i_6_), .Y(new_new_n253_));
  NOi41      g0231(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n254_));
  NA2        g0232(.A(new_new_n254_), .B(new_new_n253_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n248_), .B(new_new_n186_), .Y(new_new_n256_));
  NAi21      g0234(.An(new_new_n255_), .B(new_new_n256_), .Y(new_new_n257_));
  INV        g0235(.A(new_new_n257_), .Y(new_new_n258_));
  AOI220     g0236(.A0(new_new_n258_), .A1(new_new_n37_), .B0(new_new_n249_), .B1(new_new_n212_), .Y(new_new_n259_));
  NO2        g0237(.A(i_11_), .B(new_new_n233_), .Y(new_new_n260_));
  NOi21      g0238(.An(i_1_), .B(i_6_), .Y(new_new_n261_));
  NAi21      g0239(.An(i_3_), .B(i_7_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n245_), .B(i_9_), .Y(new_new_n263_));
  OR4        g0241(.A(new_new_n263_), .B(new_new_n262_), .C(new_new_n261_), .D(new_new_n189_), .Y(new_new_n264_));
  NO2        g0242(.A(new_new_n46_), .B(new_new_n25_), .Y(new_new_n265_));
  NO2        g0243(.A(i_12_), .B(i_3_), .Y(new_new_n266_));
  NA2        g0244(.A(new_new_n71_), .B(i_5_), .Y(new_new_n267_));
  NA2        g0245(.A(i_3_), .B(i_9_), .Y(new_new_n268_));
  NAi21      g0246(.An(i_7_), .B(i_10_), .Y(new_new_n269_));
  NO2        g0247(.A(new_new_n269_), .B(new_new_n268_), .Y(new_new_n270_));
  NA3        g0248(.A(new_new_n270_), .B(new_new_n267_), .C(new_new_n62_), .Y(new_new_n271_));
  NA2        g0249(.A(new_new_n271_), .B(new_new_n264_), .Y(new_new_n272_));
  NA3        g0250(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n273_));
  INV        g0251(.A(new_new_n144_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n245_), .B(i_13_), .Y(new_new_n275_));
  NO2        g0253(.A(new_new_n275_), .B(new_new_n73_), .Y(new_new_n276_));
  AOI220     g0254(.A0(new_new_n276_), .A1(new_new_n274_), .B0(new_new_n272_), .B1(new_new_n260_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n241_), .B(new_new_n35_), .Y(new_new_n278_));
  NA2        g0256(.A(i_12_), .B(i_6_), .Y(new_new_n279_));
  OR2        g0257(.A(i_13_), .B(i_9_), .Y(new_new_n280_));
  NO3        g0258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n46_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n251_), .B(i_2_), .Y(new_new_n282_));
  NA3        g0260(.A(new_new_n282_), .B(new_new_n281_), .C(new_new_n42_), .Y(new_new_n283_));
  NA2        g0261(.A(new_new_n260_), .B(i_9_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n267_), .B(new_new_n159_), .C(new_new_n62_), .Y(new_new_n285_));
  OAI210     g0263(.A0(new_new_n285_), .A1(new_new_n284_), .B0(new_new_n283_), .Y(new_new_n286_));
  NA2        g0264(.A(new_new_n156_), .B(new_new_n61_), .Y(new_new_n287_));
  NO3        g0265(.A(i_11_), .B(new_new_n233_), .C(new_new_n25_), .Y(new_new_n288_));
  NO2        g0266(.A(new_new_n262_), .B(i_8_), .Y(new_new_n289_));
  NO2        g0267(.A(i_6_), .B(new_new_n46_), .Y(new_new_n290_));
  NA3        g0268(.A(new_new_n290_), .B(new_new_n289_), .C(new_new_n288_), .Y(new_new_n291_));
  NO3        g0269(.A(new_new_n26_), .B(new_new_n84_), .C(i_5_), .Y(new_new_n292_));
  NA3        g0270(.A(new_new_n292_), .B(new_new_n278_), .C(new_new_n234_), .Y(new_new_n293_));
  AOI210     g0271(.A0(new_new_n293_), .A1(new_new_n291_), .B0(new_new_n287_), .Y(new_new_n294_));
  AOI210     g0272(.A0(new_new_n286_), .A1(new_new_n278_), .B0(new_new_n294_), .Y(new_new_n295_));
  NA4        g0273(.A(new_new_n295_), .B(new_new_n277_), .C(new_new_n259_), .D(new_new_n237_), .Y(new_new_n296_));
  NO3        g0274(.A(i_12_), .B(new_new_n233_), .C(new_new_n35_), .Y(new_new_n297_));
  INV        g0275(.A(new_new_n297_), .Y(new_new_n298_));
  NA2        g0276(.A(i_8_), .B(new_new_n102_), .Y(new_new_n299_));
  NOi21      g0277(.An(new_new_n165_), .B(new_new_n84_), .Y(new_new_n300_));
  NO3        g0278(.A(i_0_), .B(new_new_n44_), .C(i_1_), .Y(new_new_n301_));
  AOI220     g0279(.A0(new_new_n301_), .A1(new_new_n200_), .B0(new_new_n300_), .B1(new_new_n243_), .Y(new_new_n302_));
  NO2        g0280(.A(new_new_n302_), .B(new_new_n299_), .Y(new_new_n303_));
  NO3        g0281(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n304_));
  NO2        g0282(.A(new_new_n248_), .B(i_0_), .Y(new_new_n305_));
  AOI220     g0283(.A0(new_new_n305_), .A1(new_new_n198_), .B0(new_new_n304_), .B1(new_new_n143_), .Y(new_new_n306_));
  NA2        g0284(.A(new_new_n290_), .B(new_new_n26_), .Y(new_new_n307_));
  NO2        g0285(.A(new_new_n307_), .B(new_new_n306_), .Y(new_new_n308_));
  NA2        g0286(.A(i_0_), .B(i_1_), .Y(new_new_n309_));
  NO2        g0287(.A(new_new_n309_), .B(i_2_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n57_), .B(i_6_), .Y(new_new_n311_));
  NA3        g0289(.A(new_new_n311_), .B(new_new_n310_), .C(new_new_n165_), .Y(new_new_n312_));
  OAI210     g0290(.A0(new_new_n167_), .A1(new_new_n144_), .B0(new_new_n312_), .Y(new_new_n313_));
  NO3        g0291(.A(new_new_n313_), .B(new_new_n308_), .C(new_new_n303_), .Y(new_new_n314_));
  NO2        g0292(.A(i_3_), .B(i_10_), .Y(new_new_n315_));
  NA3        g0293(.A(new_new_n315_), .B(new_new_n37_), .C(new_new_n42_), .Y(new_new_n316_));
  NO2        g0294(.A(i_2_), .B(new_new_n102_), .Y(new_new_n317_));
  NA2        g0295(.A(i_1_), .B(new_new_n34_), .Y(new_new_n318_));
  NO2        g0296(.A(new_new_n318_), .B(i_8_), .Y(new_new_n319_));
  NOi21      g0297(.An(new_new_n225_), .B(new_new_n104_), .Y(new_new_n320_));
  NA3        g0298(.A(new_new_n320_), .B(new_new_n319_), .C(new_new_n317_), .Y(new_new_n321_));
  AN2        g0299(.A(i_3_), .B(i_10_), .Y(new_new_n322_));
  NA4        g0300(.A(new_new_n322_), .B(new_new_n202_), .C(new_new_n179_), .D(new_new_n177_), .Y(new_new_n323_));
  NO2        g0301(.A(i_5_), .B(new_new_n35_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n44_), .B(new_new_n26_), .Y(new_new_n325_));
  OR2        g0303(.A(new_new_n321_), .B(new_new_n316_), .Y(new_new_n326_));
  OAI220     g0304(.A0(new_new_n326_), .A1(i_6_), .B0(new_new_n314_), .B1(new_new_n298_), .Y(new_new_n327_));
  NO4        g0305(.A(new_new_n327_), .B(new_new_n296_), .C(new_new_n221_), .D(new_new_n170_), .Y(new_new_n328_));
  NO3        g0306(.A(new_new_n42_), .B(i_13_), .C(i_9_), .Y(new_new_n329_));
  NO2        g0307(.A(new_new_n57_), .B(new_new_n84_), .Y(new_new_n330_));
  NA2        g0308(.A(new_new_n305_), .B(new_new_n330_), .Y(new_new_n331_));
  NO3        g0309(.A(i_6_), .B(new_new_n197_), .C(i_7_), .Y(new_new_n332_));
  NA2        g0310(.A(new_new_n332_), .B(new_new_n202_), .Y(new_new_n333_));
  AOI210     g0311(.A0(new_new_n333_), .A1(new_new_n331_), .B0(new_new_n172_), .Y(new_new_n334_));
  NO2        g0312(.A(i_2_), .B(i_3_), .Y(new_new_n335_));
  OR2        g0313(.A(i_0_), .B(i_5_), .Y(new_new_n336_));
  NA2        g0314(.A(new_new_n225_), .B(new_new_n336_), .Y(new_new_n337_));
  NA4        g0315(.A(new_new_n337_), .B(new_new_n242_), .C(new_new_n335_), .D(i_1_), .Y(new_new_n338_));
  NA3        g0316(.A(new_new_n305_), .B(new_new_n300_), .C(new_new_n114_), .Y(new_new_n339_));
  NAi21      g0317(.An(i_8_), .B(i_7_), .Y(new_new_n340_));
  NO2        g0318(.A(new_new_n340_), .B(i_6_), .Y(new_new_n341_));
  NO2        g0319(.A(new_new_n159_), .B(new_new_n44_), .Y(new_new_n342_));
  NA3        g0320(.A(new_new_n342_), .B(new_new_n341_), .C(new_new_n165_), .Y(new_new_n343_));
  NA3        g0321(.A(new_new_n343_), .B(new_new_n339_), .C(new_new_n338_), .Y(new_new_n344_));
  OAI210     g0322(.A0(new_new_n344_), .A1(new_new_n334_), .B0(i_4_), .Y(new_new_n345_));
  NO2        g0323(.A(i_12_), .B(i_10_), .Y(new_new_n346_));
  NOi21      g0324(.An(i_5_), .B(i_0_), .Y(new_new_n347_));
  AOI210     g0325(.A0(i_2_), .A1(new_new_n46_), .B0(new_new_n102_), .Y(new_new_n348_));
  NO4        g0326(.A(new_new_n348_), .B(new_new_n318_), .C(new_new_n347_), .D(new_new_n130_), .Y(new_new_n349_));
  NA4        g0327(.A(new_new_n82_), .B(new_new_n34_), .C(new_new_n84_), .D(i_8_), .Y(new_new_n350_));
  NA2        g0328(.A(new_new_n349_), .B(new_new_n346_), .Y(new_new_n351_));
  NO2        g0329(.A(i_6_), .B(i_8_), .Y(new_new_n352_));
  NOi21      g0330(.An(i_0_), .B(i_2_), .Y(new_new_n353_));
  AN2        g0331(.A(new_new_n353_), .B(new_new_n352_), .Y(new_new_n354_));
  NO2        g0332(.A(i_1_), .B(i_7_), .Y(new_new_n355_));
  AO220      g0333(.A0(new_new_n355_), .A1(new_new_n354_), .B0(new_new_n341_), .B1(new_new_n243_), .Y(new_new_n356_));
  NA3        g0334(.A(new_new_n356_), .B(new_new_n39_), .C(i_5_), .Y(new_new_n357_));
  NA3        g0335(.A(new_new_n357_), .B(new_new_n351_), .C(new_new_n345_), .Y(new_new_n358_));
  NO3        g0336(.A(new_new_n241_), .B(new_new_n44_), .C(i_1_), .Y(new_new_n359_));
  NO3        g0337(.A(new_new_n340_), .B(i_2_), .C(i_1_), .Y(new_new_n360_));
  OAI210     g0338(.A0(new_new_n360_), .A1(new_new_n359_), .B0(i_6_), .Y(new_new_n361_));
  NA3        g0339(.A(new_new_n261_), .B(new_new_n317_), .C(new_new_n197_), .Y(new_new_n362_));
  AOI210     g0340(.A0(new_new_n362_), .A1(new_new_n361_), .B0(new_new_n337_), .Y(new_new_n363_));
  NOi21      g0341(.An(new_new_n155_), .B(new_new_n105_), .Y(new_new_n364_));
  NO2        g0342(.A(new_new_n364_), .B(new_new_n126_), .Y(new_new_n365_));
  OAI210     g0343(.A0(new_new_n365_), .A1(new_new_n363_), .B0(i_3_), .Y(new_new_n366_));
  INV        g0344(.A(new_new_n82_), .Y(new_new_n367_));
  NO2        g0345(.A(new_new_n309_), .B(new_new_n79_), .Y(new_new_n368_));
  NA2        g0346(.A(new_new_n368_), .B(new_new_n134_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n93_), .B(new_new_n197_), .Y(new_new_n370_));
  NA3        g0348(.A(new_new_n320_), .B(new_new_n370_), .C(new_new_n61_), .Y(new_new_n371_));
  AOI210     g0349(.A0(new_new_n371_), .A1(new_new_n369_), .B0(new_new_n367_), .Y(new_new_n372_));
  NO2        g0350(.A(new_new_n197_), .B(i_9_), .Y(new_new_n373_));
  NA3        g0351(.A(new_new_n373_), .B(new_new_n210_), .C(new_new_n159_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n374_), .B(new_new_n44_), .Y(new_new_n375_));
  NO3        g0353(.A(new_new_n375_), .B(new_new_n372_), .C(new_new_n308_), .Y(new_new_n376_));
  AOI210     g0354(.A0(new_new_n376_), .A1(new_new_n366_), .B0(new_new_n164_), .Y(new_new_n377_));
  AOI210     g0355(.A0(new_new_n358_), .A1(new_new_n329_), .B0(new_new_n377_), .Y(new_new_n378_));
  NOi32      g0356(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n379_));
  INV        g0357(.A(new_new_n379_), .Y(new_new_n380_));
  NAi21      g0358(.An(i_0_), .B(i_6_), .Y(new_new_n381_));
  NAi21      g0359(.An(i_1_), .B(i_5_), .Y(new_new_n382_));
  NA2        g0360(.A(new_new_n382_), .B(new_new_n381_), .Y(new_new_n383_));
  NA2        g0361(.A(new_new_n383_), .B(new_new_n25_), .Y(new_new_n384_));
  OAI210     g0362(.A0(new_new_n384_), .A1(new_new_n161_), .B0(new_new_n255_), .Y(new_new_n385_));
  NAi41      g0363(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n386_));
  OAI220     g0364(.A0(new_new_n386_), .A1(new_new_n382_), .B0(new_new_n228_), .B1(new_new_n161_), .Y(new_new_n387_));
  AOI210     g0365(.A0(new_new_n386_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n388_));
  NOi32      g0366(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n389_));
  NAi21      g0367(.An(i_6_), .B(i_1_), .Y(new_new_n390_));
  NA3        g0368(.A(new_new_n390_), .B(new_new_n389_), .C(new_new_n44_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(i_0_), .Y(new_new_n392_));
  OR3        g0370(.A(new_new_n392_), .B(new_new_n388_), .C(new_new_n387_), .Y(new_new_n393_));
  NO2        g0371(.A(i_1_), .B(new_new_n102_), .Y(new_new_n394_));
  NAi21      g0372(.An(i_3_), .B(i_4_), .Y(new_new_n395_));
  NO2        g0373(.A(new_new_n395_), .B(i_9_), .Y(new_new_n396_));
  AN2        g0374(.A(i_6_), .B(i_7_), .Y(new_new_n397_));
  OAI210     g0375(.A0(new_new_n397_), .A1(new_new_n394_), .B0(new_new_n396_), .Y(new_new_n398_));
  NA2        g0376(.A(i_2_), .B(i_7_), .Y(new_new_n399_));
  NO2        g0377(.A(new_new_n395_), .B(i_10_), .Y(new_new_n400_));
  NA3        g0378(.A(new_new_n400_), .B(new_new_n399_), .C(new_new_n253_), .Y(new_new_n401_));
  AOI210     g0379(.A0(new_new_n401_), .A1(new_new_n398_), .B0(new_new_n189_), .Y(new_new_n402_));
  AOI210     g0380(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n403_));
  OAI210     g0381(.A0(new_new_n403_), .A1(new_new_n192_), .B0(new_new_n400_), .Y(new_new_n404_));
  AOI220     g0382(.A0(new_new_n400_), .A1(new_new_n355_), .B0(new_new_n247_), .B1(new_new_n192_), .Y(new_new_n405_));
  AOI210     g0383(.A0(new_new_n405_), .A1(new_new_n404_), .B0(i_5_), .Y(new_new_n406_));
  NO4        g0384(.A(new_new_n406_), .B(new_new_n402_), .C(new_new_n393_), .D(new_new_n385_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n380_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n409_));
  AN2        g0387(.A(i_12_), .B(i_5_), .Y(new_new_n410_));
  NO2        g0388(.A(i_4_), .B(new_new_n26_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n411_), .B(new_new_n410_), .Y(new_new_n412_));
  NO2        g0390(.A(i_11_), .B(i_6_), .Y(new_new_n413_));
  NA3        g0391(.A(new_new_n413_), .B(new_new_n342_), .C(new_new_n233_), .Y(new_new_n414_));
  NO2        g0392(.A(new_new_n414_), .B(new_new_n412_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n251_), .B(i_5_), .Y(new_new_n416_));
  NO2        g0394(.A(i_5_), .B(i_10_), .Y(new_new_n417_));
  AOI220     g0395(.A0(new_new_n417_), .A1(new_new_n282_), .B0(new_new_n416_), .B1(new_new_n202_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n145_), .B(new_new_n43_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n418_), .Y(new_new_n420_));
  OAI210     g0398(.A0(new_new_n420_), .A1(new_new_n415_), .B0(new_new_n409_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n35_), .B(new_new_n25_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n151_), .B(new_new_n84_), .Y(new_new_n423_));
  OAI210     g0401(.A0(new_new_n423_), .A1(new_new_n415_), .B0(new_new_n422_), .Y(new_new_n424_));
  NO3        g0402(.A(new_new_n84_), .B(new_new_n46_), .C(i_9_), .Y(new_new_n425_));
  NO2        g0403(.A(i_3_), .B(new_new_n102_), .Y(new_new_n426_));
  NO2        g0404(.A(i_11_), .B(i_12_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n417_), .B(new_new_n245_), .Y(new_new_n428_));
  NA3        g0406(.A(new_new_n114_), .B(new_new_n39_), .C(i_11_), .Y(new_new_n429_));
  OAI220     g0407(.A0(new_new_n429_), .A1(new_new_n228_), .B0(new_new_n428_), .B1(new_new_n350_), .Y(new_new_n430_));
  NAi21      g0408(.An(i_13_), .B(i_0_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n431_), .B(new_new_n248_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n430_), .B(new_new_n432_), .Y(new_new_n433_));
  NA3        g0411(.A(new_new_n433_), .B(new_new_n424_), .C(new_new_n421_), .Y(new_new_n434_));
  NA2        g0412(.A(new_new_n42_), .B(new_new_n233_), .Y(new_new_n435_));
  NO3        g0413(.A(i_1_), .B(i_12_), .C(new_new_n84_), .Y(new_new_n436_));
  NO2        g0414(.A(i_0_), .B(i_11_), .Y(new_new_n437_));
  AN2        g0415(.A(i_1_), .B(i_6_), .Y(new_new_n438_));
  NOi21      g0416(.An(i_2_), .B(i_12_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n439_), .B(new_new_n438_), .Y(new_new_n440_));
  NO2        g0418(.A(new_new_n440_), .B(new_new_n1146_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n143_), .B(i_9_), .Y(new_new_n442_));
  NO2        g0420(.A(new_new_n442_), .B(i_4_), .Y(new_new_n443_));
  NA2        g0421(.A(new_new_n441_), .B(new_new_n443_), .Y(new_new_n444_));
  NAi21      g0422(.An(i_9_), .B(i_4_), .Y(new_new_n445_));
  OR2        g0423(.A(i_13_), .B(i_10_), .Y(new_new_n446_));
  NO3        g0424(.A(new_new_n446_), .B(new_new_n119_), .C(new_new_n445_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n175_), .B(new_new_n125_), .Y(new_new_n448_));
  OR2        g0426(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n449_));
  NO2        g0427(.A(new_new_n102_), .B(new_new_n25_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n297_), .B(new_new_n450_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n290_), .B(new_new_n217_), .Y(new_new_n452_));
  OAI220     g0430(.A0(new_new_n452_), .A1(new_new_n449_), .B0(new_new_n451_), .B1(new_new_n364_), .Y(new_new_n453_));
  INV        g0431(.A(new_new_n453_), .Y(new_new_n454_));
  AOI210     g0432(.A0(new_new_n454_), .A1(new_new_n444_), .B0(new_new_n26_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n339_), .B(new_new_n338_), .Y(new_new_n456_));
  AOI220     g0434(.A0(new_new_n311_), .A1(new_new_n301_), .B0(new_new_n305_), .B1(new_new_n330_), .Y(new_new_n457_));
  NO2        g0435(.A(new_new_n457_), .B(new_new_n172_), .Y(new_new_n458_));
  NO2        g0436(.A(new_new_n186_), .B(new_new_n84_), .Y(new_new_n459_));
  AOI220     g0437(.A0(new_new_n459_), .A1(new_new_n310_), .B0(new_new_n292_), .B1(new_new_n217_), .Y(new_new_n460_));
  NO2        g0438(.A(new_new_n460_), .B(new_new_n299_), .Y(new_new_n461_));
  NO3        g0439(.A(new_new_n461_), .B(new_new_n458_), .C(new_new_n456_), .Y(new_new_n462_));
  NA2        g0440(.A(new_new_n200_), .B(new_new_n97_), .Y(new_new_n463_));
  NA3        g0441(.A(new_new_n342_), .B(new_new_n165_), .C(new_new_n84_), .Y(new_new_n464_));
  AOI210     g0442(.A0(new_new_n464_), .A1(new_new_n463_), .B0(new_new_n340_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n197_), .B(i_10_), .Y(new_new_n466_));
  NA3        g0444(.A(new_new_n267_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n467_));
  NA2        g0445(.A(new_new_n311_), .B(new_new_n243_), .Y(new_new_n468_));
  OAI220     g0446(.A0(new_new_n468_), .A1(new_new_n186_), .B0(new_new_n467_), .B1(new_new_n466_), .Y(new_new_n469_));
  NO2        g0447(.A(i_3_), .B(new_new_n46_), .Y(new_new_n470_));
  NA3        g0448(.A(new_new_n355_), .B(new_new_n354_), .C(new_new_n470_), .Y(new_new_n471_));
  NA2        g0449(.A(new_new_n332_), .B(new_new_n337_), .Y(new_new_n472_));
  OAI210     g0450(.A0(new_new_n472_), .A1(new_new_n193_), .B0(new_new_n471_), .Y(new_new_n473_));
  NO3        g0451(.A(new_new_n473_), .B(new_new_n469_), .C(new_new_n465_), .Y(new_new_n474_));
  AOI210     g0452(.A0(new_new_n474_), .A1(new_new_n462_), .B0(new_new_n284_), .Y(new_new_n475_));
  NO4        g0453(.A(new_new_n475_), .B(new_new_n455_), .C(new_new_n434_), .D(new_new_n408_), .Y(new_new_n476_));
  NO2        g0454(.A(new_new_n61_), .B(i_4_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n71_), .B(i_13_), .Y(new_new_n478_));
  NA3        g0456(.A(new_new_n478_), .B(new_new_n477_), .C(i_2_), .Y(new_new_n479_));
  NO2        g0457(.A(i_10_), .B(i_9_), .Y(new_new_n480_));
  NAi21      g0458(.An(i_12_), .B(i_8_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n481_), .B(i_3_), .Y(new_new_n482_));
  NA2        g0460(.A(new_new_n482_), .B(new_new_n480_), .Y(new_new_n483_));
  NO2        g0461(.A(new_new_n44_), .B(i_4_), .Y(new_new_n484_));
  NA2        g0462(.A(new_new_n484_), .B(new_new_n105_), .Y(new_new_n485_));
  OAI220     g0463(.A0(new_new_n485_), .A1(new_new_n209_), .B0(new_new_n483_), .B1(new_new_n479_), .Y(new_new_n486_));
  NA2        g0464(.A(new_new_n325_), .B(i_0_), .Y(new_new_n487_));
  NO3        g0465(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n279_), .B(new_new_n98_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n490_));
  NA2        g0468(.A(i_8_), .B(i_9_), .Y(new_new_n491_));
  AOI210     g0469(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n492_));
  OR2        g0470(.A(new_new_n492_), .B(new_new_n491_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n297_), .B(new_new_n210_), .Y(new_new_n494_));
  OAI220     g0472(.A0(new_new_n494_), .A1(new_new_n493_), .B0(new_new_n490_), .B1(new_new_n487_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n260_), .B(new_new_n324_), .Y(new_new_n496_));
  NO3        g0474(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n497_));
  AOI210     g0475(.A0(new_new_n266_), .A1(new_new_n192_), .B0(new_new_n497_), .Y(new_new_n498_));
  NA3        g0476(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n499_));
  NA4        g0477(.A(new_new_n146_), .B(new_new_n117_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n500_));
  OAI220     g0478(.A0(new_new_n500_), .A1(new_new_n499_), .B0(new_new_n498_), .B1(new_new_n496_), .Y(new_new_n501_));
  NO3        g0479(.A(new_new_n501_), .B(new_new_n495_), .C(new_new_n486_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n310_), .B(new_new_n109_), .Y(new_new_n503_));
  OR2        g0481(.A(new_new_n503_), .B(new_new_n213_), .Y(new_new_n504_));
  OA210      g0482(.A0(new_new_n374_), .A1(new_new_n102_), .B0(new_new_n312_), .Y(new_new_n505_));
  OA220      g0483(.A0(new_new_n505_), .A1(new_new_n164_), .B0(new_new_n504_), .B1(new_new_n240_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n97_), .B(i_13_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n459_), .B(new_new_n409_), .Y(new_new_n508_));
  NO2        g0486(.A(i_2_), .B(i_13_), .Y(new_new_n509_));
  NA3        g0487(.A(new_new_n509_), .B(new_new_n163_), .C(new_new_n100_), .Y(new_new_n510_));
  OAI220     g0488(.A0(new_new_n510_), .A1(new_new_n245_), .B0(new_new_n508_), .B1(new_new_n507_), .Y(new_new_n511_));
  NO3        g0489(.A(i_4_), .B(new_new_n46_), .C(i_8_), .Y(new_new_n512_));
  NO2        g0490(.A(i_6_), .B(i_7_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n513_), .B(new_new_n512_), .Y(new_new_n514_));
  NO2        g0492(.A(i_11_), .B(i_1_), .Y(new_new_n515_));
  NO2        g0493(.A(new_new_n71_), .B(i_3_), .Y(new_new_n516_));
  OR2        g0494(.A(i_11_), .B(i_8_), .Y(new_new_n517_));
  NOi21      g0495(.An(i_2_), .B(i_7_), .Y(new_new_n518_));
  NAi31      g0496(.An(new_new_n517_), .B(new_new_n518_), .C(new_new_n516_), .Y(new_new_n519_));
  NO2        g0497(.A(new_new_n446_), .B(i_6_), .Y(new_new_n520_));
  NA3        g0498(.A(new_new_n520_), .B(new_new_n477_), .C(new_new_n73_), .Y(new_new_n521_));
  NO2        g0499(.A(new_new_n521_), .B(new_new_n519_), .Y(new_new_n522_));
  NO2        g0500(.A(i_3_), .B(new_new_n197_), .Y(new_new_n523_));
  NO2        g0501(.A(i_6_), .B(i_10_), .Y(new_new_n524_));
  NA4        g0502(.A(new_new_n524_), .B(new_new_n329_), .C(new_new_n523_), .D(new_new_n245_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n525_), .B(new_new_n157_), .Y(new_new_n526_));
  NA3        g0504(.A(new_new_n254_), .B(new_new_n174_), .C(new_new_n134_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n44_), .B(new_new_n42_), .Y(new_new_n528_));
  NO2        g0506(.A(new_new_n159_), .B(i_3_), .Y(new_new_n529_));
  NAi31      g0507(.An(new_new_n528_), .B(new_new_n529_), .C(new_new_n234_), .Y(new_new_n530_));
  NA3        g0508(.A(new_new_n422_), .B(new_new_n182_), .C(new_new_n150_), .Y(new_new_n531_));
  NA3        g0509(.A(new_new_n531_), .B(new_new_n530_), .C(new_new_n527_), .Y(new_new_n532_));
  NO4        g0510(.A(new_new_n532_), .B(new_new_n526_), .C(new_new_n522_), .D(new_new_n511_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n488_), .B(new_new_n410_), .Y(new_new_n534_));
  NA2        g0512(.A(new_new_n497_), .B(new_new_n417_), .Y(new_new_n535_));
  OAI220     g0513(.A0(new_new_n535_), .A1(new_new_n232_), .B0(new_new_n534_), .B1(new_new_n55_), .Y(new_new_n536_));
  NAi21      g0514(.An(new_new_n223_), .B(new_new_n427_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n355_), .B(new_new_n225_), .Y(new_new_n538_));
  NO2        g0516(.A(new_new_n26_), .B(i_5_), .Y(new_new_n539_));
  NO2        g0517(.A(i_0_), .B(new_new_n84_), .Y(new_new_n540_));
  NA3        g0518(.A(new_new_n540_), .B(new_new_n539_), .C(new_new_n143_), .Y(new_new_n541_));
  OR3        g0519(.A(new_new_n318_), .B(new_new_n36_), .C(new_new_n44_), .Y(new_new_n542_));
  OAI220     g0520(.A0(new_new_n542_), .A1(new_new_n541_), .B0(new_new_n538_), .B1(new_new_n537_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n27_), .B(i_10_), .Y(new_new_n544_));
  NA2        g0522(.A(new_new_n329_), .B(new_new_n247_), .Y(new_new_n545_));
  OAI220     g0523(.A0(new_new_n545_), .A1(new_new_n467_), .B0(new_new_n544_), .B1(new_new_n507_), .Y(new_new_n546_));
  NA4        g0524(.A(new_new_n322_), .B(new_new_n231_), .C(new_new_n71_), .D(new_new_n245_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n547_), .B(new_new_n514_), .Y(new_new_n548_));
  NO4        g0526(.A(new_new_n548_), .B(new_new_n546_), .C(new_new_n543_), .D(new_new_n536_), .Y(new_new_n549_));
  NA4        g0527(.A(new_new_n549_), .B(new_new_n533_), .C(new_new_n506_), .D(new_new_n502_), .Y(new_new_n550_));
  NA3        g0528(.A(new_new_n322_), .B(new_new_n179_), .C(new_new_n177_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n316_), .A1(new_new_n184_), .B0(new_new_n551_), .Y(new_new_n552_));
  AN2        g0530(.A(new_new_n301_), .B(new_new_n242_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n553_), .B(new_new_n552_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n124_), .B(new_new_n113_), .Y(new_new_n555_));
  AO220      g0533(.A0(new_new_n555_), .A1(new_new_n488_), .B0(new_new_n447_), .B1(i_6_), .Y(new_new_n556_));
  NA2        g0534(.A(new_new_n329_), .B(new_new_n166_), .Y(new_new_n557_));
  OAI210     g0535(.A0(new_new_n557_), .A1(new_new_n240_), .B0(new_new_n323_), .Y(new_new_n558_));
  AOI220     g0536(.A0(new_new_n558_), .A1(new_new_n341_), .B0(new_new_n556_), .B1(new_new_n325_), .Y(new_new_n559_));
  NA4        g0537(.A(new_new_n478_), .B(new_new_n477_), .C(new_new_n207_), .D(i_2_), .Y(new_new_n560_));
  INV        g0538(.A(new_new_n560_), .Y(new_new_n561_));
  NA2        g0539(.A(new_new_n410_), .B(new_new_n233_), .Y(new_new_n562_));
  NA2        g0540(.A(new_new_n379_), .B(new_new_n71_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n397_), .B(new_new_n389_), .Y(new_new_n564_));
  AO210      g0542(.A0(new_new_n563_), .A1(new_new_n562_), .B0(new_new_n564_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n34_), .B(i_8_), .Y(new_new_n566_));
  INV        g0544(.A(new_new_n447_), .Y(new_new_n567_));
  NA2        g0545(.A(new_new_n567_), .B(new_new_n565_), .Y(new_new_n568_));
  AOI210     g0546(.A0(new_new_n561_), .A1(new_new_n208_), .B0(new_new_n568_), .Y(new_new_n569_));
  NA2        g0547(.A(new_new_n267_), .B(new_new_n62_), .Y(new_new_n570_));
  OAI210     g0548(.A0(i_8_), .A1(new_new_n570_), .B0(new_new_n136_), .Y(new_new_n571_));
  AOI210     g0549(.A0(new_new_n198_), .A1(i_9_), .B0(new_new_n278_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n572_), .B(new_new_n203_), .Y(new_new_n573_));
  OR2        g0551(.A(new_new_n186_), .B(i_4_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n574_), .B(new_new_n84_), .Y(new_new_n575_));
  AOI220     g0553(.A0(new_new_n575_), .A1(new_new_n573_), .B0(new_new_n571_), .B1(new_new_n448_), .Y(new_new_n576_));
  NA4        g0554(.A(new_new_n576_), .B(new_new_n569_), .C(new_new_n559_), .D(new_new_n554_), .Y(new_new_n577_));
  NA2        g0555(.A(new_new_n416_), .B(new_new_n310_), .Y(new_new_n578_));
  OAI210     g0556(.A0(new_new_n412_), .A1(new_new_n171_), .B0(new_new_n578_), .Y(new_new_n579_));
  NO2        g0557(.A(i_12_), .B(new_new_n197_), .Y(new_new_n580_));
  NA2        g0558(.A(new_new_n580_), .B(new_new_n233_), .Y(new_new_n581_));
  NA3        g0559(.A(new_new_n524_), .B(new_new_n177_), .C(new_new_n27_), .Y(new_new_n582_));
  NO3        g0560(.A(new_new_n582_), .B(new_new_n581_), .C(new_new_n503_), .Y(new_new_n583_));
  NOi31      g0561(.An(new_new_n332_), .B(new_new_n446_), .C(new_new_n36_), .Y(new_new_n584_));
  OAI210     g0562(.A0(new_new_n584_), .A1(new_new_n583_), .B0(new_new_n579_), .Y(new_new_n585_));
  NO2        g0563(.A(i_8_), .B(i_7_), .Y(new_new_n586_));
  OAI210     g0564(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n587_));
  NA2        g0565(.A(new_new_n587_), .B(new_new_n231_), .Y(new_new_n588_));
  AOI220     g0566(.A0(new_new_n342_), .A1(new_new_n37_), .B0(new_new_n243_), .B1(new_new_n212_), .Y(new_new_n589_));
  OAI220     g0567(.A0(new_new_n589_), .A1(new_new_n574_), .B0(new_new_n588_), .B1(new_new_n251_), .Y(new_new_n590_));
  NA2        g0568(.A(new_new_n42_), .B(i_10_), .Y(new_new_n591_));
  NO2        g0569(.A(new_new_n591_), .B(i_6_), .Y(new_new_n592_));
  NA3        g0570(.A(new_new_n592_), .B(new_new_n590_), .C(new_new_n586_), .Y(new_new_n593_));
  AOI220     g0571(.A0(new_new_n459_), .A1(new_new_n342_), .B0(new_new_n256_), .B1(new_new_n253_), .Y(new_new_n594_));
  OAI220     g0572(.A0(new_new_n594_), .A1(new_new_n275_), .B0(new_new_n507_), .B1(new_new_n135_), .Y(new_new_n595_));
  NA2        g0573(.A(new_new_n595_), .B(new_new_n278_), .Y(new_new_n596_));
  NOi31      g0574(.An(new_new_n305_), .B(new_new_n316_), .C(new_new_n184_), .Y(new_new_n597_));
  NA3        g0575(.A(new_new_n322_), .B(new_new_n177_), .C(new_new_n97_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n229_), .B(new_new_n42_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n159_), .B(i_5_), .Y(new_new_n600_));
  NA3        g0578(.A(new_new_n600_), .B(new_new_n435_), .C(new_new_n335_), .Y(new_new_n601_));
  OAI210     g0579(.A0(new_new_n601_), .A1(new_new_n599_), .B0(new_new_n598_), .Y(new_new_n602_));
  OAI210     g0580(.A0(new_new_n602_), .A1(new_new_n597_), .B0(new_new_n497_), .Y(new_new_n603_));
  NA4        g0581(.A(new_new_n603_), .B(new_new_n596_), .C(new_new_n593_), .D(new_new_n585_), .Y(new_new_n604_));
  NA3        g0582(.A(new_new_n225_), .B(new_new_n69_), .C(new_new_n42_), .Y(new_new_n605_));
  NA2        g0583(.A(new_new_n297_), .B(new_new_n82_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n605_), .A1(new_new_n369_), .B0(new_new_n606_), .Y(new_new_n607_));
  NA2        g0585(.A(new_new_n311_), .B(new_new_n301_), .Y(new_new_n608_));
  NO2        g0586(.A(new_new_n608_), .B(new_new_n176_), .Y(new_new_n609_));
  NA2        g0587(.A(new_new_n231_), .B(new_new_n230_), .Y(new_new_n610_));
  NA2        g0588(.A(new_new_n480_), .B(new_new_n229_), .Y(new_new_n611_));
  NO2        g0589(.A(new_new_n610_), .B(new_new_n611_), .Y(new_new_n612_));
  AOI210     g0590(.A0(new_new_n390_), .A1(new_new_n44_), .B0(new_new_n394_), .Y(new_new_n613_));
  NA2        g0591(.A(i_0_), .B(new_new_n46_), .Y(new_new_n614_));
  NA3        g0592(.A(new_new_n580_), .B(new_new_n288_), .C(new_new_n614_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n613_), .B(new_new_n615_), .Y(new_new_n616_));
  NO4        g0594(.A(new_new_n616_), .B(new_new_n612_), .C(new_new_n609_), .D(new_new_n607_), .Y(new_new_n617_));
  NO4        g0595(.A(new_new_n261_), .B(new_new_n40_), .C(i_2_), .D(new_new_n46_), .Y(new_new_n618_));
  NO3        g0596(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n241_), .B(new_new_n34_), .Y(new_new_n620_));
  AN2        g0598(.A(new_new_n620_), .B(new_new_n619_), .Y(new_new_n621_));
  OA210      g0599(.A0(new_new_n621_), .A1(new_new_n618_), .B0(new_new_n379_), .Y(new_new_n622_));
  NO2        g0600(.A(new_new_n446_), .B(i_1_), .Y(new_new_n623_));
  NOi31      g0601(.An(new_new_n623_), .B(new_new_n489_), .C(new_new_n71_), .Y(new_new_n624_));
  AN4        g0602(.A(new_new_n624_), .B(new_new_n443_), .C(new_new_n539_), .D(i_2_), .Y(new_new_n625_));
  NO2        g0603(.A(new_new_n457_), .B(new_new_n180_), .Y(new_new_n626_));
  NO3        g0604(.A(new_new_n626_), .B(new_new_n625_), .C(new_new_n622_), .Y(new_new_n627_));
  NOi21      g0605(.An(i_10_), .B(i_6_), .Y(new_new_n628_));
  NO2        g0606(.A(new_new_n84_), .B(new_new_n25_), .Y(new_new_n629_));
  AOI220     g0607(.A0(new_new_n297_), .A1(new_new_n629_), .B0(new_new_n288_), .B1(new_new_n628_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n630_), .B(new_new_n487_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n332_), .B(new_new_n166_), .Y(new_new_n633_));
  AOI220     g0611(.A0(new_new_n633_), .A1(new_new_n468_), .B0(new_new_n187_), .B1(new_new_n185_), .Y(new_new_n634_));
  NO2        g0612(.A(new_new_n202_), .B(new_new_n35_), .Y(new_new_n635_));
  NOi31      g0613(.An(new_new_n147_), .B(new_new_n635_), .C(new_new_n350_), .Y(new_new_n636_));
  NO3        g0614(.A(new_new_n636_), .B(new_new_n634_), .C(new_new_n631_), .Y(new_new_n637_));
  NO2        g0615(.A(new_new_n563_), .B(new_new_n405_), .Y(new_new_n638_));
  INV        g0616(.A(new_new_n335_), .Y(new_new_n639_));
  NO2        g0617(.A(i_12_), .B(new_new_n84_), .Y(new_new_n640_));
  NA3        g0618(.A(new_new_n640_), .B(new_new_n288_), .C(new_new_n614_), .Y(new_new_n641_));
  NA3        g0619(.A(new_new_n413_), .B(new_new_n297_), .C(new_new_n225_), .Y(new_new_n642_));
  AOI210     g0620(.A0(new_new_n642_), .A1(new_new_n641_), .B0(new_new_n639_), .Y(new_new_n643_));
  NA2        g0621(.A(new_new_n177_), .B(i_0_), .Y(new_new_n644_));
  NO3        g0622(.A(new_new_n644_), .B(new_new_n361_), .C(new_new_n316_), .Y(new_new_n645_));
  OR2        g0623(.A(i_2_), .B(i_5_), .Y(new_new_n646_));
  OR2        g0624(.A(new_new_n646_), .B(new_new_n438_), .Y(new_new_n647_));
  AOI210     g0625(.A0(new_new_n399_), .A1(new_new_n253_), .B0(new_new_n202_), .Y(new_new_n648_));
  AOI210     g0626(.A0(new_new_n648_), .A1(new_new_n647_), .B0(new_new_n537_), .Y(new_new_n649_));
  NO4        g0627(.A(new_new_n649_), .B(new_new_n645_), .C(new_new_n643_), .D(new_new_n638_), .Y(new_new_n650_));
  NA4        g0628(.A(new_new_n650_), .B(new_new_n637_), .C(new_new_n627_), .D(new_new_n617_), .Y(new_new_n651_));
  NO4        g0629(.A(new_new_n651_), .B(new_new_n604_), .C(new_new_n577_), .D(new_new_n550_), .Y(new_new_n652_));
  NA4        g0630(.A(new_new_n652_), .B(new_new_n476_), .C(new_new_n378_), .D(new_new_n328_), .Y(men7));
  OAI220     g0631(.A0(new_new_n544_), .A1(new_new_n119_), .B0(new_new_n93_), .B1(new_new_n52_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n109_), .B(new_new_n90_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n411_), .B(new_new_n655_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n524_), .B(new_new_n82_), .Y(new_new_n657_));
  NA2        g0635(.A(i_11_), .B(new_new_n197_), .Y(new_new_n658_));
  NA2        g0636(.A(new_new_n145_), .B(new_new_n658_), .Y(new_new_n659_));
  OAI210     g0637(.A0(new_new_n659_), .A1(new_new_n657_), .B0(new_new_n656_), .Y(new_new_n660_));
  NA3        g0638(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n245_), .B(i_4_), .Y(new_new_n662_));
  NA2        g0640(.A(new_new_n662_), .B(i_8_), .Y(new_new_n663_));
  AOI210     g0641(.A0(new_new_n663_), .A1(new_new_n106_), .B0(new_new_n661_), .Y(new_new_n664_));
  NA2        g0642(.A(i_2_), .B(new_new_n84_), .Y(new_new_n665_));
  OAI210     g0643(.A0(new_new_n87_), .A1(new_new_n207_), .B0(new_new_n208_), .Y(new_new_n666_));
  NO2        g0644(.A(i_7_), .B(new_new_n35_), .Y(new_new_n667_));
  NA2        g0645(.A(i_4_), .B(i_8_), .Y(new_new_n668_));
  AOI210     g0646(.A0(new_new_n668_), .A1(new_new_n322_), .B0(new_new_n667_), .Y(new_new_n669_));
  OAI220     g0647(.A0(new_new_n669_), .A1(new_new_n665_), .B0(new_new_n666_), .B1(i_13_), .Y(new_new_n670_));
  NO4        g0648(.A(new_new_n670_), .B(new_new_n664_), .C(new_new_n660_), .D(new_new_n654_), .Y(new_new_n671_));
  AOI210     g0649(.A0(new_new_n130_), .A1(new_new_n60_), .B0(i_10_), .Y(new_new_n672_));
  AOI210     g0650(.A0(new_new_n672_), .A1(new_new_n245_), .B0(new_new_n163_), .Y(new_new_n673_));
  OR2        g0651(.A(i_6_), .B(i_10_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n23_), .Y(new_new_n675_));
  OR3        g0653(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n676_));
  NO3        g0654(.A(new_new_n676_), .B(i_8_), .C(new_new_n29_), .Y(new_new_n677_));
  INV        g0655(.A(new_new_n204_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n677_), .B(new_new_n675_), .Y(new_new_n679_));
  OA220      g0657(.A0(new_new_n679_), .A1(new_new_n639_), .B0(new_new_n673_), .B1(new_new_n280_), .Y(new_new_n680_));
  AOI210     g0658(.A0(new_new_n680_), .A1(new_new_n671_), .B0(new_new_n61_), .Y(new_new_n681_));
  NOi21      g0659(.An(i_11_), .B(i_7_), .Y(new_new_n682_));
  AO210      g0660(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n683_));
  NO2        g0661(.A(new_new_n683_), .B(new_new_n682_), .Y(new_new_n684_));
  NA2        g0662(.A(new_new_n684_), .B(new_new_n212_), .Y(new_new_n685_));
  NA3        g0663(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n686_));
  NAi31      g0664(.An(new_new_n686_), .B(new_new_n222_), .C(i_11_), .Y(new_new_n687_));
  AOI210     g0665(.A0(new_new_n687_), .A1(new_new_n685_), .B0(new_new_n61_), .Y(new_new_n688_));
  NA2        g0666(.A(new_new_n86_), .B(new_new_n61_), .Y(new_new_n689_));
  AO210      g0667(.A0(new_new_n689_), .A1(new_new_n405_), .B0(new_new_n38_), .Y(new_new_n690_));
  NO3        g0668(.A(new_new_n269_), .B(new_new_n214_), .C(new_new_n658_), .Y(new_new_n691_));
  OAI210     g0669(.A0(new_new_n691_), .A1(new_new_n234_), .B0(new_new_n61_), .Y(new_new_n692_));
  NA2        g0670(.A(new_new_n439_), .B(new_new_n29_), .Y(new_new_n693_));
  OR2        g0671(.A(new_new_n214_), .B(new_new_n109_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n694_), .B(new_new_n693_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n61_), .B(i_9_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(i_4_), .Y(new_new_n697_));
  NA2        g0675(.A(new_new_n697_), .B(new_new_n695_), .Y(new_new_n698_));
  NO2        g0676(.A(i_1_), .B(i_12_), .Y(new_new_n699_));
  NA3        g0677(.A(new_new_n699_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n700_));
  NA4        g0678(.A(new_new_n700_), .B(new_new_n698_), .C(new_new_n692_), .D(new_new_n690_), .Y(new_new_n701_));
  OAI210     g0679(.A0(new_new_n701_), .A1(new_new_n688_), .B0(i_6_), .Y(new_new_n702_));
  OAI210     g0680(.A0(new_new_n686_), .A1(new_new_n109_), .B0(new_new_n499_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n703_), .B(new_new_n640_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n245_), .B(new_new_n84_), .Y(new_new_n705_));
  NA3        g0683(.A(new_new_n704_), .B(new_new_n567_), .C(new_new_n490_), .Y(new_new_n706_));
  NO4        g0684(.A(new_new_n222_), .B(new_new_n130_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n707_), .B(new_new_n696_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n245_), .B(i_6_), .Y(new_new_n709_));
  NO3        g0687(.A(new_new_n674_), .B(new_new_n241_), .C(new_new_n23_), .Y(new_new_n710_));
  AOI210     g0688(.A0(i_1_), .A1(new_new_n270_), .B0(new_new_n710_), .Y(new_new_n711_));
  OAI210     g0689(.A0(new_new_n711_), .A1(new_new_n42_), .B0(new_new_n708_), .Y(new_new_n712_));
  NA3        g0690(.A(new_new_n586_), .B(i_11_), .C(new_new_n34_), .Y(new_new_n713_));
  NA3        g0691(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n714_));
  NO2        g0692(.A(new_new_n44_), .B(i_1_), .Y(new_new_n715_));
  NA3        g0693(.A(new_new_n715_), .B(new_new_n279_), .C(new_new_n42_), .Y(new_new_n716_));
  NO2        g0694(.A(new_new_n716_), .B(new_new_n714_), .Y(new_new_n717_));
  NA3        g0695(.A(new_new_n696_), .B(new_new_n335_), .C(i_6_), .Y(new_new_n718_));
  NO2        g0696(.A(new_new_n718_), .B(new_new_n23_), .Y(new_new_n719_));
  NAi21      g0697(.An(new_new_n713_), .B(new_new_n92_), .Y(new_new_n720_));
  NA2        g0698(.A(new_new_n715_), .B(new_new_n279_), .Y(new_new_n721_));
  NO2        g0699(.A(i_11_), .B(new_new_n35_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n722_), .B(new_new_n24_), .Y(new_new_n723_));
  OAI210     g0701(.A0(new_new_n723_), .A1(new_new_n721_), .B0(new_new_n720_), .Y(new_new_n724_));
  OR3        g0702(.A(new_new_n724_), .B(new_new_n719_), .C(new_new_n717_), .Y(new_new_n725_));
  NO3        g0703(.A(new_new_n725_), .B(new_new_n712_), .C(new_new_n706_), .Y(new_new_n726_));
  NO2        g0704(.A(new_new_n245_), .B(new_new_n102_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n727_), .B(new_new_n682_), .Y(new_new_n728_));
  NA2        g0706(.A(new_new_n728_), .B(i_1_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n729_), .B(new_new_n676_), .Y(new_new_n730_));
  NO2        g0708(.A(new_new_n445_), .B(new_new_n84_), .Y(new_new_n731_));
  NA2        g0709(.A(new_new_n730_), .B(new_new_n44_), .Y(new_new_n732_));
  NA2        g0710(.A(i_3_), .B(new_new_n197_), .Y(new_new_n733_));
  AOI210     g0711(.A0(new_new_n268_), .A1(new_new_n733_), .B0(new_new_n116_), .Y(new_new_n734_));
  AN2        g0712(.A(new_new_n734_), .B(new_new_n592_), .Y(new_new_n735_));
  NO2        g0713(.A(new_new_n241_), .B(new_new_n42_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n736_), .B(new_new_n325_), .C(new_new_n246_), .Y(new_new_n737_));
  NO2        g0715(.A(new_new_n119_), .B(new_new_n35_), .Y(new_new_n738_));
  NO2        g0716(.A(new_new_n738_), .B(i_6_), .Y(new_new_n739_));
  NO2        g0717(.A(new_new_n84_), .B(i_9_), .Y(new_new_n740_));
  NO2        g0718(.A(new_new_n740_), .B(new_new_n61_), .Y(new_new_n741_));
  NO2        g0719(.A(new_new_n741_), .B(new_new_n699_), .Y(new_new_n742_));
  NO4        g0720(.A(new_new_n742_), .B(new_new_n739_), .C(new_new_n737_), .D(i_4_), .Y(new_new_n743_));
  NA2        g0721(.A(i_1_), .B(i_3_), .Y(new_new_n744_));
  NO2        g0722(.A(new_new_n491_), .B(new_new_n93_), .Y(new_new_n745_));
  AOI210     g0723(.A0(new_new_n736_), .A1(new_new_n628_), .B0(new_new_n745_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n746_), .B(new_new_n744_), .Y(new_new_n747_));
  NO3        g0725(.A(new_new_n747_), .B(new_new_n743_), .C(new_new_n735_), .Y(new_new_n748_));
  NA4        g0726(.A(new_new_n748_), .B(new_new_n732_), .C(new_new_n726_), .D(new_new_n702_), .Y(new_new_n749_));
  NO3        g0727(.A(new_new_n517_), .B(i_3_), .C(i_7_), .Y(new_new_n750_));
  NOi21      g0728(.An(new_new_n750_), .B(i_10_), .Y(new_new_n751_));
  OA210      g0729(.A0(new_new_n751_), .A1(new_new_n254_), .B0(new_new_n84_), .Y(new_new_n752_));
  NA2        g0730(.A(new_new_n397_), .B(new_new_n396_), .Y(new_new_n753_));
  NA3        g0731(.A(new_new_n524_), .B(new_new_n566_), .C(new_new_n44_), .Y(new_new_n754_));
  NO3        g0732(.A(new_new_n518_), .B(new_new_n668_), .C(new_new_n84_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n755_), .B(new_new_n25_), .Y(new_new_n756_));
  NA3        g0734(.A(new_new_n163_), .B(new_new_n82_), .C(new_new_n84_), .Y(new_new_n757_));
  NA4        g0735(.A(new_new_n757_), .B(new_new_n756_), .C(new_new_n754_), .D(new_new_n753_), .Y(new_new_n758_));
  OAI210     g0736(.A0(new_new_n758_), .A1(new_new_n752_), .B0(i_1_), .Y(new_new_n759_));
  AOI210     g0737(.A0(new_new_n279_), .A1(new_new_n98_), .B0(i_1_), .Y(new_new_n760_));
  NO2        g0738(.A(new_new_n395_), .B(i_2_), .Y(new_new_n761_));
  NA2        g0739(.A(new_new_n761_), .B(new_new_n760_), .Y(new_new_n762_));
  OAI210     g0740(.A0(new_new_n718_), .A1(new_new_n481_), .B0(new_new_n762_), .Y(new_new_n763_));
  INV        g0741(.A(new_new_n763_), .Y(new_new_n764_));
  AOI210     g0742(.A0(new_new_n764_), .A1(new_new_n759_), .B0(i_13_), .Y(new_new_n765_));
  OR2        g0743(.A(i_11_), .B(i_7_), .Y(new_new_n766_));
  NA3        g0744(.A(new_new_n766_), .B(new_new_n107_), .C(new_new_n140_), .Y(new_new_n767_));
  AOI220     g0745(.A0(new_new_n509_), .A1(new_new_n163_), .B0(new_new_n484_), .B1(new_new_n140_), .Y(new_new_n768_));
  OAI210     g0746(.A0(new_new_n768_), .A1(new_new_n42_), .B0(new_new_n767_), .Y(new_new_n769_));
  NO3        g0747(.A(new_new_n518_), .B(new_new_n586_), .C(new_new_n24_), .Y(new_new_n770_));
  AOI220     g0748(.A0(new_new_n770_), .A1(new_new_n731_), .B0(new_new_n254_), .B1(new_new_n133_), .Y(new_new_n771_));
  NO2        g0749(.A(new_new_n771_), .B(new_new_n38_), .Y(new_new_n772_));
  AOI210     g0750(.A0(new_new_n769_), .A1(new_new_n352_), .B0(new_new_n772_), .Y(new_new_n773_));
  NA2        g0751(.A(new_new_n116_), .B(new_new_n109_), .Y(new_new_n774_));
  AOI220     g0752(.A0(new_new_n774_), .A1(new_new_n70_), .B0(new_new_n413_), .B1(new_new_n715_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n775_), .B(new_new_n251_), .Y(new_new_n776_));
  AOI210     g0754(.A0(new_new_n481_), .A1(new_new_n34_), .B0(i_13_), .Y(new_new_n777_));
  NOi31      g0755(.An(new_new_n777_), .B(new_new_n657_), .C(new_new_n42_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n714_), .B(new_new_n116_), .Y(new_new_n779_));
  INV        g0757(.A(new_new_n779_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n780_), .B(new_new_n69_), .Y(new_new_n781_));
  NO3        g0759(.A(new_new_n69_), .B(new_new_n30_), .C(new_new_n102_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n26_), .B(new_new_n197_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(i_7_), .Y(new_new_n784_));
  NO3        g0762(.A(new_new_n518_), .B(new_new_n245_), .C(new_new_n84_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n785_), .A1(new_new_n784_), .B0(new_new_n782_), .Y(new_new_n786_));
  AOI220     g0764(.A0(new_new_n413_), .A1(new_new_n715_), .B0(new_new_n92_), .B1(new_new_n103_), .Y(new_new_n787_));
  OAI220     g0765(.A0(new_new_n787_), .A1(new_new_n663_), .B0(new_new_n786_), .B1(new_new_n678_), .Y(new_new_n788_));
  NO4        g0766(.A(new_new_n788_), .B(new_new_n781_), .C(new_new_n778_), .D(new_new_n776_), .Y(new_new_n789_));
  OR2        g0767(.A(i_11_), .B(i_6_), .Y(new_new_n790_));
  NA3        g0768(.A(new_new_n662_), .B(new_new_n783_), .C(i_7_), .Y(new_new_n791_));
  AOI210     g0769(.A0(new_new_n791_), .A1(new_new_n780_), .B0(new_new_n790_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n103_), .B(new_new_n783_), .Y(new_new_n793_));
  NAi21      g0771(.An(i_11_), .B(i_12_), .Y(new_new_n794_));
  NOi41      g0772(.An(new_new_n112_), .B(new_new_n794_), .C(i_13_), .D(new_new_n84_), .Y(new_new_n795_));
  NO3        g0773(.A(new_new_n518_), .B(new_new_n640_), .C(new_new_n668_), .Y(new_new_n796_));
  AOI220     g0774(.A0(new_new_n796_), .A1(new_new_n329_), .B0(new_new_n795_), .B1(new_new_n793_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n797_), .Y(new_new_n798_));
  OAI210     g0776(.A0(new_new_n798_), .A1(new_new_n792_), .B0(new_new_n61_), .Y(new_new_n799_));
  NO2        g0777(.A(i_2_), .B(i_12_), .Y(new_new_n800_));
  OAI210     g0778(.A0(new_new_n672_), .A1(new_new_n394_), .B0(new_new_n800_), .Y(new_new_n801_));
  NA2        g0779(.A(i_8_), .B(new_new_n25_), .Y(new_new_n802_));
  NO3        g0780(.A(new_new_n802_), .B(new_new_n411_), .C(new_new_n662_), .Y(new_new_n803_));
  OAI210     g0781(.A0(new_new_n803_), .A1(new_new_n396_), .B0(new_new_n394_), .Y(new_new_n804_));
  NO2        g0782(.A(new_new_n130_), .B(i_2_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n805_), .B(new_new_n699_), .Y(new_new_n806_));
  NA3        g0784(.A(new_new_n806_), .B(new_new_n804_), .C(new_new_n801_), .Y(new_new_n807_));
  NA3        g0785(.A(new_new_n807_), .B(new_new_n43_), .C(new_new_n233_), .Y(new_new_n808_));
  NA4        g0786(.A(new_new_n808_), .B(new_new_n799_), .C(new_new_n789_), .D(new_new_n773_), .Y(new_new_n809_));
  OR4        g0787(.A(new_new_n809_), .B(new_new_n765_), .C(new_new_n749_), .D(new_new_n681_), .Y(men5));
  AOI210     g0788(.A0(new_new_n728_), .A1(new_new_n282_), .B0(new_new_n448_), .Y(new_new_n811_));
  NA3        g0789(.A(new_new_n24_), .B(new_new_n800_), .C(new_new_n109_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n663_), .B(i_11_), .Y(new_new_n813_));
  OAI210     g0791(.A0(new_new_n667_), .A1(new_new_n87_), .B0(new_new_n813_), .Y(new_new_n814_));
  NA4        g0792(.A(new_new_n814_), .B(new_new_n812_), .C(new_new_n811_), .D(new_new_n567_), .Y(new_new_n815_));
  NO3        g0793(.A(i_11_), .B(new_new_n245_), .C(i_13_), .Y(new_new_n816_));
  NO2        g0794(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n817_));
  NA2        g0795(.A(i_12_), .B(i_8_), .Y(new_new_n818_));
  OAI210     g0796(.A0(new_new_n44_), .A1(i_3_), .B0(new_new_n818_), .Y(new_new_n819_));
  AOI220     g0797(.A0(new_new_n335_), .A1(new_new_n632_), .B0(new_new_n819_), .B1(new_new_n817_), .Y(new_new_n820_));
  INV        g0798(.A(new_new_n820_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n821_), .B(new_new_n815_), .Y(new_new_n822_));
  INV        g0800(.A(new_new_n174_), .Y(new_new_n823_));
  INV        g0801(.A(new_new_n254_), .Y(new_new_n824_));
  OAI210     g0802(.A0(new_new_n761_), .A1(new_new_n482_), .B0(new_new_n112_), .Y(new_new_n825_));
  AOI210     g0803(.A0(new_new_n825_), .A1(new_new_n824_), .B0(new_new_n823_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n491_), .B(new_new_n26_), .Y(new_new_n827_));
  NO2        g0805(.A(new_new_n827_), .B(new_new_n450_), .Y(new_new_n828_));
  AOI210     g0806(.A0(new_new_n31_), .A1(new_new_n34_), .B0(new_new_n446_), .Y(new_new_n829_));
  AOI210     g0807(.A0(new_new_n829_), .A1(i_2_), .B0(new_new_n826_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n194_), .B(new_new_n127_), .Y(new_new_n831_));
  OAI210     g0809(.A0(new_new_n831_), .A1(new_new_n817_), .B0(i_2_), .Y(new_new_n832_));
  NO3        g0810(.A(new_new_n683_), .B(new_new_n36_), .C(new_new_n26_), .Y(new_new_n833_));
  AOI210     g0811(.A0(new_new_n173_), .A1(new_new_n87_), .B0(new_new_n833_), .Y(new_new_n834_));
  AOI210     g0812(.A0(new_new_n834_), .A1(new_new_n832_), .B0(new_new_n197_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n204_), .B(new_new_n207_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n153_), .B(new_new_n658_), .Y(new_new_n837_));
  AOI210     g0815(.A0(new_new_n837_), .A1(new_new_n836_), .B0(new_new_n399_), .Y(new_new_n838_));
  AOI210     g0816(.A0(new_new_n214_), .A1(new_new_n149_), .B0(new_new_n566_), .Y(new_new_n839_));
  OAI210     g0817(.A0(new_new_n839_), .A1(new_new_n234_), .B0(new_new_n450_), .Y(new_new_n840_));
  NA4        g0818(.A(new_new_n102_), .B(new_new_n322_), .C(new_new_n126_), .D(new_new_n40_), .Y(new_new_n841_));
  OAI210     g0819(.A0(new_new_n841_), .A1(i_11_), .B0(new_new_n840_), .Y(new_new_n842_));
  NO3        g0820(.A(new_new_n842_), .B(new_new_n838_), .C(new_new_n835_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n632_), .B(new_new_n28_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n816_), .B(new_new_n289_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n845_), .B(new_new_n844_), .Y(new_new_n846_));
  NO2        g0824(.A(new_new_n60_), .B(i_12_), .Y(new_new_n847_));
  NO2        g0825(.A(new_new_n847_), .B(new_new_n128_), .Y(new_new_n848_));
  NO2        g0826(.A(new_new_n848_), .B(new_new_n658_), .Y(new_new_n849_));
  AOI220     g0827(.A0(new_new_n849_), .A1(new_new_n34_), .B0(new_new_n846_), .B1(new_new_n44_), .Y(new_new_n850_));
  NA4        g0828(.A(new_new_n850_), .B(new_new_n843_), .C(new_new_n830_), .D(new_new_n822_), .Y(men6));
  NO3        g0829(.A(new_new_n265_), .B(new_new_n324_), .C(i_1_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n189_), .B(new_new_n141_), .Y(new_new_n853_));
  OAI210     g0831(.A0(new_new_n853_), .A1(new_new_n852_), .B0(new_new_n805_), .Y(new_new_n854_));
  NA4        g0832(.A(new_new_n417_), .B(new_new_n523_), .C(new_new_n69_), .D(new_new_n102_), .Y(new_new_n855_));
  INV        g0833(.A(new_new_n855_), .Y(new_new_n856_));
  NO2        g0834(.A(new_new_n228_), .B(new_new_n528_), .Y(new_new_n857_));
  NO2        g0835(.A(i_11_), .B(i_9_), .Y(new_new_n858_));
  AO210      g0836(.A0(new_new_n855_), .A1(new_new_n854_), .B0(i_12_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n400_), .B(new_new_n355_), .Y(new_new_n860_));
  NA2        g0838(.A(new_new_n640_), .B(new_new_n61_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n751_), .B(new_new_n69_), .Y(new_new_n862_));
  NA4        g0840(.A(new_new_n689_), .B(new_new_n862_), .C(new_new_n861_), .D(new_new_n860_), .Y(new_new_n863_));
  INV        g0841(.A(new_new_n201_), .Y(new_new_n864_));
  AOI220     g0842(.A0(new_new_n864_), .A1(new_new_n858_), .B0(new_new_n863_), .B1(new_new_n71_), .Y(new_new_n865_));
  INV        g0843(.A(new_new_n346_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n73_), .B(new_new_n133_), .Y(new_new_n867_));
  OAI210     g0845(.A0(new_new_n790_), .A1(i_5_), .B0(new_new_n126_), .Y(new_new_n868_));
  NA2        g0846(.A(new_new_n868_), .B(new_new_n44_), .Y(new_new_n869_));
  AOI210     g0847(.A0(new_new_n869_), .A1(new_new_n867_), .B0(new_new_n866_), .Y(new_new_n870_));
  NO3        g0848(.A(new_new_n261_), .B(new_new_n134_), .C(i_9_), .Y(new_new_n871_));
  NA2        g0849(.A(new_new_n871_), .B(new_new_n847_), .Y(new_new_n872_));
  AOI210     g0850(.A0(new_new_n872_), .A1(new_new_n564_), .B0(new_new_n189_), .Y(new_new_n873_));
  NO2        g0851(.A(new_new_n30_), .B(i_11_), .Y(new_new_n874_));
  NA3        g0852(.A(new_new_n874_), .B(new_new_n513_), .C(new_new_n417_), .Y(new_new_n875_));
  NAi32      g0853(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n876_));
  AOI210     g0854(.A0(new_new_n790_), .A1(new_new_n85_), .B0(new_new_n876_), .Y(new_new_n877_));
  OAI210     g0855(.A0(new_new_n750_), .A1(new_new_n620_), .B0(new_new_n619_), .Y(new_new_n878_));
  NAi31      g0856(.An(new_new_n877_), .B(new_new_n878_), .C(new_new_n875_), .Y(new_new_n879_));
  OR3        g0857(.A(new_new_n879_), .B(new_new_n873_), .C(new_new_n870_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n766_), .B(i_2_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n46_), .B(new_new_n35_), .Y(new_new_n882_));
  OAI210     g0860(.A0(new_new_n882_), .A1(new_new_n438_), .B0(new_new_n384_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n883_), .B(new_new_n881_), .Y(new_new_n884_));
  AO220      g0862(.A0(new_new_n383_), .A1(new_new_n373_), .B0(new_new_n425_), .B1(new_new_n658_), .Y(new_new_n885_));
  NA3        g0863(.A(new_new_n885_), .B(new_new_n266_), .C(i_7_), .Y(new_new_n886_));
  OR2        g0864(.A(new_new_n684_), .B(new_new_n482_), .Y(new_new_n887_));
  NA3        g0865(.A(new_new_n887_), .B(new_new_n148_), .C(new_new_n67_), .Y(new_new_n888_));
  OR2        g0866(.A(new_new_n535_), .B(new_new_n34_), .Y(new_new_n889_));
  NA4        g0867(.A(new_new_n889_), .B(new_new_n888_), .C(new_new_n886_), .D(new_new_n884_), .Y(new_new_n890_));
  OAI210     g0868(.A0(new_new_n705_), .A1(i_11_), .B0(new_new_n85_), .Y(new_new_n891_));
  AOI220     g0869(.A0(new_new_n891_), .A1(new_new_n619_), .B0(new_new_n857_), .B1(new_new_n784_), .Y(new_new_n892_));
  NA3        g0870(.A(new_new_n399_), .B(new_new_n247_), .C(new_new_n148_), .Y(new_new_n893_));
  OAI210     g0871(.A0(new_new_n425_), .A1(new_new_n208_), .B0(new_new_n68_), .Y(new_new_n894_));
  NA4        g0872(.A(new_new_n894_), .B(new_new_n893_), .C(new_new_n892_), .D(new_new_n666_), .Y(new_new_n895_));
  AO210      g0873(.A0(new_new_n566_), .A1(new_new_n44_), .B0(new_new_n86_), .Y(new_new_n896_));
  NA3        g0874(.A(new_new_n896_), .B(new_new_n524_), .C(new_new_n225_), .Y(new_new_n897_));
  AOI210     g0875(.A0(new_new_n482_), .A1(new_new_n480_), .B0(new_new_n618_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n674_), .B(new_new_n103_), .Y(new_new_n899_));
  OAI210     g0877(.A0(new_new_n899_), .A1(new_new_n113_), .B0(new_new_n437_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n253_), .B(new_new_n44_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n901_), .B(new_new_n647_), .Y(new_new_n902_));
  NA3        g0880(.A(new_new_n902_), .B(new_new_n346_), .C(i_7_), .Y(new_new_n903_));
  NA4        g0881(.A(new_new_n903_), .B(new_new_n900_), .C(new_new_n898_), .D(new_new_n897_), .Y(new_new_n904_));
  NO4        g0882(.A(new_new_n904_), .B(new_new_n895_), .C(new_new_n890_), .D(new_new_n880_), .Y(new_new_n905_));
  NA4        g0883(.A(new_new_n905_), .B(new_new_n865_), .C(new_new_n859_), .D(new_new_n407_), .Y(men3));
  NA2        g0884(.A(i_12_), .B(i_10_), .Y(new_new_n907_));
  NA2        g0885(.A(i_6_), .B(i_7_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n908_), .B(i_0_), .Y(new_new_n909_));
  NO2        g0887(.A(i_11_), .B(new_new_n245_), .Y(new_new_n910_));
  OAI210     g0888(.A0(new_new_n909_), .A1(new_new_n305_), .B0(new_new_n910_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n911_), .B(new_new_n197_), .Y(new_new_n912_));
  NO3        g0890(.A(new_new_n487_), .B(new_new_n90_), .C(new_new_n42_), .Y(new_new_n913_));
  OA210      g0891(.A0(new_new_n913_), .A1(new_new_n912_), .B0(new_new_n177_), .Y(new_new_n914_));
  NA3        g0892(.A(new_new_n893_), .B(new_new_n666_), .C(new_new_n398_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n915_), .B(new_new_n37_), .Y(new_new_n916_));
  NOi21      g0894(.An(new_new_n97_), .B(new_new_n828_), .Y(new_new_n917_));
  NO3        g0895(.A(new_new_n694_), .B(new_new_n491_), .C(new_new_n133_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n439_), .B(new_new_n43_), .Y(new_new_n919_));
  AN2        g0897(.A(new_new_n489_), .B(new_new_n53_), .Y(new_new_n920_));
  NO3        g0898(.A(new_new_n920_), .B(new_new_n918_), .C(new_new_n917_), .Y(new_new_n921_));
  AOI210     g0899(.A0(new_new_n921_), .A1(new_new_n916_), .B0(new_new_n46_), .Y(new_new_n922_));
  NO4        g0900(.A(new_new_n403_), .B(new_new_n410_), .C(new_new_n36_), .D(i_0_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n189_), .B(new_new_n628_), .Y(new_new_n924_));
  NOi21      g0902(.An(new_new_n924_), .B(new_new_n923_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n777_), .B(new_new_n740_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n353_), .B(new_new_n470_), .Y(new_new_n927_));
  OAI220     g0905(.A0(new_new_n927_), .A1(new_new_n926_), .B0(new_new_n925_), .B1(new_new_n61_), .Y(new_new_n928_));
  NOi21      g0906(.An(i_5_), .B(i_9_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n929_), .B(new_new_n478_), .Y(new_new_n930_));
  AOI210     g0908(.A0(new_new_n279_), .A1(new_new_n515_), .B0(new_new_n755_), .Y(new_new_n931_));
  NO3        g0909(.A(new_new_n442_), .B(new_new_n279_), .C(new_new_n71_), .Y(new_new_n932_));
  NO2        g0910(.A(new_new_n178_), .B(new_new_n149_), .Y(new_new_n933_));
  AOI210     g0911(.A0(new_new_n933_), .A1(new_new_n253_), .B0(new_new_n932_), .Y(new_new_n934_));
  OAI220     g0912(.A0(new_new_n934_), .A1(new_new_n184_), .B0(new_new_n931_), .B1(new_new_n930_), .Y(new_new_n935_));
  NO4        g0913(.A(new_new_n935_), .B(new_new_n928_), .C(new_new_n922_), .D(new_new_n914_), .Y(new_new_n936_));
  NOi21      g0914(.An(i_0_), .B(i_10_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n189_), .B(new_new_n24_), .Y(new_new_n938_));
  NO2        g0916(.A(new_new_n738_), .B(new_new_n655_), .Y(new_new_n939_));
  NO2        g0917(.A(new_new_n939_), .B(new_new_n938_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n329_), .B(new_new_n131_), .Y(new_new_n941_));
  NAi21      g0919(.An(new_new_n164_), .B(new_new_n470_), .Y(new_new_n942_));
  OAI220     g0920(.A0(new_new_n942_), .A1(new_new_n901_), .B0(new_new_n941_), .B1(new_new_n428_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n943_), .B(new_new_n940_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n629_), .B(i_0_), .Y(new_new_n945_));
  NO3        g0923(.A(new_new_n945_), .B(new_new_n412_), .C(new_new_n87_), .Y(new_new_n946_));
  NO4        g0924(.A(new_new_n646_), .B(new_new_n222_), .C(new_new_n446_), .D(new_new_n438_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n947_), .A1(i_11_), .B0(new_new_n946_), .Y(new_new_n948_));
  INV        g0926(.A(new_new_n513_), .Y(new_new_n949_));
  AN2        g0927(.A(new_new_n97_), .B(new_new_n252_), .Y(new_new_n950_));
  NA2        g0928(.A(new_new_n816_), .B(new_new_n347_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n524_), .A1(new_new_n87_), .B0(new_new_n56_), .Y(new_new_n952_));
  OAI220     g0930(.A0(new_new_n952_), .A1(new_new_n951_), .B0(new_new_n723_), .B1(new_new_n588_), .Y(new_new_n953_));
  NO2        g0931(.A(new_new_n263_), .B(new_new_n155_), .Y(new_new_n954_));
  NA2        g0932(.A(i_0_), .B(i_10_), .Y(new_new_n955_));
  INV        g0933(.A(new_new_n591_), .Y(new_new_n956_));
  NO4        g0934(.A(new_new_n116_), .B(new_new_n56_), .C(new_new_n733_), .D(i_5_), .Y(new_new_n957_));
  AO220      g0935(.A0(new_new_n957_), .A1(new_new_n956_), .B0(new_new_n954_), .B1(i_6_), .Y(new_new_n958_));
  AOI220     g0936(.A0(new_new_n353_), .A1(new_new_n99_), .B0(new_new_n189_), .B1(new_new_n82_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n623_), .B(i_4_), .Y(new_new_n960_));
  NA2        g0938(.A(new_new_n192_), .B(new_new_n207_), .Y(new_new_n961_));
  OAI220     g0939(.A0(new_new_n961_), .A1(new_new_n951_), .B0(new_new_n960_), .B1(new_new_n959_), .Y(new_new_n962_));
  NO4        g0940(.A(new_new_n962_), .B(new_new_n958_), .C(new_new_n953_), .D(new_new_n950_), .Y(new_new_n963_));
  NA3        g0941(.A(new_new_n963_), .B(new_new_n948_), .C(new_new_n944_), .Y(new_new_n964_));
  NO2        g0942(.A(new_new_n104_), .B(new_new_n35_), .Y(new_new_n965_));
  NA2        g0943(.A(i_11_), .B(i_9_), .Y(new_new_n966_));
  NO3        g0944(.A(i_12_), .B(new_new_n966_), .C(new_new_n665_), .Y(new_new_n967_));
  AO220      g0945(.A0(new_new_n967_), .A1(new_new_n965_), .B0(new_new_n281_), .B1(new_new_n86_), .Y(new_new_n968_));
  NO2        g0946(.A(new_new_n46_), .B(i_7_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n422_), .B(new_new_n182_), .Y(new_new_n970_));
  NAi41      g0948(.An(new_new_n276_), .B(new_new_n970_), .C(new_new_n496_), .D(new_new_n162_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n966_), .B(new_new_n71_), .Y(new_new_n972_));
  NO2        g0950(.A(new_new_n178_), .B(i_0_), .Y(new_new_n973_));
  INV        g0951(.A(new_new_n973_), .Y(new_new_n974_));
  NA2        g0952(.A(new_new_n513_), .B(new_new_n239_), .Y(new_new_n975_));
  AOI210     g0953(.A0(new_new_n397_), .A1(new_new_n39_), .B0(new_new_n436_), .Y(new_new_n976_));
  OAI220     g0954(.A0(new_new_n976_), .A1(new_new_n930_), .B0(new_new_n975_), .B1(new_new_n974_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n977_), .B(new_new_n971_), .C(new_new_n968_), .Y(new_new_n978_));
  NA2        g0956(.A(new_new_n722_), .B(new_new_n123_), .Y(new_new_n979_));
  NO2        g0957(.A(i_6_), .B(new_new_n979_), .Y(new_new_n980_));
  AOI210     g0958(.A0(new_new_n481_), .A1(new_new_n34_), .B0(i_3_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n174_), .B(new_new_n104_), .Y(new_new_n982_));
  NOi32      g0960(.An(new_new_n981_), .Bn(new_new_n192_), .C(new_new_n982_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n667_), .A1(new_new_n347_), .B0(new_new_n252_), .Y(new_new_n984_));
  NO2        g0962(.A(new_new_n984_), .B(new_new_n919_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n985_), .B(new_new_n983_), .C(new_new_n980_), .Y(new_new_n986_));
  NOi21      g0964(.An(i_7_), .B(i_5_), .Y(new_new_n987_));
  NOi31      g0965(.An(new_new_n987_), .B(new_new_n937_), .C(new_new_n794_), .Y(new_new_n988_));
  NA3        g0966(.A(new_new_n988_), .B(new_new_n411_), .C(i_6_), .Y(new_new_n989_));
  OA210      g0967(.A0(new_new_n982_), .A1(new_new_n564_), .B0(new_new_n989_), .Y(new_new_n990_));
  NO3        g0968(.A(new_new_n431_), .B(new_new_n386_), .C(new_new_n382_), .Y(new_new_n991_));
  NO2        g0969(.A(new_new_n273_), .B(new_new_n336_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n794_), .B(new_new_n268_), .Y(new_new_n993_));
  AOI210     g0971(.A0(new_new_n993_), .A1(new_new_n992_), .B0(new_new_n991_), .Y(new_new_n994_));
  NA4        g0972(.A(new_new_n994_), .B(new_new_n990_), .C(new_new_n986_), .D(new_new_n978_), .Y(new_new_n995_));
  NO2        g0973(.A(new_new_n938_), .B(new_new_n248_), .Y(new_new_n996_));
  AN2        g0974(.A(new_new_n352_), .B(new_new_n347_), .Y(new_new_n997_));
  AO220      g0975(.A0(new_new_n997_), .A1(new_new_n933_), .B0(new_new_n368_), .B1(new_new_n27_), .Y(new_new_n998_));
  OAI210     g0976(.A0(new_new_n998_), .A1(new_new_n996_), .B0(i_10_), .Y(new_new_n999_));
  NO2        g0977(.A(new_new_n907_), .B(new_new_n335_), .Y(new_new_n1000_));
  OA210      g0978(.A0(new_new_n513_), .A1(new_new_n231_), .B0(new_new_n512_), .Y(new_new_n1001_));
  OAI210     g0979(.A0(new_new_n1001_), .A1(new_new_n1000_), .B0(new_new_n972_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n512_), .B(new_new_n439_), .C(new_new_n43_), .Y(new_new_n1003_));
  OAI210     g0981(.A0(new_new_n942_), .A1(new_new_n949_), .B0(new_new_n1003_), .Y(new_new_n1004_));
  NO2        g0982(.A(new_new_n266_), .B(new_new_n44_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n972_), .B(new_new_n322_), .Y(new_new_n1006_));
  OAI210     g0984(.A0(new_new_n1005_), .A1(new_new_n191_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  AOI220     g0985(.A0(new_new_n1007_), .A1(new_new_n513_), .B0(new_new_n1004_), .B1(new_new_n71_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n882_), .B(new_new_n409_), .C(new_new_n705_), .Y(new_new_n1009_));
  NA2        g0987(.A(new_new_n93_), .B(new_new_n42_), .Y(new_new_n1010_));
  NO2        g0988(.A(new_new_n73_), .B(new_new_n818_), .Y(new_new_n1011_));
  AOI220     g0989(.A0(new_new_n1011_), .A1(new_new_n1010_), .B0(new_new_n177_), .B1(new_new_n655_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n1012_), .A1(new_new_n1009_), .B0(new_new_n45_), .Y(new_new_n1013_));
  NO3        g0991(.A(new_new_n646_), .B(new_new_n381_), .C(new_new_n24_), .Y(new_new_n1014_));
  AOI210     g0992(.A0(new_new_n770_), .A1(new_new_n600_), .B0(new_new_n1014_), .Y(new_new_n1015_));
  NAi21      g0993(.An(i_9_), .B(i_5_), .Y(new_new_n1016_));
  NO2        g0994(.A(new_new_n1016_), .B(new_new_n431_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n661_), .B(new_new_n106_), .Y(new_new_n1018_));
  AOI220     g0996(.A0(new_new_n1018_), .A1(i_0_), .B0(new_new_n1017_), .B1(new_new_n684_), .Y(new_new_n1019_));
  OAI220     g0997(.A0(new_new_n1019_), .A1(new_new_n84_), .B0(new_new_n1015_), .B1(new_new_n175_), .Y(new_new_n1020_));
  NO3        g0998(.A(new_new_n1020_), .B(new_new_n1013_), .C(new_new_n568_), .Y(new_new_n1021_));
  NA4        g0999(.A(new_new_n1021_), .B(new_new_n1008_), .C(new_new_n1002_), .D(new_new_n999_), .Y(new_new_n1022_));
  NO3        g1000(.A(new_new_n1022_), .B(new_new_n995_), .C(new_new_n964_), .Y(new_new_n1023_));
  NO2        g1001(.A(new_new_n937_), .B(new_new_n794_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n71_), .B(new_new_n42_), .Y(new_new_n1025_));
  INV        g1003(.A(new_new_n1025_), .Y(new_new_n1026_));
  NO3        g1004(.A(new_new_n106_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n1027_));
  AO220      g1005(.A0(new_new_n1027_), .A1(new_new_n1026_), .B0(new_new_n1024_), .B1(new_new_n177_), .Y(new_new_n1028_));
  AOI210     g1006(.A0(new_new_n861_), .A1(new_new_n753_), .B0(new_new_n982_), .Y(new_new_n1029_));
  AOI210     g1007(.A0(new_new_n1028_), .A1(new_new_n370_), .B0(new_new_n1029_), .Y(new_new_n1030_));
  NA2        g1008(.A(new_new_n805_), .B(new_new_n147_), .Y(new_new_n1031_));
  INV        g1009(.A(new_new_n1031_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n1032_), .B(new_new_n740_), .C(new_new_n71_), .Y(new_new_n1033_));
  NO2        g1011(.A(new_new_n878_), .B(new_new_n431_), .Y(new_new_n1034_));
  NA3        g1012(.A(new_new_n909_), .B(i_2_), .C(new_new_n46_), .Y(new_new_n1035_));
  NA2        g1013(.A(new_new_n910_), .B(i_9_), .Y(new_new_n1036_));
  AOI210     g1014(.A0(new_new_n1035_), .A1(new_new_n541_), .B0(new_new_n1036_), .Y(new_new_n1037_));
  OAI210     g1015(.A0(new_new_n253_), .A1(i_9_), .B0(new_new_n238_), .Y(new_new_n1038_));
  AOI210     g1016(.A0(new_new_n1038_), .A1(new_new_n945_), .B0(new_new_n155_), .Y(new_new_n1039_));
  NO3        g1017(.A(new_new_n1039_), .B(new_new_n1037_), .C(new_new_n1034_), .Y(new_new_n1040_));
  NA3        g1018(.A(new_new_n1040_), .B(new_new_n1033_), .C(new_new_n1030_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n997_), .B(new_new_n399_), .Y(new_new_n1042_));
  AOI210     g1020(.A0(new_new_n316_), .A1(new_new_n164_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  NA3        g1021(.A(new_new_n37_), .B(new_new_n28_), .C(new_new_n42_), .Y(new_new_n1044_));
  NA2        g1022(.A(new_new_n969_), .B(new_new_n529_), .Y(new_new_n1045_));
  AOI210     g1023(.A0(new_new_n1044_), .A1(new_new_n164_), .B0(new_new_n1045_), .Y(new_new_n1046_));
  NO2        g1024(.A(new_new_n1046_), .B(new_new_n1043_), .Y(new_new_n1047_));
  NO3        g1025(.A(new_new_n955_), .B(new_new_n929_), .C(new_new_n194_), .Y(new_new_n1048_));
  AOI220     g1026(.A0(new_new_n1048_), .A1(i_11_), .B0(new_new_n624_), .B1(new_new_n73_), .Y(new_new_n1049_));
  INV        g1027(.A(new_new_n225_), .Y(new_new_n1050_));
  OAI220     g1028(.A0(new_new_n581_), .A1(new_new_n141_), .B0(new_new_n709_), .B1(new_new_n678_), .Y(new_new_n1051_));
  NA3        g1029(.A(new_new_n1051_), .B(new_new_n426_), .C(new_new_n1050_), .Y(new_new_n1052_));
  NA3        g1030(.A(new_new_n1052_), .B(new_new_n1049_), .C(new_new_n1047_), .Y(new_new_n1053_));
  NO2        g1031(.A(new_new_n251_), .B(new_new_n93_), .Y(new_new_n1054_));
  AOI210     g1032(.A0(new_new_n1054_), .A1(new_new_n1024_), .B0(new_new_n110_), .Y(new_new_n1055_));
  AOI220     g1033(.A0(new_new_n987_), .A1(new_new_n529_), .B0(new_new_n909_), .B1(new_new_n165_), .Y(new_new_n1056_));
  NA2        g1034(.A(new_new_n373_), .B(new_new_n179_), .Y(new_new_n1057_));
  OA220      g1035(.A0(new_new_n1057_), .A1(new_new_n1056_), .B0(new_new_n1055_), .B1(i_5_), .Y(new_new_n1058_));
  AOI210     g1036(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n178_), .Y(new_new_n1059_));
  NA2        g1037(.A(new_new_n1059_), .B(new_new_n1001_), .Y(new_new_n1060_));
  NA3        g1038(.A(new_new_n675_), .B(new_new_n189_), .C(new_new_n82_), .Y(new_new_n1061_));
  NA2        g1039(.A(new_new_n1061_), .B(new_new_n598_), .Y(new_new_n1062_));
  NO3        g1040(.A(new_new_n919_), .B(new_new_n52_), .C(new_new_n46_), .Y(new_new_n1063_));
  NA3        g1041(.A(new_new_n534_), .B(new_new_n527_), .C(new_new_n510_), .Y(new_new_n1064_));
  NO3        g1042(.A(new_new_n1064_), .B(new_new_n1063_), .C(new_new_n1062_), .Y(new_new_n1065_));
  NA3        g1043(.A(new_new_n417_), .B(new_new_n174_), .C(new_new_n173_), .Y(new_new_n1066_));
  NA3        g1044(.A(new_new_n969_), .B(new_new_n305_), .C(new_new_n238_), .Y(new_new_n1067_));
  NA2        g1045(.A(new_new_n1067_), .B(new_new_n1066_), .Y(new_new_n1068_));
  NA3        g1046(.A(new_new_n417_), .B(new_new_n354_), .C(new_new_n229_), .Y(new_new_n1069_));
  INV        g1047(.A(new_new_n1069_), .Y(new_new_n1070_));
  NOi31      g1048(.An(new_new_n416_), .B(new_new_n1025_), .C(new_new_n248_), .Y(new_new_n1071_));
  NO3        g1049(.A(new_new_n966_), .B(new_new_n225_), .C(new_new_n194_), .Y(new_new_n1072_));
  NO4        g1050(.A(new_new_n1072_), .B(new_new_n1071_), .C(new_new_n1070_), .D(new_new_n1068_), .Y(new_new_n1073_));
  NA4        g1051(.A(new_new_n1073_), .B(new_new_n1065_), .C(new_new_n1060_), .D(new_new_n1058_), .Y(new_new_n1074_));
  AOI210     g1052(.A0(new_new_n623_), .A1(new_new_n580_), .B0(new_new_n677_), .Y(new_new_n1075_));
  NO3        g1053(.A(new_new_n1075_), .B(new_new_n614_), .C(new_new_n367_), .Y(new_new_n1076_));
  NO2        g1054(.A(new_new_n84_), .B(i_5_), .Y(new_new_n1077_));
  NA3        g1055(.A(new_new_n910_), .B(new_new_n111_), .C(new_new_n126_), .Y(new_new_n1078_));
  INV        g1056(.A(new_new_n1078_), .Y(new_new_n1079_));
  AOI210     g1057(.A0(new_new_n1079_), .A1(new_new_n1077_), .B0(new_new_n1076_), .Y(new_new_n1080_));
  NA3        g1058(.A(new_new_n322_), .B(i_5_), .C(new_new_n197_), .Y(new_new_n1081_));
  NAi31      g1059(.An(new_new_n250_), .B(new_new_n1081_), .C(new_new_n251_), .Y(new_new_n1082_));
  NO4        g1060(.A(new_new_n248_), .B(new_new_n216_), .C(i_0_), .D(i_12_), .Y(new_new_n1083_));
  AOI220     g1061(.A0(new_new_n1083_), .A1(new_new_n1082_), .B0(new_new_n856_), .B1(new_new_n179_), .Y(new_new_n1084_));
  BUFFER     g1062(.A(new_new_n155_), .Y(new_new_n1085_));
  NO4        g1063(.A(new_new_n1085_), .B(i_12_), .C(new_new_n713_), .D(new_new_n133_), .Y(new_new_n1086_));
  NA2        g1064(.A(new_new_n1086_), .B(new_new_n225_), .Y(new_new_n1087_));
  NA3        g1065(.A(new_new_n99_), .B(new_new_n628_), .C(i_11_), .Y(new_new_n1088_));
  NO2        g1066(.A(new_new_n1088_), .B(new_new_n157_), .Y(new_new_n1089_));
  NA2        g1067(.A(new_new_n987_), .B(new_new_n509_), .Y(new_new_n1090_));
  NA2        g1068(.A(new_new_n62_), .B(new_new_n102_), .Y(new_new_n1091_));
  OAI220     g1069(.A0(new_new_n1091_), .A1(new_new_n1081_), .B0(new_new_n1090_), .B1(new_new_n741_), .Y(new_new_n1092_));
  AOI210     g1070(.A0(new_new_n1092_), .A1(new_new_n973_), .B0(new_new_n1089_), .Y(new_new_n1093_));
  NA4        g1071(.A(new_new_n1093_), .B(new_new_n1087_), .C(new_new_n1084_), .D(new_new_n1080_), .Y(new_new_n1094_));
  NO4        g1072(.A(new_new_n1094_), .B(new_new_n1074_), .C(new_new_n1053_), .D(new_new_n1041_), .Y(new_new_n1095_));
  OAI210     g1073(.A0(new_new_n881_), .A1(new_new_n874_), .B0(new_new_n35_), .Y(new_new_n1096_));
  NA3        g1074(.A(new_new_n981_), .B(new_new_n394_), .C(i_5_), .Y(new_new_n1097_));
  NA3        g1075(.A(new_new_n1097_), .B(new_new_n1096_), .C(new_new_n673_), .Y(new_new_n1098_));
  NA2        g1076(.A(new_new_n1098_), .B(new_new_n212_), .Y(new_new_n1099_));
  AN2        g1077(.A(new_new_n766_), .B(new_new_n395_), .Y(new_new_n1100_));
  NA2        g1078(.A(new_new_n190_), .B(new_new_n192_), .Y(new_new_n1101_));
  AO210      g1079(.A0(new_new_n1100_), .A1(new_new_n31_), .B0(new_new_n1101_), .Y(new_new_n1102_));
  OAI210     g1080(.A0(new_new_n677_), .A1(new_new_n675_), .B0(new_new_n335_), .Y(new_new_n1103_));
  NAi31      g1081(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1104_));
  AOI210     g1082(.A0(new_new_n119_), .A1(new_new_n68_), .B0(new_new_n1104_), .Y(new_new_n1105_));
  NO2        g1083(.A(new_new_n1105_), .B(new_new_n710_), .Y(new_new_n1106_));
  NA3        g1084(.A(new_new_n1106_), .B(new_new_n1103_), .C(new_new_n1102_), .Y(new_new_n1107_));
  NO2        g1085(.A(new_new_n499_), .B(new_new_n279_), .Y(new_new_n1108_));
  NO4        g1086(.A(new_new_n241_), .B(new_new_n146_), .C(new_new_n744_), .D(new_new_n35_), .Y(new_new_n1109_));
  NO3        g1087(.A(new_new_n1109_), .B(new_new_n1108_), .C(new_new_n947_), .Y(new_new_n1110_));
  OAI210     g1088(.A0(new_new_n1088_), .A1(new_new_n149_), .B0(new_new_n1110_), .Y(new_new_n1111_));
  AOI210     g1089(.A0(new_new_n1107_), .A1(new_new_n46_), .B0(new_new_n1111_), .Y(new_new_n1112_));
  AOI210     g1090(.A0(new_new_n1112_), .A1(new_new_n1099_), .B0(new_new_n71_), .Y(new_new_n1113_));
  NO2        g1091(.A(new_new_n621_), .B(new_new_n406_), .Y(new_new_n1114_));
  NO2        g1092(.A(new_new_n1114_), .B(new_new_n823_), .Y(new_new_n1115_));
  OAI210     g1093(.A0(new_new_n78_), .A1(new_new_n52_), .B0(new_new_n109_), .Y(new_new_n1116_));
  NA2        g1094(.A(new_new_n1116_), .B(new_new_n74_), .Y(new_new_n1117_));
  AOI210     g1095(.A0(new_new_n1059_), .A1(new_new_n969_), .B0(new_new_n988_), .Y(new_new_n1118_));
  AOI210     g1096(.A0(new_new_n1118_), .A1(new_new_n1117_), .B0(new_new_n744_), .Y(new_new_n1119_));
  INV        g1097(.A(new_new_n55_), .Y(new_new_n1120_));
  AOI220     g1098(.A0(new_new_n1120_), .A1(new_new_n74_), .B0(new_new_n368_), .B1(new_new_n265_), .Y(new_new_n1121_));
  NO2        g1099(.A(new_new_n1121_), .B(new_new_n245_), .Y(new_new_n1122_));
  NA3        g1100(.A(new_new_n97_), .B(new_new_n324_), .C(new_new_n29_), .Y(new_new_n1123_));
  INV        g1101(.A(new_new_n1123_), .Y(new_new_n1124_));
  NO3        g1102(.A(new_new_n1124_), .B(new_new_n1122_), .C(new_new_n1119_), .Y(new_new_n1125_));
  OAI210     g1103(.A0(new_new_n281_), .A1(new_new_n160_), .B0(new_new_n87_), .Y(new_new_n1126_));
  NA3        g1104(.A(new_new_n827_), .B(new_new_n305_), .C(new_new_n78_), .Y(new_new_n1127_));
  AOI210     g1105(.A0(new_new_n1127_), .A1(new_new_n1126_), .B0(i_11_), .Y(new_new_n1128_));
  NA2        g1106(.A(new_new_n668_), .B(new_new_n222_), .Y(new_new_n1129_));
  OAI210     g1107(.A0(new_new_n1129_), .A1(new_new_n981_), .B0(new_new_n212_), .Y(new_new_n1130_));
  NA2        g1108(.A(new_new_n166_), .B(i_5_), .Y(new_new_n1131_));
  AOI210     g1109(.A0(new_new_n1130_), .A1(new_new_n836_), .B0(new_new_n1131_), .Y(new_new_n1132_));
  NO3        g1110(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n1133_));
  OAI210     g1111(.A0(new_new_n992_), .A1(new_new_n324_), .B0(new_new_n1133_), .Y(new_new_n1134_));
  NO2        g1112(.A(new_new_n1134_), .B(new_new_n794_), .Y(new_new_n1135_));
  NO4        g1113(.A(new_new_n1016_), .B(new_new_n517_), .C(new_new_n262_), .D(new_new_n261_), .Y(new_new_n1136_));
  NO2        g1114(.A(new_new_n1136_), .B(new_new_n618_), .Y(new_new_n1137_));
  NO2        g1115(.A(new_new_n877_), .B(new_new_n387_), .Y(new_new_n1138_));
  AOI210     g1116(.A0(new_new_n1138_), .A1(new_new_n1137_), .B0(new_new_n38_), .Y(new_new_n1139_));
  NO4        g1117(.A(new_new_n1139_), .B(new_new_n1135_), .C(new_new_n1132_), .D(new_new_n1128_), .Y(new_new_n1140_));
  OAI210     g1118(.A0(new_new_n1125_), .A1(i_4_), .B0(new_new_n1140_), .Y(new_new_n1141_));
  NO3        g1119(.A(new_new_n1141_), .B(new_new_n1115_), .C(new_new_n1113_), .Y(new_new_n1142_));
  NA4        g1120(.A(new_new_n1142_), .B(new_new_n1095_), .C(new_new_n1023_), .D(new_new_n936_), .Y(men4));
  INV        g1121(.A(i_5_), .Y(new_new_n1146_));
endmodule


