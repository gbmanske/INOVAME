//Benchmark atmr_max1024_476_0.5

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n393_, men_men_n394_, men_men_n395_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x8), .B(x3), .Y(ori_ori_n26_));
  NA2        o010(.A(x4), .B(x2), .Y(ori_ori_n27_));
  NO3        o011(.A(ori_ori_n27_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n28_));
  NO2        o012(.A(ori_ori_n28_), .B(ori_ori_n24_), .Y(ori_ori_n29_));
  NO2        o013(.A(x4), .B(x3), .Y(ori_ori_n30_));
  INV        o014(.A(ori_ori_n30_), .Y(ori_ori_n31_));
  NOi21      o015(.An(ori_ori_n23_), .B(ori_ori_n29_), .Y(ori00));
  NO2        o016(.A(x1), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x6), .Y(ori_ori_n34_));
  NA2        o018(.A(x4), .B(x3), .Y(ori_ori_n35_));
  NO2        o019(.A(ori_ori_n23_), .B(ori_ori_n35_), .Y(ori_ori_n36_));
  NO2        o020(.A(x2), .B(x0), .Y(ori_ori_n37_));
  INV        o021(.A(x3), .Y(ori_ori_n38_));
  NO2        o022(.A(ori_ori_n38_), .B(ori_ori_n18_), .Y(ori_ori_n39_));
  INV        o023(.A(ori_ori_n39_), .Y(ori_ori_n40_));
  INV        o024(.A(x4), .Y(ori_ori_n41_));
  OAI210     o025(.A0(ori_ori_n41_), .A1(ori_ori_n40_), .B0(ori_ori_n37_), .Y(ori_ori_n42_));
  INV        o026(.A(x4), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n44_));
  NA2        o028(.A(ori_ori_n44_), .B(x2), .Y(ori_ori_n45_));
  INV        o029(.A(ori_ori_n42_), .Y(ori_ori_n46_));
  NO2        o030(.A(ori_ori_n22_), .B(ori_ori_n33_), .Y(ori_ori_n47_));
  INV        o031(.A(x2), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n38_), .B(ori_ori_n18_), .Y(ori_ori_n50_));
  INV        o034(.A(ori_ori_n49_), .Y(ori_ori_n51_));
  OAI210     o035(.A0(ori_ori_n47_), .A1(ori_ori_n31_), .B0(ori_ori_n51_), .Y(ori_ori_n52_));
  NO3        o036(.A(ori_ori_n52_), .B(ori_ori_n46_), .C(ori_ori_n36_), .Y(ori01));
  NA2        o037(.A(ori_ori_n38_), .B(x1), .Y(ori_ori_n54_));
  INV        o038(.A(x9), .Y(ori_ori_n55_));
  NO2        o039(.A(ori_ori_n54_), .B(x5), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n25_), .B(ori_ori_n48_), .Y(ori_ori_n57_));
  NA2        o041(.A(ori_ori_n50_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  INV        o042(.A(ori_ori_n58_), .Y(ori_ori_n59_));
  NA2        o043(.A(ori_ori_n59_), .B(x4), .Y(ori_ori_n60_));
  INV        o044(.A(x0), .Y(ori_ori_n61_));
  NA2        o045(.A(x5), .B(x3), .Y(ori_ori_n62_));
  NO2        o046(.A(x8), .B(x6), .Y(ori_ori_n63_));
  NAi21      o047(.An(x4), .B(x3), .Y(ori_ori_n64_));
  INV        o048(.A(ori_ori_n64_), .Y(ori_ori_n65_));
  NO2        o049(.A(ori_ori_n65_), .B(ori_ori_n22_), .Y(ori_ori_n66_));
  NO2        o050(.A(x4), .B(x2), .Y(ori_ori_n67_));
  NO2        o051(.A(ori_ori_n66_), .B(ori_ori_n18_), .Y(ori_ori_n68_));
  NO2        o052(.A(ori_ori_n68_), .B(ori_ori_n61_), .Y(ori_ori_n69_));
  NA2        o053(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n70_));
  INV        o054(.A(x8), .Y(ori_ori_n71_));
  AOI210     o055(.A0(ori_ori_n50_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n40_), .B(ori_ori_n43_), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n74_));
  NA2        o058(.A(x4), .B(ori_ori_n38_), .Y(ori_ori_n75_));
  NO2        o059(.A(ori_ori_n75_), .B(x1), .Y(ori_ori_n76_));
  NA2        o060(.A(ori_ori_n48_), .B(x1), .Y(ori_ori_n77_));
  OAI210     o061(.A0(ori_ori_n77_), .A1(ori_ori_n35_), .B0(ori_ori_n17_), .Y(ori_ori_n78_));
  NO3        o062(.A(ori_ori_n78_), .B(ori_ori_n76_), .C(ori_ori_n74_), .Y(ori_ori_n79_));
  AO210      o063(.A0(ori_ori_n69_), .A1(ori_ori_n60_), .B0(ori_ori_n79_), .Y(ori02));
  NO2        o064(.A(x3), .B(ori_ori_n48_), .Y(ori_ori_n81_));
  NO2        o065(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n82_));
  NA2        o066(.A(ori_ori_n38_), .B(x0), .Y(ori_ori_n83_));
  INV        o067(.A(ori_ori_n83_), .Y(ori_ori_n84_));
  AOI220     o068(.A0(ori_ori_n84_), .A1(ori_ori_n82_), .B0(ori_ori_n81_), .B1(x4), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n85_), .B(x7), .Y(ori_ori_n86_));
  OR2        o070(.A(x8), .B(x0), .Y(ori_ori_n87_));
  INV        o071(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  NAi21      o072(.An(x2), .B(x8), .Y(ori_ori_n89_));
  NO2        o073(.A(x4), .B(x1), .Y(ori_ori_n90_));
  NA2        o074(.A(ori_ori_n90_), .B(x2), .Y(ori_ori_n91_));
  NO2        o075(.A(ori_ori_n91_), .B(ori_ori_n62_), .Y(ori_ori_n92_));
  NO2        o076(.A(x5), .B(ori_ori_n43_), .Y(ori_ori_n93_));
  NO2        o077(.A(x7), .B(x0), .Y(ori_ori_n94_));
  NO2        o078(.A(ori_ori_n21_), .B(ori_ori_n38_), .Y(ori_ori_n95_));
  NA2        o079(.A(x5), .B(x0), .Y(ori_ori_n96_));
  NO2        o080(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n97_));
  NA3        o081(.A(ori_ori_n97_), .B(ori_ori_n96_), .C(ori_ori_n95_), .Y(ori_ori_n98_));
  NA2        o082(.A(ori_ori_n98_), .B(ori_ori_n34_), .Y(ori_ori_n99_));
  NO3        o083(.A(ori_ori_n99_), .B(ori_ori_n92_), .C(ori_ori_n86_), .Y(ori_ori_n100_));
  NO3        o084(.A(ori_ori_n62_), .B(x4), .C(ori_ori_n24_), .Y(ori_ori_n101_));
  NA2        o085(.A(x7), .B(x3), .Y(ori_ori_n102_));
  NO2        o086(.A(ori_ori_n75_), .B(x5), .Y(ori_ori_n103_));
  NO2        o087(.A(x9), .B(x7), .Y(ori_ori_n104_));
  NOi21      o088(.An(x8), .B(x0), .Y(ori_ori_n105_));
  OA210      o089(.A0(ori_ori_n104_), .A1(x1), .B0(ori_ori_n105_), .Y(ori_ori_n106_));
  INV        o090(.A(x7), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n106_), .B(ori_ori_n103_), .Y(ori_ori_n109_));
  OAI210     o093(.A0(ori_ori_n102_), .A1(ori_ori_n45_), .B0(ori_ori_n109_), .Y(ori_ori_n110_));
  NA2        o094(.A(x5), .B(x1), .Y(ori_ori_n111_));
  INV        o095(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  AOI210     o096(.A0(ori_ori_n112_), .A1(x0), .B0(ori_ori_n34_), .Y(ori_ori_n113_));
  INV        o097(.A(x2), .Y(ori_ori_n114_));
  NA2        o098(.A(ori_ori_n114_), .B(ori_ori_n56_), .Y(ori_ori_n115_));
  NA2        o099(.A(ori_ori_n115_), .B(ori_ori_n113_), .Y(ori_ori_n116_));
  NO3        o100(.A(ori_ori_n116_), .B(ori_ori_n110_), .C(ori_ori_n101_), .Y(ori_ori_n117_));
  NO2        o101(.A(ori_ori_n117_), .B(ori_ori_n100_), .Y(ori_ori_n118_));
  NA2        o102(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n119_));
  NA2        o103(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n120_));
  NA2        o104(.A(x8), .B(x0), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n107_), .B(ori_ori_n25_), .Y(ori_ori_n122_));
  NA2        o106(.A(x2), .B(x0), .Y(ori_ori_n123_));
  NA2        o107(.A(x4), .B(x1), .Y(ori_ori_n124_));
  NAi21      o108(.An(ori_ori_n90_), .B(ori_ori_n124_), .Y(ori_ori_n125_));
  NOi21      o109(.An(ori_ori_n125_), .B(ori_ori_n123_), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n304_), .B(ori_ori_n38_), .Y(ori_ori_n127_));
  INV        o111(.A(ori_ori_n93_), .Y(ori_ori_n128_));
  NA2        o112(.A(ori_ori_n33_), .B(ori_ori_n71_), .Y(ori_ori_n129_));
  NO3        o113(.A(ori_ori_n129_), .B(ori_ori_n128_), .C(x7), .Y(ori_ori_n130_));
  NA2        o114(.A(ori_ori_n125_), .B(ori_ori_n37_), .Y(ori_ori_n131_));
  INV        o115(.A(ori_ori_n131_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n132_), .B(ori_ori_n130_), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n133_), .B(x3), .Y(ori_ori_n134_));
  NO3        o118(.A(ori_ori_n134_), .B(ori_ori_n127_), .C(ori_ori_n118_), .Y(ori03));
  NO2        o119(.A(ori_ori_n43_), .B(x3), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n137_));
  NO2        o121(.A(x5), .B(x4), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n139_));
  AN2        o123(.A(ori_ori_n137_), .B(ori_ori_n49_), .Y(ori_ori_n140_));
  INV        o124(.A(ori_ori_n140_), .Y(ori_ori_n141_));
  NA2        o125(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n142_));
  NA2        o126(.A(x9), .B(ori_ori_n48_), .Y(ori_ori_n143_));
  NO2        o127(.A(x5), .B(x1), .Y(ori_ori_n144_));
  NO2        o128(.A(ori_ori_n142_), .B(ori_ori_n119_), .Y(ori_ori_n145_));
  NO3        o129(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n146_));
  NA2        o130(.A(ori_ori_n146_), .B(ori_ori_n43_), .Y(ori_ori_n147_));
  NA2        o131(.A(ori_ori_n147_), .B(ori_ori_n141_), .Y(ori_ori_n148_));
  NO2        o132(.A(ori_ori_n43_), .B(ori_ori_n38_), .Y(ori_ori_n149_));
  NO2        o133(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n150_), .B(x6), .Y(ori_ori_n151_));
  NOi21      o135(.An(ori_ori_n67_), .B(ori_ori_n151_), .Y(ori_ori_n152_));
  NO2        o136(.A(ori_ori_n152_), .B(ori_ori_n107_), .Y(ori_ori_n153_));
  OR2        o137(.A(ori_ori_n153_), .B(ori_ori_n122_), .Y(ori_ori_n154_));
  NA2        o138(.A(ori_ori_n38_), .B(ori_ori_n48_), .Y(ori_ori_n155_));
  OAI210     o139(.A0(ori_ori_n155_), .A1(ori_ori_n25_), .B0(ori_ori_n120_), .Y(ori_ori_n156_));
  NO2        o140(.A(ori_ori_n124_), .B(x6), .Y(ori_ori_n157_));
  NA2        o141(.A(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  NA2        o142(.A(x6), .B(ori_ori_n43_), .Y(ori_ori_n159_));
  OAI210     o143(.A0(ori_ori_n88_), .A1(ori_ori_n63_), .B0(x4), .Y(ori_ori_n160_));
  AOI210     o144(.A0(ori_ori_n160_), .A1(ori_ori_n159_), .B0(ori_ori_n62_), .Y(ori_ori_n161_));
  NA3        o145(.A(ori_ori_n142_), .B(ori_ori_n93_), .C(x6), .Y(ori_ori_n162_));
  INV        o146(.A(ori_ori_n56_), .Y(ori_ori_n163_));
  NA2        o147(.A(ori_ori_n163_), .B(ori_ori_n162_), .Y(ori_ori_n164_));
  OAI210     o148(.A0(ori_ori_n164_), .A1(ori_ori_n161_), .B0(x2), .Y(ori_ori_n165_));
  NA3        o149(.A(ori_ori_n165_), .B(ori_ori_n158_), .C(ori_ori_n154_), .Y(ori_ori_n166_));
  AOI210     o150(.A0(ori_ori_n148_), .A1(x8), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  NO2        o151(.A(ori_ori_n71_), .B(x3), .Y(ori_ori_n168_));
  NA2        o152(.A(ori_ori_n168_), .B(ori_ori_n138_), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n70_), .B(ori_ori_n25_), .Y(ori_ori_n170_));
  AOI210     o154(.A0(ori_ori_n151_), .A1(ori_ori_n108_), .B0(ori_ori_n170_), .Y(ori_ori_n171_));
  AOI210     o155(.A0(ori_ori_n171_), .A1(ori_ori_n169_), .B0(x2), .Y(ori_ori_n172_));
  NA2        o156(.A(ori_ori_n55_), .B(x6), .Y(ori_ori_n173_));
  NA2        o157(.A(ori_ori_n38_), .B(ori_ori_n17_), .Y(ori_ori_n174_));
  AOI210     o158(.A0(x3), .A1(x2), .B0(ori_ori_n43_), .Y(ori_ori_n175_));
  OAI210     o159(.A0(ori_ori_n96_), .A1(x3), .B0(ori_ori_n175_), .Y(ori_ori_n176_));
  NA2        o160(.A(ori_ori_n176_), .B(x1), .Y(ori_ori_n177_));
  INV        o161(.A(ori_ori_n177_), .Y(ori_ori_n178_));
  NA2        o162(.A(x6), .B(x2), .Y(ori_ori_n179_));
  NA2        o163(.A(x4), .B(ori_ori_n178_), .Y(ori_ori_n180_));
  NA2        o164(.A(x9), .B(ori_ori_n38_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n181_), .B(x5), .Y(ori_ori_n182_));
  OR3        o166(.A(ori_ori_n182_), .B(ori_ori_n137_), .C(ori_ori_n103_), .Y(ori_ori_n183_));
  NA2        o167(.A(ori_ori_n183_), .B(ori_ori_n37_), .Y(ori_ori_n184_));
  AOI210     o168(.A0(ori_ori_n184_), .A1(ori_ori_n180_), .B0(x8), .Y(ori_ori_n185_));
  NA2        o169(.A(ori_ori_n144_), .B(ori_ori_n55_), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n186_), .B(ori_ori_n155_), .Y(ori_ori_n187_));
  NO4        o171(.A(ori_ori_n187_), .B(ori_ori_n185_), .C(x7), .D(ori_ori_n172_), .Y(ori_ori_n188_));
  OAI210     o172(.A0(x8), .A1(x6), .B0(ori_ori_n39_), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n189_), .B(ori_ori_n128_), .Y(ori_ori_n190_));
  NOi21      o174(.An(ori_ori_n179_), .B(ori_ori_n17_), .Y(ori_ori_n191_));
  NA3        o175(.A(ori_ori_n191_), .B(ori_ori_n144_), .C(ori_ori_n35_), .Y(ori_ori_n192_));
  AOI210     o176(.A0(ori_ori_n34_), .A1(ori_ori_n48_), .B0(x0), .Y(ori_ori_n193_));
  NA3        o177(.A(ori_ori_n193_), .B(ori_ori_n112_), .C(ori_ori_n31_), .Y(ori_ori_n194_));
  NA2        o178(.A(x3), .B(x2), .Y(ori_ori_n195_));
  AOI220     o179(.A0(ori_ori_n195_), .A1(ori_ori_n155_), .B0(ori_ori_n194_), .B1(ori_ori_n192_), .Y(ori_ori_n196_));
  NAi21      o180(.An(x4), .B(x0), .Y(ori_ori_n197_));
  NO3        o181(.A(ori_ori_n197_), .B(ori_ori_n39_), .C(x2), .Y(ori_ori_n198_));
  OAI210     o182(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n198_), .Y(ori_ori_n199_));
  NO2        o183(.A(ori_ori_n193_), .B(ori_ori_n191_), .Y(ori_ori_n200_));
  AOI220     o184(.A0(ori_ori_n200_), .A1(ori_ori_n65_), .B0(ori_ori_n18_), .B1(ori_ori_n30_), .Y(ori_ori_n201_));
  AOI210     o185(.A0(ori_ori_n201_), .A1(ori_ori_n199_), .B0(ori_ori_n25_), .Y(ori_ori_n202_));
  NA3        o186(.A(ori_ori_n34_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n193_), .B(ori_ori_n191_), .Y(ori_ori_n204_));
  INV        o188(.A(ori_ori_n145_), .Y(ori_ori_n205_));
  NA2        o189(.A(ori_ori_n34_), .B(ori_ori_n38_), .Y(ori_ori_n206_));
  NO2        o190(.A(ori_ori_n159_), .B(ori_ori_n205_), .Y(ori_ori_n207_));
  AO210      o191(.A0(ori_ori_n204_), .A1(ori_ori_n103_), .B0(ori_ori_n207_), .Y(ori_ori_n208_));
  NO4        o192(.A(ori_ori_n208_), .B(ori_ori_n202_), .C(ori_ori_n196_), .D(ori_ori_n190_), .Y(ori_ori_n209_));
  OAI210     o193(.A0(ori_ori_n188_), .A1(ori_ori_n167_), .B0(ori_ori_n209_), .Y(ori04));
  NO2        o194(.A(x2), .B(x1), .Y(ori_ori_n211_));
  OAI210     o195(.A0(ori_ori_n174_), .A1(ori_ori_n211_), .B0(ori_ori_n34_), .Y(ori_ori_n212_));
  NO2        o196(.A(ori_ori_n195_), .B(ori_ori_n139_), .Y(ori_ori_n213_));
  INV        o197(.A(ori_ori_n213_), .Y(ori_ori_n214_));
  NA2        o198(.A(ori_ori_n214_), .B(x6), .Y(ori_ori_n215_));
  NA2        o199(.A(ori_ori_n215_), .B(ori_ori_n212_), .Y(ori_ori_n216_));
  NO2        o200(.A(ori_ori_n143_), .B(ori_ori_n83_), .Y(ori_ori_n217_));
  NO3        o201(.A(ori_ori_n173_), .B(ori_ori_n89_), .C(ori_ori_n18_), .Y(ori_ori_n218_));
  NO2        o202(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  OAI210     o203(.A0(ori_ori_n87_), .A1(ori_ori_n77_), .B0(ori_ori_n121_), .Y(ori_ori_n220_));
  NA3        o204(.A(ori_ori_n220_), .B(x6), .C(x3), .Y(ori_ori_n221_));
  AOI210     o205(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n222_));
  OAI220     o206(.A0(ori_ori_n222_), .A1(ori_ori_n206_), .B0(ori_ori_n301_), .B1(ori_ori_n203_), .Y(ori_ori_n223_));
  INV        o207(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NA2        o208(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n225_));
  OAI210     o209(.A0(ori_ori_n77_), .A1(ori_ori_n17_), .B0(ori_ori_n225_), .Y(ori_ori_n226_));
  NA2        o210(.A(ori_ori_n226_), .B(ori_ori_n63_), .Y(ori_ori_n227_));
  NA4        o211(.A(ori_ori_n227_), .B(ori_ori_n224_), .C(ori_ori_n221_), .D(ori_ori_n219_), .Y(ori_ori_n228_));
  OAI210     o212(.A0(ori_ori_n82_), .A1(x3), .B0(ori_ori_n198_), .Y(ori_ori_n229_));
  NA2        o213(.A(ori_ori_n302_), .B(ori_ori_n67_), .Y(ori_ori_n230_));
  NA3        o214(.A(ori_ori_n230_), .B(ori_ori_n229_), .C(ori_ori_n107_), .Y(ori_ori_n231_));
  AOI210     o215(.A0(ori_ori_n228_), .A1(x4), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  INV        o216(.A(x1), .Y(ori_ori_n233_));
  XO2        o217(.A(x4), .B(x0), .Y(ori_ori_n234_));
  INV        o218(.A(x4), .Y(ori_ori_n235_));
  AOI210     o219(.A0(ori_ori_n235_), .A1(ori_ori_n233_), .B0(x3), .Y(ori_ori_n236_));
  NA2        o220(.A(ori_ori_n18_), .B(x6), .Y(ori_ori_n237_));
  NO2        o221(.A(ori_ori_n105_), .B(ori_ori_n64_), .Y(ori_ori_n238_));
  NOi21      o222(.An(ori_ori_n90_), .B(ori_ori_n26_), .Y(ori_ori_n239_));
  AOI210     o223(.A0(ori_ori_n303_), .A1(ori_ori_n238_), .B0(ori_ori_n239_), .Y(ori_ori_n240_));
  OAI210     o224(.A0(ori_ori_n197_), .A1(ori_ori_n55_), .B0(ori_ori_n240_), .Y(ori_ori_n241_));
  OAI220     o225(.A0(ori_ori_n241_), .A1(x6), .B0(ori_ori_n237_), .B1(ori_ori_n236_), .Y(ori_ori_n242_));
  AO220      o226(.A0(x7), .A1(ori_ori_n242_), .B0(ori_ori_n232_), .B1(ori_ori_n216_), .Y(ori_ori_n243_));
  AOI220     o227(.A0(ori_ori_n67_), .A1(ori_ori_n33_), .B0(ori_ori_n146_), .B1(ori_ori_n44_), .Y(ori_ori_n244_));
  NA2        o228(.A(ori_ori_n244_), .B(ori_ori_n243_), .Y(ori_ori_n245_));
  INV        o229(.A(ori_ori_n82_), .Y(ori_ori_n246_));
  NA2        o230(.A(ori_ori_n246_), .B(ori_ori_n225_), .Y(ori_ori_n247_));
  NA3        o231(.A(ori_ori_n247_), .B(ori_ori_n136_), .C(ori_ori_n107_), .Y(ori_ori_n248_));
  OAI210     o232(.A0(ori_ori_n27_), .A1(x1), .B0(ori_ori_n155_), .Y(ori_ori_n249_));
  AO220      o233(.A0(ori_ori_n249_), .A1(ori_ori_n104_), .B0(ori_ori_n81_), .B1(x4), .Y(ori_ori_n250_));
  NA3        o234(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n251_));
  NA2        o235(.A(ori_ori_n149_), .B(x0), .Y(ori_ori_n252_));
  OAI220     o236(.A0(ori_ori_n252_), .A1(ori_ori_n143_), .B0(ori_ori_n251_), .B1(x2), .Y(ori_ori_n253_));
  AOI210     o237(.A0(ori_ori_n250_), .A1(ori_ori_n88_), .B0(ori_ori_n253_), .Y(ori_ori_n254_));
  AOI210     o238(.A0(ori_ori_n254_), .A1(ori_ori_n248_), .B0(ori_ori_n25_), .Y(ori_ori_n255_));
  NA3        o239(.A(x8), .B(ori_ori_n149_), .C(x0), .Y(ori_ori_n256_));
  NAi21      o240(.An(ori_ori_n45_), .B(ori_ori_n122_), .Y(ori_ori_n257_));
  NA2        o241(.A(ori_ori_n257_), .B(ori_ori_n256_), .Y(ori_ori_n258_));
  OAI210     o242(.A0(ori_ori_n258_), .A1(ori_ori_n255_), .B0(x6), .Y(ori_ori_n259_));
  NA2        o243(.A(x7), .B(ori_ori_n149_), .Y(ori_ori_n260_));
  INV        o244(.A(x1), .Y(ori_ori_n261_));
  OAI210     o245(.A0(ori_ori_n260_), .A1(x8), .B0(ori_ori_n261_), .Y(ori_ori_n262_));
  NAi31      o246(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n263_));
  NA3        o247(.A(x0), .B(ori_ori_n102_), .C(x9), .Y(ori_ori_n264_));
  NO2        o248(.A(ori_ori_n107_), .B(x0), .Y(ori_ori_n265_));
  AOI210     o249(.A0(ori_ori_n238_), .A1(ori_ori_n107_), .B0(ori_ori_n168_), .Y(ori_ori_n266_));
  NA4        o250(.A(ori_ori_n266_), .B(x1), .C(ori_ori_n264_), .D(ori_ori_n45_), .Y(ori_ori_n267_));
  NA2        o251(.A(ori_ori_n262_), .B(ori_ori_n267_), .Y(ori_ori_n268_));
  NOi31      o252(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n269_));
  NO3        o253(.A(ori_ori_n269_), .B(x0), .C(x2), .Y(ori_ori_n270_));
  OAI210     o254(.A0(ori_ori_n197_), .A1(ori_ori_n38_), .B0(ori_ori_n234_), .Y(ori_ori_n271_));
  INV        o255(.A(ori_ori_n251_), .Y(ori_ori_n272_));
  AOI220     o256(.A0(ori_ori_n272_), .A1(ori_ori_n71_), .B0(ori_ori_n271_), .B1(ori_ori_n107_), .Y(ori_ori_n273_));
  NO2        o257(.A(ori_ori_n273_), .B(ori_ori_n48_), .Y(ori_ori_n274_));
  NO2        o258(.A(ori_ori_n274_), .B(ori_ori_n270_), .Y(ori_ori_n275_));
  AOI210     o259(.A0(ori_ori_n275_), .A1(ori_ori_n268_), .B0(ori_ori_n25_), .Y(ori_ori_n276_));
  NA4        o260(.A(ori_ori_n30_), .B(ori_ori_n71_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n277_));
  NA2        o261(.A(x1), .B(ori_ori_n175_), .Y(ori_ori_n278_));
  INV        o262(.A(ori_ori_n278_), .Y(ori_ori_n279_));
  NO2        o263(.A(ori_ori_n121_), .B(ori_ori_n35_), .Y(ori_ori_n280_));
  OAI210     o264(.A0(ori_ori_n280_), .A1(ori_ori_n279_), .B0(x7), .Y(ori_ori_n281_));
  NA2        o265(.A(ori_ori_n281_), .B(ori_ori_n277_), .Y(ori_ori_n282_));
  OAI210     o266(.A0(ori_ori_n282_), .A1(ori_ori_n276_), .B0(ori_ori_n34_), .Y(ori_ori_n283_));
  INV        o267(.A(ori_ori_n265_), .Y(ori_ori_n284_));
  NO3        o268(.A(ori_ori_n284_), .B(ori_ori_n62_), .C(x4), .Y(ori_ori_n285_));
  NA2        o269(.A(ori_ori_n174_), .B(ori_ori_n21_), .Y(ori_ori_n286_));
  NO2        o270(.A(ori_ori_n111_), .B(ori_ori_n94_), .Y(ori_ori_n287_));
  NA2        o271(.A(ori_ori_n287_), .B(ori_ori_n286_), .Y(ori_ori_n288_));
  NO2        o272(.A(ori_ori_n288_), .B(ori_ori_n27_), .Y(ori_ori_n289_));
  INV        o273(.A(ori_ori_n263_), .Y(ori_ori_n290_));
  NA2        o274(.A(ori_ori_n290_), .B(ori_ori_n122_), .Y(ori_ori_n291_));
  OAI220     o275(.A0(ori_ori_n181_), .A1(x2), .B0(ori_ori_n111_), .B1(ori_ori_n38_), .Y(ori_ori_n292_));
  NO3        o276(.A(ori_ori_n269_), .B(x3), .C(ori_ori_n48_), .Y(ori_ori_n293_));
  AOI220     o277(.A0(ori_ori_n293_), .A1(x0), .B0(ori_ori_n292_), .B1(ori_ori_n94_), .Y(ori_ori_n294_));
  AOI210     o278(.A0(ori_ori_n294_), .A1(ori_ori_n291_), .B0(ori_ori_n159_), .Y(ori_ori_n295_));
  NO3        o279(.A(ori_ori_n295_), .B(ori_ori_n289_), .C(ori_ori_n285_), .Y(ori_ori_n296_));
  NA3        o280(.A(ori_ori_n296_), .B(ori_ori_n283_), .C(ori_ori_n259_), .Y(ori_ori_n297_));
  AOI210     o281(.A0(ori_ori_n245_), .A1(ori_ori_n25_), .B0(ori_ori_n297_), .Y(ori05));
  INV        o282(.A(x2), .Y(ori_ori_n301_));
  INV        o283(.A(x6), .Y(ori_ori_n302_));
  INV        o284(.A(x2), .Y(ori_ori_n303_));
  INV        o285(.A(ori_ori_n126_), .Y(ori_ori_n304_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  INV        m005(.A(mai_mai_n19_), .Y(mai_mai_n22_));
  NA2        m006(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n23_));
  INV        m007(.A(x5), .Y(mai_mai_n24_));
  NA2        m008(.A(x8), .B(x3), .Y(mai_mai_n25_));
  NA2        m009(.A(x4), .B(x2), .Y(mai_mai_n26_));
  INV        m010(.A(mai_mai_n23_), .Y(mai_mai_n27_));
  NO2        m011(.A(x4), .B(x3), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  NOi21      m013(.An(mai_mai_n22_), .B(mai_mai_n27_), .Y(mai00));
  NO2        m014(.A(x1), .B(x0), .Y(mai_mai_n31_));
  INV        m015(.A(x6), .Y(mai_mai_n32_));
  NO2        m016(.A(mai_mai_n32_), .B(mai_mai_n24_), .Y(mai_mai_n33_));
  AN2        m017(.A(x8), .B(x7), .Y(mai_mai_n34_));
  NA3        m018(.A(mai_mai_n34_), .B(mai_mai_n33_), .C(mai_mai_n31_), .Y(mai_mai_n35_));
  NA2        m019(.A(x4), .B(x3), .Y(mai_mai_n36_));
  AOI210     m020(.A0(mai_mai_n35_), .A1(mai_mai_n22_), .B0(mai_mai_n36_), .Y(mai_mai_n37_));
  NO2        m021(.A(x2), .B(x0), .Y(mai_mai_n38_));
  INV        m022(.A(x3), .Y(mai_mai_n39_));
  NO2        m023(.A(mai_mai_n39_), .B(mai_mai_n18_), .Y(mai_mai_n40_));
  INV        m024(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(mai_mai_n33_), .B(x4), .Y(mai_mai_n42_));
  OAI210     m026(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n38_), .Y(mai_mai_n43_));
  INV        m027(.A(x4), .Y(mai_mai_n44_));
  NO2        m028(.A(mai_mai_n44_), .B(mai_mai_n17_), .Y(mai_mai_n45_));
  NA2        m029(.A(mai_mai_n45_), .B(x2), .Y(mai_mai_n46_));
  INV        m030(.A(mai_mai_n43_), .Y(mai_mai_n47_));
  NA2        m031(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n48_));
  NA2        m032(.A(mai_mai_n48_), .B(mai_mai_n31_), .Y(mai_mai_n49_));
  INV        m033(.A(x2), .Y(mai_mai_n50_));
  NO2        m034(.A(mai_mai_n50_), .B(mai_mai_n17_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n39_), .B(mai_mai_n18_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  OAI210     m037(.A0(mai_mai_n49_), .A1(mai_mai_n29_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  NO3        m038(.A(mai_mai_n54_), .B(mai_mai_n47_), .C(mai_mai_n37_), .Y(mai01));
  NA2        m039(.A(x8), .B(x7), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n39_), .B(x1), .Y(mai_mai_n57_));
  INV        m041(.A(x9), .Y(mai_mai_n58_));
  NO2        m042(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NO2        m043(.A(x7), .B(x6), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n57_), .B(x5), .Y(mai_mai_n61_));
  NO2        m045(.A(x8), .B(x2), .Y(mai_mai_n62_));
  INV        m046(.A(mai_mai_n62_), .Y(mai_mai_n63_));
  NO2        m047(.A(mai_mai_n63_), .B(x1), .Y(mai_mai_n64_));
  OA210      m048(.A0(mai_mai_n64_), .A1(mai_mai_n61_), .B0(mai_mai_n60_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n40_), .A1(mai_mai_n24_), .B0(mai_mai_n50_), .Y(mai_mai_n66_));
  OAI210     m050(.A0(mai_mai_n52_), .A1(mai_mai_n20_), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  NAi31      m051(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n67_), .B(mai_mai_n65_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n69_), .A1(mai_mai_n59_), .B0(x4), .Y(mai_mai_n70_));
  NA2        m054(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n71_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n72_));
  NA2        m056(.A(x5), .B(x3), .Y(mai_mai_n73_));
  NO3        m057(.A(mai_mai_n73_), .B(mai_mai_n60_), .C(mai_mai_n50_), .Y(mai_mai_n74_));
  NAi21      m058(.An(x4), .B(x3), .Y(mai_mai_n75_));
  INV        m059(.A(mai_mai_n75_), .Y(mai_mai_n76_));
  NO2        m060(.A(x4), .B(x2), .Y(mai_mai_n77_));
  NO2        m061(.A(mai_mai_n77_), .B(x3), .Y(mai_mai_n78_));
  NO2        m062(.A(mai_mai_n74_), .B(mai_mai_n72_), .Y(mai_mai_n79_));
  NO3        m063(.A(x6), .B(mai_mai_n39_), .C(x1), .Y(mai_mai_n80_));
  INV        m064(.A(x4), .Y(mai_mai_n81_));
  NA2        m065(.A(mai_mai_n80_), .B(mai_mai_n81_), .Y(mai_mai_n82_));
  NA2        m066(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n83_));
  NO2        m067(.A(mai_mai_n83_), .B(mai_mai_n24_), .Y(mai_mai_n84_));
  INV        m068(.A(x8), .Y(mai_mai_n85_));
  NA2        m069(.A(x2), .B(x1), .Y(mai_mai_n86_));
  NO2        m070(.A(mai_mai_n86_), .B(mai_mai_n85_), .Y(mai_mai_n87_));
  NO2        m071(.A(mai_mai_n87_), .B(mai_mai_n84_), .Y(mai_mai_n88_));
  INV        m072(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  AOI210     m073(.A0(mai_mai_n52_), .A1(mai_mai_n24_), .B0(mai_mai_n50_), .Y(mai_mai_n90_));
  OAI210     m074(.A0(mai_mai_n41_), .A1(mai_mai_n33_), .B0(mai_mai_n44_), .Y(mai_mai_n91_));
  NO3        m075(.A(mai_mai_n91_), .B(mai_mai_n90_), .C(mai_mai_n89_), .Y(mai_mai_n92_));
  NA2        m076(.A(x4), .B(mai_mai_n39_), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n44_), .B(mai_mai_n50_), .Y(mai_mai_n94_));
  OAI210     m078(.A0(mai_mai_n94_), .A1(mai_mai_n39_), .B0(mai_mai_n18_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n48_), .B(mai_mai_n95_), .Y(mai_mai_n96_));
  NO2        m080(.A(x3), .B(x2), .Y(mai_mai_n97_));
  NA2        m081(.A(mai_mai_n50_), .B(x1), .Y(mai_mai_n98_));
  OAI210     m082(.A0(mai_mai_n98_), .A1(mai_mai_n36_), .B0(mai_mai_n17_), .Y(mai_mai_n99_));
  NO4        m083(.A(mai_mai_n99_), .B(mai_mai_n97_), .C(mai_mai_n96_), .D(mai_mai_n92_), .Y(mai_mai_n100_));
  AO220      m084(.A0(mai_mai_n100_), .A1(mai_mai_n82_), .B0(mai_mai_n79_), .B1(mai_mai_n70_), .Y(mai02));
  NO2        m085(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n102_));
  NO2        m086(.A(x4), .B(x2), .Y(mai_mai_n103_));
  NO3        m087(.A(mai_mai_n387_), .B(x7), .C(x5), .Y(mai_mai_n104_));
  NA2        m088(.A(x9), .B(x2), .Y(mai_mai_n105_));
  OR2        m089(.A(x8), .B(x0), .Y(mai_mai_n106_));
  NAi21      m090(.An(x2), .B(x8), .Y(mai_mai_n107_));
  NO2        m091(.A(x4), .B(x1), .Y(mai_mai_n108_));
  NA3        m092(.A(mai_mai_n108_), .B(mai_mai_n380_), .C(mai_mai_n56_), .Y(mai_mai_n109_));
  NOi21      m093(.An(x0), .B(x1), .Y(mai_mai_n110_));
  NO3        m094(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n111_));
  NOi21      m095(.An(x0), .B(x4), .Y(mai_mai_n112_));
  NO2        m096(.A(x8), .B(mai_mai_n58_), .Y(mai_mai_n113_));
  AOI220     m097(.A0(mai_mai_n113_), .A1(mai_mai_n112_), .B0(mai_mai_n111_), .B1(mai_mai_n110_), .Y(mai_mai_n114_));
  AOI210     m098(.A0(mai_mai_n114_), .A1(mai_mai_n109_), .B0(mai_mai_n73_), .Y(mai_mai_n115_));
  NO2        m099(.A(x5), .B(mai_mai_n44_), .Y(mai_mai_n116_));
  NA2        m100(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n117_));
  OAI210     m101(.A0(x0), .A1(mai_mai_n31_), .B0(mai_mai_n116_), .Y(mai_mai_n118_));
  NAi21      m102(.An(x0), .B(x4), .Y(mai_mai_n119_));
  NO2        m103(.A(mai_mai_n119_), .B(x1), .Y(mai_mai_n120_));
  NO2        m104(.A(x7), .B(x0), .Y(mai_mai_n121_));
  NO2        m105(.A(mai_mai_n77_), .B(mai_mai_n94_), .Y(mai_mai_n122_));
  NO2        m106(.A(mai_mai_n122_), .B(x3), .Y(mai_mai_n123_));
  OAI210     m107(.A0(mai_mai_n121_), .A1(mai_mai_n120_), .B0(mai_mai_n123_), .Y(mai_mai_n124_));
  NA2        m108(.A(x5), .B(x0), .Y(mai_mai_n125_));
  NO2        m109(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n126_));
  NA3        m110(.A(mai_mai_n124_), .B(mai_mai_n118_), .C(mai_mai_n32_), .Y(mai_mai_n127_));
  NO3        m111(.A(mai_mai_n127_), .B(mai_mai_n115_), .C(mai_mai_n104_), .Y(mai_mai_n128_));
  NO3        m112(.A(mai_mai_n73_), .B(mai_mai_n71_), .C(mai_mai_n23_), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n26_), .B(mai_mai_n24_), .Y(mai_mai_n130_));
  AOI220     m114(.A0(mai_mai_n110_), .A1(mai_mai_n130_), .B0(mai_mai_n61_), .B1(mai_mai_n17_), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n131_), .B(mai_mai_n56_), .Y(mai_mai_n132_));
  NO2        m116(.A(mai_mai_n93_), .B(x5), .Y(mai_mai_n133_));
  NO2        m117(.A(x9), .B(x7), .Y(mai_mai_n134_));
  NOi21      m118(.An(x8), .B(x0), .Y(mai_mai_n135_));
  NO2        m119(.A(mai_mai_n39_), .B(x2), .Y(mai_mai_n136_));
  INV        m120(.A(x7), .Y(mai_mai_n137_));
  NA2        m121(.A(mai_mai_n137_), .B(mai_mai_n18_), .Y(mai_mai_n138_));
  AOI220     m122(.A0(mai_mai_n138_), .A1(mai_mai_n136_), .B0(mai_mai_n102_), .B1(mai_mai_n34_), .Y(mai_mai_n139_));
  NO2        m123(.A(x4), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  NA2        m124(.A(x5), .B(x1), .Y(mai_mai_n141_));
  INV        m125(.A(mai_mai_n141_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n58_), .B(mai_mai_n85_), .Y(mai_mai_n143_));
  NAi31      m127(.An(mai_mai_n73_), .B(mai_mai_n34_), .C(mai_mai_n31_), .Y(mai_mai_n144_));
  NA2        m128(.A(mai_mai_n144_), .B(x6), .Y(mai_mai_n145_));
  NO4        m129(.A(mai_mai_n145_), .B(mai_mai_n140_), .C(mai_mai_n132_), .D(mai_mai_n129_), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n146_), .B(mai_mai_n128_), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n125_), .B(mai_mai_n122_), .Y(mai_mai_n148_));
  NA2        m132(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n149_));
  NA2        m133(.A(mai_mai_n24_), .B(mai_mai_n17_), .Y(mai_mai_n150_));
  NA3        m134(.A(mai_mai_n150_), .B(mai_mai_n149_), .C(mai_mai_n23_), .Y(mai_mai_n151_));
  AN2        m135(.A(mai_mai_n151_), .B(mai_mai_n126_), .Y(mai_mai_n152_));
  NA2        m136(.A(x8), .B(x0), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n137_), .B(mai_mai_n24_), .Y(mai_mai_n154_));
  NO2        m138(.A(mai_mai_n110_), .B(x4), .Y(mai_mai_n155_));
  NA2        m139(.A(mai_mai_n155_), .B(mai_mai_n154_), .Y(mai_mai_n156_));
  AOI210     m140(.A0(mai_mai_n153_), .A1(mai_mai_n117_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NA2        m141(.A(x2), .B(x0), .Y(mai_mai_n158_));
  NA2        m142(.A(x4), .B(x1), .Y(mai_mai_n159_));
  NO2        m143(.A(x5), .B(mai_mai_n158_), .Y(mai_mai_n160_));
  NO4        m144(.A(mai_mai_n160_), .B(mai_mai_n157_), .C(mai_mai_n152_), .D(mai_mai_n148_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n161_), .B(mai_mai_n39_), .Y(mai_mai_n162_));
  NO2        m146(.A(mai_mai_n151_), .B(mai_mai_n71_), .Y(mai_mai_n163_));
  INV        m147(.A(mai_mai_n116_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n98_), .B(mai_mai_n17_), .Y(mai_mai_n165_));
  AOI210     m149(.A0(mai_mai_n31_), .A1(mai_mai_n85_), .B0(mai_mai_n165_), .Y(mai_mai_n166_));
  NO3        m150(.A(mai_mai_n166_), .B(mai_mai_n164_), .C(x7), .Y(mai_mai_n167_));
  NA2        m151(.A(mai_mai_n164_), .B(mai_mai_n38_), .Y(mai_mai_n168_));
  OAI210     m152(.A0(mai_mai_n150_), .A1(mai_mai_n122_), .B0(mai_mai_n168_), .Y(mai_mai_n169_));
  NO3        m153(.A(mai_mai_n169_), .B(mai_mai_n167_), .C(mai_mai_n163_), .Y(mai_mai_n170_));
  NO2        m154(.A(mai_mai_n170_), .B(x3), .Y(mai_mai_n171_));
  NO3        m155(.A(mai_mai_n171_), .B(mai_mai_n162_), .C(mai_mai_n147_), .Y(mai03));
  NO2        m156(.A(mai_mai_n44_), .B(x3), .Y(mai_mai_n173_));
  INV        m157(.A(x6), .Y(mai_mai_n174_));
  OAI210     m158(.A0(mai_mai_n174_), .A1(mai_mai_n17_), .B0(mai_mai_n98_), .Y(mai_mai_n175_));
  NA2        m159(.A(mai_mai_n175_), .B(mai_mai_n173_), .Y(mai_mai_n176_));
  NA2        m160(.A(x6), .B(mai_mai_n24_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n177_), .B(x4), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n179_));
  NA2        m163(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n180_));
  NO2        m164(.A(mai_mai_n180_), .B(mai_mai_n177_), .Y(mai_mai_n181_));
  NA2        m165(.A(x9), .B(mai_mai_n50_), .Y(mai_mai_n182_));
  NA2        m166(.A(mai_mai_n182_), .B(x4), .Y(mai_mai_n183_));
  INV        m167(.A(mai_mai_n177_), .Y(mai_mai_n184_));
  AOI210     m168(.A0(mai_mai_n24_), .A1(x3), .B0(mai_mai_n158_), .Y(mai_mai_n185_));
  AOI220     m169(.A0(mai_mai_n185_), .A1(mai_mai_n184_), .B0(mai_mai_n183_), .B1(mai_mai_n181_), .Y(mai_mai_n186_));
  NO2        m170(.A(x5), .B(x1), .Y(mai_mai_n187_));
  NA2        m171(.A(mai_mai_n187_), .B(mai_mai_n17_), .Y(mai_mai_n188_));
  NO2        m172(.A(mai_mai_n180_), .B(mai_mai_n149_), .Y(mai_mai_n189_));
  NA2        m173(.A(mai_mai_n385_), .B(mai_mai_n44_), .Y(mai_mai_n190_));
  NA3        m174(.A(mai_mai_n190_), .B(mai_mai_n186_), .C(mai_mai_n176_), .Y(mai_mai_n191_));
  NO2        m175(.A(mai_mai_n44_), .B(mai_mai_n39_), .Y(mai_mai_n192_));
  NO2        m176(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n193_));
  NA2        m177(.A(mai_mai_n58_), .B(mai_mai_n85_), .Y(mai_mai_n194_));
  NA3        m178(.A(mai_mai_n194_), .B(mai_mai_n193_), .C(x6), .Y(mai_mai_n195_));
  AOI210     m179(.A0(mai_mai_n195_), .A1(mai_mai_n77_), .B0(mai_mai_n137_), .Y(mai_mai_n196_));
  BUFFER     m180(.A(mai_mai_n196_), .Y(mai_mai_n197_));
  NA2        m181(.A(mai_mai_n39_), .B(mai_mai_n50_), .Y(mai_mai_n198_));
  NA2        m182(.A(mai_mai_n126_), .B(mai_mai_n84_), .Y(mai_mai_n199_));
  NA2        m183(.A(x6), .B(mai_mai_n44_), .Y(mai_mai_n200_));
  NO2        m184(.A(mai_mai_n141_), .B(mai_mai_n39_), .Y(mai_mai_n201_));
  OAI210     m185(.A0(mai_mai_n201_), .A1(mai_mai_n189_), .B0(mai_mai_n381_), .Y(mai_mai_n202_));
  NA2        m186(.A(x5), .B(mai_mai_n120_), .Y(mai_mai_n203_));
  NA2        m187(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  NA2        m188(.A(mai_mai_n204_), .B(x2), .Y(mai_mai_n205_));
  NA3        m189(.A(mai_mai_n205_), .B(mai_mai_n199_), .C(mai_mai_n197_), .Y(mai_mai_n206_));
  AOI210     m190(.A0(mai_mai_n191_), .A1(x8), .B0(mai_mai_n206_), .Y(mai_mai_n207_));
  NO2        m191(.A(mai_mai_n85_), .B(x3), .Y(mai_mai_n208_));
  NA2        m192(.A(mai_mai_n208_), .B(mai_mai_n178_), .Y(mai_mai_n209_));
  NO2        m193(.A(mai_mai_n209_), .B(x2), .Y(mai_mai_n210_));
  NO2        m194(.A(x4), .B(mai_mai_n50_), .Y(mai_mai_n211_));
  AOI220     m195(.A0(mai_mai_n178_), .A1(mai_mai_n165_), .B0(mai_mai_n211_), .B1(mai_mai_n61_), .Y(mai_mai_n212_));
  NA2        m196(.A(mai_mai_n58_), .B(x6), .Y(mai_mai_n213_));
  NA3        m197(.A(mai_mai_n24_), .B(x3), .C(x2), .Y(mai_mai_n214_));
  AOI210     m198(.A0(mai_mai_n214_), .A1(mai_mai_n125_), .B0(mai_mai_n213_), .Y(mai_mai_n215_));
  NA2        m199(.A(mai_mai_n39_), .B(mai_mai_n17_), .Y(mai_mai_n216_));
  NO2        m200(.A(mai_mai_n216_), .B(mai_mai_n24_), .Y(mai_mai_n217_));
  OAI210     m201(.A0(mai_mai_n217_), .A1(mai_mai_n215_), .B0(mai_mai_n108_), .Y(mai_mai_n218_));
  NO2        m202(.A(mai_mai_n180_), .B(x6), .Y(mai_mai_n219_));
  NA4        m203(.A(mai_mai_n389_), .B(mai_mai_n218_), .C(mai_mai_n212_), .D(mai_mai_n137_), .Y(mai_mai_n220_));
  NA2        m204(.A(x5), .B(mai_mai_n193_), .Y(mai_mai_n221_));
  NO2        m205(.A(x9), .B(x6), .Y(mai_mai_n222_));
  NO2        m206(.A(mai_mai_n125_), .B(mai_mai_n18_), .Y(mai_mai_n223_));
  NAi21      m207(.An(mai_mai_n223_), .B(mai_mai_n214_), .Y(mai_mai_n224_));
  AOI210     m208(.A0(mai_mai_n224_), .A1(mai_mai_n222_), .B0(mai_mai_n382_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n225_), .B(mai_mai_n221_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n58_), .B(x2), .Y(mai_mai_n227_));
  INV        m211(.A(mai_mai_n221_), .Y(mai_mai_n228_));
  NO3        m212(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n229_));
  NA2        m213(.A(mai_mai_n98_), .B(mai_mai_n24_), .Y(mai_mai_n230_));
  NA2        m214(.A(x6), .B(x2), .Y(mai_mai_n231_));
  NO2        m215(.A(mai_mai_n231_), .B(mai_mai_n149_), .Y(mai_mai_n232_));
  AOI210     m216(.A0(mai_mai_n230_), .A1(mai_mai_n229_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  OAI220     m217(.A0(mai_mai_n233_), .A1(mai_mai_n39_), .B0(mai_mai_n155_), .B1(mai_mai_n42_), .Y(mai_mai_n234_));
  OAI210     m218(.A0(mai_mai_n234_), .A1(mai_mai_n228_), .B0(mai_mai_n226_), .Y(mai_mai_n235_));
  NA2        m219(.A(x4), .B(x0), .Y(mai_mai_n236_));
  NA2        m220(.A(x6), .B(mai_mai_n38_), .Y(mai_mai_n237_));
  AOI210     m221(.A0(mai_mai_n237_), .A1(mai_mai_n235_), .B0(x8), .Y(mai_mai_n238_));
  NA2        m222(.A(mai_mai_n223_), .B(mai_mai_n58_), .Y(mai_mai_n239_));
  NA2        m223(.A(x0), .B(mai_mai_n20_), .Y(mai_mai_n240_));
  AOI210     m224(.A0(mai_mai_n240_), .A1(mai_mai_n239_), .B0(mai_mai_n198_), .Y(mai_mai_n241_));
  NO4        m225(.A(mai_mai_n241_), .B(mai_mai_n238_), .C(mai_mai_n220_), .D(mai_mai_n210_), .Y(mai_mai_n242_));
  NO2        m226(.A(mai_mai_n143_), .B(x1), .Y(mai_mai_n243_));
  NO2        m227(.A(x3), .B(mai_mai_n32_), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n244_), .A1(mai_mai_n219_), .B0(x2), .Y(mai_mai_n245_));
  OAI210     m229(.A0(x0), .A1(x6), .B0(mai_mai_n40_), .Y(mai_mai_n246_));
  AOI210     m230(.A0(mai_mai_n246_), .A1(mai_mai_n245_), .B0(mai_mai_n164_), .Y(mai_mai_n247_));
  NOi21      m231(.An(mai_mai_n231_), .B(mai_mai_n17_), .Y(mai_mai_n248_));
  NA3        m232(.A(mai_mai_n248_), .B(mai_mai_n187_), .C(mai_mai_n36_), .Y(mai_mai_n249_));
  AOI210     m233(.A0(mai_mai_n32_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n250_), .B(mai_mai_n142_), .Y(mai_mai_n251_));
  NA2        m235(.A(x3), .B(x2), .Y(mai_mai_n252_));
  AOI220     m236(.A0(mai_mai_n252_), .A1(mai_mai_n198_), .B0(mai_mai_n251_), .B1(mai_mai_n249_), .Y(mai_mai_n253_));
  NAi21      m237(.An(x4), .B(x0), .Y(mai_mai_n254_));
  OAI210     m238(.A0(mai_mai_n250_), .A1(mai_mai_n248_), .B0(x2), .Y(mai_mai_n255_));
  NA2        m239(.A(mai_mai_n255_), .B(mai_mai_n76_), .Y(mai_mai_n256_));
  NO2        m240(.A(mai_mai_n256_), .B(mai_mai_n24_), .Y(mai_mai_n257_));
  NA3        m241(.A(mai_mai_n32_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n258_));
  OAI210     m242(.A0(mai_mai_n250_), .A1(mai_mai_n248_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  INV        m243(.A(mai_mai_n189_), .Y(mai_mai_n260_));
  NA2        m244(.A(mai_mai_n32_), .B(mai_mai_n39_), .Y(mai_mai_n261_));
  OR2        m245(.A(mai_mai_n261_), .B(mai_mai_n236_), .Y(mai_mai_n262_));
  OAI220     m246(.A0(mai_mai_n262_), .A1(mai_mai_n141_), .B0(mai_mai_n200_), .B1(mai_mai_n260_), .Y(mai_mai_n263_));
  AO210      m247(.A0(mai_mai_n259_), .A1(mai_mai_n133_), .B0(mai_mai_n263_), .Y(mai_mai_n264_));
  NO4        m248(.A(mai_mai_n264_), .B(mai_mai_n257_), .C(mai_mai_n253_), .D(mai_mai_n247_), .Y(mai_mai_n265_));
  OAI210     m249(.A0(mai_mai_n242_), .A1(mai_mai_n207_), .B0(mai_mai_n265_), .Y(mai04));
  OAI210     m250(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n267_));
  NA3        m251(.A(mai_mai_n267_), .B(mai_mai_n229_), .C(mai_mai_n78_), .Y(mai_mai_n268_));
  NO2        m252(.A(x2), .B(x1), .Y(mai_mai_n269_));
  OAI210     m253(.A0(mai_mai_n216_), .A1(mai_mai_n269_), .B0(mai_mai_n32_), .Y(mai_mai_n270_));
  INV        m254(.A(mai_mai_n254_), .Y(mai_mai_n271_));
  OAI210     m255(.A0(mai_mai_n50_), .A1(mai_mai_n271_), .B0(mai_mai_n208_), .Y(mai_mai_n272_));
  NO2        m256(.A(mai_mai_n227_), .B(mai_mai_n83_), .Y(mai_mai_n273_));
  NO2        m257(.A(mai_mai_n252_), .B(mai_mai_n179_), .Y(mai_mai_n274_));
  NA2        m258(.A(x9), .B(x0), .Y(mai_mai_n275_));
  NO2        m259(.A(mai_mai_n83_), .B(mai_mai_n275_), .Y(mai_mai_n276_));
  OAI210     m260(.A0(mai_mai_n276_), .A1(mai_mai_n274_), .B0(mai_mai_n85_), .Y(mai_mai_n277_));
  NA3        m261(.A(mai_mai_n277_), .B(x6), .C(mai_mai_n272_), .Y(mai_mai_n278_));
  NA2        m262(.A(mai_mai_n278_), .B(mai_mai_n270_), .Y(mai_mai_n279_));
  OAI210     m263(.A0(mai_mai_n106_), .A1(mai_mai_n98_), .B0(mai_mai_n153_), .Y(mai_mai_n280_));
  NA3        m264(.A(mai_mai_n280_), .B(x6), .C(x3), .Y(mai_mai_n281_));
  NOi21      m265(.An(mai_mai_n135_), .B(mai_mai_n117_), .Y(mai_mai_n282_));
  AOI210     m266(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n283_));
  OAI220     m267(.A0(mai_mai_n283_), .A1(mai_mai_n261_), .B0(mai_mai_n227_), .B1(mai_mai_n258_), .Y(mai_mai_n284_));
  AOI210     m268(.A0(mai_mai_n282_), .A1(x6), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  NA2        m269(.A(mai_mai_n273_), .B(mai_mai_n85_), .Y(mai_mai_n286_));
  NA3        m270(.A(mai_mai_n286_), .B(mai_mai_n285_), .C(mai_mai_n281_), .Y(mai_mai_n287_));
  AOI210     m271(.A0(mai_mai_n287_), .A1(x4), .B0(x7), .Y(mai_mai_n288_));
  NA3        m272(.A(mai_mai_n271_), .B(mai_mai_n182_), .C(mai_mai_n85_), .Y(mai_mai_n289_));
  XO2        m273(.A(x4), .B(x0), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n290_), .B(mai_mai_n105_), .Y(mai_mai_n291_));
  NA2        m275(.A(mai_mai_n291_), .B(x8), .Y(mai_mai_n292_));
  AOI210     m276(.A0(mai_mai_n292_), .A1(mai_mai_n289_), .B0(x3), .Y(mai_mai_n293_));
  NO2        m277(.A(mai_mai_n85_), .B(x4), .Y(mai_mai_n294_));
  NA2        m278(.A(mai_mai_n294_), .B(mai_mai_n40_), .Y(mai_mai_n295_));
  NO3        m279(.A(mai_mai_n290_), .B(mai_mai_n143_), .C(x2), .Y(mai_mai_n296_));
  NO3        m280(.A(mai_mai_n194_), .B(mai_mai_n26_), .C(mai_mai_n23_), .Y(mai_mai_n297_));
  NO2        m281(.A(mai_mai_n297_), .B(mai_mai_n296_), .Y(mai_mai_n298_));
  NA3        m282(.A(mai_mai_n298_), .B(mai_mai_n295_), .C(x6), .Y(mai_mai_n299_));
  BUFFER     m283(.A(mai_mai_n294_), .Y(mai_mai_n300_));
  INV        m284(.A(mai_mai_n98_), .Y(mai_mai_n301_));
  NA2        m285(.A(mai_mai_n301_), .B(mai_mai_n300_), .Y(mai_mai_n302_));
  NO2        m286(.A(mai_mai_n135_), .B(mai_mai_n75_), .Y(mai_mai_n303_));
  NO2        m287(.A(mai_mai_n31_), .B(x2), .Y(mai_mai_n304_));
  NA2        m288(.A(mai_mai_n304_), .B(mai_mai_n303_), .Y(mai_mai_n305_));
  NA2        m289(.A(mai_mai_n302_), .B(mai_mai_n305_), .Y(mai_mai_n306_));
  OAI220     m290(.A0(mai_mai_n306_), .A1(x6), .B0(mai_mai_n299_), .B1(mai_mai_n293_), .Y(mai_mai_n307_));
  OAI210     m291(.A0(x6), .A1(mai_mai_n44_), .B0(mai_mai_n38_), .Y(mai_mai_n308_));
  OAI210     m292(.A0(mai_mai_n308_), .A1(mai_mai_n85_), .B0(mai_mai_n262_), .Y(mai_mai_n309_));
  AOI210     m293(.A0(mai_mai_n309_), .A1(mai_mai_n18_), .B0(mai_mai_n137_), .Y(mai_mai_n310_));
  AO220      m294(.A0(mai_mai_n310_), .A1(mai_mai_n307_), .B0(mai_mai_n288_), .B1(mai_mai_n279_), .Y(mai_mai_n311_));
  NA2        m295(.A(mai_mai_n304_), .B(x6), .Y(mai_mai_n312_));
  AOI210     m296(.A0(x6), .A1(x1), .B0(mai_mai_n136_), .Y(mai_mai_n313_));
  NA2        m297(.A(mai_mai_n294_), .B(x0), .Y(mai_mai_n314_));
  NA2        m298(.A(mai_mai_n77_), .B(x6), .Y(mai_mai_n315_));
  OAI210     m299(.A0(mai_mai_n314_), .A1(mai_mai_n313_), .B0(mai_mai_n315_), .Y(mai_mai_n316_));
  NA2        m300(.A(mai_mai_n316_), .B(mai_mai_n312_), .Y(mai_mai_n317_));
  NA3        m301(.A(mai_mai_n317_), .B(mai_mai_n311_), .C(mai_mai_n268_), .Y(mai_mai_n318_));
  NA3        m302(.A(x2), .B(mai_mai_n173_), .C(mai_mai_n137_), .Y(mai_mai_n319_));
  NO2        m303(.A(mai_mai_n386_), .B(mai_mai_n182_), .Y(mai_mai_n320_));
  INV        m304(.A(mai_mai_n320_), .Y(mai_mai_n321_));
  AOI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n319_), .B0(mai_mai_n24_), .Y(mai_mai_n322_));
  OAI210     m306(.A0(mai_mai_n173_), .A1(mai_mai_n62_), .B0(mai_mai_n179_), .Y(mai_mai_n323_));
  NA3        m307(.A(mai_mai_n388_), .B(mai_mai_n193_), .C(x8), .Y(mai_mai_n324_));
  AOI210     m308(.A0(mai_mai_n324_), .A1(mai_mai_n323_), .B0(mai_mai_n24_), .Y(mai_mai_n325_));
  AOI210     m309(.A0(mai_mai_n107_), .A1(mai_mai_n106_), .B0(mai_mai_n38_), .Y(mai_mai_n326_));
  NOi31      m310(.An(mai_mai_n326_), .B(x3), .C(mai_mai_n159_), .Y(mai_mai_n327_));
  OAI210     m311(.A0(mai_mai_n327_), .A1(mai_mai_n325_), .B0(mai_mai_n134_), .Y(mai_mai_n328_));
  NAi31      m312(.An(mai_mai_n46_), .B(mai_mai_n243_), .C(mai_mai_n154_), .Y(mai_mai_n329_));
  NA2        m313(.A(mai_mai_n329_), .B(mai_mai_n328_), .Y(mai_mai_n330_));
  OAI210     m314(.A0(mai_mai_n330_), .A1(mai_mai_n322_), .B0(x6), .Y(mai_mai_n331_));
  INV        m315(.A(mai_mai_n121_), .Y(mai_mai_n332_));
  NA3        m316(.A(mai_mai_n51_), .B(mai_mai_n34_), .C(mai_mai_n28_), .Y(mai_mai_n333_));
  AOI220     m317(.A0(mai_mai_n333_), .A1(mai_mai_n332_), .B0(mai_mai_n36_), .B1(mai_mai_n29_), .Y(mai_mai_n334_));
  AOI220     m318(.A0(mai_mai_n384_), .A1(mai_mai_n192_), .B0(mai_mai_n173_), .B1(mai_mai_n137_), .Y(mai_mai_n335_));
  AOI210     m319(.A0(mai_mai_n113_), .A1(mai_mai_n211_), .B0(x1), .Y(mai_mai_n336_));
  OAI210     m320(.A0(mai_mai_n335_), .A1(x8), .B0(mai_mai_n336_), .Y(mai_mai_n337_));
  NO4        m321(.A(x8), .B(mai_mai_n254_), .C(x9), .D(x2), .Y(mai_mai_n338_));
  NO3        m322(.A(mai_mai_n111_), .B(mai_mai_n338_), .C(mai_mai_n18_), .Y(mai_mai_n339_));
  NA2        m323(.A(mai_mai_n303_), .B(mai_mai_n137_), .Y(mai_mai_n340_));
  NA2        m324(.A(mai_mai_n340_), .B(mai_mai_n339_), .Y(mai_mai_n341_));
  OAI210     m325(.A0(mai_mai_n337_), .A1(mai_mai_n334_), .B0(mai_mai_n341_), .Y(mai_mai_n342_));
  NOi31      m326(.An(mai_mai_n384_), .B(mai_mai_n29_), .C(x8), .Y(mai_mai_n343_));
  AOI210     m327(.A0(mai_mai_n34_), .A1(x9), .B0(mai_mai_n119_), .Y(mai_mai_n344_));
  NO3        m328(.A(mai_mai_n344_), .B(mai_mai_n111_), .C(mai_mai_n39_), .Y(mai_mai_n345_));
  NO2        m329(.A(mai_mai_n56_), .B(mai_mai_n110_), .Y(mai_mai_n346_));
  NO2        m330(.A(mai_mai_n346_), .B(x3), .Y(mai_mai_n347_));
  NO3        m331(.A(mai_mai_n347_), .B(mai_mai_n345_), .C(x2), .Y(mai_mai_n348_));
  NO2        m332(.A(mai_mai_n348_), .B(mai_mai_n343_), .Y(mai_mai_n349_));
  AOI210     m333(.A0(mai_mai_n349_), .A1(mai_mai_n342_), .B0(mai_mai_n24_), .Y(mai_mai_n350_));
  NA2        m334(.A(mai_mai_n383_), .B(mai_mai_n326_), .Y(mai_mai_n351_));
  NO2        m335(.A(mai_mai_n351_), .B(mai_mai_n97_), .Y(mai_mai_n352_));
  NA2        m336(.A(mai_mai_n352_), .B(x7), .Y(mai_mai_n353_));
  NA2        m337(.A(mai_mai_n194_), .B(x7), .Y(mai_mai_n354_));
  NA3        m338(.A(mai_mai_n354_), .B(mai_mai_n136_), .C(mai_mai_n120_), .Y(mai_mai_n355_));
  NA2        m339(.A(mai_mai_n355_), .B(mai_mai_n353_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n356_), .A1(mai_mai_n350_), .B0(mai_mai_n32_), .Y(mai_mai_n357_));
  NA2        m341(.A(mai_mai_n216_), .B(mai_mai_n21_), .Y(mai_mai_n358_));
  NO2        m342(.A(mai_mai_n141_), .B(mai_mai_n121_), .Y(mai_mai_n359_));
  NA2        m343(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n360_));
  AOI210     m344(.A0(mai_mai_n360_), .A1(mai_mai_n144_), .B0(mai_mai_n26_), .Y(mai_mai_n361_));
  AOI220     m345(.A0(x3), .A1(mai_mai_n85_), .B0(mai_mai_n135_), .B1(mai_mai_n388_), .Y(mai_mai_n362_));
  NA2        m346(.A(mai_mai_n362_), .B(mai_mai_n83_), .Y(mai_mai_n363_));
  NA2        m347(.A(mai_mai_n363_), .B(mai_mai_n154_), .Y(mai_mai_n364_));
  OAI220     m348(.A0(x3), .A1(mai_mai_n63_), .B0(mai_mai_n141_), .B1(mai_mai_n39_), .Y(mai_mai_n365_));
  NA2        m349(.A(x3), .B(mai_mai_n50_), .Y(mai_mai_n366_));
  AOI210     m350(.A0(x2), .A1(mai_mai_n25_), .B0(mai_mai_n68_), .Y(mai_mai_n367_));
  OAI210     m351(.A0(mai_mai_n134_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n368_));
  AOI210     m352(.A0(x2), .A1(mai_mai_n368_), .B0(mai_mai_n367_), .Y(mai_mai_n369_));
  OAI210     m353(.A0(mai_mai_n138_), .A1(mai_mai_n366_), .B0(mai_mai_n369_), .Y(mai_mai_n370_));
  AOI220     m354(.A0(mai_mai_n370_), .A1(x0), .B0(mai_mai_n365_), .B1(mai_mai_n121_), .Y(mai_mai_n371_));
  AOI210     m355(.A0(mai_mai_n371_), .A1(mai_mai_n364_), .B0(mai_mai_n200_), .Y(mai_mai_n372_));
  INV        m356(.A(x5), .Y(mai_mai_n373_));
  NO4        m357(.A(mai_mai_n98_), .B(mai_mai_n373_), .C(mai_mai_n56_), .D(mai_mai_n29_), .Y(mai_mai_n374_));
  NO3        m358(.A(mai_mai_n374_), .B(mai_mai_n372_), .C(mai_mai_n361_), .Y(mai_mai_n375_));
  NA3        m359(.A(mai_mai_n375_), .B(mai_mai_n357_), .C(mai_mai_n331_), .Y(mai_mai_n376_));
  AOI210     m360(.A0(mai_mai_n318_), .A1(mai_mai_n24_), .B0(mai_mai_n376_), .Y(mai05));
  INV        m361(.A(mai_mai_n105_), .Y(mai_mai_n380_));
  INV        m362(.A(x6), .Y(mai_mai_n381_));
  INV        m363(.A(x4), .Y(mai_mai_n382_));
  INV        m364(.A(x4), .Y(mai_mai_n383_));
  INV        m365(.A(x0), .Y(mai_mai_n384_));
  INV        m366(.A(mai_mai_n188_), .Y(mai_mai_n385_));
  INV        m367(.A(x0), .Y(mai_mai_n386_));
  INV        m368(.A(mai_mai_n103_), .Y(mai_mai_n387_));
  INV        m369(.A(x1), .Y(mai_mai_n388_));
  INV        m370(.A(mai_mai_n130_), .Y(mai_mai_n389_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NA2        u005(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n22_));
  INV        u006(.A(x5), .Y(men_men_n23_));
  NA2        u007(.A(x7), .B(x6), .Y(men_men_n24_));
  NA2        u008(.A(x8), .B(x3), .Y(men_men_n25_));
  NA2        u009(.A(x4), .B(x2), .Y(men_men_n26_));
  NO3        u010(.A(men_men_n26_), .B(men_men_n24_), .C(men_men_n23_), .Y(men_men_n27_));
  NO2        u011(.A(men_men_n27_), .B(men_men_n22_), .Y(men_men_n28_));
  NO2        u012(.A(x4), .B(x3), .Y(men_men_n29_));
  INV        u013(.A(men_men_n29_), .Y(men_men_n30_));
  OA210      u014(.A0(men_men_n30_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n31_));
  NO2        u015(.A(men_men_n31_), .B(men_men_n28_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NA2        u018(.A(x4), .B(x3), .Y(men_men_n35_));
  NO2        u019(.A(x0), .B(men_men_n35_), .Y(men_men_n36_));
  NO2        u020(.A(x2), .B(x0), .Y(men_men_n37_));
  INV        u021(.A(x3), .Y(men_men_n38_));
  NO2        u022(.A(men_men_n38_), .B(men_men_n18_), .Y(men_men_n39_));
  INV        u023(.A(men_men_n39_), .Y(men_men_n40_));
  OAI210     u024(.A0(men_men_n23_), .A1(men_men_n40_), .B0(men_men_n37_), .Y(men_men_n41_));
  INV        u025(.A(x4), .Y(men_men_n42_));
  NO2        u026(.A(men_men_n42_), .B(men_men_n17_), .Y(men_men_n43_));
  NA2        u027(.A(men_men_n43_), .B(x2), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n20_), .B0(men_men_n41_), .Y(men_men_n45_));
  NA2        u029(.A(men_men_n20_), .B(men_men_n19_), .Y(men_men_n46_));
  INV        u030(.A(x2), .Y(men_men_n47_));
  NO2        u031(.A(men_men_n47_), .B(men_men_n17_), .Y(men_men_n48_));
  NA2        u032(.A(men_men_n38_), .B(men_men_n18_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(men_men_n48_), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n46_), .A1(men_men_n30_), .B0(men_men_n50_), .Y(men_men_n51_));
  NO3        u035(.A(men_men_n51_), .B(men_men_n45_), .C(men_men_n36_), .Y(men01));
  NA2        u036(.A(x8), .B(x7), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n38_), .B(x1), .Y(men_men_n54_));
  INV        u038(.A(x9), .Y(men_men_n55_));
  NO2        u039(.A(men_men_n55_), .B(men_men_n34_), .Y(men_men_n56_));
  INV        u040(.A(men_men_n56_), .Y(men_men_n57_));
  NO2        u041(.A(men_men_n57_), .B(men_men_n54_), .Y(men_men_n58_));
  NO2        u042(.A(x7), .B(x6), .Y(men_men_n59_));
  NO2        u043(.A(men_men_n54_), .B(x5), .Y(men_men_n60_));
  NO2        u044(.A(x8), .B(x2), .Y(men_men_n61_));
  OAI210     u045(.A0(men_men_n49_), .A1(men_men_n20_), .B0(x2), .Y(men_men_n62_));
  NAi31      u046(.An(x1), .B(x9), .C(x5), .Y(men_men_n63_));
  OAI220     u047(.A0(men_men_n63_), .A1(men_men_n38_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n64_));
  OAI210     u048(.A0(men_men_n64_), .A1(men_men_n58_), .B0(x4), .Y(men_men_n65_));
  NA2        u049(.A(men_men_n42_), .B(x2), .Y(men_men_n66_));
  OAI210     u050(.A0(men_men_n66_), .A1(men_men_n49_), .B0(x0), .Y(men_men_n67_));
  NA2        u051(.A(x5), .B(x3), .Y(men_men_n68_));
  NO2        u052(.A(x8), .B(x6), .Y(men_men_n69_));
  NO4        u053(.A(men_men_n69_), .B(men_men_n68_), .C(men_men_n59_), .D(men_men_n47_), .Y(men_men_n70_));
  NAi21      u054(.An(x4), .B(x3), .Y(men_men_n71_));
  INV        u055(.A(men_men_n71_), .Y(men_men_n72_));
  NO2        u056(.A(men_men_n72_), .B(men_men_n20_), .Y(men_men_n73_));
  NO2        u057(.A(x4), .B(x2), .Y(men_men_n74_));
  NO2        u058(.A(men_men_n74_), .B(x3), .Y(men_men_n75_));
  NO3        u059(.A(men_men_n75_), .B(men_men_n73_), .C(men_men_n18_), .Y(men_men_n76_));
  NO3        u060(.A(men_men_n76_), .B(men_men_n70_), .C(men_men_n67_), .Y(men_men_n77_));
  NO4        u061(.A(men_men_n21_), .B(x6), .C(men_men_n38_), .D(x1), .Y(men_men_n78_));
  NA2        u062(.A(men_men_n55_), .B(men_men_n42_), .Y(men_men_n79_));
  INV        u063(.A(men_men_n79_), .Y(men_men_n80_));
  OAI210     u064(.A0(men_men_n78_), .A1(men_men_n60_), .B0(men_men_n80_), .Y(men_men_n81_));
  NA2        u065(.A(x3), .B(men_men_n18_), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(men_men_n23_), .Y(men_men_n83_));
  INV        u067(.A(x8), .Y(men_men_n84_));
  NA2        u068(.A(x2), .B(x1), .Y(men_men_n85_));
  NO2        u069(.A(x2), .B(men_men_n83_), .Y(men_men_n86_));
  NO2        u070(.A(men_men_n86_), .B(men_men_n24_), .Y(men_men_n87_));
  AOI210     u071(.A0(men_men_n49_), .A1(men_men_n23_), .B0(men_men_n47_), .Y(men_men_n88_));
  NO3        u072(.A(x4), .B(men_men_n88_), .C(men_men_n87_), .Y(men_men_n89_));
  NO2        u073(.A(men_men_n42_), .B(men_men_n47_), .Y(men_men_n90_));
  OAI210     u074(.A0(men_men_n90_), .A1(men_men_n38_), .B0(men_men_n18_), .Y(men_men_n91_));
  INV        u075(.A(men_men_n91_), .Y(men_men_n92_));
  NO2        u076(.A(x3), .B(x2), .Y(men_men_n93_));
  NA3        u077(.A(men_men_n93_), .B(men_men_n24_), .C(men_men_n23_), .Y(men_men_n94_));
  AOI210     u078(.A0(x8), .A1(x6), .B0(men_men_n94_), .Y(men_men_n95_));
  NA2        u079(.A(men_men_n47_), .B(x1), .Y(men_men_n96_));
  NO4        u080(.A(x0), .B(men_men_n95_), .C(men_men_n92_), .D(men_men_n89_), .Y(men_men_n97_));
  AO220      u081(.A0(men_men_n97_), .A1(men_men_n81_), .B0(men_men_n77_), .B1(men_men_n65_), .Y(men02));
  NO2        u082(.A(x3), .B(men_men_n47_), .Y(men_men_n99_));
  NO2        u083(.A(x8), .B(men_men_n18_), .Y(men_men_n100_));
  NA2        u084(.A(men_men_n38_), .B(x0), .Y(men_men_n101_));
  OAI210     u085(.A0(men_men_n79_), .A1(x0), .B0(men_men_n101_), .Y(men_men_n102_));
  AOI220     u086(.A0(men_men_n102_), .A1(men_men_n100_), .B0(men_men_n99_), .B1(x4), .Y(men_men_n103_));
  NO3        u087(.A(men_men_n103_), .B(x7), .C(x5), .Y(men_men_n104_));
  NA2        u088(.A(x9), .B(x2), .Y(men_men_n105_));
  OR2        u089(.A(x8), .B(x0), .Y(men_men_n106_));
  INV        u090(.A(men_men_n106_), .Y(men_men_n107_));
  INV        u091(.A(x2), .Y(men_men_n108_));
  NO2        u092(.A(x4), .B(x1), .Y(men_men_n109_));
  NA3        u093(.A(men_men_n109_), .B(men_men_n106_), .C(men_men_n53_), .Y(men_men_n110_));
  NOi21      u094(.An(x0), .B(x1), .Y(men_men_n111_));
  NO3        u095(.A(x9), .B(x8), .C(x7), .Y(men_men_n112_));
  NOi21      u096(.An(x0), .B(x4), .Y(men_men_n113_));
  NAi21      u097(.An(x8), .B(x7), .Y(men_men_n114_));
  NO2        u098(.A(men_men_n110_), .B(men_men_n68_), .Y(men_men_n115_));
  NO2        u099(.A(x5), .B(men_men_n42_), .Y(men_men_n116_));
  NA2        u100(.A(x2), .B(men_men_n18_), .Y(men_men_n117_));
  AOI210     u101(.A0(men_men_n117_), .A1(men_men_n96_), .B0(men_men_n101_), .Y(men_men_n118_));
  OAI210     u102(.A0(men_men_n118_), .A1(men_men_n33_), .B0(men_men_n116_), .Y(men_men_n119_));
  NAi21      u103(.An(x0), .B(x4), .Y(men_men_n120_));
  NO2        u104(.A(men_men_n120_), .B(x1), .Y(men_men_n121_));
  NO2        u105(.A(x7), .B(x0), .Y(men_men_n122_));
  NO2        u106(.A(men_men_n74_), .B(men_men_n90_), .Y(men_men_n123_));
  NO2        u107(.A(men_men_n123_), .B(x3), .Y(men_men_n124_));
  OAI210     u108(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n124_), .Y(men_men_n125_));
  NO2        u109(.A(men_men_n21_), .B(men_men_n38_), .Y(men_men_n126_));
  NA2        u110(.A(x5), .B(x0), .Y(men_men_n127_));
  NO2        u111(.A(men_men_n42_), .B(x2), .Y(men_men_n128_));
  NA2        u112(.A(men_men_n128_), .B(men_men_n126_), .Y(men_men_n129_));
  NA4        u113(.A(men_men_n129_), .B(men_men_n125_), .C(men_men_n119_), .D(men_men_n34_), .Y(men_men_n130_));
  NO3        u114(.A(men_men_n130_), .B(men_men_n115_), .C(men_men_n104_), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n26_), .B(men_men_n23_), .Y(men_men_n132_));
  AOI220     u116(.A0(men_men_n111_), .A1(men_men_n132_), .B0(men_men_n60_), .B1(men_men_n17_), .Y(men_men_n133_));
  NO3        u117(.A(men_men_n133_), .B(men_men_n53_), .C(men_men_n55_), .Y(men_men_n134_));
  NA2        u118(.A(x7), .B(x3), .Y(men_men_n135_));
  NO2        u119(.A(men_men_n395_), .B(x5), .Y(men_men_n136_));
  NO2        u120(.A(x9), .B(x7), .Y(men_men_n137_));
  NOi21      u121(.An(x8), .B(x0), .Y(men_men_n138_));
  NO2        u122(.A(men_men_n38_), .B(x2), .Y(men_men_n139_));
  INV        u123(.A(x7), .Y(men_men_n140_));
  NA2        u124(.A(men_men_n140_), .B(men_men_n18_), .Y(men_men_n141_));
  AOI220     u125(.A0(men_men_n141_), .A1(men_men_n139_), .B0(men_men_n99_), .B1(x7), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n23_), .B(x4), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n143_), .B(men_men_n113_), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n144_), .B(men_men_n142_), .Y(men_men_n145_));
  AOI210     u129(.A0(men_men_n138_), .A1(men_men_n136_), .B0(men_men_n145_), .Y(men_men_n146_));
  OAI210     u130(.A0(men_men_n135_), .A1(men_men_n44_), .B0(men_men_n146_), .Y(men_men_n147_));
  NA2        u131(.A(x5), .B(x1), .Y(men_men_n148_));
  INV        u132(.A(men_men_n148_), .Y(men_men_n149_));
  AOI210     u133(.A0(men_men_n149_), .A1(men_men_n113_), .B0(men_men_n34_), .Y(men_men_n150_));
  NO2        u134(.A(men_men_n55_), .B(men_men_n84_), .Y(men_men_n151_));
  NAi21      u135(.An(x2), .B(x7), .Y(men_men_n152_));
  NO3        u136(.A(men_men_n152_), .B(men_men_n151_), .C(men_men_n42_), .Y(men_men_n153_));
  NA2        u137(.A(men_men_n153_), .B(men_men_n60_), .Y(men_men_n154_));
  NAi31      u138(.An(men_men_n68_), .B(x7), .C(men_men_n33_), .Y(men_men_n155_));
  NA3        u139(.A(men_men_n155_), .B(men_men_n154_), .C(men_men_n150_), .Y(men_men_n156_));
  NO3        u140(.A(men_men_n156_), .B(men_men_n147_), .C(men_men_n134_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n157_), .B(men_men_n131_), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n127_), .B(men_men_n123_), .Y(men_men_n159_));
  NA2        u143(.A(men_men_n23_), .B(men_men_n18_), .Y(men_men_n160_));
  NA2        u144(.A(men_men_n23_), .B(men_men_n17_), .Y(men_men_n161_));
  NA3        u145(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n22_), .Y(men_men_n162_));
  AN2        u146(.A(men_men_n162_), .B(men_men_n128_), .Y(men_men_n163_));
  NA2        u147(.A(x8), .B(x0), .Y(men_men_n164_));
  NO2        u148(.A(men_men_n140_), .B(men_men_n23_), .Y(men_men_n165_));
  NO2        u149(.A(men_men_n111_), .B(x4), .Y(men_men_n166_));
  NA2        u150(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  INV        u151(.A(men_men_n167_), .Y(men_men_n168_));
  NA2        u152(.A(x2), .B(x0), .Y(men_men_n169_));
  NA2        u153(.A(x4), .B(x1), .Y(men_men_n170_));
  NO3        u154(.A(men_men_n168_), .B(men_men_n163_), .C(men_men_n159_), .Y(men_men_n171_));
  NO2        u155(.A(men_men_n171_), .B(men_men_n38_), .Y(men_men_n172_));
  NO2        u156(.A(men_men_n162_), .B(men_men_n66_), .Y(men_men_n173_));
  INV        u157(.A(men_men_n116_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n161_), .B(men_men_n123_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n175_), .B(men_men_n173_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n176_), .B(x3), .Y(men_men_n177_));
  NO3        u161(.A(men_men_n177_), .B(men_men_n172_), .C(men_men_n158_), .Y(men03));
  NO2        u162(.A(men_men_n42_), .B(x3), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n47_), .B(x1), .Y(men_men_n180_));
  OAI210     u164(.A0(men_men_n180_), .A1(men_men_n23_), .B0(men_men_n56_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n181_), .B(men_men_n17_), .Y(men_men_n182_));
  NA2        u166(.A(men_men_n182_), .B(men_men_n179_), .Y(men_men_n183_));
  NO2        u167(.A(men_men_n68_), .B(x6), .Y(men_men_n184_));
  NA2        u168(.A(x6), .B(men_men_n23_), .Y(men_men_n185_));
  NO2        u169(.A(men_men_n185_), .B(x4), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n18_), .B(x0), .Y(men_men_n187_));
  AO220      u171(.A0(men_men_n187_), .A1(men_men_n186_), .B0(men_men_n184_), .B1(men_men_n48_), .Y(men_men_n188_));
  NA2        u172(.A(men_men_n188_), .B(men_men_n55_), .Y(men_men_n189_));
  NA2        u173(.A(x3), .B(men_men_n17_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n190_), .B(men_men_n185_), .Y(men_men_n191_));
  NA2        u175(.A(men_men_n185_), .B(men_men_n71_), .Y(men_men_n192_));
  AOI210     u176(.A0(men_men_n23_), .A1(x3), .B0(men_men_n169_), .Y(men_men_n193_));
  AOI210     u177(.A0(men_men_n193_), .A1(men_men_n192_), .B0(men_men_n191_), .Y(men_men_n194_));
  NO3        u178(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n195_));
  NO2        u179(.A(x5), .B(x1), .Y(men_men_n196_));
  AOI220     u180(.A0(men_men_n196_), .A1(men_men_n17_), .B0(men_men_n93_), .B1(x5), .Y(men_men_n197_));
  NO2        u181(.A(men_men_n190_), .B(men_men_n160_), .Y(men_men_n198_));
  INV        u182(.A(men_men_n198_), .Y(men_men_n199_));
  OAI210     u183(.A0(men_men_n197_), .A1(men_men_n57_), .B0(men_men_n199_), .Y(men_men_n200_));
  AOI220     u184(.A0(men_men_n200_), .A1(men_men_n42_), .B0(men_men_n195_), .B1(men_men_n116_), .Y(men_men_n201_));
  NA4        u185(.A(men_men_n201_), .B(men_men_n194_), .C(men_men_n189_), .D(men_men_n183_), .Y(men_men_n202_));
  NO2        u186(.A(men_men_n42_), .B(men_men_n38_), .Y(men_men_n203_));
  NA2        u187(.A(men_men_n203_), .B(men_men_n19_), .Y(men_men_n204_));
  NO2        u188(.A(x3), .B(men_men_n17_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n205_), .B(x6), .Y(men_men_n206_));
  NOi21      u190(.An(men_men_n74_), .B(men_men_n206_), .Y(men_men_n207_));
  NA2        u191(.A(men_men_n55_), .B(men_men_n84_), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n205_), .B(x6), .Y(men_men_n209_));
  AOI210     u193(.A0(men_men_n209_), .A1(men_men_n207_), .B0(men_men_n140_), .Y(men_men_n210_));
  AO210      u194(.A0(men_men_n210_), .A1(men_men_n204_), .B0(men_men_n165_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n38_), .B(men_men_n47_), .Y(men_men_n212_));
  NO3        u196(.A(men_men_n170_), .B(men_men_n55_), .C(x6), .Y(men_men_n213_));
  AOI220     u197(.A0(men_men_n213_), .A1(men_men_n17_), .B0(men_men_n128_), .B1(men_men_n83_), .Y(men_men_n214_));
  NA2        u198(.A(x6), .B(men_men_n42_), .Y(men_men_n215_));
  NA2        u199(.A(men_men_n69_), .B(x4), .Y(men_men_n216_));
  AOI210     u200(.A0(men_men_n216_), .A1(men_men_n215_), .B0(men_men_n68_), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n148_), .B(men_men_n38_), .Y(men_men_n218_));
  OAI210     u202(.A0(men_men_n218_), .A1(men_men_n198_), .B0(x9), .Y(men_men_n219_));
  NA2        u203(.A(men_men_n394_), .B(men_men_n121_), .Y(men_men_n220_));
  NA2        u204(.A(men_men_n116_), .B(x6), .Y(men_men_n221_));
  OAI210     u205(.A0(men_men_n84_), .A1(men_men_n34_), .B0(men_men_n60_), .Y(men_men_n222_));
  NA4        u206(.A(men_men_n222_), .B(men_men_n221_), .C(men_men_n220_), .D(men_men_n219_), .Y(men_men_n223_));
  OAI210     u207(.A0(men_men_n223_), .A1(men_men_n217_), .B0(x2), .Y(men_men_n224_));
  NA3        u208(.A(men_men_n224_), .B(men_men_n214_), .C(men_men_n211_), .Y(men_men_n225_));
  AOI210     u209(.A0(men_men_n202_), .A1(x8), .B0(men_men_n225_), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n84_), .B(x3), .Y(men_men_n227_));
  NO3        u211(.A(men_men_n82_), .B(men_men_n69_), .C(men_men_n23_), .Y(men_men_n228_));
  AOI210     u212(.A0(men_men_n206_), .A1(men_men_n143_), .B0(men_men_n228_), .Y(men_men_n229_));
  NO2        u213(.A(men_men_n229_), .B(x2), .Y(men_men_n230_));
  AOI220     u214(.A0(men_men_n186_), .A1(x0), .B0(x2), .B1(men_men_n60_), .Y(men_men_n231_));
  NA2        u215(.A(men_men_n55_), .B(x6), .Y(men_men_n232_));
  NA3        u216(.A(men_men_n23_), .B(x3), .C(x2), .Y(men_men_n233_));
  INV        u217(.A(men_men_n232_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n234_), .B(men_men_n109_), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n190_), .B(x6), .Y(men_men_n236_));
  NO2        u220(.A(men_men_n190_), .B(x6), .Y(men_men_n237_));
  NAi21      u221(.An(men_men_n151_), .B(men_men_n237_), .Y(men_men_n238_));
  NA3        u222(.A(men_men_n238_), .B(men_men_n236_), .C(men_men_n132_), .Y(men_men_n239_));
  NA4        u223(.A(men_men_n239_), .B(men_men_n235_), .C(men_men_n231_), .D(men_men_n140_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n394_), .B(men_men_n205_), .Y(men_men_n241_));
  NO2        u225(.A(men_men_n127_), .B(men_men_n18_), .Y(men_men_n242_));
  NAi21      u226(.An(men_men_n242_), .B(men_men_n233_), .Y(men_men_n243_));
  NAi21      u227(.An(x1), .B(x4), .Y(men_men_n244_));
  INV        u228(.A(x4), .Y(men_men_n245_));
  NO2        u229(.A(men_men_n245_), .B(men_men_n243_), .Y(men_men_n246_));
  NA2        u230(.A(men_men_n246_), .B(men_men_n241_), .Y(men_men_n247_));
  NA2        u231(.A(men_men_n55_), .B(x2), .Y(men_men_n248_));
  NO2        u232(.A(men_men_n248_), .B(men_men_n241_), .Y(men_men_n249_));
  NO3        u233(.A(x9), .B(x6), .C(x0), .Y(men_men_n250_));
  INV        u234(.A(men_men_n250_), .Y(men_men_n251_));
  OAI210     u235(.A0(men_men_n251_), .A1(men_men_n38_), .B0(men_men_n166_), .Y(men_men_n252_));
  OAI210     u236(.A0(men_men_n252_), .A1(men_men_n249_), .B0(men_men_n247_), .Y(men_men_n253_));
  NA2        u237(.A(x4), .B(x0), .Y(men_men_n254_));
  NO3        u238(.A(men_men_n63_), .B(men_men_n254_), .C(x6), .Y(men_men_n255_));
  AOI210     u239(.A0(men_men_n184_), .A1(men_men_n37_), .B0(men_men_n255_), .Y(men_men_n256_));
  AOI210     u240(.A0(men_men_n256_), .A1(men_men_n253_), .B0(x8), .Y(men_men_n257_));
  OAI210     u241(.A0(men_men_n242_), .A1(men_men_n196_), .B0(x6), .Y(men_men_n258_));
  INV        u242(.A(men_men_n164_), .Y(men_men_n259_));
  OAI210     u243(.A0(men_men_n259_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n260_));
  AOI210     u244(.A0(men_men_n260_), .A1(men_men_n258_), .B0(men_men_n212_), .Y(men_men_n261_));
  NO4        u245(.A(men_men_n261_), .B(men_men_n257_), .C(men_men_n240_), .D(men_men_n230_), .Y(men_men_n262_));
  OAI210     u246(.A0(men_men_n151_), .A1(men_men_n237_), .B0(x2), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n263_), .B(men_men_n174_), .Y(men_men_n264_));
  NAi21      u248(.An(x4), .B(x0), .Y(men_men_n265_));
  NO3        u249(.A(men_men_n265_), .B(men_men_n39_), .C(x2), .Y(men_men_n266_));
  OAI210     u250(.A0(x6), .A1(men_men_n18_), .B0(men_men_n266_), .Y(men_men_n267_));
  OAI220     u251(.A0(men_men_n22_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n268_));
  NO2        u252(.A(x9), .B(x8), .Y(men_men_n269_));
  NA3        u253(.A(men_men_n269_), .B(men_men_n34_), .C(men_men_n47_), .Y(men_men_n270_));
  INV        u254(.A(men_men_n270_), .Y(men_men_n271_));
  AOI220     u255(.A0(men_men_n271_), .A1(men_men_n72_), .B0(men_men_n268_), .B1(men_men_n29_), .Y(men_men_n272_));
  AOI210     u256(.A0(men_men_n272_), .A1(men_men_n267_), .B0(men_men_n23_), .Y(men_men_n273_));
  NA2        u257(.A(men_men_n34_), .B(men_men_n38_), .Y(men_men_n274_));
  OR2        u258(.A(men_men_n274_), .B(men_men_n254_), .Y(men_men_n275_));
  NO2        u259(.A(men_men_n275_), .B(men_men_n148_), .Y(men_men_n276_));
  NO3        u260(.A(men_men_n276_), .B(men_men_n273_), .C(men_men_n264_), .Y(men_men_n277_));
  OAI210     u261(.A0(men_men_n262_), .A1(men_men_n226_), .B0(men_men_n277_), .Y(men04));
  OAI210     u262(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n279_));
  NA3        u263(.A(men_men_n279_), .B(men_men_n250_), .C(men_men_n75_), .Y(men_men_n280_));
  AOI210     u264(.A0(men_men_n55_), .A1(x4), .B0(x0), .Y(men_men_n281_));
  OAI210     u265(.A0(men_men_n281_), .A1(x1), .B0(men_men_n227_), .Y(men_men_n282_));
  NO2        u266(.A(men_men_n248_), .B(men_men_n82_), .Y(men_men_n283_));
  NO2        u267(.A(men_men_n283_), .B(men_men_n34_), .Y(men_men_n284_));
  NA2        u268(.A(x9), .B(men_men_n84_), .Y(men_men_n285_));
  NA3        u269(.A(men_men_n285_), .B(men_men_n284_), .C(men_men_n282_), .Y(men_men_n286_));
  NA2        u270(.A(men_men_n286_), .B(x6), .Y(men_men_n287_));
  NO2        u271(.A(x2), .B(men_men_n18_), .Y(men_men_n288_));
  NO2        u272(.A(men_men_n288_), .B(x0), .Y(men_men_n289_));
  NA2        u273(.A(men_men_n138_), .B(men_men_n56_), .Y(men_men_n290_));
  NA3        u274(.A(x8), .B(men_men_n290_), .C(men_men_n289_), .Y(men_men_n291_));
  OAI210     u275(.A0(men_men_n100_), .A1(x3), .B0(men_men_n266_), .Y(men_men_n292_));
  NA3        u276(.A(men_men_n208_), .B(men_men_n195_), .C(men_men_n74_), .Y(men_men_n293_));
  NA3        u277(.A(men_men_n293_), .B(men_men_n292_), .C(men_men_n140_), .Y(men_men_n294_));
  AOI210     u278(.A0(men_men_n291_), .A1(x4), .B0(men_men_n294_), .Y(men_men_n295_));
  NOi21      u279(.An(x4), .B(x0), .Y(men_men_n296_));
  XO2        u280(.A(x4), .B(x0), .Y(men_men_n297_));
  OAI210     u281(.A0(men_men_n297_), .A1(men_men_n105_), .B0(men_men_n244_), .Y(men_men_n298_));
  AOI220     u282(.A0(men_men_n298_), .A1(x8), .B0(men_men_n296_), .B1(men_men_n85_), .Y(men_men_n299_));
  NO2        u283(.A(men_men_n299_), .B(x3), .Y(men_men_n300_));
  INV        u284(.A(men_men_n85_), .Y(men_men_n301_));
  NO2        u285(.A(men_men_n84_), .B(x4), .Y(men_men_n302_));
  AOI220     u286(.A0(men_men_n302_), .A1(men_men_n39_), .B0(men_men_n113_), .B1(men_men_n301_), .Y(men_men_n303_));
  NO3        u287(.A(men_men_n297_), .B(men_men_n151_), .C(x2), .Y(men_men_n304_));
  NO2        u288(.A(men_men_n26_), .B(men_men_n22_), .Y(men_men_n305_));
  NO2        u289(.A(men_men_n305_), .B(men_men_n304_), .Y(men_men_n306_));
  NA4        u290(.A(men_men_n306_), .B(men_men_n303_), .C(men_men_n204_), .D(x6), .Y(men_men_n307_));
  OAI220     u291(.A0(men_men_n265_), .A1(men_men_n82_), .B0(men_men_n169_), .B1(men_men_n84_), .Y(men_men_n308_));
  NO2        u292(.A(men_men_n38_), .B(x0), .Y(men_men_n309_));
  OR2        u293(.A(men_men_n302_), .B(men_men_n309_), .Y(men_men_n310_));
  NO2        u294(.A(men_men_n138_), .B(men_men_n96_), .Y(men_men_n311_));
  AOI220     u295(.A0(men_men_n311_), .A1(men_men_n310_), .B0(men_men_n308_), .B1(men_men_n54_), .Y(men_men_n312_));
  NOi21      u296(.An(men_men_n109_), .B(men_men_n25_), .Y(men_men_n313_));
  INV        u297(.A(men_men_n313_), .Y(men_men_n314_));
  OAI210     u298(.A0(men_men_n312_), .A1(men_men_n55_), .B0(men_men_n314_), .Y(men_men_n315_));
  OAI220     u299(.A0(men_men_n315_), .A1(x6), .B0(men_men_n307_), .B1(men_men_n300_), .Y(men_men_n316_));
  OAI210     u300(.A0(men_men_n56_), .A1(men_men_n42_), .B0(men_men_n37_), .Y(men_men_n317_));
  OAI210     u301(.A0(men_men_n317_), .A1(men_men_n84_), .B0(men_men_n275_), .Y(men_men_n318_));
  AOI210     u302(.A0(men_men_n318_), .A1(men_men_n18_), .B0(men_men_n140_), .Y(men_men_n319_));
  AO220      u303(.A0(men_men_n319_), .A1(men_men_n316_), .B0(men_men_n295_), .B1(men_men_n287_), .Y(men_men_n320_));
  NA2        u304(.A(men_men_n320_), .B(men_men_n280_), .Y(men_men_n321_));
  AOI210     u305(.A0(men_men_n180_), .A1(x8), .B0(men_men_n100_), .Y(men_men_n322_));
  INV        u306(.A(men_men_n322_), .Y(men_men_n323_));
  NA3        u307(.A(men_men_n323_), .B(men_men_n179_), .C(men_men_n140_), .Y(men_men_n324_));
  NA3        u308(.A(x7), .B(x3), .C(x0), .Y(men_men_n325_));
  NO2        u309(.A(men_men_n325_), .B(men_men_n301_), .Y(men_men_n326_));
  AOI210     u310(.A0(x4), .A1(men_men_n107_), .B0(men_men_n326_), .Y(men_men_n327_));
  AOI210     u311(.A0(men_men_n327_), .A1(men_men_n324_), .B0(men_men_n23_), .Y(men_men_n328_));
  NA3        u312(.A(men_men_n108_), .B(men_men_n203_), .C(x0), .Y(men_men_n329_));
  NA3        u313(.A(men_men_n180_), .B(men_men_n205_), .C(x8), .Y(men_men_n330_));
  AOI210     u314(.A0(men_men_n330_), .A1(x0), .B0(men_men_n23_), .Y(men_men_n331_));
  AOI210     u315(.A0(x2), .A1(men_men_n106_), .B0(men_men_n37_), .Y(men_men_n332_));
  NOi21      u316(.An(men_men_n332_), .B(men_men_n170_), .Y(men_men_n333_));
  OAI210     u317(.A0(men_men_n333_), .A1(men_men_n331_), .B0(men_men_n137_), .Y(men_men_n334_));
  NA2        u318(.A(men_men_n334_), .B(men_men_n329_), .Y(men_men_n335_));
  OAI210     u319(.A0(men_men_n335_), .A1(men_men_n328_), .B0(x6), .Y(men_men_n336_));
  OAI210     u320(.A0(men_men_n151_), .A1(men_men_n42_), .B0(men_men_n122_), .Y(men_men_n337_));
  NA3        u321(.A(men_men_n48_), .B(x7), .C(men_men_n29_), .Y(men_men_n338_));
  AOI220     u322(.A0(men_men_n338_), .A1(men_men_n337_), .B0(men_men_n35_), .B1(men_men_n30_), .Y(men_men_n339_));
  NA2        u323(.A(men_men_n179_), .B(men_men_n140_), .Y(men_men_n340_));
  OAI210     u324(.A0(men_men_n340_), .A1(x8), .B0(men_men_n393_), .Y(men_men_n341_));
  NAi31      u325(.An(x2), .B(x8), .C(x0), .Y(men_men_n342_));
  OAI210     u326(.A0(men_men_n342_), .A1(x4), .B0(men_men_n152_), .Y(men_men_n343_));
  NA3        u327(.A(men_men_n343_), .B(men_men_n135_), .C(x9), .Y(men_men_n344_));
  NO4        u328(.A(men_men_n114_), .B(men_men_n265_), .C(x9), .D(x2), .Y(men_men_n345_));
  NOi21      u329(.An(men_men_n112_), .B(men_men_n169_), .Y(men_men_n346_));
  NO3        u330(.A(men_men_n346_), .B(men_men_n345_), .C(men_men_n18_), .Y(men_men_n347_));
  NO3        u331(.A(x9), .B(men_men_n140_), .C(x0), .Y(men_men_n348_));
  NA2        u332(.A(men_men_n348_), .B(men_men_n227_), .Y(men_men_n349_));
  NA4        u333(.A(men_men_n349_), .B(men_men_n347_), .C(men_men_n344_), .D(men_men_n44_), .Y(men_men_n350_));
  OAI210     u334(.A0(men_men_n341_), .A1(men_men_n339_), .B0(men_men_n350_), .Y(men_men_n351_));
  NO2        u335(.A(men_men_n112_), .B(men_men_n38_), .Y(men_men_n352_));
  AOI220     u336(.A0(x1), .A1(men_men_n296_), .B0(men_men_n113_), .B1(x3), .Y(men_men_n353_));
  AOI210     u337(.A0(men_men_n244_), .A1(men_men_n53_), .B0(men_men_n111_), .Y(men_men_n354_));
  OAI210     u338(.A0(men_men_n354_), .A1(x3), .B0(men_men_n353_), .Y(men_men_n355_));
  NO3        u339(.A(men_men_n355_), .B(men_men_n352_), .C(x2), .Y(men_men_n356_));
  OAI220     u340(.A0(men_men_n297_), .A1(men_men_n269_), .B0(men_men_n265_), .B1(men_men_n38_), .Y(men_men_n357_));
  AOI210     u341(.A0(x9), .A1(men_men_n42_), .B0(men_men_n325_), .Y(men_men_n358_));
  AOI220     u342(.A0(men_men_n358_), .A1(men_men_n84_), .B0(men_men_n357_), .B1(men_men_n140_), .Y(men_men_n359_));
  NO2        u343(.A(men_men_n359_), .B(men_men_n47_), .Y(men_men_n360_));
  NO2        u344(.A(men_men_n360_), .B(men_men_n356_), .Y(men_men_n361_));
  AOI210     u345(.A0(men_men_n361_), .A1(men_men_n351_), .B0(men_men_n23_), .Y(men_men_n362_));
  NA4        u346(.A(men_men_n29_), .B(men_men_n84_), .C(x2), .D(men_men_n17_), .Y(men_men_n363_));
  NO3        u347(.A(men_men_n55_), .B(x4), .C(x1), .Y(men_men_n364_));
  NO3        u348(.A(men_men_n61_), .B(men_men_n18_), .C(x0), .Y(men_men_n365_));
  AOI220     u349(.A0(men_men_n365_), .A1(x4), .B0(men_men_n364_), .B1(men_men_n332_), .Y(men_men_n366_));
  NO2        u350(.A(men_men_n366_), .B(men_men_n93_), .Y(men_men_n367_));
  NO3        u351(.A(men_men_n248_), .B(men_men_n164_), .C(men_men_n35_), .Y(men_men_n368_));
  OAI210     u352(.A0(men_men_n368_), .A1(men_men_n367_), .B0(x7), .Y(men_men_n369_));
  NA2        u353(.A(men_men_n208_), .B(x7), .Y(men_men_n370_));
  NA3        u354(.A(men_men_n370_), .B(men_men_n139_), .C(men_men_n121_), .Y(men_men_n371_));
  NA3        u355(.A(men_men_n371_), .B(men_men_n369_), .C(men_men_n363_), .Y(men_men_n372_));
  OAI210     u356(.A0(men_men_n372_), .A1(men_men_n362_), .B0(men_men_n34_), .Y(men_men_n373_));
  NO2        u357(.A(men_men_n348_), .B(men_men_n187_), .Y(men_men_n374_));
  NO4        u358(.A(men_men_n374_), .B(men_men_n68_), .C(x4), .D(men_men_n47_), .Y(men_men_n375_));
  NO2        u359(.A(men_men_n155_), .B(men_men_n26_), .Y(men_men_n376_));
  AOI220     u360(.A0(men_men_n309_), .A1(men_men_n84_), .B0(men_men_n138_), .B1(men_men_n180_), .Y(men_men_n377_));
  NA3        u361(.A(men_men_n377_), .B(men_men_n342_), .C(men_men_n82_), .Y(men_men_n378_));
  NA2        u362(.A(men_men_n378_), .B(men_men_n165_), .Y(men_men_n379_));
  NA2        u363(.A(x3), .B(men_men_n47_), .Y(men_men_n380_));
  AOI210     u364(.A0(men_men_n152_), .A1(men_men_n25_), .B0(men_men_n63_), .Y(men_men_n381_));
  INV        u365(.A(men_men_n381_), .Y(men_men_n382_));
  OAI210     u366(.A0(men_men_n141_), .A1(men_men_n380_), .B0(men_men_n382_), .Y(men_men_n383_));
  NA2        u367(.A(men_men_n383_), .B(x0), .Y(men_men_n384_));
  AOI210     u368(.A0(men_men_n384_), .A1(men_men_n379_), .B0(men_men_n215_), .Y(men_men_n385_));
  NA2        u369(.A(x9), .B(x5), .Y(men_men_n386_));
  NO4        u370(.A(men_men_n96_), .B(men_men_n386_), .C(men_men_n53_), .D(men_men_n30_), .Y(men_men_n387_));
  NO4        u371(.A(men_men_n387_), .B(men_men_n385_), .C(men_men_n376_), .D(men_men_n375_), .Y(men_men_n388_));
  NA3        u372(.A(men_men_n388_), .B(men_men_n373_), .C(men_men_n336_), .Y(men_men_n389_));
  AOI210     u373(.A0(men_men_n321_), .A1(men_men_n23_), .B0(men_men_n389_), .Y(men05));
  INV        u374(.A(x1), .Y(men_men_n393_));
  INV        u375(.A(x6), .Y(men_men_n394_));
  INV        u376(.A(x4), .Y(men_men_n395_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule