// Benchmark "top" written by ABC on Thu Jun 20 14:59:19 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n140_, new_new_n141_, new_new_n142_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1057_, new_new_n1058_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  OAI210     g0067(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n89_), .Y(new_new_n90_));
  NAi21      g0068(.An(i_6_), .B(i_10_), .Y(new_new_n91_));
  NA2        g0069(.A(i_6_), .B(i_9_), .Y(new_new_n92_));
  AOI210     g0070(.A0(new_new_n92_), .A1(new_new_n91_), .B0(new_new_n64_), .Y(new_new_n93_));
  NA2        g0071(.A(i_2_), .B(i_6_), .Y(new_new_n94_));
  NO3        g0072(.A(new_new_n94_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n95_));
  NO2        g0073(.A(new_new_n95_), .B(new_new_n93_), .Y(new_new_n96_));
  AOI210     g0074(.A0(new_new_n96_), .A1(new_new_n90_), .B0(new_new_n81_), .Y(new_new_n97_));
  AN3        g0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n98_));
  NAi21      g0076(.An(i_6_), .B(i_11_), .Y(new_new_n99_));
  NO2        g0077(.A(i_5_), .B(i_8_), .Y(new_new_n100_));
  NOi21      g0078(.An(new_new_n100_), .B(new_new_n99_), .Y(new_new_n101_));
  AOI220     g0079(.A0(new_new_n101_), .A1(new_new_n63_), .B0(new_new_n98_), .B1(new_new_n32_), .Y(new_new_n102_));
  INV        g0080(.A(i_7_), .Y(new_new_n103_));
  NA2        g0081(.A(new_new_n47_), .B(new_new_n103_), .Y(new_new_n104_));
  NO2        g0082(.A(i_0_), .B(i_5_), .Y(new_new_n105_));
  NO2        g0083(.A(new_new_n105_), .B(new_new_n87_), .Y(new_new_n106_));
  NA2        g0084(.A(i_12_), .B(i_3_), .Y(new_new_n107_));
  INV        g0085(.A(new_new_n107_), .Y(new_new_n108_));
  NA3        g0086(.A(new_new_n108_), .B(new_new_n106_), .C(new_new_n104_), .Y(new_new_n109_));
  NAi21      g0087(.An(i_7_), .B(i_11_), .Y(new_new_n110_));
  AN2        g0088(.A(i_2_), .B(i_10_), .Y(new_new_n111_));
  NO2        g0089(.A(new_new_n111_), .B(i_7_), .Y(new_new_n112_));
  OR2        g0090(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n113_));
  NO2        g0091(.A(i_8_), .B(new_new_n103_), .Y(new_new_n114_));
  NO3        g0092(.A(new_new_n114_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n115_));
  NA2        g0093(.A(i_12_), .B(i_7_), .Y(new_new_n116_));
  NO2        g0094(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n117_));
  NA2        g0095(.A(new_new_n117_), .B(i_0_), .Y(new_new_n118_));
  NA2        g0096(.A(i_11_), .B(i_12_), .Y(new_new_n119_));
  OAI210     g0097(.A0(new_new_n118_), .A1(new_new_n116_), .B0(new_new_n119_), .Y(new_new_n120_));
  NO2        g0098(.A(new_new_n120_), .B(new_new_n115_), .Y(new_new_n121_));
  NA3        g0099(.A(new_new_n121_), .B(new_new_n109_), .C(new_new_n102_), .Y(new_new_n122_));
  NOi21      g0100(.An(i_1_), .B(i_5_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n123_), .B(i_11_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n125_));
  NA2        g0103(.A(i_7_), .B(new_new_n25_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NO2        g0105(.A(new_new_n127_), .B(new_new_n47_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n92_), .B(new_new_n91_), .Y(new_new_n129_));
  NAi21      g0107(.An(i_3_), .B(i_8_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n130_), .B(new_new_n63_), .Y(new_new_n131_));
  NOi31      g0109(.An(new_new_n131_), .B(new_new_n129_), .C(new_new_n128_), .Y(new_new_n132_));
  NO2        g0110(.A(i_1_), .B(new_new_n87_), .Y(new_new_n133_));
  NO2        g0111(.A(i_6_), .B(i_5_), .Y(new_new_n134_));
  NA2        g0112(.A(new_new_n134_), .B(i_3_), .Y(new_new_n135_));
  AO210      g0113(.A0(new_new_n135_), .A1(new_new_n48_), .B0(new_new_n133_), .Y(new_new_n136_));
  OAI220     g0114(.A0(new_new_n136_), .A1(new_new_n110_), .B0(new_new_n132_), .B1(new_new_n124_), .Y(new_new_n137_));
  NO3        g0115(.A(new_new_n137_), .B(new_new_n122_), .C(new_new_n97_), .Y(new_new_n138_));
  NA3        g0116(.A(new_new_n138_), .B(new_new_n80_), .C(new_new_n57_), .Y(men2));
  NO2        g0117(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n140_));
  NA2        g0118(.A(i_6_), .B(new_new_n25_), .Y(new_new_n141_));
  NA2        g0119(.A(new_new_n141_), .B(new_new_n140_), .Y(new_new_n142_));
  NA4        g0120(.A(new_new_n142_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(men0));
  AN2        g0121(.A(i_8_), .B(i_7_), .Y(new_new_n144_));
  NA2        g0122(.A(new_new_n144_), .B(i_6_), .Y(new_new_n145_));
  NO2        g0123(.A(i_12_), .B(i_13_), .Y(new_new_n146_));
  NAi21      g0124(.An(i_5_), .B(i_11_), .Y(new_new_n147_));
  NOi21      g0125(.An(new_new_n146_), .B(new_new_n147_), .Y(new_new_n148_));
  NO2        g0126(.A(i_0_), .B(i_1_), .Y(new_new_n149_));
  NA2        g0127(.A(i_2_), .B(i_3_), .Y(new_new_n150_));
  NO2        g0128(.A(new_new_n150_), .B(i_4_), .Y(new_new_n151_));
  NA3        g0129(.A(new_new_n151_), .B(new_new_n149_), .C(new_new_n148_), .Y(new_new_n152_));
  AN2        g0130(.A(new_new_n146_), .B(new_new_n84_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(new_new_n27_), .Y(new_new_n154_));
  NA2        g0132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n156_));
  NA2        g0134(.A(new_new_n156_), .B(new_new_n36_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n158_));
  OR2        g0136(.A(i_0_), .B(i_1_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n160_));
  NAi32      g0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n161_));
  NAi21      g0139(.An(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NOi21      g0140(.An(i_4_), .B(i_10_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n40_), .Y(new_new_n164_));
  NO2        g0142(.A(i_3_), .B(i_5_), .Y(new_new_n165_));
  NO3        g0143(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  OAI210     g0145(.A0(new_new_n167_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n168_));
  NO2        g0146(.A(new_new_n168_), .B(new_new_n158_), .Y(new_new_n169_));
  AOI210     g0147(.A0(new_new_n169_), .A1(new_new_n152_), .B0(new_new_n145_), .Y(new_new_n170_));
  NA3        g0148(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n171_));
  NA2        g0149(.A(i_3_), .B(new_new_n49_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_4_), .B(i_9_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_11_), .B(i_13_), .Y(new_new_n174_));
  NA2        g0152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  OR2        g0153(.A(new_new_n175_), .B(new_new_n172_), .Y(new_new_n176_));
  NO2        g0154(.A(i_4_), .B(i_5_), .Y(new_new_n177_));
  NAi21      g0155(.An(i_12_), .B(i_11_), .Y(new_new_n178_));
  NO2        g0156(.A(new_new_n178_), .B(i_13_), .Y(new_new_n179_));
  NA3        g0157(.A(new_new_n179_), .B(new_new_n177_), .C(new_new_n84_), .Y(new_new_n180_));
  AOI210     g0158(.A0(new_new_n180_), .A1(new_new_n176_), .B0(new_new_n171_), .Y(new_new_n181_));
  NO2        g0159(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n36_), .B(i_5_), .Y(new_new_n183_));
  NA2        g0161(.A(i_3_), .B(i_5_), .Y(new_new_n184_));
  NO2        g0162(.A(new_new_n74_), .B(i_5_), .Y(new_new_n185_));
  NO2        g0163(.A(i_13_), .B(i_10_), .Y(new_new_n186_));
  NA3        g0164(.A(new_new_n186_), .B(new_new_n185_), .C(new_new_n45_), .Y(new_new_n187_));
  NO2        g0165(.A(i_2_), .B(i_1_), .Y(new_new_n188_));
  NA2        g0166(.A(new_new_n188_), .B(i_3_), .Y(new_new_n189_));
  NAi21      g0167(.An(i_4_), .B(i_12_), .Y(new_new_n190_));
  NO4        g0168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n187_), .D(new_new_n25_), .Y(new_new_n191_));
  NO2        g0169(.A(new_new_n191_), .B(new_new_n181_), .Y(new_new_n192_));
  INV        g0170(.A(i_8_), .Y(new_new_n193_));
  NO2        g0171(.A(new_new_n193_), .B(i_7_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(i_6_), .Y(new_new_n195_));
  NO3        g0173(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(new_new_n114_), .Y(new_new_n197_));
  NO3        g0175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n198_));
  NA3        g0176(.A(new_new_n198_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n199_));
  NO3        g0177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n200_));
  OAI210     g0178(.A0(new_new_n98_), .A1(i_12_), .B0(new_new_n200_), .Y(new_new_n201_));
  AOI210     g0179(.A0(new_new_n201_), .A1(new_new_n199_), .B0(new_new_n197_), .Y(new_new_n202_));
  NO2        g0180(.A(i_3_), .B(i_8_), .Y(new_new_n203_));
  NO3        g0181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(new_new_n203_), .C(new_new_n40_), .Y(new_new_n205_));
  NO2        g0183(.A(new_new_n105_), .B(new_new_n59_), .Y(new_new_n206_));
  INV        g0184(.A(new_new_n206_), .Y(new_new_n207_));
  NO2        g0185(.A(i_13_), .B(i_9_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(i_6_), .C(new_new_n193_), .Y(new_new_n209_));
  NAi21      g0187(.An(i_12_), .B(i_3_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n45_), .B(i_5_), .Y(new_new_n211_));
  NO3        g0189(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n212_));
  NA3        g0190(.A(new_new_n212_), .B(new_new_n211_), .C(i_10_), .Y(new_new_n213_));
  OAI220     g0191(.A0(new_new_n213_), .A1(new_new_n209_), .B0(new_new_n207_), .B1(new_new_n205_), .Y(new_new_n214_));
  AOI210     g0192(.A0(new_new_n214_), .A1(i_7_), .B0(new_new_n202_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(i_4_), .B0(new_new_n195_), .B1(new_new_n192_), .Y(new_new_n216_));
  NAi21      g0194(.An(i_12_), .B(i_7_), .Y(new_new_n217_));
  NA3        g0195(.A(i_13_), .B(new_new_n193_), .C(i_10_), .Y(new_new_n218_));
  NA2        g0196(.A(i_0_), .B(i_5_), .Y(new_new_n219_));
  NAi31      g0197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n36_), .B(i_13_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n223_));
  NA3        g0201(.A(new_new_n223_), .B(new_new_n222_), .C(new_new_n221_), .Y(new_new_n224_));
  INV        g0202(.A(i_13_), .Y(new_new_n225_));
  NO2        g0203(.A(i_12_), .B(new_new_n225_), .Y(new_new_n226_));
  NA3        g0204(.A(new_new_n226_), .B(new_new_n198_), .C(new_new_n196_), .Y(new_new_n227_));
  OAI210     g0205(.A0(new_new_n224_), .A1(new_new_n220_), .B0(new_new_n227_), .Y(new_new_n228_));
  NA2        g0206(.A(new_new_n228_), .B(new_new_n144_), .Y(new_new_n229_));
  NO2        g0207(.A(i_12_), .B(new_new_n37_), .Y(new_new_n230_));
  NO2        g0208(.A(new_new_n184_), .B(i_4_), .Y(new_new_n231_));
  NA2        g0209(.A(new_new_n231_), .B(new_new_n230_), .Y(new_new_n232_));
  OR2        g0210(.A(i_8_), .B(i_7_), .Y(new_new_n233_));
  NO2        g0211(.A(new_new_n233_), .B(new_new_n87_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n54_), .B(i_1_), .Y(new_new_n235_));
  INV        g0213(.A(i_12_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n45_), .B(new_new_n236_), .Y(new_new_n237_));
  NO3        g0215(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n238_));
  NA2        g0216(.A(i_2_), .B(i_1_), .Y(new_new_n239_));
  NO3        g0217(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n240_));
  NAi21      g0218(.An(i_4_), .B(i_3_), .Y(new_new_n241_));
  NO2        g0219(.A(i_0_), .B(i_6_), .Y(new_new_n242_));
  NOi41      g0220(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(new_new_n243_), .B(new_new_n242_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n239_), .B(new_new_n184_), .Y(new_new_n245_));
  NAi21      g0223(.An(new_new_n244_), .B(new_new_n245_), .Y(new_new_n246_));
  INV        g0224(.A(new_new_n246_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n247_), .B(new_new_n40_), .Y(new_new_n248_));
  NO2        g0226(.A(i_11_), .B(new_new_n225_), .Y(new_new_n249_));
  NOi21      g0227(.An(i_1_), .B(i_6_), .Y(new_new_n250_));
  NAi21      g0228(.An(i_3_), .B(i_7_), .Y(new_new_n251_));
  NA2        g0229(.A(new_new_n236_), .B(i_9_), .Y(new_new_n252_));
  OR4        g0230(.A(new_new_n252_), .B(new_new_n251_), .C(new_new_n250_), .D(new_new_n185_), .Y(new_new_n253_));
  NO2        g0231(.A(i_12_), .B(i_3_), .Y(new_new_n254_));
  NA2        g0232(.A(new_new_n74_), .B(i_5_), .Y(new_new_n255_));
  NA2        g0233(.A(i_3_), .B(i_9_), .Y(new_new_n256_));
  NAi21      g0234(.An(i_7_), .B(i_10_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n257_), .B(new_new_n256_), .Y(new_new_n258_));
  NA3        g0236(.A(new_new_n258_), .B(new_new_n255_), .C(new_new_n65_), .Y(new_new_n259_));
  NA2        g0237(.A(new_new_n259_), .B(new_new_n253_), .Y(new_new_n260_));
  NA3        g0238(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n261_));
  INV        g0239(.A(new_new_n145_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n236_), .B(i_13_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n263_), .B(new_new_n76_), .Y(new_new_n264_));
  AOI220     g0242(.A0(new_new_n264_), .A1(new_new_n262_), .B0(new_new_n260_), .B1(new_new_n249_), .Y(new_new_n265_));
  NA2        g0243(.A(i_12_), .B(i_6_), .Y(new_new_n266_));
  OR2        g0244(.A(i_13_), .B(i_9_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n241_), .B(i_2_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n249_), .B(i_9_), .Y(new_new_n269_));
  NO3        g0247(.A(i_11_), .B(new_new_n225_), .C(new_new_n25_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n251_), .B(i_8_), .Y(new_new_n271_));
  NO2        g0249(.A(i_6_), .B(new_new_n49_), .Y(new_new_n272_));
  NA3        g0250(.A(new_new_n265_), .B(new_new_n248_), .C(new_new_n229_), .Y(new_new_n273_));
  NO3        g0251(.A(i_12_), .B(new_new_n225_), .C(new_new_n37_), .Y(new_new_n274_));
  INV        g0252(.A(new_new_n274_), .Y(new_new_n275_));
  NO3        g0253(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n276_));
  NO3        g0254(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n277_));
  NO2        g0255(.A(new_new_n239_), .B(i_0_), .Y(new_new_n278_));
  AOI220     g0256(.A0(new_new_n278_), .A1(new_new_n194_), .B0(new_new_n277_), .B1(new_new_n144_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n272_), .B(new_new_n26_), .Y(new_new_n280_));
  NO2        g0258(.A(new_new_n280_), .B(new_new_n279_), .Y(new_new_n281_));
  NA2        g0259(.A(i_0_), .B(i_1_), .Y(new_new_n282_));
  NO2        g0260(.A(new_new_n282_), .B(i_2_), .Y(new_new_n283_));
  NO2        g0261(.A(new_new_n60_), .B(i_6_), .Y(new_new_n284_));
  NA3        g0262(.A(new_new_n284_), .B(new_new_n283_), .C(new_new_n165_), .Y(new_new_n285_));
  OAI210     g0263(.A0(new_new_n167_), .A1(new_new_n145_), .B0(new_new_n285_), .Y(new_new_n286_));
  NO2        g0264(.A(new_new_n286_), .B(new_new_n281_), .Y(new_new_n287_));
  NO2        g0265(.A(i_3_), .B(i_10_), .Y(new_new_n288_));
  NA3        g0266(.A(new_new_n288_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n289_));
  NO2        g0267(.A(i_2_), .B(new_new_n103_), .Y(new_new_n290_));
  NA2        g0268(.A(i_1_), .B(new_new_n36_), .Y(new_new_n291_));
  NO2        g0269(.A(new_new_n291_), .B(i_8_), .Y(new_new_n292_));
  NA2        g0270(.A(new_new_n292_), .B(new_new_n290_), .Y(new_new_n293_));
  AN2        g0271(.A(i_3_), .B(i_10_), .Y(new_new_n294_));
  NA4        g0272(.A(new_new_n294_), .B(new_new_n198_), .C(new_new_n179_), .D(new_new_n177_), .Y(new_new_n295_));
  NO2        g0273(.A(i_5_), .B(new_new_n37_), .Y(new_new_n296_));
  NO2        g0274(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n297_));
  OR2        g0275(.A(new_new_n293_), .B(new_new_n289_), .Y(new_new_n298_));
  OAI220     g0276(.A0(new_new_n298_), .A1(i_6_), .B0(new_new_n287_), .B1(new_new_n275_), .Y(new_new_n299_));
  NO4        g0277(.A(new_new_n299_), .B(new_new_n273_), .C(new_new_n216_), .D(new_new_n170_), .Y(new_new_n300_));
  NO3        g0278(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n302_));
  NA2        g0280(.A(new_new_n278_), .B(new_new_n302_), .Y(new_new_n303_));
  NO3        g0281(.A(i_6_), .B(new_new_n193_), .C(i_7_), .Y(new_new_n304_));
  NA2        g0282(.A(new_new_n304_), .B(new_new_n198_), .Y(new_new_n305_));
  AOI210     g0283(.A0(new_new_n305_), .A1(new_new_n303_), .B0(new_new_n172_), .Y(new_new_n306_));
  NO2        g0284(.A(i_2_), .B(i_3_), .Y(new_new_n307_));
  OR2        g0285(.A(i_0_), .B(i_5_), .Y(new_new_n308_));
  NA2        g0286(.A(new_new_n219_), .B(new_new_n308_), .Y(new_new_n309_));
  NAi21      g0287(.An(i_8_), .B(i_7_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n310_), .B(i_6_), .Y(new_new_n311_));
  NO2        g0289(.A(new_new_n159_), .B(new_new_n47_), .Y(new_new_n312_));
  NA3        g0290(.A(new_new_n312_), .B(new_new_n311_), .C(new_new_n165_), .Y(new_new_n313_));
  INV        g0291(.A(new_new_n313_), .Y(new_new_n314_));
  OAI210     g0292(.A0(new_new_n314_), .A1(new_new_n306_), .B0(i_4_), .Y(new_new_n315_));
  NO2        g0293(.A(i_12_), .B(i_10_), .Y(new_new_n316_));
  NOi21      g0294(.An(i_5_), .B(i_0_), .Y(new_new_n317_));
  AOI210     g0295(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n103_), .Y(new_new_n318_));
  NO4        g0296(.A(new_new_n318_), .B(new_new_n291_), .C(new_new_n317_), .D(new_new_n130_), .Y(new_new_n319_));
  NA4        g0297(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n319_), .B(new_new_n316_), .Y(new_new_n321_));
  NO2        g0299(.A(i_6_), .B(i_8_), .Y(new_new_n322_));
  NOi21      g0300(.An(i_0_), .B(i_2_), .Y(new_new_n323_));
  AN2        g0301(.A(new_new_n323_), .B(new_new_n322_), .Y(new_new_n324_));
  NO2        g0302(.A(i_1_), .B(i_7_), .Y(new_new_n325_));
  AO220      g0303(.A0(new_new_n325_), .A1(new_new_n324_), .B0(new_new_n311_), .B1(new_new_n235_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n327_));
  NA3        g0305(.A(new_new_n327_), .B(new_new_n321_), .C(new_new_n315_), .Y(new_new_n328_));
  NA3        g0306(.A(new_new_n250_), .B(new_new_n290_), .C(new_new_n193_), .Y(new_new_n329_));
  NO2        g0307(.A(new_new_n329_), .B(new_new_n309_), .Y(new_new_n330_));
  NOi21      g0308(.An(new_new_n155_), .B(new_new_n106_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n331_), .B(new_new_n126_), .Y(new_new_n332_));
  OAI210     g0310(.A0(new_new_n332_), .A1(new_new_n330_), .B0(i_3_), .Y(new_new_n333_));
  INV        g0311(.A(new_new_n85_), .Y(new_new_n334_));
  NO2        g0312(.A(new_new_n282_), .B(new_new_n82_), .Y(new_new_n335_));
  NA2        g0313(.A(new_new_n335_), .B(new_new_n134_), .Y(new_new_n336_));
  NO2        g0314(.A(new_new_n94_), .B(new_new_n193_), .Y(new_new_n337_));
  NA3        g0315(.A(new_new_n219_), .B(new_new_n337_), .C(new_new_n64_), .Y(new_new_n338_));
  AOI210     g0316(.A0(new_new_n338_), .A1(new_new_n336_), .B0(new_new_n334_), .Y(new_new_n339_));
  NO2        g0317(.A(new_new_n193_), .B(i_9_), .Y(new_new_n340_));
  NA2        g0318(.A(new_new_n340_), .B(new_new_n206_), .Y(new_new_n341_));
  NO2        g0319(.A(new_new_n341_), .B(new_new_n47_), .Y(new_new_n342_));
  NO3        g0320(.A(new_new_n342_), .B(new_new_n339_), .C(new_new_n281_), .Y(new_new_n343_));
  AOI210     g0321(.A0(new_new_n343_), .A1(new_new_n333_), .B0(new_new_n164_), .Y(new_new_n344_));
  AOI210     g0322(.A0(new_new_n328_), .A1(new_new_n301_), .B0(new_new_n344_), .Y(new_new_n345_));
  NOi32      g0323(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n346_));
  INV        g0324(.A(new_new_n346_), .Y(new_new_n347_));
  NAi21      g0325(.An(i_0_), .B(i_6_), .Y(new_new_n348_));
  NAi21      g0326(.An(i_1_), .B(i_5_), .Y(new_new_n349_));
  NA2        g0327(.A(new_new_n349_), .B(new_new_n348_), .Y(new_new_n350_));
  NA2        g0328(.A(new_new_n350_), .B(new_new_n25_), .Y(new_new_n351_));
  OAI210     g0329(.A0(new_new_n351_), .A1(new_new_n161_), .B0(new_new_n244_), .Y(new_new_n352_));
  NAi41      g0330(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n353_));
  OAI220     g0331(.A0(new_new_n353_), .A1(new_new_n349_), .B0(new_new_n220_), .B1(new_new_n161_), .Y(new_new_n354_));
  AOI210     g0332(.A0(new_new_n353_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n355_));
  NOi32      g0333(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n356_));
  NAi21      g0334(.An(i_6_), .B(i_1_), .Y(new_new_n357_));
  NA3        g0335(.A(new_new_n357_), .B(new_new_n356_), .C(new_new_n47_), .Y(new_new_n358_));
  NO2        g0336(.A(new_new_n358_), .B(i_0_), .Y(new_new_n359_));
  OR3        g0337(.A(new_new_n359_), .B(new_new_n355_), .C(new_new_n354_), .Y(new_new_n360_));
  NO2        g0338(.A(i_1_), .B(new_new_n103_), .Y(new_new_n361_));
  NAi21      g0339(.An(i_3_), .B(i_4_), .Y(new_new_n362_));
  NO2        g0340(.A(new_new_n362_), .B(i_9_), .Y(new_new_n363_));
  AN2        g0341(.A(i_6_), .B(i_7_), .Y(new_new_n364_));
  OAI210     g0342(.A0(new_new_n364_), .A1(new_new_n361_), .B0(new_new_n363_), .Y(new_new_n365_));
  NA2        g0343(.A(i_2_), .B(i_7_), .Y(new_new_n366_));
  NO2        g0344(.A(new_new_n362_), .B(i_10_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n366_), .C(new_new_n242_), .Y(new_new_n368_));
  AOI210     g0346(.A0(new_new_n368_), .A1(new_new_n365_), .B0(new_new_n185_), .Y(new_new_n369_));
  AOI210     g0347(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n370_));
  OAI210     g0348(.A0(new_new_n370_), .A1(new_new_n188_), .B0(new_new_n367_), .Y(new_new_n371_));
  AOI220     g0349(.A0(new_new_n367_), .A1(new_new_n325_), .B0(new_new_n238_), .B1(new_new_n188_), .Y(new_new_n372_));
  AOI210     g0350(.A0(new_new_n372_), .A1(new_new_n371_), .B0(i_5_), .Y(new_new_n373_));
  NO4        g0351(.A(new_new_n373_), .B(new_new_n369_), .C(new_new_n360_), .D(new_new_n352_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n374_), .B(new_new_n347_), .Y(new_new_n375_));
  NO2        g0353(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n376_));
  AN2        g0354(.A(i_12_), .B(i_5_), .Y(new_new_n377_));
  NO2        g0355(.A(i_4_), .B(new_new_n26_), .Y(new_new_n378_));
  NA2        g0356(.A(new_new_n378_), .B(new_new_n377_), .Y(new_new_n379_));
  NO2        g0357(.A(i_11_), .B(i_6_), .Y(new_new_n380_));
  NA3        g0358(.A(new_new_n380_), .B(new_new_n312_), .C(new_new_n225_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n381_), .B(new_new_n379_), .Y(new_new_n382_));
  NO2        g0360(.A(new_new_n241_), .B(i_5_), .Y(new_new_n383_));
  NO2        g0361(.A(i_5_), .B(i_10_), .Y(new_new_n384_));
  AOI220     g0362(.A0(new_new_n384_), .A1(new_new_n268_), .B0(new_new_n383_), .B1(new_new_n198_), .Y(new_new_n385_));
  NA2        g0363(.A(new_new_n146_), .B(new_new_n46_), .Y(new_new_n386_));
  NO2        g0364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n382_), .B0(new_new_n376_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n152_), .B(new_new_n87_), .Y(new_new_n390_));
  OAI210     g0368(.A0(new_new_n390_), .A1(new_new_n382_), .B0(new_new_n389_), .Y(new_new_n391_));
  NO3        g0369(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n392_));
  NO2        g0370(.A(i_3_), .B(new_new_n103_), .Y(new_new_n393_));
  NO2        g0371(.A(i_11_), .B(i_12_), .Y(new_new_n394_));
  NA2        g0372(.A(new_new_n384_), .B(new_new_n236_), .Y(new_new_n395_));
  NA3        g0373(.A(new_new_n114_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n396_));
  OAI220     g0374(.A0(new_new_n396_), .A1(new_new_n220_), .B0(new_new_n395_), .B1(new_new_n320_), .Y(new_new_n397_));
  NAi21      g0375(.An(i_13_), .B(i_0_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n398_), .B(new_new_n239_), .Y(new_new_n399_));
  NA2        g0377(.A(new_new_n397_), .B(new_new_n399_), .Y(new_new_n400_));
  NA3        g0378(.A(new_new_n400_), .B(new_new_n391_), .C(new_new_n388_), .Y(new_new_n401_));
  NA2        g0379(.A(new_new_n45_), .B(new_new_n225_), .Y(new_new_n402_));
  NO3        g0380(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n403_));
  NO2        g0381(.A(i_0_), .B(i_11_), .Y(new_new_n404_));
  INV        g0382(.A(i_5_), .Y(new_new_n405_));
  AN2        g0383(.A(i_1_), .B(i_6_), .Y(new_new_n406_));
  NOi21      g0384(.An(i_2_), .B(i_12_), .Y(new_new_n407_));
  NA2        g0385(.A(new_new_n407_), .B(new_new_n406_), .Y(new_new_n408_));
  NO2        g0386(.A(new_new_n408_), .B(new_new_n405_), .Y(new_new_n409_));
  NA2        g0387(.A(new_new_n144_), .B(i_9_), .Y(new_new_n410_));
  NO2        g0388(.A(new_new_n410_), .B(i_4_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n409_), .B(new_new_n411_), .Y(new_new_n412_));
  NAi21      g0390(.An(i_9_), .B(i_4_), .Y(new_new_n413_));
  OR2        g0391(.A(i_13_), .B(i_10_), .Y(new_new_n414_));
  NO3        g0392(.A(new_new_n414_), .B(new_new_n119_), .C(new_new_n413_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n175_), .B(new_new_n125_), .Y(new_new_n416_));
  OR2        g0394(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n103_), .B(new_new_n25_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n274_), .B(new_new_n418_), .Y(new_new_n419_));
  NA2        g0397(.A(new_new_n272_), .B(new_new_n212_), .Y(new_new_n420_));
  OAI220     g0398(.A0(new_new_n420_), .A1(new_new_n417_), .B0(new_new_n419_), .B1(new_new_n331_), .Y(new_new_n421_));
  INV        g0399(.A(new_new_n421_), .Y(new_new_n422_));
  AOI210     g0400(.A0(new_new_n422_), .A1(new_new_n412_), .B0(new_new_n26_), .Y(new_new_n423_));
  AOI220     g0401(.A0(new_new_n284_), .A1(new_new_n276_), .B0(new_new_n278_), .B1(new_new_n302_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(new_new_n172_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n184_), .B(new_new_n87_), .Y(new_new_n426_));
  INV        g0404(.A(new_new_n425_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n196_), .B(new_new_n98_), .Y(new_new_n428_));
  NA3        g0406(.A(new_new_n312_), .B(new_new_n165_), .C(new_new_n87_), .Y(new_new_n429_));
  AOI210     g0407(.A0(new_new_n429_), .A1(new_new_n428_), .B0(new_new_n310_), .Y(new_new_n430_));
  NA2        g0408(.A(new_new_n193_), .B(i_10_), .Y(new_new_n431_));
  NA3        g0409(.A(new_new_n255_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n433_));
  NO2        g0411(.A(i_3_), .B(new_new_n49_), .Y(new_new_n434_));
  NA3        g0412(.A(new_new_n325_), .B(new_new_n324_), .C(new_new_n434_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n304_), .B(new_new_n309_), .Y(new_new_n436_));
  OAI210     g0414(.A0(new_new_n436_), .A1(new_new_n189_), .B0(new_new_n435_), .Y(new_new_n437_));
  NO3        g0415(.A(new_new_n437_), .B(new_new_n433_), .C(new_new_n430_), .Y(new_new_n438_));
  AOI210     g0416(.A0(new_new_n438_), .A1(new_new_n427_), .B0(new_new_n269_), .Y(new_new_n439_));
  NO4        g0417(.A(new_new_n439_), .B(new_new_n423_), .C(new_new_n401_), .D(new_new_n375_), .Y(new_new_n440_));
  NO2        g0418(.A(new_new_n64_), .B(i_4_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n74_), .B(i_13_), .Y(new_new_n442_));
  NO2        g0420(.A(i_10_), .B(i_9_), .Y(new_new_n443_));
  NAi21      g0421(.An(i_12_), .B(i_8_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n444_), .B(i_3_), .Y(new_new_n445_));
  NO2        g0423(.A(new_new_n47_), .B(i_4_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n446_), .B(new_new_n106_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n447_), .B(new_new_n205_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n297_), .B(i_0_), .Y(new_new_n449_));
  NO3        g0427(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n450_));
  NA2        g0428(.A(new_new_n266_), .B(new_new_n99_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n451_), .B(new_new_n450_), .Y(new_new_n452_));
  NA2        g0430(.A(i_8_), .B(i_9_), .Y(new_new_n453_));
  AOI210     g0431(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n454_));
  OR2        g0432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n274_), .B(new_new_n206_), .Y(new_new_n456_));
  OAI220     g0434(.A0(new_new_n456_), .A1(new_new_n455_), .B0(new_new_n452_), .B1(new_new_n449_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n249_), .B(new_new_n296_), .Y(new_new_n458_));
  NO3        g0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n459_));
  INV        g0437(.A(new_new_n459_), .Y(new_new_n460_));
  NA3        g0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n461_));
  NA4        g0439(.A(new_new_n147_), .B(new_new_n117_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n461_), .B0(new_new_n460_), .B1(new_new_n458_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n463_), .B(new_new_n457_), .C(new_new_n448_), .Y(new_new_n464_));
  NA2        g0442(.A(new_new_n283_), .B(new_new_n110_), .Y(new_new_n465_));
  OR2        g0443(.A(new_new_n465_), .B(new_new_n209_), .Y(new_new_n466_));
  OA210      g0444(.A0(new_new_n341_), .A1(new_new_n103_), .B0(new_new_n285_), .Y(new_new_n467_));
  OA220      g0445(.A0(new_new_n467_), .A1(new_new_n164_), .B0(new_new_n466_), .B1(new_new_n232_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n98_), .B(i_13_), .Y(new_new_n469_));
  NA2        g0447(.A(new_new_n426_), .B(new_new_n376_), .Y(new_new_n470_));
  NO2        g0448(.A(i_2_), .B(i_13_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n470_), .B(new_new_n469_), .Y(new_new_n472_));
  NO3        g0450(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n473_));
  NO2        g0451(.A(i_6_), .B(i_7_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NO2        g0453(.A(i_11_), .B(i_1_), .Y(new_new_n476_));
  NO2        g0454(.A(new_new_n74_), .B(i_3_), .Y(new_new_n477_));
  OR2        g0455(.A(i_11_), .B(i_8_), .Y(new_new_n478_));
  NOi21      g0456(.An(i_2_), .B(i_7_), .Y(new_new_n479_));
  NAi31      g0457(.An(new_new_n478_), .B(new_new_n479_), .C(new_new_n477_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n414_), .B(i_6_), .Y(new_new_n481_));
  NA3        g0459(.A(new_new_n481_), .B(new_new_n441_), .C(new_new_n76_), .Y(new_new_n482_));
  NO2        g0460(.A(new_new_n482_), .B(new_new_n480_), .Y(new_new_n483_));
  NO2        g0461(.A(i_3_), .B(new_new_n193_), .Y(new_new_n484_));
  NO2        g0462(.A(i_6_), .B(i_10_), .Y(new_new_n485_));
  NA4        g0463(.A(new_new_n485_), .B(new_new_n301_), .C(new_new_n484_), .D(new_new_n236_), .Y(new_new_n486_));
  NO2        g0464(.A(new_new_n486_), .B(new_new_n157_), .Y(new_new_n487_));
  NA3        g0465(.A(new_new_n243_), .B(new_new_n174_), .C(new_new_n134_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n489_));
  NO2        g0467(.A(new_new_n159_), .B(i_3_), .Y(new_new_n490_));
  NAi31      g0468(.An(new_new_n489_), .B(new_new_n490_), .C(new_new_n226_), .Y(new_new_n491_));
  NA3        g0469(.A(new_new_n389_), .B(new_new_n182_), .C(new_new_n151_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n492_), .B(new_new_n491_), .C(new_new_n488_), .Y(new_new_n493_));
  NO4        g0471(.A(new_new_n493_), .B(new_new_n487_), .C(new_new_n483_), .D(new_new_n472_), .Y(new_new_n494_));
  NA2        g0472(.A(new_new_n450_), .B(new_new_n377_), .Y(new_new_n495_));
  NA2        g0473(.A(new_new_n459_), .B(new_new_n384_), .Y(new_new_n496_));
  NO2        g0474(.A(new_new_n496_), .B(new_new_n224_), .Y(new_new_n497_));
  NAi21      g0475(.An(new_new_n218_), .B(new_new_n394_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n325_), .B(new_new_n219_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n26_), .B(i_5_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n499_), .B(new_new_n498_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n27_), .B(i_10_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n301_), .B(new_new_n238_), .Y(new_new_n503_));
  OAI220     g0481(.A0(new_new_n503_), .A1(new_new_n432_), .B0(new_new_n502_), .B1(new_new_n469_), .Y(new_new_n504_));
  NA4        g0482(.A(new_new_n294_), .B(new_new_n223_), .C(new_new_n74_), .D(new_new_n236_), .Y(new_new_n505_));
  NO2        g0483(.A(new_new_n505_), .B(new_new_n475_), .Y(new_new_n506_));
  NO4        g0484(.A(new_new_n506_), .B(new_new_n504_), .C(new_new_n501_), .D(new_new_n497_), .Y(new_new_n507_));
  NA4        g0485(.A(new_new_n507_), .B(new_new_n494_), .C(new_new_n468_), .D(new_new_n464_), .Y(new_new_n508_));
  NA3        g0486(.A(new_new_n294_), .B(new_new_n179_), .C(new_new_n177_), .Y(new_new_n509_));
  OAI210     g0487(.A0(new_new_n289_), .A1(new_new_n183_), .B0(new_new_n509_), .Y(new_new_n510_));
  AN2        g0488(.A(new_new_n276_), .B(new_new_n234_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n511_), .B(new_new_n510_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n124_), .B(new_new_n113_), .Y(new_new_n513_));
  AN2        g0491(.A(new_new_n513_), .B(new_new_n450_), .Y(new_new_n514_));
  NA2        g0492(.A(new_new_n301_), .B(new_new_n166_), .Y(new_new_n515_));
  OAI210     g0493(.A0(new_new_n515_), .A1(new_new_n232_), .B0(new_new_n295_), .Y(new_new_n516_));
  AOI220     g0494(.A0(new_new_n516_), .A1(new_new_n311_), .B0(new_new_n514_), .B1(new_new_n297_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n377_), .B(new_new_n225_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n346_), .B(new_new_n74_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n364_), .B(new_new_n356_), .Y(new_new_n520_));
  OR2        g0498(.A(new_new_n518_), .B(new_new_n520_), .Y(new_new_n521_));
  NO2        g0499(.A(new_new_n36_), .B(i_8_), .Y(new_new_n522_));
  NAi41      g0500(.An(new_new_n519_), .B(new_new_n485_), .C(new_new_n522_), .D(new_new_n47_), .Y(new_new_n523_));
  AOI210     g0501(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n415_), .Y(new_new_n524_));
  NA3        g0502(.A(new_new_n524_), .B(new_new_n523_), .C(new_new_n521_), .Y(new_new_n525_));
  INV        g0503(.A(new_new_n525_), .Y(new_new_n526_));
  NA2        g0504(.A(new_new_n255_), .B(new_new_n65_), .Y(new_new_n527_));
  OAI210     g0505(.A0(i_8_), .A1(new_new_n527_), .B0(new_new_n136_), .Y(new_new_n528_));
  NO2        g0506(.A(i_7_), .B(new_new_n199_), .Y(new_new_n529_));
  OR2        g0507(.A(new_new_n184_), .B(i_4_), .Y(new_new_n530_));
  NO2        g0508(.A(new_new_n530_), .B(new_new_n87_), .Y(new_new_n531_));
  AOI220     g0509(.A0(new_new_n531_), .A1(new_new_n529_), .B0(new_new_n528_), .B1(new_new_n416_), .Y(new_new_n532_));
  NA4        g0510(.A(new_new_n532_), .B(new_new_n526_), .C(new_new_n517_), .D(new_new_n512_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n383_), .B(new_new_n283_), .Y(new_new_n534_));
  OAI210     g0512(.A0(new_new_n379_), .A1(new_new_n171_), .B0(new_new_n534_), .Y(new_new_n535_));
  NO2        g0513(.A(i_12_), .B(new_new_n193_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n536_), .B(new_new_n225_), .Y(new_new_n537_));
  NO3        g0515(.A(new_new_n1058_), .B(new_new_n537_), .C(new_new_n465_), .Y(new_new_n538_));
  NOi31      g0516(.An(new_new_n304_), .B(new_new_n414_), .C(new_new_n38_), .Y(new_new_n539_));
  OAI210     g0517(.A0(new_new_n539_), .A1(new_new_n538_), .B0(new_new_n535_), .Y(new_new_n540_));
  NO2        g0518(.A(i_8_), .B(i_7_), .Y(new_new_n541_));
  AOI220     g0519(.A0(new_new_n312_), .A1(new_new_n40_), .B0(new_new_n235_), .B1(new_new_n208_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n542_), .B(new_new_n530_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n45_), .B(i_10_), .Y(new_new_n544_));
  NO2        g0522(.A(new_new_n544_), .B(i_6_), .Y(new_new_n545_));
  NA3        g0523(.A(new_new_n545_), .B(new_new_n543_), .C(new_new_n541_), .Y(new_new_n546_));
  NOi31      g0524(.An(new_new_n278_), .B(new_new_n289_), .C(new_new_n183_), .Y(new_new_n547_));
  NA3        g0525(.A(new_new_n294_), .B(new_new_n177_), .C(new_new_n98_), .Y(new_new_n548_));
  NO2        g0526(.A(new_new_n221_), .B(new_new_n45_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n159_), .B(i_5_), .Y(new_new_n550_));
  NA3        g0528(.A(new_new_n550_), .B(new_new_n402_), .C(new_new_n307_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n551_), .A1(new_new_n549_), .B0(new_new_n548_), .Y(new_new_n552_));
  OAI210     g0530(.A0(new_new_n552_), .A1(new_new_n547_), .B0(new_new_n459_), .Y(new_new_n553_));
  NA3        g0531(.A(new_new_n553_), .B(new_new_n546_), .C(new_new_n540_), .Y(new_new_n554_));
  NA3        g0532(.A(new_new_n219_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n274_), .B(new_new_n85_), .Y(new_new_n556_));
  AOI210     g0534(.A0(new_new_n555_), .A1(new_new_n336_), .B0(new_new_n556_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n284_), .B(new_new_n276_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n558_), .B(new_new_n176_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n560_));
  NA2        g0538(.A(new_new_n443_), .B(new_new_n221_), .Y(new_new_n561_));
  NO2        g0539(.A(new_new_n560_), .B(new_new_n561_), .Y(new_new_n562_));
  AOI210     g0540(.A0(new_new_n357_), .A1(new_new_n47_), .B0(new_new_n361_), .Y(new_new_n563_));
  NA2        g0541(.A(i_0_), .B(new_new_n49_), .Y(new_new_n564_));
  NA3        g0542(.A(new_new_n536_), .B(new_new_n270_), .C(new_new_n564_), .Y(new_new_n565_));
  NO2        g0543(.A(new_new_n563_), .B(new_new_n565_), .Y(new_new_n566_));
  NO4        g0544(.A(new_new_n566_), .B(new_new_n562_), .C(new_new_n559_), .D(new_new_n557_), .Y(new_new_n567_));
  NO4        g0545(.A(new_new_n250_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n568_));
  NO3        g0546(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n569_));
  NO2        g0547(.A(new_new_n233_), .B(new_new_n36_), .Y(new_new_n570_));
  AN2        g0548(.A(new_new_n570_), .B(new_new_n569_), .Y(new_new_n571_));
  OA210      g0549(.A0(new_new_n571_), .A1(new_new_n568_), .B0(new_new_n346_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n414_), .B(i_1_), .Y(new_new_n573_));
  NOi31      g0551(.An(new_new_n573_), .B(new_new_n451_), .C(new_new_n74_), .Y(new_new_n574_));
  AN4        g0552(.A(new_new_n574_), .B(new_new_n411_), .C(new_new_n500_), .D(i_2_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n424_), .B(new_new_n180_), .Y(new_new_n576_));
  NO3        g0554(.A(new_new_n576_), .B(new_new_n575_), .C(new_new_n572_), .Y(new_new_n577_));
  NOi21      g0555(.An(i_10_), .B(i_6_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n579_));
  AOI220     g0557(.A0(new_new_n274_), .A1(new_new_n579_), .B0(new_new_n270_), .B1(new_new_n578_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n580_), .B(new_new_n449_), .Y(new_new_n581_));
  NO2        g0559(.A(new_new_n116_), .B(new_new_n23_), .Y(new_new_n582_));
  NOi31      g0560(.An(new_new_n148_), .B(i_10_), .C(new_new_n320_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n583_), .B(new_new_n581_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n519_), .B(new_new_n372_), .Y(new_new_n585_));
  INV        g0563(.A(new_new_n307_), .Y(new_new_n586_));
  NO2        g0564(.A(i_12_), .B(new_new_n87_), .Y(new_new_n587_));
  NA3        g0565(.A(new_new_n587_), .B(new_new_n270_), .C(new_new_n564_), .Y(new_new_n588_));
  NA3        g0566(.A(new_new_n380_), .B(new_new_n274_), .C(new_new_n219_), .Y(new_new_n589_));
  AOI210     g0567(.A0(new_new_n589_), .A1(new_new_n588_), .B0(new_new_n586_), .Y(new_new_n590_));
  OR2        g0568(.A(i_2_), .B(i_5_), .Y(new_new_n591_));
  OR2        g0569(.A(new_new_n591_), .B(new_new_n406_), .Y(new_new_n592_));
  AOI210     g0570(.A0(new_new_n366_), .A1(new_new_n242_), .B0(new_new_n198_), .Y(new_new_n593_));
  AOI210     g0571(.A0(new_new_n593_), .A1(new_new_n592_), .B0(new_new_n498_), .Y(new_new_n594_));
  NO3        g0572(.A(new_new_n594_), .B(new_new_n590_), .C(new_new_n585_), .Y(new_new_n595_));
  NA4        g0573(.A(new_new_n595_), .B(new_new_n584_), .C(new_new_n577_), .D(new_new_n567_), .Y(new_new_n596_));
  NO4        g0574(.A(new_new_n596_), .B(new_new_n554_), .C(new_new_n533_), .D(new_new_n508_), .Y(new_new_n597_));
  NA4        g0575(.A(new_new_n597_), .B(new_new_n440_), .C(new_new_n345_), .D(new_new_n300_), .Y(men7));
  NO2        g0576(.A(new_new_n94_), .B(new_new_n55_), .Y(new_new_n599_));
  NA2        g0577(.A(new_new_n485_), .B(new_new_n85_), .Y(new_new_n600_));
  NA2        g0578(.A(i_11_), .B(new_new_n193_), .Y(new_new_n601_));
  NA3        g0579(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n236_), .B(i_4_), .Y(new_new_n603_));
  NA2        g0581(.A(new_new_n603_), .B(i_8_), .Y(new_new_n604_));
  NO2        g0582(.A(new_new_n107_), .B(new_new_n602_), .Y(new_new_n605_));
  NA2        g0583(.A(i_2_), .B(new_new_n87_), .Y(new_new_n606_));
  OAI210     g0584(.A0(new_new_n88_), .A1(new_new_n203_), .B0(new_new_n204_), .Y(new_new_n607_));
  NO2        g0585(.A(i_7_), .B(new_new_n37_), .Y(new_new_n608_));
  NA2        g0586(.A(i_4_), .B(i_8_), .Y(new_new_n609_));
  AOI210     g0587(.A0(new_new_n609_), .A1(new_new_n294_), .B0(new_new_n608_), .Y(new_new_n610_));
  OAI220     g0588(.A0(new_new_n610_), .A1(new_new_n606_), .B0(new_new_n607_), .B1(i_13_), .Y(new_new_n611_));
  NO3        g0589(.A(new_new_n611_), .B(new_new_n605_), .C(new_new_n599_), .Y(new_new_n612_));
  AOI210     g0590(.A0(new_new_n130_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n613_));
  AOI210     g0591(.A0(new_new_n613_), .A1(new_new_n236_), .B0(new_new_n163_), .Y(new_new_n614_));
  OR2        g0592(.A(i_6_), .B(i_10_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n615_), .B(new_new_n23_), .Y(new_new_n616_));
  OR3        g0594(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n617_));
  NO3        g0595(.A(new_new_n617_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n618_));
  INV        g0596(.A(new_new_n200_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n618_), .B(new_new_n616_), .Y(new_new_n620_));
  OA220      g0598(.A0(new_new_n620_), .A1(new_new_n586_), .B0(new_new_n614_), .B1(new_new_n267_), .Y(new_new_n621_));
  AOI210     g0599(.A0(new_new_n621_), .A1(new_new_n612_), .B0(new_new_n64_), .Y(new_new_n622_));
  NOi21      g0600(.An(i_11_), .B(i_7_), .Y(new_new_n623_));
  AO210      g0601(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n624_), .B(new_new_n623_), .Y(new_new_n625_));
  NA2        g0603(.A(new_new_n625_), .B(new_new_n208_), .Y(new_new_n626_));
  NA3        g0604(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n627_));
  NAi31      g0605(.An(new_new_n627_), .B(new_new_n217_), .C(i_11_), .Y(new_new_n628_));
  AOI210     g0606(.A0(new_new_n628_), .A1(new_new_n626_), .B0(new_new_n64_), .Y(new_new_n629_));
  OR2        g0607(.A(new_new_n372_), .B(new_new_n41_), .Y(new_new_n630_));
  NO3        g0608(.A(new_new_n257_), .B(new_new_n210_), .C(new_new_n601_), .Y(new_new_n631_));
  OAI210     g0609(.A0(new_new_n631_), .A1(new_new_n226_), .B0(new_new_n64_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n407_), .B(new_new_n31_), .Y(new_new_n633_));
  OR2        g0611(.A(new_new_n210_), .B(new_new_n110_), .Y(new_new_n634_));
  NA2        g0612(.A(new_new_n634_), .B(new_new_n633_), .Y(new_new_n635_));
  NO2        g0613(.A(new_new_n64_), .B(i_9_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n636_), .B(i_4_), .Y(new_new_n637_));
  NA2        g0615(.A(new_new_n637_), .B(new_new_n635_), .Y(new_new_n638_));
  NO2        g0616(.A(i_1_), .B(i_12_), .Y(new_new_n639_));
  NA3        g0617(.A(new_new_n639_), .B(new_new_n111_), .C(new_new_n24_), .Y(new_new_n640_));
  BUFFER     g0618(.A(new_new_n640_), .Y(new_new_n641_));
  NA4        g0619(.A(new_new_n641_), .B(new_new_n638_), .C(new_new_n632_), .D(new_new_n630_), .Y(new_new_n642_));
  OAI210     g0620(.A0(new_new_n642_), .A1(new_new_n629_), .B0(i_6_), .Y(new_new_n643_));
  NO2        g0621(.A(new_new_n627_), .B(new_new_n110_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n644_), .B(new_new_n587_), .Y(new_new_n645_));
  NO2        g0623(.A(new_new_n236_), .B(new_new_n87_), .Y(new_new_n646_));
  NO2        g0624(.A(new_new_n646_), .B(i_11_), .Y(new_new_n647_));
  NA2        g0625(.A(new_new_n645_), .B(new_new_n452_), .Y(new_new_n648_));
  NO4        g0626(.A(new_new_n217_), .B(new_new_n130_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n649_), .B(new_new_n636_), .Y(new_new_n650_));
  NA2        g0628(.A(new_new_n236_), .B(i_6_), .Y(new_new_n651_));
  NO3        g0629(.A(new_new_n615_), .B(new_new_n233_), .C(new_new_n23_), .Y(new_new_n652_));
  AOI210     g0630(.A0(i_1_), .A1(new_new_n258_), .B0(new_new_n652_), .Y(new_new_n653_));
  OAI210     g0631(.A0(new_new_n653_), .A1(new_new_n45_), .B0(new_new_n650_), .Y(new_new_n654_));
  NA3        g0632(.A(new_new_n541_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n655_));
  INV        g0633(.A(i_2_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n140_), .B(i_9_), .Y(new_new_n657_));
  NA3        g0635(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n47_), .B(i_1_), .Y(new_new_n659_));
  NA3        g0637(.A(new_new_n659_), .B(new_new_n266_), .C(new_new_n45_), .Y(new_new_n660_));
  OAI220     g0638(.A0(new_new_n660_), .A1(new_new_n658_), .B0(new_new_n657_), .B1(new_new_n656_), .Y(new_new_n661_));
  AOI210     g0639(.A0(new_new_n476_), .A1(new_new_n418_), .B0(new_new_n240_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n662_), .B(new_new_n606_), .Y(new_new_n663_));
  NAi21      g0641(.An(new_new_n655_), .B(new_new_n93_), .Y(new_new_n664_));
  NO2        g0642(.A(i_11_), .B(new_new_n37_), .Y(new_new_n665_));
  INV        g0643(.A(new_new_n664_), .Y(new_new_n666_));
  OR3        g0644(.A(new_new_n666_), .B(new_new_n663_), .C(new_new_n661_), .Y(new_new_n667_));
  NO3        g0645(.A(new_new_n667_), .B(new_new_n654_), .C(new_new_n648_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n236_), .B(new_new_n103_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n669_), .B(new_new_n623_), .Y(new_new_n670_));
  NA2        g0648(.A(new_new_n670_), .B(i_1_), .Y(new_new_n671_));
  NO2        g0649(.A(new_new_n671_), .B(new_new_n617_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n413_), .B(new_new_n87_), .Y(new_new_n673_));
  NA2        g0651(.A(new_new_n672_), .B(new_new_n47_), .Y(new_new_n674_));
  NA2        g0652(.A(i_3_), .B(new_new_n193_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n675_), .B(new_new_n116_), .Y(new_new_n676_));
  AN2        g0654(.A(new_new_n676_), .B(new_new_n545_), .Y(new_new_n677_));
  NO2        g0655(.A(new_new_n233_), .B(new_new_n45_), .Y(new_new_n678_));
  NO3        g0656(.A(new_new_n678_), .B(new_new_n297_), .C(new_new_n237_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n119_), .B(new_new_n37_), .Y(new_new_n680_));
  NO2        g0658(.A(new_new_n680_), .B(i_6_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n87_), .B(i_9_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n682_), .B(new_new_n64_), .Y(new_new_n683_));
  NO2        g0661(.A(new_new_n683_), .B(new_new_n639_), .Y(new_new_n684_));
  NO4        g0662(.A(new_new_n684_), .B(new_new_n681_), .C(new_new_n679_), .D(i_4_), .Y(new_new_n685_));
  NA2        g0663(.A(i_1_), .B(i_3_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n453_), .B(new_new_n94_), .Y(new_new_n687_));
  AOI210     g0665(.A0(new_new_n678_), .A1(new_new_n578_), .B0(new_new_n687_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(new_new_n686_), .Y(new_new_n689_));
  NO3        g0667(.A(new_new_n689_), .B(new_new_n685_), .C(new_new_n677_), .Y(new_new_n690_));
  NA4        g0668(.A(new_new_n690_), .B(new_new_n674_), .C(new_new_n668_), .D(new_new_n643_), .Y(new_new_n691_));
  NO3        g0669(.A(new_new_n478_), .B(i_3_), .C(i_7_), .Y(new_new_n692_));
  NOi21      g0670(.An(new_new_n692_), .B(i_10_), .Y(new_new_n693_));
  OA210      g0671(.A0(new_new_n693_), .A1(new_new_n243_), .B0(new_new_n87_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n364_), .B(new_new_n363_), .Y(new_new_n695_));
  NA3        g0673(.A(new_new_n485_), .B(new_new_n522_), .C(new_new_n47_), .Y(new_new_n696_));
  NO3        g0674(.A(new_new_n479_), .B(new_new_n609_), .C(new_new_n87_), .Y(new_new_n697_));
  NA2        g0675(.A(new_new_n697_), .B(new_new_n25_), .Y(new_new_n698_));
  NA3        g0676(.A(new_new_n163_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n699_));
  NA4        g0677(.A(new_new_n699_), .B(new_new_n698_), .C(new_new_n696_), .D(new_new_n695_), .Y(new_new_n700_));
  OAI210     g0678(.A0(new_new_n700_), .A1(new_new_n694_), .B0(i_1_), .Y(new_new_n701_));
  AOI210     g0679(.A0(new_new_n266_), .A1(new_new_n99_), .B0(i_1_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n362_), .B(i_2_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n703_), .B(new_new_n702_), .Y(new_new_n704_));
  AOI210     g0682(.A0(new_new_n704_), .A1(new_new_n701_), .B0(i_13_), .Y(new_new_n705_));
  OR2        g0683(.A(i_11_), .B(i_7_), .Y(new_new_n706_));
  NA3        g0684(.A(new_new_n706_), .B(new_new_n108_), .C(new_new_n140_), .Y(new_new_n707_));
  AOI220     g0685(.A0(new_new_n471_), .A1(new_new_n163_), .B0(new_new_n446_), .B1(new_new_n140_), .Y(new_new_n708_));
  OAI210     g0686(.A0(new_new_n708_), .A1(new_new_n45_), .B0(new_new_n707_), .Y(new_new_n709_));
  AOI210     g0687(.A0(new_new_n658_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n710_));
  NO2        g0688(.A(new_new_n479_), .B(new_new_n24_), .Y(new_new_n711_));
  AOI220     g0689(.A0(new_new_n711_), .A1(new_new_n673_), .B0(new_new_n243_), .B1(new_new_n133_), .Y(new_new_n712_));
  OAI220     g0690(.A0(new_new_n712_), .A1(new_new_n41_), .B0(new_new_n1057_), .B1(new_new_n94_), .Y(new_new_n713_));
  AOI210     g0691(.A0(new_new_n709_), .A1(new_new_n322_), .B0(new_new_n713_), .Y(new_new_n714_));
  NA2        g0692(.A(new_new_n380_), .B(new_new_n659_), .Y(new_new_n715_));
  NO2        g0693(.A(new_new_n715_), .B(new_new_n241_), .Y(new_new_n716_));
  AOI210     g0694(.A0(new_new_n444_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n717_));
  NOi31      g0695(.An(new_new_n717_), .B(new_new_n600_), .C(new_new_n45_), .Y(new_new_n718_));
  NA2        g0696(.A(new_new_n129_), .B(i_13_), .Y(new_new_n719_));
  NO2        g0697(.A(new_new_n658_), .B(new_new_n116_), .Y(new_new_n720_));
  INV        g0698(.A(new_new_n720_), .Y(new_new_n721_));
  OAI220     g0699(.A0(new_new_n721_), .A1(new_new_n72_), .B0(new_new_n719_), .B1(new_new_n702_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n26_), .B(new_new_n193_), .Y(new_new_n723_));
  NA2        g0701(.A(new_new_n723_), .B(i_7_), .Y(new_new_n724_));
  NO3        g0702(.A(new_new_n479_), .B(new_new_n236_), .C(new_new_n87_), .Y(new_new_n725_));
  NA2        g0703(.A(new_new_n725_), .B(new_new_n724_), .Y(new_new_n726_));
  AOI220     g0704(.A0(new_new_n380_), .A1(new_new_n659_), .B0(new_new_n93_), .B1(new_new_n104_), .Y(new_new_n727_));
  OAI220     g0705(.A0(new_new_n727_), .A1(new_new_n604_), .B0(new_new_n726_), .B1(new_new_n619_), .Y(new_new_n728_));
  NO4        g0706(.A(new_new_n728_), .B(new_new_n722_), .C(new_new_n718_), .D(new_new_n716_), .Y(new_new_n729_));
  OR2        g0707(.A(i_11_), .B(i_6_), .Y(new_new_n730_));
  NA3        g0708(.A(new_new_n603_), .B(new_new_n723_), .C(i_7_), .Y(new_new_n731_));
  AOI210     g0709(.A0(new_new_n731_), .A1(new_new_n721_), .B0(new_new_n730_), .Y(new_new_n732_));
  NA3        g0710(.A(new_new_n407_), .B(new_new_n608_), .C(new_new_n99_), .Y(new_new_n733_));
  NA2        g0711(.A(new_new_n647_), .B(i_13_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n104_), .B(new_new_n723_), .Y(new_new_n735_));
  NAi21      g0713(.An(i_11_), .B(i_12_), .Y(new_new_n736_));
  NOi41      g0714(.An(new_new_n112_), .B(new_new_n736_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n737_));
  NO3        g0715(.A(new_new_n479_), .B(new_new_n587_), .C(new_new_n609_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n738_), .A1(new_new_n301_), .B0(new_new_n737_), .B1(new_new_n735_), .Y(new_new_n739_));
  NA3        g0717(.A(new_new_n739_), .B(new_new_n734_), .C(new_new_n733_), .Y(new_new_n740_));
  OAI210     g0718(.A0(new_new_n740_), .A1(new_new_n732_), .B0(new_new_n64_), .Y(new_new_n741_));
  NO2        g0719(.A(i_2_), .B(i_12_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n361_), .B(new_new_n742_), .Y(new_new_n743_));
  NA2        g0721(.A(i_8_), .B(new_new_n25_), .Y(new_new_n744_));
  NO3        g0722(.A(new_new_n744_), .B(new_new_n378_), .C(new_new_n603_), .Y(new_new_n745_));
  OAI210     g0723(.A0(new_new_n745_), .A1(new_new_n363_), .B0(new_new_n361_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n130_), .B(i_2_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n746_), .B(new_new_n743_), .Y(new_new_n748_));
  NA3        g0726(.A(new_new_n748_), .B(new_new_n46_), .C(new_new_n225_), .Y(new_new_n749_));
  NA4        g0727(.A(new_new_n749_), .B(new_new_n741_), .C(new_new_n729_), .D(new_new_n714_), .Y(new_new_n750_));
  OR4        g0728(.A(new_new_n750_), .B(new_new_n705_), .C(new_new_n691_), .D(new_new_n622_), .Y(men5));
  NA2        g0729(.A(new_new_n670_), .B(new_new_n268_), .Y(new_new_n752_));
  AN2        g0730(.A(new_new_n24_), .B(i_10_), .Y(new_new_n753_));
  NA3        g0731(.A(new_new_n753_), .B(new_new_n742_), .C(new_new_n110_), .Y(new_new_n754_));
  NO2        g0732(.A(new_new_n604_), .B(i_11_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n88_), .B(new_new_n755_), .Y(new_new_n756_));
  NA3        g0734(.A(new_new_n756_), .B(new_new_n754_), .C(new_new_n752_), .Y(new_new_n757_));
  NO3        g0735(.A(i_11_), .B(new_new_n236_), .C(i_13_), .Y(new_new_n758_));
  NO2        g0736(.A(new_new_n126_), .B(new_new_n23_), .Y(new_new_n759_));
  NA2        g0737(.A(i_12_), .B(i_8_), .Y(new_new_n760_));
  OAI210     g0738(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n760_), .Y(new_new_n761_));
  INV        g0739(.A(new_new_n443_), .Y(new_new_n762_));
  AOI220     g0740(.A0(new_new_n307_), .A1(new_new_n582_), .B0(new_new_n761_), .B1(new_new_n759_), .Y(new_new_n763_));
  INV        g0741(.A(new_new_n763_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n764_), .B(new_new_n757_), .Y(new_new_n765_));
  INV        g0743(.A(new_new_n174_), .Y(new_new_n766_));
  INV        g0744(.A(new_new_n243_), .Y(new_new_n767_));
  OAI210     g0745(.A0(new_new_n703_), .A1(new_new_n445_), .B0(new_new_n112_), .Y(new_new_n768_));
  AOI210     g0746(.A0(new_new_n768_), .A1(new_new_n767_), .B0(new_new_n766_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n453_), .B(new_new_n26_), .Y(new_new_n770_));
  NO2        g0748(.A(new_new_n770_), .B(new_new_n418_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(i_2_), .Y(new_new_n772_));
  INV        g0750(.A(new_new_n772_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n414_), .Y(new_new_n774_));
  AOI210     g0752(.A0(new_new_n774_), .A1(new_new_n773_), .B0(new_new_n769_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n190_), .B(new_new_n127_), .Y(new_new_n776_));
  OAI210     g0754(.A0(new_new_n776_), .A1(new_new_n759_), .B0(i_2_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n175_), .Y(new_new_n778_));
  NO3        g0756(.A(new_new_n624_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n779_));
  AOI210     g0757(.A0(new_new_n778_), .A1(new_new_n88_), .B0(new_new_n779_), .Y(new_new_n780_));
  AOI210     g0758(.A0(new_new_n780_), .A1(new_new_n777_), .B0(new_new_n193_), .Y(new_new_n781_));
  OA210      g0759(.A0(new_new_n625_), .A1(new_new_n128_), .B0(i_13_), .Y(new_new_n782_));
  NA2        g0760(.A(new_new_n200_), .B(new_new_n203_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n153_), .B(new_new_n601_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n784_), .A1(new_new_n783_), .B0(new_new_n366_), .Y(new_new_n785_));
  AOI210     g0763(.A0(new_new_n210_), .A1(new_new_n150_), .B0(new_new_n522_), .Y(new_new_n786_));
  NA2        g0764(.A(new_new_n786_), .B(new_new_n418_), .Y(new_new_n787_));
  NO2        g0765(.A(new_new_n104_), .B(new_new_n45_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n290_), .Y(new_new_n789_));
  NA4        g0767(.A(new_new_n789_), .B(new_new_n294_), .C(new_new_n126_), .D(new_new_n43_), .Y(new_new_n790_));
  OAI210     g0768(.A0(new_new_n790_), .A1(new_new_n788_), .B0(new_new_n787_), .Y(new_new_n791_));
  NO4        g0769(.A(new_new_n791_), .B(new_new_n785_), .C(new_new_n782_), .D(new_new_n781_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n582_), .B(new_new_n28_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n758_), .B(new_new_n271_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n794_), .B(new_new_n793_), .Y(new_new_n795_));
  NO2        g0773(.A(new_new_n63_), .B(i_12_), .Y(new_new_n796_));
  NO2        g0774(.A(new_new_n796_), .B(new_new_n128_), .Y(new_new_n797_));
  NO2        g0775(.A(new_new_n797_), .B(new_new_n601_), .Y(new_new_n798_));
  AOI220     g0776(.A0(new_new_n798_), .A1(new_new_n36_), .B0(new_new_n795_), .B1(new_new_n47_), .Y(new_new_n799_));
  NA4        g0777(.A(new_new_n799_), .B(new_new_n792_), .C(new_new_n775_), .D(new_new_n765_), .Y(men6));
  NA4        g0778(.A(new_new_n384_), .B(new_new_n484_), .C(new_new_n72_), .D(new_new_n103_), .Y(new_new_n801_));
  INV        g0779(.A(new_new_n801_), .Y(new_new_n802_));
  NO2        g0780(.A(new_new_n220_), .B(new_new_n489_), .Y(new_new_n803_));
  NO2        g0781(.A(i_11_), .B(i_9_), .Y(new_new_n804_));
  NO2        g0782(.A(new_new_n802_), .B(new_new_n317_), .Y(new_new_n805_));
  OR2        g0783(.A(new_new_n805_), .B(i_12_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n367_), .B(new_new_n325_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n587_), .B(new_new_n64_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n693_), .B(new_new_n72_), .Y(new_new_n809_));
  NA3        g0787(.A(new_new_n809_), .B(new_new_n808_), .C(new_new_n807_), .Y(new_new_n810_));
  INV        g0788(.A(new_new_n197_), .Y(new_new_n811_));
  AOI220     g0789(.A0(new_new_n811_), .A1(new_new_n804_), .B0(new_new_n810_), .B1(new_new_n74_), .Y(new_new_n812_));
  INV        g0790(.A(new_new_n316_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n76_), .B(new_new_n133_), .Y(new_new_n814_));
  INV        g0792(.A(new_new_n126_), .Y(new_new_n815_));
  NA2        g0793(.A(new_new_n815_), .B(new_new_n47_), .Y(new_new_n816_));
  AOI210     g0794(.A0(new_new_n816_), .A1(new_new_n814_), .B0(new_new_n813_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n250_), .B(i_9_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n818_), .B(new_new_n796_), .Y(new_new_n819_));
  AOI210     g0797(.A0(new_new_n819_), .A1(new_new_n520_), .B0(new_new_n185_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n32_), .B(i_11_), .Y(new_new_n821_));
  NA3        g0799(.A(new_new_n821_), .B(new_new_n474_), .C(new_new_n384_), .Y(new_new_n822_));
  NAi32      g0800(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n823_));
  NO2        g0801(.A(new_new_n730_), .B(new_new_n823_), .Y(new_new_n824_));
  NAi21      g0802(.An(new_new_n824_), .B(new_new_n822_), .Y(new_new_n825_));
  OR3        g0803(.A(new_new_n825_), .B(new_new_n820_), .C(new_new_n817_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n706_), .B(i_2_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n828_));
  NO2        g0806(.A(new_new_n828_), .B(new_new_n406_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n829_), .B(new_new_n827_), .Y(new_new_n830_));
  AO220      g0808(.A0(new_new_n350_), .A1(new_new_n340_), .B0(new_new_n392_), .B1(new_new_n601_), .Y(new_new_n831_));
  NA3        g0809(.A(new_new_n831_), .B(new_new_n254_), .C(i_7_), .Y(new_new_n832_));
  BUFFER     g0810(.A(new_new_n625_), .Y(new_new_n833_));
  NA3        g0811(.A(new_new_n833_), .B(new_new_n149_), .C(new_new_n70_), .Y(new_new_n834_));
  AO210      g0812(.A0(new_new_n496_), .A1(new_new_n762_), .B0(new_new_n36_), .Y(new_new_n835_));
  NA4        g0813(.A(new_new_n835_), .B(new_new_n834_), .C(new_new_n832_), .D(new_new_n830_), .Y(new_new_n836_));
  NO2        g0814(.A(new_new_n646_), .B(i_11_), .Y(new_new_n837_));
  AOI220     g0815(.A0(new_new_n837_), .A1(new_new_n569_), .B0(new_new_n803_), .B1(new_new_n724_), .Y(new_new_n838_));
  NA3        g0816(.A(new_new_n366_), .B(new_new_n238_), .C(new_new_n149_), .Y(new_new_n839_));
  NA2        g0817(.A(new_new_n392_), .B(new_new_n71_), .Y(new_new_n840_));
  NA4        g0818(.A(new_new_n840_), .B(new_new_n839_), .C(new_new_n838_), .D(new_new_n607_), .Y(new_new_n841_));
  AOI210     g0819(.A0(new_new_n445_), .A1(new_new_n443_), .B0(new_new_n568_), .Y(new_new_n842_));
  NO2        g0820(.A(new_new_n615_), .B(new_new_n104_), .Y(new_new_n843_));
  OAI210     g0821(.A0(new_new_n843_), .A1(new_new_n113_), .B0(new_new_n404_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n242_), .B(new_new_n47_), .Y(new_new_n845_));
  INV        g0823(.A(new_new_n592_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n846_), .B(new_new_n316_), .C(i_7_), .Y(new_new_n847_));
  NA3        g0825(.A(new_new_n847_), .B(new_new_n844_), .C(new_new_n842_), .Y(new_new_n848_));
  NO4        g0826(.A(new_new_n848_), .B(new_new_n841_), .C(new_new_n836_), .D(new_new_n826_), .Y(new_new_n849_));
  NA4        g0827(.A(new_new_n849_), .B(new_new_n812_), .C(new_new_n806_), .D(new_new_n374_), .Y(men3));
  NA2        g0828(.A(i_12_), .B(i_10_), .Y(new_new_n851_));
  NA2        g0829(.A(i_6_), .B(i_7_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n852_), .B(i_0_), .Y(new_new_n853_));
  NO2        g0831(.A(i_11_), .B(new_new_n236_), .Y(new_new_n854_));
  NA3        g0832(.A(new_new_n839_), .B(new_new_n607_), .C(new_new_n365_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n855_), .B(new_new_n40_), .Y(new_new_n856_));
  NOi21      g0834(.An(new_new_n98_), .B(new_new_n771_), .Y(new_new_n857_));
  NO3        g0835(.A(new_new_n634_), .B(new_new_n453_), .C(new_new_n133_), .Y(new_new_n858_));
  AN2        g0836(.A(new_new_n451_), .B(new_new_n56_), .Y(new_new_n859_));
  NO3        g0837(.A(new_new_n859_), .B(new_new_n858_), .C(new_new_n857_), .Y(new_new_n860_));
  AOI210     g0838(.A0(new_new_n860_), .A1(new_new_n856_), .B0(new_new_n49_), .Y(new_new_n861_));
  NO4        g0839(.A(new_new_n370_), .B(new_new_n377_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n862_));
  NA2        g0840(.A(new_new_n185_), .B(new_new_n578_), .Y(new_new_n863_));
  NOi21      g0841(.An(new_new_n863_), .B(new_new_n862_), .Y(new_new_n864_));
  NO2        g0842(.A(new_new_n864_), .B(new_new_n64_), .Y(new_new_n865_));
  NOi21      g0843(.An(i_5_), .B(i_9_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n866_), .B(new_new_n442_), .Y(new_new_n867_));
  BUFFER     g0845(.A(new_new_n266_), .Y(new_new_n868_));
  AOI210     g0846(.A0(new_new_n868_), .A1(new_new_n476_), .B0(new_new_n697_), .Y(new_new_n869_));
  NO3        g0847(.A(new_new_n410_), .B(new_new_n266_), .C(new_new_n74_), .Y(new_new_n870_));
  NO2        g0848(.A(new_new_n178_), .B(new_new_n150_), .Y(new_new_n871_));
  AOI210     g0849(.A0(new_new_n871_), .A1(new_new_n242_), .B0(new_new_n870_), .Y(new_new_n872_));
  OAI220     g0850(.A0(new_new_n872_), .A1(new_new_n183_), .B0(new_new_n869_), .B1(new_new_n867_), .Y(new_new_n873_));
  NO3        g0851(.A(new_new_n873_), .B(new_new_n865_), .C(new_new_n861_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n185_), .B(new_new_n24_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n301_), .B(new_new_n131_), .Y(new_new_n876_));
  NAi21      g0854(.An(new_new_n164_), .B(new_new_n434_), .Y(new_new_n877_));
  OAI220     g0855(.A0(new_new_n877_), .A1(new_new_n845_), .B0(new_new_n876_), .B1(new_new_n395_), .Y(new_new_n878_));
  INV        g0856(.A(new_new_n878_), .Y(new_new_n879_));
  NO2        g0857(.A(new_new_n384_), .B(new_new_n282_), .Y(new_new_n880_));
  NA2        g0858(.A(new_new_n880_), .B(new_new_n720_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n579_), .B(i_0_), .Y(new_new_n882_));
  NO3        g0860(.A(new_new_n882_), .B(new_new_n379_), .C(new_new_n88_), .Y(new_new_n883_));
  NO4        g0861(.A(new_new_n591_), .B(new_new_n217_), .C(new_new_n414_), .D(new_new_n406_), .Y(new_new_n884_));
  AOI210     g0862(.A0(new_new_n884_), .A1(i_11_), .B0(new_new_n883_), .Y(new_new_n885_));
  INV        g0863(.A(new_new_n474_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n758_), .B(new_new_n317_), .Y(new_new_n887_));
  AOI210     g0865(.A0(new_new_n485_), .A1(new_new_n88_), .B0(new_new_n59_), .Y(new_new_n888_));
  NO2        g0866(.A(new_new_n888_), .B(new_new_n887_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n252_), .B(new_new_n155_), .Y(new_new_n890_));
  NA2        g0868(.A(i_0_), .B(i_10_), .Y(new_new_n891_));
  INV        g0869(.A(new_new_n544_), .Y(new_new_n892_));
  NO4        g0870(.A(new_new_n116_), .B(new_new_n59_), .C(new_new_n675_), .D(i_5_), .Y(new_new_n893_));
  AO220      g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n890_), .B1(i_6_), .Y(new_new_n894_));
  AOI220     g0872(.A0(new_new_n323_), .A1(new_new_n100_), .B0(new_new_n185_), .B1(new_new_n85_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n573_), .B(i_4_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n188_), .B(new_new_n203_), .Y(new_new_n897_));
  OAI220     g0875(.A0(new_new_n897_), .A1(new_new_n887_), .B0(new_new_n896_), .B1(new_new_n895_), .Y(new_new_n898_));
  NO3        g0876(.A(new_new_n898_), .B(new_new_n894_), .C(new_new_n889_), .Y(new_new_n899_));
  NA4        g0877(.A(new_new_n899_), .B(new_new_n885_), .C(new_new_n881_), .D(new_new_n879_), .Y(new_new_n900_));
  NO2        g0878(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n901_));
  NA2        g0879(.A(i_11_), .B(i_9_), .Y(new_new_n902_));
  NO3        g0880(.A(i_12_), .B(new_new_n902_), .C(new_new_n606_), .Y(new_new_n903_));
  AN2        g0881(.A(new_new_n903_), .B(new_new_n901_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n49_), .B(i_7_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n389_), .B(new_new_n182_), .Y(new_new_n906_));
  NA2        g0884(.A(new_new_n906_), .B(new_new_n162_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n902_), .B(new_new_n74_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n178_), .B(i_0_), .Y(new_new_n909_));
  INV        g0887(.A(new_new_n909_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n474_), .B(new_new_n231_), .Y(new_new_n911_));
  AOI210     g0889(.A0(new_new_n364_), .A1(new_new_n42_), .B0(new_new_n403_), .Y(new_new_n912_));
  OAI220     g0890(.A0(new_new_n912_), .A1(new_new_n867_), .B0(new_new_n911_), .B1(new_new_n910_), .Y(new_new_n913_));
  NO3        g0891(.A(new_new_n913_), .B(new_new_n907_), .C(new_new_n904_), .Y(new_new_n914_));
  NA2        g0892(.A(new_new_n665_), .B(new_new_n123_), .Y(new_new_n915_));
  NO2        g0893(.A(i_6_), .B(new_new_n915_), .Y(new_new_n916_));
  AOI210     g0894(.A0(new_new_n444_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n917_));
  NA2        g0895(.A(new_new_n174_), .B(new_new_n105_), .Y(new_new_n918_));
  NOi32      g0896(.An(new_new_n917_), .Bn(new_new_n188_), .C(new_new_n918_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n919_), .B(new_new_n916_), .Y(new_new_n920_));
  NOi21      g0898(.An(i_7_), .B(i_5_), .Y(new_new_n921_));
  NOi31      g0899(.An(new_new_n921_), .B(i_0_), .C(new_new_n736_), .Y(new_new_n922_));
  NA3        g0900(.A(new_new_n922_), .B(new_new_n378_), .C(i_6_), .Y(new_new_n923_));
  OA210      g0901(.A0(new_new_n918_), .A1(new_new_n520_), .B0(new_new_n923_), .Y(new_new_n924_));
  NO3        g0902(.A(new_new_n398_), .B(new_new_n353_), .C(new_new_n349_), .Y(new_new_n925_));
  NO2        g0903(.A(new_new_n261_), .B(new_new_n308_), .Y(new_new_n926_));
  NO2        g0904(.A(new_new_n736_), .B(new_new_n256_), .Y(new_new_n927_));
  AOI210     g0905(.A0(new_new_n927_), .A1(new_new_n926_), .B0(new_new_n925_), .Y(new_new_n928_));
  NA4        g0906(.A(new_new_n928_), .B(new_new_n924_), .C(new_new_n920_), .D(new_new_n914_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n875_), .B(new_new_n239_), .Y(new_new_n930_));
  AN2        g0908(.A(new_new_n322_), .B(new_new_n317_), .Y(new_new_n931_));
  AN2        g0909(.A(new_new_n931_), .B(new_new_n871_), .Y(new_new_n932_));
  OAI210     g0910(.A0(new_new_n932_), .A1(new_new_n930_), .B0(i_10_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n851_), .B(new_new_n307_), .Y(new_new_n934_));
  NA2        g0912(.A(new_new_n934_), .B(new_new_n908_), .Y(new_new_n935_));
  NA3        g0913(.A(new_new_n473_), .B(new_new_n407_), .C(new_new_n46_), .Y(new_new_n936_));
  OAI210     g0914(.A0(new_new_n877_), .A1(new_new_n886_), .B0(new_new_n936_), .Y(new_new_n937_));
  NO2        g0915(.A(new_new_n254_), .B(new_new_n47_), .Y(new_new_n938_));
  NA2        g0916(.A(new_new_n908_), .B(new_new_n294_), .Y(new_new_n939_));
  OAI210     g0917(.A0(new_new_n938_), .A1(new_new_n187_), .B0(new_new_n939_), .Y(new_new_n940_));
  AOI220     g0918(.A0(new_new_n940_), .A1(new_new_n474_), .B0(new_new_n937_), .B1(new_new_n74_), .Y(new_new_n941_));
  NA3        g0919(.A(new_new_n828_), .B(new_new_n376_), .C(new_new_n646_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n942_), .B(new_new_n48_), .Y(new_new_n943_));
  NO3        g0921(.A(new_new_n591_), .B(new_new_n348_), .C(new_new_n24_), .Y(new_new_n944_));
  AOI210     g0922(.A0(new_new_n711_), .A1(new_new_n550_), .B0(new_new_n944_), .Y(new_new_n945_));
  NAi21      g0923(.An(i_9_), .B(i_5_), .Y(new_new_n946_));
  NO2        g0924(.A(new_new_n946_), .B(new_new_n398_), .Y(new_new_n947_));
  NA2        g0925(.A(new_new_n947_), .B(new_new_n625_), .Y(new_new_n948_));
  OAI220     g0926(.A0(new_new_n948_), .A1(new_new_n87_), .B0(new_new_n945_), .B1(new_new_n175_), .Y(new_new_n949_));
  NO3        g0927(.A(new_new_n949_), .B(new_new_n943_), .C(new_new_n525_), .Y(new_new_n950_));
  NA4        g0928(.A(new_new_n950_), .B(new_new_n941_), .C(new_new_n935_), .D(new_new_n933_), .Y(new_new_n951_));
  NO3        g0929(.A(new_new_n951_), .B(new_new_n929_), .C(new_new_n900_), .Y(new_new_n952_));
  NO2        g0930(.A(i_0_), .B(new_new_n736_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n954_));
  INV        g0932(.A(new_new_n954_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n107_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n956_));
  AO220      g0934(.A0(new_new_n956_), .A1(new_new_n955_), .B0(new_new_n953_), .B1(new_new_n177_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n808_), .B(new_new_n918_), .Y(new_new_n958_));
  AOI210     g0936(.A0(new_new_n957_), .A1(new_new_n337_), .B0(new_new_n958_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n747_), .B(new_new_n148_), .Y(new_new_n960_));
  INV        g0938(.A(new_new_n960_), .Y(new_new_n961_));
  NA3        g0939(.A(new_new_n961_), .B(new_new_n682_), .C(new_new_n74_), .Y(new_new_n962_));
  OAI210     g0940(.A0(new_new_n242_), .A1(i_9_), .B0(new_new_n230_), .Y(new_new_n963_));
  AOI210     g0941(.A0(new_new_n963_), .A1(new_new_n882_), .B0(new_new_n155_), .Y(new_new_n964_));
  INV        g0942(.A(new_new_n964_), .Y(new_new_n965_));
  NA3        g0943(.A(new_new_n965_), .B(new_new_n962_), .C(new_new_n959_), .Y(new_new_n966_));
  NA2        g0944(.A(new_new_n931_), .B(new_new_n366_), .Y(new_new_n967_));
  AOI210     g0945(.A0(new_new_n289_), .A1(new_new_n164_), .B0(new_new_n967_), .Y(new_new_n968_));
  NA3        g0946(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n905_), .B(new_new_n490_), .Y(new_new_n970_));
  AOI210     g0948(.A0(new_new_n969_), .A1(new_new_n164_), .B0(new_new_n970_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n971_), .B(new_new_n968_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n891_), .B(new_new_n866_), .C(new_new_n190_), .Y(new_new_n973_));
  AOI220     g0951(.A0(new_new_n973_), .A1(i_11_), .B0(new_new_n574_), .B1(new_new_n76_), .Y(new_new_n974_));
  NO3        g0952(.A(new_new_n211_), .B(new_new_n377_), .C(i_0_), .Y(new_new_n975_));
  OAI210     g0953(.A0(new_new_n975_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n976_));
  INV        g0954(.A(new_new_n219_), .Y(new_new_n977_));
  OAI220     g0955(.A0(new_new_n537_), .A1(new_new_n141_), .B0(new_new_n651_), .B1(new_new_n619_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n978_), .B(new_new_n393_), .C(new_new_n977_), .Y(new_new_n979_));
  NA4        g0957(.A(new_new_n979_), .B(new_new_n976_), .C(new_new_n974_), .D(new_new_n972_), .Y(new_new_n980_));
  AOI220     g0958(.A0(new_new_n921_), .A1(new_new_n490_), .B0(new_new_n853_), .B1(new_new_n165_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n340_), .B(new_new_n179_), .Y(new_new_n982_));
  OR2        g0960(.A(new_new_n982_), .B(new_new_n981_), .Y(new_new_n983_));
  NA3        g0961(.A(new_new_n616_), .B(new_new_n185_), .C(new_new_n85_), .Y(new_new_n984_));
  NA2        g0962(.A(new_new_n984_), .B(new_new_n548_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n495_), .B(new_new_n488_), .Y(new_new_n986_));
  NO2        g0964(.A(new_new_n986_), .B(new_new_n985_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n384_), .B(new_new_n174_), .C(new_new_n173_), .Y(new_new_n988_));
  INV        g0966(.A(new_new_n988_), .Y(new_new_n989_));
  NA3        g0967(.A(new_new_n384_), .B(new_new_n324_), .C(new_new_n221_), .Y(new_new_n990_));
  INV        g0968(.A(new_new_n990_), .Y(new_new_n991_));
  NOi31      g0969(.An(new_new_n383_), .B(new_new_n954_), .C(new_new_n239_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n902_), .B(new_new_n219_), .C(new_new_n190_), .Y(new_new_n993_));
  NO4        g0971(.A(new_new_n993_), .B(new_new_n992_), .C(new_new_n991_), .D(new_new_n989_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n994_), .B(new_new_n987_), .C(new_new_n983_), .Y(new_new_n995_));
  INV        g0973(.A(new_new_n618_), .Y(new_new_n996_));
  NO3        g0974(.A(new_new_n996_), .B(new_new_n564_), .C(new_new_n334_), .Y(new_new_n997_));
  NO2        g0975(.A(new_new_n87_), .B(i_5_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n854_), .B(new_new_n111_), .C(new_new_n126_), .Y(new_new_n999_));
  INV        g0977(.A(new_new_n999_), .Y(new_new_n1000_));
  AOI210     g0978(.A0(new_new_n1000_), .A1(new_new_n998_), .B0(new_new_n997_), .Y(new_new_n1001_));
  NA3        g0979(.A(new_new_n294_), .B(i_5_), .C(new_new_n193_), .Y(new_new_n1002_));
  NAi31      g0980(.An(new_new_n240_), .B(new_new_n1002_), .C(new_new_n241_), .Y(new_new_n1003_));
  NO4        g0981(.A(new_new_n239_), .B(new_new_n211_), .C(i_0_), .D(i_12_), .Y(new_new_n1004_));
  AOI220     g0982(.A0(new_new_n1004_), .A1(new_new_n1003_), .B0(new_new_n802_), .B1(new_new_n179_), .Y(new_new_n1005_));
  AN2        g0983(.A(new_new_n891_), .B(new_new_n155_), .Y(new_new_n1006_));
  NO4        g0984(.A(new_new_n1006_), .B(i_12_), .C(new_new_n655_), .D(new_new_n133_), .Y(new_new_n1007_));
  NA2        g0985(.A(new_new_n1007_), .B(new_new_n219_), .Y(new_new_n1008_));
  NA3        g0986(.A(new_new_n100_), .B(new_new_n578_), .C(i_11_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n1009_), .B(new_new_n157_), .Y(new_new_n1010_));
  NA2        g0988(.A(new_new_n921_), .B(new_new_n471_), .Y(new_new_n1011_));
  NA2        g0989(.A(new_new_n65_), .B(new_new_n103_), .Y(new_new_n1012_));
  OAI220     g0990(.A0(new_new_n1012_), .A1(new_new_n1002_), .B0(new_new_n1011_), .B1(new_new_n683_), .Y(new_new_n1013_));
  AOI210     g0991(.A0(new_new_n1013_), .A1(new_new_n909_), .B0(new_new_n1010_), .Y(new_new_n1014_));
  NA4        g0992(.A(new_new_n1014_), .B(new_new_n1008_), .C(new_new_n1005_), .D(new_new_n1001_), .Y(new_new_n1015_));
  NO4        g0993(.A(new_new_n1015_), .B(new_new_n995_), .C(new_new_n980_), .D(new_new_n966_), .Y(new_new_n1016_));
  OAI210     g0994(.A0(new_new_n827_), .A1(new_new_n821_), .B0(new_new_n37_), .Y(new_new_n1017_));
  NA2        g0995(.A(new_new_n1017_), .B(new_new_n614_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n1018_), .B(new_new_n208_), .Y(new_new_n1019_));
  AN2        g0997(.A(new_new_n706_), .B(new_new_n362_), .Y(new_new_n1020_));
  NA2        g0998(.A(new_new_n186_), .B(new_new_n188_), .Y(new_new_n1021_));
  AO210      g0999(.A0(new_new_n1020_), .A1(new_new_n33_), .B0(new_new_n1021_), .Y(new_new_n1022_));
  OAI210     g1000(.A0(new_new_n618_), .A1(new_new_n616_), .B0(new_new_n307_), .Y(new_new_n1023_));
  NAi31      g1001(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1024_));
  AOI210     g1002(.A0(new_new_n119_), .A1(new_new_n71_), .B0(new_new_n1024_), .Y(new_new_n1025_));
  NO2        g1003(.A(new_new_n1025_), .B(new_new_n652_), .Y(new_new_n1026_));
  NA3        g1004(.A(new_new_n1026_), .B(new_new_n1023_), .C(new_new_n1022_), .Y(new_new_n1027_));
  NO2        g1005(.A(new_new_n461_), .B(new_new_n266_), .Y(new_new_n1028_));
  NO4        g1006(.A(new_new_n233_), .B(new_new_n147_), .C(new_new_n686_), .D(new_new_n37_), .Y(new_new_n1029_));
  NO3        g1007(.A(new_new_n1029_), .B(new_new_n1028_), .C(new_new_n884_), .Y(new_new_n1030_));
  OAI210     g1008(.A0(new_new_n1009_), .A1(new_new_n150_), .B0(new_new_n1030_), .Y(new_new_n1031_));
  AOI210     g1009(.A0(new_new_n1027_), .A1(new_new_n49_), .B0(new_new_n1031_), .Y(new_new_n1032_));
  AOI210     g1010(.A0(new_new_n1032_), .A1(new_new_n1019_), .B0(new_new_n74_), .Y(new_new_n1033_));
  NO2        g1011(.A(new_new_n571_), .B(new_new_n373_), .Y(new_new_n1034_));
  NO2        g1012(.A(new_new_n1034_), .B(new_new_n766_), .Y(new_new_n1035_));
  NA3        g1013(.A(new_new_n98_), .B(new_new_n296_), .C(new_new_n31_), .Y(new_new_n1036_));
  NA2        g1014(.A(new_new_n160_), .B(new_new_n88_), .Y(new_new_n1037_));
  NA3        g1015(.A(new_new_n770_), .B(new_new_n278_), .C(new_new_n81_), .Y(new_new_n1038_));
  AOI210     g1016(.A0(new_new_n1038_), .A1(new_new_n1037_), .B0(i_11_), .Y(new_new_n1039_));
  NA2        g1017(.A(new_new_n609_), .B(new_new_n217_), .Y(new_new_n1040_));
  OAI210     g1018(.A0(new_new_n1040_), .A1(new_new_n917_), .B0(new_new_n208_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n166_), .B(i_5_), .Y(new_new_n1042_));
  NO2        g1020(.A(new_new_n1041_), .B(new_new_n1042_), .Y(new_new_n1043_));
  NO3        g1021(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1044_));
  OAI210     g1022(.A0(new_new_n926_), .A1(new_new_n296_), .B0(new_new_n1044_), .Y(new_new_n1045_));
  NO2        g1023(.A(new_new_n1045_), .B(new_new_n736_), .Y(new_new_n1046_));
  NO4        g1024(.A(new_new_n946_), .B(new_new_n478_), .C(new_new_n251_), .D(new_new_n250_), .Y(new_new_n1047_));
  NO2        g1025(.A(new_new_n1047_), .B(new_new_n568_), .Y(new_new_n1048_));
  INV        g1026(.A(new_new_n354_), .Y(new_new_n1049_));
  AOI210     g1027(.A0(new_new_n1049_), .A1(new_new_n1048_), .B0(new_new_n41_), .Y(new_new_n1050_));
  NO4        g1028(.A(new_new_n1050_), .B(new_new_n1046_), .C(new_new_n1043_), .D(new_new_n1039_), .Y(new_new_n1051_));
  OAI210     g1029(.A0(new_new_n1036_), .A1(i_4_), .B0(new_new_n1051_), .Y(new_new_n1052_));
  NO3        g1030(.A(new_new_n1052_), .B(new_new_n1035_), .C(new_new_n1033_), .Y(new_new_n1053_));
  NA4        g1031(.A(new_new_n1053_), .B(new_new_n1016_), .C(new_new_n952_), .D(new_new_n874_), .Y(men4));
  INV        g1032(.A(new_new_n710_), .Y(new_new_n1057_));
  INV        g1033(.A(new_new_n485_), .Y(new_new_n1058_));
endmodule


