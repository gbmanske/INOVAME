//Benchmark atmr_9sym_175_0.25

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, ori00, mai00, men00;
  ONE        o0(.Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  INV        m006(.A(i_4_), .Y(mai_mai_n17_));
  NA2        m007(.A(i_0_), .B(mai_mai_n17_), .Y(mai_mai_n18_));
  INV        m008(.A(i_7_), .Y(mai_mai_n19_));
  NA3        m009(.A(i_6_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n20_));
  NOi21      m010(.An(i_8_), .B(i_6_), .Y(mai_mai_n21_));
  NA2        m011(.A(mai_mai_n21_), .B(i_5_), .Y(mai_mai_n22_));
  AOI210     m012(.A0(mai_mai_n22_), .A1(mai_mai_n20_), .B0(mai_mai_n18_), .Y(mai_mai_n23_));
  NA2        m013(.A(mai_mai_n23_), .B(mai_mai_n11_), .Y(mai_mai_n24_));
  NA2        m014(.A(i_0_), .B(mai_mai_n13_), .Y(mai_mai_n25_));
  NA2        m015(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n26_));
  NO2        m016(.A(i_2_), .B(i_4_), .Y(mai_mai_n27_));
  NA3        m017(.A(mai_mai_n27_), .B(i_6_), .C(i_8_), .Y(mai_mai_n28_));
  AOI210     m018(.A0(mai_mai_n26_), .A1(mai_mai_n25_), .B0(mai_mai_n28_), .Y(mai_mai_n29_));
  INV        m019(.A(i_2_), .Y(mai_mai_n30_));
  NOi21      m020(.An(i_5_), .B(i_0_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_6_), .B(i_8_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_7_), .B(i_1_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_5_), .B(i_6_), .Y(mai_mai_n34_));
  AOI220     m024(.A0(mai_mai_n34_), .A1(mai_mai_n33_), .B0(mai_mai_n32_), .B1(mai_mai_n31_), .Y(mai_mai_n35_));
  NO3        m025(.A(mai_mai_n35_), .B(mai_mai_n30_), .C(i_4_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_0_), .B(i_4_), .Y(mai_mai_n37_));
  XO2        m027(.A(i_1_), .B(i_3_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_7_), .B(i_5_), .Y(mai_mai_n39_));
  AN3        m029(.A(mai_mai_n39_), .B(mai_mai_n38_), .C(mai_mai_n37_), .Y(mai_mai_n40_));
  INV        m030(.A(i_1_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_3_), .B(i_0_), .Y(mai_mai_n42_));
  NA2        m032(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA3        m033(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n44_));
  AOI210     m034(.A0(mai_mai_n44_), .A1(mai_mai_n20_), .B0(mai_mai_n43_), .Y(mai_mai_n45_));
  NO4        m035(.A(mai_mai_n45_), .B(mai_mai_n40_), .C(mai_mai_n36_), .D(mai_mai_n29_), .Y(mai_mai_n46_));
  NOi21      m036(.An(i_4_), .B(i_0_), .Y(mai_mai_n47_));
  AOI210     m037(.A0(mai_mai_n47_), .A1(mai_mai_n21_), .B0(mai_mai_n14_), .Y(mai_mai_n48_));
  NA2        m038(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_2_), .B(i_8_), .Y(mai_mai_n50_));
  NO3        m040(.A(mai_mai_n50_), .B(mai_mai_n47_), .C(mai_mai_n37_), .Y(mai_mai_n51_));
  NO3        m041(.A(mai_mai_n51_), .B(mai_mai_n49_), .C(mai_mai_n48_), .Y(mai_mai_n52_));
  INV        m042(.A(mai_mai_n52_), .Y(mai_mai_n53_));
  NOi31      m043(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n54_));
  NOi21      m044(.An(i_4_), .B(i_3_), .Y(mai_mai_n55_));
  NOi21      m045(.An(i_1_), .B(i_4_), .Y(mai_mai_n56_));
  OAI210     m046(.A0(mai_mai_n56_), .A1(mai_mai_n55_), .B0(mai_mai_n50_), .Y(mai_mai_n57_));
  INV        m047(.A(mai_mai_n57_), .Y(mai_mai_n58_));
  AN2        m048(.A(i_8_), .B(i_7_), .Y(mai_mai_n59_));
  NA2        m049(.A(mai_mai_n59_), .B(mai_mai_n12_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_8_), .B(i_7_), .Y(mai_mai_n61_));
  NA3        m051(.A(mai_mai_n61_), .B(mai_mai_n55_), .C(i_6_), .Y(mai_mai_n62_));
  OAI210     m052(.A0(mai_mai_n60_), .A1(mai_mai_n49_), .B0(mai_mai_n62_), .Y(mai_mai_n63_));
  AOI220     m053(.A0(mai_mai_n63_), .A1(mai_mai_n30_), .B0(mai_mai_n58_), .B1(mai_mai_n34_), .Y(mai_mai_n64_));
  NA4        m054(.A(mai_mai_n64_), .B(mai_mai_n53_), .C(mai_mai_n46_), .D(mai_mai_n24_), .Y(mai_mai_n65_));
  NA2        m055(.A(i_8_), .B(mai_mai_n19_), .Y(mai_mai_n66_));
  AOI220     m056(.A0(mai_mai_n42_), .A1(i_1_), .B0(mai_mai_n38_), .B1(i_2_), .Y(mai_mai_n67_));
  NOi21      m057(.An(i_1_), .B(i_2_), .Y(mai_mai_n68_));
  NA3        m058(.A(mai_mai_n68_), .B(mai_mai_n47_), .C(i_6_), .Y(mai_mai_n69_));
  OAI210     m059(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n69_), .Y(mai_mai_n70_));
  NA2        m060(.A(mai_mai_n70_), .B(mai_mai_n13_), .Y(mai_mai_n71_));
  NA3        m061(.A(mai_mai_n61_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n72_));
  INV        m062(.A(mai_mai_n72_), .Y(mai_mai_n73_));
  NA2        m063(.A(mai_mai_n73_), .B(mai_mai_n55_), .Y(mai_mai_n74_));
  NA2        m064(.A(mai_mai_n74_), .B(mai_mai_n71_), .Y(mai_mai_n75_));
  NA2        m065(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n76_));
  NOi21      m066(.An(i_7_), .B(i_8_), .Y(mai_mai_n77_));
  NA2        m067(.A(mai_mai_n77_), .B(mai_mai_n12_), .Y(mai_mai_n78_));
  OAI210     m068(.A0(mai_mai_n78_), .A1(mai_mai_n11_), .B0(mai_mai_n76_), .Y(mai_mai_n79_));
  NA2        m069(.A(mai_mai_n79_), .B(mai_mai_n68_), .Y(mai_mai_n80_));
  AOI220     m070(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n16_), .B1(mai_mai_n30_), .Y(mai_mai_n81_));
  NA3        m071(.A(mai_mai_n17_), .B(i_5_), .C(i_7_), .Y(mai_mai_n82_));
  NO2        m072(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n83_));
  INV        m073(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  NAi21      m074(.An(i_6_), .B(i_0_), .Y(mai_mai_n85_));
  NA3        m075(.A(mai_mai_n56_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n86_));
  NOi21      m076(.An(i_4_), .B(i_6_), .Y(mai_mai_n87_));
  NOi21      m077(.An(i_5_), .B(i_3_), .Y(mai_mai_n88_));
  NA3        m078(.A(mai_mai_n88_), .B(mai_mai_n68_), .C(mai_mai_n87_), .Y(mai_mai_n89_));
  OAI210     m079(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n68_), .B(mai_mai_n32_), .Y(mai_mai_n91_));
  NOi21      m081(.An(mai_mai_n39_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  NO2        m082(.A(mai_mai_n92_), .B(mai_mai_n90_), .Y(mai_mai_n93_));
  NOi21      m083(.An(i_6_), .B(i_1_), .Y(mai_mai_n94_));
  AOI220     m084(.A0(mai_mai_n94_), .A1(i_7_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n95_));
  NOi31      m085(.An(mai_mai_n47_), .B(mai_mai_n95_), .C(i_2_), .Y(mai_mai_n96_));
  INV        m086(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NA4        m087(.A(mai_mai_n97_), .B(mai_mai_n93_), .C(mai_mai_n84_), .D(mai_mai_n80_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n50_), .B(mai_mai_n14_), .Y(mai_mai_n99_));
  NA3        m089(.A(mai_mai_n32_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n100_));
  NA3        m090(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(mai_mai_n91_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n101_), .B(mai_mai_n37_), .Y(mai_mai_n102_));
  NA2        m092(.A(mai_mai_n55_), .B(mai_mai_n33_), .Y(mai_mai_n103_));
  AOI210     m093(.A0(mai_mai_n103_), .A1(mai_mai_n72_), .B0(mai_mai_n26_), .Y(mai_mai_n104_));
  NA3        m094(.A(mai_mai_n61_), .B(mai_mai_n54_), .C(i_6_), .Y(mai_mai_n105_));
  INV        m095(.A(mai_mai_n105_), .Y(mai_mai_n106_));
  NOi21      m096(.An(i_0_), .B(i_2_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n107_), .B(mai_mai_n33_), .C(mai_mai_n87_), .Y(mai_mai_n108_));
  NA3        m098(.A(mai_mai_n47_), .B(mai_mai_n39_), .C(mai_mai_n16_), .Y(mai_mai_n109_));
  NA3        m099(.A(mai_mai_n107_), .B(mai_mai_n55_), .C(mai_mai_n32_), .Y(mai_mai_n110_));
  NA3        m100(.A(mai_mai_n110_), .B(mai_mai_n109_), .C(mai_mai_n108_), .Y(mai_mai_n111_));
  NA4        m101(.A(mai_mai_n54_), .B(i_6_), .C(mai_mai_n13_), .D(i_7_), .Y(mai_mai_n112_));
  INV        m102(.A(mai_mai_n112_), .Y(mai_mai_n113_));
  NO4        m103(.A(mai_mai_n113_), .B(mai_mai_n111_), .C(mai_mai_n106_), .D(mai_mai_n104_), .Y(mai_mai_n114_));
  NA2        m104(.A(mai_mai_n77_), .B(mai_mai_n12_), .Y(mai_mai_n115_));
  NA3        m105(.A(i_2_), .B(i_1_), .C(mai_mai_n13_), .Y(mai_mai_n116_));
  NA2        m106(.A(mai_mai_n47_), .B(i_3_), .Y(mai_mai_n117_));
  AOI210     m107(.A0(mai_mai_n117_), .A1(mai_mai_n116_), .B0(mai_mai_n115_), .Y(mai_mai_n118_));
  NA3        m108(.A(mai_mai_n107_), .B(mai_mai_n61_), .C(mai_mai_n87_), .Y(mai_mai_n119_));
  INV        m109(.A(mai_mai_n119_), .Y(mai_mai_n120_));
  NA4        m110(.A(mai_mai_n88_), .B(mai_mai_n59_), .C(mai_mai_n41_), .D(mai_mai_n17_), .Y(mai_mai_n121_));
  NA3        m111(.A(mai_mai_n50_), .B(mai_mai_n31_), .C(mai_mai_n14_), .Y(mai_mai_n122_));
  NA2        m112(.A(mai_mai_n122_), .B(mai_mai_n121_), .Y(mai_mai_n123_));
  NO3        m113(.A(mai_mai_n123_), .B(mai_mai_n120_), .C(mai_mai_n118_), .Y(mai_mai_n124_));
  NA3        m114(.A(mai_mai_n124_), .B(mai_mai_n114_), .C(mai_mai_n102_), .Y(mai_mai_n125_));
  OR4        m115(.A(mai_mai_n125_), .B(mai_mai_n98_), .C(mai_mai_n75_), .D(mai_mai_n65_), .Y(mai00));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  NOi21      u014(.An(i_1_), .B(i_8_), .Y(men_men_n25_));
  AOI220     u015(.A0(men_men_n25_), .A1(i_2_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n26_));
  NO2        u016(.A(men_men_n26_), .B(men_men_n22_), .Y(men_men_n27_));
  AOI210     u017(.A0(men_men_n27_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n28_));
  NA2        u018(.A(i_0_), .B(men_men_n14_), .Y(men_men_n29_));
  NA2        u019(.A(men_men_n17_), .B(i_5_), .Y(men_men_n30_));
  NO2        u020(.A(i_2_), .B(i_4_), .Y(men_men_n31_));
  INV        u021(.A(i_2_), .Y(men_men_n32_));
  NOi21      u022(.An(i_6_), .B(i_8_), .Y(men_men_n33_));
  NOi21      u023(.An(i_5_), .B(i_6_), .Y(men_men_n34_));
  NOi21      u024(.An(i_0_), .B(i_4_), .Y(men_men_n35_));
  INV        u025(.A(i_1_), .Y(men_men_n36_));
  NOi21      u026(.An(i_3_), .B(i_0_), .Y(men_men_n37_));
  INV        u027(.A(i_8_), .Y(men_men_n38_));
  NA2        u028(.A(i_1_), .B(men_men_n11_), .Y(men_men_n39_));
  NO4        u029(.A(men_men_n39_), .B(men_men_n29_), .C(i_2_), .D(men_men_n38_), .Y(men_men_n40_));
  NOi21      u030(.An(i_4_), .B(i_0_), .Y(men_men_n41_));
  NOi21      u031(.An(i_2_), .B(i_8_), .Y(men_men_n42_));
  INV        u032(.A(men_men_n40_), .Y(men_men_n43_));
  NOi31      u033(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n44_));
  NA2        u034(.A(men_men_n44_), .B(i_0_), .Y(men_men_n45_));
  NOi21      u035(.An(i_4_), .B(i_3_), .Y(men_men_n46_));
  NOi21      u036(.An(i_1_), .B(i_4_), .Y(men_men_n47_));
  OAI210     u037(.A0(men_men_n47_), .A1(men_men_n46_), .B0(men_men_n42_), .Y(men_men_n48_));
  NA2        u038(.A(men_men_n48_), .B(men_men_n45_), .Y(men_men_n49_));
  AN2        u039(.A(i_8_), .B(i_7_), .Y(men_men_n50_));
  NOi21      u040(.An(i_8_), .B(i_7_), .Y(men_men_n51_));
  NA2        u041(.A(men_men_n49_), .B(men_men_n34_), .Y(men_men_n52_));
  NA3        u042(.A(men_men_n52_), .B(men_men_n43_), .C(men_men_n28_), .Y(men_men_n53_));
  NA2        u043(.A(i_8_), .B(i_7_), .Y(men_men_n54_));
  NO3        u044(.A(men_men_n54_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n55_));
  NOi21      u045(.An(i_1_), .B(i_2_), .Y(men_men_n56_));
  NA2        u046(.A(men_men_n55_), .B(men_men_n14_), .Y(men_men_n57_));
  NA3        u047(.A(men_men_n25_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n58_));
  INV        u048(.A(men_men_n58_), .Y(men_men_n59_));
  NOi32      u049(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(i_3_), .Y(men_men_n61_));
  NA3        u051(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n62_));
  NA2        u052(.A(men_men_n62_), .B(men_men_n61_), .Y(men_men_n63_));
  NO2        u053(.A(i_0_), .B(i_4_), .Y(men_men_n64_));
  AOI220     u054(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n59_), .B1(men_men_n46_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(men_men_n57_), .Y(men_men_n66_));
  NAi21      u056(.An(i_3_), .B(i_6_), .Y(men_men_n67_));
  NO3        u057(.A(men_men_n67_), .B(i_0_), .C(men_men_n38_), .Y(men_men_n68_));
  NOi21      u058(.An(i_7_), .B(i_8_), .Y(men_men_n69_));
  NOi31      u059(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n70_));
  AOI210     u060(.A0(men_men_n69_), .A1(men_men_n12_), .B0(men_men_n70_), .Y(men_men_n71_));
  NO2        u061(.A(men_men_n71_), .B(men_men_n11_), .Y(men_men_n72_));
  OAI210     u062(.A0(men_men_n72_), .A1(men_men_n68_), .B0(men_men_n56_), .Y(men_men_n73_));
  NA3        u063(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n74_));
  AOI210     u064(.A0(men_men_n22_), .A1(men_men_n39_), .B0(men_men_n74_), .Y(men_men_n75_));
  OAI210     u065(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n76_));
  NA3        u066(.A(men_men_n54_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n77_));
  NO2        u067(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NO2        u068(.A(men_men_n78_), .B(men_men_n75_), .Y(men_men_n79_));
  NA3        u069(.A(men_men_n51_), .B(men_men_n32_), .C(i_3_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n36_), .B(i_6_), .Y(men_men_n81_));
  AOI210     u071(.A0(men_men_n81_), .A1(men_men_n22_), .B0(men_men_n80_), .Y(men_men_n82_));
  NOi21      u072(.An(i_2_), .B(i_1_), .Y(men_men_n83_));
  AN3        u073(.A(men_men_n69_), .B(men_men_n83_), .C(men_men_n41_), .Y(men_men_n84_));
  NAi21      u074(.An(i_6_), .B(i_0_), .Y(men_men_n85_));
  NOi21      u075(.An(i_4_), .B(i_6_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n56_), .B(men_men_n33_), .Y(men_men_n87_));
  NO2        u077(.A(men_men_n84_), .B(men_men_n82_), .Y(men_men_n88_));
  NA2        u078(.A(men_men_n51_), .B(men_men_n12_), .Y(men_men_n89_));
  NA2        u079(.A(men_men_n33_), .B(men_men_n14_), .Y(men_men_n90_));
  NOi21      u080(.An(i_3_), .B(i_1_), .Y(men_men_n91_));
  NA2        u081(.A(men_men_n91_), .B(i_4_), .Y(men_men_n92_));
  AOI210     u082(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n92_), .Y(men_men_n93_));
  AOI220     u083(.A0(men_men_n69_), .A1(men_men_n14_), .B0(men_men_n86_), .B1(men_men_n23_), .Y(men_men_n94_));
  NOi31      u084(.An(men_men_n37_), .B(men_men_n94_), .C(men_men_n32_), .Y(men_men_n95_));
  NO2        u085(.A(men_men_n95_), .B(men_men_n93_), .Y(men_men_n96_));
  NA4        u086(.A(men_men_n96_), .B(men_men_n88_), .C(men_men_n79_), .D(men_men_n73_), .Y(men_men_n97_));
  NA2        u087(.A(men_men_n42_), .B(men_men_n15_), .Y(men_men_n98_));
  NOi31      u088(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n99_));
  NOi31      u089(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n100_));
  OAI210     u090(.A0(men_men_n100_), .A1(men_men_n99_), .B0(i_7_), .Y(men_men_n101_));
  NA3        u091(.A(men_men_n101_), .B(men_men_n98_), .C(men_men_n87_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n102_), .B(men_men_n35_), .Y(men_men_n103_));
  NA4        u093(.A(men_men_n50_), .B(men_men_n83_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n104_));
  NAi31      u094(.An(men_men_n85_), .B(men_men_n69_), .C(men_men_n83_), .Y(men_men_n105_));
  NA3        u095(.A(men_men_n51_), .B(men_men_n44_), .C(i_6_), .Y(men_men_n106_));
  NA3        u096(.A(men_men_n106_), .B(men_men_n105_), .C(men_men_n104_), .Y(men_men_n107_));
  NOi32      u097(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n108_));
  NA2        u098(.A(men_men_n108_), .B(men_men_n99_), .Y(men_men_n109_));
  INV        u099(.A(men_men_n109_), .Y(men_men_n110_));
  NA4        u100(.A(men_men_n47_), .B(men_men_n34_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n111_));
  NA4        u101(.A(men_men_n47_), .B(men_men_n37_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n112_));
  NA2        u102(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NO3        u103(.A(men_men_n113_), .B(men_men_n110_), .C(men_men_n107_), .Y(men_men_n114_));
  NOi21      u104(.An(i_5_), .B(i_2_), .Y(men_men_n115_));
  AOI220     u105(.A0(men_men_n115_), .A1(men_men_n69_), .B0(men_men_n50_), .B1(men_men_n31_), .Y(men_men_n116_));
  AOI210     u106(.A0(men_men_n116_), .A1(men_men_n98_), .B0(men_men_n81_), .Y(men_men_n117_));
  NO4        u107(.A(i_2_), .B(men_men_n21_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n118_));
  NA2        u108(.A(i_2_), .B(i_4_), .Y(men_men_n119_));
  AOI210     u109(.A0(men_men_n85_), .A1(men_men_n67_), .B0(men_men_n119_), .Y(men_men_n120_));
  NO2        u110(.A(i_8_), .B(i_7_), .Y(men_men_n121_));
  OA210      u111(.A0(men_men_n120_), .A1(men_men_n118_), .B0(men_men_n121_), .Y(men_men_n122_));
  NA4        u112(.A(men_men_n91_), .B(i_0_), .C(i_5_), .D(men_men_n23_), .Y(men_men_n123_));
  NO2        u113(.A(men_men_n123_), .B(i_4_), .Y(men_men_n124_));
  NO3        u114(.A(men_men_n124_), .B(men_men_n122_), .C(men_men_n117_), .Y(men_men_n125_));
  NO2        u115(.A(men_men_n80_), .B(men_men_n30_), .Y(men_men_n126_));
  NA3        u116(.A(men_men_n70_), .B(men_men_n91_), .C(i_0_), .Y(men_men_n127_));
  NOi31      u117(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n128_));
  OAI210     u118(.A0(men_men_n108_), .A1(men_men_n60_), .B0(men_men_n128_), .Y(men_men_n129_));
  NA2        u119(.A(men_men_n129_), .B(men_men_n127_), .Y(men_men_n130_));
  NO2        u120(.A(men_men_n130_), .B(men_men_n126_), .Y(men_men_n131_));
  NA4        u121(.A(men_men_n131_), .B(men_men_n125_), .C(men_men_n114_), .D(men_men_n103_), .Y(men_men_n132_));
  OR4        u122(.A(men_men_n132_), .B(men_men_n97_), .C(men_men_n66_), .D(men_men_n53_), .Y(men00));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule