// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n121_, new_new_n122_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n548_, new_new_n549_, new_new_n550_,
    new_new_n551_, new_new_n552_, new_new_n553_, new_new_n554_,
    new_new_n555_, new_new_n556_, new_new_n557_, new_new_n558_,
    new_new_n559_, new_new_n560_, new_new_n561_, new_new_n562_,
    new_new_n563_, new_new_n564_, new_new_n565_, new_new_n566_,
    new_new_n567_, new_new_n568_, new_new_n569_, new_new_n570_,
    new_new_n571_, new_new_n572_, new_new_n573_, new_new_n574_,
    new_new_n575_, new_new_n576_, new_new_n577_, new_new_n578_,
    new_new_n579_, new_new_n580_, new_new_n581_, new_new_n582_,
    new_new_n583_, new_new_n584_, new_new_n585_, new_new_n586_,
    new_new_n588_, new_new_n589_, new_new_n590_, new_new_n591_,
    new_new_n592_, new_new_n593_, new_new_n594_, new_new_n595_,
    new_new_n596_, new_new_n597_, new_new_n598_, new_new_n599_,
    new_new_n600_, new_new_n601_, new_new_n602_, new_new_n603_,
    new_new_n604_, new_new_n605_, new_new_n606_, new_new_n607_,
    new_new_n608_, new_new_n609_, new_new_n610_, new_new_n611_,
    new_new_n612_, new_new_n613_, new_new_n614_, new_new_n615_,
    new_new_n616_, new_new_n617_, new_new_n618_, new_new_n619_,
    new_new_n620_, new_new_n621_, new_new_n622_, new_new_n623_,
    new_new_n624_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(mai1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  OAI210     g027(.A0(new_new_n49_), .A1(i_3_), .B0(new_new_n47_), .Y(new_new_n50_));
  AOI210     g028(.A0(new_new_n50_), .A1(new_new_n46_), .B0(new_new_n45_), .Y(new_new_n51_));
  NA2        g029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NO2        g031(.A(new_new_n53_), .B(new_new_n52_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n51_), .B(new_new_n44_), .Y(new_new_n55_));
  NA3        g033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  OAI210     g036(.A0(new_new_n58_), .A1(new_new_n57_), .B0(new_new_n56_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g039(.A(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n61_), .B(new_new_n31_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n64_), .B(new_new_n60_), .Y(new_new_n65_));
  NA2        g043(.A(new_new_n49_), .B(i_2_), .Y(new_new_n66_));
  AOI210     g044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n67_));
  NA2        g045(.A(i_1_), .B(i_6_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n25_), .Y(new_new_n69_));
  INV        g047(.A(i_0_), .Y(new_new_n70_));
  NAi21      g048(.An(i_5_), .B(i_10_), .Y(new_new_n71_));
  NA2        g049(.A(i_5_), .B(i_9_), .Y(new_new_n72_));
  AOI210     g050(.A0(new_new_n72_), .A1(new_new_n71_), .B0(new_new_n70_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n69_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n74_), .Y(new_new_n75_));
  OAI210     g053(.A0(new_new_n75_), .A1(new_new_n65_), .B0(i_0_), .Y(new_new_n76_));
  NA2        g054(.A(i_12_), .B(i_5_), .Y(new_new_n77_));
  NO2        g055(.A(i_3_), .B(i_9_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n78_), .B(new_new_n62_), .Y(new_new_n80_));
  INV        g058(.A(i_6_), .Y(new_new_n81_));
  NA2        g059(.A(new_new_n80_), .B(i_2_), .Y(new_new_n82_));
  NAi21      g060(.An(i_6_), .B(i_10_), .Y(new_new_n83_));
  NA2        g061(.A(i_6_), .B(i_9_), .Y(new_new_n84_));
  AOI210     g062(.A0(new_new_n84_), .A1(new_new_n83_), .B0(new_new_n62_), .Y(new_new_n85_));
  NA2        g063(.A(i_2_), .B(i_6_), .Y(new_new_n86_));
  NO3        g064(.A(new_new_n86_), .B(new_new_n48_), .C(new_new_n25_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n87_), .B(new_new_n85_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n88_), .A1(new_new_n82_), .B0(new_new_n77_), .Y(new_new_n89_));
  NAi21      g067(.An(i_6_), .B(i_11_), .Y(new_new_n90_));
  INV        g068(.A(i_7_), .Y(new_new_n91_));
  NO2        g069(.A(i_0_), .B(i_5_), .Y(new_new_n92_));
  NAi21      g070(.An(i_7_), .B(i_11_), .Y(new_new_n93_));
  NO3        g071(.A(new_new_n93_), .B(new_new_n83_), .C(new_new_n52_), .Y(new_new_n94_));
  AN2        g072(.A(i_2_), .B(i_10_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(i_7_), .Y(new_new_n96_));
  OR2        g074(.A(new_new_n77_), .B(new_new_n57_), .Y(new_new_n97_));
  NO3        g075(.A(i_7_), .B(new_new_n97_), .C(new_new_n96_), .Y(new_new_n98_));
  NA2        g076(.A(i_12_), .B(i_7_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n100_), .B(i_0_), .Y(new_new_n101_));
  NA2        g079(.A(i_11_), .B(i_12_), .Y(new_new_n102_));
  OAI210     g080(.A0(new_new_n101_), .A1(new_new_n99_), .B0(new_new_n102_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n103_), .B(new_new_n98_), .Y(new_new_n104_));
  NAi21      g082(.An(new_new_n94_), .B(new_new_n104_), .Y(new_new_n105_));
  NOi21      g083(.An(i_1_), .B(i_5_), .Y(new_new_n106_));
  NA2        g084(.A(new_new_n106_), .B(i_11_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n91_), .B(new_new_n37_), .Y(new_new_n108_));
  NA2        g086(.A(i_7_), .B(new_new_n25_), .Y(new_new_n109_));
  NA2        g087(.A(new_new_n109_), .B(new_new_n108_), .Y(new_new_n110_));
  NO2        g088(.A(new_new_n110_), .B(new_new_n45_), .Y(new_new_n111_));
  NA2        g089(.A(new_new_n84_), .B(new_new_n83_), .Y(new_new_n112_));
  NAi21      g090(.An(i_3_), .B(i_8_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n113_), .B(new_new_n61_), .Y(new_new_n114_));
  NOi31      g092(.An(new_new_n114_), .B(new_new_n112_), .C(new_new_n111_), .Y(new_new_n115_));
  NO2        g093(.A(i_1_), .B(new_new_n81_), .Y(new_new_n116_));
  NO2        g094(.A(i_6_), .B(i_5_), .Y(new_new_n117_));
  OAI220     g095(.A0(new_new_n46_), .A1(new_new_n93_), .B0(new_new_n115_), .B1(new_new_n107_), .Y(new_new_n118_));
  NO3        g096(.A(new_new_n118_), .B(new_new_n105_), .C(new_new_n89_), .Y(new_new_n119_));
  NA3        g097(.A(new_new_n119_), .B(new_new_n76_), .C(new_new_n55_), .Y(mai2));
  NO2        g098(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n773_), .B(new_new_n121_), .Y(new_new_n122_));
  NA4        g100(.A(new_new_n122_), .B(new_new_n74_), .C(new_new_n66_), .D(new_new_n30_), .Y(mai0));
  AN2        g101(.A(i_8_), .B(i_7_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(i_6_), .Y(new_new_n125_));
  NO2        g103(.A(i_12_), .B(i_13_), .Y(new_new_n126_));
  NAi21      g104(.An(i_5_), .B(i_11_), .Y(new_new_n127_));
  NOi21      g105(.An(new_new_n126_), .B(new_new_n127_), .Y(new_new_n128_));
  NO2        g106(.A(i_0_), .B(i_1_), .Y(new_new_n129_));
  NA2        g107(.A(i_2_), .B(i_3_), .Y(new_new_n130_));
  NO2        g108(.A(new_new_n130_), .B(i_4_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(new_new_n128_), .Y(new_new_n132_));
  AN2        g110(.A(new_new_n126_), .B(new_new_n78_), .Y(new_new_n133_));
  NA2        g111(.A(i_1_), .B(i_5_), .Y(new_new_n134_));
  NO3        g112(.A(new_new_n778_), .B(new_new_n134_), .C(new_new_n26_), .Y(new_new_n135_));
  OR2        g113(.A(i_0_), .B(i_1_), .Y(new_new_n136_));
  NO3        g114(.A(new_new_n136_), .B(new_new_n77_), .C(i_13_), .Y(new_new_n137_));
  NAi32      g115(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n138_));
  NAi21      g116(.An(new_new_n138_), .B(new_new_n137_), .Y(new_new_n139_));
  NOi21      g117(.An(i_4_), .B(i_10_), .Y(new_new_n140_));
  NA2        g118(.A(new_new_n140_), .B(new_new_n39_), .Y(new_new_n141_));
  NO2        g119(.A(i_3_), .B(i_5_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n137_), .B(new_new_n135_), .Y(new_new_n143_));
  AOI210     g121(.A0(new_new_n143_), .A1(new_new_n132_), .B0(new_new_n125_), .Y(new_new_n144_));
  NOi21      g122(.An(i_4_), .B(i_9_), .Y(new_new_n145_));
  NOi21      g123(.An(i_11_), .B(i_13_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(new_new_n145_), .Y(new_new_n147_));
  NO2        g125(.A(i_4_), .B(i_5_), .Y(new_new_n148_));
  NAi21      g126(.An(i_12_), .B(i_11_), .Y(new_new_n149_));
  NO2        g127(.A(new_new_n149_), .B(i_13_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n70_), .B(new_new_n62_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n36_), .B(i_5_), .Y(new_new_n152_));
  NAi31      g130(.An(new_new_n152_), .B(new_new_n133_), .C(i_11_), .Y(new_new_n153_));
  NA2        g131(.A(i_3_), .B(i_5_), .Y(new_new_n154_));
  AOI210     g132(.A0(new_new_n147_), .A1(new_new_n153_), .B0(new_new_n62_), .Y(new_new_n155_));
  NO2        g133(.A(new_new_n70_), .B(i_5_), .Y(new_new_n156_));
  NO2        g134(.A(i_13_), .B(i_10_), .Y(new_new_n157_));
  NA3        g135(.A(new_new_n157_), .B(new_new_n156_), .C(new_new_n43_), .Y(new_new_n158_));
  NO2        g136(.A(i_2_), .B(i_1_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n159_), .B(i_3_), .Y(new_new_n160_));
  NAi21      g138(.An(i_4_), .B(i_12_), .Y(new_new_n161_));
  NO3        g139(.A(new_new_n161_), .B(new_new_n158_), .C(new_new_n25_), .Y(new_new_n162_));
  NO2        g140(.A(new_new_n162_), .B(new_new_n155_), .Y(new_new_n163_));
  INV        g141(.A(i_8_), .Y(new_new_n164_));
  NA2        g142(.A(i_8_), .B(i_6_), .Y(new_new_n165_));
  NO3        g143(.A(i_3_), .B(new_new_n81_), .C(new_new_n47_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(i_7_), .Y(new_new_n167_));
  NO3        g145(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n168_));
  NA3        g146(.A(new_new_n168_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n169_));
  NO3        g147(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n169_), .B(new_new_n167_), .Y(new_new_n171_));
  NO3        g149(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n172_));
  NA2        g150(.A(new_new_n172_), .B(new_new_n39_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n92_), .B(new_new_n57_), .Y(new_new_n174_));
  NO2        g152(.A(i_13_), .B(i_9_), .Y(new_new_n175_));
  NA3        g153(.A(new_new_n175_), .B(i_6_), .C(new_new_n164_), .Y(new_new_n176_));
  NAi21      g154(.An(i_12_), .B(i_3_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n43_), .B(i_5_), .Y(new_new_n178_));
  OAI210     g156(.A0(new_new_n57_), .A1(new_new_n173_), .B0(new_new_n176_), .Y(new_new_n179_));
  AOI210     g157(.A0(new_new_n179_), .A1(i_7_), .B0(new_new_n171_), .Y(new_new_n180_));
  OAI220     g158(.A0(new_new_n180_), .A1(i_4_), .B0(new_new_n165_), .B1(new_new_n163_), .Y(new_new_n181_));
  NAi21      g159(.An(i_12_), .B(i_7_), .Y(new_new_n182_));
  NA3        g160(.A(i_13_), .B(new_new_n164_), .C(i_10_), .Y(new_new_n183_));
  NO2        g161(.A(new_new_n183_), .B(new_new_n182_), .Y(new_new_n184_));
  NA2        g162(.A(i_0_), .B(i_5_), .Y(new_new_n185_));
  INV        g163(.A(new_new_n160_), .Y(new_new_n186_));
  NAi31      g164(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n45_), .B(new_new_n62_), .Y(new_new_n188_));
  INV        g166(.A(i_13_), .Y(new_new_n189_));
  NO2        g167(.A(i_12_), .B(new_new_n189_), .Y(new_new_n190_));
  NA2        g168(.A(new_new_n190_), .B(new_new_n166_), .Y(new_new_n191_));
  INV        g169(.A(new_new_n191_), .Y(new_new_n192_));
  AOI220     g170(.A0(new_new_n192_), .A1(new_new_n124_), .B0(new_new_n186_), .B1(new_new_n184_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n154_), .B(i_4_), .Y(new_new_n194_));
  NA2        g172(.A(new_new_n194_), .B(i_10_), .Y(new_new_n195_));
  OR2        g173(.A(i_8_), .B(i_7_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n52_), .B(i_1_), .Y(new_new_n197_));
  INV        g175(.A(i_12_), .Y(new_new_n198_));
  NO3        g176(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n199_));
  NA2        g177(.A(i_2_), .B(i_1_), .Y(new_new_n200_));
  NO3        g178(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n201_));
  NAi21      g179(.An(i_4_), .B(i_3_), .Y(new_new_n202_));
  NO2        g180(.A(i_0_), .B(i_6_), .Y(new_new_n203_));
  NOi41      g181(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n204_));
  NO2        g182(.A(i_11_), .B(new_new_n189_), .Y(new_new_n205_));
  NAi21      g183(.An(i_3_), .B(i_7_), .Y(new_new_n206_));
  NA2        g184(.A(new_new_n198_), .B(i_9_), .Y(new_new_n207_));
  OR3        g185(.A(new_new_n207_), .B(new_new_n206_), .C(i_1_), .Y(new_new_n208_));
  NO2        g186(.A(i_12_), .B(i_3_), .Y(new_new_n209_));
  INV        g187(.A(new_new_n208_), .Y(new_new_n210_));
  NA2        g188(.A(new_new_n210_), .B(new_new_n205_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n196_), .B(new_new_n37_), .Y(new_new_n212_));
  NA2        g190(.A(i_12_), .B(i_6_), .Y(new_new_n213_));
  OR2        g191(.A(i_13_), .B(i_9_), .Y(new_new_n214_));
  NO3        g192(.A(new_new_n214_), .B(new_new_n213_), .C(new_new_n47_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n202_), .B(i_2_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n205_), .B(i_9_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n62_), .B(new_new_n217_), .Y(new_new_n218_));
  NA2        g196(.A(i_2_), .B(new_new_n62_), .Y(new_new_n219_));
  NO3        g197(.A(i_11_), .B(new_new_n189_), .C(new_new_n25_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n206_), .B(i_8_), .Y(new_new_n221_));
  NA2        g199(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n222_));
  NA3        g200(.A(i_3_), .B(new_new_n212_), .C(new_new_n190_), .Y(new_new_n223_));
  AOI210     g201(.A0(new_new_n223_), .A1(new_new_n222_), .B0(new_new_n219_), .Y(new_new_n224_));
  AOI210     g202(.A0(new_new_n218_), .A1(new_new_n212_), .B0(new_new_n224_), .Y(new_new_n225_));
  NA3        g203(.A(new_new_n225_), .B(new_new_n211_), .C(new_new_n193_), .Y(new_new_n226_));
  NO3        g204(.A(i_12_), .B(new_new_n189_), .C(new_new_n37_), .Y(new_new_n227_));
  INV        g205(.A(new_new_n227_), .Y(new_new_n228_));
  INV        g206(.A(i_8_), .Y(new_new_n229_));
  NO3        g207(.A(i_0_), .B(new_new_n45_), .C(i_1_), .Y(new_new_n230_));
  AOI220     g208(.A0(new_new_n230_), .A1(new_new_n166_), .B0(new_new_n142_), .B1(new_new_n197_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n231_), .B(new_new_n229_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n200_), .B(i_0_), .Y(new_new_n233_));
  NO2        g211(.A(i_6_), .B(i_0_), .Y(new_new_n234_));
  NA2        g212(.A(i_0_), .B(i_1_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n235_), .B(i_2_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n58_), .B(i_6_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  OAI210     g216(.A0(i_3_), .A1(new_new_n125_), .B0(new_new_n238_), .Y(new_new_n239_));
  NO3        g217(.A(new_new_n239_), .B(new_new_n234_), .C(new_new_n232_), .Y(new_new_n240_));
  NO2        g218(.A(i_3_), .B(i_10_), .Y(new_new_n241_));
  NA3        g219(.A(new_new_n241_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n242_));
  NA2        g220(.A(i_1_), .B(i_7_), .Y(new_new_n243_));
  AN2        g221(.A(i_3_), .B(i_10_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n150_), .B(new_new_n148_), .Y(new_new_n245_));
  OR2        g223(.A(new_new_n243_), .B(new_new_n242_), .Y(new_new_n246_));
  OAI220     g224(.A0(new_new_n246_), .A1(i_6_), .B0(new_new_n240_), .B1(new_new_n228_), .Y(new_new_n247_));
  NO4        g225(.A(new_new_n247_), .B(new_new_n226_), .C(new_new_n181_), .D(new_new_n144_), .Y(new_new_n248_));
  NO3        g226(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n249_));
  NO3        g227(.A(i_6_), .B(new_new_n164_), .C(i_7_), .Y(new_new_n250_));
  NO2        g228(.A(i_2_), .B(i_3_), .Y(new_new_n251_));
  OR2        g229(.A(i_0_), .B(i_5_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n185_), .B(new_new_n252_), .Y(new_new_n253_));
  NA3        g231(.A(new_new_n771_), .B(new_new_n251_), .C(i_1_), .Y(new_new_n254_));
  INV        g232(.A(i_6_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n136_), .B(new_new_n45_), .Y(new_new_n256_));
  INV        g234(.A(new_new_n256_), .Y(new_new_n257_));
  NA3        g235(.A(new_new_n257_), .B(new_new_n200_), .C(new_new_n254_), .Y(new_new_n258_));
  OAI210     g236(.A0(new_new_n258_), .A1(new_new_n250_), .B0(i_4_), .Y(new_new_n259_));
  NO2        g237(.A(i_12_), .B(i_10_), .Y(new_new_n260_));
  NOi21      g238(.An(i_5_), .B(i_0_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n769_), .B(new_new_n113_), .Y(new_new_n262_));
  INV        g240(.A(new_new_n262_), .Y(new_new_n263_));
  NO2        g241(.A(i_6_), .B(i_8_), .Y(new_new_n264_));
  NO2        g242(.A(i_1_), .B(i_7_), .Y(new_new_n265_));
  NA3        g243(.A(new_new_n264_), .B(i_4_), .C(i_5_), .Y(new_new_n266_));
  NA3        g244(.A(new_new_n266_), .B(new_new_n263_), .C(new_new_n259_), .Y(new_new_n267_));
  OAI210     g245(.A0(i_7_), .A1(i_2_), .B0(i_6_), .Y(new_new_n268_));
  NA2        g246(.A(i_0_), .B(new_new_n117_), .Y(new_new_n269_));
  AOI210     g247(.A0(new_new_n164_), .A1(new_new_n253_), .B0(new_new_n141_), .Y(new_new_n270_));
  AOI210     g248(.A0(new_new_n267_), .A1(new_new_n249_), .B0(new_new_n270_), .Y(new_new_n271_));
  NOi32      g249(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n272_));
  INV        g250(.A(new_new_n272_), .Y(new_new_n273_));
  NAi21      g251(.An(i_1_), .B(i_5_), .Y(new_new_n274_));
  NA2        g252(.A(new_new_n274_), .B(i_0_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n275_), .B(new_new_n25_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(new_new_n138_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n138_), .B(new_new_n136_), .Y(new_new_n278_));
  NOi32      g256(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n279_), .B(new_new_n45_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(i_0_), .Y(new_new_n281_));
  OR2        g259(.A(new_new_n281_), .B(new_new_n278_), .Y(new_new_n282_));
  NO2        g260(.A(i_1_), .B(new_new_n91_), .Y(new_new_n283_));
  NAi21      g261(.An(i_3_), .B(i_4_), .Y(new_new_n284_));
  NO2        g262(.A(new_new_n284_), .B(i_9_), .Y(new_new_n285_));
  NA2        g263(.A(i_7_), .B(new_new_n285_), .Y(new_new_n286_));
  NA2        g264(.A(i_2_), .B(i_7_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n284_), .B(i_10_), .Y(new_new_n288_));
  NA3        g266(.A(new_new_n288_), .B(new_new_n287_), .C(new_new_n203_), .Y(new_new_n289_));
  AOI210     g267(.A0(new_new_n289_), .A1(new_new_n286_), .B0(new_new_n156_), .Y(new_new_n290_));
  AOI210     g268(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n291_));
  OAI210     g269(.A0(new_new_n291_), .A1(new_new_n159_), .B0(new_new_n288_), .Y(new_new_n292_));
  AOI220     g270(.A0(new_new_n288_), .A1(new_new_n265_), .B0(new_new_n199_), .B1(new_new_n159_), .Y(new_new_n293_));
  AOI210     g271(.A0(new_new_n293_), .A1(new_new_n292_), .B0(i_5_), .Y(new_new_n294_));
  NO4        g272(.A(new_new_n294_), .B(new_new_n290_), .C(new_new_n282_), .D(new_new_n277_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n295_), .B(new_new_n273_), .Y(new_new_n296_));
  AN2        g274(.A(i_12_), .B(i_5_), .Y(new_new_n297_));
  NA2        g275(.A(i_3_), .B(new_new_n297_), .Y(new_new_n298_));
  NO2        g276(.A(i_11_), .B(i_6_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n136_), .B(new_new_n298_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n202_), .B(i_5_), .Y(new_new_n301_));
  NO2        g279(.A(i_5_), .B(i_10_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n300_), .B(i_9_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n304_));
  NO3        g282(.A(new_new_n81_), .B(new_new_n47_), .C(i_9_), .Y(new_new_n305_));
  NO2        g283(.A(i_11_), .B(i_12_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n302_), .B(new_new_n198_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n91_), .B(new_new_n187_), .Y(new_new_n308_));
  NO2        g286(.A(i_13_), .B(new_new_n200_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n308_), .B(new_new_n309_), .Y(new_new_n310_));
  NA3        g288(.A(new_new_n310_), .B(new_new_n132_), .C(new_new_n303_), .Y(new_new_n311_));
  NO2        g289(.A(i_0_), .B(i_11_), .Y(new_new_n312_));
  AN2        g290(.A(i_1_), .B(i_6_), .Y(new_new_n313_));
  OR2        g291(.A(i_13_), .B(i_10_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n147_), .B(new_new_n108_), .Y(new_new_n315_));
  BUFFER     g293(.A(new_new_n183_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n91_), .B(new_new_n25_), .Y(new_new_n317_));
  NA2        g295(.A(new_new_n227_), .B(new_new_n317_), .Y(new_new_n318_));
  OAI220     g296(.A0(i_6_), .A1(new_new_n316_), .B0(new_new_n318_), .B1(new_new_n92_), .Y(new_new_n319_));
  INV        g297(.A(new_new_n319_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(new_new_n26_), .Y(new_new_n321_));
  INV        g299(.A(new_new_n254_), .Y(new_new_n322_));
  AOI220     g300(.A0(new_new_n237_), .A1(new_new_n230_), .B0(new_new_n233_), .B1(i_7_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n323_), .B(i_5_), .Y(new_new_n324_));
  NO2        g302(.A(i_2_), .B(new_new_n229_), .Y(new_new_n325_));
  NO3        g303(.A(new_new_n325_), .B(new_new_n324_), .C(new_new_n322_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n166_), .B(i_1_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(i_8_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n63_), .B(i_2_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n237_), .B(new_new_n197_), .Y(new_new_n330_));
  OAI220     g308(.A0(new_new_n330_), .A1(new_new_n154_), .B0(new_new_n329_), .B1(new_new_n774_), .Y(new_new_n331_));
  NA3        g309(.A(new_new_n265_), .B(new_new_n264_), .C(i_5_), .Y(new_new_n332_));
  INV        g310(.A(new_new_n332_), .Y(new_new_n333_));
  NO3        g311(.A(new_new_n333_), .B(new_new_n331_), .C(new_new_n328_), .Y(new_new_n334_));
  AOI210     g312(.A0(new_new_n334_), .A1(new_new_n326_), .B0(new_new_n217_), .Y(new_new_n335_));
  NO4        g313(.A(new_new_n335_), .B(new_new_n321_), .C(new_new_n311_), .D(new_new_n296_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n70_), .B(i_13_), .Y(new_new_n337_));
  NO2        g315(.A(i_10_), .B(i_9_), .Y(new_new_n338_));
  NAi21      g316(.An(i_12_), .B(i_8_), .Y(new_new_n339_));
  NO2        g317(.A(new_new_n339_), .B(i_3_), .Y(new_new_n340_));
  NO3        g318(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n213_), .B(new_new_n90_), .Y(new_new_n342_));
  NA2        g320(.A(i_8_), .B(i_9_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n227_), .B(new_new_n174_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n344_), .B(new_new_n343_), .Y(new_new_n345_));
  NO3        g323(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n346_));
  NA3        g324(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n100_), .B(new_new_n23_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n347_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(new_new_n345_), .Y(new_new_n350_));
  OR2        g328(.A(new_new_n176_), .B(new_new_n195_), .Y(new_new_n351_));
  NO2        g329(.A(i_2_), .B(i_13_), .Y(new_new_n352_));
  NO3        g330(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n353_));
  NO2        g331(.A(i_6_), .B(i_7_), .Y(new_new_n354_));
  NO2        g332(.A(i_11_), .B(i_1_), .Y(new_new_n355_));
  NAi31      g333(.An(i_11_), .B(i_2_), .C(i_0_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n314_), .B(i_6_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n357_), .B(i_1_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n358_), .B(new_new_n356_), .Y(new_new_n359_));
  NO2        g337(.A(i_6_), .B(i_10_), .Y(new_new_n360_));
  INV        g338(.A(new_new_n359_), .Y(new_new_n361_));
  NAi21      g339(.An(new_new_n183_), .B(new_new_n306_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n265_), .B(new_new_n185_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n26_), .B(i_5_), .Y(new_new_n364_));
  NA3        g342(.A(i_6_), .B(new_new_n364_), .C(new_new_n124_), .Y(new_new_n365_));
  OR3        g343(.A(new_new_n769_), .B(new_new_n38_), .C(new_new_n45_), .Y(new_new_n366_));
  OAI220     g344(.A0(new_new_n366_), .A1(new_new_n365_), .B0(new_new_n363_), .B1(new_new_n362_), .Y(new_new_n367_));
  NA2        g345(.A(new_new_n249_), .B(new_new_n199_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n368_), .B(new_new_n329_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(new_new_n367_), .Y(new_new_n370_));
  NA4        g348(.A(new_new_n370_), .B(new_new_n361_), .C(new_new_n351_), .D(new_new_n350_), .Y(new_new_n371_));
  AN2        g349(.A(i_5_), .B(new_new_n341_), .Y(new_new_n372_));
  OAI210     g350(.A0(new_new_n70_), .A1(new_new_n195_), .B0(new_new_n245_), .Y(new_new_n373_));
  AOI220     g351(.A0(new_new_n373_), .A1(new_new_n255_), .B0(new_new_n372_), .B1(i_3_), .Y(new_new_n374_));
  NA3        g352(.A(new_new_n337_), .B(i_1_), .C(i_2_), .Y(new_new_n375_));
  INV        g353(.A(new_new_n375_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n297_), .B(new_new_n189_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n272_), .B(new_new_n70_), .Y(new_new_n378_));
  NA2        g356(.A(i_7_), .B(new_new_n279_), .Y(new_new_n379_));
  AO210      g357(.A0(new_new_n378_), .A1(new_new_n377_), .B0(new_new_n379_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n36_), .B(i_8_), .Y(new_new_n381_));
  NAi41      g359(.An(new_new_n378_), .B(new_new_n360_), .C(new_new_n381_), .D(new_new_n45_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n382_), .B(new_new_n380_), .Y(new_new_n383_));
  AOI210     g361(.A0(new_new_n376_), .A1(new_new_n172_), .B0(new_new_n383_), .Y(new_new_n384_));
  NO2        g362(.A(i_7_), .B(new_new_n169_), .Y(new_new_n385_));
  AOI220     g363(.A0(i_3_), .A1(new_new_n385_), .B0(new_new_n766_), .B1(new_new_n315_), .Y(new_new_n386_));
  NA3        g364(.A(new_new_n386_), .B(new_new_n384_), .C(new_new_n374_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n301_), .B(new_new_n236_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n298_), .B(new_new_n388_), .Y(new_new_n389_));
  NO2        g367(.A(i_12_), .B(new_new_n164_), .Y(new_new_n390_));
  OAI210     g368(.A0(new_new_n250_), .A1(new_new_n390_), .B0(new_new_n389_), .Y(new_new_n391_));
  NO2        g369(.A(i_8_), .B(i_7_), .Y(new_new_n392_));
  INV        g370(.A(new_new_n188_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n43_), .B(i_10_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n394_), .B(i_6_), .Y(new_new_n395_));
  NA3        g373(.A(new_new_n395_), .B(i_3_), .C(new_new_n392_), .Y(new_new_n396_));
  NA2        g374(.A(i_5_), .B(new_new_n203_), .Y(new_new_n397_));
  INV        g375(.A(new_new_n397_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n398_), .B(new_new_n212_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n242_), .B(new_new_n152_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n244_), .B(new_new_n148_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n780_), .B(new_new_n251_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n402_), .B(new_new_n401_), .Y(new_new_n403_));
  OAI210     g381(.A0(new_new_n403_), .A1(new_new_n400_), .B0(new_new_n346_), .Y(new_new_n404_));
  NA4        g382(.A(new_new_n404_), .B(new_new_n399_), .C(new_new_n396_), .D(new_new_n391_), .Y(new_new_n405_));
  NA3        g383(.A(new_new_n185_), .B(new_new_n68_), .C(new_new_n43_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n227_), .B(new_new_n79_), .Y(new_new_n407_));
  AOI210     g385(.A0(new_new_n406_), .A1(new_new_n269_), .B0(new_new_n407_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n390_), .B(new_new_n220_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n91_), .B(new_new_n409_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n410_), .B(new_new_n408_), .Y(new_new_n411_));
  NO4        g389(.A(i_1_), .B(new_new_n41_), .C(i_2_), .D(new_new_n47_), .Y(new_new_n412_));
  NO3        g390(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n196_), .B(new_new_n36_), .Y(new_new_n414_));
  AN2        g392(.A(new_new_n414_), .B(new_new_n413_), .Y(new_new_n415_));
  OA210      g393(.A0(new_new_n415_), .A1(new_new_n412_), .B0(new_new_n272_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n314_), .B(i_1_), .Y(new_new_n417_));
  NOi31      g395(.An(new_new_n417_), .B(new_new_n342_), .C(new_new_n70_), .Y(new_new_n418_));
  AN4        g396(.A(new_new_n418_), .B(new_new_n124_), .C(new_new_n364_), .D(i_2_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n419_), .B(new_new_n416_), .Y(new_new_n420_));
  NOi21      g398(.An(i_10_), .B(i_6_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n99_), .B(new_new_n23_), .Y(new_new_n422_));
  INV        g400(.A(new_new_n250_), .Y(new_new_n423_));
  AOI220     g401(.A0(new_new_n423_), .A1(new_new_n330_), .B0(new_new_n147_), .B1(new_new_n153_), .Y(new_new_n424_));
  INV        g402(.A(new_new_n424_), .Y(new_new_n425_));
  INV        g403(.A(new_new_n251_), .Y(new_new_n426_));
  NO2        g404(.A(i_12_), .B(new_new_n81_), .Y(new_new_n427_));
  NA2        g405(.A(new_new_n427_), .B(new_new_n220_), .Y(new_new_n428_));
  NA3        g406(.A(new_new_n299_), .B(new_new_n227_), .C(new_new_n185_), .Y(new_new_n429_));
  AOI210     g407(.A0(new_new_n429_), .A1(new_new_n428_), .B0(new_new_n426_), .Y(new_new_n430_));
  NO3        g408(.A(i_4_), .B(new_new_n268_), .C(new_new_n242_), .Y(new_new_n431_));
  OR2        g409(.A(i_5_), .B(new_new_n313_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n432_), .B(new_new_n362_), .Y(new_new_n433_));
  NO3        g411(.A(new_new_n433_), .B(new_new_n431_), .C(new_new_n430_), .Y(new_new_n434_));
  NA4        g412(.A(new_new_n434_), .B(new_new_n425_), .C(new_new_n420_), .D(new_new_n411_), .Y(new_new_n435_));
  NO4        g413(.A(new_new_n435_), .B(new_new_n405_), .C(new_new_n387_), .D(new_new_n371_), .Y(new_new_n436_));
  NA4        g414(.A(new_new_n436_), .B(new_new_n336_), .C(new_new_n271_), .D(new_new_n248_), .Y(mai7));
  NO2        g415(.A(new_new_n93_), .B(new_new_n83_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n360_), .B(new_new_n79_), .Y(new_new_n439_));
  NA2        g417(.A(i_11_), .B(new_new_n164_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n198_), .B(i_4_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n441_), .B(i_8_), .Y(new_new_n442_));
  INV        g420(.A(i_2_), .Y(new_new_n443_));
  INV        g421(.A(new_new_n172_), .Y(new_new_n444_));
  NO2        g422(.A(i_7_), .B(new_new_n37_), .Y(new_new_n445_));
  NA2        g423(.A(i_4_), .B(i_8_), .Y(new_new_n446_));
  INV        g424(.A(new_new_n438_), .Y(new_new_n447_));
  OR2        g425(.A(i_6_), .B(i_10_), .Y(new_new_n448_));
  NO2        g426(.A(new_new_n448_), .B(new_new_n23_), .Y(new_new_n449_));
  OR3        g427(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n450_));
  NO3        g428(.A(new_new_n450_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n451_));
  INV        g429(.A(new_new_n170_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n451_), .B(new_new_n449_), .Y(new_new_n453_));
  OA220      g431(.A0(new_new_n453_), .A1(new_new_n426_), .B0(new_new_n764_), .B1(new_new_n214_), .Y(new_new_n454_));
  AOI210     g432(.A0(new_new_n454_), .A1(new_new_n447_), .B0(new_new_n62_), .Y(new_new_n455_));
  NOi21      g433(.An(i_11_), .B(i_7_), .Y(new_new_n456_));
  AO210      g434(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n457_), .B(new_new_n456_), .Y(new_new_n458_));
  NA3        g436(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n459_));
  NAi31      g437(.An(new_new_n459_), .B(new_new_n182_), .C(i_11_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n460_), .B(new_new_n62_), .Y(new_new_n461_));
  AO210      g439(.A0(i_8_), .A1(new_new_n293_), .B0(new_new_n40_), .Y(new_new_n462_));
  NO3        g440(.A(i_7_), .B(new_new_n177_), .C(new_new_n440_), .Y(new_new_n463_));
  OAI210     g441(.A0(new_new_n463_), .A1(new_new_n190_), .B0(new_new_n62_), .Y(new_new_n464_));
  NA2        g442(.A(i_2_), .B(new_new_n31_), .Y(new_new_n465_));
  OR2        g443(.A(new_new_n177_), .B(new_new_n93_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n466_), .B(new_new_n465_), .Y(new_new_n467_));
  INV        g445(.A(i_4_), .Y(new_new_n468_));
  NA2        g446(.A(new_new_n468_), .B(new_new_n467_), .Y(new_new_n469_));
  NO2        g447(.A(i_1_), .B(i_12_), .Y(new_new_n470_));
  NA3        g448(.A(new_new_n470_), .B(new_new_n95_), .C(new_new_n24_), .Y(new_new_n471_));
  NA4        g449(.A(new_new_n471_), .B(new_new_n469_), .C(new_new_n464_), .D(new_new_n462_), .Y(new_new_n472_));
  OAI210     g450(.A0(new_new_n472_), .A1(new_new_n461_), .B0(i_6_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n459_), .B(new_new_n93_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n474_), .B(new_new_n427_), .Y(new_new_n475_));
  NO2        g453(.A(i_6_), .B(i_11_), .Y(new_new_n476_));
  INV        g454(.A(new_new_n475_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n392_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n478_));
  NA2        g456(.A(new_new_n121_), .B(i_9_), .Y(new_new_n479_));
  NA3        g457(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n480_));
  NA3        g458(.A(i_2_), .B(new_new_n213_), .C(new_new_n43_), .Y(new_new_n481_));
  OAI220     g459(.A0(new_new_n481_), .A1(new_new_n480_), .B0(new_new_n479_), .B1(new_new_n763_), .Y(new_new_n482_));
  AOI210     g460(.A0(new_new_n355_), .A1(new_new_n317_), .B0(new_new_n201_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n443_), .Y(new_new_n484_));
  NO2        g462(.A(i_11_), .B(new_new_n37_), .Y(new_new_n485_));
  NA2        g463(.A(new_new_n485_), .B(new_new_n24_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n486_), .B(new_new_n45_), .Y(new_new_n487_));
  OR3        g465(.A(new_new_n487_), .B(new_new_n484_), .C(new_new_n482_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n488_), .B(new_new_n477_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n198_), .B(new_new_n91_), .Y(new_new_n490_));
  NO2        g468(.A(new_new_n490_), .B(new_new_n456_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n491_), .B(i_1_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n492_), .B(new_new_n450_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n45_), .Y(new_new_n494_));
  NA2        g472(.A(i_3_), .B(new_new_n164_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n495_), .B(new_new_n99_), .Y(new_new_n496_));
  AN2        g474(.A(new_new_n496_), .B(new_new_n395_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n81_), .B(i_9_), .Y(new_new_n498_));
  NA2        g476(.A(i_1_), .B(i_3_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n86_), .B(new_new_n499_), .Y(new_new_n500_));
  NO2        g478(.A(new_new_n500_), .B(new_new_n497_), .Y(new_new_n501_));
  NA4        g479(.A(new_new_n501_), .B(new_new_n494_), .C(new_new_n489_), .D(new_new_n473_), .Y(new_new_n502_));
  NO3        g480(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n503_));
  OR2        g481(.A(new_new_n503_), .B(new_new_n204_), .Y(new_new_n504_));
  NA3        g482(.A(new_new_n360_), .B(new_new_n381_), .C(new_new_n45_), .Y(new_new_n505_));
  NA2        g483(.A(i_6_), .B(new_new_n25_), .Y(new_new_n506_));
  NA2        g484(.A(new_new_n506_), .B(new_new_n505_), .Y(new_new_n507_));
  OAI210     g485(.A0(new_new_n507_), .A1(new_new_n504_), .B0(i_1_), .Y(new_new_n508_));
  AOI210     g486(.A0(new_new_n213_), .A1(new_new_n90_), .B0(i_1_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n284_), .B(i_2_), .Y(new_new_n510_));
  NA2        g488(.A(new_new_n510_), .B(new_new_n509_), .Y(new_new_n511_));
  AOI210     g489(.A0(new_new_n511_), .A1(new_new_n508_), .B0(i_13_), .Y(new_new_n512_));
  NA2        g490(.A(i_12_), .B(new_new_n121_), .Y(new_new_n513_));
  AOI220     g491(.A0(new_new_n352_), .A1(new_new_n140_), .B0(i_2_), .B1(new_new_n121_), .Y(new_new_n514_));
  OAI210     g492(.A0(new_new_n514_), .A1(new_new_n43_), .B0(new_new_n513_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n53_), .B(new_new_n86_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n515_), .A1(new_new_n264_), .B0(new_new_n516_), .Y(new_new_n517_));
  AOI220     g495(.A0(i_12_), .A1(new_new_n69_), .B0(new_new_n299_), .B1(i_2_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(new_new_n202_), .Y(new_new_n519_));
  AOI210     g497(.A0(new_new_n339_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n520_));
  NOi31      g498(.An(new_new_n520_), .B(new_new_n439_), .C(new_new_n43_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n112_), .B(i_13_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n480_), .B(new_new_n99_), .Y(new_new_n523_));
  INV        g501(.A(new_new_n523_), .Y(new_new_n524_));
  OAI220     g502(.A0(new_new_n524_), .A1(new_new_n68_), .B0(new_new_n522_), .B1(new_new_n509_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n198_), .B(new_new_n81_), .Y(new_new_n526_));
  INV        g504(.A(new_new_n526_), .Y(new_new_n527_));
  AOI210     g505(.A0(new_new_n299_), .A1(i_2_), .B0(new_new_n85_), .Y(new_new_n528_));
  OAI220     g506(.A0(new_new_n528_), .A1(new_new_n442_), .B0(new_new_n527_), .B1(new_new_n452_), .Y(new_new_n529_));
  NO4        g507(.A(new_new_n529_), .B(new_new_n525_), .C(new_new_n521_), .D(new_new_n519_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n524_), .B(i_11_), .Y(new_new_n531_));
  NA2        g509(.A(i_2_), .B(new_new_n445_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n476_), .B(i_13_), .Y(new_new_n533_));
  NAi21      g511(.An(i_11_), .B(i_12_), .Y(new_new_n534_));
  NOi41      g512(.An(new_new_n96_), .B(new_new_n534_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n427_), .B(new_new_n446_), .Y(new_new_n536_));
  AOI210     g514(.A0(new_new_n536_), .A1(new_new_n249_), .B0(new_new_n535_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n537_), .B(new_new_n533_), .C(new_new_n532_), .Y(new_new_n538_));
  OAI210     g516(.A0(new_new_n538_), .A1(new_new_n531_), .B0(new_new_n62_), .Y(new_new_n539_));
  NO3        g517(.A(i_9_), .B(i_3_), .C(new_new_n441_), .Y(new_new_n540_));
  NA2        g518(.A(new_new_n540_), .B(new_new_n283_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n113_), .B(i_2_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n542_), .B(new_new_n470_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n543_), .B(new_new_n541_), .Y(new_new_n544_));
  NA3        g522(.A(new_new_n544_), .B(new_new_n44_), .C(new_new_n189_), .Y(new_new_n545_));
  NA4        g523(.A(new_new_n545_), .B(new_new_n539_), .C(new_new_n530_), .D(new_new_n517_), .Y(new_new_n546_));
  OR4        g524(.A(new_new_n546_), .B(new_new_n512_), .C(new_new_n502_), .D(new_new_n455_), .Y(mai5));
  NA2        g525(.A(new_new_n491_), .B(new_new_n216_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n442_), .B(i_11_), .Y(new_new_n549_));
  INV        g527(.A(new_new_n549_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n550_), .B(new_new_n548_), .Y(new_new_n551_));
  NO3        g529(.A(i_11_), .B(new_new_n198_), .C(i_13_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n553_));
  NA2        g531(.A(i_12_), .B(i_8_), .Y(new_new_n554_));
  NA2        g532(.A(i_12_), .B(new_new_n553_), .Y(new_new_n555_));
  INV        g533(.A(new_new_n555_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n556_), .B(new_new_n551_), .Y(new_new_n557_));
  INV        g535(.A(new_new_n146_), .Y(new_new_n558_));
  INV        g536(.A(new_new_n204_), .Y(new_new_n559_));
  OAI210     g537(.A0(new_new_n510_), .A1(new_new_n340_), .B0(new_new_n96_), .Y(new_new_n560_));
  AOI210     g538(.A0(new_new_n560_), .A1(new_new_n559_), .B0(new_new_n558_), .Y(new_new_n561_));
  INV        g539(.A(new_new_n317_), .Y(new_new_n562_));
  NA2        g540(.A(new_new_n562_), .B(i_2_), .Y(new_new_n563_));
  INV        g541(.A(new_new_n563_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n314_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n565_), .A1(new_new_n564_), .B0(new_new_n561_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n161_), .B(new_new_n110_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n567_), .B(i_2_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n568_), .B(new_new_n164_), .Y(new_new_n569_));
  OA210      g547(.A0(new_new_n458_), .A1(new_new_n111_), .B0(i_13_), .Y(new_new_n570_));
  INV        g548(.A(new_new_n170_), .Y(new_new_n571_));
  INV        g549(.A(new_new_n133_), .Y(new_new_n572_));
  AOI210     g550(.A0(new_new_n572_), .A1(new_new_n571_), .B0(new_new_n287_), .Y(new_new_n573_));
  AOI210     g551(.A0(new_new_n177_), .A1(new_new_n130_), .B0(new_new_n381_), .Y(new_new_n574_));
  NA2        g552(.A(new_new_n574_), .B(new_new_n317_), .Y(new_new_n575_));
  NO2        g553(.A(i_2_), .B(new_new_n43_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n244_), .B(new_new_n41_), .Y(new_new_n577_));
  OAI210     g555(.A0(new_new_n577_), .A1(new_new_n576_), .B0(new_new_n575_), .Y(new_new_n578_));
  NO4        g556(.A(new_new_n578_), .B(new_new_n573_), .C(new_new_n570_), .D(new_new_n569_), .Y(new_new_n579_));
  INV        g557(.A(new_new_n422_), .Y(new_new_n580_));
  NA2        g558(.A(new_new_n552_), .B(new_new_n221_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n581_), .B(new_new_n580_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n61_), .B(i_12_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n583_), .B(new_new_n111_), .Y(new_new_n584_));
  NO2        g562(.A(new_new_n584_), .B(new_new_n440_), .Y(new_new_n585_));
  AOI220     g563(.A0(new_new_n585_), .A1(new_new_n36_), .B0(new_new_n582_), .B1(new_new_n45_), .Y(new_new_n586_));
  NA4        g564(.A(new_new_n586_), .B(new_new_n579_), .C(new_new_n566_), .D(new_new_n557_), .Y(mai6));
  NA2        g565(.A(new_new_n25_), .B(new_new_n542_), .Y(new_new_n588_));
  NA3        g566(.A(new_new_n302_), .B(i_8_), .C(new_new_n68_), .Y(new_new_n589_));
  INV        g567(.A(new_new_n589_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n187_), .B(i_2_), .Y(new_new_n591_));
  INV        g569(.A(i_9_), .Y(new_new_n592_));
  NO2        g570(.A(new_new_n590_), .B(new_new_n261_), .Y(new_new_n593_));
  AO210      g571(.A0(new_new_n593_), .A1(new_new_n588_), .B0(i_12_), .Y(new_new_n594_));
  NA2        g572(.A(new_new_n288_), .B(new_new_n265_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n427_), .B(new_new_n62_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n596_), .B(new_new_n595_), .Y(new_new_n597_));
  INV        g575(.A(new_new_n167_), .Y(new_new_n598_));
  AOI220     g576(.A0(new_new_n598_), .A1(new_new_n592_), .B0(new_new_n597_), .B1(new_new_n70_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n767_), .B(new_new_n583_), .Y(new_new_n600_));
  AOI210     g578(.A0(new_new_n600_), .A1(new_new_n379_), .B0(new_new_n156_), .Y(new_new_n601_));
  NA3        g579(.A(new_new_n770_), .B(new_new_n354_), .C(new_new_n302_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n414_), .B(new_new_n413_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n603_), .B(new_new_n602_), .Y(new_new_n604_));
  OR2        g582(.A(new_new_n604_), .B(new_new_n601_), .Y(new_new_n605_));
  NO2        g583(.A(i_11_), .B(i_2_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n47_), .B(new_new_n37_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n607_), .B(new_new_n313_), .Y(new_new_n608_));
  NA2        g586(.A(new_new_n608_), .B(new_new_n606_), .Y(new_new_n609_));
  NA3        g587(.A(new_new_n772_), .B(new_new_n209_), .C(i_7_), .Y(new_new_n610_));
  BUFFER     g588(.A(new_new_n340_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n611_), .B(new_new_n129_), .Y(new_new_n612_));
  NA3        g590(.A(new_new_n612_), .B(new_new_n610_), .C(new_new_n609_), .Y(new_new_n613_));
  AOI210     g591(.A0(new_new_n765_), .A1(new_new_n413_), .B0(new_new_n591_), .Y(new_new_n614_));
  NA2        g592(.A(new_new_n199_), .B(new_new_n129_), .Y(new_new_n615_));
  OAI210     g593(.A0(new_new_n305_), .A1(new_new_n172_), .B0(new_new_n67_), .Y(new_new_n616_));
  NA4        g594(.A(new_new_n616_), .B(new_new_n615_), .C(new_new_n614_), .D(new_new_n444_), .Y(new_new_n617_));
  NA3        g595(.A(new_new_n381_), .B(new_new_n360_), .C(new_new_n185_), .Y(new_new_n618_));
  AOI210     g596(.A0(new_new_n340_), .A1(new_new_n338_), .B0(new_new_n412_), .Y(new_new_n619_));
  INV        g597(.A(new_new_n312_), .Y(new_new_n620_));
  INV        g598(.A(new_new_n432_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n621_), .B(new_new_n260_), .C(i_7_), .Y(new_new_n622_));
  NA4        g600(.A(new_new_n622_), .B(new_new_n620_), .C(new_new_n619_), .D(new_new_n618_), .Y(new_new_n623_));
  NO4        g601(.A(new_new_n623_), .B(new_new_n617_), .C(new_new_n613_), .D(new_new_n605_), .Y(new_new_n624_));
  NA4        g602(.A(new_new_n624_), .B(new_new_n599_), .C(new_new_n594_), .D(new_new_n295_), .Y(mai3));
  NA2        g603(.A(i_12_), .B(i_10_), .Y(new_new_n626_));
  NO2        g604(.A(i_11_), .B(new_new_n198_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n233_), .B(new_new_n627_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n164_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n83_), .B(new_new_n43_), .Y(new_new_n630_));
  OA210      g608(.A0(new_new_n630_), .A1(new_new_n629_), .B0(new_new_n148_), .Y(new_new_n631_));
  NO3        g609(.A(new_new_n466_), .B(new_new_n343_), .C(new_new_n116_), .Y(new_new_n632_));
  NA2        g610(.A(i_2_), .B(new_new_n44_), .Y(new_new_n633_));
  AN2        g611(.A(new_new_n342_), .B(new_new_n54_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n634_), .B(new_new_n632_), .Y(new_new_n635_));
  INV        g613(.A(new_new_n635_), .Y(new_new_n636_));
  NO3        g614(.A(new_new_n291_), .B(new_new_n38_), .C(i_0_), .Y(new_new_n637_));
  NO2        g615(.A(new_new_n779_), .B(new_new_n62_), .Y(new_new_n638_));
  NOi21      g616(.An(i_5_), .B(i_9_), .Y(new_new_n639_));
  NA2        g617(.A(new_new_n639_), .B(new_new_n337_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n149_), .B(new_new_n130_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(new_new_n203_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n642_), .B(new_new_n152_), .Y(new_new_n643_));
  NO4        g621(.A(new_new_n643_), .B(new_new_n638_), .C(new_new_n636_), .D(new_new_n631_), .Y(new_new_n644_));
  NA2        g622(.A(new_new_n156_), .B(new_new_n24_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n102_), .B(new_new_n645_), .Y(new_new_n646_));
  NA2        g624(.A(new_new_n249_), .B(new_new_n114_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n647_), .B(new_new_n307_), .Y(new_new_n648_));
  NO2        g626(.A(new_new_n648_), .B(new_new_n646_), .Y(new_new_n649_));
  NA2        g627(.A(i_6_), .B(i_0_), .Y(new_new_n650_));
  NO4        g628(.A(i_5_), .B(new_new_n182_), .C(new_new_n314_), .D(new_new_n313_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n651_), .B(i_11_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n552_), .B(new_new_n261_), .Y(new_new_n653_));
  OAI220     g631(.A0(i_6_), .A1(new_new_n653_), .B0(new_new_n486_), .B1(new_new_n393_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n207_), .B(new_new_n134_), .Y(new_new_n655_));
  NA2        g633(.A(i_0_), .B(i_10_), .Y(new_new_n656_));
  NO4        g634(.A(new_new_n99_), .B(new_new_n57_), .C(new_new_n495_), .D(i_5_), .Y(new_new_n657_));
  AO220      g635(.A0(new_new_n657_), .A1(i_0_), .B0(new_new_n655_), .B1(i_6_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n658_), .B(new_new_n654_), .Y(new_new_n659_));
  NA3        g637(.A(new_new_n659_), .B(new_new_n652_), .C(new_new_n649_), .Y(new_new_n660_));
  NA2        g638(.A(i_11_), .B(i_9_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n304_), .B(new_new_n151_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n662_), .B(new_new_n139_), .Y(new_new_n663_));
  NO2        g641(.A(new_new_n661_), .B(new_new_n70_), .Y(new_new_n664_));
  NO2        g642(.A(new_new_n149_), .B(i_0_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n354_), .B(new_new_n194_), .Y(new_new_n666_));
  OAI220     g644(.A0(i_12_), .A1(new_new_n640_), .B0(new_new_n666_), .B1(new_new_n149_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n667_), .B(new_new_n663_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n485_), .B(new_new_n106_), .Y(new_new_n669_));
  NO2        g647(.A(i_6_), .B(new_new_n669_), .Y(new_new_n670_));
  AOI210     g648(.A0(new_new_n339_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n146_), .B(new_new_n92_), .Y(new_new_n672_));
  NOi32      g650(.An(new_new_n671_), .Bn(new_new_n159_), .C(new_new_n672_), .Y(new_new_n673_));
  NO2        g651(.A(new_new_n37_), .B(new_new_n633_), .Y(new_new_n674_));
  NO3        g652(.A(new_new_n674_), .B(new_new_n673_), .C(new_new_n670_), .Y(new_new_n675_));
  NOi31      g653(.An(i_7_), .B(i_0_), .C(new_new_n534_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n675_), .B(new_new_n668_), .Y(new_new_n677_));
  INV        g655(.A(new_new_n626_), .Y(new_new_n678_));
  OA210      g656(.A0(new_new_n354_), .A1(new_new_n188_), .B0(new_new_n353_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n678_), .B(new_new_n664_), .Y(new_new_n680_));
  NA3        g658(.A(new_new_n353_), .B(i_2_), .C(new_new_n44_), .Y(new_new_n681_));
  INV        g659(.A(new_new_n681_), .Y(new_new_n682_));
  INV        g660(.A(new_new_n158_), .Y(new_new_n683_));
  AOI220     g661(.A0(new_new_n683_), .A1(new_new_n354_), .B0(new_new_n682_), .B1(new_new_n70_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n86_), .B(new_new_n43_), .Y(new_new_n685_));
  NO2        g663(.A(new_new_n72_), .B(new_new_n554_), .Y(new_new_n686_));
  NA2        g664(.A(new_new_n686_), .B(new_new_n685_), .Y(new_new_n687_));
  NO2        g665(.A(new_new_n687_), .B(new_new_n46_), .Y(new_new_n688_));
  NO3        g666(.A(i_5_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n689_));
  INV        g667(.A(new_new_n689_), .Y(new_new_n690_));
  NO2        g668(.A(new_new_n690_), .B(new_new_n147_), .Y(new_new_n691_));
  NO3        g669(.A(new_new_n691_), .B(new_new_n688_), .C(new_new_n383_), .Y(new_new_n692_));
  NA3        g670(.A(new_new_n692_), .B(new_new_n684_), .C(new_new_n680_), .Y(new_new_n693_));
  NO3        g671(.A(new_new_n693_), .B(new_new_n677_), .C(new_new_n660_), .Y(new_new_n694_));
  NO2        g672(.A(i_0_), .B(new_new_n534_), .Y(new_new_n695_));
  NO2        g673(.A(new_new_n596_), .B(new_new_n672_), .Y(new_new_n696_));
  INV        g674(.A(new_new_n696_), .Y(new_new_n697_));
  NA3        g675(.A(new_new_n128_), .B(new_new_n498_), .C(new_new_n70_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n627_), .B(i_9_), .Y(new_new_n699_));
  AOI210     g677(.A0(new_new_n775_), .A1(new_new_n365_), .B0(new_new_n699_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n203_), .B(i_10_), .Y(new_new_n701_));
  AOI210     g679(.A0(new_new_n701_), .A1(new_new_n650_), .B0(new_new_n134_), .Y(new_new_n702_));
  NO2        g680(.A(new_new_n702_), .B(new_new_n700_), .Y(new_new_n703_));
  NA3        g681(.A(new_new_n703_), .B(new_new_n698_), .C(new_new_n697_), .Y(new_new_n704_));
  NO2        g682(.A(new_new_n141_), .B(new_new_n768_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n705_), .Y(new_new_n706_));
  NA2        g684(.A(new_new_n418_), .B(new_new_n72_), .Y(new_new_n707_));
  NO3        g685(.A(new_new_n178_), .B(new_new_n297_), .C(i_0_), .Y(new_new_n708_));
  OAI210     g686(.A0(new_new_n708_), .A1(new_new_n73_), .B0(i_13_), .Y(new_new_n709_));
  NA3        g687(.A(new_new_n709_), .B(new_new_n707_), .C(new_new_n706_), .Y(new_new_n710_));
  AOI210     g688(.A0(i_6_), .A1(new_new_n695_), .B0(new_new_n94_), .Y(new_new_n711_));
  BUFFER     g689(.A(new_new_n711_), .Y(new_new_n712_));
  AOI210     g690(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n149_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n713_), .B(new_new_n679_), .Y(new_new_n714_));
  NOi31      g692(.An(new_new_n301_), .B(i_11_), .C(new_new_n200_), .Y(new_new_n715_));
  NO3        g693(.A(new_new_n661_), .B(new_new_n185_), .C(new_new_n161_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n716_), .B(new_new_n715_), .Y(new_new_n717_));
  NA3        g695(.A(new_new_n717_), .B(new_new_n714_), .C(new_new_n712_), .Y(new_new_n718_));
  NAi21      g696(.An(new_new_n201_), .B(new_new_n202_), .Y(new_new_n719_));
  NO4        g697(.A(new_new_n200_), .B(new_new_n178_), .C(i_0_), .D(i_12_), .Y(new_new_n720_));
  AOI220     g698(.A0(new_new_n720_), .A1(new_new_n719_), .B0(new_new_n590_), .B1(new_new_n150_), .Y(new_new_n721_));
  AN2        g699(.A(new_new_n656_), .B(new_new_n134_), .Y(new_new_n722_));
  NO4        g700(.A(new_new_n722_), .B(i_12_), .C(new_new_n478_), .D(new_new_n116_), .Y(new_new_n723_));
  INV        g701(.A(new_new_n723_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n421_), .B(i_11_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n725_), .B(new_new_n778_), .Y(new_new_n726_));
  NA2        g704(.A(i_7_), .B(new_new_n352_), .Y(new_new_n727_));
  OAI220     g705(.A0(i_6_), .A1(new_new_n776_), .B0(new_new_n727_), .B1(i_1_), .Y(new_new_n728_));
  AOI210     g706(.A0(new_new_n728_), .A1(new_new_n665_), .B0(new_new_n726_), .Y(new_new_n729_));
  NA3        g707(.A(new_new_n729_), .B(new_new_n724_), .C(new_new_n721_), .Y(new_new_n730_));
  NO4        g708(.A(new_new_n730_), .B(new_new_n718_), .C(new_new_n710_), .D(new_new_n704_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n770_), .B(new_new_n37_), .Y(new_new_n732_));
  NA2        g710(.A(new_new_n732_), .B(new_new_n764_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n733_), .B(new_new_n175_), .Y(new_new_n734_));
  OAI210     g712(.A0(new_new_n451_), .A1(new_new_n449_), .B0(new_new_n251_), .Y(new_new_n735_));
  INV        g713(.A(new_new_n735_), .Y(new_new_n736_));
  NO4        g714(.A(new_new_n196_), .B(new_new_n127_), .C(new_new_n499_), .D(new_new_n37_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n737_), .B(new_new_n651_), .Y(new_new_n738_));
  NA2        g716(.A(new_new_n725_), .B(new_new_n738_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n736_), .A1(new_new_n47_), .B0(new_new_n739_), .Y(new_new_n740_));
  AOI210     g718(.A0(new_new_n740_), .A1(new_new_n734_), .B0(new_new_n70_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n415_), .B(new_new_n294_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n742_), .B(new_new_n558_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n93_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n744_), .B(new_new_n73_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n713_), .A1(new_new_n777_), .B0(new_new_n676_), .Y(new_new_n746_));
  AOI210     g724(.A0(new_new_n746_), .A1(new_new_n745_), .B0(new_new_n499_), .Y(new_new_n747_));
  INV        g725(.A(new_new_n56_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n748_), .B(new_new_n73_), .Y(new_new_n749_));
  NO2        g727(.A(new_new_n749_), .B(new_new_n198_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n750_), .B(new_new_n747_), .Y(new_new_n751_));
  NO3        g729(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n752_));
  INV        g730(.A(new_new_n752_), .Y(new_new_n753_));
  NO2        g731(.A(new_new_n753_), .B(new_new_n534_), .Y(new_new_n754_));
  INV        g732(.A(new_new_n412_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n755_), .B(new_new_n40_), .Y(new_new_n756_));
  NO3        g734(.A(new_new_n756_), .B(new_new_n754_), .C(new_new_n215_), .Y(new_new_n757_));
  OAI210     g735(.A0(new_new_n751_), .A1(i_4_), .B0(new_new_n757_), .Y(new_new_n758_));
  NO3        g736(.A(new_new_n758_), .B(new_new_n743_), .C(new_new_n741_), .Y(new_new_n759_));
  NA4        g737(.A(new_new_n759_), .B(new_new_n731_), .C(new_new_n694_), .D(new_new_n644_), .Y(mai4));
  INV        g738(.A(i_2_), .Y(new_new_n763_));
  INV        g739(.A(new_new_n140_), .Y(new_new_n764_));
  INV        g740(.A(i_11_), .Y(new_new_n765_));
  INV        g741(.A(new_new_n116_), .Y(new_new_n766_));
  INV        g742(.A(i_9_), .Y(new_new_n767_));
  INV        g743(.A(new_new_n261_), .Y(new_new_n768_));
  INV        g744(.A(i_1_), .Y(new_new_n769_));
  INV        g745(.A(i_11_), .Y(new_new_n770_));
  INV        g746(.A(i_7_), .Y(new_new_n771_));
  INV        g747(.A(i_9_), .Y(new_new_n772_));
  INV        g748(.A(i_6_), .Y(new_new_n773_));
  INV        g749(.A(i_10_), .Y(new_new_n774_));
  INV        g750(.A(i_6_), .Y(new_new_n775_));
  INV        g751(.A(i_10_), .Y(new_new_n776_));
  INV        g752(.A(i_7_), .Y(new_new_n777_));
  INV        g753(.A(i_2_), .Y(new_new_n778_));
  INV        g754(.A(new_new_n637_), .Y(new_new_n779_));
  INV        g755(.A(i_0_), .Y(new_new_n780_));
endmodule


