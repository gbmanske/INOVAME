//Benchmark atmr_misex3_1774_0.0313

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1244_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1287_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1493_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1504_, men_men_n1505_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(g), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(g), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(g), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO4        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NA2        o0031(.A(g), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NAi21      o0032(.An(i), .B(h), .Y(ori_ori_n61_));
  NAi31      o0033(.An(i), .B(l), .C(j), .Y(ori_ori_n62_));
  OAI220     o0034(.A0(ori_ori_n62_), .A1(ori_ori_n49_), .B0(ori_ori_n61_), .B1(ori_ori_n44_), .Y(ori_ori_n63_));
  NAi31      o0035(.An(ori_ori_n60_), .B(ori_ori_n63_), .C(ori_ori_n58_), .Y(ori_ori_n64_));
  NAi41      o0036(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n65_));
  NA2        o0037(.A(g), .B(f), .Y(ori_ori_n66_));
  NO2        o0038(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NAi21      o0039(.An(i), .B(j), .Y(ori_ori_n68_));
  NAi32      o0040(.An(n), .Bn(k), .C(m), .Y(ori_ori_n69_));
  NAi31      o0041(.An(l), .B(m), .C(k), .Y(ori_ori_n70_));
  NAi21      o0042(.An(e), .B(h), .Y(ori_ori_n71_));
  NAi41      o0043(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n72_));
  INV        o0044(.A(m), .Y(ori_ori_n73_));
  NOi21      o0045(.An(k), .B(l), .Y(ori_ori_n74_));
  NA2        o0046(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  AN4        o0047(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n76_));
  NOi31      o0048(.An(h), .B(g), .C(f), .Y(ori_ori_n77_));
  NAi32      o0049(.An(m), .Bn(k), .C(j), .Y(ori_ori_n78_));
  NOi32      o0050(.An(h), .Bn(g), .C(f), .Y(ori_ori_n79_));
  INV        o0051(.A(ori_ori_n64_), .Y(ori_ori_n80_));
  INV        o0052(.A(n), .Y(ori_ori_n81_));
  NOi32      o0053(.An(e), .Bn(b), .C(d), .Y(ori_ori_n82_));
  NA2        o0054(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n83_));
  INV        o0055(.A(j), .Y(ori_ori_n84_));
  AN3        o0056(.A(m), .B(k), .C(i), .Y(ori_ori_n85_));
  NA3        o0057(.A(ori_ori_n85_), .B(ori_ori_n84_), .C(g), .Y(ori_ori_n86_));
  NO2        o0058(.A(ori_ori_n86_), .B(f), .Y(ori_ori_n87_));
  NAi32      o0059(.An(g), .Bn(f), .C(h), .Y(ori_ori_n88_));
  NAi31      o0060(.An(j), .B(m), .C(l), .Y(ori_ori_n89_));
  NO2        o0061(.A(ori_ori_n89_), .B(ori_ori_n88_), .Y(ori_ori_n90_));
  NA2        o0062(.A(m), .B(l), .Y(ori_ori_n91_));
  NAi31      o0063(.An(k), .B(j), .C(g), .Y(ori_ori_n92_));
  NO3        o0064(.A(ori_ori_n92_), .B(ori_ori_n91_), .C(f), .Y(ori_ori_n93_));
  AN2        o0065(.A(j), .B(g), .Y(ori_ori_n94_));
  NOi32      o0066(.An(m), .Bn(l), .C(i), .Y(ori_ori_n95_));
  NOi21      o0067(.An(g), .B(i), .Y(ori_ori_n96_));
  NOi32      o0068(.An(m), .Bn(j), .C(k), .Y(ori_ori_n97_));
  AOI220     o0069(.A0(ori_ori_n97_), .A1(ori_ori_n96_), .B0(ori_ori_n95_), .B1(ori_ori_n94_), .Y(ori_ori_n98_));
  NO2        o0070(.A(ori_ori_n98_), .B(f), .Y(ori_ori_n99_));
  NO3        o0071(.A(ori_ori_n99_), .B(ori_ori_n90_), .C(ori_ori_n87_), .Y(ori_ori_n100_));
  NAi41      o0072(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n101_));
  AN2        o0073(.A(e), .B(b), .Y(ori_ori_n102_));
  NOi31      o0074(.An(c), .B(h), .C(f), .Y(ori_ori_n103_));
  NA2        o0075(.A(ori_ori_n103_), .B(ori_ori_n102_), .Y(ori_ori_n104_));
  NO2        o0076(.A(ori_ori_n104_), .B(ori_ori_n101_), .Y(ori_ori_n105_));
  NOi21      o0077(.An(g), .B(f), .Y(ori_ori_n106_));
  NOi21      o0078(.An(i), .B(h), .Y(ori_ori_n107_));
  NA3        o0079(.A(ori_ori_n107_), .B(ori_ori_n106_), .C(ori_ori_n36_), .Y(ori_ori_n108_));
  INV        o0080(.A(a), .Y(ori_ori_n109_));
  NA2        o0081(.A(ori_ori_n102_), .B(ori_ori_n109_), .Y(ori_ori_n110_));
  INV        o0082(.A(l), .Y(ori_ori_n111_));
  NOi21      o0083(.An(m), .B(n), .Y(ori_ori_n112_));
  AN2        o0084(.A(k), .B(h), .Y(ori_ori_n113_));
  NO2        o0085(.A(ori_ori_n108_), .B(ori_ori_n83_), .Y(ori_ori_n114_));
  INV        o0086(.A(b), .Y(ori_ori_n115_));
  NA2        o0087(.A(l), .B(j), .Y(ori_ori_n116_));
  AN2        o0088(.A(k), .B(i), .Y(ori_ori_n117_));
  NA2        o0089(.A(g), .B(e), .Y(ori_ori_n118_));
  NOi32      o0090(.An(c), .Bn(a), .C(d), .Y(ori_ori_n119_));
  NA2        o0091(.A(ori_ori_n119_), .B(ori_ori_n112_), .Y(ori_ori_n120_));
  NO2        o0092(.A(ori_ori_n114_), .B(ori_ori_n105_), .Y(ori_ori_n121_));
  OAI210     o0093(.A0(ori_ori_n100_), .A1(ori_ori_n83_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  NOi31      o0094(.An(k), .B(m), .C(j), .Y(ori_ori_n123_));
  NA3        o0095(.A(ori_ori_n123_), .B(ori_ori_n77_), .C(ori_ori_n76_), .Y(ori_ori_n124_));
  NOi31      o0096(.An(k), .B(m), .C(i), .Y(ori_ori_n125_));
  NA3        o0097(.A(ori_ori_n125_), .B(ori_ori_n79_), .C(ori_ori_n76_), .Y(ori_ori_n126_));
  NA2        o0098(.A(ori_ori_n126_), .B(ori_ori_n124_), .Y(ori_ori_n127_));
  NOi32      o0099(.An(f), .Bn(b), .C(e), .Y(ori_ori_n128_));
  NAi21      o0100(.An(g), .B(h), .Y(ori_ori_n129_));
  NAi21      o0101(.An(m), .B(n), .Y(ori_ori_n130_));
  NAi21      o0102(.An(j), .B(k), .Y(ori_ori_n131_));
  NO3        o0103(.A(ori_ori_n131_), .B(ori_ori_n130_), .C(ori_ori_n129_), .Y(ori_ori_n132_));
  NAi41      o0104(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n133_));
  NAi31      o0105(.An(j), .B(k), .C(h), .Y(ori_ori_n134_));
  NO3        o0106(.A(ori_ori_n134_), .B(ori_ori_n133_), .C(ori_ori_n130_), .Y(ori_ori_n135_));
  AOI210     o0107(.A0(ori_ori_n132_), .A1(ori_ori_n128_), .B0(ori_ori_n135_), .Y(ori_ori_n136_));
  NO2        o0108(.A(k), .B(j), .Y(ori_ori_n137_));
  NO2        o0109(.A(ori_ori_n137_), .B(ori_ori_n130_), .Y(ori_ori_n138_));
  AN2        o0110(.A(k), .B(j), .Y(ori_ori_n139_));
  NAi21      o0111(.An(c), .B(b), .Y(ori_ori_n140_));
  NA2        o0112(.A(f), .B(d), .Y(ori_ori_n141_));
  NO4        o0113(.A(ori_ori_n141_), .B(ori_ori_n140_), .C(ori_ori_n139_), .D(ori_ori_n129_), .Y(ori_ori_n142_));
  NA2        o0114(.A(h), .B(c), .Y(ori_ori_n143_));
  NAi31      o0115(.An(f), .B(e), .C(b), .Y(ori_ori_n144_));
  NA2        o0116(.A(ori_ori_n142_), .B(ori_ori_n138_), .Y(ori_ori_n145_));
  NA2        o0117(.A(d), .B(b), .Y(ori_ori_n146_));
  NAi21      o0118(.An(e), .B(f), .Y(ori_ori_n147_));
  NO2        o0119(.A(ori_ori_n147_), .B(ori_ori_n146_), .Y(ori_ori_n148_));
  NA2        o0120(.A(b), .B(a), .Y(ori_ori_n149_));
  NAi21      o0121(.An(e), .B(g), .Y(ori_ori_n150_));
  NAi21      o0122(.An(c), .B(d), .Y(ori_ori_n151_));
  NAi31      o0123(.An(l), .B(k), .C(h), .Y(ori_ori_n152_));
  NO2        o0124(.A(ori_ori_n130_), .B(ori_ori_n152_), .Y(ori_ori_n153_));
  NA2        o0125(.A(ori_ori_n153_), .B(ori_ori_n148_), .Y(ori_ori_n154_));
  NAi41      o0126(.An(ori_ori_n127_), .B(ori_ori_n154_), .C(ori_ori_n145_), .D(ori_ori_n136_), .Y(ori_ori_n155_));
  NAi31      o0127(.An(e), .B(f), .C(b), .Y(ori_ori_n156_));
  NOi21      o0128(.An(g), .B(d), .Y(ori_ori_n157_));
  NO2        o0129(.A(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  NOi21      o0130(.An(h), .B(i), .Y(ori_ori_n159_));
  NOi21      o0131(.An(k), .B(m), .Y(ori_ori_n160_));
  NA3        o0132(.A(ori_ori_n160_), .B(ori_ori_n159_), .C(n), .Y(ori_ori_n161_));
  NOi21      o0133(.An(ori_ori_n158_), .B(ori_ori_n161_), .Y(ori_ori_n162_));
  NOi21      o0134(.An(h), .B(g), .Y(ori_ori_n163_));
  NO2        o0135(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n164_));
  NAi31      o0136(.An(l), .B(j), .C(h), .Y(ori_ori_n165_));
  NO2        o0137(.A(ori_ori_n165_), .B(ori_ori_n49_), .Y(ori_ori_n166_));
  NA2        o0138(.A(ori_ori_n166_), .B(ori_ori_n67_), .Y(ori_ori_n167_));
  NOi32      o0139(.An(n), .Bn(k), .C(m), .Y(ori_ori_n168_));
  INV        o0140(.A(ori_ori_n167_), .Y(ori_ori_n169_));
  NAi31      o0141(.An(d), .B(f), .C(c), .Y(ori_ori_n170_));
  NAi31      o0142(.An(e), .B(f), .C(c), .Y(ori_ori_n171_));
  NA2        o0143(.A(ori_ori_n171_), .B(ori_ori_n170_), .Y(ori_ori_n172_));
  NA2        o0144(.A(j), .B(h), .Y(ori_ori_n173_));
  OR3        o0145(.A(n), .B(m), .C(k), .Y(ori_ori_n174_));
  NO2        o0146(.A(ori_ori_n174_), .B(ori_ori_n173_), .Y(ori_ori_n175_));
  NAi32      o0147(.An(m), .Bn(k), .C(n), .Y(ori_ori_n176_));
  NO2        o0148(.A(ori_ori_n176_), .B(ori_ori_n173_), .Y(ori_ori_n177_));
  AOI220     o0149(.A0(ori_ori_n177_), .A1(ori_ori_n158_), .B0(ori_ori_n175_), .B1(ori_ori_n172_), .Y(ori_ori_n178_));
  NO2        o0150(.A(n), .B(m), .Y(ori_ori_n179_));
  NA2        o0151(.A(ori_ori_n179_), .B(ori_ori_n50_), .Y(ori_ori_n180_));
  NAi21      o0152(.An(f), .B(e), .Y(ori_ori_n181_));
  NA2        o0153(.A(d), .B(c), .Y(ori_ori_n182_));
  NO2        o0154(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n183_));
  NOi21      o0155(.An(ori_ori_n183_), .B(ori_ori_n180_), .Y(ori_ori_n184_));
  NAi21      o0156(.An(d), .B(c), .Y(ori_ori_n185_));
  NAi31      o0157(.An(m), .B(n), .C(b), .Y(ori_ori_n186_));
  NA2        o0158(.A(k), .B(i), .Y(ori_ori_n187_));
  NAi21      o0159(.An(h), .B(f), .Y(ori_ori_n188_));
  NO2        o0160(.A(ori_ori_n188_), .B(ori_ori_n187_), .Y(ori_ori_n189_));
  NO2        o0161(.A(ori_ori_n186_), .B(ori_ori_n151_), .Y(ori_ori_n190_));
  NA2        o0162(.A(ori_ori_n190_), .B(ori_ori_n189_), .Y(ori_ori_n191_));
  NOi32      o0163(.An(f), .Bn(c), .C(d), .Y(ori_ori_n192_));
  NOi32      o0164(.An(f), .Bn(c), .C(e), .Y(ori_ori_n193_));
  NO2        o0165(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NO3        o0166(.A(n), .B(m), .C(j), .Y(ori_ori_n195_));
  NA2        o0167(.A(ori_ori_n195_), .B(ori_ori_n113_), .Y(ori_ori_n196_));
  AO210      o0168(.A0(ori_ori_n196_), .A1(ori_ori_n180_), .B0(ori_ori_n194_), .Y(ori_ori_n197_));
  NAi41      o0169(.An(ori_ori_n184_), .B(ori_ori_n197_), .C(ori_ori_n191_), .D(ori_ori_n178_), .Y(ori_ori_n198_));
  OR4        o0170(.A(ori_ori_n198_), .B(ori_ori_n169_), .C(ori_ori_n162_), .D(ori_ori_n155_), .Y(ori_ori_n199_));
  NO4        o0171(.A(ori_ori_n199_), .B(ori_ori_n122_), .C(ori_ori_n80_), .D(ori_ori_n55_), .Y(ori_ori_n200_));
  NA3        o0172(.A(m), .B(ori_ori_n111_), .C(j), .Y(ori_ori_n201_));
  NAi31      o0173(.An(n), .B(h), .C(g), .Y(ori_ori_n202_));
  NO2        o0174(.A(ori_ori_n202_), .B(ori_ori_n201_), .Y(ori_ori_n203_));
  NOi32      o0175(.An(m), .Bn(k), .C(l), .Y(ori_ori_n204_));
  NA3        o0176(.A(ori_ori_n204_), .B(ori_ori_n84_), .C(g), .Y(ori_ori_n205_));
  NO2        o0177(.A(ori_ori_n205_), .B(n), .Y(ori_ori_n206_));
  NOi21      o0178(.An(k), .B(j), .Y(ori_ori_n207_));
  NA4        o0179(.A(ori_ori_n207_), .B(ori_ori_n112_), .C(i), .D(g), .Y(ori_ori_n208_));
  AN2        o0180(.A(i), .B(g), .Y(ori_ori_n209_));
  NA3        o0181(.A(ori_ori_n74_), .B(ori_ori_n209_), .C(ori_ori_n112_), .Y(ori_ori_n210_));
  NA2        o0182(.A(ori_ori_n210_), .B(ori_ori_n208_), .Y(ori_ori_n211_));
  NO2        o0183(.A(ori_ori_n211_), .B(ori_ori_n203_), .Y(ori_ori_n212_));
  NAi41      o0184(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n213_));
  INV        o0185(.A(ori_ori_n213_), .Y(ori_ori_n214_));
  INV        o0186(.A(f), .Y(ori_ori_n215_));
  INV        o0187(.A(g), .Y(ori_ori_n216_));
  NOi31      o0188(.An(i), .B(j), .C(h), .Y(ori_ori_n217_));
  NOi21      o0189(.An(l), .B(m), .Y(ori_ori_n218_));
  NA2        o0190(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  NO3        o0191(.A(ori_ori_n219_), .B(ori_ori_n216_), .C(ori_ori_n215_), .Y(ori_ori_n220_));
  NA2        o0192(.A(ori_ori_n220_), .B(ori_ori_n214_), .Y(ori_ori_n221_));
  OAI210     o0193(.A0(ori_ori_n212_), .A1(ori_ori_n32_), .B0(ori_ori_n221_), .Y(ori_ori_n222_));
  NOi21      o0194(.An(n), .B(m), .Y(ori_ori_n223_));
  NOi32      o0195(.An(l), .Bn(i), .C(j), .Y(ori_ori_n224_));
  NA2        o0196(.A(ori_ori_n224_), .B(ori_ori_n223_), .Y(ori_ori_n225_));
  NAi21      o0197(.An(j), .B(h), .Y(ori_ori_n226_));
  XN2        o0198(.A(i), .B(h), .Y(ori_ori_n227_));
  NA2        o0199(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  NOi31      o0200(.An(k), .B(n), .C(m), .Y(ori_ori_n229_));
  NOi31      o0201(.An(ori_ori_n229_), .B(ori_ori_n182_), .C(ori_ori_n181_), .Y(ori_ori_n230_));
  NA2        o0202(.A(ori_ori_n230_), .B(ori_ori_n228_), .Y(ori_ori_n231_));
  NAi31      o0203(.An(f), .B(e), .C(c), .Y(ori_ori_n232_));
  NO4        o0204(.A(ori_ori_n232_), .B(ori_ori_n174_), .C(ori_ori_n173_), .D(ori_ori_n59_), .Y(ori_ori_n233_));
  NA4        o0205(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n234_));
  NAi32      o0206(.An(m), .Bn(i), .C(k), .Y(ori_ori_n235_));
  NO3        o0207(.A(ori_ori_n235_), .B(ori_ori_n88_), .C(ori_ori_n234_), .Y(ori_ori_n236_));
  INV        o0208(.A(k), .Y(ori_ori_n237_));
  NO2        o0209(.A(ori_ori_n236_), .B(ori_ori_n233_), .Y(ori_ori_n238_));
  NAi21      o0210(.An(n), .B(a), .Y(ori_ori_n239_));
  NO2        o0211(.A(ori_ori_n239_), .B(ori_ori_n146_), .Y(ori_ori_n240_));
  NAi41      o0212(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n241_), .B(e), .Y(ori_ori_n242_));
  NA2        o0214(.A(ori_ori_n242_), .B(ori_ori_n240_), .Y(ori_ori_n243_));
  AN3        o0215(.A(ori_ori_n243_), .B(ori_ori_n238_), .C(ori_ori_n231_), .Y(ori_ori_n244_));
  OR2        o0216(.A(h), .B(g), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(ori_ori_n101_), .Y(ori_ori_n246_));
  NA2        o0218(.A(ori_ori_n246_), .B(ori_ori_n128_), .Y(ori_ori_n247_));
  NAi41      o0219(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n248_));
  NO2        o0220(.A(ori_ori_n248_), .B(ori_ori_n215_), .Y(ori_ori_n249_));
  NA2        o0221(.A(ori_ori_n160_), .B(ori_ori_n107_), .Y(ori_ori_n250_));
  NAi21      o0222(.An(ori_ori_n250_), .B(ori_ori_n249_), .Y(ori_ori_n251_));
  NO2        o0223(.A(n), .B(a), .Y(ori_ori_n252_));
  NAi31      o0224(.An(ori_ori_n241_), .B(ori_ori_n252_), .C(ori_ori_n102_), .Y(ori_ori_n253_));
  AN2        o0225(.A(ori_ori_n253_), .B(ori_ori_n251_), .Y(ori_ori_n254_));
  NAi21      o0226(.An(h), .B(i), .Y(ori_ori_n255_));
  NA2        o0227(.A(ori_ori_n179_), .B(k), .Y(ori_ori_n256_));
  NO2        o0228(.A(ori_ori_n256_), .B(ori_ori_n255_), .Y(ori_ori_n257_));
  NA2        o0229(.A(ori_ori_n257_), .B(ori_ori_n192_), .Y(ori_ori_n258_));
  NA3        o0230(.A(ori_ori_n258_), .B(ori_ori_n254_), .C(ori_ori_n247_), .Y(ori_ori_n259_));
  NOi21      o0231(.An(g), .B(e), .Y(ori_ori_n260_));
  NO2        o0232(.A(ori_ori_n72_), .B(ori_ori_n73_), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n261_), .B(ori_ori_n260_), .Y(ori_ori_n262_));
  NOi32      o0234(.An(l), .Bn(j), .C(i), .Y(ori_ori_n263_));
  AOI210     o0235(.A0(ori_ori_n74_), .A1(ori_ori_n84_), .B0(ori_ori_n263_), .Y(ori_ori_n264_));
  NO2        o0236(.A(ori_ori_n255_), .B(ori_ori_n44_), .Y(ori_ori_n265_));
  NAi21      o0237(.An(f), .B(g), .Y(ori_ori_n266_));
  NO2        o0238(.A(ori_ori_n266_), .B(ori_ori_n65_), .Y(ori_ori_n267_));
  NA2        o0239(.A(ori_ori_n265_), .B(ori_ori_n67_), .Y(ori_ori_n268_));
  OAI210     o0240(.A0(ori_ori_n264_), .A1(ori_ori_n262_), .B0(ori_ori_n268_), .Y(ori_ori_n269_));
  NO2        o0241(.A(ori_ori_n131_), .B(ori_ori_n49_), .Y(ori_ori_n270_));
  NOi41      o0242(.An(ori_ori_n244_), .B(ori_ori_n269_), .C(ori_ori_n259_), .D(ori_ori_n222_), .Y(ori_ori_n271_));
  NO4        o0243(.A(ori_ori_n203_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n272_));
  NO2        o0244(.A(ori_ori_n272_), .B(ori_ori_n110_), .Y(ori_ori_n273_));
  NA3        o0245(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n274_));
  NAi21      o0246(.An(h), .B(g), .Y(ori_ori_n275_));
  OR4        o0247(.A(ori_ori_n275_), .B(ori_ori_n274_), .C(ori_ori_n225_), .D(e), .Y(ori_ori_n276_));
  NAi31      o0248(.An(g), .B(k), .C(h), .Y(ori_ori_n277_));
  NAi31      o0249(.An(e), .B(d), .C(a), .Y(ori_ori_n278_));
  INV        o0250(.A(ori_ori_n276_), .Y(ori_ori_n279_));
  NA3        o0251(.A(ori_ori_n160_), .B(ori_ori_n159_), .C(ori_ori_n81_), .Y(ori_ori_n280_));
  NO2        o0252(.A(ori_ori_n280_), .B(ori_ori_n194_), .Y(ori_ori_n281_));
  INV        o0253(.A(ori_ori_n281_), .Y(ori_ori_n282_));
  NA3        o0254(.A(e), .B(c), .C(b), .Y(ori_ori_n283_));
  NO2        o0255(.A(ori_ori_n60_), .B(ori_ori_n283_), .Y(ori_ori_n284_));
  NAi32      o0256(.An(k), .Bn(i), .C(j), .Y(ori_ori_n285_));
  NAi31      o0257(.An(h), .B(l), .C(i), .Y(ori_ori_n286_));
  NA3        o0258(.A(ori_ori_n286_), .B(ori_ori_n285_), .C(ori_ori_n165_), .Y(ori_ori_n287_));
  NOi21      o0259(.An(ori_ori_n287_), .B(ori_ori_n49_), .Y(ori_ori_n288_));
  OAI210     o0260(.A0(ori_ori_n267_), .A1(ori_ori_n284_), .B0(ori_ori_n288_), .Y(ori_ori_n289_));
  NAi21      o0261(.An(l), .B(k), .Y(ori_ori_n290_));
  NO2        o0262(.A(ori_ori_n290_), .B(ori_ori_n49_), .Y(ori_ori_n291_));
  NOi21      o0263(.An(l), .B(j), .Y(ori_ori_n292_));
  NA2        o0264(.A(ori_ori_n163_), .B(ori_ori_n292_), .Y(ori_ori_n293_));
  NAi32      o0265(.An(j), .Bn(h), .C(i), .Y(ori_ori_n294_));
  NAi21      o0266(.An(m), .B(l), .Y(ori_ori_n295_));
  NO3        o0267(.A(ori_ori_n295_), .B(ori_ori_n294_), .C(ori_ori_n81_), .Y(ori_ori_n296_));
  NA2        o0268(.A(h), .B(g), .Y(ori_ori_n297_));
  NA2        o0269(.A(ori_ori_n168_), .B(ori_ori_n45_), .Y(ori_ori_n298_));
  NO2        o0270(.A(ori_ori_n298_), .B(ori_ori_n297_), .Y(ori_ori_n299_));
  NA2        o0271(.A(ori_ori_n299_), .B(ori_ori_n164_), .Y(ori_ori_n300_));
  NA3        o0272(.A(ori_ori_n300_), .B(ori_ori_n289_), .C(ori_ori_n282_), .Y(ori_ori_n301_));
  NO2        o0273(.A(ori_ori_n144_), .B(d), .Y(ori_ori_n302_));
  NA2        o0274(.A(ori_ori_n302_), .B(ori_ori_n53_), .Y(ori_ori_n303_));
  NO2        o0275(.A(ori_ori_n104_), .B(ori_ori_n101_), .Y(ori_ori_n304_));
  NAi32      o0276(.An(n), .Bn(m), .C(l), .Y(ori_ori_n305_));
  NO2        o0277(.A(ori_ori_n305_), .B(ori_ori_n294_), .Y(ori_ori_n306_));
  NA2        o0278(.A(ori_ori_n306_), .B(ori_ori_n183_), .Y(ori_ori_n307_));
  NO2        o0279(.A(ori_ori_n120_), .B(ori_ori_n115_), .Y(ori_ori_n308_));
  NAi31      o0280(.An(k), .B(l), .C(j), .Y(ori_ori_n309_));
  OAI210     o0281(.A0(ori_ori_n290_), .A1(j), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  NOi21      o0282(.An(ori_ori_n310_), .B(ori_ori_n118_), .Y(ori_ori_n311_));
  NA2        o0283(.A(ori_ori_n311_), .B(ori_ori_n308_), .Y(ori_ori_n312_));
  NA3        o0284(.A(ori_ori_n312_), .B(ori_ori_n307_), .C(ori_ori_n303_), .Y(ori_ori_n313_));
  NO4        o0285(.A(ori_ori_n313_), .B(ori_ori_n301_), .C(ori_ori_n279_), .D(ori_ori_n273_), .Y(ori_ori_n314_));
  NA2        o0286(.A(ori_ori_n257_), .B(ori_ori_n193_), .Y(ori_ori_n315_));
  NAi21      o0287(.An(m), .B(k), .Y(ori_ori_n316_));
  NO2        o0288(.A(ori_ori_n227_), .B(ori_ori_n316_), .Y(ori_ori_n317_));
  NAi41      o0289(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n318_));
  NO2        o0290(.A(ori_ori_n318_), .B(ori_ori_n150_), .Y(ori_ori_n319_));
  NA2        o0291(.A(ori_ori_n319_), .B(ori_ori_n317_), .Y(ori_ori_n320_));
  NAi31      o0292(.An(i), .B(l), .C(h), .Y(ori_ori_n321_));
  NO4        o0293(.A(ori_ori_n321_), .B(ori_ori_n150_), .C(ori_ori_n72_), .D(ori_ori_n73_), .Y(ori_ori_n322_));
  NA2        o0294(.A(e), .B(c), .Y(ori_ori_n323_));
  NO3        o0295(.A(ori_ori_n323_), .B(n), .C(d), .Y(ori_ori_n324_));
  NOi21      o0296(.An(f), .B(h), .Y(ori_ori_n325_));
  NAi31      o0297(.An(d), .B(e), .C(b), .Y(ori_ori_n326_));
  NAi31      o0298(.An(ori_ori_n322_), .B(ori_ori_n320_), .C(ori_ori_n315_), .Y(ori_ori_n327_));
  NO4        o0299(.A(ori_ori_n318_), .B(ori_ori_n78_), .C(ori_ori_n71_), .D(ori_ori_n216_), .Y(ori_ori_n328_));
  NA2        o0300(.A(ori_ori_n252_), .B(ori_ori_n102_), .Y(ori_ori_n329_));
  OR2        o0301(.A(ori_ori_n329_), .B(ori_ori_n205_), .Y(ori_ori_n330_));
  NOi31      o0302(.An(l), .B(n), .C(m), .Y(ori_ori_n331_));
  NA2        o0303(.A(ori_ori_n331_), .B(ori_ori_n217_), .Y(ori_ori_n332_));
  NO2        o0304(.A(ori_ori_n332_), .B(ori_ori_n194_), .Y(ori_ori_n333_));
  NAi32      o0305(.An(ori_ori_n333_), .Bn(ori_ori_n328_), .C(ori_ori_n330_), .Y(ori_ori_n334_));
  NAi32      o0306(.An(m), .Bn(j), .C(k), .Y(ori_ori_n335_));
  NAi41      o0307(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n336_));
  NOi31      o0308(.An(j), .B(m), .C(k), .Y(ori_ori_n337_));
  NO2        o0309(.A(ori_ori_n123_), .B(ori_ori_n337_), .Y(ori_ori_n338_));
  AN3        o0310(.A(h), .B(g), .C(f), .Y(ori_ori_n339_));
  NOi32      o0311(.An(m), .Bn(j), .C(l), .Y(ori_ori_n340_));
  NO2        o0312(.A(ori_ori_n340_), .B(ori_ori_n95_), .Y(ori_ori_n341_));
  NO2        o0313(.A(ori_ori_n295_), .B(ori_ori_n294_), .Y(ori_ori_n342_));
  NA2        o0314(.A(ori_ori_n249_), .B(ori_ori_n342_), .Y(ori_ori_n343_));
  NA2        o0315(.A(ori_ori_n235_), .B(ori_ori_n78_), .Y(ori_ori_n344_));
  NA3        o0316(.A(ori_ori_n344_), .B(ori_ori_n339_), .C(ori_ori_n214_), .Y(ori_ori_n345_));
  NA2        o0317(.A(ori_ori_n345_), .B(ori_ori_n343_), .Y(ori_ori_n346_));
  NA3        o0318(.A(h), .B(g), .C(f), .Y(ori_ori_n347_));
  NO2        o0319(.A(ori_ori_n347_), .B(ori_ori_n75_), .Y(ori_ori_n348_));
  NA2        o0320(.A(ori_ori_n163_), .B(e), .Y(ori_ori_n349_));
  NO2        o0321(.A(ori_ori_n349_), .B(ori_ori_n41_), .Y(ori_ori_n350_));
  NOi32      o0322(.An(j), .Bn(g), .C(i), .Y(ori_ori_n351_));
  NA3        o0323(.A(ori_ori_n351_), .B(ori_ori_n290_), .C(ori_ori_n112_), .Y(ori_ori_n352_));
  AO210      o0324(.A0(ori_ori_n110_), .A1(ori_ori_n32_), .B0(ori_ori_n352_), .Y(ori_ori_n353_));
  NOi32      o0325(.An(e), .Bn(b), .C(a), .Y(ori_ori_n354_));
  AN2        o0326(.A(l), .B(j), .Y(ori_ori_n355_));
  NO2        o0327(.A(ori_ori_n316_), .B(ori_ori_n355_), .Y(ori_ori_n356_));
  NO3        o0328(.A(ori_ori_n318_), .B(ori_ori_n71_), .C(ori_ori_n216_), .Y(ori_ori_n357_));
  NA3        o0329(.A(ori_ori_n210_), .B(ori_ori_n208_), .C(ori_ori_n35_), .Y(ori_ori_n358_));
  AOI220     o0330(.A0(ori_ori_n358_), .A1(ori_ori_n354_), .B0(ori_ori_n357_), .B1(ori_ori_n356_), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n326_), .B(n), .Y(ori_ori_n360_));
  NA2        o0332(.A(ori_ori_n209_), .B(k), .Y(ori_ori_n361_));
  NA3        o0333(.A(m), .B(ori_ori_n111_), .C(ori_ori_n215_), .Y(ori_ori_n362_));
  NA4        o0334(.A(ori_ori_n204_), .B(ori_ori_n84_), .C(g), .D(ori_ori_n215_), .Y(ori_ori_n363_));
  OAI210     o0335(.A0(ori_ori_n362_), .A1(ori_ori_n361_), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  NAi41      o0336(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n365_));
  NA2        o0337(.A(ori_ori_n51_), .B(ori_ori_n112_), .Y(ori_ori_n366_));
  NO2        o0338(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n367_));
  AOI220     o0339(.A0(ori_ori_n367_), .A1(b), .B0(ori_ori_n364_), .B1(ori_ori_n360_), .Y(ori_ori_n368_));
  NA3        o0340(.A(ori_ori_n368_), .B(ori_ori_n359_), .C(ori_ori_n353_), .Y(ori_ori_n369_));
  NO4        o0341(.A(ori_ori_n369_), .B(ori_ori_n346_), .C(ori_ori_n334_), .D(ori_ori_n327_), .Y(ori_ori_n370_));
  NA4        o0342(.A(ori_ori_n370_), .B(ori_ori_n314_), .C(ori_ori_n271_), .D(ori_ori_n200_), .Y(ori10));
  NA3        o0343(.A(m), .B(k), .C(i), .Y(ori_ori_n372_));
  NO3        o0344(.A(ori_ori_n372_), .B(j), .C(ori_ori_n216_), .Y(ori_ori_n373_));
  NOi21      o0345(.An(e), .B(f), .Y(ori_ori_n374_));
  NAi31      o0346(.An(b), .B(f), .C(c), .Y(ori_ori_n375_));
  INV        o0347(.A(ori_ori_n375_), .Y(ori_ori_n376_));
  NOi32      o0348(.An(k), .Bn(h), .C(j), .Y(ori_ori_n377_));
  NA2        o0349(.A(ori_ori_n377_), .B(ori_ori_n223_), .Y(ori_ori_n378_));
  NA2        o0350(.A(ori_ori_n161_), .B(ori_ori_n378_), .Y(ori_ori_n379_));
  NA2        o0351(.A(ori_ori_n379_), .B(ori_ori_n376_), .Y(ori_ori_n380_));
  AN2        o0352(.A(j), .B(h), .Y(ori_ori_n381_));
  NO3        o0353(.A(n), .B(m), .C(k), .Y(ori_ori_n382_));
  NA2        o0354(.A(ori_ori_n382_), .B(ori_ori_n381_), .Y(ori_ori_n383_));
  NO3        o0355(.A(ori_ori_n383_), .B(ori_ori_n151_), .C(ori_ori_n215_), .Y(ori_ori_n384_));
  OR2        o0356(.A(m), .B(k), .Y(ori_ori_n385_));
  NO2        o0357(.A(ori_ori_n173_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  NA4        o0358(.A(n), .B(f), .C(c), .D(ori_ori_n115_), .Y(ori_ori_n387_));
  NOi21      o0359(.An(ori_ori_n386_), .B(ori_ori_n387_), .Y(ori_ori_n388_));
  NOi32      o0360(.An(d), .Bn(a), .C(c), .Y(ori_ori_n389_));
  NA2        o0361(.A(ori_ori_n389_), .B(ori_ori_n181_), .Y(ori_ori_n390_));
  NAi21      o0362(.An(i), .B(g), .Y(ori_ori_n391_));
  NAi31      o0363(.An(k), .B(m), .C(j), .Y(ori_ori_n392_));
  NO3        o0364(.A(ori_ori_n392_), .B(ori_ori_n391_), .C(n), .Y(ori_ori_n393_));
  NOi21      o0365(.An(ori_ori_n393_), .B(ori_ori_n390_), .Y(ori_ori_n394_));
  NO3        o0366(.A(ori_ori_n394_), .B(ori_ori_n388_), .C(ori_ori_n384_), .Y(ori_ori_n395_));
  NO2        o0367(.A(ori_ori_n387_), .B(ori_ori_n295_), .Y(ori_ori_n396_));
  NOi32      o0368(.An(f), .Bn(d), .C(c), .Y(ori_ori_n397_));
  AOI220     o0369(.A0(ori_ori_n397_), .A1(ori_ori_n306_), .B0(ori_ori_n396_), .B1(ori_ori_n217_), .Y(ori_ori_n398_));
  NA3        o0370(.A(ori_ori_n398_), .B(ori_ori_n395_), .C(ori_ori_n380_), .Y(ori_ori_n399_));
  NO2        o0371(.A(ori_ori_n59_), .B(ori_ori_n115_), .Y(ori_ori_n400_));
  NA2        o0372(.A(ori_ori_n252_), .B(ori_ori_n400_), .Y(ori_ori_n401_));
  INV        o0373(.A(e), .Y(ori_ori_n402_));
  NA2        o0374(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n403_));
  OAI220     o0375(.A0(ori_ori_n403_), .A1(ori_ori_n201_), .B0(ori_ori_n205_), .B1(ori_ori_n402_), .Y(ori_ori_n404_));
  AN2        o0376(.A(g), .B(e), .Y(ori_ori_n405_));
  NA3        o0377(.A(ori_ori_n405_), .B(ori_ori_n204_), .C(i), .Y(ori_ori_n406_));
  OAI210     o0378(.A0(ori_ori_n86_), .A1(ori_ori_n402_), .B0(ori_ori_n406_), .Y(ori_ori_n407_));
  NO2        o0379(.A(ori_ori_n98_), .B(ori_ori_n402_), .Y(ori_ori_n408_));
  NO3        o0380(.A(ori_ori_n408_), .B(ori_ori_n407_), .C(ori_ori_n404_), .Y(ori_ori_n409_));
  NOi32      o0381(.An(h), .Bn(e), .C(g), .Y(ori_ori_n410_));
  NA3        o0382(.A(ori_ori_n410_), .B(ori_ori_n292_), .C(m), .Y(ori_ori_n411_));
  NOi21      o0383(.An(g), .B(h), .Y(ori_ori_n412_));
  AN3        o0384(.A(m), .B(l), .C(i), .Y(ori_ori_n413_));
  NA3        o0385(.A(ori_ori_n413_), .B(ori_ori_n412_), .C(e), .Y(ori_ori_n414_));
  AN3        o0386(.A(h), .B(g), .C(e), .Y(ori_ori_n415_));
  NA2        o0387(.A(ori_ori_n415_), .B(ori_ori_n95_), .Y(ori_ori_n416_));
  AN3        o0388(.A(ori_ori_n416_), .B(ori_ori_n414_), .C(ori_ori_n411_), .Y(ori_ori_n417_));
  AOI210     o0389(.A0(ori_ori_n417_), .A1(ori_ori_n409_), .B0(ori_ori_n401_), .Y(ori_ori_n418_));
  NA3        o0390(.A(ori_ori_n389_), .B(ori_ori_n181_), .C(ori_ori_n81_), .Y(ori_ori_n419_));
  NAi31      o0391(.An(b), .B(c), .C(a), .Y(ori_ori_n420_));
  NO2        o0392(.A(ori_ori_n420_), .B(n), .Y(ori_ori_n421_));
  NA2        o0393(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n422_));
  NO2        o0394(.A(ori_ori_n422_), .B(ori_ori_n147_), .Y(ori_ori_n423_));
  NA2        o0395(.A(ori_ori_n423_), .B(ori_ori_n421_), .Y(ori_ori_n424_));
  INV        o0396(.A(ori_ori_n424_), .Y(ori_ori_n425_));
  NO3        o0397(.A(ori_ori_n425_), .B(ori_ori_n418_), .C(ori_ori_n399_), .Y(ori_ori_n426_));
  NA2        o0398(.A(i), .B(g), .Y(ori_ori_n427_));
  NOi21      o0399(.An(d), .B(c), .Y(ori_ori_n428_));
  NA3        o0400(.A(i), .B(g), .C(f), .Y(ori_ori_n429_));
  OR2        o0401(.A(n), .B(m), .Y(ori_ori_n430_));
  NO2        o0402(.A(ori_ori_n430_), .B(ori_ori_n152_), .Y(ori_ori_n431_));
  NO2        o0403(.A(ori_ori_n182_), .B(ori_ori_n147_), .Y(ori_ori_n432_));
  OAI210     o0404(.A0(ori_ori_n431_), .A1(ori_ori_n175_), .B0(ori_ori_n432_), .Y(ori_ori_n433_));
  INV        o0405(.A(ori_ori_n366_), .Y(ori_ori_n434_));
  NA3        o0406(.A(ori_ori_n434_), .B(ori_ori_n354_), .C(d), .Y(ori_ori_n435_));
  NO2        o0407(.A(ori_ori_n420_), .B(ori_ori_n49_), .Y(ori_ori_n436_));
  NO3        o0408(.A(ori_ori_n66_), .B(ori_ori_n111_), .C(e), .Y(ori_ori_n437_));
  NAi21      o0409(.An(k), .B(j), .Y(ori_ori_n438_));
  NA3        o0410(.A(i), .B(ori_ori_n437_), .C(ori_ori_n436_), .Y(ori_ori_n439_));
  NAi21      o0411(.An(e), .B(d), .Y(ori_ori_n440_));
  INV        o0412(.A(ori_ori_n440_), .Y(ori_ori_n441_));
  NO2        o0413(.A(ori_ori_n256_), .B(ori_ori_n215_), .Y(ori_ori_n442_));
  NA3        o0414(.A(ori_ori_n442_), .B(ori_ori_n441_), .C(ori_ori_n228_), .Y(ori_ori_n443_));
  NA4        o0415(.A(ori_ori_n443_), .B(ori_ori_n439_), .C(ori_ori_n435_), .D(ori_ori_n433_), .Y(ori_ori_n444_));
  NO2        o0416(.A(ori_ori_n332_), .B(ori_ori_n215_), .Y(ori_ori_n445_));
  NA2        o0417(.A(ori_ori_n445_), .B(ori_ori_n441_), .Y(ori_ori_n446_));
  NOi31      o0418(.An(n), .B(m), .C(k), .Y(ori_ori_n447_));
  AOI220     o0419(.A0(ori_ori_n447_), .A1(ori_ori_n381_), .B0(ori_ori_n223_), .B1(ori_ori_n50_), .Y(ori_ori_n448_));
  NAi31      o0420(.An(g), .B(f), .C(c), .Y(ori_ori_n449_));
  OR3        o0421(.A(ori_ori_n449_), .B(ori_ori_n448_), .C(e), .Y(ori_ori_n450_));
  NA3        o0422(.A(ori_ori_n450_), .B(ori_ori_n446_), .C(ori_ori_n307_), .Y(ori_ori_n451_));
  NO3        o0423(.A(ori_ori_n451_), .B(ori_ori_n444_), .C(ori_ori_n269_), .Y(ori_ori_n452_));
  NOi32      o0424(.An(c), .Bn(a), .C(b), .Y(ori_ori_n453_));
  NA2        o0425(.A(ori_ori_n453_), .B(ori_ori_n112_), .Y(ori_ori_n454_));
  INV        o0426(.A(ori_ori_n277_), .Y(ori_ori_n455_));
  AN2        o0427(.A(e), .B(d), .Y(ori_ori_n456_));
  NA2        o0428(.A(ori_ori_n456_), .B(ori_ori_n455_), .Y(ori_ori_n457_));
  INV        o0429(.A(ori_ori_n147_), .Y(ori_ori_n458_));
  NO2        o0430(.A(ori_ori_n129_), .B(ori_ori_n41_), .Y(ori_ori_n459_));
  NO2        o0431(.A(ori_ori_n66_), .B(e), .Y(ori_ori_n460_));
  NOi31      o0432(.An(j), .B(k), .C(i), .Y(ori_ori_n461_));
  NOi21      o0433(.An(ori_ori_n165_), .B(ori_ori_n461_), .Y(ori_ori_n462_));
  NA3        o0434(.A(ori_ori_n321_), .B(ori_ori_n462_), .C(ori_ori_n264_), .Y(ori_ori_n463_));
  AOI220     o0435(.A0(ori_ori_n463_), .A1(ori_ori_n460_), .B0(ori_ori_n459_), .B1(ori_ori_n458_), .Y(ori_ori_n464_));
  AOI210     o0436(.A0(ori_ori_n464_), .A1(ori_ori_n457_), .B0(ori_ori_n454_), .Y(ori_ori_n465_));
  NO2        o0437(.A(ori_ori_n211_), .B(ori_ori_n206_), .Y(ori_ori_n466_));
  NOi21      o0438(.An(a), .B(b), .Y(ori_ori_n467_));
  NA3        o0439(.A(e), .B(d), .C(c), .Y(ori_ori_n468_));
  NAi21      o0440(.An(ori_ori_n468_), .B(ori_ori_n467_), .Y(ori_ori_n469_));
  NO2        o0441(.A(ori_ori_n419_), .B(ori_ori_n205_), .Y(ori_ori_n470_));
  NOi21      o0442(.An(ori_ori_n469_), .B(ori_ori_n470_), .Y(ori_ori_n471_));
  AOI210     o0443(.A0(ori_ori_n272_), .A1(ori_ori_n466_), .B0(ori_ori_n471_), .Y(ori_ori_n472_));
  NO4        o0444(.A(ori_ori_n188_), .B(ori_ori_n101_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n473_));
  NA2        o0445(.A(ori_ori_n376_), .B(ori_ori_n153_), .Y(ori_ori_n474_));
  OR2        o0446(.A(k), .B(j), .Y(ori_ori_n475_));
  NA2        o0447(.A(l), .B(k), .Y(ori_ori_n476_));
  NA3        o0448(.A(ori_ori_n476_), .B(ori_ori_n475_), .C(ori_ori_n223_), .Y(ori_ori_n477_));
  AOI210     o0449(.A0(ori_ori_n235_), .A1(ori_ori_n335_), .B0(ori_ori_n81_), .Y(ori_ori_n478_));
  NOi21      o0450(.An(ori_ori_n477_), .B(ori_ori_n478_), .Y(ori_ori_n479_));
  OR3        o0451(.A(ori_ori_n479_), .B(ori_ori_n143_), .C(ori_ori_n133_), .Y(ori_ori_n480_));
  NA2        o0452(.A(ori_ori_n126_), .B(ori_ori_n124_), .Y(ori_ori_n481_));
  NO3        o0453(.A(ori_ori_n419_), .B(ori_ori_n89_), .C(ori_ori_n129_), .Y(ori_ori_n482_));
  NO3        o0454(.A(ori_ori_n482_), .B(ori_ori_n481_), .C(ori_ori_n322_), .Y(ori_ori_n483_));
  NA3        o0455(.A(ori_ori_n483_), .B(ori_ori_n480_), .C(ori_ori_n474_), .Y(ori_ori_n484_));
  NO4        o0456(.A(ori_ori_n484_), .B(ori_ori_n473_), .C(ori_ori_n472_), .D(ori_ori_n465_), .Y(ori_ori_n485_));
  NOi21      o0457(.An(d), .B(e), .Y(ori_ori_n486_));
  NO2        o0458(.A(ori_ori_n188_), .B(ori_ori_n56_), .Y(ori_ori_n487_));
  NAi31      o0459(.An(j), .B(l), .C(i), .Y(ori_ori_n488_));
  INV        o0460(.A(ori_ori_n101_), .Y(ori_ori_n489_));
  NA3        o0461(.A(ori_ori_n489_), .B(ori_ori_n487_), .C(ori_ori_n486_), .Y(ori_ori_n490_));
  NO3        o0462(.A(ori_ori_n390_), .B(ori_ori_n341_), .C(ori_ori_n202_), .Y(ori_ori_n491_));
  NO2        o0463(.A(ori_ori_n390_), .B(ori_ori_n366_), .Y(ori_ori_n492_));
  NO4        o0464(.A(ori_ori_n492_), .B(ori_ori_n491_), .C(ori_ori_n184_), .D(ori_ori_n304_), .Y(ori_ori_n493_));
  NA3        o0465(.A(ori_ori_n493_), .B(ori_ori_n490_), .C(ori_ori_n244_), .Y(ori_ori_n494_));
  OAI210     o0466(.A0(ori_ori_n125_), .A1(ori_ori_n123_), .B0(n), .Y(ori_ori_n495_));
  NO2        o0467(.A(ori_ori_n495_), .B(ori_ori_n129_), .Y(ori_ori_n496_));
  OR2        o0468(.A(ori_ori_n296_), .B(ori_ori_n246_), .Y(ori_ori_n497_));
  OA210      o0469(.A0(ori_ori_n497_), .A1(ori_ori_n496_), .B0(ori_ori_n193_), .Y(ori_ori_n498_));
  XO2        o0470(.A(i), .B(h), .Y(ori_ori_n499_));
  NA3        o0471(.A(ori_ori_n499_), .B(ori_ori_n160_), .C(n), .Y(ori_ori_n500_));
  NAi41      o0472(.An(ori_ori_n296_), .B(ori_ori_n500_), .C(ori_ori_n448_), .D(ori_ori_n378_), .Y(ori_ori_n501_));
  NOi32      o0473(.An(ori_ori_n501_), .Bn(ori_ori_n460_), .C(ori_ori_n274_), .Y(ori_ori_n502_));
  NAi31      o0474(.An(c), .B(f), .C(d), .Y(ori_ori_n503_));
  AOI210     o0475(.A0(ori_ori_n280_), .A1(ori_ori_n196_), .B0(ori_ori_n503_), .Y(ori_ori_n504_));
  INV        o0476(.A(ori_ori_n504_), .Y(ori_ori_n505_));
  NA2        o0477(.A(ori_ori_n229_), .B(ori_ori_n107_), .Y(ori_ori_n506_));
  AOI210     o0478(.A0(ori_ori_n506_), .A1(ori_ori_n180_), .B0(ori_ori_n503_), .Y(ori_ori_n507_));
  AOI210     o0479(.A0(ori_ori_n352_), .A1(ori_ori_n35_), .B0(ori_ori_n469_), .Y(ori_ori_n508_));
  NO2        o0480(.A(ori_ori_n508_), .B(ori_ori_n507_), .Y(ori_ori_n509_));
  AO220      o0481(.A0(ori_ori_n288_), .A1(ori_ori_n267_), .B0(ori_ori_n166_), .B1(ori_ori_n67_), .Y(ori_ori_n510_));
  NA3        o0482(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n511_));
  NAi31      o0483(.An(ori_ori_n510_), .B(ori_ori_n509_), .C(ori_ori_n505_), .Y(ori_ori_n512_));
  NO4        o0484(.A(ori_ori_n512_), .B(ori_ori_n502_), .C(ori_ori_n498_), .D(ori_ori_n494_), .Y(ori_ori_n513_));
  NA4        o0485(.A(ori_ori_n513_), .B(ori_ori_n485_), .C(ori_ori_n452_), .D(ori_ori_n426_), .Y(ori11));
  NO2        o0486(.A(ori_ori_n72_), .B(f), .Y(ori_ori_n515_));
  NA2        o0487(.A(j), .B(g), .Y(ori_ori_n516_));
  NAi31      o0488(.An(i), .B(m), .C(l), .Y(ori_ori_n517_));
  NA3        o0489(.A(m), .B(k), .C(j), .Y(ori_ori_n518_));
  OAI220     o0490(.A0(ori_ori_n518_), .A1(ori_ori_n129_), .B0(ori_ori_n517_), .B1(ori_ori_n516_), .Y(ori_ori_n519_));
  NA2        o0491(.A(ori_ori_n519_), .B(ori_ori_n515_), .Y(ori_ori_n520_));
  NOi32      o0492(.An(e), .Bn(b), .C(f), .Y(ori_ori_n521_));
  NA2        o0493(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n522_));
  NO2        o0494(.A(ori_ori_n522_), .B(ori_ori_n298_), .Y(ori_ori_n523_));
  NAi31      o0495(.An(d), .B(e), .C(a), .Y(ori_ori_n524_));
  NO2        o0496(.A(ori_ori_n524_), .B(n), .Y(ori_ori_n525_));
  AOI220     o0497(.A0(ori_ori_n525_), .A1(ori_ori_n99_), .B0(ori_ori_n523_), .B1(ori_ori_n521_), .Y(ori_ori_n526_));
  NAi41      o0498(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n527_));
  AN2        o0499(.A(ori_ori_n527_), .B(ori_ori_n365_), .Y(ori_ori_n528_));
  AOI210     o0500(.A0(ori_ori_n528_), .A1(ori_ori_n390_), .B0(ori_ori_n275_), .Y(ori_ori_n529_));
  NA2        o0501(.A(j), .B(i), .Y(ori_ori_n530_));
  NAi31      o0502(.An(n), .B(m), .C(k), .Y(ori_ori_n531_));
  NO3        o0503(.A(ori_ori_n531_), .B(ori_ori_n530_), .C(ori_ori_n111_), .Y(ori_ori_n532_));
  NO4        o0504(.A(n), .B(d), .C(ori_ori_n115_), .D(a), .Y(ori_ori_n533_));
  OR2        o0505(.A(n), .B(c), .Y(ori_ori_n534_));
  NO2        o0506(.A(ori_ori_n534_), .B(ori_ori_n149_), .Y(ori_ori_n535_));
  NO2        o0507(.A(ori_ori_n535_), .B(ori_ori_n533_), .Y(ori_ori_n536_));
  NOi32      o0508(.An(g), .Bn(f), .C(i), .Y(ori_ori_n537_));
  AOI220     o0509(.A0(ori_ori_n537_), .A1(ori_ori_n97_), .B0(ori_ori_n519_), .B1(f), .Y(ori_ori_n538_));
  NO2        o0510(.A(ori_ori_n277_), .B(ori_ori_n49_), .Y(ori_ori_n539_));
  NO2        o0511(.A(ori_ori_n538_), .B(ori_ori_n536_), .Y(ori_ori_n540_));
  AOI210     o0512(.A0(ori_ori_n532_), .A1(ori_ori_n529_), .B0(ori_ori_n540_), .Y(ori_ori_n541_));
  NA2        o0513(.A(ori_ori_n139_), .B(ori_ori_n34_), .Y(ori_ori_n542_));
  OAI220     o0514(.A0(ori_ori_n542_), .A1(m), .B0(ori_ori_n522_), .B1(ori_ori_n235_), .Y(ori_ori_n543_));
  NOi41      o0515(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n544_));
  NAi32      o0516(.An(e), .Bn(b), .C(c), .Y(ori_ori_n545_));
  OR2        o0517(.A(ori_ori_n545_), .B(ori_ori_n81_), .Y(ori_ori_n546_));
  AN2        o0518(.A(ori_ori_n336_), .B(ori_ori_n318_), .Y(ori_ori_n547_));
  NA2        o0519(.A(ori_ori_n547_), .B(ori_ori_n546_), .Y(ori_ori_n548_));
  OA210      o0520(.A0(ori_ori_n548_), .A1(ori_ori_n544_), .B0(ori_ori_n543_), .Y(ori_ori_n549_));
  OAI220     o0521(.A0(ori_ori_n392_), .A1(ori_ori_n391_), .B0(ori_ori_n517_), .B1(ori_ori_n516_), .Y(ori_ori_n550_));
  NAi31      o0522(.An(d), .B(c), .C(a), .Y(ori_ori_n551_));
  NO2        o0523(.A(ori_ori_n551_), .B(n), .Y(ori_ori_n552_));
  NA3        o0524(.A(ori_ori_n552_), .B(ori_ori_n550_), .C(e), .Y(ori_ori_n553_));
  INV        o0525(.A(ori_ori_n553_), .Y(ori_ori_n554_));
  NO2        o0526(.A(ori_ori_n278_), .B(n), .Y(ori_ori_n555_));
  NO2        o0527(.A(ori_ori_n421_), .B(ori_ori_n555_), .Y(ori_ori_n556_));
  NA2        o0528(.A(ori_ori_n550_), .B(f), .Y(ori_ori_n557_));
  NAi32      o0529(.An(d), .Bn(a), .C(b), .Y(ori_ori_n558_));
  NO2        o0530(.A(ori_ori_n558_), .B(ori_ori_n49_), .Y(ori_ori_n559_));
  NA2        o0531(.A(h), .B(f), .Y(ori_ori_n560_));
  NO2        o0532(.A(ori_ori_n560_), .B(ori_ori_n92_), .Y(ori_ori_n561_));
  NA2        o0533(.A(ori_ori_n561_), .B(ori_ori_n559_), .Y(ori_ori_n562_));
  OAI210     o0534(.A0(ori_ori_n557_), .A1(ori_ori_n556_), .B0(ori_ori_n562_), .Y(ori_ori_n563_));
  NO2        o0535(.A(ori_ori_n146_), .B(c), .Y(ori_ori_n564_));
  NA3        o0536(.A(f), .B(d), .C(b), .Y(ori_ori_n565_));
  NO4        o0537(.A(ori_ori_n565_), .B(ori_ori_n176_), .C(ori_ori_n173_), .D(g), .Y(ori_ori_n566_));
  NO4        o0538(.A(ori_ori_n566_), .B(ori_ori_n563_), .C(ori_ori_n554_), .D(ori_ori_n549_), .Y(ori_ori_n567_));
  AN4        o0539(.A(ori_ori_n567_), .B(ori_ori_n541_), .C(ori_ori_n526_), .D(ori_ori_n520_), .Y(ori_ori_n568_));
  INV        o0540(.A(k), .Y(ori_ori_n569_));
  NA3        o0541(.A(l), .B(ori_ori_n569_), .C(i), .Y(ori_ori_n570_));
  INV        o0542(.A(ori_ori_n570_), .Y(ori_ori_n571_));
  NAi32      o0543(.An(h), .Bn(f), .C(g), .Y(ori_ori_n572_));
  NAi41      o0544(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n573_));
  OAI210     o0545(.A0(ori_ori_n524_), .A1(n), .B0(ori_ori_n573_), .Y(ori_ori_n574_));
  NA2        o0546(.A(ori_ori_n574_), .B(m), .Y(ori_ori_n575_));
  NAi31      o0547(.An(h), .B(g), .C(f), .Y(ori_ori_n576_));
  OR3        o0548(.A(ori_ori_n576_), .B(ori_ori_n278_), .C(ori_ori_n49_), .Y(ori_ori_n577_));
  NA4        o0549(.A(ori_ori_n412_), .B(ori_ori_n119_), .C(ori_ori_n112_), .D(e), .Y(ori_ori_n578_));
  AN2        o0550(.A(ori_ori_n578_), .B(ori_ori_n577_), .Y(ori_ori_n579_));
  OA210      o0551(.A0(ori_ori_n575_), .A1(ori_ori_n572_), .B0(ori_ori_n579_), .Y(ori_ori_n580_));
  NO3        o0552(.A(ori_ori_n572_), .B(ori_ori_n72_), .C(ori_ori_n73_), .Y(ori_ori_n581_));
  NO4        o0553(.A(ori_ori_n576_), .B(ori_ori_n534_), .C(ori_ori_n149_), .D(ori_ori_n73_), .Y(ori_ori_n582_));
  OR2        o0554(.A(ori_ori_n582_), .B(ori_ori_n581_), .Y(ori_ori_n583_));
  NAi21      o0555(.An(ori_ori_n583_), .B(ori_ori_n580_), .Y(ori_ori_n584_));
  NAi31      o0556(.An(f), .B(h), .C(g), .Y(ori_ori_n585_));
  NOi32      o0557(.An(b), .Bn(a), .C(c), .Y(ori_ori_n586_));
  NOi41      o0558(.An(ori_ori_n586_), .B(ori_ori_n347_), .C(ori_ori_n69_), .D(ori_ori_n116_), .Y(ori_ori_n587_));
  NOi32      o0559(.An(d), .Bn(a), .C(e), .Y(ori_ori_n588_));
  NA2        o0560(.A(ori_ori_n588_), .B(ori_ori_n112_), .Y(ori_ori_n589_));
  NO2        o0561(.A(n), .B(c), .Y(ori_ori_n590_));
  NA3        o0562(.A(ori_ori_n590_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n591_));
  NAi32      o0563(.An(n), .Bn(f), .C(m), .Y(ori_ori_n592_));
  NA3        o0564(.A(ori_ori_n592_), .B(ori_ori_n591_), .C(ori_ori_n589_), .Y(ori_ori_n593_));
  NOi32      o0565(.An(e), .Bn(a), .C(d), .Y(ori_ori_n594_));
  AOI210     o0566(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n594_), .Y(ori_ori_n595_));
  AOI210     o0567(.A0(ori_ori_n595_), .A1(ori_ori_n215_), .B0(ori_ori_n542_), .Y(ori_ori_n596_));
  AOI210     o0568(.A0(ori_ori_n596_), .A1(ori_ori_n593_), .B0(ori_ori_n587_), .Y(ori_ori_n597_));
  OAI210     o0569(.A0(ori_ori_n251_), .A1(ori_ori_n84_), .B0(ori_ori_n597_), .Y(ori_ori_n598_));
  AOI210     o0570(.A0(ori_ori_n584_), .A1(ori_ori_n571_), .B0(ori_ori_n598_), .Y(ori_ori_n599_));
  NO3        o0571(.A(ori_ori_n316_), .B(ori_ori_n61_), .C(n), .Y(ori_ori_n600_));
  NA3        o0572(.A(ori_ori_n503_), .B(ori_ori_n171_), .C(ori_ori_n170_), .Y(ori_ori_n601_));
  NA2        o0573(.A(ori_ori_n449_), .B(ori_ori_n232_), .Y(ori_ori_n602_));
  OR2        o0574(.A(ori_ori_n602_), .B(ori_ori_n601_), .Y(ori_ori_n603_));
  NA2        o0575(.A(ori_ori_n603_), .B(ori_ori_n600_), .Y(ori_ori_n604_));
  NO2        o0576(.A(ori_ori_n604_), .B(ori_ori_n84_), .Y(ori_ori_n605_));
  NA3        o0577(.A(ori_ori_n544_), .B(ori_ori_n337_), .C(ori_ori_n46_), .Y(ori_ori_n606_));
  NOi32      o0578(.An(e), .Bn(c), .C(f), .Y(ori_ori_n607_));
  NOi21      o0579(.An(f), .B(g), .Y(ori_ori_n608_));
  NO2        o0580(.A(ori_ori_n608_), .B(ori_ori_n213_), .Y(ori_ori_n609_));
  AOI220     o0581(.A0(ori_ori_n609_), .A1(ori_ori_n386_), .B0(ori_ori_n607_), .B1(ori_ori_n175_), .Y(ori_ori_n610_));
  NA3        o0582(.A(ori_ori_n610_), .B(ori_ori_n606_), .C(ori_ori_n178_), .Y(ori_ori_n611_));
  AOI210     o0583(.A0(ori_ori_n528_), .A1(ori_ori_n390_), .B0(ori_ori_n297_), .Y(ori_ori_n612_));
  NOi21      o0584(.An(j), .B(l), .Y(ori_ori_n613_));
  NAi21      o0585(.An(k), .B(h), .Y(ori_ori_n614_));
  NO2        o0586(.A(ori_ori_n614_), .B(ori_ori_n266_), .Y(ori_ori_n615_));
  NA2        o0587(.A(ori_ori_n615_), .B(ori_ori_n613_), .Y(ori_ori_n616_));
  OR2        o0588(.A(ori_ori_n616_), .B(ori_ori_n575_), .Y(ori_ori_n617_));
  NOi31      o0589(.An(m), .B(n), .C(k), .Y(ori_ori_n618_));
  NA2        o0590(.A(ori_ori_n613_), .B(ori_ori_n618_), .Y(ori_ori_n619_));
  AOI210     o0591(.A0(ori_ori_n390_), .A1(ori_ori_n365_), .B0(ori_ori_n297_), .Y(ori_ori_n620_));
  NAi21      o0592(.An(ori_ori_n619_), .B(ori_ori_n620_), .Y(ori_ori_n621_));
  NO2        o0593(.A(ori_ori_n278_), .B(ori_ori_n49_), .Y(ori_ori_n622_));
  NO2        o0594(.A(ori_ori_n309_), .B(ori_ori_n585_), .Y(ori_ori_n623_));
  NO2        o0595(.A(ori_ori_n524_), .B(ori_ori_n49_), .Y(ori_ori_n624_));
  AOI220     o0596(.A0(ori_ori_n624_), .A1(ori_ori_n623_), .B0(ori_ori_n622_), .B1(ori_ori_n561_), .Y(ori_ori_n625_));
  NA3        o0597(.A(ori_ori_n625_), .B(ori_ori_n621_), .C(ori_ori_n617_), .Y(ori_ori_n626_));
  NA2        o0598(.A(ori_ori_n107_), .B(ori_ori_n36_), .Y(ori_ori_n627_));
  NO2        o0599(.A(k), .B(ori_ori_n216_), .Y(ori_ori_n628_));
  INV        o0600(.A(ori_ori_n354_), .Y(ori_ori_n629_));
  NO2        o0601(.A(ori_ori_n629_), .B(n), .Y(ori_ori_n630_));
  NAi31      o0602(.An(ori_ori_n627_), .B(ori_ori_n630_), .C(ori_ori_n628_), .Y(ori_ori_n631_));
  NO2        o0603(.A(ori_ori_n522_), .B(ori_ori_n176_), .Y(ori_ori_n632_));
  NA3        o0604(.A(ori_ori_n545_), .B(ori_ori_n274_), .C(ori_ori_n144_), .Y(ori_ori_n633_));
  NA2        o0605(.A(ori_ori_n499_), .B(ori_ori_n160_), .Y(ori_ori_n634_));
  NO3        o0606(.A(ori_ori_n387_), .B(ori_ori_n634_), .C(ori_ori_n84_), .Y(ori_ori_n635_));
  AOI210     o0607(.A0(ori_ori_n633_), .A1(ori_ori_n632_), .B0(ori_ori_n635_), .Y(ori_ori_n636_));
  AN3        o0608(.A(f), .B(d), .C(b), .Y(ori_ori_n637_));
  OAI210     o0609(.A0(ori_ori_n637_), .A1(ori_ori_n128_), .B0(n), .Y(ori_ori_n638_));
  NA3        o0610(.A(ori_ori_n499_), .B(ori_ori_n160_), .C(ori_ori_n216_), .Y(ori_ori_n639_));
  AOI210     o0611(.A0(ori_ori_n638_), .A1(ori_ori_n234_), .B0(ori_ori_n639_), .Y(ori_ori_n640_));
  NAi31      o0612(.An(m), .B(n), .C(k), .Y(ori_ori_n641_));
  INV        o0613(.A(ori_ori_n253_), .Y(ori_ori_n642_));
  OAI210     o0614(.A0(ori_ori_n642_), .A1(ori_ori_n640_), .B0(j), .Y(ori_ori_n643_));
  NA3        o0615(.A(ori_ori_n643_), .B(ori_ori_n636_), .C(ori_ori_n631_), .Y(ori_ori_n644_));
  NO4        o0616(.A(ori_ori_n644_), .B(ori_ori_n626_), .C(ori_ori_n611_), .D(ori_ori_n605_), .Y(ori_ori_n645_));
  NAi31      o0617(.An(g), .B(h), .C(f), .Y(ori_ori_n646_));
  OR3        o0618(.A(ori_ori_n646_), .B(ori_ori_n278_), .C(n), .Y(ori_ori_n647_));
  OA210      o0619(.A0(ori_ori_n524_), .A1(n), .B0(ori_ori_n573_), .Y(ori_ori_n648_));
  NA3        o0620(.A(ori_ori_n410_), .B(ori_ori_n119_), .C(ori_ori_n81_), .Y(ori_ori_n649_));
  OAI210     o0621(.A0(ori_ori_n648_), .A1(ori_ori_n88_), .B0(ori_ori_n649_), .Y(ori_ori_n650_));
  NOi21      o0622(.An(ori_ori_n647_), .B(ori_ori_n650_), .Y(ori_ori_n651_));
  NO2        o0623(.A(ori_ori_n651_), .B(ori_ori_n518_), .Y(ori_ori_n652_));
  NO3        o0624(.A(g), .B(ori_ori_n215_), .C(ori_ori_n56_), .Y(ori_ori_n653_));
  NAi21      o0625(.An(h), .B(j), .Y(ori_ori_n654_));
  NO2        o0626(.A(ori_ori_n506_), .B(ori_ori_n84_), .Y(ori_ori_n655_));
  OAI210     o0627(.A0(ori_ori_n655_), .A1(ori_ori_n386_), .B0(ori_ori_n653_), .Y(ori_ori_n656_));
  OR2        o0628(.A(ori_ori_n72_), .B(ori_ori_n73_), .Y(ori_ori_n657_));
  NA2        o0629(.A(ori_ori_n586_), .B(ori_ori_n339_), .Y(ori_ori_n658_));
  OA220      o0630(.A0(ori_ori_n619_), .A1(ori_ori_n658_), .B0(ori_ori_n616_), .B1(ori_ori_n657_), .Y(ori_ori_n659_));
  NA3        o0631(.A(ori_ori_n515_), .B(ori_ori_n97_), .C(ori_ori_n96_), .Y(ori_ori_n660_));
  AN2        o0632(.A(h), .B(f), .Y(ori_ori_n661_));
  NA2        o0633(.A(ori_ori_n661_), .B(ori_ori_n37_), .Y(ori_ori_n662_));
  NA2        o0634(.A(ori_ori_n97_), .B(ori_ori_n46_), .Y(ori_ori_n663_));
  OAI220     o0635(.A0(ori_ori_n663_), .A1(ori_ori_n329_), .B0(ori_ori_n662_), .B1(ori_ori_n454_), .Y(ori_ori_n664_));
  AOI210     o0636(.A0(ori_ori_n558_), .A1(ori_ori_n420_), .B0(ori_ori_n49_), .Y(ori_ori_n665_));
  INV        o0637(.A(ori_ori_n664_), .Y(ori_ori_n666_));
  NA4        o0638(.A(ori_ori_n666_), .B(ori_ori_n660_), .C(ori_ori_n659_), .D(ori_ori_n656_), .Y(ori_ori_n667_));
  NA2        o0639(.A(ori_ori_n130_), .B(ori_ori_n49_), .Y(ori_ori_n668_));
  NA2        o0640(.A(ori_ori_n354_), .B(ori_ori_n112_), .Y(ori_ori_n669_));
  OA220      o0641(.A0(ori_ori_n669_), .A1(ori_ori_n542_), .B0(ori_ori_n352_), .B1(ori_ori_n110_), .Y(ori_ori_n670_));
  INV        o0642(.A(ori_ori_n670_), .Y(ori_ori_n671_));
  NO3        o0643(.A(ori_ori_n397_), .B(ori_ori_n193_), .C(ori_ori_n192_), .Y(ori_ori_n672_));
  NA2        o0644(.A(ori_ori_n672_), .B(ori_ori_n232_), .Y(ori_ori_n673_));
  NA3        o0645(.A(ori_ori_n673_), .B(ori_ori_n257_), .C(j), .Y(ori_ori_n674_));
  NO3        o0646(.A(ori_ori_n449_), .B(ori_ori_n173_), .C(i), .Y(ori_ori_n675_));
  NA2        o0647(.A(ori_ori_n453_), .B(ori_ori_n81_), .Y(ori_ori_n676_));
  NA2        o0648(.A(ori_ori_n674_), .B(ori_ori_n395_), .Y(ori_ori_n677_));
  NO4        o0649(.A(ori_ori_n677_), .B(ori_ori_n671_), .C(ori_ori_n667_), .D(ori_ori_n652_), .Y(ori_ori_n678_));
  NA4        o0650(.A(ori_ori_n678_), .B(ori_ori_n645_), .C(ori_ori_n599_), .D(ori_ori_n568_), .Y(ori08));
  NO2        o0651(.A(k), .B(h), .Y(ori_ori_n680_));
  AO210      o0652(.A0(ori_ori_n255_), .A1(ori_ori_n438_), .B0(ori_ori_n680_), .Y(ori_ori_n681_));
  NO2        o0653(.A(ori_ori_n681_), .B(ori_ori_n295_), .Y(ori_ori_n682_));
  NA2        o0654(.A(ori_ori_n607_), .B(ori_ori_n81_), .Y(ori_ori_n683_));
  NA2        o0655(.A(ori_ori_n683_), .B(ori_ori_n449_), .Y(ori_ori_n684_));
  AOI210     o0656(.A0(ori_ori_n684_), .A1(ori_ori_n682_), .B0(ori_ori_n482_), .Y(ori_ori_n685_));
  NA2        o0657(.A(ori_ori_n81_), .B(ori_ori_n109_), .Y(ori_ori_n686_));
  NO2        o0658(.A(ori_ori_n686_), .B(ori_ori_n57_), .Y(ori_ori_n687_));
  NO4        o0659(.A(ori_ori_n372_), .B(ori_ori_n111_), .C(j), .D(ori_ori_n216_), .Y(ori_ori_n688_));
  NA2        o0660(.A(ori_ori_n688_), .B(ori_ori_n687_), .Y(ori_ori_n689_));
  AOI210     o0661(.A0(ori_ori_n565_), .A1(ori_ori_n156_), .B0(ori_ori_n81_), .Y(ori_ori_n690_));
  NA4        o0662(.A(ori_ori_n218_), .B(ori_ori_n139_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n691_));
  AN2        o0663(.A(l), .B(k), .Y(ori_ori_n692_));
  NA4        o0664(.A(ori_ori_n692_), .B(ori_ori_n107_), .C(ori_ori_n73_), .D(ori_ori_n216_), .Y(ori_ori_n693_));
  OAI210     o0665(.A0(ori_ori_n691_), .A1(g), .B0(ori_ori_n693_), .Y(ori_ori_n694_));
  NA2        o0666(.A(ori_ori_n694_), .B(ori_ori_n690_), .Y(ori_ori_n695_));
  NA4        o0667(.A(ori_ori_n695_), .B(ori_ori_n689_), .C(ori_ori_n685_), .D(ori_ori_n343_), .Y(ori_ori_n696_));
  AN2        o0668(.A(ori_ori_n525_), .B(ori_ori_n93_), .Y(ori_ori_n697_));
  NO2        o0669(.A(ori_ori_n38_), .B(ori_ori_n215_), .Y(ori_ori_n698_));
  AOI220     o0670(.A0(ori_ori_n609_), .A1(ori_ori_n342_), .B0(ori_ori_n698_), .B1(ori_ori_n555_), .Y(ori_ori_n699_));
  NAi21      o0671(.An(ori_ori_n697_), .B(ori_ori_n699_), .Y(ori_ori_n700_));
  NO2        o0672(.A(ori_ori_n528_), .B(ori_ori_n35_), .Y(ori_ori_n701_));
  INV        o0673(.A(ori_ori_n701_), .Y(ori_ori_n702_));
  NO3        o0674(.A(ori_ori_n316_), .B(ori_ori_n129_), .C(ori_ori_n41_), .Y(ori_ori_n703_));
  NAi21      o0675(.An(ori_ori_n703_), .B(ori_ori_n693_), .Y(ori_ori_n704_));
  NA2        o0676(.A(ori_ori_n681_), .B(ori_ori_n134_), .Y(ori_ori_n705_));
  AOI220     o0677(.A0(ori_ori_n705_), .A1(ori_ori_n396_), .B0(ori_ori_n704_), .B1(ori_ori_n76_), .Y(ori_ori_n706_));
  OAI210     o0678(.A0(ori_ori_n702_), .A1(ori_ori_n84_), .B0(ori_ori_n706_), .Y(ori_ori_n707_));
  NA2        o0679(.A(ori_ori_n354_), .B(ori_ori_n43_), .Y(ori_ori_n708_));
  NA3        o0680(.A(ori_ori_n673_), .B(ori_ori_n331_), .C(ori_ori_n377_), .Y(ori_ori_n709_));
  NA3        o0681(.A(m), .B(l), .C(k), .Y(ori_ori_n710_));
  AOI210     o0682(.A0(ori_ori_n649_), .A1(ori_ori_n647_), .B0(ori_ori_n710_), .Y(ori_ori_n711_));
  NA3        o0683(.A(ori_ori_n112_), .B(k), .C(ori_ori_n84_), .Y(ori_ori_n712_));
  INV        o0684(.A(ori_ori_n711_), .Y(ori_ori_n713_));
  NA3        o0685(.A(ori_ori_n713_), .B(ori_ori_n709_), .C(ori_ori_n708_), .Y(ori_ori_n714_));
  NO4        o0686(.A(ori_ori_n714_), .B(ori_ori_n707_), .C(ori_ori_n700_), .D(ori_ori_n696_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n609_), .B(ori_ori_n386_), .Y(ori_ori_n716_));
  NOi31      o0688(.An(g), .B(h), .C(f), .Y(ori_ori_n717_));
  NA2        o0689(.A(ori_ori_n624_), .B(ori_ori_n717_), .Y(ori_ori_n718_));
  AO210      o0690(.A0(ori_ori_n718_), .A1(ori_ori_n577_), .B0(ori_ori_n530_), .Y(ori_ori_n719_));
  NO3        o0691(.A(ori_ori_n390_), .B(ori_ori_n516_), .C(h), .Y(ori_ori_n720_));
  NA2        o0692(.A(ori_ori_n720_), .B(ori_ori_n112_), .Y(ori_ori_n721_));
  NA4        o0693(.A(ori_ori_n721_), .B(ori_ori_n719_), .C(ori_ori_n716_), .D(ori_ori_n254_), .Y(ori_ori_n722_));
  NA2        o0694(.A(ori_ori_n692_), .B(ori_ori_n73_), .Y(ori_ori_n723_));
  NO4        o0695(.A(ori_ori_n672_), .B(ori_ori_n173_), .C(n), .D(i), .Y(ori_ori_n724_));
  NOi21      o0696(.An(h), .B(j), .Y(ori_ori_n725_));
  NA2        o0697(.A(ori_ori_n725_), .B(f), .Y(ori_ori_n726_));
  NO2        o0698(.A(ori_ori_n726_), .B(ori_ori_n248_), .Y(ori_ori_n727_));
  NO3        o0699(.A(ori_ori_n727_), .B(ori_ori_n724_), .C(ori_ori_n675_), .Y(ori_ori_n728_));
  OAI220     o0700(.A0(ori_ori_n728_), .A1(ori_ori_n723_), .B0(ori_ori_n579_), .B1(ori_ori_n62_), .Y(ori_ori_n729_));
  AOI210     o0701(.A0(ori_ori_n722_), .A1(l), .B0(ori_ori_n729_), .Y(ori_ori_n730_));
  NO2        o0702(.A(j), .B(i), .Y(ori_ori_n731_));
  NA3        o0703(.A(ori_ori_n731_), .B(ori_ori_n79_), .C(l), .Y(ori_ori_n732_));
  NA2        o0704(.A(ori_ori_n731_), .B(ori_ori_n33_), .Y(ori_ori_n733_));
  NA2        o0705(.A(ori_ori_n415_), .B(ori_ori_n119_), .Y(ori_ori_n734_));
  OA220      o0706(.A0(ori_ori_n734_), .A1(ori_ori_n733_), .B0(ori_ori_n732_), .B1(ori_ori_n575_), .Y(ori_ori_n735_));
  NO3        o0707(.A(ori_ori_n151_), .B(ori_ori_n49_), .C(ori_ori_n109_), .Y(ori_ori_n736_));
  NO3        o0708(.A(ori_ori_n534_), .B(ori_ori_n149_), .C(ori_ori_n73_), .Y(ori_ori_n737_));
  NO3        o0709(.A(ori_ori_n476_), .B(ori_ori_n429_), .C(j), .Y(ori_ori_n738_));
  NA2        o0710(.A(ori_ori_n737_), .B(ori_ori_n738_), .Y(ori_ori_n739_));
  OAI210     o0711(.A0(ori_ori_n718_), .A1(ori_ori_n62_), .B0(ori_ori_n739_), .Y(ori_ori_n740_));
  AOI210     o0712(.A0(ori_ori_n521_), .A1(n), .B0(ori_ori_n544_), .Y(ori_ori_n741_));
  NA2        o0713(.A(ori_ori_n741_), .B(ori_ori_n547_), .Y(ori_ori_n742_));
  NO3        o0714(.A(ori_ori_n173_), .B(ori_ori_n385_), .C(ori_ori_n111_), .Y(ori_ori_n743_));
  AOI220     o0715(.A0(ori_ori_n743_), .A1(ori_ori_n249_), .B0(ori_ori_n602_), .B1(ori_ori_n306_), .Y(ori_ori_n744_));
  INV        o0716(.A(ori_ori_n744_), .Y(ori_ori_n745_));
  NO2        o0717(.A(ori_ori_n295_), .B(ori_ori_n134_), .Y(ori_ori_n746_));
  AOI220     o0718(.A0(ori_ori_n746_), .A1(ori_ori_n609_), .B0(ori_ori_n703_), .B1(ori_ori_n690_), .Y(ori_ori_n747_));
  NO2        o0719(.A(ori_ori_n710_), .B(ori_ori_n88_), .Y(ori_ori_n748_));
  NA2        o0720(.A(ori_ori_n748_), .B(ori_ori_n574_), .Y(ori_ori_n749_));
  NO2        o0721(.A(ori_ori_n576_), .B(ori_ori_n116_), .Y(ori_ori_n750_));
  OAI210     o0722(.A0(ori_ori_n750_), .A1(ori_ori_n738_), .B0(ori_ori_n665_), .Y(ori_ori_n751_));
  NA3        o0723(.A(ori_ori_n751_), .B(ori_ori_n749_), .C(ori_ori_n747_), .Y(ori_ori_n752_));
  OR3        o0724(.A(ori_ori_n752_), .B(ori_ori_n745_), .C(ori_ori_n740_), .Y(ori_ori_n753_));
  NA3        o0725(.A(ori_ori_n741_), .B(ori_ori_n547_), .C(ori_ori_n546_), .Y(ori_ori_n754_));
  NA4        o0726(.A(ori_ori_n754_), .B(ori_ori_n218_), .C(ori_ori_n438_), .D(ori_ori_n34_), .Y(ori_ori_n755_));
  NO4        o0727(.A(ori_ori_n476_), .B(ori_ori_n427_), .C(j), .D(f), .Y(ori_ori_n756_));
  OAI220     o0728(.A0(ori_ori_n691_), .A1(ori_ori_n683_), .B0(ori_ori_n329_), .B1(ori_ori_n38_), .Y(ori_ori_n757_));
  AOI210     o0729(.A0(ori_ori_n756_), .A1(ori_ori_n261_), .B0(ori_ori_n757_), .Y(ori_ori_n758_));
  NA3        o0730(.A(ori_ori_n537_), .B(ori_ori_n292_), .C(h), .Y(ori_ori_n759_));
  NO2        o0731(.A(ori_ori_n89_), .B(ori_ori_n47_), .Y(ori_ori_n760_));
  OAI220     o0732(.A0(ori_ori_n759_), .A1(ori_ori_n591_), .B0(ori_ori_n732_), .B1(ori_ori_n657_), .Y(ori_ori_n761_));
  AOI210     o0733(.A0(ori_ori_n760_), .A1(ori_ori_n630_), .B0(ori_ori_n761_), .Y(ori_ori_n762_));
  NA3        o0734(.A(ori_ori_n762_), .B(ori_ori_n758_), .C(ori_ori_n755_), .Y(ori_ori_n763_));
  BUFFER     o0735(.A(ori_ori_n748_), .Y(ori_ori_n764_));
  AOI220     o0736(.A0(ori_ori_n764_), .A1(ori_ori_n240_), .B0(ori_ori_n738_), .B1(ori_ori_n622_), .Y(ori_ori_n765_));
  NO2        o0737(.A(ori_ori_n648_), .B(ori_ori_n73_), .Y(ori_ori_n766_));
  AOI210     o0738(.A0(ori_ori_n756_), .A1(ori_ori_n766_), .B0(ori_ori_n333_), .Y(ori_ori_n767_));
  OAI210     o0739(.A0(ori_ori_n710_), .A1(ori_ori_n646_), .B0(ori_ori_n511_), .Y(ori_ori_n768_));
  NA3        o0740(.A(ori_ori_n252_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n769_));
  AOI220     o0741(.A0(ori_ori_n590_), .A1(ori_ori_n29_), .B0(ori_ori_n453_), .B1(ori_ori_n81_), .Y(ori_ori_n770_));
  NA2        o0742(.A(ori_ori_n770_), .B(ori_ori_n769_), .Y(ori_ori_n771_));
  NA2        o0743(.A(ori_ori_n771_), .B(ori_ori_n768_), .Y(ori_ori_n772_));
  NA3        o0744(.A(ori_ori_n772_), .B(ori_ori_n767_), .C(ori_ori_n765_), .Y(ori_ori_n773_));
  NOi41      o0745(.An(ori_ori_n735_), .B(ori_ori_n773_), .C(ori_ori_n763_), .D(ori_ori_n753_), .Y(ori_ori_n774_));
  OR2        o0746(.A(ori_ori_n691_), .B(ori_ori_n234_), .Y(ori_ori_n775_));
  NO3        o0747(.A(ori_ori_n338_), .B(ori_ori_n297_), .C(ori_ori_n111_), .Y(ori_ori_n776_));
  NA2        o0748(.A(ori_ori_n776_), .B(ori_ori_n742_), .Y(ori_ori_n777_));
  NO3        o0749(.A(ori_ori_n516_), .B(ori_ori_n91_), .C(h), .Y(ori_ori_n778_));
  NA2        o0750(.A(ori_ori_n778_), .B(ori_ori_n687_), .Y(ori_ori_n779_));
  NA4        o0751(.A(ori_ori_n779_), .B(ori_ori_n777_), .C(ori_ori_n775_), .D(ori_ori_n398_), .Y(ori_ori_n780_));
  OR2        o0752(.A(ori_ori_n646_), .B(ori_ori_n89_), .Y(ori_ori_n781_));
  NOi31      o0753(.An(b), .B(d), .C(a), .Y(ori_ori_n782_));
  NO2        o0754(.A(ori_ori_n782_), .B(ori_ori_n588_), .Y(ori_ori_n783_));
  NO2        o0755(.A(ori_ori_n783_), .B(n), .Y(ori_ori_n784_));
  NOi21      o0756(.An(ori_ori_n770_), .B(ori_ori_n784_), .Y(ori_ori_n785_));
  OAI220     o0757(.A0(ori_ori_n785_), .A1(ori_ori_n781_), .B0(ori_ori_n759_), .B1(ori_ori_n589_), .Y(ori_ori_n786_));
  NO2        o0758(.A(ori_ori_n545_), .B(ori_ori_n81_), .Y(ori_ori_n787_));
  NO3        o0759(.A(ori_ori_n608_), .B(ori_ori_n326_), .C(ori_ori_n116_), .Y(ori_ori_n788_));
  NOi21      o0760(.An(ori_ori_n788_), .B(ori_ori_n161_), .Y(ori_ori_n789_));
  AOI210     o0761(.A0(ori_ori_n776_), .A1(ori_ori_n787_), .B0(ori_ori_n789_), .Y(ori_ori_n790_));
  OAI210     o0762(.A0(ori_ori_n691_), .A1(ori_ori_n387_), .B0(ori_ori_n790_), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n672_), .B(n), .Y(ori_ori_n792_));
  AOI220     o0764(.A0(ori_ori_n746_), .A1(ori_ori_n653_), .B0(ori_ori_n792_), .B1(ori_ori_n682_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n323_), .B(ori_ori_n239_), .Y(ori_ori_n794_));
  OAI210     o0766(.A0(ori_ori_n93_), .A1(ori_ori_n90_), .B0(ori_ori_n794_), .Y(ori_ori_n795_));
  NA2        o0767(.A(ori_ori_n119_), .B(ori_ori_n81_), .Y(ori_ori_n796_));
  INV        o0768(.A(ori_ori_n795_), .Y(ori_ori_n797_));
  NO2        o0769(.A(ori_ori_n275_), .B(i), .Y(ori_ori_n798_));
  OAI210     o0770(.A0(ori_ori_n582_), .A1(ori_ori_n581_), .B0(ori_ori_n355_), .Y(ori_ori_n799_));
  NAi31      o0771(.An(ori_ori_n797_), .B(ori_ori_n799_), .C(ori_ori_n793_), .Y(ori_ori_n800_));
  NO4        o0772(.A(ori_ori_n800_), .B(ori_ori_n791_), .C(ori_ori_n786_), .D(ori_ori_n780_), .Y(ori_ori_n801_));
  NA4        o0773(.A(ori_ori_n801_), .B(ori_ori_n774_), .C(ori_ori_n730_), .D(ori_ori_n715_), .Y(ori09));
  INV        o0774(.A(ori_ori_n120_), .Y(ori_ori_n803_));
  NA2        o0775(.A(f), .B(e), .Y(ori_ori_n804_));
  NO2        o0776(.A(ori_ori_n227_), .B(ori_ori_n111_), .Y(ori_ori_n805_));
  NA2        o0777(.A(ori_ori_n805_), .B(g), .Y(ori_ori_n806_));
  NA3        o0778(.A(ori_ori_n309_), .B(ori_ori_n462_), .C(ori_ori_n264_), .Y(ori_ori_n807_));
  AOI210     o0779(.A0(ori_ori_n807_), .A1(g), .B0(ori_ori_n459_), .Y(ori_ori_n808_));
  AOI210     o0780(.A0(ori_ori_n808_), .A1(ori_ori_n806_), .B0(ori_ori_n804_), .Y(ori_ori_n809_));
  NA2        o0781(.A(ori_ori_n431_), .B(e), .Y(ori_ori_n810_));
  NO2        o0782(.A(ori_ori_n810_), .B(ori_ori_n503_), .Y(ori_ori_n811_));
  AOI210     o0783(.A0(ori_ori_n809_), .A1(ori_ori_n803_), .B0(ori_ori_n811_), .Y(ori_ori_n812_));
  NO2        o0784(.A(ori_ori_n205_), .B(ori_ori_n215_), .Y(ori_ori_n813_));
  NA3        o0785(.A(m), .B(l), .C(i), .Y(ori_ori_n814_));
  OAI220     o0786(.A0(ori_ori_n576_), .A1(ori_ori_n814_), .B0(ori_ori_n347_), .B1(ori_ori_n517_), .Y(ori_ori_n815_));
  NA4        o0787(.A(ori_ori_n85_), .B(ori_ori_n84_), .C(g), .D(f), .Y(ori_ori_n816_));
  NAi21      o0788(.An(ori_ori_n815_), .B(ori_ori_n816_), .Y(ori_ori_n817_));
  OR2        o0789(.A(ori_ori_n817_), .B(ori_ori_n813_), .Y(ori_ori_n818_));
  NA3        o0790(.A(ori_ori_n781_), .B(ori_ori_n557_), .C(ori_ori_n511_), .Y(ori_ori_n819_));
  OA210      o0791(.A0(ori_ori_n819_), .A1(ori_ori_n818_), .B0(ori_ori_n784_), .Y(ori_ori_n820_));
  INV        o0792(.A(ori_ori_n336_), .Y(ori_ori_n821_));
  NO2        o0793(.A(ori_ori_n125_), .B(ori_ori_n123_), .Y(ori_ori_n822_));
  INV        o0794(.A(ori_ori_n337_), .Y(ori_ori_n823_));
  AOI210     o0795(.A0(ori_ori_n823_), .A1(ori_ori_n822_), .B0(ori_ori_n585_), .Y(ori_ori_n824_));
  NA2        o0796(.A(ori_ori_n769_), .B(ori_ori_n329_), .Y(ori_ori_n825_));
  NA2        o0797(.A(ori_ori_n339_), .B(ori_ori_n340_), .Y(ori_ori_n826_));
  OAI210     o0798(.A0(ori_ori_n205_), .A1(ori_ori_n215_), .B0(ori_ori_n826_), .Y(ori_ori_n827_));
  AOI220     o0799(.A0(ori_ori_n827_), .A1(ori_ori_n825_), .B0(ori_ori_n824_), .B1(ori_ori_n821_), .Y(ori_ori_n828_));
  NA2        o0800(.A(ori_ori_n681_), .B(ori_ori_n134_), .Y(ori_ori_n829_));
  NA3        o0801(.A(ori_ori_n829_), .B(ori_ori_n190_), .C(ori_ori_n31_), .Y(ori_ori_n830_));
  NA3        o0802(.A(ori_ori_n830_), .B(ori_ori_n828_), .C(ori_ori_n610_), .Y(ori_ori_n831_));
  NO2        o0803(.A(ori_ori_n572_), .B(ori_ori_n488_), .Y(ori_ori_n832_));
  NOi21      o0804(.An(f), .B(d), .Y(ori_ori_n833_));
  NA2        o0805(.A(ori_ori_n833_), .B(m), .Y(ori_ori_n834_));
  NO2        o0806(.A(ori_ori_n834_), .B(ori_ori_n52_), .Y(ori_ori_n835_));
  NOi32      o0807(.An(g), .Bn(f), .C(d), .Y(ori_ori_n836_));
  NA4        o0808(.A(ori_ori_n836_), .B(ori_ori_n590_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n837_));
  NA2        o0809(.A(ori_ori_n835_), .B(ori_ori_n535_), .Y(ori_ori_n838_));
  AN2        o0810(.A(f), .B(d), .Y(ori_ori_n839_));
  NA3        o0811(.A(ori_ori_n467_), .B(ori_ori_n839_), .C(ori_ori_n81_), .Y(ori_ori_n840_));
  NO3        o0812(.A(ori_ori_n840_), .B(ori_ori_n73_), .C(ori_ori_n216_), .Y(ori_ori_n841_));
  NAi21      o0813(.An(ori_ori_n481_), .B(ori_ori_n838_), .Y(ori_ori_n842_));
  NO2        o0814(.A(ori_ori_n641_), .B(ori_ori_n326_), .Y(ori_ori_n843_));
  INV        o0815(.A(ori_ori_n236_), .Y(ori_ori_n844_));
  NA2        o0816(.A(ori_ori_n588_), .B(ori_ori_n81_), .Y(ori_ori_n845_));
  NO2        o0817(.A(ori_ori_n826_), .B(ori_ori_n845_), .Y(ori_ori_n846_));
  NA3        o0818(.A(ori_ori_n160_), .B(ori_ori_n107_), .C(ori_ori_n106_), .Y(ori_ori_n847_));
  OAI220     o0819(.A0(ori_ori_n840_), .A1(ori_ori_n422_), .B0(ori_ori_n336_), .B1(ori_ori_n847_), .Y(ori_ori_n848_));
  NO3        o0820(.A(ori_ori_n848_), .B(ori_ori_n846_), .C(ori_ori_n304_), .Y(ori_ori_n849_));
  NA2        o0821(.A(c), .B(ori_ori_n115_), .Y(ori_ori_n850_));
  NO2        o0822(.A(ori_ori_n850_), .B(ori_ori_n402_), .Y(ori_ori_n851_));
  NA3        o0823(.A(ori_ori_n851_), .B(ori_ori_n501_), .C(f), .Y(ori_ori_n852_));
  OR2        o0824(.A(ori_ori_n646_), .B(ori_ori_n531_), .Y(ori_ori_n853_));
  INV        o0825(.A(ori_ori_n853_), .Y(ori_ori_n854_));
  NA2        o0826(.A(ori_ori_n783_), .B(ori_ori_n110_), .Y(ori_ori_n855_));
  NA2        o0827(.A(ori_ori_n855_), .B(ori_ori_n854_), .Y(ori_ori_n856_));
  NA4        o0828(.A(ori_ori_n856_), .B(ori_ori_n852_), .C(ori_ori_n849_), .D(ori_ori_n844_), .Y(ori_ori_n857_));
  NO4        o0829(.A(ori_ori_n857_), .B(ori_ori_n842_), .C(ori_ori_n831_), .D(ori_ori_n820_), .Y(ori_ori_n858_));
  NA2        o0830(.A(ori_ori_n111_), .B(j), .Y(ori_ori_n859_));
  NO2        o0831(.A(ori_ori_n329_), .B(ori_ori_n816_), .Y(ori_ori_n860_));
  NO2        o0832(.A(ori_ori_n134_), .B(ori_ori_n130_), .Y(ori_ori_n861_));
  NO2        o0833(.A(ori_ori_n232_), .B(ori_ori_n226_), .Y(ori_ori_n862_));
  AOI220     o0834(.A0(ori_ori_n862_), .A1(ori_ori_n229_), .B0(ori_ori_n302_), .B1(ori_ori_n861_), .Y(ori_ori_n863_));
  NO2        o0835(.A(ori_ori_n422_), .B(ori_ori_n804_), .Y(ori_ori_n864_));
  NA2        o0836(.A(ori_ori_n864_), .B(ori_ori_n552_), .Y(ori_ori_n865_));
  NA2        o0837(.A(ori_ori_n865_), .B(ori_ori_n863_), .Y(ori_ori_n866_));
  NA2        o0838(.A(e), .B(d), .Y(ori_ori_n867_));
  OAI220     o0839(.A0(ori_ori_n867_), .A1(c), .B0(ori_ori_n323_), .B1(d), .Y(ori_ori_n868_));
  NA3        o0840(.A(ori_ori_n868_), .B(ori_ori_n442_), .C(ori_ori_n499_), .Y(ori_ori_n869_));
  AOI210     o0841(.A0(ori_ori_n506_), .A1(ori_ori_n180_), .B0(ori_ori_n232_), .Y(ori_ori_n870_));
  AOI210     o0842(.A0(ori_ori_n609_), .A1(ori_ori_n342_), .B0(ori_ori_n870_), .Y(ori_ori_n871_));
  NA2        o0843(.A(ori_ori_n285_), .B(ori_ori_n165_), .Y(ori_ori_n872_));
  NA2        o0844(.A(ori_ori_n841_), .B(ori_ori_n872_), .Y(ori_ori_n873_));
  NA3        o0845(.A(ori_ori_n873_), .B(ori_ori_n871_), .C(ori_ori_n869_), .Y(ori_ori_n874_));
  NO3        o0846(.A(ori_ori_n874_), .B(ori_ori_n866_), .C(ori_ori_n860_), .Y(ori_ori_n875_));
  OR2        o0847(.A(ori_ori_n683_), .B(ori_ori_n219_), .Y(ori_ori_n876_));
  NO2        o0848(.A(ori_ori_n608_), .B(ori_ori_n61_), .Y(ori_ori_n877_));
  AOI220     o0849(.A0(ori_ori_n877_), .A1(ori_ori_n843_), .B0(ori_ori_n600_), .B1(ori_ori_n607_), .Y(ori_ori_n878_));
  OAI210     o0850(.A0(ori_ori_n810_), .A1(ori_ori_n170_), .B0(ori_ori_n878_), .Y(ori_ori_n879_));
  OAI210     o0851(.A0(ori_ori_n805_), .A1(ori_ori_n872_), .B0(ori_ori_n836_), .Y(ori_ori_n880_));
  NO2        o0852(.A(ori_ori_n880_), .B(ori_ori_n591_), .Y(ori_ori_n881_));
  AOI210     o0853(.A0(ori_ori_n117_), .A1(ori_ori_n116_), .B0(ori_ori_n263_), .Y(ori_ori_n882_));
  NO2        o0854(.A(ori_ori_n882_), .B(ori_ori_n837_), .Y(ori_ori_n883_));
  AO210      o0855(.A0(ori_ori_n825_), .A1(ori_ori_n815_), .B0(ori_ori_n883_), .Y(ori_ori_n884_));
  NOi31      o0856(.An(ori_ori_n535_), .B(ori_ori_n834_), .C(ori_ori_n293_), .Y(ori_ori_n885_));
  NO4        o0857(.A(ori_ori_n885_), .B(ori_ori_n884_), .C(ori_ori_n881_), .D(ori_ori_n879_), .Y(ori_ori_n886_));
  AO220      o0858(.A0(ori_ori_n442_), .A1(ori_ori_n725_), .B0(ori_ori_n175_), .B1(f), .Y(ori_ori_n887_));
  OAI210     o0859(.A0(ori_ori_n887_), .A1(ori_ori_n445_), .B0(ori_ori_n868_), .Y(ori_ori_n888_));
  NO2        o0860(.A(ori_ori_n429_), .B(ori_ori_n70_), .Y(ori_ori_n889_));
  OAI210     o0861(.A0(ori_ori_n819_), .A1(ori_ori_n889_), .B0(ori_ori_n687_), .Y(ori_ori_n890_));
  AN4        o0862(.A(ori_ori_n890_), .B(ori_ori_n888_), .C(ori_ori_n886_), .D(ori_ori_n876_), .Y(ori_ori_n891_));
  NA4        o0863(.A(ori_ori_n891_), .B(ori_ori_n875_), .C(ori_ori_n858_), .D(ori_ori_n812_), .Y(ori12));
  NO2        o0864(.A(ori_ori_n440_), .B(c), .Y(ori_ori_n893_));
  NO4        o0865(.A(ori_ori_n430_), .B(ori_ori_n255_), .C(ori_ori_n569_), .D(ori_ori_n216_), .Y(ori_ori_n894_));
  NA2        o0866(.A(ori_ori_n894_), .B(ori_ori_n893_), .Y(ori_ori_n895_));
  NA2        o0867(.A(ori_ori_n535_), .B(ori_ori_n889_), .Y(ori_ori_n896_));
  NO2        o0868(.A(ori_ori_n440_), .B(ori_ori_n115_), .Y(ori_ori_n897_));
  NO2        o0869(.A(ori_ori_n822_), .B(ori_ori_n347_), .Y(ori_ori_n898_));
  NO2        o0870(.A(ori_ori_n646_), .B(ori_ori_n372_), .Y(ori_ori_n899_));
  AOI220     o0871(.A0(ori_ori_n899_), .A1(ori_ori_n533_), .B0(ori_ori_n898_), .B1(ori_ori_n897_), .Y(ori_ori_n900_));
  NA3        o0872(.A(ori_ori_n900_), .B(ori_ori_n896_), .C(ori_ori_n895_), .Y(ori_ori_n901_));
  AOI210     o0873(.A0(ori_ori_n235_), .A1(ori_ori_n335_), .B0(ori_ori_n202_), .Y(ori_ori_n902_));
  OR2        o0874(.A(ori_ori_n902_), .B(ori_ori_n894_), .Y(ori_ori_n903_));
  AOI210     o0875(.A0(ori_ori_n332_), .A1(ori_ori_n383_), .B0(ori_ori_n216_), .Y(ori_ori_n904_));
  OAI210     o0876(.A0(ori_ori_n904_), .A1(ori_ori_n903_), .B0(ori_ori_n397_), .Y(ori_ori_n905_));
  NO2        o0877(.A(ori_ori_n627_), .B(ori_ori_n266_), .Y(ori_ori_n906_));
  NO2        o0878(.A(ori_ori_n576_), .B(ori_ori_n814_), .Y(ori_ori_n907_));
  AOI220     o0879(.A0(ori_ori_n907_), .A1(ori_ori_n555_), .B0(ori_ori_n794_), .B1(ori_ori_n906_), .Y(ori_ori_n908_));
  NO2        o0880(.A(ori_ori_n151_), .B(ori_ori_n239_), .Y(ori_ori_n909_));
  NA2        o0881(.A(ori_ori_n908_), .B(ori_ori_n905_), .Y(ori_ori_n910_));
  OR2        o0882(.A(ori_ori_n324_), .B(ori_ori_n897_), .Y(ori_ori_n911_));
  NA2        o0883(.A(ori_ori_n911_), .B(ori_ori_n348_), .Y(ori_ori_n912_));
  NA4        o0884(.A(ori_ori_n431_), .B(ori_ori_n428_), .C(ori_ori_n181_), .D(g), .Y(ori_ori_n913_));
  NA2        o0885(.A(ori_ori_n913_), .B(ori_ori_n912_), .Y(ori_ori_n914_));
  NO3        o0886(.A(ori_ori_n651_), .B(ori_ori_n89_), .C(ori_ori_n45_), .Y(ori_ori_n915_));
  NO4        o0887(.A(ori_ori_n915_), .B(ori_ori_n914_), .C(ori_ori_n910_), .D(ori_ori_n901_), .Y(ori_ori_n916_));
  NA2        o0888(.A(ori_ori_n545_), .B(ori_ori_n144_), .Y(ori_ori_n917_));
  NOi21      o0889(.An(ori_ori_n34_), .B(ori_ori_n641_), .Y(ori_ori_n918_));
  NA2        o0890(.A(ori_ori_n918_), .B(ori_ori_n917_), .Y(ori_ori_n919_));
  OAI210     o0891(.A0(ori_ori_n253_), .A1(ori_ori_n45_), .B0(ori_ori_n919_), .Y(ori_ori_n920_));
  INV        o0892(.A(ori_ori_n320_), .Y(ori_ori_n921_));
  NO2        o0893(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n922_));
  NO2        o0894(.A(ori_ori_n495_), .B(ori_ori_n297_), .Y(ori_ori_n923_));
  INV        o0895(.A(ori_ori_n923_), .Y(ori_ori_n924_));
  NO2        o0896(.A(ori_ori_n924_), .B(ori_ori_n144_), .Y(ori_ori_n925_));
  INV        o0897(.A(ori_ori_n359_), .Y(ori_ori_n926_));
  NO4        o0898(.A(ori_ori_n926_), .B(ori_ori_n925_), .C(ori_ori_n921_), .D(ori_ori_n920_), .Y(ori_ori_n927_));
  NA2        o0899(.A(ori_ori_n342_), .B(g), .Y(ori_ori_n928_));
  NA2        o0900(.A(ori_ori_n163_), .B(i), .Y(ori_ori_n929_));
  NA2        o0901(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n930_));
  OAI220     o0902(.A0(ori_ori_n930_), .A1(ori_ori_n201_), .B0(ori_ori_n929_), .B1(ori_ori_n89_), .Y(ori_ori_n931_));
  INV        o0903(.A(ori_ori_n931_), .Y(ori_ori_n932_));
  NA2        o0904(.A(ori_ori_n545_), .B(ori_ori_n375_), .Y(ori_ori_n933_));
  AOI210     o0905(.A0(ori_ori_n933_), .A1(n), .B0(ori_ori_n544_), .Y(ori_ori_n934_));
  OAI220     o0906(.A0(ori_ori_n934_), .A1(ori_ori_n928_), .B0(ori_ori_n932_), .B1(ori_ori_n329_), .Y(ori_ori_n935_));
  NO2        o0907(.A(ori_ori_n646_), .B(ori_ori_n488_), .Y(ori_ori_n936_));
  NA3        o0908(.A(ori_ori_n339_), .B(ori_ori_n613_), .C(i), .Y(ori_ori_n937_));
  OAI210     o0909(.A0(ori_ori_n429_), .A1(ori_ori_n309_), .B0(ori_ori_n937_), .Y(ori_ori_n938_));
  OAI220     o0910(.A0(ori_ori_n938_), .A1(ori_ori_n936_), .B0(ori_ori_n665_), .B1(ori_ori_n737_), .Y(ori_ori_n939_));
  NA2        o0911(.A(ori_ori_n594_), .B(ori_ori_n112_), .Y(ori_ori_n940_));
  OR3        o0912(.A(ori_ori_n309_), .B(ori_ori_n427_), .C(f), .Y(ori_ori_n941_));
  NA3        o0913(.A(ori_ori_n613_), .B(ori_ori_n79_), .C(i), .Y(ori_ori_n942_));
  OA220      o0914(.A0(ori_ori_n942_), .A1(ori_ori_n940_), .B0(ori_ori_n941_), .B1(ori_ori_n575_), .Y(ori_ori_n943_));
  NA3        o0915(.A(ori_ori_n325_), .B(ori_ori_n117_), .C(g), .Y(ori_ori_n944_));
  AOI210     o0916(.A0(ori_ori_n662_), .A1(ori_ori_n944_), .B0(m), .Y(ori_ori_n945_));
  OAI210     o0917(.A0(ori_ori_n945_), .A1(ori_ori_n898_), .B0(ori_ori_n324_), .Y(ori_ori_n946_));
  NA2        o0918(.A(ori_ori_n676_), .B(ori_ori_n845_), .Y(ori_ori_n947_));
  INV        o0919(.A(ori_ori_n816_), .Y(ori_ori_n948_));
  INV        o0920(.A(ori_ori_n942_), .Y(ori_ori_n949_));
  AOI220     o0921(.A0(ori_ori_n949_), .A1(ori_ori_n261_), .B0(ori_ori_n948_), .B1(ori_ori_n947_), .Y(ori_ori_n950_));
  NA4        o0922(.A(ori_ori_n950_), .B(ori_ori_n946_), .C(ori_ori_n943_), .D(ori_ori_n939_), .Y(ori_ori_n951_));
  NO2        o0923(.A(ori_ori_n372_), .B(ori_ori_n88_), .Y(ori_ori_n952_));
  OAI210     o0924(.A0(ori_ori_n952_), .A1(ori_ori_n906_), .B0(ori_ori_n240_), .Y(ori_ori_n953_));
  NA2        o0925(.A(ori_ori_n650_), .B(ori_ori_n85_), .Y(ori_ori_n954_));
  NO2        o0926(.A(ori_ori_n448_), .B(ori_ori_n216_), .Y(ori_ori_n955_));
  AOI220     o0927(.A0(ori_ori_n955_), .A1(ori_ori_n376_), .B0(ori_ori_n911_), .B1(ori_ori_n220_), .Y(ori_ori_n956_));
  AOI220     o0928(.A0(ori_ori_n899_), .A1(ori_ori_n909_), .B0(ori_ori_n574_), .B1(ori_ori_n87_), .Y(ori_ori_n957_));
  NA4        o0929(.A(ori_ori_n957_), .B(ori_ori_n956_), .C(ori_ori_n954_), .D(ori_ori_n953_), .Y(ori_ori_n958_));
  NA2        o0930(.A(ori_ori_n948_), .B(ori_ori_n533_), .Y(ori_ori_n959_));
  AOI210     o0931(.A0(ori_ori_n414_), .A1(ori_ori_n406_), .B0(ori_ori_n796_), .Y(ori_ori_n960_));
  OAI210     o0932(.A0(ori_ori_n362_), .A1(ori_ori_n361_), .B0(ori_ori_n108_), .Y(ori_ori_n961_));
  AOI210     o0933(.A0(ori_ori_n961_), .A1(ori_ori_n525_), .B0(ori_ori_n960_), .Y(ori_ori_n962_));
  NA2        o0934(.A(ori_ori_n945_), .B(ori_ori_n897_), .Y(ori_ori_n963_));
  NO3        o0935(.A(ori_ori_n859_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n964_));
  NA2        o0936(.A(ori_ori_n964_), .B(ori_ori_n612_), .Y(ori_ori_n965_));
  NA4        o0937(.A(ori_ori_n965_), .B(ori_ori_n963_), .C(ori_ori_n962_), .D(ori_ori_n959_), .Y(ori_ori_n966_));
  NO4        o0938(.A(ori_ori_n966_), .B(ori_ori_n958_), .C(ori_ori_n951_), .D(ori_ori_n935_), .Y(ori_ori_n967_));
  NAi31      o0939(.An(ori_ori_n140_), .B(ori_ori_n415_), .C(n), .Y(ori_ori_n968_));
  NO2        o0940(.A(ori_ori_n123_), .B(ori_ori_n337_), .Y(ori_ori_n969_));
  NO2        o0941(.A(ori_ori_n969_), .B(ori_ori_n968_), .Y(ori_ori_n970_));
  NO3        o0942(.A(ori_ori_n275_), .B(ori_ori_n140_), .C(ori_ori_n402_), .Y(ori_ori_n971_));
  AOI210     o0943(.A0(ori_ori_n971_), .A1(ori_ori_n489_), .B0(ori_ori_n970_), .Y(ori_ori_n972_));
  NA2        o0944(.A(ori_ori_n482_), .B(i), .Y(ori_ori_n973_));
  NA2        o0945(.A(ori_ori_n973_), .B(ori_ori_n972_), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n232_), .B(ori_ori_n171_), .Y(ori_ori_n975_));
  NO3        o0947(.A(ori_ori_n306_), .B(ori_ori_n431_), .C(ori_ori_n175_), .Y(ori_ori_n976_));
  NOi31      o0948(.An(ori_ori_n975_), .B(ori_ori_n976_), .C(ori_ori_n216_), .Y(ori_ori_n977_));
  NAi21      o0949(.An(ori_ori_n545_), .B(ori_ori_n955_), .Y(ori_ori_n978_));
  NA2        o0950(.A(ori_ori_n473_), .B(g), .Y(ori_ori_n979_));
  NA2        o0951(.A(ori_ori_n979_), .B(ori_ori_n978_), .Y(ori_ori_n980_));
  OAI220     o0952(.A0(ori_ori_n968_), .A1(ori_ori_n235_), .B0(ori_ori_n937_), .B1(ori_ori_n589_), .Y(ori_ori_n981_));
  NO2        o0953(.A(ori_ori_n647_), .B(ori_ori_n372_), .Y(ori_ori_n982_));
  NA2        o0954(.A(ori_ori_n902_), .B(ori_ori_n893_), .Y(ori_ori_n983_));
  NO3        o0955(.A(ori_ori_n534_), .B(ori_ori_n149_), .C(ori_ori_n215_), .Y(ori_ori_n984_));
  OAI210     o0956(.A0(ori_ori_n984_), .A1(ori_ori_n515_), .B0(ori_ori_n373_), .Y(ori_ori_n985_));
  OAI220     o0957(.A0(ori_ori_n899_), .A1(ori_ori_n907_), .B0(ori_ori_n535_), .B1(ori_ori_n421_), .Y(ori_ori_n986_));
  NA4        o0958(.A(ori_ori_n986_), .B(ori_ori_n985_), .C(ori_ori_n983_), .D(ori_ori_n606_), .Y(ori_ori_n987_));
  OAI210     o0959(.A0(ori_ori_n902_), .A1(ori_ori_n894_), .B0(ori_ori_n975_), .Y(ori_ori_n988_));
  NA3        o0960(.A(ori_ori_n933_), .B(ori_ori_n478_), .C(ori_ori_n46_), .Y(ori_ori_n989_));
  INV        o0961(.A(ori_ori_n328_), .Y(ori_ori_n990_));
  NA4        o0962(.A(ori_ori_n990_), .B(ori_ori_n989_), .C(ori_ori_n988_), .D(ori_ori_n276_), .Y(ori_ori_n991_));
  OR4        o0963(.A(ori_ori_n991_), .B(ori_ori_n987_), .C(ori_ori_n982_), .D(ori_ori_n981_), .Y(ori_ori_n992_));
  NO4        o0964(.A(ori_ori_n992_), .B(ori_ori_n980_), .C(ori_ori_n977_), .D(ori_ori_n974_), .Y(ori_ori_n993_));
  NA4        o0965(.A(ori_ori_n993_), .B(ori_ori_n967_), .C(ori_ori_n927_), .D(ori_ori_n916_), .Y(ori13));
  NAi32      o0966(.An(d), .Bn(c), .C(e), .Y(ori_ori_n995_));
  NA2        o0967(.A(ori_ori_n139_), .B(ori_ori_n45_), .Y(ori_ori_n996_));
  NO4        o0968(.A(ori_ori_n996_), .B(ori_ori_n995_), .C(ori_ori_n576_), .D(ori_ori_n305_), .Y(ori_ori_n997_));
  NA2        o0969(.A(ori_ori_n405_), .B(ori_ori_n215_), .Y(ori_ori_n998_));
  AN2        o0970(.A(d), .B(c), .Y(ori_ori_n999_));
  NA2        o0971(.A(ori_ori_n999_), .B(ori_ori_n115_), .Y(ori_ori_n1000_));
  NA2        o0972(.A(ori_ori_n486_), .B(c), .Y(ori_ori_n1001_));
  NO4        o0973(.A(ori_ori_n996_), .B(ori_ori_n572_), .C(ori_ori_n1001_), .D(ori_ori_n305_), .Y(ori_ori_n1002_));
  OR2        o0974(.A(ori_ori_n1002_), .B(ori_ori_n997_), .Y(ori_ori_n1003_));
  NAi32      o0975(.An(f), .Bn(e), .C(c), .Y(ori_ori_n1004_));
  NO2        o0976(.A(ori_ori_n1001_), .B(ori_ori_n305_), .Y(ori_ori_n1005_));
  NO2        o0977(.A(j), .B(ori_ori_n45_), .Y(ori_ori_n1006_));
  NA2        o0978(.A(ori_ori_n615_), .B(ori_ori_n1006_), .Y(ori_ori_n1007_));
  NOi21      o0979(.An(ori_ori_n1005_), .B(ori_ori_n1007_), .Y(ori_ori_n1008_));
  NOi41      o0980(.An(n), .B(m), .C(i), .D(h), .Y(ori_ori_n1009_));
  NA3        o0981(.A(k), .B(j), .C(i), .Y(ori_ori_n1010_));
  NA3        o0982(.A(ori_ori_n456_), .B(ori_ori_n331_), .C(ori_ori_n56_), .Y(ori_ori_n1011_));
  NO2        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1007_), .Y(ori_ori_n1012_));
  NO3        o0984(.A(ori_ori_n1011_), .B(ori_ori_n572_), .C(ori_ori_n438_), .Y(ori_ori_n1013_));
  OR2        o0985(.A(ori_ori_n1013_), .B(ori_ori_n1012_), .Y(ori_ori_n1014_));
  OR3        o0986(.A(ori_ori_n1014_), .B(ori_ori_n1008_), .C(ori_ori_n1003_), .Y(ori02));
  OR3        o0987(.A(n), .B(m), .C(i), .Y(ori_ori_n1016_));
  NOi31      o0988(.An(e), .B(d), .C(c), .Y(ori_ori_n1017_));
  INV        o0989(.A(ori_ori_n997_), .Y(ori_ori_n1018_));
  AN3        o0990(.A(g), .B(f), .C(c), .Y(ori_ori_n1019_));
  NO3        o0991(.A(ori_ori_n1011_), .B(ori_ori_n996_), .C(ori_ori_n572_), .Y(ori_ori_n1020_));
  INV        o0992(.A(ori_ori_n1020_), .Y(ori_ori_n1021_));
  NA3        o0993(.A(l), .B(k), .C(j), .Y(ori_ori_n1022_));
  NA2        o0994(.A(i), .B(h), .Y(ori_ori_n1023_));
  NO3        o0995(.A(ori_ori_n1023_), .B(ori_ori_n1022_), .C(ori_ori_n130_), .Y(ori_ori_n1024_));
  NO3        o0996(.A(ori_ori_n141_), .B(ori_ori_n283_), .C(ori_ori_n216_), .Y(ori_ori_n1025_));
  AOI210     o0997(.A0(ori_ori_n1025_), .A1(ori_ori_n1024_), .B0(ori_ori_n1008_), .Y(ori_ori_n1026_));
  NA3        o0998(.A(c), .B(b), .C(a), .Y(ori_ori_n1027_));
  INV        o0999(.A(ori_ori_n1012_), .Y(ori_ori_n1028_));
  AN3        o1000(.A(ori_ori_n1028_), .B(ori_ori_n1026_), .C(ori_ori_n1021_), .Y(ori_ori_n1029_));
  NA2        o1001(.A(ori_ori_n1029_), .B(ori_ori_n1018_), .Y(ori03));
  NA4        o1002(.A(ori_ori_n85_), .B(ori_ori_n84_), .C(g), .D(ori_ori_n215_), .Y(ori_ori_n1031_));
  INV        o1003(.A(ori_ori_n1031_), .Y(ori_ori_n1032_));
  NO2        o1004(.A(ori_ori_n1032_), .B(ori_ori_n961_), .Y(ori_ori_n1033_));
  NOi41      o1005(.An(ori_ori_n781_), .B(ori_ori_n827_), .C(ori_ori_n817_), .D(ori_ori_n698_), .Y(ori_ori_n1034_));
  OAI220     o1006(.A0(ori_ori_n1034_), .A1(ori_ori_n676_), .B0(ori_ori_n1033_), .B1(ori_ori_n573_), .Y(ori_ori_n1035_));
  NOi31      o1007(.An(i), .B(k), .C(j), .Y(ori_ori_n1036_));
  NA4        o1008(.A(ori_ori_n1036_), .B(ori_ori_n1017_), .C(ori_ori_n339_), .D(ori_ori_n331_), .Y(ori_ori_n1037_));
  OAI210     o1009(.A0(ori_ori_n796_), .A1(ori_ori_n416_), .B0(ori_ori_n1037_), .Y(ori_ori_n1038_));
  NOi31      o1010(.An(m), .B(n), .C(f), .Y(ori_ori_n1039_));
  NA2        o1011(.A(ori_ori_n1039_), .B(ori_ori_n51_), .Y(ori_ori_n1040_));
  AN2        o1012(.A(e), .B(c), .Y(ori_ori_n1041_));
  NA2        o1013(.A(ori_ori_n1041_), .B(a), .Y(ori_ori_n1042_));
  OAI220     o1014(.A0(ori_ori_n1042_), .A1(ori_ori_n1040_), .B0(ori_ori_n853_), .B1(ori_ori_n420_), .Y(ori_ori_n1043_));
  NA2        o1015(.A(ori_ori_n499_), .B(l), .Y(ori_ori_n1044_));
  NO3        o1016(.A(ori_ori_n1043_), .B(ori_ori_n1038_), .C(ori_ori_n960_), .Y(ori_ori_n1045_));
  NO2        o1017(.A(ori_ori_n283_), .B(a), .Y(ori_ori_n1046_));
  INV        o1018(.A(ori_ori_n997_), .Y(ori_ori_n1047_));
  NO2        o1019(.A(ori_ori_n84_), .B(g), .Y(ori_ori_n1048_));
  NA2        o1020(.A(ori_ori_n1047_), .B(ori_ori_n1045_), .Y(ori_ori_n1049_));
  NO4        o1021(.A(ori_ori_n1049_), .B(ori_ori_n1035_), .C(ori_ori_n797_), .D(ori_ori_n554_), .Y(ori_ori_n1050_));
  NA2        o1022(.A(c), .B(b), .Y(ori_ori_n1051_));
  NO2        o1023(.A(ori_ori_n686_), .B(ori_ori_n1051_), .Y(ori_ori_n1052_));
  OAI210     o1024(.A0(ori_ori_n834_), .A1(ori_ori_n808_), .B0(ori_ori_n409_), .Y(ori_ori_n1053_));
  OAI210     o1025(.A0(ori_ori_n1053_), .A1(ori_ori_n835_), .B0(ori_ori_n1052_), .Y(ori_ori_n1054_));
  NAi21      o1026(.An(ori_ori_n417_), .B(ori_ori_n1052_), .Y(ori_ori_n1055_));
  NA3        o1027(.A(ori_ori_n421_), .B(ori_ori_n550_), .C(f), .Y(ori_ori_n1056_));
  OAI210     o1028(.A0(ori_ori_n539_), .A1(ori_ori_n39_), .B0(ori_ori_n1046_), .Y(ori_ori_n1057_));
  NA3        o1029(.A(ori_ori_n1057_), .B(ori_ori_n1056_), .C(ori_ori_n1055_), .Y(ori_ori_n1058_));
  INV        o1030(.A(ori_ori_n264_), .Y(ori_ori_n1059_));
  OAI210     o1031(.A0(ori_ori_n1059_), .A1(ori_ori_n287_), .B0(g), .Y(ori_ori_n1060_));
  NAi21      o1032(.An(f), .B(d), .Y(ori_ori_n1061_));
  NO2        o1033(.A(ori_ori_n1061_), .B(ori_ori_n1027_), .Y(ori_ori_n1062_));
  INV        o1034(.A(ori_ori_n1062_), .Y(ori_ori_n1063_));
  NO2        o1035(.A(ori_ori_n1060_), .B(ori_ori_n1063_), .Y(ori_ori_n1064_));
  AOI210     o1036(.A0(ori_ori_n1064_), .A1(ori_ori_n112_), .B0(ori_ori_n1058_), .Y(ori_ori_n1065_));
  NA2        o1037(.A(ori_ori_n459_), .B(ori_ori_n458_), .Y(ori_ori_n1066_));
  NO2        o1038(.A(ori_ori_n182_), .B(ori_ori_n239_), .Y(ori_ori_n1067_));
  NA2        o1039(.A(ori_ori_n1067_), .B(m), .Y(ori_ori_n1068_));
  NA3        o1040(.A(ori_ori_n882_), .B(ori_ori_n1044_), .C(ori_ori_n462_), .Y(ori_ori_n1069_));
  OAI210     o1041(.A0(ori_ori_n1069_), .A1(ori_ori_n310_), .B0(ori_ori_n460_), .Y(ori_ori_n1070_));
  AOI210     o1042(.A0(ori_ori_n1070_), .A1(ori_ori_n1066_), .B0(ori_ori_n1068_), .Y(ori_ori_n1071_));
  NA2        o1043(.A(ori_ori_n552_), .B(ori_ori_n404_), .Y(ori_ori_n1072_));
  NA2        o1044(.A(ori_ori_n159_), .B(ori_ori_n33_), .Y(ori_ori_n1073_));
  NO2        o1045(.A(ori_ori_n1073_), .B(ori_ori_n216_), .Y(ori_ori_n1074_));
  OAI210     o1046(.A0(ori_ori_n1074_), .A1(ori_ori_n434_), .B0(ori_ori_n1062_), .Y(ori_ori_n1075_));
  NO2        o1047(.A(ori_ori_n366_), .B(ori_ori_n365_), .Y(ori_ori_n1076_));
  NA2        o1048(.A(ori_ori_n1067_), .B(ori_ori_n423_), .Y(ori_ori_n1077_));
  NAi41      o1049(.An(ori_ori_n1076_), .B(ori_ori_n1077_), .C(ori_ori_n1075_), .D(ori_ori_n1072_), .Y(ori_ori_n1078_));
  NO2        o1050(.A(ori_ori_n1078_), .B(ori_ori_n1071_), .Y(ori_ori_n1079_));
  NA4        o1051(.A(ori_ori_n1079_), .B(ori_ori_n1065_), .C(ori_ori_n1054_), .D(ori_ori_n1050_), .Y(ori00));
  AOI210     o1052(.A0(ori_ori_n864_), .A1(ori_ori_n909_), .B0(ori_ori_n1038_), .Y(ori_ori_n1081_));
  NO2        o1053(.A(ori_ori_n1020_), .B(ori_ori_n697_), .Y(ori_ori_n1082_));
  NA3        o1054(.A(ori_ori_n1082_), .B(ori_ori_n1081_), .C(ori_ori_n962_), .Y(ori_ori_n1083_));
  NA2        o1055(.A(ori_ori_n501_), .B(f), .Y(ori_ori_n1084_));
  OAI210     o1056(.A0(ori_ori_n969_), .A1(ori_ori_n40_), .B0(ori_ori_n634_), .Y(ori_ori_n1085_));
  NA3        o1057(.A(ori_ori_n1085_), .B(ori_ori_n260_), .C(n), .Y(ori_ori_n1086_));
  AOI210     o1058(.A0(ori_ori_n1086_), .A1(ori_ori_n1084_), .B0(ori_ori_n1000_), .Y(ori_ori_n1087_));
  NO3        o1059(.A(ori_ori_n1087_), .B(ori_ori_n1083_), .C(ori_ori_n1008_), .Y(ori_ori_n1088_));
  NA3        o1060(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1089_));
  NO2        o1061(.A(ori_ori_n1076_), .B(ori_ori_n885_), .Y(ori_ori_n1090_));
  NO4        o1062(.A(ori_ori_n479_), .B(ori_ori_n349_), .C(ori_ori_n1051_), .D(ori_ori_n59_), .Y(ori_ori_n1091_));
  NA3        o1063(.A(ori_ori_n377_), .B(ori_ori_n223_), .C(g), .Y(ori_ori_n1092_));
  OA220      o1064(.A0(ori_ori_n1092_), .A1(ori_ori_n1089_), .B0(ori_ori_n378_), .B1(ori_ori_n133_), .Y(ori_ori_n1093_));
  NO2        o1065(.A(h), .B(g), .Y(ori_ori_n1094_));
  OAI220     o1066(.A0(ori_ori_n517_), .A1(ori_ori_n585_), .B0(ori_ori_n89_), .B1(ori_ori_n88_), .Y(ori_ori_n1095_));
  NA2        o1067(.A(ori_ori_n1095_), .B(ori_ori_n525_), .Y(ori_ori_n1096_));
  AOI220     o1068(.A0(ori_ori_n317_), .A1(ori_ori_n249_), .B0(ori_ori_n177_), .B1(ori_ori_n148_), .Y(ori_ori_n1097_));
  NA3        o1069(.A(ori_ori_n1097_), .B(ori_ori_n1096_), .C(ori_ori_n1093_), .Y(ori_ori_n1098_));
  NO3        o1070(.A(ori_ori_n1098_), .B(ori_ori_n1091_), .C(ori_ori_n269_), .Y(ori_ori_n1099_));
  INV        o1071(.A(ori_ori_n322_), .Y(ori_ori_n1100_));
  AOI210     o1072(.A0(ori_ori_n249_), .A1(ori_ori_n342_), .B0(ori_ori_n566_), .Y(ori_ori_n1101_));
  NA3        o1073(.A(ori_ori_n1101_), .B(ori_ori_n1100_), .C(ori_ori_n154_), .Y(ori_ori_n1102_));
  NO2        o1074(.A(ori_ori_n241_), .B(ori_ori_n181_), .Y(ori_ori_n1103_));
  NA2        o1075(.A(ori_ori_n1103_), .B(ori_ori_n421_), .Y(ori_ori_n1104_));
  NA2        o1076(.A(ori_ori_n179_), .B(ori_ori_n111_), .Y(ori_ori_n1105_));
  NAi31      o1077(.An(ori_ori_n186_), .B(ori_ori_n832_), .C(ori_ori_n456_), .Y(ori_ori_n1106_));
  NA2        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1104_), .Y(ori_ori_n1107_));
  NO4        o1079(.A(ori_ori_n1002_), .B(ori_ori_n1107_), .C(ori_ori_n1102_), .D(ori_ori_n510_), .Y(ori_ori_n1108_));
  AN3        o1080(.A(ori_ori_n1108_), .B(ori_ori_n1099_), .C(ori_ori_n1090_), .Y(ori_ori_n1109_));
  NA2        o1081(.A(ori_ori_n525_), .B(ori_ori_n99_), .Y(ori_ori_n1110_));
  NA3        o1082(.A(ori_ori_n1039_), .B(ori_ori_n594_), .C(ori_ori_n455_), .Y(ori_ori_n1111_));
  NA4        o1083(.A(ori_ori_n1111_), .B(ori_ori_n553_), .C(ori_ori_n1110_), .D(ori_ori_n243_), .Y(ori_ori_n1112_));
  NA2        o1084(.A(ori_ori_n1032_), .B(ori_ori_n525_), .Y(ori_ori_n1113_));
  NA4        o1085(.A(ori_ori_n637_), .B(ori_ori_n207_), .C(ori_ori_n223_), .D(ori_ori_n163_), .Y(ori_ori_n1114_));
  NA2        o1086(.A(ori_ori_n1114_), .B(ori_ori_n1113_), .Y(ori_ori_n1115_));
  OAI210     o1087(.A0(ori_ori_n454_), .A1(ori_ori_n118_), .B0(ori_ori_n837_), .Y(ori_ori_n1116_));
  AOI220     o1088(.A0(ori_ori_n1116_), .A1(ori_ori_n1069_), .B0(ori_ori_n552_), .B1(ori_ori_n404_), .Y(ori_ori_n1117_));
  NA2        o1089(.A(n), .B(e), .Y(ori_ori_n1118_));
  NO2        o1090(.A(ori_ori_n1118_), .B(ori_ori_n146_), .Y(ori_ori_n1119_));
  OAI210     o1091(.A0(ori_ori_n350_), .A1(ori_ori_n311_), .B0(ori_ori_n436_), .Y(ori_ori_n1120_));
  NA2        o1092(.A(ori_ori_n1120_), .B(ori_ori_n1117_), .Y(ori_ori_n1121_));
  NA2        o1093(.A(ori_ori_n1119_), .B(ori_ori_n824_), .Y(ori_ori_n1122_));
  AOI220     o1094(.A0(ori_ori_n918_), .A1(ori_ori_n564_), .B0(ori_ori_n637_), .B1(ori_ori_n246_), .Y(ori_ori_n1123_));
  NO2        o1095(.A(ori_ori_n68_), .B(h), .Y(ori_ori_n1124_));
  NA3        o1096(.A(ori_ori_n1123_), .B(ori_ori_n1122_), .C(ori_ori_n838_), .Y(ori_ori_n1125_));
  NO4        o1097(.A(ori_ori_n1125_), .B(ori_ori_n1121_), .C(ori_ori_n1115_), .D(ori_ori_n1112_), .Y(ori_ori_n1126_));
  NA2        o1098(.A(ori_ori_n809_), .B(ori_ori_n736_), .Y(ori_ori_n1127_));
  NA4        o1099(.A(ori_ori_n1127_), .B(ori_ori_n1126_), .C(ori_ori_n1109_), .D(ori_ori_n1088_), .Y(ori01));
  AN2        o1100(.A(ori_ori_n985_), .B(ori_ori_n983_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(ori_ori_n470_), .B(ori_ori_n281_), .Y(ori_ori_n1130_));
  NA2        o1102(.A(ori_ori_n388_), .B(i), .Y(ori_ori_n1131_));
  NA3        o1103(.A(ori_ori_n1131_), .B(ori_ori_n1130_), .C(ori_ori_n1129_), .Y(ori_ori_n1132_));
  NA2        o1104(.A(ori_ori_n574_), .B(ori_ori_n87_), .Y(ori_ori_n1133_));
  NA2        o1105(.A(ori_ori_n545_), .B(ori_ori_n274_), .Y(ori_ori_n1134_));
  NA2        o1106(.A(ori_ori_n923_), .B(ori_ori_n1134_), .Y(ori_ori_n1135_));
  NA4        o1107(.A(ori_ori_n1135_), .B(ori_ori_n1133_), .C(ori_ori_n878_), .D(ori_ori_n330_), .Y(ori_ori_n1136_));
  NA2        o1108(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1137_));
  NA2        o1109(.A(ori_ori_n692_), .B(ori_ori_n94_), .Y(ori_ori_n1138_));
  NO2        o1110(.A(ori_ori_n1138_), .B(ori_ori_n1137_), .Y(ori_ori_n1139_));
  OAI210     o1111(.A0(ori_ori_n759_), .A1(ori_ori_n589_), .B0(ori_ori_n1114_), .Y(ori_ori_n1140_));
  AOI210     o1112(.A0(ori_ori_n1139_), .A1(ori_ori_n622_), .B0(ori_ori_n1140_), .Y(ori_ori_n1141_));
  INV        o1113(.A(ori_ori_n117_), .Y(ori_ori_n1142_));
  NAi31      o1114(.An(ori_ori_n162_), .B(ori_ori_n1141_), .C(ori_ori_n863_), .Y(ori_ori_n1143_));
  NO2        o1115(.A(ori_ori_n664_), .B(ori_ori_n504_), .Y(ori_ori_n1144_));
  NA4        o1116(.A(ori_ori_n692_), .B(ori_ori_n94_), .C(ori_ori_n45_), .D(ori_ori_n215_), .Y(ori_ori_n1145_));
  OA220      o1117(.A0(ori_ori_n1145_), .A1(ori_ori_n657_), .B0(ori_ori_n196_), .B1(ori_ori_n194_), .Y(ori_ori_n1146_));
  NA3        o1118(.A(ori_ori_n1146_), .B(ori_ori_n1144_), .C(ori_ori_n136_), .Y(ori_ori_n1147_));
  NO4        o1119(.A(ori_ori_n1147_), .B(ori_ori_n1143_), .C(ori_ori_n1136_), .D(ori_ori_n1132_), .Y(ori_ori_n1148_));
  NA2        o1120(.A(ori_ori_n299_), .B(ori_ori_n521_), .Y(ori_ori_n1149_));
  AOI210     o1121(.A0(ori_ori_n205_), .A1(ori_ori_n86_), .B0(ori_ori_n215_), .Y(ori_ori_n1150_));
  OAI210     o1122(.A0(ori_ori_n784_), .A1(ori_ori_n421_), .B0(ori_ori_n1150_), .Y(ori_ori_n1151_));
  AN3        o1123(.A(m), .B(l), .C(k), .Y(ori_ori_n1152_));
  OAI210     o1124(.A0(ori_ori_n351_), .A1(ori_ori_n34_), .B0(ori_ori_n1152_), .Y(ori_ori_n1153_));
  NA2        o1125(.A(ori_ori_n204_), .B(ori_ori_n34_), .Y(ori_ori_n1154_));
  AO210      o1126(.A0(ori_ori_n1154_), .A1(ori_ori_n1153_), .B0(ori_ori_n329_), .Y(ori_ori_n1155_));
  NA3        o1127(.A(ori_ori_n1155_), .B(ori_ori_n1151_), .C(ori_ori_n1149_), .Y(ori_ori_n1156_));
  AOI210     o1128(.A0(ori_ori_n583_), .A1(ori_ori_n117_), .B0(ori_ori_n587_), .Y(ori_ori_n1157_));
  OAI210     o1129(.A0(ori_ori_n1142_), .A1(ori_ori_n580_), .B0(ori_ori_n1157_), .Y(ori_ori_n1158_));
  NA2        o1130(.A(ori_ori_n280_), .B(ori_ori_n196_), .Y(ori_ori_n1159_));
  NA2        o1131(.A(ori_ori_n1159_), .B(ori_ori_n653_), .Y(ori_ori_n1160_));
  NO3        o1132(.A(ori_ori_n796_), .B(ori_ori_n205_), .C(ori_ori_n402_), .Y(ori_ori_n1161_));
  INV        o1133(.A(ori_ori_n1161_), .Y(ori_ori_n1162_));
  NA2        o1134(.A(ori_ori_n1139_), .B(ori_ori_n665_), .Y(ori_ori_n1163_));
  NA4        o1135(.A(ori_ori_n1163_), .B(ori_ori_n1162_), .C(ori_ori_n1160_), .D(ori_ori_n762_), .Y(ori_ori_n1164_));
  NO3        o1136(.A(ori_ori_n1164_), .B(ori_ori_n1158_), .C(ori_ori_n1156_), .Y(ori_ori_n1165_));
  NA2        o1137(.A(ori_ori_n496_), .B(ori_ori_n58_), .Y(ori_ori_n1166_));
  OR3        o1138(.A(ori_ori_n1138_), .B(ori_ori_n591_), .C(ori_ori_n1137_), .Y(ori_ori_n1167_));
  NO2        o1139(.A(ori_ori_n1145_), .B(ori_ori_n940_), .Y(ori_ori_n1168_));
  NO2        o1140(.A(ori_ori_n208_), .B(ori_ori_n110_), .Y(ori_ori_n1169_));
  NO2        o1141(.A(ori_ori_n1169_), .B(ori_ori_n1168_), .Y(ori_ori_n1170_));
  NA4        o1142(.A(ori_ori_n1170_), .B(ori_ori_n1167_), .C(ori_ori_n1166_), .D(ori_ori_n735_), .Y(ori_ori_n1171_));
  NO2        o1143(.A(ori_ori_n929_), .B(ori_ori_n234_), .Y(ori_ori_n1172_));
  NO2        o1144(.A(ori_ori_n930_), .B(ori_ori_n547_), .Y(ori_ori_n1173_));
  OAI210     o1145(.A0(ori_ori_n1173_), .A1(ori_ori_n1172_), .B0(ori_ori_n337_), .Y(ori_ori_n1174_));
  NA2        o1146(.A(ori_ori_n561_), .B(ori_ori_n559_), .Y(ori_ori_n1175_));
  NA2        o1147(.A(ori_ori_n1175_), .B(ori_ori_n659_), .Y(ori_ori_n1176_));
  OR2        o1148(.A(ori_ori_n1092_), .B(ori_ori_n1089_), .Y(ori_ori_n1177_));
  NO2        o1149(.A(ori_ori_n363_), .B(ori_ori_n72_), .Y(ori_ori_n1178_));
  INV        o1150(.A(ori_ori_n1178_), .Y(ori_ori_n1179_));
  NA3        o1151(.A(ori_ori_n1179_), .B(ori_ori_n1177_), .C(ori_ori_n380_), .Y(ori_ori_n1180_));
  NOi41      o1152(.An(ori_ori_n1174_), .B(ori_ori_n1180_), .C(ori_ori_n1176_), .D(ori_ori_n1171_), .Y(ori_ori_n1181_));
  NO2        o1153(.A(ori_ori_n129_), .B(ori_ori_n45_), .Y(ori_ori_n1182_));
  NO2        o1154(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1183_));
  AO220      o1155(.A0(ori_ori_n1183_), .A1(ori_ori_n609_), .B0(ori_ori_n1182_), .B1(ori_ori_n690_), .Y(ori_ori_n1184_));
  NA2        o1156(.A(ori_ori_n1184_), .B(ori_ori_n337_), .Y(ori_ori_n1185_));
  INV        o1157(.A(ori_ori_n133_), .Y(ori_ori_n1186_));
  NO3        o1158(.A(ori_ori_n1023_), .B(ori_ori_n176_), .C(ori_ori_n84_), .Y(ori_ori_n1187_));
  NA2        o1159(.A(ori_ori_n1187_), .B(ori_ori_n1186_), .Y(ori_ori_n1188_));
  NA2        o1160(.A(ori_ori_n1188_), .B(ori_ori_n1185_), .Y(ori_ori_n1189_));
  NO2        o1161(.A(ori_ori_n602_), .B(ori_ori_n601_), .Y(ori_ori_n1190_));
  NO4        o1162(.A(ori_ori_n1023_), .B(ori_ori_n1190_), .C(ori_ori_n174_), .D(ori_ori_n84_), .Y(ori_ori_n1191_));
  NO3        o1163(.A(ori_ori_n1191_), .B(ori_ori_n1189_), .C(ori_ori_n626_), .Y(ori_ori_n1192_));
  NA4        o1164(.A(ori_ori_n1192_), .B(ori_ori_n1181_), .C(ori_ori_n1165_), .D(ori_ori_n1148_), .Y(ori06));
  NO2        o1165(.A(ori_ori_n403_), .B(ori_ori_n551_), .Y(ori_ori_n1194_));
  NA2        o1166(.A(ori_ori_n270_), .B(ori_ori_n1194_), .Y(ori_ori_n1195_));
  NO2        o1167(.A(ori_ori_n226_), .B(ori_ori_n101_), .Y(ori_ori_n1196_));
  OAI210     o1168(.A0(ori_ori_n1196_), .A1(ori_ori_n1187_), .B0(ori_ori_n376_), .Y(ori_ori_n1197_));
  NO3        o1169(.A(ori_ori_n586_), .B(ori_ori_n782_), .C(ori_ori_n588_), .Y(ori_ori_n1198_));
  OR2        o1170(.A(ori_ori_n1198_), .B(ori_ori_n853_), .Y(ori_ori_n1199_));
  NA4        o1171(.A(ori_ori_n1199_), .B(ori_ori_n1197_), .C(ori_ori_n1195_), .D(ori_ori_n1174_), .Y(ori_ori_n1200_));
  NO3        o1172(.A(ori_ori_n1200_), .B(ori_ori_n1176_), .C(ori_ori_n259_), .Y(ori_ori_n1201_));
  NO2        o1173(.A(ori_ori_n297_), .B(ori_ori_n45_), .Y(ori_ori_n1202_));
  AOI210     o1174(.A0(ori_ori_n1202_), .A1(ori_ori_n544_), .B0(ori_ori_n1172_), .Y(ori_ori_n1203_));
  AOI210     o1175(.A0(ori_ori_n1202_), .A1(ori_ori_n548_), .B0(ori_ori_n1184_), .Y(ori_ori_n1204_));
  AOI210     o1176(.A0(ori_ori_n1204_), .A1(ori_ori_n1203_), .B0(ori_ori_n335_), .Y(ori_ori_n1205_));
  OAI210     o1177(.A0(ori_ori_n86_), .A1(ori_ori_n40_), .B0(ori_ori_n663_), .Y(ori_ori_n1206_));
  NA2        o1178(.A(ori_ori_n1206_), .B(ori_ori_n630_), .Y(ori_ori_n1207_));
  NO2        o1179(.A(ori_ori_n506_), .B(ori_ori_n171_), .Y(ori_ori_n1208_));
  NOi21      o1180(.An(ori_ori_n135_), .B(ori_ori_n45_), .Y(ori_ori_n1209_));
  NO2        o1181(.A(ori_ori_n595_), .B(ori_ori_n1040_), .Y(ori_ori_n1210_));
  NO2        o1182(.A(ori_ori_n449_), .B(ori_ori_n250_), .Y(ori_ori_n1211_));
  NO4        o1183(.A(ori_ori_n1211_), .B(ori_ori_n1210_), .C(ori_ori_n1209_), .D(ori_ori_n1208_), .Y(ori_ori_n1212_));
  INV        o1184(.A(ori_ori_n587_), .Y(ori_ori_n1213_));
  NA3        o1185(.A(ori_ori_n1213_), .B(ori_ori_n1212_), .C(ori_ori_n1207_), .Y(ori_ori_n1214_));
  NO2        o1186(.A(ori_ori_n726_), .B(ori_ori_n361_), .Y(ori_ori_n1215_));
  NO3        o1187(.A(ori_ori_n665_), .B(ori_ori_n737_), .C(ori_ori_n622_), .Y(ori_ori_n1216_));
  NOi21      o1188(.An(ori_ori_n1215_), .B(ori_ori_n1216_), .Y(ori_ori_n1217_));
  AN2        o1189(.A(ori_ori_n918_), .B(ori_ori_n633_), .Y(ori_ori_n1218_));
  NO4        o1190(.A(ori_ori_n1218_), .B(ori_ori_n1217_), .C(ori_ori_n1214_), .D(ori_ori_n1205_), .Y(ori_ori_n1219_));
  NO2        o1191(.A(ori_ori_n712_), .B(ori_ori_n47_), .Y(ori_ori_n1220_));
  NA2        o1192(.A(ori_ori_n354_), .B(ori_ori_n1220_), .Y(ori_ori_n1221_));
  NO3        o1193(.A(ori_ori_n245_), .B(ori_ori_n101_), .C(ori_ori_n283_), .Y(ori_ori_n1222_));
  OAI220     o1194(.A0(ori_ori_n683_), .A1(ori_ori_n250_), .B0(ori_ori_n503_), .B1(ori_ori_n506_), .Y(ori_ori_n1223_));
  INV        o1195(.A(k), .Y(ori_ori_n1224_));
  NO3        o1196(.A(ori_ori_n1224_), .B(ori_ori_n585_), .C(j), .Y(ori_ori_n1225_));
  NOi21      o1197(.An(ori_ori_n1225_), .B(ori_ori_n657_), .Y(ori_ori_n1226_));
  NO4        o1198(.A(ori_ori_n1226_), .B(ori_ori_n1223_), .C(ori_ori_n1222_), .D(ori_ori_n1043_), .Y(ori_ori_n1227_));
  NA3        o1199(.A(ori_ori_n1227_), .B(ori_ori_n1221_), .C(ori_ori_n1123_), .Y(ori_ori_n1228_));
  OR3        o1200(.A(ori_ori_n1198_), .B(ori_ori_n759_), .C(ori_ori_n531_), .Y(ori_ori_n1229_));
  AOI210     o1201(.A0(ori_ori_n561_), .A1(ori_ori_n436_), .B0(ori_ori_n367_), .Y(ori_ori_n1230_));
  NA2        o1202(.A(ori_ori_n1225_), .B(ori_ori_n766_), .Y(ori_ori_n1231_));
  NA3        o1203(.A(ori_ori_n1231_), .B(ori_ori_n1230_), .C(ori_ori_n1229_), .Y(ori_ori_n1232_));
  AN2        o1204(.A(ori_ori_n894_), .B(ori_ori_n893_), .Y(ori_ori_n1233_));
  NO3        o1205(.A(ori_ori_n1233_), .B(ori_ori_n492_), .C(ori_ori_n473_), .Y(ori_ori_n1234_));
  INV        o1206(.A(ori_ori_n1234_), .Y(ori_ori_n1235_));
  NAi21      o1207(.An(j), .B(i), .Y(ori_ori_n1236_));
  NO4        o1208(.A(ori_ori_n1190_), .B(ori_ori_n1236_), .C(ori_ori_n430_), .D(ori_ori_n237_), .Y(ori_ori_n1237_));
  NO4        o1209(.A(ori_ori_n1237_), .B(ori_ori_n1235_), .C(ori_ori_n1232_), .D(ori_ori_n1228_), .Y(ori_ori_n1238_));
  NA4        o1210(.A(ori_ori_n1238_), .B(ori_ori_n1219_), .C(ori_ori_n1201_), .D(ori_ori_n1192_), .Y(ori07));
  NOi21      o1211(.An(j), .B(k), .Y(ori_ori_n1240_));
  NA4        o1212(.A(ori_ori_n179_), .B(ori_ori_n107_), .C(ori_ori_n1240_), .D(f), .Y(ori_ori_n1241_));
  NAi32      o1213(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1242_));
  NO3        o1214(.A(ori_ori_n1242_), .B(g), .C(f), .Y(ori_ori_n1243_));
  INV        o1215(.A(ori_ori_n1243_), .Y(ori_ori_n1244_));
  NAi21      o1216(.An(f), .B(c), .Y(ori_ori_n1245_));
  OR2        o1217(.A(e), .B(d), .Y(ori_ori_n1246_));
  NO2        o1218(.A(ori_ori_n614_), .B(ori_ori_n323_), .Y(ori_ori_n1247_));
  NA3        o1219(.A(ori_ori_n1247_), .B(ori_ori_n1006_), .C(ori_ori_n179_), .Y(ori_ori_n1248_));
  NOi31      o1220(.An(n), .B(m), .C(b), .Y(ori_ori_n1249_));
  NA3        o1221(.A(ori_ori_n1248_), .B(ori_ori_n1244_), .C(ori_ori_n1241_), .Y(ori_ori_n1250_));
  NOi41      o1222(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1251_));
  NO2        o1223(.A(k), .B(i), .Y(ori_ori_n1252_));
  NA3        o1224(.A(ori_ori_n1252_), .B(ori_ori_n862_), .C(ori_ori_n179_), .Y(ori_ori_n1253_));
  NA2        o1225(.A(ori_ori_n84_), .B(ori_ori_n45_), .Y(ori_ori_n1254_));
  NO2        o1226(.A(ori_ori_n1004_), .B(ori_ori_n430_), .Y(ori_ori_n1255_));
  NA3        o1227(.A(ori_ori_n1255_), .B(ori_ori_n1254_), .C(ori_ori_n216_), .Y(ori_ori_n1256_));
  NO2        o1228(.A(ori_ori_n1010_), .B(ori_ori_n305_), .Y(ori_ori_n1257_));
  NA2        o1229(.A(ori_ori_n532_), .B(ori_ori_n79_), .Y(ori_ori_n1258_));
  NA2        o1230(.A(ori_ori_n1124_), .B(ori_ori_n291_), .Y(ori_ori_n1259_));
  NA4        o1231(.A(ori_ori_n1259_), .B(ori_ori_n1258_), .C(ori_ori_n1256_), .D(ori_ori_n1253_), .Y(ori_ori_n1260_));
  NO2        o1232(.A(ori_ori_n1260_), .B(ori_ori_n1250_), .Y(ori_ori_n1261_));
  NO3        o1233(.A(e), .B(d), .C(c), .Y(ori_ori_n1262_));
  NO2        o1234(.A(ori_ori_n130_), .B(ori_ori_n216_), .Y(ori_ori_n1263_));
  NA2        o1235(.A(ori_ori_n1263_), .B(ori_ori_n1262_), .Y(ori_ori_n1264_));
  INV        o1236(.A(ori_ori_n1264_), .Y(ori_ori_n1265_));
  OR2        o1237(.A(h), .B(f), .Y(ori_ori_n1266_));
  NO3        o1238(.A(n), .B(m), .C(i), .Y(ori_ori_n1267_));
  OAI210     o1239(.A0(ori_ori_n1041_), .A1(ori_ori_n157_), .B0(ori_ori_n1267_), .Y(ori_ori_n1268_));
  NO2        o1240(.A(ori_ori_n1268_), .B(ori_ori_n1266_), .Y(ori_ori_n1269_));
  NA3        o1241(.A(ori_ori_n680_), .B(ori_ori_n668_), .C(ori_ori_n111_), .Y(ori_ori_n1270_));
  NO2        o1242(.A(ori_ori_n1270_), .B(ori_ori_n45_), .Y(ori_ori_n1271_));
  NO2        o1243(.A(l), .B(k), .Y(ori_ori_n1272_));
  NO3        o1244(.A(ori_ori_n430_), .B(d), .C(c), .Y(ori_ori_n1273_));
  NO3        o1245(.A(ori_ori_n1271_), .B(ori_ori_n1269_), .C(ori_ori_n1265_), .Y(ori_ori_n1274_));
  NO2        o1246(.A(ori_ori_n147_), .B(h), .Y(ori_ori_n1275_));
  NO2        o1247(.A(g), .B(c), .Y(ori_ori_n1276_));
  NO2        o1248(.A(ori_ori_n440_), .B(a), .Y(ori_ori_n1277_));
  NA2        o1249(.A(ori_ori_n1277_), .B(ori_ori_n112_), .Y(ori_ori_n1278_));
  NA2        o1250(.A(ori_ori_n137_), .B(ori_ori_n223_), .Y(ori_ori_n1279_));
  NO2        o1251(.A(ori_ori_n1279_), .B(ori_ori_n1405_), .Y(ori_ori_n1280_));
  NO2        o1252(.A(ori_ori_n733_), .B(ori_ori_n188_), .Y(ori_ori_n1281_));
  NOi31      o1253(.An(m), .B(n), .C(b), .Y(ori_ori_n1282_));
  NOi31      o1254(.An(f), .B(d), .C(c), .Y(ori_ori_n1283_));
  NA2        o1255(.A(ori_ori_n1283_), .B(ori_ori_n1282_), .Y(ori_ori_n1284_));
  INV        o1256(.A(ori_ori_n1284_), .Y(ori_ori_n1285_));
  NO3        o1257(.A(ori_ori_n1285_), .B(ori_ori_n1281_), .C(ori_ori_n1280_), .Y(ori_ori_n1286_));
  NA2        o1258(.A(ori_ori_n1019_), .B(ori_ori_n456_), .Y(ori_ori_n1287_));
  NO2        o1259(.A(ori_ori_n1287_), .B(ori_ori_n430_), .Y(ori_ori_n1288_));
  NO3        o1260(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1289_));
  NO2        o1261(.A(ori_ori_n1009_), .B(ori_ori_n1288_), .Y(ori_ori_n1290_));
  AN3        o1262(.A(ori_ori_n1290_), .B(ori_ori_n1286_), .C(ori_ori_n1278_), .Y(ori_ori_n1291_));
  NA2        o1263(.A(ori_ori_n1249_), .B(ori_ori_n374_), .Y(ori_ori_n1292_));
  INV        o1264(.A(ori_ori_n1292_), .Y(ori_ori_n1293_));
  NA2        o1265(.A(ori_ori_n1273_), .B(ori_ori_n217_), .Y(ori_ori_n1294_));
  NA2        o1266(.A(ori_ori_n1024_), .B(ori_ori_n1287_), .Y(ori_ori_n1295_));
  NAi31      o1267(.An(ori_ori_n1293_), .B(ori_ori_n1295_), .C(ori_ori_n1294_), .Y(ori_ori_n1296_));
  NO4        o1268(.A(ori_ori_n130_), .B(g), .C(f), .D(e), .Y(ori_ori_n1297_));
  NA2        o1269(.A(ori_ori_n195_), .B(ori_ori_n96_), .Y(ori_ori_n1298_));
  NO2        o1270(.A(ori_ori_n1246_), .B(ori_ori_n1245_), .Y(ori_ori_n1299_));
  AOI210     o1271(.A0(ori_ori_n30_), .A1(h), .B0(ori_ori_n1299_), .Y(ori_ori_n1300_));
  NO2        o1272(.A(ori_ori_n1300_), .B(ori_ori_n1016_), .Y(ori_ori_n1301_));
  NA2        o1273(.A(ori_ori_n1251_), .B(ori_ori_n1272_), .Y(ori_ori_n1302_));
  INV        o1274(.A(ori_ori_n1302_), .Y(ori_ori_n1303_));
  OR3        o1275(.A(ori_ori_n531_), .B(ori_ori_n530_), .C(ori_ori_n111_), .Y(ori_ori_n1304_));
  NA2        o1276(.A(ori_ori_n1039_), .B(ori_ori_n402_), .Y(ori_ori_n1305_));
  NO2        o1277(.A(ori_ori_n1305_), .B(ori_ori_n428_), .Y(ori_ori_n1306_));
  AO210      o1278(.A0(ori_ori_n1306_), .A1(ori_ori_n115_), .B0(ori_ori_n1303_), .Y(ori_ori_n1307_));
  NO3        o1279(.A(ori_ori_n1307_), .B(ori_ori_n1301_), .C(ori_ori_n1296_), .Y(ori_ori_n1308_));
  NA4        o1280(.A(ori_ori_n1308_), .B(ori_ori_n1291_), .C(ori_ori_n1274_), .D(ori_ori_n1261_), .Y(ori_ori_n1309_));
  NO2        o1281(.A(ori_ori_n1051_), .B(ori_ori_n109_), .Y(ori_ori_n1310_));
  NA2        o1282(.A(ori_ori_n374_), .B(ori_ori_n56_), .Y(ori_ori_n1311_));
  NA2        o1283(.A(ori_ori_n217_), .B(ori_ori_n179_), .Y(ori_ori_n1312_));
  AOI210     o1284(.A0(ori_ori_n1312_), .A1(ori_ori_n1105_), .B0(ori_ori_n1311_), .Y(ori_ori_n1313_));
  NO2        o1285(.A(ori_ori_n385_), .B(j), .Y(ori_ori_n1314_));
  NA2        o1286(.A(ori_ori_n1289_), .B(ori_ori_n1039_), .Y(ori_ori_n1315_));
  INV        o1287(.A(ori_ori_n1315_), .Y(ori_ori_n1316_));
  NA3        o1288(.A(g), .B(ori_ori_n1314_), .C(ori_ori_n159_), .Y(ori_ori_n1317_));
  INV        o1289(.A(ori_ori_n1317_), .Y(ori_ori_n1318_));
  NO3        o1290(.A(ori_ori_n726_), .B(ori_ori_n174_), .C(ori_ori_n405_), .Y(ori_ori_n1319_));
  NO3        o1291(.A(ori_ori_n1319_), .B(ori_ori_n1318_), .C(ori_ori_n1316_), .Y(ori_ori_n1320_));
  AOI210     o1292(.A0(ori_ori_n1312_), .A1(ori_ori_n1298_), .B0(ori_ori_n1004_), .Y(ori_ori_n1321_));
  OR2        o1293(.A(n), .B(i), .Y(ori_ori_n1322_));
  NA2        o1294(.A(ori_ori_n1322_), .B(ori_ori_n49_), .Y(ori_ori_n1323_));
  AOI220     o1295(.A0(ori_ori_n1323_), .A1(ori_ori_n1094_), .B0(ori_ori_n798_), .B1(ori_ori_n195_), .Y(ori_ori_n1324_));
  INV        o1296(.A(ori_ori_n1324_), .Y(ori_ori_n1325_));
  NO2        o1297(.A(ori_ori_n654_), .B(ori_ori_n176_), .Y(ori_ori_n1326_));
  NO3        o1298(.A(ori_ori_n1326_), .B(ori_ori_n1325_), .C(ori_ori_n1321_), .Y(ori_ori_n1327_));
  NO3        o1299(.A(ori_ori_n1027_), .B(ori_ori_n1246_), .C(ori_ori_n49_), .Y(ori_ori_n1328_));
  NO2        o1300(.A(ori_ori_n1016_), .B(h), .Y(ori_ori_n1329_));
  NA3        o1301(.A(ori_ori_n1329_), .B(d), .C(ori_ori_n998_), .Y(ori_ori_n1330_));
  NO2        o1302(.A(ori_ori_n1330_), .B(c), .Y(ori_ori_n1331_));
  NA3        o1303(.A(ori_ori_n1310_), .B(ori_ori_n456_), .C(f), .Y(ori_ori_n1332_));
  NA2        o1304(.A(ori_ori_n179_), .B(ori_ori_n111_), .Y(ori_ori_n1333_));
  NO2        o1305(.A(ori_ori_n1404_), .B(ori_ori_n1332_), .Y(ori_ori_n1334_));
  NO2        o1306(.A(ori_ori_n1236_), .B(ori_ori_n174_), .Y(ori_ori_n1335_));
  NOi21      o1307(.An(d), .B(f), .Y(ori_ori_n1336_));
  NO3        o1308(.A(ori_ori_n1283_), .B(ori_ori_n1336_), .C(ori_ori_n40_), .Y(ori_ori_n1337_));
  NA2        o1309(.A(ori_ori_n1337_), .B(ori_ori_n1335_), .Y(ori_ori_n1338_));
  INV        o1310(.A(ori_ori_n1338_), .Y(ori_ori_n1339_));
  NO3        o1311(.A(ori_ori_n1339_), .B(ori_ori_n1334_), .C(ori_ori_n1331_), .Y(ori_ori_n1340_));
  NA4        o1312(.A(ori_ori_n1340_), .B(ori_ori_n1327_), .C(ori_ori_n1320_), .D(ori_ori_n1406_), .Y(ori_ori_n1341_));
  NA2        o1313(.A(h), .B(ori_ori_n1257_), .Y(ori_ori_n1342_));
  OAI210     o1314(.A0(ori_ori_n1297_), .A1(ori_ori_n1249_), .B0(ori_ori_n850_), .Y(ori_ori_n1343_));
  NO2        o1315(.A(ori_ori_n995_), .B(ori_ori_n130_), .Y(ori_ori_n1344_));
  NA2        o1316(.A(ori_ori_n1344_), .B(ori_ori_n608_), .Y(ori_ori_n1345_));
  NA3        o1317(.A(ori_ori_n1345_), .B(ori_ori_n1343_), .C(ori_ori_n1342_), .Y(ori_ori_n1346_));
  NA2        o1318(.A(ori_ori_n1276_), .B(ori_ori_n1336_), .Y(ori_ori_n1347_));
  NO2        o1319(.A(ori_ori_n1347_), .B(m), .Y(ori_ori_n1348_));
  NO2        o1320(.A(ori_ori_n151_), .B(ori_ori_n181_), .Y(ori_ori_n1349_));
  OAI210     o1321(.A0(ori_ori_n1349_), .A1(ori_ori_n109_), .B0(ori_ori_n1282_), .Y(ori_ori_n1350_));
  INV        o1322(.A(ori_ori_n1350_), .Y(ori_ori_n1351_));
  NO3        o1323(.A(ori_ori_n1351_), .B(ori_ori_n1348_), .C(ori_ori_n1346_), .Y(ori_ori_n1352_));
  NO2        o1324(.A(ori_ori_n1245_), .B(e), .Y(ori_ori_n1353_));
  NA2        o1325(.A(ori_ori_n1353_), .B(ori_ori_n400_), .Y(ori_ori_n1354_));
  BUFFER     o1326(.A(ori_ori_n130_), .Y(ori_ori_n1355_));
  NO2        o1327(.A(ori_ori_n1355_), .B(ori_ori_n1354_), .Y(ori_ori_n1356_));
  NO2        o1328(.A(ori_ori_n1304_), .B(ori_ori_n347_), .Y(ori_ori_n1357_));
  NO2        o1329(.A(ori_ori_n1357_), .B(ori_ori_n1356_), .Y(ori_ori_n1358_));
  NO2        o1330(.A(ori_ori_n181_), .B(c), .Y(ori_ori_n1359_));
  OAI210     o1331(.A0(ori_ori_n1359_), .A1(ori_ori_n1353_), .B0(ori_ori_n179_), .Y(ori_ori_n1360_));
  AOI210     o1332(.A0(ori_ori_n522_), .A1(ori_ori_n361_), .B0(ori_ori_n1360_), .Y(ori_ori_n1361_));
  INV        o1333(.A(ori_ori_n530_), .Y(ori_ori_n1362_));
  AOI210     o1334(.A0(ori_ori_n1362_), .A1(ori_ori_n1273_), .B0(ori_ori_n1328_), .Y(ori_ori_n1363_));
  INV        o1335(.A(ori_ori_n1048_), .Y(ori_ori_n1364_));
  OAI210     o1336(.A0(ori_ori_n1364_), .A1(ori_ori_n69_), .B0(ori_ori_n1363_), .Y(ori_ori_n1365_));
  INV        o1337(.A(ori_ori_n103_), .Y(ori_ori_n1366_));
  OR2        o1338(.A(ori_ori_n1366_), .B(ori_ori_n530_), .Y(ori_ori_n1367_));
  NO2        o1339(.A(ori_ori_n1367_), .B(ori_ori_n174_), .Y(ori_ori_n1368_));
  NA3        o1340(.A(ori_ori_n1025_), .B(ori_ori_n1022_), .C(ori_ori_n223_), .Y(ori_ori_n1369_));
  NO2        o1341(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1370_));
  INV        o1342(.A(ori_ori_n475_), .Y(ori_ori_n1371_));
  NA2        o1343(.A(ori_ori_n1371_), .B(ori_ori_n1370_), .Y(ori_ori_n1372_));
  NO2        o1344(.A(m), .B(i), .Y(ori_ori_n1373_));
  BUFFER     o1345(.A(ori_ori_n1373_), .Y(ori_ori_n1374_));
  NA2        o1346(.A(ori_ori_n1374_), .B(ori_ori_n1275_), .Y(ori_ori_n1375_));
  NA3        o1347(.A(ori_ori_n1375_), .B(ori_ori_n1372_), .C(ori_ori_n1369_), .Y(ori_ori_n1376_));
  NO4        o1348(.A(ori_ori_n1376_), .B(ori_ori_n1368_), .C(ori_ori_n1365_), .D(ori_ori_n1361_), .Y(ori_ori_n1377_));
  NA3        o1349(.A(ori_ori_n1377_), .B(ori_ori_n1358_), .C(ori_ori_n1352_), .Y(ori_ori_n1378_));
  NA3        o1350(.A(ori_ori_n922_), .B(ori_ori_n137_), .C(ori_ori_n46_), .Y(ori_ori_n1379_));
  INV        o1351(.A(ori_ori_n1379_), .Y(ori_ori_n1380_));
  INV        o1352(.A(ori_ori_n185_), .Y(ori_ori_n1381_));
  NA2        o1353(.A(ori_ori_n1381_), .B(ori_ori_n1329_), .Y(ori_ori_n1382_));
  NO2        o1354(.A(ori_ori_n71_), .B(c), .Y(ori_ori_n1383_));
  NA2        o1355(.A(ori_ori_n1335_), .B(ori_ori_n1383_), .Y(ori_ori_n1384_));
  NA2        o1356(.A(ori_ori_n1384_), .B(ori_ori_n1382_), .Y(ori_ori_n1385_));
  NO2        o1357(.A(ori_ori_n1385_), .B(ori_ori_n1380_), .Y(ori_ori_n1386_));
  AOI210     o1358(.A0(ori_ori_n157_), .A1(ori_ori_n56_), .B0(ori_ori_n1353_), .Y(ori_ori_n1387_));
  NO2        o1359(.A(ori_ori_n1387_), .B(ori_ori_n1333_), .Y(ori_ori_n1388_));
  INV        o1360(.A(ori_ori_n1388_), .Y(ori_ori_n1389_));
  AOI220     o1361(.A0(ori_ori_n1373_), .A1(ori_ori_n628_), .B0(ori_ori_n1006_), .B1(ori_ori_n160_), .Y(ori_ori_n1390_));
  NOi31      o1362(.An(ori_ori_n30_), .B(ori_ori_n1390_), .C(n), .Y(ori_ori_n1391_));
  INV        o1363(.A(ori_ori_n1391_), .Y(ori_ori_n1392_));
  NO2        o1364(.A(ori_ori_n1305_), .B(d), .Y(ori_ori_n1393_));
  INV        o1365(.A(ori_ori_n1393_), .Y(ori_ori_n1394_));
  NA4        o1366(.A(ori_ori_n1394_), .B(ori_ori_n1392_), .C(ori_ori_n1389_), .D(ori_ori_n1386_), .Y(ori_ori_n1395_));
  OR4        o1367(.A(ori_ori_n1395_), .B(ori_ori_n1378_), .C(ori_ori_n1341_), .D(ori_ori_n1309_), .Y(ori04));
  NO2        o1368(.A(ori_ori_n1254_), .B(ori_ori_n88_), .Y(ori_ori_n1397_));
  NA2        o1369(.A(ori_ori_n1397_), .B(ori_ori_n1005_), .Y(ori_ori_n1398_));
  INV        o1370(.A(ori_ori_n1398_), .Y(ori_ori_n1399_));
  NO3        o1371(.A(ori_ori_n1399_), .B(ori_ori_n1013_), .C(ori_ori_n1003_), .Y(ori_ori_n1400_));
  NA3        o1372(.A(ori_ori_n1400_), .B(ori_ori_n1037_), .C(ori_ori_n1029_), .Y(ori05));
  INV        o1373(.A(ori_ori_n112_), .Y(ori_ori_n1404_));
  INV        o1374(.A(h), .Y(ori_ori_n1405_));
  INV        o1375(.A(ori_ori_n1313_), .Y(ori_ori_n1406_));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  INV        m0015(.A(i), .Y(mai_mai_n44_));
  AN2        m0016(.A(h), .B(g), .Y(mai_mai_n45_));
  NA2        m0017(.A(mai_mai_n45_), .B(mai_mai_n44_), .Y(mai_mai_n46_));
  NAi21      m0018(.An(n), .B(m), .Y(mai_mai_n47_));
  NOi32      m0019(.An(k), .Bn(h), .C(l), .Y(mai_mai_n48_));
  NOi32      m0020(.An(k), .Bn(h), .C(g), .Y(mai_mai_n49_));
  INV        m0021(.A(mai_mai_n49_), .Y(mai_mai_n50_));
  NO2        m0022(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n43_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n32_), .Y(mai_mai_n53_));
  INV        m0025(.A(c), .Y(mai_mai_n54_));
  NA2        m0026(.A(e), .B(b), .Y(mai_mai_n55_));
  NO2        m0027(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  INV        m0028(.A(d), .Y(mai_mai_n57_));
  NAi21      m0029(.An(i), .B(h), .Y(mai_mai_n58_));
  NAi31      m0030(.An(i), .B(l), .C(j), .Y(mai_mai_n59_));
  NAi41      m0031(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n60_));
  NA2        m0032(.A(g), .B(f), .Y(mai_mai_n61_));
  NO2        m0033(.A(mai_mai_n61_), .B(mai_mai_n60_), .Y(mai_mai_n62_));
  NAi21      m0034(.An(i), .B(j), .Y(mai_mai_n63_));
  NAi32      m0035(.An(n), .Bn(k), .C(m), .Y(mai_mai_n64_));
  NO2        m0036(.A(mai_mai_n64_), .B(mai_mai_n63_), .Y(mai_mai_n65_));
  NAi31      m0037(.An(l), .B(m), .C(k), .Y(mai_mai_n66_));
  NAi41      m0038(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n67_));
  NA2        m0039(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n68_));
  INV        m0040(.A(m), .Y(mai_mai_n69_));
  NOi21      m0041(.An(k), .B(l), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n70_), .B(mai_mai_n69_), .Y(mai_mai_n71_));
  AN4        m0043(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n72_));
  NOi31      m0044(.An(h), .B(g), .C(f), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NAi32      m0046(.An(m), .Bn(k), .C(j), .Y(mai_mai_n75_));
  NOi32      m0047(.An(h), .Bn(g), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n72_), .Y(mai_mai_n77_));
  OA220      m0049(.A0(mai_mai_n77_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .B1(mai_mai_n71_), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n68_), .Y(mai_mai_n79_));
  INV        m0051(.A(n), .Y(mai_mai_n80_));
  NOi32      m0052(.An(e), .Bn(b), .C(d), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  INV        m0054(.A(j), .Y(mai_mai_n83_));
  AN3        m0055(.A(m), .B(k), .C(i), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n85_));
  NAi32      m0057(.An(g), .Bn(f), .C(h), .Y(mai_mai_n86_));
  NAi31      m0058(.An(j), .B(m), .C(l), .Y(mai_mai_n87_));
  NO2        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .Y(mai_mai_n88_));
  NA2        m0060(.A(m), .B(l), .Y(mai_mai_n89_));
  NAi31      m0061(.An(k), .B(j), .C(g), .Y(mai_mai_n90_));
  NO3        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(f), .Y(mai_mai_n91_));
  AN2        m0063(.A(j), .B(g), .Y(mai_mai_n92_));
  NOi32      m0064(.An(m), .Bn(l), .C(i), .Y(mai_mai_n93_));
  NOi21      m0065(.An(g), .B(i), .Y(mai_mai_n94_));
  NOi32      m0066(.An(m), .Bn(j), .C(k), .Y(mai_mai_n95_));
  NO2        m0067(.A(mai_mai_n91_), .B(mai_mai_n88_), .Y(mai_mai_n96_));
  NAi41      m0068(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n97_));
  AN2        m0069(.A(e), .B(b), .Y(mai_mai_n98_));
  NOi31      m0070(.An(c), .B(h), .C(f), .Y(mai_mai_n99_));
  NA2        m0071(.A(mai_mai_n99_), .B(mai_mai_n98_), .Y(mai_mai_n100_));
  NO2        m0072(.A(mai_mai_n100_), .B(mai_mai_n97_), .Y(mai_mai_n101_));
  NOi21      m0073(.An(g), .B(f), .Y(mai_mai_n102_));
  NOi21      m0074(.An(i), .B(h), .Y(mai_mai_n103_));
  NA3        m0075(.A(mai_mai_n103_), .B(mai_mai_n102_), .C(mai_mai_n36_), .Y(mai_mai_n104_));
  INV        m0076(.A(a), .Y(mai_mai_n105_));
  NA2        m0077(.A(mai_mai_n98_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  INV        m0078(.A(l), .Y(mai_mai_n107_));
  NOi21      m0079(.An(m), .B(n), .Y(mai_mai_n108_));
  AN2        m0080(.A(k), .B(h), .Y(mai_mai_n109_));
  NO2        m0081(.A(mai_mai_n104_), .B(mai_mai_n82_), .Y(mai_mai_n110_));
  INV        m0082(.A(b), .Y(mai_mai_n111_));
  NA2        m0083(.A(l), .B(j), .Y(mai_mai_n112_));
  AN2        m0084(.A(k), .B(i), .Y(mai_mai_n113_));
  NA2        m0085(.A(mai_mai_n113_), .B(mai_mai_n112_), .Y(mai_mai_n114_));
  NA2        m0086(.A(g), .B(e), .Y(mai_mai_n115_));
  NOi32      m0087(.An(c), .Bn(a), .C(d), .Y(mai_mai_n116_));
  NA2        m0088(.A(mai_mai_n116_), .B(mai_mai_n108_), .Y(mai_mai_n117_));
  NO4        m0089(.A(mai_mai_n117_), .B(mai_mai_n115_), .C(mai_mai_n114_), .D(mai_mai_n111_), .Y(mai_mai_n118_));
  NO3        m0090(.A(mai_mai_n118_), .B(mai_mai_n110_), .C(mai_mai_n101_), .Y(mai_mai_n119_));
  OAI210     m0091(.A0(mai_mai_n96_), .A1(mai_mai_n82_), .B0(mai_mai_n119_), .Y(mai_mai_n120_));
  NOi31      m0092(.An(k), .B(m), .C(j), .Y(mai_mai_n121_));
  NA3        m0093(.A(mai_mai_n121_), .B(mai_mai_n73_), .C(mai_mai_n72_), .Y(mai_mai_n122_));
  NOi31      m0094(.An(k), .B(m), .C(i), .Y(mai_mai_n123_));
  INV        m0095(.A(mai_mai_n122_), .Y(mai_mai_n124_));
  NOi32      m0096(.An(f), .Bn(b), .C(e), .Y(mai_mai_n125_));
  NAi21      m0097(.An(g), .B(h), .Y(mai_mai_n126_));
  NAi21      m0098(.An(m), .B(n), .Y(mai_mai_n127_));
  NAi21      m0099(.An(j), .B(k), .Y(mai_mai_n128_));
  NO3        m0100(.A(mai_mai_n128_), .B(mai_mai_n127_), .C(mai_mai_n126_), .Y(mai_mai_n129_));
  NAi41      m0101(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n130_));
  NAi31      m0102(.An(j), .B(k), .C(h), .Y(mai_mai_n131_));
  NO3        m0103(.A(mai_mai_n131_), .B(mai_mai_n130_), .C(mai_mai_n127_), .Y(mai_mai_n132_));
  AOI210     m0104(.A0(mai_mai_n129_), .A1(mai_mai_n125_), .B0(mai_mai_n132_), .Y(mai_mai_n133_));
  NO2        m0105(.A(k), .B(j), .Y(mai_mai_n134_));
  AN2        m0106(.A(k), .B(j), .Y(mai_mai_n135_));
  NAi21      m0107(.An(c), .B(b), .Y(mai_mai_n136_));
  NA2        m0108(.A(f), .B(d), .Y(mai_mai_n137_));
  NA2        m0109(.A(h), .B(c), .Y(mai_mai_n138_));
  NAi31      m0110(.An(f), .B(e), .C(b), .Y(mai_mai_n139_));
  NA2        m0111(.A(d), .B(b), .Y(mai_mai_n140_));
  NAi21      m0112(.An(e), .B(f), .Y(mai_mai_n141_));
  NO2        m0113(.A(mai_mai_n141_), .B(mai_mai_n140_), .Y(mai_mai_n142_));
  NA2        m0114(.A(b), .B(a), .Y(mai_mai_n143_));
  NAi21      m0115(.An(e), .B(g), .Y(mai_mai_n144_));
  NAi21      m0116(.An(c), .B(d), .Y(mai_mai_n145_));
  NAi31      m0117(.An(l), .B(k), .C(h), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n127_), .B(mai_mai_n146_), .Y(mai_mai_n147_));
  NA2        m0119(.A(mai_mai_n147_), .B(mai_mai_n142_), .Y(mai_mai_n148_));
  NAi31      m0120(.An(mai_mai_n124_), .B(mai_mai_n148_), .C(mai_mai_n133_), .Y(mai_mai_n149_));
  NAi31      m0121(.An(e), .B(f), .C(b), .Y(mai_mai_n150_));
  NOi21      m0122(.An(g), .B(d), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  NOi21      m0124(.An(h), .B(i), .Y(mai_mai_n153_));
  NOi21      m0125(.An(k), .B(m), .Y(mai_mai_n154_));
  NA3        m0126(.A(mai_mai_n154_), .B(mai_mai_n153_), .C(n), .Y(mai_mai_n155_));
  NOi21      m0127(.An(mai_mai_n152_), .B(mai_mai_n155_), .Y(mai_mai_n156_));
  NOi21      m0128(.An(h), .B(g), .Y(mai_mai_n157_));
  NO2        m0129(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NOi32      m0131(.An(n), .Bn(k), .C(m), .Y(mai_mai_n160_));
  NA2        m0132(.A(l), .B(i), .Y(mai_mai_n161_));
  NA2        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n162_), .B(mai_mai_n159_), .Y(mai_mai_n163_));
  NAi31      m0135(.An(d), .B(f), .C(c), .Y(mai_mai_n164_));
  NAi31      m0136(.An(e), .B(f), .C(c), .Y(mai_mai_n165_));
  NA2        m0137(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  NA2        m0138(.A(j), .B(h), .Y(mai_mai_n167_));
  OR3        m0139(.A(n), .B(m), .C(k), .Y(mai_mai_n168_));
  NO2        m0140(.A(mai_mai_n168_), .B(mai_mai_n167_), .Y(mai_mai_n169_));
  NAi32      m0141(.An(m), .Bn(k), .C(n), .Y(mai_mai_n170_));
  NO2        m0142(.A(mai_mai_n170_), .B(mai_mai_n167_), .Y(mai_mai_n171_));
  AOI220     m0143(.A0(mai_mai_n171_), .A1(mai_mai_n152_), .B0(mai_mai_n169_), .B1(mai_mai_n166_), .Y(mai_mai_n172_));
  NO2        m0144(.A(n), .B(m), .Y(mai_mai_n173_));
  NA2        m0145(.A(mai_mai_n173_), .B(mai_mai_n48_), .Y(mai_mai_n174_));
  NAi21      m0146(.An(f), .B(e), .Y(mai_mai_n175_));
  NA2        m0147(.A(d), .B(c), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  NOi21      m0149(.An(mai_mai_n177_), .B(mai_mai_n174_), .Y(mai_mai_n178_));
  NAi21      m0150(.An(d), .B(c), .Y(mai_mai_n179_));
  NAi31      m0151(.An(m), .B(n), .C(b), .Y(mai_mai_n180_));
  NA2        m0152(.A(k), .B(i), .Y(mai_mai_n181_));
  NAi21      m0153(.An(h), .B(f), .Y(mai_mai_n182_));
  NO2        m0154(.A(mai_mai_n182_), .B(mai_mai_n181_), .Y(mai_mai_n183_));
  NO2        m0155(.A(mai_mai_n180_), .B(mai_mai_n145_), .Y(mai_mai_n184_));
  NA2        m0156(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  NOi32      m0157(.An(f), .Bn(c), .C(d), .Y(mai_mai_n186_));
  NOi32      m0158(.An(f), .Bn(c), .C(e), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n187_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  NO3        m0160(.A(n), .B(m), .C(j), .Y(mai_mai_n189_));
  NA2        m0161(.A(mai_mai_n189_), .B(mai_mai_n109_), .Y(mai_mai_n190_));
  AO210      m0162(.A0(mai_mai_n190_), .A1(mai_mai_n174_), .B0(mai_mai_n188_), .Y(mai_mai_n191_));
  NAi41      m0163(.An(mai_mai_n178_), .B(mai_mai_n191_), .C(mai_mai_n185_), .D(mai_mai_n172_), .Y(mai_mai_n192_));
  OR4        m0164(.A(mai_mai_n192_), .B(mai_mai_n163_), .C(mai_mai_n156_), .D(mai_mai_n149_), .Y(mai_mai_n193_));
  NO4        m0165(.A(mai_mai_n193_), .B(mai_mai_n120_), .C(mai_mai_n79_), .D(mai_mai_n53_), .Y(mai_mai_n194_));
  NA3        m0166(.A(m), .B(mai_mai_n107_), .C(j), .Y(mai_mai_n195_));
  NAi31      m0167(.An(n), .B(h), .C(g), .Y(mai_mai_n196_));
  NO2        m0168(.A(mai_mai_n196_), .B(mai_mai_n195_), .Y(mai_mai_n197_));
  NOi32      m0169(.An(m), .Bn(k), .C(l), .Y(mai_mai_n198_));
  NA3        m0170(.A(mai_mai_n198_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n199_));
  NO2        m0171(.A(mai_mai_n199_), .B(n), .Y(mai_mai_n200_));
  AN2        m0172(.A(i), .B(g), .Y(mai_mai_n201_));
  NA3        m0173(.A(mai_mai_n70_), .B(mai_mai_n201_), .C(mai_mai_n108_), .Y(mai_mai_n202_));
  INV        m0174(.A(mai_mai_n200_), .Y(mai_mai_n203_));
  NAi41      m0175(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n204_));
  INV        m0176(.A(mai_mai_n204_), .Y(mai_mai_n205_));
  INV        m0177(.A(f), .Y(mai_mai_n206_));
  INV        m0178(.A(g), .Y(mai_mai_n207_));
  NOi31      m0179(.An(i), .B(j), .C(h), .Y(mai_mai_n208_));
  NOi21      m0180(.An(l), .B(m), .Y(mai_mai_n209_));
  NA2        m0181(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  NO3        m0182(.A(mai_mai_n210_), .B(mai_mai_n207_), .C(mai_mai_n206_), .Y(mai_mai_n211_));
  NA2        m0183(.A(mai_mai_n211_), .B(mai_mai_n205_), .Y(mai_mai_n212_));
  OAI210     m0184(.A0(mai_mai_n203_), .A1(mai_mai_n32_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  NOi21      m0185(.An(n), .B(m), .Y(mai_mai_n214_));
  NOi32      m0186(.An(l), .Bn(i), .C(j), .Y(mai_mai_n215_));
  NA2        m0187(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n216_));
  OA220      m0188(.A0(mai_mai_n216_), .A1(mai_mai_n100_), .B0(mai_mai_n75_), .B1(mai_mai_n74_), .Y(mai_mai_n217_));
  NAi21      m0189(.An(j), .B(h), .Y(mai_mai_n218_));
  XN2        m0190(.A(i), .B(h), .Y(mai_mai_n219_));
  NA2        m0191(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  NOi31      m0192(.An(k), .B(n), .C(m), .Y(mai_mai_n221_));
  NOi31      m0193(.An(mai_mai_n221_), .B(mai_mai_n176_), .C(mai_mai_n175_), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n220_), .Y(mai_mai_n223_));
  NAi31      m0195(.An(f), .B(e), .C(c), .Y(mai_mai_n224_));
  NO4        m0196(.A(mai_mai_n224_), .B(mai_mai_n168_), .C(mai_mai_n167_), .D(mai_mai_n57_), .Y(mai_mai_n225_));
  NA3        m0197(.A(e), .B(c), .C(b), .Y(mai_mai_n226_));
  NAi32      m0198(.An(m), .Bn(i), .C(k), .Y(mai_mai_n227_));
  INV        m0199(.A(k), .Y(mai_mai_n228_));
  INV        m0200(.A(mai_mai_n225_), .Y(mai_mai_n229_));
  NAi21      m0201(.An(n), .B(a), .Y(mai_mai_n230_));
  NO2        m0202(.A(mai_mai_n230_), .B(mai_mai_n140_), .Y(mai_mai_n231_));
  NAi41      m0203(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n232_));
  NO2        m0204(.A(mai_mai_n232_), .B(e), .Y(mai_mai_n233_));
  NO3        m0205(.A(mai_mai_n141_), .B(mai_mai_n90_), .C(mai_mai_n89_), .Y(mai_mai_n234_));
  OAI210     m0206(.A0(mai_mai_n234_), .A1(mai_mai_n233_), .B0(mai_mai_n231_), .Y(mai_mai_n235_));
  AN4        m0207(.A(mai_mai_n235_), .B(mai_mai_n229_), .C(mai_mai_n223_), .D(mai_mai_n217_), .Y(mai_mai_n236_));
  OR2        m0208(.A(h), .B(g), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n237_), .B(mai_mai_n97_), .Y(mai_mai_n238_));
  NA2        m0210(.A(mai_mai_n238_), .B(mai_mai_n125_), .Y(mai_mai_n239_));
  NAi41      m0211(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n240_), .B(mai_mai_n206_), .Y(mai_mai_n241_));
  NA2        m0213(.A(mai_mai_n154_), .B(mai_mai_n103_), .Y(mai_mai_n242_));
  NAi21      m0214(.An(mai_mai_n242_), .B(mai_mai_n241_), .Y(mai_mai_n243_));
  NO2        m0215(.A(n), .B(a), .Y(mai_mai_n244_));
  NAi31      m0216(.An(mai_mai_n232_), .B(mai_mai_n244_), .C(mai_mai_n98_), .Y(mai_mai_n245_));
  AN2        m0217(.A(mai_mai_n245_), .B(mai_mai_n243_), .Y(mai_mai_n246_));
  NAi21      m0218(.An(h), .B(i), .Y(mai_mai_n247_));
  NA2        m0219(.A(mai_mai_n173_), .B(k), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n248_), .B(mai_mai_n247_), .Y(mai_mai_n249_));
  NA2        m0221(.A(mai_mai_n249_), .B(mai_mai_n186_), .Y(mai_mai_n250_));
  NA3        m0222(.A(mai_mai_n250_), .B(mai_mai_n246_), .C(mai_mai_n239_), .Y(mai_mai_n251_));
  NOi21      m0223(.An(g), .B(e), .Y(mai_mai_n252_));
  NO2        m0224(.A(mai_mai_n67_), .B(mai_mai_n69_), .Y(mai_mai_n253_));
  NOi32      m0225(.An(l), .Bn(j), .C(i), .Y(mai_mai_n254_));
  AOI210     m0226(.A0(mai_mai_n70_), .A1(mai_mai_n83_), .B0(mai_mai_n254_), .Y(mai_mai_n255_));
  NAi21      m0227(.An(f), .B(g), .Y(mai_mai_n256_));
  NO2        m0228(.A(mai_mai_n256_), .B(mai_mai_n60_), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n64_), .B(mai_mai_n112_), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n258_), .B(mai_mai_n257_), .Y(mai_mai_n259_));
  INV        m0231(.A(mai_mai_n259_), .Y(mai_mai_n260_));
  NO3        m0232(.A(mai_mai_n128_), .B(mai_mai_n47_), .C(mai_mai_n44_), .Y(mai_mai_n261_));
  NOi41      m0233(.An(mai_mai_n236_), .B(mai_mai_n260_), .C(mai_mai_n251_), .D(mai_mai_n213_), .Y(mai_mai_n262_));
  NO3        m0234(.A(mai_mai_n197_), .B(mai_mai_n43_), .C(mai_mai_n39_), .Y(mai_mai_n263_));
  NO2        m0235(.A(mai_mai_n263_), .B(mai_mai_n106_), .Y(mai_mai_n264_));
  NA3        m0236(.A(mai_mai_n57_), .B(c), .C(b), .Y(mai_mai_n265_));
  NAi21      m0237(.An(h), .B(g), .Y(mai_mai_n266_));
  NO2        m0238(.A(mai_mai_n242_), .B(mai_mai_n256_), .Y(mai_mai_n267_));
  NAi31      m0239(.An(g), .B(k), .C(h), .Y(mai_mai_n268_));
  NO3        m0240(.A(mai_mai_n127_), .B(mai_mai_n268_), .C(l), .Y(mai_mai_n269_));
  NAi31      m0241(.An(e), .B(d), .C(a), .Y(mai_mai_n270_));
  NA2        m0242(.A(mai_mai_n269_), .B(mai_mai_n125_), .Y(mai_mai_n271_));
  INV        m0243(.A(mai_mai_n271_), .Y(mai_mai_n272_));
  NA4        m0244(.A(mai_mai_n154_), .B(mai_mai_n76_), .C(mai_mai_n72_), .D(mai_mai_n112_), .Y(mai_mai_n273_));
  NA3        m0245(.A(mai_mai_n154_), .B(mai_mai_n153_), .C(mai_mai_n80_), .Y(mai_mai_n274_));
  NO2        m0246(.A(mai_mai_n274_), .B(mai_mai_n188_), .Y(mai_mai_n275_));
  NOi21      m0247(.An(mai_mai_n273_), .B(mai_mai_n275_), .Y(mai_mai_n276_));
  NA3        m0248(.A(e), .B(c), .C(b), .Y(mai_mai_n277_));
  NAi32      m0249(.An(k), .Bn(i), .C(j), .Y(mai_mai_n278_));
  NAi21      m0250(.An(l), .B(k), .Y(mai_mai_n279_));
  NO2        m0251(.A(mai_mai_n279_), .B(mai_mai_n47_), .Y(mai_mai_n280_));
  NOi21      m0252(.An(l), .B(j), .Y(mai_mai_n281_));
  NA2        m0253(.A(mai_mai_n157_), .B(mai_mai_n281_), .Y(mai_mai_n282_));
  NA3        m0254(.A(mai_mai_n113_), .B(mai_mai_n112_), .C(g), .Y(mai_mai_n283_));
  OR3        m0255(.A(mai_mai_n67_), .B(mai_mai_n69_), .C(e), .Y(mai_mai_n284_));
  AOI210     m0256(.A0(mai_mai_n283_), .A1(mai_mai_n282_), .B0(mai_mai_n284_), .Y(mai_mai_n285_));
  INV        m0257(.A(mai_mai_n285_), .Y(mai_mai_n286_));
  NAi32      m0258(.An(j), .Bn(h), .C(i), .Y(mai_mai_n287_));
  NAi21      m0259(.An(m), .B(l), .Y(mai_mai_n288_));
  NO3        m0260(.A(mai_mai_n288_), .B(mai_mai_n287_), .C(mai_mai_n80_), .Y(mai_mai_n289_));
  NA2        m0261(.A(h), .B(g), .Y(mai_mai_n290_));
  NA2        m0262(.A(mai_mai_n289_), .B(mai_mai_n158_), .Y(mai_mai_n291_));
  NA3        m0263(.A(mai_mai_n291_), .B(mai_mai_n286_), .C(mai_mai_n276_), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n139_), .B(d), .Y(mai_mai_n293_));
  NA2        m0265(.A(mai_mai_n293_), .B(mai_mai_n51_), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n100_), .B(mai_mai_n97_), .Y(mai_mai_n295_));
  NAi32      m0267(.An(n), .Bn(m), .C(l), .Y(mai_mai_n296_));
  NO2        m0268(.A(mai_mai_n296_), .B(mai_mai_n287_), .Y(mai_mai_n297_));
  NA2        m0269(.A(mai_mai_n297_), .B(mai_mai_n177_), .Y(mai_mai_n298_));
  NO2        m0270(.A(mai_mai_n117_), .B(mai_mai_n111_), .Y(mai_mai_n299_));
  NAi31      m0271(.An(k), .B(l), .C(j), .Y(mai_mai_n300_));
  OAI210     m0272(.A0(mai_mai_n279_), .A1(j), .B0(mai_mai_n300_), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n298_), .B(mai_mai_n294_), .Y(mai_mai_n302_));
  NO4        m0274(.A(mai_mai_n302_), .B(mai_mai_n292_), .C(mai_mai_n272_), .D(mai_mai_n264_), .Y(mai_mai_n303_));
  NA2        m0275(.A(mai_mai_n249_), .B(mai_mai_n187_), .Y(mai_mai_n304_));
  NAi21      m0276(.An(m), .B(k), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n219_), .B(mai_mai_n305_), .Y(mai_mai_n306_));
  NAi41      m0278(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n307_), .B(mai_mai_n144_), .Y(mai_mai_n308_));
  NA2        m0280(.A(mai_mai_n308_), .B(mai_mai_n306_), .Y(mai_mai_n309_));
  NAi31      m0281(.An(i), .B(l), .C(h), .Y(mai_mai_n310_));
  NO4        m0282(.A(mai_mai_n310_), .B(mai_mai_n144_), .C(mai_mai_n67_), .D(mai_mai_n69_), .Y(mai_mai_n311_));
  NA2        m0283(.A(e), .B(c), .Y(mai_mai_n312_));
  NO3        m0284(.A(mai_mai_n312_), .B(n), .C(d), .Y(mai_mai_n313_));
  NOi21      m0285(.An(f), .B(h), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n314_), .B(mai_mai_n113_), .Y(mai_mai_n315_));
  NO2        m0287(.A(mai_mai_n315_), .B(mai_mai_n207_), .Y(mai_mai_n316_));
  NAi31      m0288(.An(d), .B(e), .C(b), .Y(mai_mai_n317_));
  NO2        m0289(.A(mai_mai_n127_), .B(mai_mai_n317_), .Y(mai_mai_n318_));
  NA2        m0290(.A(mai_mai_n318_), .B(mai_mai_n316_), .Y(mai_mai_n319_));
  NAi41      m0291(.An(mai_mai_n311_), .B(mai_mai_n319_), .C(mai_mai_n309_), .D(mai_mai_n304_), .Y(mai_mai_n320_));
  NA2        m0292(.A(mai_mai_n244_), .B(mai_mai_n98_), .Y(mai_mai_n321_));
  OR2        m0293(.A(mai_mai_n321_), .B(mai_mai_n199_), .Y(mai_mai_n322_));
  NOi31      m0294(.An(l), .B(n), .C(m), .Y(mai_mai_n323_));
  NA2        m0295(.A(mai_mai_n323_), .B(mai_mai_n208_), .Y(mai_mai_n324_));
  NO2        m0296(.A(mai_mai_n324_), .B(mai_mai_n188_), .Y(mai_mai_n325_));
  NAi21      m0297(.An(mai_mai_n325_), .B(mai_mai_n322_), .Y(mai_mai_n326_));
  NAi32      m0298(.An(m), .Bn(j), .C(k), .Y(mai_mai_n327_));
  NAi41      m0299(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n328_));
  OAI210     m0300(.A0(mai_mai_n204_), .A1(mai_mai_n327_), .B0(mai_mai_n328_), .Y(mai_mai_n329_));
  NOi31      m0301(.An(j), .B(m), .C(k), .Y(mai_mai_n330_));
  NO2        m0302(.A(mai_mai_n121_), .B(mai_mai_n330_), .Y(mai_mai_n331_));
  AN3        m0303(.A(h), .B(g), .C(f), .Y(mai_mai_n332_));
  NAi31      m0304(.An(mai_mai_n331_), .B(mai_mai_n332_), .C(mai_mai_n329_), .Y(mai_mai_n333_));
  NOi32      m0305(.An(m), .Bn(j), .C(l), .Y(mai_mai_n334_));
  NO2        m0306(.A(mai_mai_n334_), .B(mai_mai_n93_), .Y(mai_mai_n335_));
  NAi32      m0307(.An(mai_mai_n335_), .Bn(mai_mai_n196_), .C(mai_mai_n293_), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n288_), .B(mai_mai_n287_), .Y(mai_mai_n337_));
  NO2        m0309(.A(mai_mai_n210_), .B(g), .Y(mai_mai_n338_));
  NO2        m0310(.A(mai_mai_n150_), .B(mai_mai_n80_), .Y(mai_mai_n339_));
  AOI220     m0311(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n241_), .B1(mai_mai_n337_), .Y(mai_mai_n340_));
  NA2        m0312(.A(mai_mai_n227_), .B(mai_mai_n75_), .Y(mai_mai_n341_));
  NA3        m0313(.A(mai_mai_n341_), .B(mai_mai_n332_), .C(mai_mai_n205_), .Y(mai_mai_n342_));
  NA4        m0314(.A(mai_mai_n342_), .B(mai_mai_n340_), .C(mai_mai_n336_), .D(mai_mai_n333_), .Y(mai_mai_n343_));
  NA3        m0315(.A(h), .B(g), .C(f), .Y(mai_mai_n344_));
  NO2        m0316(.A(mai_mai_n344_), .B(mai_mai_n71_), .Y(mai_mai_n345_));
  NA2        m0317(.A(mai_mai_n328_), .B(mai_mai_n204_), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n157_), .B(e), .Y(mai_mai_n347_));
  NO2        m0319(.A(mai_mai_n347_), .B(mai_mai_n41_), .Y(mai_mai_n348_));
  AOI220     m0320(.A0(mai_mai_n348_), .A1(mai_mai_n299_), .B0(mai_mai_n346_), .B1(mai_mai_n345_), .Y(mai_mai_n349_));
  NOi32      m0321(.An(j), .Bn(g), .C(i), .Y(mai_mai_n350_));
  NA3        m0322(.A(mai_mai_n350_), .B(mai_mai_n279_), .C(mai_mai_n108_), .Y(mai_mai_n351_));
  AO210      m0323(.A0(mai_mai_n106_), .A1(mai_mai_n32_), .B0(mai_mai_n351_), .Y(mai_mai_n352_));
  NOi32      m0324(.An(e), .Bn(b), .C(a), .Y(mai_mai_n353_));
  AN2        m0325(.A(l), .B(j), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n202_), .B(mai_mai_n35_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n355_), .B(mai_mai_n353_), .Y(mai_mai_n356_));
  NO2        m0328(.A(mai_mai_n317_), .B(n), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n201_), .B(k), .Y(mai_mai_n358_));
  NA3        m0330(.A(m), .B(mai_mai_n107_), .C(mai_mai_n206_), .Y(mai_mai_n359_));
  NA4        m0331(.A(mai_mai_n198_), .B(mai_mai_n83_), .C(g), .D(mai_mai_n206_), .Y(mai_mai_n360_));
  OAI210     m0332(.A0(mai_mai_n359_), .A1(mai_mai_n358_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  NAi41      m0333(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n362_));
  NA2        m0334(.A(mai_mai_n49_), .B(mai_mai_n108_), .Y(mai_mai_n363_));
  NA2        m0335(.A(mai_mai_n361_), .B(mai_mai_n357_), .Y(mai_mai_n364_));
  NA4        m0336(.A(mai_mai_n364_), .B(mai_mai_n356_), .C(mai_mai_n352_), .D(mai_mai_n349_), .Y(mai_mai_n365_));
  NO4        m0337(.A(mai_mai_n365_), .B(mai_mai_n343_), .C(mai_mai_n326_), .D(mai_mai_n320_), .Y(mai_mai_n366_));
  NA4        m0338(.A(mai_mai_n366_), .B(mai_mai_n303_), .C(mai_mai_n262_), .D(mai_mai_n194_), .Y(mai10));
  NA3        m0339(.A(m), .B(k), .C(i), .Y(mai_mai_n368_));
  NO3        m0340(.A(mai_mai_n368_), .B(j), .C(mai_mai_n207_), .Y(mai_mai_n369_));
  NOi21      m0341(.An(e), .B(f), .Y(mai_mai_n370_));
  NO4        m0342(.A(mai_mai_n145_), .B(mai_mai_n370_), .C(n), .D(mai_mai_n105_), .Y(mai_mai_n371_));
  NAi31      m0343(.An(b), .B(f), .C(c), .Y(mai_mai_n372_));
  INV        m0344(.A(mai_mai_n372_), .Y(mai_mai_n373_));
  NOi32      m0345(.An(k), .Bn(h), .C(j), .Y(mai_mai_n374_));
  NA2        m0346(.A(mai_mai_n374_), .B(mai_mai_n214_), .Y(mai_mai_n375_));
  NA2        m0347(.A(mai_mai_n155_), .B(mai_mai_n375_), .Y(mai_mai_n376_));
  AOI220     m0348(.A0(mai_mai_n376_), .A1(mai_mai_n373_), .B0(mai_mai_n371_), .B1(mai_mai_n369_), .Y(mai_mai_n377_));
  AN2        m0349(.A(j), .B(h), .Y(mai_mai_n378_));
  NO3        m0350(.A(n), .B(m), .C(k), .Y(mai_mai_n379_));
  NA2        m0351(.A(mai_mai_n379_), .B(mai_mai_n378_), .Y(mai_mai_n380_));
  NO3        m0352(.A(mai_mai_n380_), .B(mai_mai_n145_), .C(mai_mai_n206_), .Y(mai_mai_n381_));
  OR2        m0353(.A(m), .B(k), .Y(mai_mai_n382_));
  NO2        m0354(.A(mai_mai_n167_), .B(mai_mai_n382_), .Y(mai_mai_n383_));
  NA4        m0355(.A(n), .B(f), .C(c), .D(mai_mai_n111_), .Y(mai_mai_n384_));
  NOi21      m0356(.An(mai_mai_n383_), .B(mai_mai_n384_), .Y(mai_mai_n385_));
  NOi32      m0357(.An(d), .Bn(a), .C(c), .Y(mai_mai_n386_));
  NA2        m0358(.A(mai_mai_n386_), .B(mai_mai_n175_), .Y(mai_mai_n387_));
  NAi21      m0359(.An(i), .B(g), .Y(mai_mai_n388_));
  NAi31      m0360(.An(k), .B(m), .C(j), .Y(mai_mai_n389_));
  NO3        m0361(.A(mai_mai_n389_), .B(mai_mai_n388_), .C(n), .Y(mai_mai_n390_));
  NO2        m0362(.A(mai_mai_n385_), .B(mai_mai_n381_), .Y(mai_mai_n391_));
  NO2        m0363(.A(mai_mai_n384_), .B(mai_mai_n288_), .Y(mai_mai_n392_));
  NOi32      m0364(.An(f), .Bn(d), .C(c), .Y(mai_mai_n393_));
  AOI220     m0365(.A0(mai_mai_n393_), .A1(mai_mai_n297_), .B0(mai_mai_n392_), .B1(mai_mai_n208_), .Y(mai_mai_n394_));
  NA3        m0366(.A(mai_mai_n394_), .B(mai_mai_n391_), .C(mai_mai_n377_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n57_), .B(mai_mai_n111_), .Y(mai_mai_n396_));
  NA2        m0368(.A(mai_mai_n244_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  INV        m0369(.A(e), .Y(mai_mai_n398_));
  NA2        m0370(.A(mai_mai_n45_), .B(e), .Y(mai_mai_n399_));
  OAI220     m0371(.A0(mai_mai_n399_), .A1(mai_mai_n195_), .B0(mai_mai_n199_), .B1(mai_mai_n398_), .Y(mai_mai_n400_));
  AN2        m0372(.A(g), .B(e), .Y(mai_mai_n401_));
  INV        m0373(.A(mai_mai_n400_), .Y(mai_mai_n402_));
  NOi32      m0374(.An(h), .Bn(e), .C(g), .Y(mai_mai_n403_));
  NA3        m0375(.A(mai_mai_n403_), .B(mai_mai_n281_), .C(m), .Y(mai_mai_n404_));
  NOi21      m0376(.An(g), .B(h), .Y(mai_mai_n405_));
  AN3        m0377(.A(m), .B(l), .C(i), .Y(mai_mai_n406_));
  AN3        m0378(.A(h), .B(g), .C(e), .Y(mai_mai_n407_));
  AOI210     m0379(.A0(mai_mai_n404_), .A1(mai_mai_n402_), .B0(mai_mai_n397_), .Y(mai_mai_n408_));
  NA3        m0380(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n409_));
  NO2        m0381(.A(mai_mai_n409_), .B(mai_mai_n397_), .Y(mai_mai_n410_));
  NA3        m0382(.A(mai_mai_n386_), .B(mai_mai_n175_), .C(mai_mai_n80_), .Y(mai_mai_n411_));
  NAi31      m0383(.An(b), .B(c), .C(a), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n412_), .B(n), .Y(mai_mai_n413_));
  NA2        m0385(.A(mai_mai_n49_), .B(m), .Y(mai_mai_n414_));
  NO2        m0386(.A(mai_mai_n414_), .B(mai_mai_n141_), .Y(mai_mai_n415_));
  NA2        m0387(.A(mai_mai_n415_), .B(mai_mai_n413_), .Y(mai_mai_n416_));
  INV        m0388(.A(mai_mai_n416_), .Y(mai_mai_n417_));
  NO4        m0389(.A(mai_mai_n417_), .B(mai_mai_n410_), .C(mai_mai_n408_), .D(mai_mai_n395_), .Y(mai_mai_n418_));
  NA2        m0390(.A(i), .B(g), .Y(mai_mai_n419_));
  NO3        m0391(.A(mai_mai_n270_), .B(mai_mai_n419_), .C(c), .Y(mai_mai_n420_));
  NOi21      m0392(.An(a), .B(n), .Y(mai_mai_n421_));
  NOi21      m0393(.An(d), .B(c), .Y(mai_mai_n422_));
  NA2        m0394(.A(mai_mai_n422_), .B(mai_mai_n421_), .Y(mai_mai_n423_));
  NA3        m0395(.A(i), .B(g), .C(f), .Y(mai_mai_n424_));
  OR2        m0396(.A(mai_mai_n424_), .B(mai_mai_n66_), .Y(mai_mai_n425_));
  NA3        m0397(.A(mai_mai_n406_), .B(mai_mai_n405_), .C(mai_mai_n175_), .Y(mai_mai_n426_));
  AOI210     m0398(.A0(mai_mai_n426_), .A1(mai_mai_n425_), .B0(mai_mai_n423_), .Y(mai_mai_n427_));
  AOI210     m0399(.A0(mai_mai_n420_), .A1(mai_mai_n280_), .B0(mai_mai_n427_), .Y(mai_mai_n428_));
  OR2        m0400(.A(n), .B(m), .Y(mai_mai_n429_));
  NO2        m0401(.A(mai_mai_n429_), .B(mai_mai_n146_), .Y(mai_mai_n430_));
  NO2        m0402(.A(mai_mai_n176_), .B(mai_mai_n141_), .Y(mai_mai_n431_));
  OAI210     m0403(.A0(mai_mai_n430_), .A1(mai_mai_n169_), .B0(mai_mai_n431_), .Y(mai_mai_n432_));
  INV        m0404(.A(mai_mai_n363_), .Y(mai_mai_n433_));
  NA3        m0405(.A(mai_mai_n433_), .B(mai_mai_n353_), .C(d), .Y(mai_mai_n434_));
  NO2        m0406(.A(mai_mai_n412_), .B(mai_mai_n47_), .Y(mai_mai_n435_));
  NO3        m0407(.A(mai_mai_n61_), .B(mai_mai_n107_), .C(e), .Y(mai_mai_n436_));
  NAi21      m0408(.An(k), .B(j), .Y(mai_mai_n437_));
  NA2        m0409(.A(mai_mai_n247_), .B(mai_mai_n437_), .Y(mai_mai_n438_));
  NA3        m0410(.A(mai_mai_n438_), .B(mai_mai_n436_), .C(mai_mai_n435_), .Y(mai_mai_n439_));
  NAi21      m0411(.An(e), .B(d), .Y(mai_mai_n440_));
  INV        m0412(.A(mai_mai_n440_), .Y(mai_mai_n441_));
  NO2        m0413(.A(mai_mai_n248_), .B(mai_mai_n206_), .Y(mai_mai_n442_));
  NA3        m0414(.A(mai_mai_n442_), .B(mai_mai_n441_), .C(mai_mai_n220_), .Y(mai_mai_n443_));
  NA4        m0415(.A(mai_mai_n443_), .B(mai_mai_n439_), .C(mai_mai_n434_), .D(mai_mai_n432_), .Y(mai_mai_n444_));
  NO2        m0416(.A(mai_mai_n324_), .B(mai_mai_n206_), .Y(mai_mai_n445_));
  NA2        m0417(.A(mai_mai_n445_), .B(mai_mai_n441_), .Y(mai_mai_n446_));
  NOi31      m0418(.An(n), .B(m), .C(k), .Y(mai_mai_n447_));
  AOI220     m0419(.A0(mai_mai_n447_), .A1(mai_mai_n378_), .B0(mai_mai_n214_), .B1(mai_mai_n48_), .Y(mai_mai_n448_));
  NAi31      m0420(.An(g), .B(f), .C(c), .Y(mai_mai_n449_));
  OR3        m0421(.A(mai_mai_n449_), .B(mai_mai_n448_), .C(e), .Y(mai_mai_n450_));
  NA3        m0422(.A(mai_mai_n450_), .B(mai_mai_n446_), .C(mai_mai_n298_), .Y(mai_mai_n451_));
  NOi41      m0423(.An(mai_mai_n428_), .B(mai_mai_n451_), .C(mai_mai_n444_), .D(mai_mai_n260_), .Y(mai_mai_n452_));
  NOi32      m0424(.An(c), .Bn(a), .C(b), .Y(mai_mai_n453_));
  NA2        m0425(.A(mai_mai_n453_), .B(mai_mai_n108_), .Y(mai_mai_n454_));
  INV        m0426(.A(mai_mai_n268_), .Y(mai_mai_n455_));
  AN2        m0427(.A(e), .B(d), .Y(mai_mai_n456_));
  NA2        m0428(.A(mai_mai_n456_), .B(mai_mai_n455_), .Y(mai_mai_n457_));
  NO2        m0429(.A(mai_mai_n126_), .B(mai_mai_n41_), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n61_), .B(e), .Y(mai_mai_n459_));
  NA3        m0431(.A(mai_mai_n310_), .B(mai_mai_n255_), .C(mai_mai_n114_), .Y(mai_mai_n460_));
  NA2        m0432(.A(mai_mai_n460_), .B(mai_mai_n459_), .Y(mai_mai_n461_));
  AOI210     m0433(.A0(mai_mai_n461_), .A1(mai_mai_n457_), .B0(mai_mai_n454_), .Y(mai_mai_n462_));
  INV        m0434(.A(mai_mai_n200_), .Y(mai_mai_n463_));
  NOi21      m0435(.An(a), .B(b), .Y(mai_mai_n464_));
  NA3        m0436(.A(e), .B(d), .C(c), .Y(mai_mai_n465_));
  NAi21      m0437(.An(mai_mai_n465_), .B(mai_mai_n464_), .Y(mai_mai_n466_));
  NO2        m0438(.A(mai_mai_n411_), .B(mai_mai_n199_), .Y(mai_mai_n467_));
  NOi21      m0439(.An(mai_mai_n466_), .B(mai_mai_n467_), .Y(mai_mai_n468_));
  AOI210     m0440(.A0(mai_mai_n263_), .A1(mai_mai_n463_), .B0(mai_mai_n468_), .Y(mai_mai_n469_));
  NO4        m0441(.A(mai_mai_n182_), .B(mai_mai_n97_), .C(mai_mai_n54_), .D(b), .Y(mai_mai_n470_));
  NA2        m0442(.A(mai_mai_n373_), .B(mai_mai_n147_), .Y(mai_mai_n471_));
  OR2        m0443(.A(k), .B(j), .Y(mai_mai_n472_));
  NA2        m0444(.A(l), .B(k), .Y(mai_mai_n473_));
  NA3        m0445(.A(mai_mai_n473_), .B(mai_mai_n472_), .C(mai_mai_n214_), .Y(mai_mai_n474_));
  AOI210     m0446(.A0(mai_mai_n227_), .A1(mai_mai_n327_), .B0(mai_mai_n80_), .Y(mai_mai_n475_));
  NOi21      m0447(.An(mai_mai_n474_), .B(mai_mai_n475_), .Y(mai_mai_n476_));
  OR3        m0448(.A(mai_mai_n476_), .B(mai_mai_n138_), .C(mai_mai_n130_), .Y(mai_mai_n477_));
  NA2        m0449(.A(mai_mai_n273_), .B(mai_mai_n122_), .Y(mai_mai_n478_));
  NA2        m0450(.A(mai_mai_n386_), .B(mai_mai_n108_), .Y(mai_mai_n479_));
  NO4        m0451(.A(mai_mai_n479_), .B(mai_mai_n90_), .C(mai_mai_n107_), .D(e), .Y(mai_mai_n480_));
  NO3        m0452(.A(mai_mai_n411_), .B(mai_mai_n87_), .C(mai_mai_n126_), .Y(mai_mai_n481_));
  NO4        m0453(.A(mai_mai_n481_), .B(mai_mai_n480_), .C(mai_mai_n478_), .D(mai_mai_n311_), .Y(mai_mai_n482_));
  NA3        m0454(.A(mai_mai_n482_), .B(mai_mai_n477_), .C(mai_mai_n471_), .Y(mai_mai_n483_));
  NO4        m0455(.A(mai_mai_n483_), .B(mai_mai_n470_), .C(mai_mai_n469_), .D(mai_mai_n462_), .Y(mai_mai_n484_));
  NA2        m0456(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n485_));
  NOi21      m0457(.An(d), .B(e), .Y(mai_mai_n486_));
  NO2        m0458(.A(mai_mai_n182_), .B(mai_mai_n54_), .Y(mai_mai_n487_));
  NAi31      m0459(.An(j), .B(l), .C(i), .Y(mai_mai_n488_));
  OAI210     m0460(.A0(mai_mai_n488_), .A1(mai_mai_n127_), .B0(mai_mai_n97_), .Y(mai_mai_n489_));
  NA3        m0461(.A(mai_mai_n489_), .B(mai_mai_n487_), .C(mai_mai_n486_), .Y(mai_mai_n490_));
  NO3        m0462(.A(mai_mai_n387_), .B(mai_mai_n335_), .C(mai_mai_n196_), .Y(mai_mai_n491_));
  NO2        m0463(.A(mai_mai_n387_), .B(mai_mai_n363_), .Y(mai_mai_n492_));
  NO4        m0464(.A(mai_mai_n492_), .B(mai_mai_n491_), .C(mai_mai_n178_), .D(mai_mai_n295_), .Y(mai_mai_n493_));
  NA4        m0465(.A(mai_mai_n493_), .B(mai_mai_n490_), .C(mai_mai_n485_), .D(mai_mai_n236_), .Y(mai_mai_n494_));
  OAI210     m0466(.A0(mai_mai_n123_), .A1(mai_mai_n121_), .B0(n), .Y(mai_mai_n495_));
  NO2        m0467(.A(mai_mai_n495_), .B(mai_mai_n126_), .Y(mai_mai_n496_));
  BUFFER     m0468(.A(mai_mai_n238_), .Y(mai_mai_n497_));
  OA210      m0469(.A0(mai_mai_n497_), .A1(mai_mai_n496_), .B0(mai_mai_n187_), .Y(mai_mai_n498_));
  XO2        m0470(.A(i), .B(h), .Y(mai_mai_n499_));
  NA3        m0471(.A(mai_mai_n499_), .B(mai_mai_n154_), .C(n), .Y(mai_mai_n500_));
  NAi41      m0472(.An(mai_mai_n289_), .B(mai_mai_n500_), .C(mai_mai_n448_), .D(mai_mai_n375_), .Y(mai_mai_n501_));
  NOi32      m0473(.An(mai_mai_n501_), .Bn(mai_mai_n459_), .C(mai_mai_n265_), .Y(mai_mai_n502_));
  NAi31      m0474(.An(c), .B(f), .C(d), .Y(mai_mai_n503_));
  AOI210     m0475(.A0(mai_mai_n274_), .A1(mai_mai_n190_), .B0(mai_mai_n503_), .Y(mai_mai_n504_));
  NOi21      m0476(.An(mai_mai_n78_), .B(mai_mai_n504_), .Y(mai_mai_n505_));
  NA3        m0477(.A(mai_mai_n371_), .B(mai_mai_n93_), .C(mai_mai_n92_), .Y(mai_mai_n506_));
  NA2        m0478(.A(mai_mai_n221_), .B(mai_mai_n103_), .Y(mai_mai_n507_));
  AOI210     m0479(.A0(mai_mai_n507_), .A1(mai_mai_n174_), .B0(mai_mai_n503_), .Y(mai_mai_n508_));
  AOI210     m0480(.A0(mai_mai_n351_), .A1(mai_mai_n35_), .B0(mai_mai_n466_), .Y(mai_mai_n509_));
  NOi31      m0481(.An(mai_mai_n506_), .B(mai_mai_n509_), .C(mai_mai_n508_), .Y(mai_mai_n510_));
  NA3        m0482(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n511_), .B(mai_mai_n423_), .Y(mai_mai_n512_));
  NO2        m0484(.A(mai_mai_n512_), .B(mai_mai_n285_), .Y(mai_mai_n513_));
  NA3        m0485(.A(mai_mai_n513_), .B(mai_mai_n510_), .C(mai_mai_n505_), .Y(mai_mai_n514_));
  NO4        m0486(.A(mai_mai_n514_), .B(mai_mai_n502_), .C(mai_mai_n498_), .D(mai_mai_n494_), .Y(mai_mai_n515_));
  NA4        m0487(.A(mai_mai_n515_), .B(mai_mai_n484_), .C(mai_mai_n452_), .D(mai_mai_n418_), .Y(mai11));
  NO2        m0488(.A(mai_mai_n67_), .B(f), .Y(mai_mai_n517_));
  NA2        m0489(.A(j), .B(g), .Y(mai_mai_n518_));
  NAi31      m0490(.An(i), .B(m), .C(l), .Y(mai_mai_n519_));
  NA3        m0491(.A(m), .B(k), .C(j), .Y(mai_mai_n520_));
  OAI220     m0492(.A0(mai_mai_n520_), .A1(mai_mai_n126_), .B0(mai_mai_n519_), .B1(mai_mai_n518_), .Y(mai_mai_n521_));
  NOi32      m0493(.An(e), .Bn(b), .C(f), .Y(mai_mai_n522_));
  NA2        m0494(.A(mai_mai_n254_), .B(mai_mai_n108_), .Y(mai_mai_n523_));
  NA2        m0495(.A(mai_mai_n45_), .B(j), .Y(mai_mai_n524_));
  NAi31      m0496(.An(d), .B(e), .C(a), .Y(mai_mai_n525_));
  NO2        m0497(.A(mai_mai_n525_), .B(n), .Y(mai_mai_n526_));
  NAi41      m0498(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n527_));
  AN2        m0499(.A(mai_mai_n527_), .B(mai_mai_n362_), .Y(mai_mai_n528_));
  AOI210     m0500(.A0(mai_mai_n528_), .A1(mai_mai_n387_), .B0(mai_mai_n266_), .Y(mai_mai_n529_));
  NA2        m0501(.A(j), .B(i), .Y(mai_mai_n530_));
  NAi31      m0502(.An(n), .B(m), .C(k), .Y(mai_mai_n531_));
  NO3        m0503(.A(mai_mai_n531_), .B(mai_mai_n530_), .C(mai_mai_n107_), .Y(mai_mai_n532_));
  NO4        m0504(.A(n), .B(d), .C(mai_mai_n111_), .D(a), .Y(mai_mai_n533_));
  OR2        m0505(.A(n), .B(c), .Y(mai_mai_n534_));
  NO2        m0506(.A(mai_mai_n534_), .B(mai_mai_n143_), .Y(mai_mai_n535_));
  NO2        m0507(.A(mai_mai_n535_), .B(mai_mai_n533_), .Y(mai_mai_n536_));
  NOi32      m0508(.An(g), .Bn(f), .C(i), .Y(mai_mai_n537_));
  NA2        m0509(.A(mai_mai_n521_), .B(f), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n268_), .B(mai_mai_n47_), .Y(mai_mai_n539_));
  NO2        m0511(.A(mai_mai_n538_), .B(mai_mai_n536_), .Y(mai_mai_n540_));
  AOI210     m0512(.A0(mai_mai_n532_), .A1(mai_mai_n529_), .B0(mai_mai_n540_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n135_), .B(mai_mai_n34_), .Y(mai_mai_n542_));
  OAI220     m0514(.A0(mai_mai_n542_), .A1(m), .B0(mai_mai_n524_), .B1(mai_mai_n227_), .Y(mai_mai_n543_));
  NOi41      m0515(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n544_));
  NAi32      m0516(.An(e), .Bn(b), .C(c), .Y(mai_mai_n545_));
  OR2        m0517(.A(mai_mai_n545_), .B(mai_mai_n80_), .Y(mai_mai_n546_));
  AN2        m0518(.A(mai_mai_n328_), .B(mai_mai_n307_), .Y(mai_mai_n547_));
  NA2        m0519(.A(mai_mai_n547_), .B(mai_mai_n546_), .Y(mai_mai_n548_));
  OA210      m0520(.A0(mai_mai_n548_), .A1(mai_mai_n544_), .B0(mai_mai_n543_), .Y(mai_mai_n549_));
  OAI220     m0521(.A0(mai_mai_n389_), .A1(mai_mai_n388_), .B0(mai_mai_n519_), .B1(mai_mai_n518_), .Y(mai_mai_n550_));
  NO3        m0522(.A(mai_mai_n59_), .B(mai_mai_n47_), .C(mai_mai_n207_), .Y(mai_mai_n551_));
  NO2        m0523(.A(mai_mai_n224_), .B(mai_mai_n105_), .Y(mai_mai_n552_));
  OAI210     m0524(.A0(mai_mai_n551_), .A1(mai_mai_n390_), .B0(mai_mai_n552_), .Y(mai_mai_n553_));
  INV        m0525(.A(mai_mai_n553_), .Y(mai_mai_n554_));
  INV        m0526(.A(mai_mai_n413_), .Y(mai_mai_n555_));
  NA2        m0527(.A(mai_mai_n550_), .B(f), .Y(mai_mai_n556_));
  NAi32      m0528(.An(d), .Bn(a), .C(b), .Y(mai_mai_n557_));
  NO2        m0529(.A(mai_mai_n557_), .B(mai_mai_n47_), .Y(mai_mai_n558_));
  NA2        m0530(.A(h), .B(f), .Y(mai_mai_n559_));
  NO2        m0531(.A(mai_mai_n559_), .B(mai_mai_n90_), .Y(mai_mai_n560_));
  NO3        m0532(.A(mai_mai_n170_), .B(mai_mai_n167_), .C(g), .Y(mai_mai_n561_));
  AOI220     m0533(.A0(mai_mai_n561_), .A1(mai_mai_n56_), .B0(mai_mai_n560_), .B1(mai_mai_n558_), .Y(mai_mai_n562_));
  OAI210     m0534(.A0(mai_mai_n556_), .A1(mai_mai_n555_), .B0(mai_mai_n562_), .Y(mai_mai_n563_));
  AN3        m0535(.A(j), .B(h), .C(g), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n140_), .B(c), .Y(mai_mai_n565_));
  NA3        m0537(.A(mai_mai_n565_), .B(mai_mai_n564_), .C(mai_mai_n447_), .Y(mai_mai_n566_));
  NA3        m0538(.A(f), .B(d), .C(b), .Y(mai_mai_n567_));
  INV        m0539(.A(mai_mai_n566_), .Y(mai_mai_n568_));
  NO4        m0540(.A(mai_mai_n568_), .B(mai_mai_n563_), .C(mai_mai_n554_), .D(mai_mai_n549_), .Y(mai_mai_n569_));
  AN2        m0541(.A(mai_mai_n569_), .B(mai_mai_n541_), .Y(mai_mai_n570_));
  INV        m0542(.A(k), .Y(mai_mai_n571_));
  NA3        m0543(.A(l), .B(mai_mai_n571_), .C(i), .Y(mai_mai_n572_));
  INV        m0544(.A(mai_mai_n572_), .Y(mai_mai_n573_));
  NA4        m0545(.A(mai_mai_n386_), .B(mai_mai_n405_), .C(mai_mai_n175_), .D(mai_mai_n108_), .Y(mai_mai_n574_));
  NAi32      m0546(.An(h), .Bn(f), .C(g), .Y(mai_mai_n575_));
  NAi41      m0547(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n576_));
  OAI210     m0548(.A0(mai_mai_n525_), .A1(n), .B0(mai_mai_n576_), .Y(mai_mai_n577_));
  NA2        m0549(.A(mai_mai_n577_), .B(m), .Y(mai_mai_n578_));
  NAi31      m0550(.An(h), .B(g), .C(f), .Y(mai_mai_n579_));
  NA4        m0551(.A(mai_mai_n405_), .B(mai_mai_n116_), .C(mai_mai_n108_), .D(e), .Y(mai_mai_n580_));
  OA210      m0552(.A0(mai_mai_n578_), .A1(mai_mai_n575_), .B0(mai_mai_n580_), .Y(mai_mai_n581_));
  NA2        m0553(.A(mai_mai_n581_), .B(mai_mai_n574_), .Y(mai_mai_n582_));
  NAi31      m0554(.An(f), .B(h), .C(g), .Y(mai_mai_n583_));
  NO4        m0555(.A(mai_mai_n300_), .B(mai_mai_n583_), .C(mai_mai_n67_), .D(mai_mai_n69_), .Y(mai_mai_n584_));
  NOi32      m0556(.An(b), .Bn(a), .C(c), .Y(mai_mai_n585_));
  NOi32      m0557(.An(d), .Bn(a), .C(e), .Y(mai_mai_n586_));
  NO2        m0558(.A(n), .B(c), .Y(mai_mai_n587_));
  NA3        m0559(.A(mai_mai_n587_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n588_));
  NAi32      m0560(.An(n), .Bn(f), .C(m), .Y(mai_mai_n589_));
  NOi32      m0561(.An(e), .Bn(a), .C(d), .Y(mai_mai_n590_));
  AOI210     m0562(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n590_), .Y(mai_mai_n591_));
  AOI210     m0563(.A0(mai_mai_n591_), .A1(mai_mai_n206_), .B0(mai_mai_n542_), .Y(mai_mai_n592_));
  AOI210     m0564(.A0(mai_mai_n592_), .A1(mai_mai_n1493_), .B0(mai_mai_n584_), .Y(mai_mai_n593_));
  OAI210     m0565(.A0(mai_mai_n243_), .A1(mai_mai_n83_), .B0(mai_mai_n593_), .Y(mai_mai_n594_));
  AOI210     m0566(.A0(mai_mai_n582_), .A1(mai_mai_n573_), .B0(mai_mai_n594_), .Y(mai_mai_n595_));
  NO3        m0567(.A(mai_mai_n305_), .B(mai_mai_n58_), .C(n), .Y(mai_mai_n596_));
  NA3        m0568(.A(mai_mai_n503_), .B(mai_mai_n165_), .C(mai_mai_n164_), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n449_), .B(mai_mai_n224_), .Y(mai_mai_n598_));
  OR2        m0570(.A(mai_mai_n598_), .B(mai_mai_n597_), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n70_), .B(mai_mai_n108_), .Y(mai_mai_n600_));
  NO2        m0572(.A(mai_mai_n600_), .B(mai_mai_n44_), .Y(mai_mai_n601_));
  AOI220     m0573(.A0(mai_mai_n601_), .A1(mai_mai_n529_), .B0(mai_mai_n599_), .B1(mai_mai_n596_), .Y(mai_mai_n602_));
  NO2        m0574(.A(mai_mai_n602_), .B(mai_mai_n83_), .Y(mai_mai_n603_));
  NA3        m0575(.A(mai_mai_n544_), .B(mai_mai_n330_), .C(mai_mai_n45_), .Y(mai_mai_n604_));
  NOi32      m0576(.An(e), .Bn(c), .C(f), .Y(mai_mai_n605_));
  NOi21      m0577(.An(f), .B(g), .Y(mai_mai_n606_));
  NO2        m0578(.A(mai_mai_n606_), .B(mai_mai_n204_), .Y(mai_mai_n607_));
  AOI220     m0579(.A0(mai_mai_n607_), .A1(mai_mai_n383_), .B0(mai_mai_n605_), .B1(mai_mai_n169_), .Y(mai_mai_n608_));
  NA3        m0580(.A(mai_mai_n608_), .B(mai_mai_n604_), .C(mai_mai_n172_), .Y(mai_mai_n609_));
  AOI210     m0581(.A0(mai_mai_n528_), .A1(mai_mai_n387_), .B0(mai_mai_n290_), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n610_), .B(mai_mai_n258_), .Y(mai_mai_n611_));
  NAi21      m0583(.An(k), .B(h), .Y(mai_mai_n612_));
  NO2        m0584(.A(mai_mai_n612_), .B(mai_mai_n256_), .Y(mai_mai_n613_));
  NOi31      m0585(.An(m), .B(n), .C(k), .Y(mai_mai_n614_));
  NA2        m0586(.A(j), .B(mai_mai_n614_), .Y(mai_mai_n615_));
  AOI210     m0587(.A0(mai_mai_n387_), .A1(mai_mai_n362_), .B0(mai_mai_n290_), .Y(mai_mai_n616_));
  NAi21      m0588(.An(mai_mai_n615_), .B(mai_mai_n616_), .Y(mai_mai_n617_));
  NA2        m0589(.A(mai_mai_n617_), .B(mai_mai_n611_), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n103_), .B(mai_mai_n36_), .Y(mai_mai_n619_));
  NO2        m0591(.A(k), .B(mai_mai_n207_), .Y(mai_mai_n620_));
  INV        m0592(.A(mai_mai_n353_), .Y(mai_mai_n621_));
  NO2        m0593(.A(mai_mai_n621_), .B(n), .Y(mai_mai_n622_));
  NAi31      m0594(.An(mai_mai_n619_), .B(mai_mai_n622_), .C(mai_mai_n620_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n524_), .B(mai_mai_n170_), .Y(mai_mai_n624_));
  NA3        m0596(.A(mai_mai_n545_), .B(mai_mai_n265_), .C(mai_mai_n139_), .Y(mai_mai_n625_));
  NA2        m0597(.A(mai_mai_n499_), .B(mai_mai_n154_), .Y(mai_mai_n626_));
  NO3        m0598(.A(mai_mai_n384_), .B(mai_mai_n626_), .C(mai_mai_n83_), .Y(mai_mai_n627_));
  AOI210     m0599(.A0(mai_mai_n625_), .A1(mai_mai_n624_), .B0(mai_mai_n627_), .Y(mai_mai_n628_));
  AN3        m0600(.A(f), .B(d), .C(b), .Y(mai_mai_n629_));
  OAI210     m0601(.A0(mai_mai_n629_), .A1(mai_mai_n125_), .B0(n), .Y(mai_mai_n630_));
  NA3        m0602(.A(mai_mai_n499_), .B(mai_mai_n154_), .C(mai_mai_n207_), .Y(mai_mai_n631_));
  AOI210     m0603(.A0(mai_mai_n630_), .A1(mai_mai_n226_), .B0(mai_mai_n631_), .Y(mai_mai_n632_));
  NAi31      m0604(.An(m), .B(n), .C(k), .Y(mai_mai_n633_));
  OR2        m0605(.A(mai_mai_n130_), .B(mai_mai_n58_), .Y(mai_mai_n634_));
  OAI210     m0606(.A0(mai_mai_n634_), .A1(mai_mai_n633_), .B0(mai_mai_n245_), .Y(mai_mai_n635_));
  OAI210     m0607(.A0(mai_mai_n635_), .A1(mai_mai_n632_), .B0(j), .Y(mai_mai_n636_));
  NA3        m0608(.A(mai_mai_n636_), .B(mai_mai_n628_), .C(mai_mai_n623_), .Y(mai_mai_n637_));
  NO4        m0609(.A(mai_mai_n637_), .B(mai_mai_n618_), .C(mai_mai_n609_), .D(mai_mai_n603_), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n371_), .B(mai_mai_n157_), .Y(mai_mai_n639_));
  NAi31      m0611(.An(g), .B(h), .C(f), .Y(mai_mai_n640_));
  OA210      m0612(.A0(mai_mai_n525_), .A1(n), .B0(mai_mai_n576_), .Y(mai_mai_n641_));
  NO2        m0613(.A(mai_mai_n641_), .B(mai_mai_n86_), .Y(mai_mai_n642_));
  INV        m0614(.A(mai_mai_n642_), .Y(mai_mai_n643_));
  AOI210     m0615(.A0(mai_mai_n643_), .A1(mai_mai_n639_), .B0(mai_mai_n520_), .Y(mai_mai_n644_));
  NO3        m0616(.A(g), .B(mai_mai_n206_), .C(mai_mai_n54_), .Y(mai_mai_n645_));
  NAi21      m0617(.An(h), .B(j), .Y(mai_mai_n646_));
  NA2        m0618(.A(mai_mai_n383_), .B(mai_mai_n645_), .Y(mai_mai_n647_));
  OR2        m0619(.A(mai_mai_n67_), .B(mai_mai_n69_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n517_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n649_));
  AN2        m0621(.A(h), .B(f), .Y(mai_mai_n650_));
  NA2        m0622(.A(mai_mai_n650_), .B(mai_mai_n37_), .Y(mai_mai_n651_));
  NA2        m0623(.A(mai_mai_n95_), .B(mai_mai_n45_), .Y(mai_mai_n652_));
  OAI220     m0624(.A0(mai_mai_n652_), .A1(mai_mai_n321_), .B0(mai_mai_n651_), .B1(mai_mai_n454_), .Y(mai_mai_n653_));
  AOI210     m0625(.A0(mai_mai_n557_), .A1(mai_mai_n412_), .B0(mai_mai_n47_), .Y(mai_mai_n654_));
  OAI220     m0626(.A0(mai_mai_n579_), .A1(mai_mai_n572_), .B0(mai_mai_n315_), .B1(mai_mai_n518_), .Y(mai_mai_n655_));
  AOI210     m0627(.A0(mai_mai_n655_), .A1(mai_mai_n654_), .B0(mai_mai_n653_), .Y(mai_mai_n656_));
  NA3        m0628(.A(mai_mai_n656_), .B(mai_mai_n649_), .C(mai_mai_n647_), .Y(mai_mai_n657_));
  NO2        m0629(.A(mai_mai_n247_), .B(f), .Y(mai_mai_n658_));
  NO2        m0630(.A(mai_mai_n606_), .B(mai_mai_n58_), .Y(mai_mai_n659_));
  NO3        m0631(.A(mai_mai_n659_), .B(mai_mai_n658_), .C(mai_mai_n34_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n318_), .B(mai_mai_n135_), .Y(mai_mai_n661_));
  NA2        m0633(.A(mai_mai_n127_), .B(mai_mai_n47_), .Y(mai_mai_n662_));
  NA2        m0634(.A(mai_mai_n662_), .B(mai_mai_n522_), .Y(mai_mai_n663_));
  OA220      m0635(.A0(mai_mai_n663_), .A1(mai_mai_n542_), .B0(mai_mai_n351_), .B1(mai_mai_n106_), .Y(mai_mai_n664_));
  OAI210     m0636(.A0(mai_mai_n661_), .A1(mai_mai_n660_), .B0(mai_mai_n664_), .Y(mai_mai_n665_));
  NO3        m0637(.A(mai_mai_n393_), .B(mai_mai_n187_), .C(mai_mai_n186_), .Y(mai_mai_n666_));
  NA2        m0638(.A(mai_mai_n666_), .B(mai_mai_n224_), .Y(mai_mai_n667_));
  NA3        m0639(.A(mai_mai_n667_), .B(mai_mai_n249_), .C(j), .Y(mai_mai_n668_));
  NO3        m0640(.A(mai_mai_n449_), .B(mai_mai_n167_), .C(i), .Y(mai_mai_n669_));
  NA2        m0641(.A(mai_mai_n453_), .B(mai_mai_n80_), .Y(mai_mai_n670_));
  NO4        m0642(.A(mai_mai_n520_), .B(mai_mai_n670_), .C(mai_mai_n126_), .D(mai_mai_n206_), .Y(mai_mai_n671_));
  INV        m0643(.A(mai_mai_n671_), .Y(mai_mai_n672_));
  NA4        m0644(.A(mai_mai_n672_), .B(mai_mai_n668_), .C(mai_mai_n506_), .D(mai_mai_n391_), .Y(mai_mai_n673_));
  NO4        m0645(.A(mai_mai_n673_), .B(mai_mai_n665_), .C(mai_mai_n657_), .D(mai_mai_n644_), .Y(mai_mai_n674_));
  NA4        m0646(.A(mai_mai_n674_), .B(mai_mai_n638_), .C(mai_mai_n595_), .D(mai_mai_n570_), .Y(mai08));
  NO2        m0647(.A(k), .B(h), .Y(mai_mai_n676_));
  AO210      m0648(.A0(mai_mai_n247_), .A1(mai_mai_n437_), .B0(mai_mai_n676_), .Y(mai_mai_n677_));
  NO2        m0649(.A(mai_mai_n677_), .B(mai_mai_n288_), .Y(mai_mai_n678_));
  NA2        m0650(.A(mai_mai_n605_), .B(mai_mai_n80_), .Y(mai_mai_n679_));
  NA2        m0651(.A(mai_mai_n679_), .B(mai_mai_n449_), .Y(mai_mai_n680_));
  AOI210     m0652(.A0(mai_mai_n680_), .A1(mai_mai_n678_), .B0(mai_mai_n481_), .Y(mai_mai_n681_));
  NA2        m0653(.A(mai_mai_n80_), .B(mai_mai_n105_), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n682_), .B(mai_mai_n55_), .Y(mai_mai_n683_));
  NA2        m0655(.A(mai_mai_n567_), .B(mai_mai_n226_), .Y(mai_mai_n684_));
  NA2        m0656(.A(mai_mai_n684_), .B(mai_mai_n338_), .Y(mai_mai_n685_));
  AOI210     m0657(.A0(mai_mai_n567_), .A1(mai_mai_n150_), .B0(mai_mai_n80_), .Y(mai_mai_n686_));
  NA4        m0658(.A(mai_mai_n209_), .B(mai_mai_n135_), .C(mai_mai_n44_), .D(h), .Y(mai_mai_n687_));
  AN2        m0659(.A(l), .B(k), .Y(mai_mai_n688_));
  NA3        m0660(.A(mai_mai_n685_), .B(mai_mai_n681_), .C(mai_mai_n340_), .Y(mai_mai_n689_));
  NO4        m0661(.A(mai_mai_n167_), .B(mai_mai_n382_), .C(mai_mai_n107_), .D(g), .Y(mai_mai_n690_));
  AOI210     m0662(.A0(mai_mai_n690_), .A1(mai_mai_n684_), .B0(mai_mai_n512_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n607_), .B(mai_mai_n337_), .Y(mai_mai_n692_));
  NA2        m0664(.A(mai_mai_n692_), .B(mai_mai_n691_), .Y(mai_mai_n693_));
  NO2        m0665(.A(mai_mai_n528_), .B(mai_mai_n35_), .Y(mai_mai_n694_));
  OAI210     m0666(.A0(mai_mai_n545_), .A1(mai_mai_n46_), .B0(mai_mai_n634_), .Y(mai_mai_n695_));
  NO2        m0667(.A(mai_mai_n473_), .B(mai_mai_n127_), .Y(mai_mai_n696_));
  AOI210     m0668(.A0(mai_mai_n696_), .A1(mai_mai_n695_), .B0(mai_mai_n694_), .Y(mai_mai_n697_));
  NO3        m0669(.A(mai_mai_n305_), .B(mai_mai_n126_), .C(mai_mai_n41_), .Y(mai_mai_n698_));
  BUFFER     m0670(.A(mai_mai_n698_), .Y(mai_mai_n699_));
  NA2        m0671(.A(mai_mai_n677_), .B(mai_mai_n131_), .Y(mai_mai_n700_));
  AOI220     m0672(.A0(mai_mai_n700_), .A1(mai_mai_n392_), .B0(mai_mai_n699_), .B1(mai_mai_n72_), .Y(mai_mai_n701_));
  OAI210     m0673(.A0(mai_mai_n697_), .A1(mai_mai_n83_), .B0(mai_mai_n701_), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n353_), .B(mai_mai_n43_), .Y(mai_mai_n703_));
  NA3        m0675(.A(mai_mai_n667_), .B(mai_mai_n323_), .C(mai_mai_n374_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n688_), .B(mai_mai_n214_), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n705_), .B(mai_mai_n317_), .Y(mai_mai_n706_));
  AOI210     m0678(.A0(mai_mai_n706_), .A1(mai_mai_n658_), .B0(mai_mai_n480_), .Y(mai_mai_n707_));
  NA3        m0679(.A(m), .B(l), .C(k), .Y(mai_mai_n708_));
  NO2        m0680(.A(mai_mai_n527_), .B(mai_mai_n266_), .Y(mai_mai_n709_));
  NOi21      m0681(.An(mai_mai_n709_), .B(mai_mai_n523_), .Y(mai_mai_n710_));
  NA4        m0682(.A(mai_mai_n108_), .B(l), .C(k), .D(mai_mai_n83_), .Y(mai_mai_n711_));
  NA3        m0683(.A(mai_mai_n116_), .B(mai_mai_n401_), .C(i), .Y(mai_mai_n712_));
  NO2        m0684(.A(mai_mai_n712_), .B(mai_mai_n711_), .Y(mai_mai_n713_));
  NO2        m0685(.A(mai_mai_n713_), .B(mai_mai_n710_), .Y(mai_mai_n714_));
  NA4        m0686(.A(mai_mai_n714_), .B(mai_mai_n707_), .C(mai_mai_n704_), .D(mai_mai_n703_), .Y(mai_mai_n715_));
  NO4        m0687(.A(mai_mai_n715_), .B(mai_mai_n702_), .C(mai_mai_n693_), .D(mai_mai_n689_), .Y(mai_mai_n716_));
  NA2        m0688(.A(mai_mai_n607_), .B(mai_mai_n383_), .Y(mai_mai_n717_));
  NO3        m0689(.A(mai_mai_n387_), .B(mai_mai_n518_), .C(h), .Y(mai_mai_n718_));
  AOI210     m0690(.A0(mai_mai_n718_), .A1(mai_mai_n108_), .B0(mai_mai_n492_), .Y(mai_mai_n719_));
  NA3        m0691(.A(mai_mai_n719_), .B(mai_mai_n717_), .C(mai_mai_n246_), .Y(mai_mai_n720_));
  NA2        m0692(.A(mai_mai_n688_), .B(mai_mai_n69_), .Y(mai_mai_n721_));
  NO4        m0693(.A(mai_mai_n666_), .B(mai_mai_n167_), .C(n), .D(i), .Y(mai_mai_n722_));
  NOi21      m0694(.An(h), .B(j), .Y(mai_mai_n723_));
  NA2        m0695(.A(mai_mai_n723_), .B(f), .Y(mai_mai_n724_));
  NO2        m0696(.A(mai_mai_n724_), .B(mai_mai_n240_), .Y(mai_mai_n725_));
  NO3        m0697(.A(mai_mai_n725_), .B(mai_mai_n722_), .C(mai_mai_n669_), .Y(mai_mai_n726_));
  NO2        m0698(.A(mai_mai_n726_), .B(mai_mai_n721_), .Y(mai_mai_n727_));
  AOI210     m0699(.A0(mai_mai_n720_), .A1(l), .B0(mai_mai_n727_), .Y(mai_mai_n728_));
  NO2        m0700(.A(j), .B(i), .Y(mai_mai_n729_));
  NA3        m0701(.A(mai_mai_n729_), .B(mai_mai_n76_), .C(l), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n729_), .B(mai_mai_n33_), .Y(mai_mai_n731_));
  OR2        m0703(.A(mai_mai_n730_), .B(mai_mai_n578_), .Y(mai_mai_n732_));
  NO3        m0704(.A(mai_mai_n145_), .B(mai_mai_n47_), .C(mai_mai_n105_), .Y(mai_mai_n733_));
  NO3        m0705(.A(mai_mai_n473_), .B(mai_mai_n424_), .C(j), .Y(mai_mai_n734_));
  NA2        m0706(.A(mai_mai_n733_), .B(mai_mai_n734_), .Y(mai_mai_n735_));
  INV        m0707(.A(mai_mai_n735_), .Y(mai_mai_n736_));
  NA2        m0708(.A(k), .B(j), .Y(mai_mai_n737_));
  NO3        m0709(.A(mai_mai_n288_), .B(mai_mai_n737_), .C(mai_mai_n40_), .Y(mai_mai_n738_));
  AOI210     m0710(.A0(mai_mai_n522_), .A1(n), .B0(mai_mai_n544_), .Y(mai_mai_n739_));
  NA2        m0711(.A(mai_mai_n739_), .B(mai_mai_n547_), .Y(mai_mai_n740_));
  AN3        m0712(.A(mai_mai_n740_), .B(mai_mai_n738_), .C(mai_mai_n94_), .Y(mai_mai_n741_));
  NO3        m0713(.A(mai_mai_n167_), .B(mai_mai_n382_), .C(mai_mai_n107_), .Y(mai_mai_n742_));
  AOI220     m0714(.A0(mai_mai_n742_), .A1(mai_mai_n241_), .B0(mai_mai_n598_), .B1(mai_mai_n297_), .Y(mai_mai_n743_));
  NAi31      m0715(.An(mai_mai_n591_), .B(mai_mai_n88_), .C(mai_mai_n80_), .Y(mai_mai_n744_));
  NA2        m0716(.A(mai_mai_n744_), .B(mai_mai_n743_), .Y(mai_mai_n745_));
  NO2        m0717(.A(mai_mai_n288_), .B(mai_mai_n131_), .Y(mai_mai_n746_));
  AOI220     m0718(.A0(mai_mai_n746_), .A1(mai_mai_n607_), .B0(mai_mai_n698_), .B1(mai_mai_n686_), .Y(mai_mai_n747_));
  NO2        m0719(.A(mai_mai_n708_), .B(mai_mai_n86_), .Y(mai_mai_n748_));
  NA2        m0720(.A(mai_mai_n748_), .B(mai_mai_n577_), .Y(mai_mai_n749_));
  NO2        m0721(.A(mai_mai_n579_), .B(mai_mai_n112_), .Y(mai_mai_n750_));
  OAI210     m0722(.A0(mai_mai_n750_), .A1(mai_mai_n734_), .B0(mai_mai_n654_), .Y(mai_mai_n751_));
  NA3        m0723(.A(mai_mai_n751_), .B(mai_mai_n749_), .C(mai_mai_n747_), .Y(mai_mai_n752_));
  OR4        m0724(.A(mai_mai_n752_), .B(mai_mai_n745_), .C(mai_mai_n741_), .D(mai_mai_n736_), .Y(mai_mai_n753_));
  NA3        m0725(.A(mai_mai_n739_), .B(mai_mai_n547_), .C(mai_mai_n546_), .Y(mai_mai_n754_));
  NA4        m0726(.A(mai_mai_n754_), .B(mai_mai_n209_), .C(mai_mai_n437_), .D(mai_mai_n34_), .Y(mai_mai_n755_));
  NO4        m0727(.A(mai_mai_n473_), .B(mai_mai_n419_), .C(j), .D(f), .Y(mai_mai_n756_));
  OAI220     m0728(.A0(mai_mai_n687_), .A1(mai_mai_n679_), .B0(mai_mai_n321_), .B1(mai_mai_n38_), .Y(mai_mai_n757_));
  AOI210     m0729(.A0(mai_mai_n756_), .A1(mai_mai_n253_), .B0(mai_mai_n757_), .Y(mai_mai_n758_));
  NA3        m0730(.A(mai_mai_n537_), .B(mai_mai_n281_), .C(h), .Y(mai_mai_n759_));
  NOi21      m0731(.An(mai_mai_n654_), .B(mai_mai_n759_), .Y(mai_mai_n760_));
  NO2        m0732(.A(mai_mai_n730_), .B(mai_mai_n648_), .Y(mai_mai_n761_));
  INV        m0733(.A(mai_mai_n761_), .Y(mai_mai_n762_));
  NAi41      m0734(.An(mai_mai_n760_), .B(mai_mai_n762_), .C(mai_mai_n758_), .D(mai_mai_n755_), .Y(mai_mai_n763_));
  OR2        m0735(.A(mai_mai_n748_), .B(mai_mai_n91_), .Y(mai_mai_n764_));
  NA2        m0736(.A(mai_mai_n764_), .B(mai_mai_n231_), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n641_), .B(mai_mai_n69_), .Y(mai_mai_n766_));
  AOI210     m0738(.A0(mai_mai_n756_), .A1(mai_mai_n766_), .B0(mai_mai_n325_), .Y(mai_mai_n767_));
  OAI210     m0739(.A0(mai_mai_n708_), .A1(mai_mai_n640_), .B0(mai_mai_n511_), .Y(mai_mai_n768_));
  NA3        m0740(.A(mai_mai_n244_), .B(mai_mai_n57_), .C(b), .Y(mai_mai_n769_));
  AOI220     m0741(.A0(mai_mai_n587_), .A1(mai_mai_n29_), .B0(mai_mai_n453_), .B1(mai_mai_n80_), .Y(mai_mai_n770_));
  NA2        m0742(.A(mai_mai_n770_), .B(mai_mai_n769_), .Y(mai_mai_n771_));
  NO2        m0743(.A(mai_mai_n759_), .B(mai_mai_n479_), .Y(mai_mai_n772_));
  AOI210     m0744(.A0(mai_mai_n771_), .A1(mai_mai_n768_), .B0(mai_mai_n772_), .Y(mai_mai_n773_));
  NA3        m0745(.A(mai_mai_n773_), .B(mai_mai_n767_), .C(mai_mai_n765_), .Y(mai_mai_n774_));
  NOi41      m0746(.An(mai_mai_n732_), .B(mai_mai_n774_), .C(mai_mai_n763_), .D(mai_mai_n753_), .Y(mai_mai_n775_));
  NO3        m0747(.A(mai_mai_n331_), .B(mai_mai_n290_), .C(mai_mai_n107_), .Y(mai_mai_n776_));
  NA2        m0748(.A(mai_mai_n776_), .B(mai_mai_n740_), .Y(mai_mai_n777_));
  NA2        m0749(.A(mai_mai_n45_), .B(mai_mai_n54_), .Y(mai_mai_n778_));
  NO3        m0750(.A(mai_mai_n778_), .B(mai_mai_n731_), .C(mai_mai_n270_), .Y(mai_mai_n779_));
  INV        m0751(.A(mai_mai_n779_), .Y(mai_mai_n780_));
  NA3        m0752(.A(mai_mai_n780_), .B(mai_mai_n777_), .C(mai_mai_n394_), .Y(mai_mai_n781_));
  OR2        m0753(.A(mai_mai_n640_), .B(mai_mai_n87_), .Y(mai_mai_n782_));
  NOi31      m0754(.An(b), .B(d), .C(a), .Y(mai_mai_n783_));
  NO2        m0755(.A(mai_mai_n783_), .B(mai_mai_n586_), .Y(mai_mai_n784_));
  NO2        m0756(.A(mai_mai_n784_), .B(n), .Y(mai_mai_n785_));
  NO2        m0757(.A(mai_mai_n545_), .B(mai_mai_n80_), .Y(mai_mai_n786_));
  NA2        m0758(.A(mai_mai_n776_), .B(mai_mai_n786_), .Y(mai_mai_n787_));
  OAI210     m0759(.A0(mai_mai_n687_), .A1(mai_mai_n384_), .B0(mai_mai_n787_), .Y(mai_mai_n788_));
  NO2        m0760(.A(mai_mai_n666_), .B(n), .Y(mai_mai_n789_));
  AOI220     m0761(.A0(mai_mai_n746_), .A1(mai_mai_n645_), .B0(mai_mai_n789_), .B1(mai_mai_n678_), .Y(mai_mai_n790_));
  NO2        m0762(.A(mai_mai_n312_), .B(mai_mai_n230_), .Y(mai_mai_n791_));
  OAI210     m0763(.A0(mai_mai_n91_), .A1(mai_mai_n88_), .B0(mai_mai_n791_), .Y(mai_mai_n792_));
  NA2        m0764(.A(mai_mai_n116_), .B(mai_mai_n80_), .Y(mai_mai_n793_));
  AOI210     m0765(.A0(mai_mai_n409_), .A1(mai_mai_n404_), .B0(mai_mai_n793_), .Y(mai_mai_n794_));
  NAi21      m0766(.An(mai_mai_n794_), .B(mai_mai_n792_), .Y(mai_mai_n795_));
  NA2        m0767(.A(mai_mai_n706_), .B(mai_mai_n34_), .Y(mai_mai_n796_));
  NAi21      m0768(.An(mai_mai_n711_), .B(mai_mai_n420_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n266_), .B(i), .Y(mai_mai_n798_));
  NA2        m0770(.A(mai_mai_n690_), .B(mai_mai_n339_), .Y(mai_mai_n799_));
  AN2        m0771(.A(mai_mai_n799_), .B(mai_mai_n797_), .Y(mai_mai_n800_));
  NAi41      m0772(.An(mai_mai_n795_), .B(mai_mai_n800_), .C(mai_mai_n796_), .D(mai_mai_n790_), .Y(mai_mai_n801_));
  NO3        m0773(.A(mai_mai_n801_), .B(mai_mai_n788_), .C(mai_mai_n781_), .Y(mai_mai_n802_));
  NA4        m0774(.A(mai_mai_n802_), .B(mai_mai_n775_), .C(mai_mai_n728_), .D(mai_mai_n716_), .Y(mai09));
  INV        m0775(.A(mai_mai_n117_), .Y(mai_mai_n804_));
  NA2        m0776(.A(f), .B(e), .Y(mai_mai_n805_));
  NO2        m0777(.A(mai_mai_n219_), .B(mai_mai_n107_), .Y(mai_mai_n806_));
  NA2        m0778(.A(mai_mai_n806_), .B(g), .Y(mai_mai_n807_));
  NA3        m0779(.A(mai_mai_n300_), .B(mai_mai_n255_), .C(mai_mai_n114_), .Y(mai_mai_n808_));
  AOI210     m0780(.A0(mai_mai_n808_), .A1(g), .B0(mai_mai_n458_), .Y(mai_mai_n809_));
  AOI210     m0781(.A0(mai_mai_n809_), .A1(mai_mai_n807_), .B0(mai_mai_n805_), .Y(mai_mai_n810_));
  NA2        m0782(.A(mai_mai_n430_), .B(e), .Y(mai_mai_n811_));
  NO2        m0783(.A(mai_mai_n811_), .B(mai_mai_n503_), .Y(mai_mai_n812_));
  AOI210     m0784(.A0(mai_mai_n810_), .A1(mai_mai_n804_), .B0(mai_mai_n812_), .Y(mai_mai_n813_));
  NO2        m0785(.A(mai_mai_n199_), .B(mai_mai_n206_), .Y(mai_mai_n814_));
  NA3        m0786(.A(m), .B(l), .C(i), .Y(mai_mai_n815_));
  OAI220     m0787(.A0(mai_mai_n579_), .A1(mai_mai_n815_), .B0(mai_mai_n344_), .B1(mai_mai_n519_), .Y(mai_mai_n816_));
  NAi21      m0788(.An(mai_mai_n816_), .B(mai_mai_n425_), .Y(mai_mai_n817_));
  OR2        m0789(.A(mai_mai_n817_), .B(mai_mai_n814_), .Y(mai_mai_n818_));
  NA3        m0790(.A(mai_mai_n782_), .B(mai_mai_n556_), .C(mai_mai_n511_), .Y(mai_mai_n819_));
  OA210      m0791(.A0(mai_mai_n819_), .A1(mai_mai_n818_), .B0(mai_mai_n785_), .Y(mai_mai_n820_));
  INV        m0792(.A(mai_mai_n328_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n123_), .B(mai_mai_n121_), .Y(mai_mai_n822_));
  NOi31      m0794(.An(k), .B(m), .C(l), .Y(mai_mai_n823_));
  NO2        m0795(.A(mai_mai_n330_), .B(mai_mai_n823_), .Y(mai_mai_n824_));
  AOI210     m0796(.A0(mai_mai_n824_), .A1(mai_mai_n822_), .B0(mai_mai_n583_), .Y(mai_mai_n825_));
  NA2        m0797(.A(mai_mai_n769_), .B(mai_mai_n321_), .Y(mai_mai_n826_));
  NA2        m0798(.A(mai_mai_n332_), .B(mai_mai_n334_), .Y(mai_mai_n827_));
  OAI210     m0799(.A0(mai_mai_n199_), .A1(mai_mai_n206_), .B0(mai_mai_n827_), .Y(mai_mai_n828_));
  AOI220     m0800(.A0(mai_mai_n828_), .A1(mai_mai_n826_), .B0(mai_mai_n825_), .B1(mai_mai_n821_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n161_), .B(mai_mai_n109_), .Y(mai_mai_n830_));
  NA3        m0802(.A(mai_mai_n830_), .B(mai_mai_n677_), .C(mai_mai_n131_), .Y(mai_mai_n831_));
  NA3        m0803(.A(mai_mai_n831_), .B(mai_mai_n184_), .C(mai_mai_n31_), .Y(mai_mai_n832_));
  NA4        m0804(.A(mai_mai_n832_), .B(mai_mai_n829_), .C(mai_mai_n608_), .D(mai_mai_n78_), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n575_), .B(mai_mai_n488_), .Y(mai_mai_n834_));
  NA2        m0806(.A(mai_mai_n834_), .B(mai_mai_n184_), .Y(mai_mai_n835_));
  NOi21      m0807(.An(f), .B(d), .Y(mai_mai_n836_));
  NA2        m0808(.A(mai_mai_n836_), .B(m), .Y(mai_mai_n837_));
  NO2        m0809(.A(mai_mai_n837_), .B(mai_mai_n50_), .Y(mai_mai_n838_));
  NOi32      m0810(.An(g), .Bn(f), .C(d), .Y(mai_mai_n839_));
  NA4        m0811(.A(mai_mai_n839_), .B(mai_mai_n587_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n840_));
  NOi21      m0812(.An(mai_mai_n301_), .B(mai_mai_n840_), .Y(mai_mai_n841_));
  AOI210     m0813(.A0(mai_mai_n838_), .A1(mai_mai_n535_), .B0(mai_mai_n841_), .Y(mai_mai_n842_));
  NA3        m0814(.A(mai_mai_n300_), .B(mai_mai_n255_), .C(mai_mai_n114_), .Y(mai_mai_n843_));
  AN2        m0815(.A(f), .B(d), .Y(mai_mai_n844_));
  NA3        m0816(.A(mai_mai_n464_), .B(mai_mai_n844_), .C(mai_mai_n80_), .Y(mai_mai_n845_));
  NO3        m0817(.A(mai_mai_n845_), .B(mai_mai_n69_), .C(mai_mai_n207_), .Y(mai_mai_n846_));
  NO2        m0818(.A(mai_mai_n278_), .B(mai_mai_n54_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n843_), .B(mai_mai_n846_), .Y(mai_mai_n848_));
  NAi41      m0820(.An(mai_mai_n478_), .B(mai_mai_n848_), .C(mai_mai_n842_), .D(mai_mai_n835_), .Y(mai_mai_n849_));
  NO4        m0821(.A(mai_mai_n606_), .B(mai_mai_n127_), .C(mai_mai_n317_), .D(mai_mai_n146_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n633_), .B(mai_mai_n317_), .Y(mai_mai_n851_));
  AN2        m0823(.A(mai_mai_n851_), .B(mai_mai_n658_), .Y(mai_mai_n852_));
  NO2        m0824(.A(mai_mai_n852_), .B(mai_mai_n850_), .Y(mai_mai_n853_));
  NA2        m0825(.A(mai_mai_n586_), .B(mai_mai_n80_), .Y(mai_mai_n854_));
  NA3        m0826(.A(mai_mai_n154_), .B(mai_mai_n103_), .C(mai_mai_n102_), .Y(mai_mai_n855_));
  OAI220     m0827(.A0(mai_mai_n845_), .A1(mai_mai_n414_), .B0(mai_mai_n328_), .B1(mai_mai_n855_), .Y(mai_mai_n856_));
  NOi31      m0828(.An(mai_mai_n217_), .B(mai_mai_n856_), .C(mai_mai_n295_), .Y(mai_mai_n857_));
  NA2        m0829(.A(c), .B(mai_mai_n111_), .Y(mai_mai_n858_));
  NO2        m0830(.A(mai_mai_n858_), .B(mai_mai_n398_), .Y(mai_mai_n859_));
  NA3        m0831(.A(mai_mai_n859_), .B(mai_mai_n501_), .C(f), .Y(mai_mai_n860_));
  OR2        m0832(.A(mai_mai_n640_), .B(mai_mai_n531_), .Y(mai_mai_n861_));
  INV        m0833(.A(mai_mai_n861_), .Y(mai_mai_n862_));
  NA2        m0834(.A(mai_mai_n784_), .B(mai_mai_n106_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n863_), .B(mai_mai_n862_), .Y(mai_mai_n864_));
  NA4        m0836(.A(mai_mai_n864_), .B(mai_mai_n860_), .C(mai_mai_n857_), .D(mai_mai_n853_), .Y(mai_mai_n865_));
  NO4        m0837(.A(mai_mai_n865_), .B(mai_mai_n849_), .C(mai_mai_n833_), .D(mai_mai_n820_), .Y(mai_mai_n866_));
  OR2        m0838(.A(mai_mai_n845_), .B(mai_mai_n69_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n107_), .B(j), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n806_), .B(g), .Y(mai_mai_n869_));
  AOI210     m0841(.A0(mai_mai_n869_), .A1(mai_mai_n282_), .B0(mai_mai_n867_), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n224_), .B(mai_mai_n218_), .Y(mai_mai_n871_));
  NA2        m0843(.A(mai_mai_n871_), .B(mai_mai_n221_), .Y(mai_mai_n872_));
  INV        m0844(.A(mai_mai_n872_), .Y(mai_mai_n873_));
  NA2        m0845(.A(e), .B(d), .Y(mai_mai_n874_));
  OAI220     m0846(.A0(mai_mai_n874_), .A1(c), .B0(mai_mai_n312_), .B1(d), .Y(mai_mai_n875_));
  NA3        m0847(.A(mai_mai_n875_), .B(mai_mai_n442_), .C(mai_mai_n499_), .Y(mai_mai_n876_));
  AOI210     m0848(.A0(mai_mai_n507_), .A1(mai_mai_n174_), .B0(mai_mai_n224_), .Y(mai_mai_n877_));
  AOI210     m0849(.A0(mai_mai_n607_), .A1(mai_mai_n337_), .B0(mai_mai_n877_), .Y(mai_mai_n878_));
  NA3        m0850(.A(mai_mai_n160_), .B(mai_mai_n81_), .C(mai_mai_n34_), .Y(mai_mai_n879_));
  NA3        m0851(.A(mai_mai_n879_), .B(mai_mai_n878_), .C(mai_mai_n876_), .Y(mai_mai_n880_));
  NO3        m0852(.A(mai_mai_n880_), .B(mai_mai_n873_), .C(mai_mai_n870_), .Y(mai_mai_n881_));
  NA2        m0853(.A(mai_mai_n821_), .B(mai_mai_n31_), .Y(mai_mai_n882_));
  AO210      m0854(.A0(mai_mai_n882_), .A1(mai_mai_n679_), .B0(mai_mai_n210_), .Y(mai_mai_n883_));
  OAI220     m0855(.A0(mai_mai_n606_), .A1(mai_mai_n58_), .B0(mai_mai_n290_), .B1(j), .Y(mai_mai_n884_));
  AOI220     m0856(.A0(mai_mai_n884_), .A1(mai_mai_n851_), .B0(mai_mai_n596_), .B1(mai_mai_n605_), .Y(mai_mai_n885_));
  OAI210     m0857(.A0(mai_mai_n811_), .A1(mai_mai_n164_), .B0(mai_mai_n885_), .Y(mai_mai_n886_));
  AOI210     m0858(.A0(mai_mai_n113_), .A1(mai_mai_n112_), .B0(mai_mai_n254_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n887_), .B(mai_mai_n840_), .Y(mai_mai_n888_));
  BUFFER     m0860(.A(mai_mai_n888_), .Y(mai_mai_n889_));
  NOi31      m0861(.An(mai_mai_n535_), .B(mai_mai_n837_), .C(mai_mai_n282_), .Y(mai_mai_n890_));
  NO3        m0862(.A(mai_mai_n890_), .B(mai_mai_n889_), .C(mai_mai_n886_), .Y(mai_mai_n891_));
  AO220      m0863(.A0(mai_mai_n442_), .A1(mai_mai_n723_), .B0(mai_mai_n169_), .B1(f), .Y(mai_mai_n892_));
  OAI210     m0864(.A0(mai_mai_n892_), .A1(mai_mai_n445_), .B0(mai_mai_n875_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n819_), .B(mai_mai_n683_), .Y(mai_mai_n894_));
  AN4        m0866(.A(mai_mai_n894_), .B(mai_mai_n893_), .C(mai_mai_n891_), .D(mai_mai_n883_), .Y(mai_mai_n895_));
  NA4        m0867(.A(mai_mai_n895_), .B(mai_mai_n881_), .C(mai_mai_n866_), .D(mai_mai_n813_), .Y(mai12));
  NO2        m0868(.A(mai_mai_n440_), .B(c), .Y(mai_mai_n897_));
  NO4        m0869(.A(mai_mai_n429_), .B(mai_mai_n247_), .C(mai_mai_n571_), .D(mai_mai_n207_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n898_), .B(mai_mai_n897_), .Y(mai_mai_n899_));
  NO2        m0871(.A(mai_mai_n440_), .B(mai_mai_n111_), .Y(mai_mai_n900_));
  NO2        m0872(.A(mai_mai_n822_), .B(mai_mai_n344_), .Y(mai_mai_n901_));
  NO2        m0873(.A(mai_mai_n640_), .B(mai_mai_n368_), .Y(mai_mai_n902_));
  AOI220     m0874(.A0(mai_mai_n902_), .A1(mai_mai_n533_), .B0(mai_mai_n901_), .B1(mai_mai_n900_), .Y(mai_mai_n903_));
  NA3        m0875(.A(mai_mai_n903_), .B(mai_mai_n899_), .C(mai_mai_n428_), .Y(mai_mai_n904_));
  AOI210     m0876(.A0(mai_mai_n227_), .A1(mai_mai_n327_), .B0(mai_mai_n196_), .Y(mai_mai_n905_));
  OR2        m0877(.A(mai_mai_n905_), .B(mai_mai_n898_), .Y(mai_mai_n906_));
  AOI210     m0878(.A0(mai_mai_n324_), .A1(mai_mai_n380_), .B0(mai_mai_n207_), .Y(mai_mai_n907_));
  OAI210     m0879(.A0(mai_mai_n907_), .A1(mai_mai_n906_), .B0(mai_mai_n393_), .Y(mai_mai_n908_));
  NO2        m0880(.A(mai_mai_n619_), .B(mai_mai_n256_), .Y(mai_mai_n909_));
  NO2        m0881(.A(mai_mai_n579_), .B(mai_mai_n815_), .Y(mai_mai_n910_));
  NA2        m0882(.A(mai_mai_n791_), .B(mai_mai_n909_), .Y(mai_mai_n911_));
  NO2        m0883(.A(mai_mai_n145_), .B(mai_mai_n230_), .Y(mai_mai_n912_));
  NA3        m0884(.A(mai_mai_n912_), .B(mai_mai_n233_), .C(i), .Y(mai_mai_n913_));
  NA3        m0885(.A(mai_mai_n913_), .B(mai_mai_n911_), .C(mai_mai_n908_), .Y(mai_mai_n914_));
  OR2        m0886(.A(mai_mai_n313_), .B(mai_mai_n900_), .Y(mai_mai_n915_));
  NA2        m0887(.A(mai_mai_n915_), .B(mai_mai_n345_), .Y(mai_mai_n916_));
  NO3        m0888(.A(mai_mai_n127_), .B(mai_mai_n146_), .C(mai_mai_n207_), .Y(mai_mai_n917_));
  NA2        m0889(.A(mai_mai_n917_), .B(mai_mai_n522_), .Y(mai_mai_n918_));
  NA4        m0890(.A(mai_mai_n430_), .B(mai_mai_n422_), .C(mai_mai_n175_), .D(g), .Y(mai_mai_n919_));
  NA3        m0891(.A(mai_mai_n919_), .B(mai_mai_n918_), .C(mai_mai_n916_), .Y(mai_mai_n920_));
  NO3        m0892(.A(mai_mai_n920_), .B(mai_mai_n914_), .C(mai_mai_n904_), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n576_), .B(mai_mai_n67_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n545_), .B(mai_mai_n139_), .Y(mai_mai_n924_));
  NOi21      m0896(.An(mai_mai_n34_), .B(mai_mai_n633_), .Y(mai_mai_n925_));
  AOI220     m0897(.A0(mai_mai_n925_), .A1(mai_mai_n924_), .B0(mai_mai_n923_), .B1(mai_mai_n922_), .Y(mai_mai_n926_));
  OAI210     m0898(.A0(mai_mai_n245_), .A1(mai_mai_n44_), .B0(mai_mai_n926_), .Y(mai_mai_n927_));
  NA2        m0899(.A(mai_mai_n420_), .B(mai_mai_n258_), .Y(mai_mai_n928_));
  NO3        m0900(.A(mai_mai_n793_), .B(mai_mai_n85_), .C(mai_mai_n398_), .Y(mai_mai_n929_));
  NAi31      m0901(.An(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n309_), .Y(mai_mai_n930_));
  NO2        m0902(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n931_));
  NO2        m0903(.A(mai_mai_n495_), .B(mai_mai_n290_), .Y(mai_mai_n932_));
  INV        m0904(.A(mai_mai_n932_), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n933_), .B(mai_mai_n139_), .Y(mai_mai_n934_));
  NA2        m0906(.A(mai_mai_n614_), .B(mai_mai_n354_), .Y(mai_mai_n935_));
  OAI210     m0907(.A0(mai_mai_n712_), .A1(mai_mai_n935_), .B0(mai_mai_n356_), .Y(mai_mai_n936_));
  NO4        m0908(.A(mai_mai_n936_), .B(mai_mai_n934_), .C(mai_mai_n930_), .D(mai_mai_n927_), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n337_), .B(g), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n157_), .B(i), .Y(mai_mai_n939_));
  NA2        m0911(.A(mai_mai_n45_), .B(i), .Y(mai_mai_n940_));
  OAI220     m0912(.A0(mai_mai_n940_), .A1(mai_mai_n195_), .B0(mai_mai_n939_), .B1(mai_mai_n87_), .Y(mai_mai_n941_));
  AOI210     m0913(.A0(mai_mai_n406_), .A1(mai_mai_n37_), .B0(mai_mai_n941_), .Y(mai_mai_n942_));
  NO2        m0914(.A(mai_mai_n139_), .B(mai_mai_n80_), .Y(mai_mai_n943_));
  OR2        m0915(.A(mai_mai_n943_), .B(mai_mai_n544_), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n545_), .B(mai_mai_n372_), .Y(mai_mai_n945_));
  AOI210     m0917(.A0(mai_mai_n945_), .A1(n), .B0(mai_mai_n944_), .Y(mai_mai_n946_));
  OAI220     m0918(.A0(mai_mai_n946_), .A1(mai_mai_n938_), .B0(mai_mai_n942_), .B1(mai_mai_n321_), .Y(mai_mai_n947_));
  OR3        m0919(.A(mai_mai_n300_), .B(mai_mai_n419_), .C(f), .Y(mai_mai_n948_));
  NA3        m0920(.A(mai_mai_n314_), .B(mai_mai_n113_), .C(g), .Y(mai_mai_n949_));
  AOI210     m0921(.A0(mai_mai_n651_), .A1(mai_mai_n949_), .B0(m), .Y(mai_mai_n950_));
  OAI210     m0922(.A0(mai_mai_n950_), .A1(mai_mai_n901_), .B0(mai_mai_n313_), .Y(mai_mai_n951_));
  NA2        m0923(.A(mai_mai_n670_), .B(mai_mai_n854_), .Y(mai_mai_n952_));
  INV        m0924(.A(mai_mai_n425_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n215_), .B(mai_mai_n73_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n954_), .B(mai_mai_n948_), .Y(mai_mai_n955_));
  AOI220     m0927(.A0(mai_mai_n955_), .A1(mai_mai_n253_), .B0(mai_mai_n953_), .B1(mai_mai_n952_), .Y(mai_mai_n956_));
  NA2        m0928(.A(mai_mai_n956_), .B(mai_mai_n951_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n642_), .B(mai_mai_n84_), .Y(mai_mai_n958_));
  NO2        m0930(.A(mai_mai_n448_), .B(mai_mai_n207_), .Y(mai_mai_n959_));
  AOI220     m0931(.A0(mai_mai_n959_), .A1(mai_mai_n373_), .B0(mai_mai_n915_), .B1(mai_mai_n211_), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n960_), .B(mai_mai_n958_), .Y(mai_mai_n961_));
  OAI210     m0933(.A0(mai_mai_n953_), .A1(mai_mai_n910_), .B0(mai_mai_n533_), .Y(mai_mai_n962_));
  OAI210     m0934(.A0(mai_mai_n359_), .A1(mai_mai_n358_), .B0(mai_mai_n104_), .Y(mai_mai_n963_));
  NA2        m0935(.A(mai_mai_n963_), .B(mai_mai_n526_), .Y(mai_mai_n964_));
  NA2        m0936(.A(mai_mai_n950_), .B(mai_mai_n900_), .Y(mai_mai_n965_));
  NO3        m0937(.A(mai_mai_n868_), .B(mai_mai_n47_), .C(mai_mai_n44_), .Y(mai_mai_n966_));
  AOI220     m0938(.A0(mai_mai_n966_), .A1(mai_mai_n610_), .B0(mai_mai_n624_), .B1(mai_mai_n522_), .Y(mai_mai_n967_));
  NA4        m0939(.A(mai_mai_n967_), .B(mai_mai_n965_), .C(mai_mai_n964_), .D(mai_mai_n962_), .Y(mai_mai_n968_));
  NO4        m0940(.A(mai_mai_n968_), .B(mai_mai_n961_), .C(mai_mai_n957_), .D(mai_mai_n947_), .Y(mai_mai_n969_));
  NAi31      m0941(.An(mai_mai_n136_), .B(mai_mai_n407_), .C(n), .Y(mai_mai_n970_));
  NO3        m0942(.A(mai_mai_n121_), .B(mai_mai_n330_), .C(mai_mai_n823_), .Y(mai_mai_n971_));
  NO2        m0943(.A(mai_mai_n971_), .B(mai_mai_n970_), .Y(mai_mai_n972_));
  NO3        m0944(.A(mai_mai_n266_), .B(mai_mai_n136_), .C(mai_mai_n398_), .Y(mai_mai_n973_));
  AOI210     m0945(.A0(mai_mai_n973_), .A1(mai_mai_n489_), .B0(mai_mai_n972_), .Y(mai_mai_n974_));
  NA2        m0946(.A(mai_mai_n481_), .B(i), .Y(mai_mai_n975_));
  NA2        m0947(.A(mai_mai_n975_), .B(mai_mai_n974_), .Y(mai_mai_n976_));
  NA2        m0948(.A(mai_mai_n224_), .B(mai_mai_n165_), .Y(mai_mai_n977_));
  NO3        m0949(.A(mai_mai_n297_), .B(mai_mai_n430_), .C(mai_mai_n169_), .Y(mai_mai_n978_));
  NOi31      m0950(.An(mai_mai_n977_), .B(mai_mai_n978_), .C(mai_mai_n207_), .Y(mai_mai_n979_));
  NAi21      m0951(.An(mai_mai_n545_), .B(mai_mai_n959_), .Y(mai_mai_n980_));
  NA2        m0952(.A(mai_mai_n423_), .B(mai_mai_n854_), .Y(mai_mai_n981_));
  NO3        m0953(.A(mai_mai_n424_), .B(mai_mai_n300_), .C(mai_mai_n69_), .Y(mai_mai_n982_));
  AOI220     m0954(.A0(mai_mai_n982_), .A1(mai_mai_n981_), .B0(mai_mai_n470_), .B1(g), .Y(mai_mai_n983_));
  NA2        m0955(.A(mai_mai_n983_), .B(mai_mai_n980_), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n905_), .B(mai_mai_n897_), .Y(mai_mai_n985_));
  NO3        m0957(.A(mai_mai_n534_), .B(mai_mai_n143_), .C(mai_mai_n206_), .Y(mai_mai_n986_));
  OAI210     m0958(.A0(mai_mai_n986_), .A1(mai_mai_n517_), .B0(mai_mai_n369_), .Y(mai_mai_n987_));
  OAI220     m0959(.A0(mai_mai_n902_), .A1(mai_mai_n910_), .B0(mai_mai_n535_), .B1(mai_mai_n413_), .Y(mai_mai_n988_));
  NA4        m0960(.A(mai_mai_n988_), .B(mai_mai_n987_), .C(mai_mai_n985_), .D(mai_mai_n604_), .Y(mai_mai_n989_));
  OAI210     m0961(.A0(mai_mai_n905_), .A1(mai_mai_n898_), .B0(mai_mai_n977_), .Y(mai_mai_n990_));
  NA3        m0962(.A(mai_mai_n945_), .B(mai_mai_n475_), .C(mai_mai_n45_), .Y(mai_mai_n991_));
  NA2        m0963(.A(mai_mai_n371_), .B(mai_mai_n369_), .Y(mai_mai_n992_));
  NA3        m0964(.A(mai_mai_n992_), .B(mai_mai_n991_), .C(mai_mai_n990_), .Y(mai_mai_n993_));
  OR2        m0965(.A(mai_mai_n993_), .B(mai_mai_n989_), .Y(mai_mai_n994_));
  NO4        m0966(.A(mai_mai_n994_), .B(mai_mai_n984_), .C(mai_mai_n979_), .D(mai_mai_n976_), .Y(mai_mai_n995_));
  NA4        m0967(.A(mai_mai_n995_), .B(mai_mai_n969_), .C(mai_mai_n937_), .D(mai_mai_n921_), .Y(mai13));
  INV        m0968(.A(mai_mai_n45_), .Y(mai_mai_n997_));
  AN2        m0969(.A(c), .B(b), .Y(mai_mai_n998_));
  NA3        m0970(.A(mai_mai_n244_), .B(mai_mai_n998_), .C(m), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n486_), .B(f), .Y(mai_mai_n1000_));
  NO4        m0972(.A(mai_mai_n1000_), .B(mai_mai_n999_), .C(mai_mai_n997_), .D(mai_mai_n572_), .Y(mai_mai_n1001_));
  NA2        m0973(.A(mai_mai_n258_), .B(mai_mai_n998_), .Y(mai_mai_n1002_));
  NO4        m0974(.A(mai_mai_n1002_), .B(mai_mai_n1000_), .C(mai_mai_n939_), .D(a), .Y(mai_mai_n1003_));
  NAi32      m0975(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1004_));
  NA2        m0976(.A(mai_mai_n135_), .B(mai_mai_n44_), .Y(mai_mai_n1005_));
  NO4        m0977(.A(mai_mai_n1005_), .B(mai_mai_n1004_), .C(mai_mai_n579_), .D(mai_mai_n296_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n646_), .B(mai_mai_n218_), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n401_), .B(mai_mai_n206_), .Y(mai_mai_n1008_));
  AN2        m0980(.A(d), .B(c), .Y(mai_mai_n1009_));
  NA2        m0981(.A(mai_mai_n1009_), .B(mai_mai_n111_), .Y(mai_mai_n1010_));
  NO4        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1008_), .C(mai_mai_n170_), .D(mai_mai_n161_), .Y(mai_mai_n1011_));
  NA2        m0983(.A(mai_mai_n486_), .B(c), .Y(mai_mai_n1012_));
  NO4        m0984(.A(mai_mai_n1005_), .B(mai_mai_n575_), .C(mai_mai_n1012_), .D(mai_mai_n296_), .Y(mai_mai_n1013_));
  AO210      m0985(.A0(mai_mai_n1011_), .A1(mai_mai_n1007_), .B0(mai_mai_n1013_), .Y(mai_mai_n1014_));
  OR4        m0986(.A(mai_mai_n1014_), .B(mai_mai_n1006_), .C(mai_mai_n1003_), .D(mai_mai_n1001_), .Y(mai_mai_n1015_));
  NAi32      m0987(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1016_));
  NO2        m0988(.A(mai_mai_n1016_), .B(mai_mai_n140_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n1017_), .B(g), .Y(mai_mai_n1018_));
  OR3        m0990(.A(mai_mai_n218_), .B(mai_mai_n170_), .C(mai_mai_n161_), .Y(mai_mai_n1019_));
  NO2        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1018_), .Y(mai_mai_n1020_));
  NO2        m0992(.A(mai_mai_n1012_), .B(mai_mai_n296_), .Y(mai_mai_n1021_));
  NO2        m0993(.A(j), .B(mai_mai_n44_), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n613_), .B(mai_mai_n1022_), .Y(mai_mai_n1023_));
  NOi21      m0995(.An(mai_mai_n1021_), .B(mai_mai_n1023_), .Y(mai_mai_n1024_));
  NO2        m0996(.A(mai_mai_n737_), .B(mai_mai_n107_), .Y(mai_mai_n1025_));
  NOi41      m0997(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n1026_), .B(mai_mai_n1025_), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n1027_), .B(mai_mai_n1018_), .Y(mai_mai_n1028_));
  OR3        m1000(.A(e), .B(d), .C(c), .Y(mai_mai_n1029_));
  NA3        m1001(.A(k), .B(j), .C(i), .Y(mai_mai_n1030_));
  NO3        m1002(.A(mai_mai_n1030_), .B(mai_mai_n296_), .C(mai_mai_n86_), .Y(mai_mai_n1031_));
  NOi21      m1003(.An(mai_mai_n1031_), .B(mai_mai_n1029_), .Y(mai_mai_n1032_));
  OR4        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1028_), .C(mai_mai_n1024_), .D(mai_mai_n1020_), .Y(mai_mai_n1033_));
  NA3        m1005(.A(mai_mai_n456_), .B(mai_mai_n323_), .C(mai_mai_n54_), .Y(mai_mai_n1034_));
  NO2        m1006(.A(mai_mai_n1034_), .B(mai_mai_n1023_), .Y(mai_mai_n1035_));
  NO4        m1007(.A(mai_mai_n1034_), .B(mai_mai_n575_), .C(mai_mai_n437_), .D(mai_mai_n44_), .Y(mai_mai_n1036_));
  NO2        m1008(.A(f), .B(c), .Y(mai_mai_n1037_));
  NOi21      m1009(.An(mai_mai_n1037_), .B(mai_mai_n429_), .Y(mai_mai_n1038_));
  NA2        m1010(.A(mai_mai_n1038_), .B(mai_mai_n57_), .Y(mai_mai_n1039_));
  OR2        m1011(.A(k), .B(i), .Y(mai_mai_n1040_));
  NO3        m1012(.A(mai_mai_n1040_), .B(mai_mai_n237_), .C(l), .Y(mai_mai_n1041_));
  NOi31      m1013(.An(mai_mai_n1041_), .B(mai_mai_n1039_), .C(j), .Y(mai_mai_n1042_));
  OR3        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1036_), .C(mai_mai_n1035_), .Y(mai_mai_n1043_));
  OR3        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1033_), .C(mai_mai_n1015_), .Y(mai02));
  OR2        m1016(.A(l), .B(k), .Y(mai_mai_n1045_));
  OR3        m1017(.A(h), .B(g), .C(f), .Y(mai_mai_n1046_));
  OR3        m1018(.A(n), .B(m), .C(i), .Y(mai_mai_n1047_));
  NO4        m1019(.A(mai_mai_n1047_), .B(mai_mai_n1046_), .C(mai_mai_n1045_), .D(mai_mai_n1029_), .Y(mai_mai_n1048_));
  NO2        m1020(.A(d), .B(c), .Y(mai_mai_n1049_));
  AOI210     m1021(.A0(mai_mai_n1031_), .A1(mai_mai_n1049_), .B0(mai_mai_n1006_), .Y(mai_mai_n1050_));
  AN3        m1022(.A(g), .B(f), .C(c), .Y(mai_mai_n1051_));
  NA3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n456_), .C(h), .Y(mai_mai_n1052_));
  OR2        m1024(.A(mai_mai_n1030_), .B(mai_mai_n296_), .Y(mai_mai_n1053_));
  OR2        m1025(.A(mai_mai_n1053_), .B(mai_mai_n1052_), .Y(mai_mai_n1054_));
  NO3        m1026(.A(mai_mai_n1034_), .B(mai_mai_n1005_), .C(mai_mai_n575_), .Y(mai_mai_n1055_));
  NO2        m1027(.A(mai_mai_n1055_), .B(mai_mai_n1020_), .Y(mai_mai_n1056_));
  NA3        m1028(.A(l), .B(k), .C(j), .Y(mai_mai_n1057_));
  NA2        m1029(.A(i), .B(h), .Y(mai_mai_n1058_));
  NO3        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1057_), .C(mai_mai_n127_), .Y(mai_mai_n1059_));
  NO3        m1031(.A(mai_mai_n137_), .B(mai_mai_n277_), .C(mai_mai_n207_), .Y(mai_mai_n1060_));
  AOI210     m1032(.A0(mai_mai_n1060_), .A1(mai_mai_n1059_), .B0(mai_mai_n1024_), .Y(mai_mai_n1061_));
  NA3        m1033(.A(c), .B(b), .C(a), .Y(mai_mai_n1062_));
  NO3        m1034(.A(mai_mai_n1062_), .B(mai_mai_n874_), .C(mai_mai_n206_), .Y(mai_mai_n1063_));
  NO4        m1035(.A(mai_mai_n1030_), .B(mai_mai_n290_), .C(mai_mai_n47_), .D(mai_mai_n107_), .Y(mai_mai_n1064_));
  AOI210     m1036(.A0(mai_mai_n1064_), .A1(mai_mai_n1063_), .B0(mai_mai_n1035_), .Y(mai_mai_n1065_));
  AN4        m1037(.A(mai_mai_n1065_), .B(mai_mai_n1061_), .C(mai_mai_n1056_), .D(mai_mai_n1054_), .Y(mai_mai_n1066_));
  NO2        m1038(.A(mai_mai_n1010_), .B(mai_mai_n1008_), .Y(mai_mai_n1067_));
  NA2        m1039(.A(mai_mai_n1027_), .B(mai_mai_n1019_), .Y(mai_mai_n1068_));
  AOI210     m1040(.A0(mai_mai_n1068_), .A1(mai_mai_n1067_), .B0(mai_mai_n1001_), .Y(mai_mai_n1069_));
  NAi41      m1041(.An(mai_mai_n1048_), .B(mai_mai_n1069_), .C(mai_mai_n1066_), .D(mai_mai_n1050_), .Y(mai03));
  NO2        m1042(.A(mai_mai_n519_), .B(mai_mai_n583_), .Y(mai_mai_n1071_));
  NA4        m1043(.A(mai_mai_n564_), .B(m), .C(mai_mai_n107_), .D(mai_mai_n206_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n1072_), .B(mai_mai_n360_), .Y(mai_mai_n1073_));
  NO3        m1045(.A(mai_mai_n1073_), .B(mai_mai_n1071_), .C(mai_mai_n963_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n828_), .B(mai_mai_n817_), .Y(mai_mai_n1075_));
  OAI220     m1047(.A0(mai_mai_n1075_), .A1(mai_mai_n670_), .B0(mai_mai_n1074_), .B1(mai_mai_n576_), .Y(mai_mai_n1076_));
  NOi31      m1048(.An(m), .B(n), .C(f), .Y(mai_mai_n1077_));
  NA2        m1049(.A(mai_mai_n1077_), .B(mai_mai_n49_), .Y(mai_mai_n1078_));
  AN2        m1050(.A(e), .B(c), .Y(mai_mai_n1079_));
  NA2        m1051(.A(mai_mai_n1079_), .B(a), .Y(mai_mai_n1080_));
  OAI220     m1052(.A0(mai_mai_n1080_), .A1(mai_mai_n1078_), .B0(mai_mai_n861_), .B1(mai_mai_n412_), .Y(mai_mai_n1081_));
  NA2        m1053(.A(mai_mai_n499_), .B(l), .Y(mai_mai_n1082_));
  NOi31      m1054(.An(mai_mai_n839_), .B(mai_mai_n999_), .C(mai_mai_n1082_), .Y(mai_mai_n1083_));
  NO2        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1081_), .Y(mai_mai_n1084_));
  NO2        m1056(.A(mai_mai_n277_), .B(a), .Y(mai_mai_n1085_));
  INV        m1057(.A(mai_mai_n1006_), .Y(mai_mai_n1086_));
  NO2        m1058(.A(mai_mai_n1058_), .B(mai_mai_n473_), .Y(mai_mai_n1087_));
  NO2        m1059(.A(mai_mai_n83_), .B(g), .Y(mai_mai_n1088_));
  AOI210     m1060(.A0(mai_mai_n1088_), .A1(mai_mai_n1087_), .B0(mai_mai_n1041_), .Y(mai_mai_n1089_));
  OR2        m1061(.A(mai_mai_n1089_), .B(mai_mai_n1039_), .Y(mai_mai_n1090_));
  NA3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1086_), .C(mai_mai_n1084_), .Y(mai_mai_n1091_));
  NO4        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1076_), .C(mai_mai_n795_), .D(mai_mai_n554_), .Y(mai_mai_n1092_));
  NA2        m1064(.A(c), .B(b), .Y(mai_mai_n1093_));
  NO2        m1065(.A(mai_mai_n682_), .B(mai_mai_n1093_), .Y(mai_mai_n1094_));
  OAI210     m1066(.A0(mai_mai_n837_), .A1(mai_mai_n809_), .B0(mai_mai_n402_), .Y(mai_mai_n1095_));
  OAI210     m1067(.A0(mai_mai_n1095_), .A1(mai_mai_n838_), .B0(mai_mai_n1094_), .Y(mai_mai_n1096_));
  NAi21      m1068(.An(mai_mai_n404_), .B(mai_mai_n1094_), .Y(mai_mai_n1097_));
  NA3        m1069(.A(mai_mai_n413_), .B(mai_mai_n550_), .C(f), .Y(mai_mai_n1098_));
  OAI210     m1070(.A0(mai_mai_n539_), .A1(mai_mai_n39_), .B0(mai_mai_n1085_), .Y(mai_mai_n1099_));
  NA3        m1071(.A(mai_mai_n1099_), .B(mai_mai_n1098_), .C(mai_mai_n1097_), .Y(mai_mai_n1100_));
  INV        m1072(.A(mai_mai_n114_), .Y(mai_mai_n1101_));
  NA2        m1073(.A(mai_mai_n1101_), .B(g), .Y(mai_mai_n1102_));
  NAi21      m1074(.An(f), .B(d), .Y(mai_mai_n1103_));
  NO2        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1062_), .Y(mai_mai_n1104_));
  INV        m1076(.A(mai_mai_n1104_), .Y(mai_mai_n1105_));
  AOI210     m1077(.A0(mai_mai_n1102_), .A1(mai_mai_n282_), .B0(mai_mai_n1105_), .Y(mai_mai_n1106_));
  AOI210     m1078(.A0(mai_mai_n1106_), .A1(mai_mai_n108_), .B0(mai_mai_n1100_), .Y(mai_mai_n1107_));
  NA2        m1079(.A(mai_mai_n887_), .B(mai_mai_n1082_), .Y(mai_mai_n1108_));
  NA2        m1080(.A(mai_mai_n153_), .B(mai_mai_n33_), .Y(mai_mai_n1109_));
  AOI210     m1081(.A0(mai_mai_n935_), .A1(mai_mai_n1109_), .B0(mai_mai_n207_), .Y(mai_mai_n1110_));
  NA2        m1082(.A(mai_mai_n1110_), .B(mai_mai_n1104_), .Y(mai_mai_n1111_));
  INV        m1083(.A(mai_mai_n929_), .Y(mai_mai_n1112_));
  NA2        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1111_), .Y(mai_mai_n1113_));
  INV        m1085(.A(mai_mai_n1113_), .Y(mai_mai_n1114_));
  NA4        m1086(.A(mai_mai_n1114_), .B(mai_mai_n1107_), .C(mai_mai_n1096_), .D(mai_mai_n1092_), .Y(mai00));
  AOI210     m1087(.A0(mai_mai_n289_), .A1(mai_mai_n207_), .B0(mai_mai_n269_), .Y(mai_mai_n1116_));
  NO2        m1088(.A(mai_mai_n1116_), .B(mai_mai_n567_), .Y(mai_mai_n1117_));
  NO2        m1089(.A(mai_mai_n1055_), .B(mai_mai_n929_), .Y(mai_mai_n1118_));
  NA2        m1090(.A(mai_mai_n1118_), .B(mai_mai_n964_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n501_), .B(f), .Y(mai_mai_n1120_));
  OAI210     m1092(.A0(mai_mai_n971_), .A1(mai_mai_n40_), .B0(mai_mai_n626_), .Y(mai_mai_n1121_));
  NA3        m1093(.A(mai_mai_n1121_), .B(mai_mai_n252_), .C(n), .Y(mai_mai_n1122_));
  AOI210     m1094(.A0(mai_mai_n1122_), .A1(mai_mai_n1120_), .B0(mai_mai_n1010_), .Y(mai_mai_n1123_));
  NO4        m1095(.A(mai_mai_n1123_), .B(mai_mai_n1119_), .C(mai_mai_n1117_), .D(mai_mai_n1033_), .Y(mai_mai_n1124_));
  NA3        m1096(.A(mai_mai_n160_), .B(mai_mai_n45_), .C(mai_mai_n44_), .Y(mai_mai_n1125_));
  NA3        m1097(.A(d), .B(mai_mai_n54_), .C(b), .Y(mai_mai_n1126_));
  NOi31      m1098(.An(n), .B(m), .C(i), .Y(mai_mai_n1127_));
  NA3        m1099(.A(mai_mai_n1127_), .B(mai_mai_n629_), .C(mai_mai_n49_), .Y(mai_mai_n1128_));
  OAI210     m1100(.A0(mai_mai_n1126_), .A1(mai_mai_n1125_), .B0(mai_mai_n1128_), .Y(mai_mai_n1129_));
  INV        m1101(.A(mai_mai_n566_), .Y(mai_mai_n1130_));
  NO3        m1102(.A(mai_mai_n1130_), .B(mai_mai_n1129_), .C(mai_mai_n890_), .Y(mai_mai_n1131_));
  NO4        m1103(.A(mai_mai_n476_), .B(mai_mai_n347_), .C(mai_mai_n1093_), .D(mai_mai_n57_), .Y(mai_mai_n1132_));
  NA3        m1104(.A(mai_mai_n374_), .B(mai_mai_n214_), .C(g), .Y(mai_mai_n1133_));
  OA220      m1105(.A0(mai_mai_n1133_), .A1(mai_mai_n1126_), .B0(mai_mai_n375_), .B1(mai_mai_n130_), .Y(mai_mai_n1134_));
  NO2        m1106(.A(h), .B(g), .Y(mai_mai_n1135_));
  NA4        m1107(.A(mai_mai_n489_), .B(mai_mai_n456_), .C(mai_mai_n1135_), .D(mai_mai_n998_), .Y(mai_mai_n1136_));
  OAI220     m1108(.A0(mai_mai_n519_), .A1(mai_mai_n583_), .B0(mai_mai_n87_), .B1(mai_mai_n86_), .Y(mai_mai_n1137_));
  AOI220     m1109(.A0(mai_mai_n1137_), .A1(mai_mai_n526_), .B0(mai_mai_n917_), .B1(mai_mai_n565_), .Y(mai_mai_n1138_));
  AOI220     m1110(.A0(mai_mai_n306_), .A1(mai_mai_n241_), .B0(mai_mai_n171_), .B1(mai_mai_n142_), .Y(mai_mai_n1139_));
  NA4        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1138_), .C(mai_mai_n1136_), .D(mai_mai_n1134_), .Y(mai_mai_n1140_));
  NO3        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1132_), .C(mai_mai_n260_), .Y(mai_mai_n1141_));
  INV        m1113(.A(mai_mai_n311_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n241_), .B(mai_mai_n337_), .Y(mai_mai_n1143_));
  NA3        m1115(.A(mai_mai_n1143_), .B(mai_mai_n1142_), .C(mai_mai_n148_), .Y(mai_mai_n1144_));
  NA3        m1116(.A(mai_mai_n173_), .B(mai_mai_n107_), .C(g), .Y(mai_mai_n1145_));
  NA3        m1117(.A(mai_mai_n456_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1146_));
  NOi31      m1118(.An(mai_mai_n847_), .B(mai_mai_n1146_), .C(mai_mai_n1145_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n268_), .B(mai_mai_n69_), .Y(mai_mai_n1148_));
  NO3        m1120(.A(mai_mai_n412_), .B(mai_mai_n805_), .C(n), .Y(mai_mai_n1149_));
  AOI210     m1121(.A0(mai_mai_n1149_), .A1(mai_mai_n1148_), .B0(mai_mai_n1048_), .Y(mai_mai_n1150_));
  NAi31      m1122(.An(mai_mai_n1013_), .B(mai_mai_n1150_), .C(mai_mai_n68_), .Y(mai_mai_n1151_));
  NO3        m1123(.A(mai_mai_n1151_), .B(mai_mai_n1147_), .C(mai_mai_n1144_), .Y(mai_mai_n1152_));
  AN3        m1124(.A(mai_mai_n1152_), .B(mai_mai_n1141_), .C(mai_mai_n1131_), .Y(mai_mai_n1153_));
  NA3        m1125(.A(mai_mai_n1077_), .B(mai_mai_n590_), .C(mai_mai_n455_), .Y(mai_mai_n1154_));
  NA2        m1126(.A(mai_mai_n1154_), .B(mai_mai_n235_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n1073_), .B(mai_mai_n526_), .Y(mai_mai_n1156_));
  NA2        m1128(.A(mai_mai_n1156_), .B(mai_mai_n286_), .Y(mai_mai_n1157_));
  OAI210     m1129(.A0(mai_mai_n454_), .A1(mai_mai_n115_), .B0(mai_mai_n840_), .Y(mai_mai_n1158_));
  NA2        m1130(.A(mai_mai_n1158_), .B(mai_mai_n1108_), .Y(mai_mai_n1159_));
  OR4        m1131(.A(mai_mai_n1010_), .B(mai_mai_n266_), .C(mai_mai_n216_), .D(e), .Y(mai_mai_n1160_));
  NO2        m1132(.A(mai_mai_n210_), .B(mai_mai_n207_), .Y(mai_mai_n1161_));
  NA2        m1133(.A(n), .B(e), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n1162_), .B(mai_mai_n140_), .Y(mai_mai_n1163_));
  AOI220     m1135(.A0(mai_mai_n1163_), .A1(mai_mai_n267_), .B0(mai_mai_n821_), .B1(mai_mai_n1161_), .Y(mai_mai_n1164_));
  NA3        m1136(.A(mai_mai_n1164_), .B(mai_mai_n1160_), .C(mai_mai_n1159_), .Y(mai_mai_n1165_));
  AOI210     m1137(.A0(mai_mai_n1163_), .A1(mai_mai_n825_), .B0(mai_mai_n794_), .Y(mai_mai_n1166_));
  AOI220     m1138(.A0(mai_mai_n925_), .A1(mai_mai_n565_), .B0(mai_mai_n629_), .B1(mai_mai_n238_), .Y(mai_mai_n1167_));
  NO2        m1139(.A(mai_mai_n63_), .B(h), .Y(mai_mai_n1168_));
  NO3        m1140(.A(mai_mai_n1010_), .B(mai_mai_n1008_), .C(mai_mai_n705_), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n1045_), .B(mai_mai_n127_), .Y(mai_mai_n1170_));
  AN2        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1060_), .Y(mai_mai_n1171_));
  OAI210     m1143(.A0(mai_mai_n1171_), .A1(mai_mai_n1169_), .B0(mai_mai_n1168_), .Y(mai_mai_n1172_));
  NA4        m1144(.A(mai_mai_n1172_), .B(mai_mai_n1167_), .C(mai_mai_n1166_), .D(mai_mai_n842_), .Y(mai_mai_n1173_));
  NO4        m1145(.A(mai_mai_n1173_), .B(mai_mai_n1165_), .C(mai_mai_n1157_), .D(mai_mai_n1155_), .Y(mai_mai_n1174_));
  NA2        m1146(.A(mai_mai_n810_), .B(mai_mai_n733_), .Y(mai_mai_n1175_));
  NA4        m1147(.A(mai_mai_n1175_), .B(mai_mai_n1174_), .C(mai_mai_n1153_), .D(mai_mai_n1124_), .Y(mai01));
  AN2        m1148(.A(mai_mai_n987_), .B(mai_mai_n985_), .Y(mai_mai_n1177_));
  NO4        m1149(.A(mai_mai_n779_), .B(mai_mai_n772_), .C(mai_mai_n467_), .D(mai_mai_n275_), .Y(mai_mai_n1178_));
  NA2        m1150(.A(mai_mai_n385_), .B(i), .Y(mai_mai_n1179_));
  NA3        m1151(.A(mai_mai_n1179_), .B(mai_mai_n1178_), .C(mai_mai_n1177_), .Y(mai_mai_n1180_));
  NA2        m1152(.A(mai_mai_n545_), .B(mai_mai_n265_), .Y(mai_mai_n1181_));
  NA2        m1153(.A(mai_mai_n932_), .B(mai_mai_n1181_), .Y(mai_mai_n1182_));
  NA3        m1154(.A(mai_mai_n1182_), .B(mai_mai_n885_), .C(mai_mai_n322_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n44_), .B(f), .Y(mai_mai_n1184_));
  NA2        m1156(.A(mai_mai_n688_), .B(mai_mai_n92_), .Y(mai_mai_n1185_));
  NO2        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1184_), .Y(mai_mai_n1186_));
  INV        m1158(.A(mai_mai_n113_), .Y(mai_mai_n1187_));
  OA220      m1159(.A0(mai_mai_n1187_), .A1(mai_mai_n574_), .B0(mai_mai_n641_), .B1(mai_mai_n360_), .Y(mai_mai_n1188_));
  NAi31      m1160(.An(mai_mai_n156_), .B(mai_mai_n1188_), .C(mai_mai_n872_), .Y(mai_mai_n1189_));
  NO3        m1161(.A(mai_mai_n760_), .B(mai_mai_n653_), .C(mai_mai_n504_), .Y(mai_mai_n1190_));
  OR2        m1162(.A(mai_mai_n190_), .B(mai_mai_n188_), .Y(mai_mai_n1191_));
  NA3        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1190_), .C(mai_mai_n133_), .Y(mai_mai_n1192_));
  NO4        m1164(.A(mai_mai_n1192_), .B(mai_mai_n1189_), .C(mai_mai_n1183_), .D(mai_mai_n1180_), .Y(mai_mai_n1193_));
  INV        m1165(.A(mai_mai_n1133_), .Y(mai_mai_n1194_));
  NA2        m1166(.A(mai_mai_n1194_), .B(mai_mai_n522_), .Y(mai_mai_n1195_));
  NA2        m1167(.A(mai_mai_n528_), .B(mai_mai_n387_), .Y(mai_mai_n1196_));
  NOi21      m1168(.An(mai_mai_n551_), .B(mai_mai_n571_), .Y(mai_mai_n1197_));
  NA2        m1169(.A(mai_mai_n1197_), .B(mai_mai_n1196_), .Y(mai_mai_n1198_));
  NO2        m1170(.A(mai_mai_n199_), .B(mai_mai_n206_), .Y(mai_mai_n1199_));
  OAI210     m1171(.A0(mai_mai_n785_), .A1(mai_mai_n413_), .B0(mai_mai_n1199_), .Y(mai_mai_n1200_));
  NA3        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1198_), .C(mai_mai_n1195_), .Y(mai_mai_n1201_));
  INV        m1173(.A(mai_mai_n584_), .Y(mai_mai_n1202_));
  OAI210     m1174(.A0(mai_mai_n1187_), .A1(mai_mai_n581_), .B0(mai_mai_n1202_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n274_), .B(mai_mai_n190_), .Y(mai_mai_n1204_));
  NA2        m1176(.A(mai_mai_n1204_), .B(mai_mai_n645_), .Y(mai_mai_n1205_));
  INV        m1177(.A(mai_mai_n929_), .Y(mai_mai_n1206_));
  OAI210     m1178(.A0(mai_mai_n1186_), .A1(mai_mai_n316_), .B0(mai_mai_n654_), .Y(mai_mai_n1207_));
  NA4        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1206_), .C(mai_mai_n1205_), .D(mai_mai_n762_), .Y(mai_mai_n1208_));
  NO3        m1180(.A(mai_mai_n1208_), .B(mai_mai_n1203_), .C(mai_mai_n1201_), .Y(mai_mai_n1209_));
  NA3        m1181(.A(mai_mai_n587_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1210_));
  NO2        m1182(.A(mai_mai_n1210_), .B(mai_mai_n199_), .Y(mai_mai_n1211_));
  AOI210     m1183(.A0(mai_mai_n496_), .A1(mai_mai_n56_), .B0(mai_mai_n1211_), .Y(mai_mai_n1212_));
  OR3        m1184(.A(mai_mai_n1185_), .B(mai_mai_n588_), .C(mai_mai_n1184_), .Y(mai_mai_n1213_));
  INV        m1185(.A(mai_mai_n1129_), .Y(mai_mai_n1214_));
  NA4        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1213_), .C(mai_mai_n1212_), .D(mai_mai_n732_), .Y(mai_mai_n1215_));
  NO2        m1187(.A(mai_mai_n939_), .B(mai_mai_n226_), .Y(mai_mai_n1216_));
  NO2        m1188(.A(mai_mai_n940_), .B(mai_mai_n547_), .Y(mai_mai_n1217_));
  OAI210     m1189(.A0(mai_mai_n1217_), .A1(mai_mai_n1216_), .B0(mai_mai_n330_), .Y(mai_mai_n1218_));
  NA2        m1190(.A(mai_mai_n560_), .B(mai_mai_n558_), .Y(mai_mai_n1219_));
  NO3        m1191(.A(mai_mai_n75_), .B(mai_mai_n290_), .C(mai_mai_n44_), .Y(mai_mai_n1220_));
  NA2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n544_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n1221_), .B(mai_mai_n1219_), .Y(mai_mai_n1222_));
  OR2        m1194(.A(mai_mai_n1133_), .B(mai_mai_n1126_), .Y(mai_mai_n1223_));
  NA2        m1195(.A(mai_mai_n1220_), .B(mai_mai_n786_), .Y(mai_mai_n1224_));
  NA3        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1223_), .C(mai_mai_n377_), .Y(mai_mai_n1225_));
  NOi41      m1197(.An(mai_mai_n1218_), .B(mai_mai_n1225_), .C(mai_mai_n1222_), .D(mai_mai_n1215_), .Y(mai_mai_n1226_));
  NO2        m1198(.A(mai_mai_n126_), .B(mai_mai_n44_), .Y(mai_mai_n1227_));
  NO2        m1199(.A(mai_mai_n44_), .B(mai_mai_n40_), .Y(mai_mai_n1228_));
  AO220      m1200(.A0(mai_mai_n1228_), .A1(mai_mai_n607_), .B0(mai_mai_n1227_), .B1(mai_mai_n686_), .Y(mai_mai_n1229_));
  NA2        m1201(.A(mai_mai_n1229_), .B(mai_mai_n330_), .Y(mai_mai_n1230_));
  INV        m1202(.A(mai_mai_n130_), .Y(mai_mai_n1231_));
  NO3        m1203(.A(mai_mai_n1058_), .B(mai_mai_n170_), .C(mai_mai_n83_), .Y(mai_mai_n1232_));
  AOI220     m1204(.A0(mai_mai_n1232_), .A1(mai_mai_n1231_), .B0(mai_mai_n1220_), .B1(mai_mai_n943_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n1233_), .B(mai_mai_n1230_), .Y(mai_mai_n1234_));
  NO2        m1206(.A(mai_mai_n598_), .B(mai_mai_n597_), .Y(mai_mai_n1235_));
  NO4        m1207(.A(mai_mai_n1058_), .B(mai_mai_n1235_), .C(mai_mai_n168_), .D(mai_mai_n83_), .Y(mai_mai_n1236_));
  NO3        m1208(.A(mai_mai_n1236_), .B(mai_mai_n1234_), .C(mai_mai_n618_), .Y(mai_mai_n1237_));
  NA4        m1209(.A(mai_mai_n1237_), .B(mai_mai_n1226_), .C(mai_mai_n1209_), .D(mai_mai_n1193_), .Y(mai06));
  NO2        m1210(.A(mai_mai_n218_), .B(mai_mai_n97_), .Y(mai_mai_n1239_));
  OAI210     m1211(.A0(mai_mai_n1239_), .A1(mai_mai_n1232_), .B0(mai_mai_n373_), .Y(mai_mai_n1240_));
  NO2        m1212(.A(mai_mai_n585_), .B(mai_mai_n783_), .Y(mai_mai_n1241_));
  OR2        m1213(.A(mai_mai_n1241_), .B(mai_mai_n861_), .Y(mai_mai_n1242_));
  NA3        m1214(.A(mai_mai_n1242_), .B(mai_mai_n1240_), .C(mai_mai_n1218_), .Y(mai_mai_n1243_));
  NO3        m1215(.A(mai_mai_n1243_), .B(mai_mai_n1222_), .C(mai_mai_n251_), .Y(mai_mai_n1244_));
  NO2        m1216(.A(mai_mai_n290_), .B(mai_mai_n44_), .Y(mai_mai_n1245_));
  AOI210     m1217(.A0(mai_mai_n1245_), .A1(mai_mai_n944_), .B0(mai_mai_n1216_), .Y(mai_mai_n1246_));
  AOI210     m1218(.A0(mai_mai_n1245_), .A1(mai_mai_n548_), .B0(mai_mai_n1229_), .Y(mai_mai_n1247_));
  AOI210     m1219(.A0(mai_mai_n1247_), .A1(mai_mai_n1246_), .B0(mai_mai_n327_), .Y(mai_mai_n1248_));
  INV        m1220(.A(mai_mai_n652_), .Y(mai_mai_n1249_));
  NA2        m1221(.A(mai_mai_n1249_), .B(mai_mai_n622_), .Y(mai_mai_n1250_));
  NO2        m1222(.A(mai_mai_n507_), .B(mai_mai_n165_), .Y(mai_mai_n1251_));
  NOi21      m1223(.An(mai_mai_n132_), .B(mai_mai_n44_), .Y(mai_mai_n1252_));
  NO2        m1224(.A(mai_mai_n591_), .B(mai_mai_n1078_), .Y(mai_mai_n1253_));
  OAI210     m1225(.A0(mai_mai_n449_), .A1(mai_mai_n242_), .B0(mai_mai_n879_), .Y(mai_mai_n1254_));
  NO4        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1253_), .C(mai_mai_n1252_), .D(mai_mai_n1251_), .Y(mai_mai_n1255_));
  INV        m1227(.A(mai_mai_n584_), .Y(mai_mai_n1256_));
  NA3        m1228(.A(mai_mai_n1256_), .B(mai_mai_n1255_), .C(mai_mai_n1250_), .Y(mai_mai_n1257_));
  NO2        m1229(.A(mai_mai_n724_), .B(mai_mai_n358_), .Y(mai_mai_n1258_));
  AN2        m1230(.A(mai_mai_n925_), .B(mai_mai_n625_), .Y(mai_mai_n1259_));
  NO3        m1231(.A(mai_mai_n1259_), .B(mai_mai_n1257_), .C(mai_mai_n1248_), .Y(mai_mai_n1260_));
  NO2        m1232(.A(mai_mai_n778_), .B(mai_mai_n270_), .Y(mai_mai_n1261_));
  OAI220     m1233(.A0(mai_mai_n711_), .A1(mai_mai_n46_), .B0(mai_mai_n218_), .B1(mai_mai_n600_), .Y(mai_mai_n1262_));
  OAI210     m1234(.A0(mai_mai_n270_), .A1(c), .B0(mai_mai_n621_), .Y(mai_mai_n1263_));
  AOI220     m1235(.A0(mai_mai_n1263_), .A1(mai_mai_n1262_), .B0(mai_mai_n1261_), .B1(mai_mai_n261_), .Y(mai_mai_n1264_));
  OAI220     m1236(.A0(mai_mai_n679_), .A1(mai_mai_n242_), .B0(mai_mai_n503_), .B1(mai_mai_n507_), .Y(mai_mai_n1265_));
  OAI210     m1237(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1266_));
  NO3        m1238(.A(mai_mai_n1266_), .B(mai_mai_n583_), .C(j), .Y(mai_mai_n1267_));
  NOi21      m1239(.An(mai_mai_n1267_), .B(mai_mai_n648_), .Y(mai_mai_n1268_));
  NO3        m1240(.A(mai_mai_n1268_), .B(mai_mai_n1265_), .C(mai_mai_n1081_), .Y(mai_mai_n1269_));
  NA4        m1241(.A(mai_mai_n770_), .B(mai_mai_n769_), .C(mai_mai_n423_), .D(mai_mai_n854_), .Y(mai_mai_n1270_));
  NAi31      m1242(.An(mai_mai_n724_), .B(mai_mai_n1270_), .C(mai_mai_n198_), .Y(mai_mai_n1271_));
  NA4        m1243(.A(mai_mai_n1271_), .B(mai_mai_n1269_), .C(mai_mai_n1264_), .D(mai_mai_n1167_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n453_), .B(mai_mai_n386_), .Y(mai_mai_n1273_));
  OR3        m1245(.A(mai_mai_n1273_), .B(mai_mai_n759_), .C(mai_mai_n531_), .Y(mai_mai_n1274_));
  NA2        m1246(.A(mai_mai_n1267_), .B(mai_mai_n766_), .Y(mai_mai_n1275_));
  NA2        m1247(.A(mai_mai_n1275_), .B(mai_mai_n1274_), .Y(mai_mai_n1276_));
  NA2        m1248(.A(mai_mai_n1258_), .B(mai_mai_n733_), .Y(mai_mai_n1277_));
  AN2        m1249(.A(mai_mai_n898_), .B(mai_mai_n897_), .Y(mai_mai_n1278_));
  NO4        m1250(.A(mai_mai_n1278_), .B(mai_mai_n852_), .C(mai_mai_n492_), .D(mai_mai_n470_), .Y(mai_mai_n1279_));
  NA3        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1277_), .C(mai_mai_n1224_), .Y(mai_mai_n1280_));
  NAi21      m1252(.An(j), .B(i), .Y(mai_mai_n1281_));
  NO4        m1253(.A(mai_mai_n1235_), .B(mai_mai_n1281_), .C(mai_mai_n429_), .D(mai_mai_n228_), .Y(mai_mai_n1282_));
  NO4        m1254(.A(mai_mai_n1282_), .B(mai_mai_n1280_), .C(mai_mai_n1276_), .D(mai_mai_n1272_), .Y(mai_mai_n1283_));
  NA4        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1260_), .C(mai_mai_n1244_), .D(mai_mai_n1237_), .Y(mai07));
  NOi21      m1256(.An(j), .B(k), .Y(mai_mai_n1285_));
  NA4        m1257(.A(mai_mai_n173_), .B(mai_mai_n103_), .C(mai_mai_n1285_), .D(f), .Y(mai_mai_n1286_));
  NAi32      m1258(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1287_));
  NO3        m1259(.A(mai_mai_n1287_), .B(g), .C(f), .Y(mai_mai_n1288_));
  OAI210     m1260(.A0(mai_mai_n310_), .A1(mai_mai_n472_), .B0(mai_mai_n1288_), .Y(mai_mai_n1289_));
  NAi21      m1261(.An(f), .B(c), .Y(mai_mai_n1290_));
  OR2        m1262(.A(e), .B(d), .Y(mai_mai_n1291_));
  OAI220     m1263(.A0(mai_mai_n1291_), .A1(mai_mai_n1290_), .B0(mai_mai_n612_), .B1(mai_mai_n312_), .Y(mai_mai_n1292_));
  NA3        m1264(.A(mai_mai_n1292_), .B(mai_mai_n1022_), .C(mai_mai_n173_), .Y(mai_mai_n1293_));
  NOi31      m1265(.An(n), .B(m), .C(b), .Y(mai_mai_n1294_));
  NO3        m1266(.A(mai_mai_n127_), .B(mai_mai_n437_), .C(h), .Y(mai_mai_n1295_));
  NA3        m1267(.A(mai_mai_n1293_), .B(mai_mai_n1289_), .C(mai_mai_n1286_), .Y(mai_mai_n1296_));
  NOi41      m1268(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1297_));
  NA3        m1269(.A(mai_mai_n1297_), .B(mai_mai_n844_), .C(mai_mai_n401_), .Y(mai_mai_n1298_));
  NOi21      m1270(.An(h), .B(k), .Y(mai_mai_n1299_));
  NO2        m1271(.A(mai_mai_n1298_), .B(mai_mai_n54_), .Y(mai_mai_n1300_));
  NO2        m1272(.A(k), .B(i), .Y(mai_mai_n1301_));
  NA3        m1273(.A(mai_mai_n1301_), .B(mai_mai_n871_), .C(mai_mai_n173_), .Y(mai_mai_n1302_));
  NA2        m1274(.A(mai_mai_n83_), .B(mai_mai_n44_), .Y(mai_mai_n1303_));
  NO2        m1275(.A(mai_mai_n1016_), .B(mai_mai_n429_), .Y(mai_mai_n1304_));
  NA3        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1303_), .C(mai_mai_n207_), .Y(mai_mai_n1305_));
  NO2        m1277(.A(mai_mai_n1030_), .B(mai_mai_n296_), .Y(mai_mai_n1306_));
  NA2        m1278(.A(mai_mai_n532_), .B(mai_mai_n76_), .Y(mai_mai_n1307_));
  NA2        m1279(.A(mai_mai_n1168_), .B(mai_mai_n280_), .Y(mai_mai_n1308_));
  NA4        m1280(.A(mai_mai_n1308_), .B(mai_mai_n1307_), .C(mai_mai_n1305_), .D(mai_mai_n1302_), .Y(mai_mai_n1309_));
  NO3        m1281(.A(mai_mai_n1309_), .B(mai_mai_n1300_), .C(mai_mai_n1296_), .Y(mai_mai_n1310_));
  NO3        m1282(.A(e), .B(d), .C(c), .Y(mai_mai_n1311_));
  OAI210     m1283(.A0(mai_mai_n127_), .A1(mai_mai_n207_), .B0(mai_mai_n589_), .Y(mai_mai_n1312_));
  NA2        m1284(.A(mai_mai_n1312_), .B(mai_mai_n1311_), .Y(mai_mai_n1313_));
  INV        m1285(.A(mai_mai_n1313_), .Y(mai_mai_n1314_));
  OR2        m1286(.A(h), .B(f), .Y(mai_mai_n1315_));
  NO3        m1287(.A(n), .B(m), .C(i), .Y(mai_mai_n1316_));
  OAI210     m1288(.A0(mai_mai_n1079_), .A1(mai_mai_n151_), .B0(mai_mai_n1316_), .Y(mai_mai_n1317_));
  NO2        m1289(.A(mai_mai_n1317_), .B(mai_mai_n1315_), .Y(mai_mai_n1318_));
  NA3        m1290(.A(mai_mai_n676_), .B(mai_mai_n662_), .C(mai_mai_n107_), .Y(mai_mai_n1319_));
  NA3        m1291(.A(mai_mai_n1294_), .B(mai_mai_n1025_), .C(mai_mai_n650_), .Y(mai_mai_n1320_));
  AOI210     m1292(.A0(mai_mai_n1320_), .A1(mai_mai_n1319_), .B0(mai_mai_n44_), .Y(mai_mai_n1321_));
  NA2        m1293(.A(mai_mai_n1316_), .B(mai_mai_n620_), .Y(mai_mai_n1322_));
  NO2        m1294(.A(l), .B(k), .Y(mai_mai_n1323_));
  NOi41      m1295(.An(mai_mai_n537_), .B(mai_mai_n1323_), .C(mai_mai_n465_), .D(mai_mai_n429_), .Y(mai_mai_n1324_));
  NO3        m1296(.A(mai_mai_n429_), .B(d), .C(c), .Y(mai_mai_n1325_));
  NO4        m1297(.A(mai_mai_n1324_), .B(mai_mai_n1321_), .C(mai_mai_n1318_), .D(mai_mai_n1314_), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n141_), .B(h), .Y(mai_mai_n1327_));
  NO2        m1299(.A(mai_mai_n1040_), .B(l), .Y(mai_mai_n1328_));
  NO2        m1300(.A(g), .B(c), .Y(mai_mai_n1329_));
  NA3        m1301(.A(mai_mai_n1329_), .B(mai_mai_n137_), .C(mai_mai_n181_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n1330_), .B(mai_mai_n1328_), .Y(mai_mai_n1331_));
  NA2        m1303(.A(mai_mai_n1331_), .B(mai_mai_n173_), .Y(mai_mai_n1332_));
  NA2        m1304(.A(mai_mai_n1299_), .B(mai_mai_n1040_), .Y(mai_mai_n1333_));
  NO2        m1305(.A(mai_mai_n440_), .B(a), .Y(mai_mai_n1334_));
  NA3        m1306(.A(mai_mai_n1334_), .B(mai_mai_n1333_), .C(mai_mai_n108_), .Y(mai_mai_n1335_));
  NO2        m1307(.A(i), .B(h), .Y(mai_mai_n1336_));
  NA2        m1308(.A(mai_mai_n1336_), .B(mai_mai_n214_), .Y(mai_mai_n1337_));
  AOI210     m1309(.A0(mai_mai_n1103_), .A1(h), .B0(mai_mai_n403_), .Y(mai_mai_n1338_));
  NA2        m1310(.A(mai_mai_n134_), .B(mai_mai_n214_), .Y(mai_mai_n1339_));
  AOI210     m1311(.A0(mai_mai_n252_), .A1(mai_mai_n111_), .B0(mai_mai_n522_), .Y(mai_mai_n1340_));
  OAI220     m1312(.A0(mai_mai_n1340_), .A1(mai_mai_n1337_), .B0(mai_mai_n1339_), .B1(mai_mai_n1338_), .Y(mai_mai_n1341_));
  NO2        m1313(.A(mai_mai_n731_), .B(mai_mai_n182_), .Y(mai_mai_n1342_));
  NOi31      m1314(.An(m), .B(n), .C(b), .Y(mai_mai_n1343_));
  NOi31      m1315(.An(f), .B(d), .C(c), .Y(mai_mai_n1344_));
  NA2        m1316(.A(mai_mai_n1344_), .B(mai_mai_n1343_), .Y(mai_mai_n1345_));
  INV        m1317(.A(mai_mai_n1345_), .Y(mai_mai_n1346_));
  NO3        m1318(.A(mai_mai_n1346_), .B(mai_mai_n1342_), .C(mai_mai_n1341_), .Y(mai_mai_n1347_));
  NA2        m1319(.A(mai_mai_n1051_), .B(mai_mai_n456_), .Y(mai_mai_n1348_));
  NO4        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1025_), .C(mai_mai_n429_), .D(mai_mai_n44_), .Y(mai_mai_n1349_));
  OAI210     m1321(.A0(mai_mai_n176_), .A1(mai_mai_n518_), .B0(mai_mai_n1026_), .Y(mai_mai_n1350_));
  NO3        m1322(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1351_));
  INV        m1323(.A(mai_mai_n1350_), .Y(mai_mai_n1352_));
  NO2        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1349_), .Y(mai_mai_n1353_));
  AN4        m1325(.A(mai_mai_n1353_), .B(mai_mai_n1347_), .C(mai_mai_n1335_), .D(mai_mai_n1332_), .Y(mai_mai_n1354_));
  NA2        m1326(.A(mai_mai_n1294_), .B(mai_mai_n370_), .Y(mai_mai_n1355_));
  NO2        m1327(.A(mai_mai_n1355_), .B(mai_mai_n1007_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n182_), .B(b), .Y(mai_mai_n1357_));
  AOI220     m1329(.A0(mai_mai_n1127_), .A1(mai_mai_n1357_), .B0(mai_mai_n1059_), .B1(mai_mai_n1348_), .Y(mai_mai_n1358_));
  NAi21      m1330(.An(mai_mai_n1356_), .B(mai_mai_n1358_), .Y(mai_mai_n1359_));
  NO4        m1331(.A(mai_mai_n127_), .B(g), .C(f), .D(e), .Y(mai_mai_n1360_));
  NA3        m1332(.A(mai_mai_n1301_), .B(mai_mai_n281_), .C(h), .Y(mai_mai_n1361_));
  OR2        m1333(.A(e), .B(a), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1291_), .B(mai_mai_n1290_), .Y(mai_mai_n1363_));
  AOI210     m1335(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1363_), .Y(mai_mai_n1364_));
  NO2        m1336(.A(mai_mai_n1364_), .B(mai_mai_n1047_), .Y(mai_mai_n1365_));
  NA2        m1337(.A(mai_mai_n1297_), .B(mai_mai_n1323_), .Y(mai_mai_n1366_));
  INV        m1338(.A(mai_mai_n1366_), .Y(mai_mai_n1367_));
  OR3        m1339(.A(mai_mai_n531_), .B(mai_mai_n530_), .C(mai_mai_n107_), .Y(mai_mai_n1368_));
  NA2        m1340(.A(mai_mai_n1077_), .B(mai_mai_n398_), .Y(mai_mai_n1369_));
  OAI220     m1341(.A0(mai_mai_n1369_), .A1(mai_mai_n422_), .B0(mai_mai_n1368_), .B1(mai_mai_n290_), .Y(mai_mai_n1370_));
  AO210      m1342(.A0(mai_mai_n1370_), .A1(mai_mai_n111_), .B0(mai_mai_n1367_), .Y(mai_mai_n1371_));
  NO3        m1343(.A(mai_mai_n1371_), .B(mai_mai_n1365_), .C(mai_mai_n1359_), .Y(mai_mai_n1372_));
  NA4        m1344(.A(mai_mai_n1372_), .B(mai_mai_n1354_), .C(mai_mai_n1326_), .D(mai_mai_n1310_), .Y(mai_mai_n1373_));
  NO2        m1345(.A(mai_mai_n1093_), .B(mai_mai_n105_), .Y(mai_mai_n1374_));
  NA2        m1346(.A(mai_mai_n370_), .B(mai_mai_n54_), .Y(mai_mai_n1375_));
  AOI210     m1347(.A0(mai_mai_n1375_), .A1(mai_mai_n1016_), .B0(mai_mai_n1322_), .Y(mai_mai_n1376_));
  NA2        m1348(.A(mai_mai_n208_), .B(mai_mai_n173_), .Y(mai_mai_n1377_));
  AOI210     m1349(.A0(mai_mai_n1377_), .A1(mai_mai_n1145_), .B0(mai_mai_n1375_), .Y(mai_mai_n1378_));
  NO2        m1350(.A(mai_mai_n1052_), .B(mai_mai_n1047_), .Y(mai_mai_n1379_));
  NO3        m1351(.A(mai_mai_n1379_), .B(mai_mai_n1378_), .C(mai_mai_n1376_), .Y(mai_mai_n1380_));
  NO2        m1352(.A(mai_mai_n382_), .B(j), .Y(mai_mai_n1381_));
  NA3        m1353(.A(mai_mai_n1351_), .B(mai_mai_n1291_), .C(mai_mai_n1077_), .Y(mai_mai_n1382_));
  NAi41      m1354(.An(mai_mai_n1336_), .B(mai_mai_n1038_), .C(mai_mai_n161_), .D(mai_mai_n144_), .Y(mai_mai_n1383_));
  NA2        m1355(.A(mai_mai_n1383_), .B(mai_mai_n1382_), .Y(mai_mai_n1384_));
  NA3        m1356(.A(g), .B(mai_mai_n1381_), .C(mai_mai_n153_), .Y(mai_mai_n1385_));
  INV        m1357(.A(mai_mai_n1385_), .Y(mai_mai_n1386_));
  NO2        m1358(.A(mai_mai_n724_), .B(mai_mai_n168_), .Y(mai_mai_n1387_));
  NO3        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1386_), .C(mai_mai_n1384_), .Y(mai_mai_n1388_));
  NO3        m1360(.A(mai_mai_n1047_), .B(mai_mai_n571_), .C(g), .Y(mai_mai_n1389_));
  NOi21      m1361(.An(mai_mai_n1377_), .B(mai_mai_n1389_), .Y(mai_mai_n1390_));
  NO2        m1362(.A(mai_mai_n1390_), .B(mai_mai_n1016_), .Y(mai_mai_n1391_));
  OR2        m1363(.A(n), .B(i), .Y(mai_mai_n1392_));
  OAI210     m1364(.A0(mai_mai_n1392_), .A1(mai_mai_n1037_), .B0(mai_mai_n47_), .Y(mai_mai_n1393_));
  AOI220     m1365(.A0(mai_mai_n1393_), .A1(mai_mai_n1135_), .B0(mai_mai_n798_), .B1(mai_mai_n189_), .Y(mai_mai_n1394_));
  INV        m1366(.A(mai_mai_n1394_), .Y(mai_mai_n1395_));
  OAI220     m1367(.A0(mai_mai_n646_), .A1(g), .B0(mai_mai_n218_), .B1(c), .Y(mai_mai_n1396_));
  AOI210     m1368(.A0(mai_mai_n1357_), .A1(mai_mai_n41_), .B0(mai_mai_n1396_), .Y(mai_mai_n1397_));
  NO2        m1369(.A(mai_mai_n127_), .B(l), .Y(mai_mai_n1398_));
  NO2        m1370(.A(mai_mai_n218_), .B(k), .Y(mai_mai_n1399_));
  OAI210     m1371(.A0(mai_mai_n1399_), .A1(mai_mai_n1336_), .B0(mai_mai_n1398_), .Y(mai_mai_n1400_));
  OAI220     m1372(.A0(mai_mai_n1400_), .A1(mai_mai_n31_), .B0(mai_mai_n1397_), .B1(mai_mai_n170_), .Y(mai_mai_n1401_));
  NO3        m1373(.A(mai_mai_n1368_), .B(mai_mai_n456_), .C(mai_mai_n344_), .Y(mai_mai_n1402_));
  NO4        m1374(.A(mai_mai_n1402_), .B(mai_mai_n1401_), .C(mai_mai_n1395_), .D(mai_mai_n1391_), .Y(mai_mai_n1403_));
  NO3        m1375(.A(mai_mai_n1062_), .B(mai_mai_n1291_), .C(mai_mai_n47_), .Y(mai_mai_n1404_));
  NO2        m1376(.A(mai_mai_n1047_), .B(h), .Y(mai_mai_n1405_));
  NA3        m1377(.A(mai_mai_n1405_), .B(d), .C(mai_mai_n1008_), .Y(mai_mai_n1406_));
  NO2        m1378(.A(mai_mai_n1406_), .B(c), .Y(mai_mai_n1407_));
  NA3        m1379(.A(mai_mai_n1374_), .B(mai_mai_n456_), .C(f), .Y(mai_mai_n1408_));
  NA2        m1380(.A(mai_mai_n173_), .B(mai_mai_n107_), .Y(mai_mai_n1409_));
  NO2        m1381(.A(mai_mai_n1285_), .B(mai_mai_n42_), .Y(mai_mai_n1410_));
  AOI210     m1382(.A0(mai_mai_n108_), .A1(mai_mai_n40_), .B0(mai_mai_n1410_), .Y(mai_mai_n1411_));
  NO2        m1383(.A(mai_mai_n1411_), .B(mai_mai_n1408_), .Y(mai_mai_n1412_));
  NOi21      m1384(.An(d), .B(f), .Y(mai_mai_n1413_));
  NO2        m1385(.A(mai_mai_n1291_), .B(f), .Y(mai_mai_n1414_));
  NA2        m1386(.A(mai_mai_n1334_), .B(mai_mai_n1410_), .Y(mai_mai_n1415_));
  INV        m1387(.A(mai_mai_n1415_), .Y(mai_mai_n1416_));
  NO3        m1388(.A(mai_mai_n1416_), .B(mai_mai_n1412_), .C(mai_mai_n1407_), .Y(mai_mai_n1417_));
  NA4        m1389(.A(mai_mai_n1417_), .B(mai_mai_n1403_), .C(mai_mai_n1388_), .D(mai_mai_n1380_), .Y(mai_mai_n1418_));
  NO3        m1390(.A(mai_mai_n1051_), .B(mai_mai_n1037_), .C(mai_mai_n40_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n456_), .B(mai_mai_n290_), .Y(mai_mai_n1420_));
  OAI210     m1392(.A0(mai_mai_n1420_), .A1(mai_mai_n1419_), .B0(mai_mai_n1306_), .Y(mai_mai_n1421_));
  OAI210     m1393(.A0(mai_mai_n1360_), .A1(mai_mai_n1294_), .B0(mai_mai_n858_), .Y(mai_mai_n1422_));
  NO2        m1394(.A(mai_mai_n1004_), .B(mai_mai_n127_), .Y(mai_mai_n1423_));
  NA2        m1395(.A(mai_mai_n1423_), .B(mai_mai_n606_), .Y(mai_mai_n1424_));
  NA3        m1396(.A(mai_mai_n1424_), .B(mai_mai_n1422_), .C(mai_mai_n1421_), .Y(mai_mai_n1425_));
  NA2        m1397(.A(mai_mai_n1329_), .B(mai_mai_n1413_), .Y(mai_mai_n1426_));
  NO2        m1398(.A(mai_mai_n1426_), .B(m), .Y(mai_mai_n1427_));
  NA3        m1399(.A(mai_mai_n1060_), .B(mai_mai_n103_), .C(mai_mai_n214_), .Y(mai_mai_n1428_));
  NO2        m1400(.A(mai_mai_n145_), .B(mai_mai_n175_), .Y(mai_mai_n1429_));
  OAI210     m1401(.A0(mai_mai_n1429_), .A1(mai_mai_n105_), .B0(mai_mai_n1343_), .Y(mai_mai_n1430_));
  NA2        m1402(.A(mai_mai_n1430_), .B(mai_mai_n1428_), .Y(mai_mai_n1431_));
  NO3        m1403(.A(mai_mai_n1431_), .B(mai_mai_n1427_), .C(mai_mai_n1425_), .Y(mai_mai_n1432_));
  NO2        m1404(.A(mai_mai_n1290_), .B(e), .Y(mai_mai_n1433_));
  NA2        m1405(.A(mai_mai_n1433_), .B(mai_mai_n396_), .Y(mai_mai_n1434_));
  NA2        m1406(.A(mai_mai_n1088_), .B(mai_mai_n614_), .Y(mai_mai_n1435_));
  OR3        m1407(.A(mai_mai_n1399_), .B(mai_mai_n1168_), .C(mai_mai_n127_), .Y(mai_mai_n1436_));
  OAI220     m1408(.A0(mai_mai_n1436_), .A1(mai_mai_n1434_), .B0(mai_mai_n1435_), .B1(mai_mai_n431_), .Y(mai_mai_n1437_));
  NO3        m1409(.A(mai_mai_n1368_), .B(mai_mai_n344_), .C(a), .Y(mai_mai_n1438_));
  NO2        m1410(.A(mai_mai_n1438_), .B(mai_mai_n1437_), .Y(mai_mai_n1439_));
  NO2        m1411(.A(mai_mai_n175_), .B(c), .Y(mai_mai_n1440_));
  OAI210     m1412(.A0(mai_mai_n1440_), .A1(mai_mai_n1433_), .B0(mai_mai_n173_), .Y(mai_mai_n1441_));
  AOI220     m1413(.A0(mai_mai_n1441_), .A1(mai_mai_n1039_), .B0(mai_mai_n524_), .B1(mai_mai_n358_), .Y(mai_mai_n1442_));
  AOI210     m1414(.A0(i), .A1(mai_mai_n1325_), .B0(mai_mai_n1404_), .Y(mai_mai_n1443_));
  NO2        m1415(.A(mai_mai_n1362_), .B(f), .Y(mai_mai_n1444_));
  AOI210     m1416(.A0(mai_mai_n1088_), .A1(a), .B0(mai_mai_n1444_), .Y(mai_mai_n1445_));
  OAI220     m1417(.A0(mai_mai_n1445_), .A1(mai_mai_n64_), .B0(mai_mai_n1443_), .B1(mai_mai_n206_), .Y(mai_mai_n1446_));
  AOI210     m1418(.A0(mai_mai_n874_), .A1(mai_mai_n405_), .B0(mai_mai_n99_), .Y(mai_mai_n1447_));
  OR2        m1419(.A(mai_mai_n1447_), .B(mai_mai_n530_), .Y(mai_mai_n1448_));
  NA2        m1420(.A(mai_mai_n1444_), .B(mai_mai_n1303_), .Y(mai_mai_n1449_));
  OAI220     m1421(.A0(mai_mai_n1449_), .A1(mai_mai_n47_), .B0(mai_mai_n1448_), .B1(mai_mai_n168_), .Y(mai_mai_n1450_));
  NA4        m1422(.A(mai_mai_n1060_), .B(mai_mai_n1057_), .C(mai_mai_n214_), .D(mai_mai_n63_), .Y(mai_mai_n1451_));
  NA2        m1423(.A(mai_mai_n1295_), .B(mai_mai_n176_), .Y(mai_mai_n1452_));
  NO2        m1424(.A(mai_mai_n47_), .B(l), .Y(mai_mai_n1453_));
  OAI210     m1425(.A0(mai_mai_n1362_), .A1(mai_mai_n836_), .B0(mai_mai_n472_), .Y(mai_mai_n1454_));
  OAI210     m1426(.A0(mai_mai_n1454_), .A1(mai_mai_n1063_), .B0(mai_mai_n1453_), .Y(mai_mai_n1455_));
  NO2        m1427(.A(mai_mai_n247_), .B(g), .Y(mai_mai_n1456_));
  NO2        m1428(.A(m), .B(i), .Y(mai_mai_n1457_));
  BUFFER     m1429(.A(mai_mai_n1457_), .Y(mai_mai_n1458_));
  AOI220     m1430(.A0(mai_mai_n1458_), .A1(mai_mai_n1327_), .B0(mai_mai_n1038_), .B1(mai_mai_n1456_), .Y(mai_mai_n1459_));
  NA4        m1431(.A(mai_mai_n1459_), .B(mai_mai_n1455_), .C(mai_mai_n1452_), .D(mai_mai_n1451_), .Y(mai_mai_n1460_));
  NO4        m1432(.A(mai_mai_n1460_), .B(mai_mai_n1450_), .C(mai_mai_n1446_), .D(mai_mai_n1442_), .Y(mai_mai_n1461_));
  NA3        m1433(.A(mai_mai_n1461_), .B(mai_mai_n1439_), .C(mai_mai_n1432_), .Y(mai_mai_n1462_));
  NA3        m1434(.A(mai_mai_n931_), .B(mai_mai_n134_), .C(mai_mai_n45_), .Y(mai_mai_n1463_));
  AOI210     m1435(.A0(mai_mai_n142_), .A1(c), .B0(mai_mai_n1463_), .Y(mai_mai_n1464_));
  INV        m1436(.A(mai_mai_n179_), .Y(mai_mai_n1465_));
  NA2        m1437(.A(mai_mai_n1465_), .B(mai_mai_n1405_), .Y(mai_mai_n1466_));
  OR2        m1438(.A(mai_mai_n128_), .B(mai_mai_n1355_), .Y(mai_mai_n1467_));
  NA2        m1439(.A(mai_mai_n1467_), .B(mai_mai_n1466_), .Y(mai_mai_n1468_));
  NO2        m1440(.A(mai_mai_n1468_), .B(mai_mai_n1464_), .Y(mai_mai_n1469_));
  AOI210     m1441(.A0(mai_mai_n151_), .A1(mai_mai_n54_), .B0(mai_mai_n1433_), .Y(mai_mai_n1470_));
  NO2        m1442(.A(mai_mai_n1470_), .B(mai_mai_n1409_), .Y(mai_mai_n1471_));
  INV        m1443(.A(mai_mai_n1471_), .Y(mai_mai_n1472_));
  AN2        m1444(.A(mai_mai_n1060_), .B(mai_mai_n1045_), .Y(mai_mai_n1473_));
  NA2        m1445(.A(mai_mai_n1473_), .B(mai_mai_n1127_), .Y(mai_mai_n1474_));
  NO2        m1446(.A(mai_mai_n1408_), .B(mai_mai_n64_), .Y(mai_mai_n1475_));
  NA2        m1447(.A(mai_mai_n57_), .B(a), .Y(mai_mai_n1476_));
  NO2        m1448(.A(mai_mai_n1301_), .B(mai_mai_n113_), .Y(mai_mai_n1477_));
  OAI220     m1449(.A0(mai_mai_n1477_), .A1(mai_mai_n1355_), .B0(mai_mai_n1369_), .B1(mai_mai_n1476_), .Y(mai_mai_n1478_));
  NO2        m1450(.A(mai_mai_n1478_), .B(mai_mai_n1475_), .Y(mai_mai_n1479_));
  NA4        m1451(.A(mai_mai_n1479_), .B(mai_mai_n1474_), .C(mai_mai_n1472_), .D(mai_mai_n1469_), .Y(mai_mai_n1480_));
  OR4        m1452(.A(mai_mai_n1480_), .B(mai_mai_n1462_), .C(mai_mai_n1418_), .D(mai_mai_n1373_), .Y(mai04));
  NOi31      m1453(.An(mai_mai_n1360_), .B(mai_mai_n1361_), .C(mai_mai_n1010_), .Y(mai_mai_n1482_));
  NA2        m1454(.A(mai_mai_n1414_), .B(mai_mai_n798_), .Y(mai_mai_n1483_));
  NO3        m1455(.A(mai_mai_n1483_), .B(mai_mai_n999_), .C(mai_mai_n473_), .Y(mai_mai_n1484_));
  OR3        m1456(.A(mai_mai_n1484_), .B(mai_mai_n1482_), .C(mai_mai_n1028_), .Y(mai_mai_n1485_));
  NO3        m1457(.A(mai_mai_n1303_), .B(mai_mai_n86_), .C(k), .Y(mai_mai_n1486_));
  AOI210     m1458(.A0(mai_mai_n1486_), .A1(mai_mai_n1021_), .B0(mai_mai_n1147_), .Y(mai_mai_n1487_));
  NA2        m1459(.A(mai_mai_n1487_), .B(mai_mai_n1172_), .Y(mai_mai_n1488_));
  NO4        m1460(.A(mai_mai_n1488_), .B(mai_mai_n1485_), .C(mai_mai_n1036_), .D(mai_mai_n1015_), .Y(mai_mai_n1489_));
  NA3        m1461(.A(mai_mai_n1489_), .B(mai_mai_n1090_), .C(mai_mai_n1066_), .Y(mai05));
  INV        m1462(.A(mai_mai_n589_), .Y(mai_mai_n1493_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi31      u0013(.An(n), .B(m), .C(l), .Y(men_men_n42_));
  INV        u0014(.A(i), .Y(men_men_n43_));
  AN2        u0015(.A(h), .B(g), .Y(men_men_n44_));
  NA2        u0016(.A(men_men_n44_), .B(men_men_n43_), .Y(men_men_n45_));
  NO2        u0017(.A(men_men_n45_), .B(men_men_n42_), .Y(men_men_n46_));
  NAi21      u0018(.An(n), .B(m), .Y(men_men_n47_));
  NOi32      u0019(.An(k), .Bn(h), .C(l), .Y(men_men_n48_));
  NOi32      u0020(.An(k), .Bn(h), .C(g), .Y(men_men_n49_));
  INV        u0021(.A(men_men_n49_), .Y(men_men_n50_));
  NO2        u0022(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n51_));
  NO3        u0023(.A(men_men_n51_), .B(men_men_n46_), .C(men_men_n39_), .Y(men_men_n52_));
  AOI210     u0024(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n53_));
  INV        u0025(.A(c), .Y(men_men_n54_));
  NA2        u0026(.A(e), .B(b), .Y(men_men_n55_));
  NO2        u0027(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  INV        u0028(.A(d), .Y(men_men_n57_));
  NA3        u0029(.A(g), .B(men_men_n57_), .C(a), .Y(men_men_n58_));
  NAi21      u0030(.An(i), .B(h), .Y(men_men_n59_));
  NAi31      u0031(.An(i), .B(l), .C(j), .Y(men_men_n60_));
  OAI220     u0032(.A0(men_men_n60_), .A1(men_men_n47_), .B0(men_men_n59_), .B1(men_men_n42_), .Y(men_men_n61_));
  NAi31      u0033(.An(men_men_n58_), .B(men_men_n61_), .C(men_men_n56_), .Y(men_men_n62_));
  NAi41      u0034(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n63_));
  NA2        u0035(.A(g), .B(f), .Y(men_men_n64_));
  NO2        u0036(.A(men_men_n64_), .B(men_men_n63_), .Y(men_men_n65_));
  NAi21      u0037(.An(i), .B(j), .Y(men_men_n66_));
  NAi32      u0038(.An(n), .Bn(k), .C(m), .Y(men_men_n67_));
  NO2        u0039(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n68_));
  NAi31      u0040(.An(l), .B(m), .C(k), .Y(men_men_n69_));
  NAi21      u0041(.An(e), .B(h), .Y(men_men_n70_));
  NAi41      u0042(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n71_));
  NA2        u0043(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n72_));
  INV        u0044(.A(m), .Y(men_men_n73_));
  NOi21      u0045(.An(k), .B(l), .Y(men_men_n74_));
  NA2        u0046(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n75_));
  AN4        u0047(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n76_));
  NOi31      u0048(.An(h), .B(g), .C(f), .Y(men_men_n77_));
  NA2        u0049(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NAi32      u0050(.An(m), .Bn(k), .C(j), .Y(men_men_n79_));
  NOi32      u0051(.An(h), .Bn(g), .C(f), .Y(men_men_n80_));
  NA2        u0052(.A(men_men_n80_), .B(men_men_n76_), .Y(men_men_n81_));
  OA220      u0053(.A0(men_men_n81_), .A1(men_men_n79_), .B0(men_men_n78_), .B1(men_men_n75_), .Y(men_men_n82_));
  NA3        u0054(.A(men_men_n82_), .B(men_men_n72_), .C(men_men_n62_), .Y(men_men_n83_));
  INV        u0055(.A(n), .Y(men_men_n84_));
  NOi32      u0056(.An(e), .Bn(b), .C(d), .Y(men_men_n85_));
  NA2        u0057(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n86_));
  INV        u0058(.A(j), .Y(men_men_n87_));
  AN3        u0059(.A(m), .B(k), .C(i), .Y(men_men_n88_));
  NA3        u0060(.A(men_men_n88_), .B(men_men_n87_), .C(g), .Y(men_men_n89_));
  NO2        u0061(.A(men_men_n89_), .B(f), .Y(men_men_n90_));
  NAi32      u0062(.An(g), .Bn(f), .C(h), .Y(men_men_n91_));
  NAi31      u0063(.An(j), .B(m), .C(l), .Y(men_men_n92_));
  NO2        u0064(.A(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  NA2        u0065(.A(m), .B(l), .Y(men_men_n94_));
  NAi31      u0066(.An(k), .B(j), .C(g), .Y(men_men_n95_));
  NO3        u0067(.A(men_men_n95_), .B(men_men_n94_), .C(f), .Y(men_men_n96_));
  AN2        u0068(.A(j), .B(g), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(l), .C(i), .Y(men_men_n98_));
  NOi21      u0070(.An(g), .B(i), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(j), .C(k), .Y(men_men_n100_));
  AOI220     u0072(.A0(men_men_n100_), .A1(men_men_n99_), .B0(men_men_n98_), .B1(men_men_n97_), .Y(men_men_n101_));
  NO2        u0073(.A(men_men_n101_), .B(f), .Y(men_men_n102_));
  NO3        u0074(.A(men_men_n102_), .B(men_men_n96_), .C(men_men_n90_), .Y(men_men_n103_));
  NAi41      u0075(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n104_));
  AN2        u0076(.A(e), .B(b), .Y(men_men_n105_));
  NOi31      u0077(.An(c), .B(h), .C(f), .Y(men_men_n106_));
  NA2        u0078(.A(men_men_n106_), .B(men_men_n105_), .Y(men_men_n107_));
  NO2        u0079(.A(men_men_n107_), .B(men_men_n104_), .Y(men_men_n108_));
  NOi21      u0080(.An(i), .B(h), .Y(men_men_n109_));
  INV        u0081(.A(a), .Y(men_men_n110_));
  NA2        u0082(.A(men_men_n105_), .B(men_men_n110_), .Y(men_men_n111_));
  INV        u0083(.A(l), .Y(men_men_n112_));
  NOi21      u0084(.An(m), .B(n), .Y(men_men_n113_));
  AN2        u0085(.A(k), .B(h), .Y(men_men_n114_));
  INV        u0086(.A(b), .Y(men_men_n115_));
  NA2        u0087(.A(l), .B(j), .Y(men_men_n116_));
  AN2        u0088(.A(k), .B(i), .Y(men_men_n117_));
  NA2        u0089(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u0090(.A(g), .B(e), .Y(men_men_n119_));
  NOi32      u0091(.An(c), .Bn(a), .C(d), .Y(men_men_n120_));
  NA2        u0092(.A(men_men_n120_), .B(men_men_n113_), .Y(men_men_n121_));
  NO4        u0093(.A(men_men_n121_), .B(men_men_n119_), .C(men_men_n118_), .D(men_men_n115_), .Y(men_men_n122_));
  NO2        u0094(.A(men_men_n122_), .B(men_men_n108_), .Y(men_men_n123_));
  OAI210     u0095(.A0(men_men_n103_), .A1(men_men_n86_), .B0(men_men_n123_), .Y(men_men_n124_));
  NOi31      u0096(.An(k), .B(m), .C(j), .Y(men_men_n125_));
  NOi31      u0097(.An(k), .B(m), .C(i), .Y(men_men_n126_));
  NA3        u0098(.A(men_men_n126_), .B(men_men_n80_), .C(men_men_n76_), .Y(men_men_n127_));
  INV        u0099(.A(men_men_n127_), .Y(men_men_n128_));
  NOi32      u0100(.An(f), .Bn(b), .C(e), .Y(men_men_n129_));
  NAi21      u0101(.An(g), .B(h), .Y(men_men_n130_));
  NAi21      u0102(.An(m), .B(n), .Y(men_men_n131_));
  NAi21      u0103(.An(j), .B(k), .Y(men_men_n132_));
  NAi41      u0104(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n133_));
  NAi31      u0105(.An(j), .B(k), .C(h), .Y(men_men_n134_));
  NO2        u0106(.A(k), .B(j), .Y(men_men_n135_));
  NO2        u0107(.A(men_men_n135_), .B(men_men_n131_), .Y(men_men_n136_));
  AN2        u0108(.A(k), .B(j), .Y(men_men_n137_));
  NAi21      u0109(.An(c), .B(b), .Y(men_men_n138_));
  NA2        u0110(.A(f), .B(d), .Y(men_men_n139_));
  NO4        u0111(.A(men_men_n139_), .B(men_men_n138_), .C(men_men_n137_), .D(men_men_n130_), .Y(men_men_n140_));
  NAi31      u0112(.An(f), .B(e), .C(b), .Y(men_men_n141_));
  NA2        u0113(.A(men_men_n140_), .B(men_men_n136_), .Y(men_men_n142_));
  NA2        u0114(.A(d), .B(b), .Y(men_men_n143_));
  NAi21      u0115(.An(e), .B(f), .Y(men_men_n144_));
  NA2        u0116(.A(b), .B(a), .Y(men_men_n145_));
  NAi21      u0117(.An(e), .B(g), .Y(men_men_n146_));
  NAi21      u0118(.An(c), .B(d), .Y(men_men_n147_));
  NAi31      u0119(.An(l), .B(k), .C(h), .Y(men_men_n148_));
  NO2        u0120(.A(men_men_n131_), .B(men_men_n148_), .Y(men_men_n149_));
  NAi21      u0121(.An(men_men_n128_), .B(men_men_n142_), .Y(men_men_n150_));
  NAi31      u0122(.An(e), .B(f), .C(b), .Y(men_men_n151_));
  NO2        u0123(.A(g), .B(men_men_n151_), .Y(men_men_n152_));
  NOi21      u0124(.An(h), .B(i), .Y(men_men_n153_));
  NOi21      u0125(.An(k), .B(m), .Y(men_men_n154_));
  NA3        u0126(.A(men_men_n154_), .B(men_men_n153_), .C(n), .Y(men_men_n155_));
  NOi21      u0127(.An(men_men_n152_), .B(men_men_n155_), .Y(men_men_n156_));
  NOi21      u0128(.An(h), .B(g), .Y(men_men_n157_));
  NO2        u0129(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n158_));
  NA2        u0130(.A(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NAi31      u0131(.An(l), .B(j), .C(h), .Y(men_men_n160_));
  NO2        u0132(.A(men_men_n160_), .B(men_men_n47_), .Y(men_men_n161_));
  NA2        u0133(.A(men_men_n161_), .B(men_men_n65_), .Y(men_men_n162_));
  NOi32      u0134(.An(n), .Bn(k), .C(m), .Y(men_men_n163_));
  NA2        u0135(.A(l), .B(i), .Y(men_men_n164_));
  NA2        u0136(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OAI210     u0137(.A0(men_men_n165_), .A1(men_men_n159_), .B0(men_men_n162_), .Y(men_men_n166_));
  NAi31      u0138(.An(d), .B(f), .C(c), .Y(men_men_n167_));
  NAi31      u0139(.An(e), .B(f), .C(c), .Y(men_men_n168_));
  NA2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  NA2        u0141(.A(j), .B(h), .Y(men_men_n170_));
  OR3        u0142(.A(n), .B(m), .C(k), .Y(men_men_n171_));
  NO2        u0143(.A(men_men_n171_), .B(men_men_n170_), .Y(men_men_n172_));
  NAi32      u0144(.An(m), .Bn(k), .C(n), .Y(men_men_n173_));
  NO2        u0145(.A(men_men_n173_), .B(men_men_n170_), .Y(men_men_n174_));
  AOI220     u0146(.A0(men_men_n174_), .A1(men_men_n152_), .B0(men_men_n172_), .B1(men_men_n169_), .Y(men_men_n175_));
  NO2        u0147(.A(n), .B(m), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n48_), .Y(men_men_n177_));
  NAi21      u0149(.An(f), .B(e), .Y(men_men_n178_));
  NA2        u0150(.A(d), .B(c), .Y(men_men_n179_));
  NAi31      u0151(.An(m), .B(n), .C(b), .Y(men_men_n180_));
  NA2        u0152(.A(k), .B(i), .Y(men_men_n181_));
  NAi21      u0153(.An(h), .B(f), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n180_), .B(men_men_n147_), .Y(men_men_n184_));
  NA2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NOi32      u0157(.An(f), .Bn(c), .C(d), .Y(men_men_n186_));
  NOi32      u0158(.An(f), .Bn(c), .C(e), .Y(men_men_n187_));
  NO2        u0159(.A(men_men_n187_), .B(men_men_n186_), .Y(men_men_n188_));
  NO3        u0160(.A(n), .B(m), .C(j), .Y(men_men_n189_));
  NA2        u0161(.A(men_men_n189_), .B(men_men_n114_), .Y(men_men_n190_));
  AO210      u0162(.A0(men_men_n190_), .A1(men_men_n177_), .B0(men_men_n188_), .Y(men_men_n191_));
  NA3        u0163(.A(men_men_n191_), .B(men_men_n185_), .C(men_men_n175_), .Y(men_men_n192_));
  OR4        u0164(.A(men_men_n192_), .B(men_men_n166_), .C(men_men_n156_), .D(men_men_n150_), .Y(men_men_n193_));
  NO4        u0165(.A(men_men_n193_), .B(men_men_n124_), .C(men_men_n83_), .D(men_men_n53_), .Y(men_men_n194_));
  NA3        u0166(.A(m), .B(men_men_n112_), .C(j), .Y(men_men_n195_));
  NAi31      u0167(.An(n), .B(h), .C(g), .Y(men_men_n196_));
  NO2        u0168(.A(men_men_n196_), .B(men_men_n195_), .Y(men_men_n197_));
  NOi32      u0169(.An(m), .Bn(k), .C(l), .Y(men_men_n198_));
  NA3        u0170(.A(men_men_n198_), .B(men_men_n87_), .C(g), .Y(men_men_n199_));
  NO2        u0171(.A(men_men_n199_), .B(n), .Y(men_men_n200_));
  NOi21      u0172(.An(k), .B(j), .Y(men_men_n201_));
  NA4        u0173(.A(men_men_n201_), .B(men_men_n113_), .C(i), .D(g), .Y(men_men_n202_));
  AN2        u0174(.A(i), .B(g), .Y(men_men_n203_));
  NA3        u0175(.A(men_men_n74_), .B(men_men_n203_), .C(men_men_n113_), .Y(men_men_n204_));
  NA2        u0176(.A(men_men_n204_), .B(men_men_n202_), .Y(men_men_n205_));
  NO3        u0177(.A(men_men_n205_), .B(men_men_n200_), .C(men_men_n197_), .Y(men_men_n206_));
  NAi41      u0178(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n207_));
  INV        u0179(.A(men_men_n207_), .Y(men_men_n208_));
  INV        u0180(.A(f), .Y(men_men_n209_));
  INV        u0181(.A(g), .Y(men_men_n210_));
  NOi31      u0182(.An(i), .B(j), .C(h), .Y(men_men_n211_));
  NOi21      u0183(.An(l), .B(m), .Y(men_men_n212_));
  NA2        u0184(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  NO2        u0185(.A(men_men_n206_), .B(men_men_n32_), .Y(men_men_n214_));
  NOi21      u0186(.An(n), .B(m), .Y(men_men_n215_));
  NOi32      u0187(.An(l), .Bn(i), .C(j), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  OA220      u0189(.A0(men_men_n217_), .A1(men_men_n107_), .B0(men_men_n79_), .B1(men_men_n78_), .Y(men_men_n218_));
  NAi21      u0190(.An(j), .B(h), .Y(men_men_n219_));
  XN2        u0191(.A(i), .B(h), .Y(men_men_n220_));
  NA2        u0192(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n221_));
  NOi31      u0193(.An(k), .B(n), .C(m), .Y(men_men_n222_));
  NOi31      u0194(.An(men_men_n222_), .B(men_men_n179_), .C(men_men_n178_), .Y(men_men_n223_));
  NA2        u0195(.A(men_men_n223_), .B(men_men_n221_), .Y(men_men_n224_));
  NAi31      u0196(.An(f), .B(e), .C(c), .Y(men_men_n225_));
  NO4        u0197(.A(men_men_n225_), .B(men_men_n171_), .C(men_men_n170_), .D(men_men_n57_), .Y(men_men_n226_));
  NA4        u0198(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n227_));
  NAi32      u0199(.An(m), .Bn(i), .C(k), .Y(men_men_n228_));
  NO3        u0200(.A(men_men_n228_), .B(men_men_n91_), .C(men_men_n227_), .Y(men_men_n229_));
  INV        u0201(.A(k), .Y(men_men_n230_));
  NO2        u0202(.A(men_men_n229_), .B(men_men_n226_), .Y(men_men_n231_));
  NAi21      u0203(.An(n), .B(a), .Y(men_men_n232_));
  NO2        u0204(.A(men_men_n232_), .B(men_men_n143_), .Y(men_men_n233_));
  NAi41      u0205(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n234_));
  NO2        u0206(.A(men_men_n234_), .B(e), .Y(men_men_n235_));
  NO3        u0207(.A(men_men_n144_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n236_));
  OAI210     u0208(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n233_), .Y(men_men_n237_));
  AN4        u0209(.A(men_men_n237_), .B(men_men_n231_), .C(men_men_n224_), .D(men_men_n218_), .Y(men_men_n238_));
  OR2        u0210(.A(h), .B(g), .Y(men_men_n239_));
  NO2        u0211(.A(men_men_n239_), .B(men_men_n104_), .Y(men_men_n240_));
  NA2        u0212(.A(men_men_n240_), .B(men_men_n129_), .Y(men_men_n241_));
  NA2        u0213(.A(men_men_n154_), .B(men_men_n109_), .Y(men_men_n242_));
  NO2        u0214(.A(n), .B(a), .Y(men_men_n243_));
  NAi31      u0215(.An(men_men_n234_), .B(men_men_n243_), .C(men_men_n105_), .Y(men_men_n244_));
  NAi21      u0216(.An(h), .B(i), .Y(men_men_n245_));
  NA2        u0217(.A(men_men_n176_), .B(k), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(men_men_n245_), .Y(men_men_n247_));
  NA2        u0219(.A(men_men_n247_), .B(men_men_n186_), .Y(men_men_n248_));
  NA3        u0220(.A(men_men_n248_), .B(men_men_n244_), .C(men_men_n241_), .Y(men_men_n249_));
  NOi21      u0221(.An(g), .B(e), .Y(men_men_n250_));
  NO2        u0222(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n251_));
  NA2        u0223(.A(men_men_n251_), .B(men_men_n250_), .Y(men_men_n252_));
  NOi32      u0224(.An(l), .Bn(j), .C(i), .Y(men_men_n253_));
  AOI210     u0225(.A0(men_men_n74_), .A1(men_men_n87_), .B0(men_men_n253_), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n245_), .B(men_men_n42_), .Y(men_men_n255_));
  NAi21      u0227(.An(f), .B(g), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n63_), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n67_), .B(men_men_n116_), .Y(men_men_n258_));
  AOI220     u0230(.A0(men_men_n258_), .A1(men_men_n257_), .B0(men_men_n255_), .B1(men_men_n65_), .Y(men_men_n259_));
  OAI210     u0231(.A0(men_men_n254_), .A1(men_men_n252_), .B0(men_men_n259_), .Y(men_men_n260_));
  NO3        u0232(.A(men_men_n132_), .B(men_men_n47_), .C(men_men_n43_), .Y(men_men_n261_));
  NOi41      u0233(.An(men_men_n238_), .B(men_men_n260_), .C(men_men_n249_), .D(men_men_n214_), .Y(men_men_n262_));
  NO3        u0234(.A(men_men_n197_), .B(men_men_n46_), .C(men_men_n39_), .Y(men_men_n263_));
  NO2        u0235(.A(men_men_n263_), .B(men_men_n111_), .Y(men_men_n264_));
  NA3        u0236(.A(men_men_n57_), .B(c), .C(b), .Y(men_men_n265_));
  NAi21      u0237(.An(h), .B(g), .Y(men_men_n266_));
  OR4        u0238(.A(men_men_n266_), .B(men_men_n265_), .C(men_men_n217_), .D(e), .Y(men_men_n267_));
  NO2        u0239(.A(men_men_n242_), .B(men_men_n256_), .Y(men_men_n268_));
  NAi31      u0240(.An(g), .B(k), .C(h), .Y(men_men_n269_));
  NO3        u0241(.A(men_men_n131_), .B(men_men_n269_), .C(l), .Y(men_men_n270_));
  NAi31      u0242(.An(e), .B(d), .C(a), .Y(men_men_n271_));
  NA2        u0243(.A(men_men_n270_), .B(men_men_n129_), .Y(men_men_n272_));
  NA2        u0244(.A(men_men_n272_), .B(men_men_n267_), .Y(men_men_n273_));
  NA4        u0245(.A(men_men_n154_), .B(men_men_n80_), .C(men_men_n76_), .D(men_men_n116_), .Y(men_men_n274_));
  NA3        u0246(.A(men_men_n154_), .B(men_men_n153_), .C(men_men_n84_), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n275_), .B(men_men_n188_), .Y(men_men_n276_));
  NOi21      u0248(.An(men_men_n274_), .B(men_men_n276_), .Y(men_men_n277_));
  NA3        u0249(.A(e), .B(c), .C(b), .Y(men_men_n278_));
  NO2        u0250(.A(men_men_n58_), .B(men_men_n278_), .Y(men_men_n279_));
  NAi32      u0251(.An(k), .Bn(i), .C(j), .Y(men_men_n280_));
  NAi31      u0252(.An(h), .B(l), .C(i), .Y(men_men_n281_));
  NA3        u0253(.A(men_men_n281_), .B(men_men_n280_), .C(men_men_n160_), .Y(men_men_n282_));
  NOi21      u0254(.An(men_men_n282_), .B(men_men_n47_), .Y(men_men_n283_));
  OAI210     u0255(.A0(men_men_n257_), .A1(men_men_n279_), .B0(men_men_n283_), .Y(men_men_n284_));
  NAi21      u0256(.An(l), .B(k), .Y(men_men_n285_));
  NO2        u0257(.A(men_men_n285_), .B(men_men_n47_), .Y(men_men_n286_));
  NOi21      u0258(.An(l), .B(j), .Y(men_men_n287_));
  NA2        u0259(.A(men_men_n157_), .B(men_men_n287_), .Y(men_men_n288_));
  NA3        u0260(.A(men_men_n117_), .B(men_men_n116_), .C(g), .Y(men_men_n289_));
  OR3        u0261(.A(men_men_n71_), .B(men_men_n73_), .C(e), .Y(men_men_n290_));
  AOI210     u0262(.A0(men_men_n289_), .A1(men_men_n288_), .B0(men_men_n290_), .Y(men_men_n291_));
  INV        u0263(.A(men_men_n291_), .Y(men_men_n292_));
  NAi32      u0264(.An(j), .Bn(h), .C(i), .Y(men_men_n293_));
  NAi21      u0265(.An(m), .B(l), .Y(men_men_n294_));
  NO3        u0266(.A(men_men_n294_), .B(men_men_n293_), .C(men_men_n84_), .Y(men_men_n295_));
  NA2        u0267(.A(h), .B(g), .Y(men_men_n296_));
  NA2        u0268(.A(men_men_n163_), .B(men_men_n43_), .Y(men_men_n297_));
  NO2        u0269(.A(men_men_n297_), .B(men_men_n296_), .Y(men_men_n298_));
  OAI210     u0270(.A0(men_men_n298_), .A1(men_men_n295_), .B0(men_men_n158_), .Y(men_men_n299_));
  NA4        u0271(.A(men_men_n299_), .B(men_men_n292_), .C(men_men_n284_), .D(men_men_n277_), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n141_), .B(d), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n301_), .B(men_men_n51_), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n107_), .B(men_men_n104_), .Y(men_men_n303_));
  NAi32      u0275(.An(n), .Bn(m), .C(l), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n304_), .B(men_men_n293_), .Y(men_men_n305_));
  NO2        u0277(.A(men_men_n121_), .B(men_men_n115_), .Y(men_men_n306_));
  NAi31      u0278(.An(k), .B(l), .C(j), .Y(men_men_n307_));
  OAI210     u0279(.A0(men_men_n285_), .A1(j), .B0(men_men_n307_), .Y(men_men_n308_));
  NOi21      u0280(.An(men_men_n308_), .B(men_men_n119_), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n309_), .B(men_men_n306_), .Y(men_men_n310_));
  NA2        u0282(.A(men_men_n310_), .B(men_men_n302_), .Y(men_men_n311_));
  NO4        u0283(.A(men_men_n311_), .B(men_men_n300_), .C(men_men_n273_), .D(men_men_n264_), .Y(men_men_n312_));
  NA2        u0284(.A(men_men_n247_), .B(men_men_n187_), .Y(men_men_n313_));
  NAi21      u0285(.An(m), .B(k), .Y(men_men_n314_));
  NO2        u0286(.A(men_men_n220_), .B(men_men_n314_), .Y(men_men_n315_));
  NAi41      u0287(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n316_));
  NO2        u0288(.A(men_men_n316_), .B(men_men_n146_), .Y(men_men_n317_));
  NA2        u0289(.A(men_men_n317_), .B(men_men_n315_), .Y(men_men_n318_));
  NAi31      u0290(.An(i), .B(l), .C(h), .Y(men_men_n319_));
  NA2        u0291(.A(e), .B(c), .Y(men_men_n320_));
  NO3        u0292(.A(men_men_n320_), .B(n), .C(d), .Y(men_men_n321_));
  NOi21      u0293(.An(f), .B(h), .Y(men_men_n322_));
  NA2        u0294(.A(men_men_n322_), .B(men_men_n117_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n323_), .B(men_men_n210_), .Y(men_men_n324_));
  NAi31      u0296(.An(d), .B(e), .C(b), .Y(men_men_n325_));
  NO2        u0297(.A(men_men_n131_), .B(men_men_n325_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n324_), .Y(men_men_n327_));
  NA3        u0299(.A(men_men_n327_), .B(men_men_n318_), .C(men_men_n313_), .Y(men_men_n328_));
  NO4        u0300(.A(men_men_n316_), .B(men_men_n79_), .C(men_men_n70_), .D(men_men_n210_), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n243_), .B(men_men_n105_), .Y(men_men_n330_));
  OR2        u0302(.A(men_men_n330_), .B(men_men_n199_), .Y(men_men_n331_));
  NOi31      u0303(.An(l), .B(n), .C(m), .Y(men_men_n332_));
  NAi21      u0304(.An(men_men_n329_), .B(men_men_n331_), .Y(men_men_n333_));
  NAi32      u0305(.An(m), .Bn(j), .C(k), .Y(men_men_n334_));
  NAi41      u0306(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n335_));
  OAI210     u0307(.A0(men_men_n207_), .A1(men_men_n334_), .B0(men_men_n335_), .Y(men_men_n336_));
  NOi31      u0308(.An(j), .B(m), .C(k), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n125_), .B(men_men_n337_), .Y(men_men_n338_));
  AN3        u0310(.A(h), .B(g), .C(f), .Y(men_men_n339_));
  NAi31      u0311(.An(men_men_n338_), .B(men_men_n339_), .C(men_men_n336_), .Y(men_men_n340_));
  NOi32      u0312(.An(m), .Bn(j), .C(l), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n341_), .B(men_men_n98_), .Y(men_men_n342_));
  NAi32      u0314(.An(men_men_n342_), .Bn(men_men_n196_), .C(men_men_n301_), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n294_), .B(men_men_n293_), .Y(men_men_n344_));
  NO2        u0316(.A(men_men_n213_), .B(g), .Y(men_men_n345_));
  NO2        u0317(.A(men_men_n151_), .B(men_men_n84_), .Y(men_men_n346_));
  NA2        u0318(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n228_), .B(men_men_n79_), .Y(men_men_n348_));
  NA3        u0320(.A(men_men_n348_), .B(men_men_n339_), .C(men_men_n208_), .Y(men_men_n349_));
  NA4        u0321(.A(men_men_n349_), .B(men_men_n347_), .C(men_men_n343_), .D(men_men_n340_), .Y(men_men_n350_));
  NA3        u0322(.A(h), .B(g), .C(f), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n351_), .B(men_men_n75_), .Y(men_men_n352_));
  NA2        u0324(.A(men_men_n335_), .B(men_men_n207_), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n157_), .B(e), .Y(men_men_n354_));
  NO2        u0326(.A(men_men_n354_), .B(men_men_n41_), .Y(men_men_n355_));
  AOI220     u0327(.A0(men_men_n355_), .A1(men_men_n306_), .B0(men_men_n353_), .B1(men_men_n352_), .Y(men_men_n356_));
  NOi32      u0328(.An(j), .Bn(g), .C(i), .Y(men_men_n357_));
  NA3        u0329(.A(men_men_n357_), .B(men_men_n285_), .C(men_men_n113_), .Y(men_men_n358_));
  OR2        u0330(.A(men_men_n111_), .B(men_men_n358_), .Y(men_men_n359_));
  NOi32      u0331(.An(e), .Bn(b), .C(a), .Y(men_men_n360_));
  AN2        u0332(.A(l), .B(j), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n314_), .B(men_men_n361_), .Y(men_men_n362_));
  NO3        u0334(.A(men_men_n316_), .B(men_men_n70_), .C(men_men_n210_), .Y(men_men_n363_));
  NA3        u0335(.A(men_men_n204_), .B(men_men_n202_), .C(men_men_n35_), .Y(men_men_n364_));
  AOI220     u0336(.A0(men_men_n364_), .A1(men_men_n360_), .B0(men_men_n363_), .B1(men_men_n362_), .Y(men_men_n365_));
  NA2        u0337(.A(men_men_n203_), .B(k), .Y(men_men_n366_));
  NA3        u0338(.A(m), .B(men_men_n112_), .C(men_men_n209_), .Y(men_men_n367_));
  NA4        u0339(.A(men_men_n198_), .B(men_men_n87_), .C(g), .D(men_men_n209_), .Y(men_men_n368_));
  NAi41      u0340(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n369_));
  NA2        u0341(.A(men_men_n49_), .B(men_men_n113_), .Y(men_men_n370_));
  NO2        u0342(.A(men_men_n370_), .B(men_men_n369_), .Y(men_men_n371_));
  NA2        u0343(.A(men_men_n371_), .B(b), .Y(men_men_n372_));
  NA4        u0344(.A(men_men_n372_), .B(men_men_n365_), .C(men_men_n359_), .D(men_men_n356_), .Y(men_men_n373_));
  NO4        u0345(.A(men_men_n373_), .B(men_men_n350_), .C(men_men_n333_), .D(men_men_n328_), .Y(men_men_n374_));
  NA4        u0346(.A(men_men_n374_), .B(men_men_n312_), .C(men_men_n262_), .D(men_men_n194_), .Y(men10));
  NA3        u0347(.A(m), .B(k), .C(i), .Y(men_men_n376_));
  NO3        u0348(.A(men_men_n376_), .B(j), .C(men_men_n210_), .Y(men_men_n377_));
  NOi21      u0349(.An(e), .B(f), .Y(men_men_n378_));
  NO4        u0350(.A(men_men_n147_), .B(men_men_n378_), .C(n), .D(men_men_n110_), .Y(men_men_n379_));
  NAi31      u0351(.An(b), .B(f), .C(c), .Y(men_men_n380_));
  INV        u0352(.A(men_men_n380_), .Y(men_men_n381_));
  NOi32      u0353(.An(k), .Bn(h), .C(j), .Y(men_men_n382_));
  NA2        u0354(.A(men_men_n382_), .B(men_men_n215_), .Y(men_men_n383_));
  NA2        u0355(.A(men_men_n155_), .B(men_men_n383_), .Y(men_men_n384_));
  AOI220     u0356(.A0(men_men_n384_), .A1(men_men_n381_), .B0(men_men_n379_), .B1(men_men_n377_), .Y(men_men_n385_));
  AN2        u0357(.A(j), .B(h), .Y(men_men_n386_));
  NO3        u0358(.A(n), .B(m), .C(k), .Y(men_men_n387_));
  NA2        u0359(.A(men_men_n387_), .B(men_men_n386_), .Y(men_men_n388_));
  NO3        u0360(.A(men_men_n388_), .B(men_men_n147_), .C(men_men_n209_), .Y(men_men_n389_));
  OR2        u0361(.A(m), .B(k), .Y(men_men_n390_));
  NO2        u0362(.A(men_men_n170_), .B(men_men_n390_), .Y(men_men_n391_));
  NA4        u0363(.A(n), .B(f), .C(c), .D(men_men_n115_), .Y(men_men_n392_));
  NOi21      u0364(.An(men_men_n391_), .B(men_men_n392_), .Y(men_men_n393_));
  NOi32      u0365(.An(d), .Bn(a), .C(c), .Y(men_men_n394_));
  NA2        u0366(.A(men_men_n394_), .B(men_men_n178_), .Y(men_men_n395_));
  NAi21      u0367(.An(i), .B(g), .Y(men_men_n396_));
  NAi31      u0368(.An(k), .B(m), .C(j), .Y(men_men_n397_));
  NO3        u0369(.A(men_men_n397_), .B(men_men_n396_), .C(n), .Y(men_men_n398_));
  NOi21      u0370(.An(men_men_n398_), .B(men_men_n395_), .Y(men_men_n399_));
  NO3        u0371(.A(men_men_n399_), .B(men_men_n393_), .C(men_men_n389_), .Y(men_men_n400_));
  NO2        u0372(.A(men_men_n392_), .B(men_men_n294_), .Y(men_men_n401_));
  NOi32      u0373(.An(f), .Bn(d), .C(c), .Y(men_men_n402_));
  AOI220     u0374(.A0(men_men_n402_), .A1(men_men_n305_), .B0(men_men_n401_), .B1(men_men_n211_), .Y(men_men_n403_));
  NA3        u0375(.A(men_men_n403_), .B(men_men_n400_), .C(men_men_n385_), .Y(men_men_n404_));
  NO2        u0376(.A(men_men_n57_), .B(men_men_n115_), .Y(men_men_n405_));
  NA2        u0377(.A(men_men_n243_), .B(men_men_n405_), .Y(men_men_n406_));
  INV        u0378(.A(e), .Y(men_men_n407_));
  NA2        u0379(.A(men_men_n44_), .B(e), .Y(men_men_n408_));
  OAI220     u0380(.A0(men_men_n408_), .A1(men_men_n195_), .B0(men_men_n199_), .B1(men_men_n407_), .Y(men_men_n409_));
  AN2        u0381(.A(g), .B(e), .Y(men_men_n410_));
  NA3        u0382(.A(men_men_n410_), .B(men_men_n198_), .C(i), .Y(men_men_n411_));
  OAI210     u0383(.A0(men_men_n89_), .A1(men_men_n407_), .B0(men_men_n411_), .Y(men_men_n412_));
  NO2        u0384(.A(men_men_n101_), .B(men_men_n407_), .Y(men_men_n413_));
  NO3        u0385(.A(men_men_n413_), .B(men_men_n412_), .C(men_men_n409_), .Y(men_men_n414_));
  NOi32      u0386(.An(h), .Bn(e), .C(g), .Y(men_men_n415_));
  NA3        u0387(.A(men_men_n415_), .B(men_men_n287_), .C(m), .Y(men_men_n416_));
  NOi21      u0388(.An(g), .B(h), .Y(men_men_n417_));
  AN3        u0389(.A(m), .B(l), .C(i), .Y(men_men_n418_));
  NA3        u0390(.A(men_men_n418_), .B(men_men_n417_), .C(e), .Y(men_men_n419_));
  AN3        u0391(.A(h), .B(g), .C(e), .Y(men_men_n420_));
  NA2        u0392(.A(men_men_n420_), .B(men_men_n98_), .Y(men_men_n421_));
  AN2        u0393(.A(men_men_n421_), .B(men_men_n419_), .Y(men_men_n422_));
  AOI210     u0394(.A0(men_men_n422_), .A1(men_men_n414_), .B0(men_men_n406_), .Y(men_men_n423_));
  NA3        u0395(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n424_), .B(men_men_n406_), .Y(men_men_n425_));
  NAi31      u0397(.An(b), .B(c), .C(a), .Y(men_men_n426_));
  NO2        u0398(.A(men_men_n426_), .B(n), .Y(men_men_n427_));
  NA2        u0399(.A(men_men_n49_), .B(m), .Y(men_men_n428_));
  NO2        u0400(.A(men_men_n428_), .B(men_men_n144_), .Y(men_men_n429_));
  NA2        u0401(.A(men_men_n429_), .B(men_men_n427_), .Y(men_men_n430_));
  INV        u0402(.A(men_men_n430_), .Y(men_men_n431_));
  NO4        u0403(.A(men_men_n431_), .B(men_men_n425_), .C(men_men_n423_), .D(men_men_n404_), .Y(men_men_n432_));
  NA2        u0404(.A(i), .B(g), .Y(men_men_n433_));
  NO3        u0405(.A(men_men_n271_), .B(men_men_n433_), .C(c), .Y(men_men_n434_));
  NOi21      u0406(.An(a), .B(n), .Y(men_men_n435_));
  NOi21      u0407(.An(d), .B(c), .Y(men_men_n436_));
  NA2        u0408(.A(men_men_n436_), .B(men_men_n435_), .Y(men_men_n437_));
  NA3        u0409(.A(i), .B(g), .C(f), .Y(men_men_n438_));
  OR2        u0410(.A(men_men_n438_), .B(men_men_n69_), .Y(men_men_n439_));
  NA3        u0411(.A(men_men_n418_), .B(men_men_n417_), .C(men_men_n178_), .Y(men_men_n440_));
  AOI210     u0412(.A0(men_men_n440_), .A1(men_men_n439_), .B0(men_men_n437_), .Y(men_men_n441_));
  AOI210     u0413(.A0(men_men_n434_), .A1(men_men_n286_), .B0(men_men_n441_), .Y(men_men_n442_));
  OR2        u0414(.A(n), .B(m), .Y(men_men_n443_));
  NO2        u0415(.A(men_men_n443_), .B(men_men_n148_), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n179_), .B(men_men_n144_), .Y(men_men_n445_));
  OAI210     u0417(.A0(men_men_n444_), .A1(men_men_n172_), .B0(men_men_n445_), .Y(men_men_n446_));
  INV        u0418(.A(men_men_n370_), .Y(men_men_n447_));
  NA3        u0419(.A(men_men_n447_), .B(men_men_n360_), .C(d), .Y(men_men_n448_));
  NO2        u0420(.A(men_men_n426_), .B(men_men_n47_), .Y(men_men_n449_));
  NAi21      u0421(.An(k), .B(j), .Y(men_men_n450_));
  NAi21      u0422(.An(e), .B(d), .Y(men_men_n451_));
  INV        u0423(.A(men_men_n451_), .Y(men_men_n452_));
  NO2        u0424(.A(men_men_n246_), .B(men_men_n209_), .Y(men_men_n453_));
  NA3        u0425(.A(men_men_n453_), .B(men_men_n452_), .C(men_men_n221_), .Y(men_men_n454_));
  NA3        u0426(.A(men_men_n454_), .B(men_men_n448_), .C(men_men_n446_), .Y(men_men_n455_));
  NOi31      u0427(.An(n), .B(m), .C(k), .Y(men_men_n456_));
  AOI220     u0428(.A0(men_men_n456_), .A1(men_men_n386_), .B0(men_men_n215_), .B1(men_men_n48_), .Y(men_men_n457_));
  NAi31      u0429(.An(g), .B(f), .C(c), .Y(men_men_n458_));
  OR3        u0430(.A(men_men_n458_), .B(men_men_n457_), .C(e), .Y(men_men_n459_));
  INV        u0431(.A(men_men_n459_), .Y(men_men_n460_));
  NOi41      u0432(.An(men_men_n442_), .B(men_men_n460_), .C(men_men_n455_), .D(men_men_n260_), .Y(men_men_n461_));
  NOi32      u0433(.An(c), .Bn(a), .C(b), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n462_), .B(men_men_n113_), .Y(men_men_n463_));
  INV        u0435(.A(men_men_n269_), .Y(men_men_n464_));
  AN2        u0436(.A(e), .B(d), .Y(men_men_n465_));
  NA2        u0437(.A(men_men_n465_), .B(men_men_n464_), .Y(men_men_n466_));
  INV        u0438(.A(men_men_n144_), .Y(men_men_n467_));
  NO2        u0439(.A(men_men_n130_), .B(men_men_n41_), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n64_), .B(e), .Y(men_men_n469_));
  NOi31      u0441(.An(j), .B(k), .C(i), .Y(men_men_n470_));
  NOi21      u0442(.An(men_men_n160_), .B(men_men_n470_), .Y(men_men_n471_));
  NA4        u0443(.A(men_men_n319_), .B(men_men_n471_), .C(men_men_n254_), .D(men_men_n118_), .Y(men_men_n472_));
  AOI220     u0444(.A0(men_men_n472_), .A1(men_men_n469_), .B0(men_men_n468_), .B1(men_men_n467_), .Y(men_men_n473_));
  AOI210     u0445(.A0(men_men_n473_), .A1(men_men_n466_), .B0(men_men_n463_), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n205_), .B(men_men_n200_), .Y(men_men_n475_));
  NOi21      u0447(.An(a), .B(b), .Y(men_men_n476_));
  NA3        u0448(.A(e), .B(d), .C(c), .Y(men_men_n477_));
  NAi21      u0449(.An(men_men_n477_), .B(men_men_n476_), .Y(men_men_n478_));
  AOI210     u0450(.A0(men_men_n263_), .A1(men_men_n475_), .B0(men_men_n478_), .Y(men_men_n479_));
  NO4        u0451(.A(men_men_n182_), .B(men_men_n104_), .C(men_men_n54_), .D(b), .Y(men_men_n480_));
  NA2        u0452(.A(men_men_n381_), .B(men_men_n149_), .Y(men_men_n481_));
  OR2        u0453(.A(k), .B(j), .Y(men_men_n482_));
  NA2        u0454(.A(l), .B(k), .Y(men_men_n483_));
  AOI210     u0455(.A0(men_men_n228_), .A1(men_men_n334_), .B0(men_men_n84_), .Y(men_men_n484_));
  NA2        u0456(.A(men_men_n274_), .B(men_men_n127_), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n394_), .B(men_men_n113_), .Y(men_men_n486_));
  NO4        u0458(.A(men_men_n486_), .B(men_men_n95_), .C(men_men_n112_), .D(e), .Y(men_men_n487_));
  NO2        u0459(.A(men_men_n487_), .B(men_men_n485_), .Y(men_men_n488_));
  NA2        u0460(.A(men_men_n488_), .B(men_men_n481_), .Y(men_men_n489_));
  NO4        u0461(.A(men_men_n489_), .B(men_men_n480_), .C(men_men_n479_), .D(men_men_n474_), .Y(men_men_n490_));
  NA2        u0462(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n491_));
  NAi31      u0463(.An(j), .B(l), .C(i), .Y(men_men_n492_));
  OAI210     u0464(.A0(men_men_n492_), .A1(men_men_n131_), .B0(men_men_n104_), .Y(men_men_n493_));
  NO3        u0465(.A(men_men_n395_), .B(men_men_n342_), .C(men_men_n196_), .Y(men_men_n494_));
  NO2        u0466(.A(men_men_n395_), .B(men_men_n370_), .Y(men_men_n495_));
  NO3        u0467(.A(men_men_n495_), .B(men_men_n494_), .C(men_men_n303_), .Y(men_men_n496_));
  NA3        u0468(.A(men_men_n496_), .B(men_men_n491_), .C(men_men_n238_), .Y(men_men_n497_));
  OAI210     u0469(.A0(men_men_n126_), .A1(men_men_n125_), .B0(n), .Y(men_men_n498_));
  NO2        u0470(.A(men_men_n498_), .B(men_men_n130_), .Y(men_men_n499_));
  OR2        u0471(.A(men_men_n295_), .B(men_men_n240_), .Y(men_men_n500_));
  OA210      u0472(.A0(men_men_n500_), .A1(men_men_n499_), .B0(men_men_n187_), .Y(men_men_n501_));
  XO2        u0473(.A(i), .B(h), .Y(men_men_n502_));
  NA3        u0474(.A(men_men_n502_), .B(men_men_n154_), .C(n), .Y(men_men_n503_));
  NAi41      u0475(.An(men_men_n295_), .B(men_men_n503_), .C(men_men_n457_), .D(men_men_n383_), .Y(men_men_n504_));
  NOi32      u0476(.An(men_men_n504_), .Bn(men_men_n469_), .C(men_men_n265_), .Y(men_men_n505_));
  NAi31      u0477(.An(c), .B(f), .C(d), .Y(men_men_n506_));
  AOI210     u0478(.A0(men_men_n275_), .A1(men_men_n190_), .B0(men_men_n506_), .Y(men_men_n507_));
  NOi21      u0479(.An(men_men_n82_), .B(men_men_n507_), .Y(men_men_n508_));
  NA3        u0480(.A(men_men_n379_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n509_));
  NA2        u0481(.A(men_men_n222_), .B(men_men_n109_), .Y(men_men_n510_));
  AOI210     u0482(.A0(men_men_n510_), .A1(men_men_n177_), .B0(men_men_n506_), .Y(men_men_n511_));
  NOi21      u0483(.An(men_men_n509_), .B(men_men_n511_), .Y(men_men_n512_));
  AO220      u0484(.A0(men_men_n283_), .A1(men_men_n257_), .B0(men_men_n161_), .B1(men_men_n65_), .Y(men_men_n513_));
  NA3        u0485(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n514_));
  NO2        u0486(.A(men_men_n514_), .B(men_men_n437_), .Y(men_men_n515_));
  NO2        u0487(.A(men_men_n515_), .B(men_men_n291_), .Y(men_men_n516_));
  NAi41      u0488(.An(men_men_n513_), .B(men_men_n516_), .C(men_men_n512_), .D(men_men_n508_), .Y(men_men_n517_));
  NO4        u0489(.A(men_men_n517_), .B(men_men_n505_), .C(men_men_n501_), .D(men_men_n497_), .Y(men_men_n518_));
  NA4        u0490(.A(men_men_n518_), .B(men_men_n490_), .C(men_men_n461_), .D(men_men_n432_), .Y(men11));
  NO2        u0491(.A(men_men_n71_), .B(f), .Y(men_men_n520_));
  NA2        u0492(.A(j), .B(g), .Y(men_men_n521_));
  NAi31      u0493(.An(i), .B(m), .C(l), .Y(men_men_n522_));
  NA3        u0494(.A(m), .B(k), .C(j), .Y(men_men_n523_));
  OAI220     u0495(.A0(men_men_n523_), .A1(men_men_n130_), .B0(men_men_n522_), .B1(men_men_n521_), .Y(men_men_n524_));
  NA2        u0496(.A(men_men_n524_), .B(men_men_n520_), .Y(men_men_n525_));
  NOi32      u0497(.An(e), .Bn(b), .C(f), .Y(men_men_n526_));
  NA2        u0498(.A(men_men_n253_), .B(men_men_n113_), .Y(men_men_n527_));
  NA2        u0499(.A(men_men_n44_), .B(j), .Y(men_men_n528_));
  NO2        u0500(.A(men_men_n528_), .B(men_men_n297_), .Y(men_men_n529_));
  NAi31      u0501(.An(d), .B(e), .C(a), .Y(men_men_n530_));
  NO2        u0502(.A(men_men_n530_), .B(n), .Y(men_men_n531_));
  AOI220     u0503(.A0(men_men_n531_), .A1(men_men_n102_), .B0(men_men_n529_), .B1(men_men_n526_), .Y(men_men_n532_));
  NAi41      u0504(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n533_));
  AN2        u0505(.A(men_men_n533_), .B(men_men_n369_), .Y(men_men_n534_));
  AOI210     u0506(.A0(men_men_n534_), .A1(men_men_n395_), .B0(men_men_n266_), .Y(men_men_n535_));
  NA2        u0507(.A(j), .B(i), .Y(men_men_n536_));
  NAi31      u0508(.An(n), .B(m), .C(k), .Y(men_men_n537_));
  NO3        u0509(.A(men_men_n537_), .B(men_men_n536_), .C(men_men_n112_), .Y(men_men_n538_));
  NO4        u0510(.A(n), .B(d), .C(men_men_n115_), .D(a), .Y(men_men_n539_));
  OR2        u0511(.A(n), .B(c), .Y(men_men_n540_));
  NO2        u0512(.A(men_men_n540_), .B(men_men_n145_), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(men_men_n539_), .Y(men_men_n542_));
  NOi32      u0514(.An(g), .Bn(f), .C(i), .Y(men_men_n543_));
  AOI220     u0515(.A0(men_men_n543_), .A1(men_men_n100_), .B0(men_men_n524_), .B1(f), .Y(men_men_n544_));
  NO2        u0516(.A(men_men_n269_), .B(men_men_n47_), .Y(men_men_n545_));
  NO2        u0517(.A(men_men_n544_), .B(men_men_n542_), .Y(men_men_n546_));
  INV        u0518(.A(men_men_n546_), .Y(men_men_n547_));
  NA2        u0519(.A(men_men_n137_), .B(men_men_n34_), .Y(men_men_n548_));
  OAI220     u0520(.A0(men_men_n548_), .A1(m), .B0(men_men_n528_), .B1(men_men_n228_), .Y(men_men_n549_));
  NOi41      u0521(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n550_));
  NAi32      u0522(.An(e), .Bn(b), .C(c), .Y(men_men_n551_));
  OR2        u0523(.A(men_men_n551_), .B(men_men_n84_), .Y(men_men_n552_));
  AN2        u0524(.A(men_men_n335_), .B(men_men_n316_), .Y(men_men_n553_));
  NA2        u0525(.A(men_men_n553_), .B(men_men_n552_), .Y(men_men_n554_));
  OA210      u0526(.A0(men_men_n554_), .A1(men_men_n550_), .B0(men_men_n549_), .Y(men_men_n555_));
  OAI220     u0527(.A0(men_men_n397_), .A1(men_men_n396_), .B0(men_men_n522_), .B1(men_men_n521_), .Y(men_men_n556_));
  NAi31      u0528(.An(d), .B(c), .C(a), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n557_), .B(n), .Y(men_men_n558_));
  NA3        u0530(.A(men_men_n558_), .B(men_men_n556_), .C(e), .Y(men_men_n559_));
  NO3        u0531(.A(men_men_n60_), .B(men_men_n47_), .C(men_men_n210_), .Y(men_men_n560_));
  NO2        u0532(.A(men_men_n225_), .B(men_men_n110_), .Y(men_men_n561_));
  OAI210     u0533(.A0(men_men_n560_), .A1(men_men_n398_), .B0(men_men_n561_), .Y(men_men_n562_));
  NA2        u0534(.A(men_men_n562_), .B(men_men_n559_), .Y(men_men_n563_));
  NO2        u0535(.A(men_men_n271_), .B(n), .Y(men_men_n564_));
  NO2        u0536(.A(men_men_n427_), .B(men_men_n564_), .Y(men_men_n565_));
  NA2        u0537(.A(men_men_n556_), .B(f), .Y(men_men_n566_));
  NAi32      u0538(.An(d), .Bn(a), .C(b), .Y(men_men_n567_));
  NA2        u0539(.A(h), .B(f), .Y(men_men_n568_));
  NO2        u0540(.A(men_men_n568_), .B(men_men_n95_), .Y(men_men_n569_));
  NO3        u0541(.A(men_men_n173_), .B(men_men_n170_), .C(g), .Y(men_men_n570_));
  NA2        u0542(.A(men_men_n570_), .B(men_men_n56_), .Y(men_men_n571_));
  OAI210     u0543(.A0(men_men_n566_), .A1(men_men_n565_), .B0(men_men_n571_), .Y(men_men_n572_));
  AN3        u0544(.A(j), .B(h), .C(g), .Y(men_men_n573_));
  NO2        u0545(.A(men_men_n143_), .B(c), .Y(men_men_n574_));
  NA3        u0546(.A(men_men_n574_), .B(men_men_n573_), .C(men_men_n456_), .Y(men_men_n575_));
  NA3        u0547(.A(f), .B(d), .C(b), .Y(men_men_n576_));
  NO4        u0548(.A(men_men_n576_), .B(men_men_n173_), .C(men_men_n170_), .D(g), .Y(men_men_n577_));
  NAi21      u0549(.An(men_men_n577_), .B(men_men_n575_), .Y(men_men_n578_));
  NO4        u0550(.A(men_men_n578_), .B(men_men_n572_), .C(men_men_n563_), .D(men_men_n555_), .Y(men_men_n579_));
  AN4        u0551(.A(men_men_n579_), .B(men_men_n547_), .C(men_men_n532_), .D(men_men_n525_), .Y(men_men_n580_));
  INV        u0552(.A(k), .Y(men_men_n581_));
  NA3        u0553(.A(l), .B(men_men_n581_), .C(i), .Y(men_men_n582_));
  INV        u0554(.A(men_men_n582_), .Y(men_men_n583_));
  NA4        u0555(.A(men_men_n394_), .B(men_men_n417_), .C(men_men_n178_), .D(men_men_n113_), .Y(men_men_n584_));
  NAi32      u0556(.An(h), .Bn(f), .C(g), .Y(men_men_n585_));
  NAi41      u0557(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n586_));
  OAI210     u0558(.A0(men_men_n530_), .A1(n), .B0(men_men_n586_), .Y(men_men_n587_));
  NA2        u0559(.A(men_men_n587_), .B(m), .Y(men_men_n588_));
  NAi31      u0560(.An(h), .B(g), .C(f), .Y(men_men_n589_));
  OR3        u0561(.A(men_men_n589_), .B(men_men_n271_), .C(men_men_n47_), .Y(men_men_n590_));
  NA4        u0562(.A(men_men_n417_), .B(men_men_n120_), .C(men_men_n113_), .D(e), .Y(men_men_n591_));
  AN2        u0563(.A(men_men_n591_), .B(men_men_n590_), .Y(men_men_n592_));
  OA210      u0564(.A0(men_men_n588_), .A1(men_men_n585_), .B0(men_men_n592_), .Y(men_men_n593_));
  NO3        u0565(.A(men_men_n585_), .B(men_men_n71_), .C(men_men_n73_), .Y(men_men_n594_));
  NO4        u0566(.A(men_men_n589_), .B(men_men_n540_), .C(men_men_n145_), .D(men_men_n73_), .Y(men_men_n595_));
  OR2        u0567(.A(men_men_n595_), .B(men_men_n594_), .Y(men_men_n596_));
  NAi31      u0568(.An(men_men_n596_), .B(men_men_n593_), .C(men_men_n584_), .Y(men_men_n597_));
  NAi31      u0569(.An(f), .B(h), .C(g), .Y(men_men_n598_));
  NO4        u0570(.A(men_men_n307_), .B(men_men_n598_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n599_));
  NOi32      u0571(.An(b), .Bn(a), .C(c), .Y(men_men_n600_));
  NOi41      u0572(.An(men_men_n600_), .B(men_men_n351_), .C(men_men_n67_), .D(men_men_n116_), .Y(men_men_n601_));
  OR2        u0573(.A(men_men_n601_), .B(men_men_n599_), .Y(men_men_n602_));
  NOi32      u0574(.An(d), .Bn(a), .C(e), .Y(men_men_n603_));
  NA2        u0575(.A(men_men_n603_), .B(men_men_n113_), .Y(men_men_n604_));
  NO2        u0576(.A(n), .B(c), .Y(men_men_n605_));
  NA3        u0577(.A(men_men_n605_), .B(men_men_n29_), .C(m), .Y(men_men_n606_));
  NA2        u0578(.A(men_men_n606_), .B(men_men_n604_), .Y(men_men_n607_));
  NOi32      u0579(.An(e), .Bn(a), .C(d), .Y(men_men_n608_));
  AOI210     u0580(.A0(men_men_n29_), .A1(d), .B0(men_men_n608_), .Y(men_men_n609_));
  AOI210     u0581(.A0(men_men_n609_), .A1(men_men_n209_), .B0(men_men_n548_), .Y(men_men_n610_));
  AOI210     u0582(.A0(men_men_n610_), .A1(men_men_n607_), .B0(men_men_n602_), .Y(men_men_n611_));
  INV        u0583(.A(men_men_n611_), .Y(men_men_n612_));
  AOI210     u0584(.A0(men_men_n597_), .A1(men_men_n583_), .B0(men_men_n612_), .Y(men_men_n613_));
  NO3        u0585(.A(men_men_n314_), .B(men_men_n59_), .C(n), .Y(men_men_n614_));
  NA3        u0586(.A(men_men_n506_), .B(men_men_n168_), .C(men_men_n167_), .Y(men_men_n615_));
  NA2        u0587(.A(men_men_n458_), .B(men_men_n225_), .Y(men_men_n616_));
  OR2        u0588(.A(men_men_n616_), .B(men_men_n615_), .Y(men_men_n617_));
  NA2        u0589(.A(men_men_n74_), .B(men_men_n113_), .Y(men_men_n618_));
  NO2        u0590(.A(men_men_n618_), .B(men_men_n43_), .Y(men_men_n619_));
  AOI220     u0591(.A0(men_men_n619_), .A1(men_men_n535_), .B0(men_men_n617_), .B1(men_men_n614_), .Y(men_men_n620_));
  NO2        u0592(.A(men_men_n620_), .B(men_men_n87_), .Y(men_men_n621_));
  NA3        u0593(.A(men_men_n550_), .B(men_men_n337_), .C(men_men_n44_), .Y(men_men_n622_));
  NOi32      u0594(.An(e), .Bn(c), .C(f), .Y(men_men_n623_));
  NOi21      u0595(.An(f), .B(g), .Y(men_men_n624_));
  NO2        u0596(.A(men_men_n624_), .B(men_men_n207_), .Y(men_men_n625_));
  AOI220     u0597(.A0(men_men_n625_), .A1(men_men_n391_), .B0(men_men_n623_), .B1(men_men_n172_), .Y(men_men_n626_));
  NA3        u0598(.A(men_men_n626_), .B(men_men_n622_), .C(men_men_n175_), .Y(men_men_n627_));
  AOI210     u0599(.A0(men_men_n534_), .A1(men_men_n395_), .B0(men_men_n296_), .Y(men_men_n628_));
  NA2        u0600(.A(men_men_n628_), .B(men_men_n258_), .Y(men_men_n629_));
  NOi21      u0601(.An(j), .B(l), .Y(men_men_n630_));
  NAi21      u0602(.An(k), .B(h), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n631_), .B(men_men_n256_), .Y(men_men_n632_));
  NA2        u0604(.A(men_men_n632_), .B(men_men_n630_), .Y(men_men_n633_));
  OR2        u0605(.A(men_men_n633_), .B(men_men_n588_), .Y(men_men_n634_));
  NOi31      u0606(.An(m), .B(n), .C(k), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n630_), .B(men_men_n635_), .Y(men_men_n636_));
  NO2        u0608(.A(men_men_n271_), .B(men_men_n47_), .Y(men_men_n637_));
  NO2        u0609(.A(men_men_n307_), .B(men_men_n598_), .Y(men_men_n638_));
  NO2        u0610(.A(men_men_n530_), .B(men_men_n47_), .Y(men_men_n639_));
  AOI220     u0611(.A0(men_men_n639_), .A1(men_men_n638_), .B0(men_men_n637_), .B1(men_men_n569_), .Y(men_men_n640_));
  NA3        u0612(.A(men_men_n640_), .B(men_men_n634_), .C(men_men_n629_), .Y(men_men_n641_));
  NA2        u0613(.A(men_men_n109_), .B(men_men_n36_), .Y(men_men_n642_));
  INV        u0614(.A(men_men_n360_), .Y(men_men_n643_));
  NO2        u0615(.A(men_men_n643_), .B(n), .Y(men_men_n644_));
  NO2        u0616(.A(men_men_n528_), .B(men_men_n173_), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n551_), .B(men_men_n265_), .C(men_men_n141_), .Y(men_men_n646_));
  NA2        u0618(.A(men_men_n502_), .B(men_men_n154_), .Y(men_men_n647_));
  NO3        u0619(.A(men_men_n392_), .B(men_men_n647_), .C(men_men_n87_), .Y(men_men_n648_));
  AOI210     u0620(.A0(men_men_n646_), .A1(men_men_n645_), .B0(men_men_n648_), .Y(men_men_n649_));
  AN3        u0621(.A(f), .B(d), .C(b), .Y(men_men_n650_));
  OAI210     u0622(.A0(men_men_n650_), .A1(men_men_n129_), .B0(n), .Y(men_men_n651_));
  NA3        u0623(.A(men_men_n502_), .B(men_men_n154_), .C(men_men_n210_), .Y(men_men_n652_));
  AOI210     u0624(.A0(men_men_n651_), .A1(men_men_n227_), .B0(men_men_n652_), .Y(men_men_n653_));
  NAi31      u0625(.An(m), .B(n), .C(k), .Y(men_men_n654_));
  OR2        u0626(.A(men_men_n133_), .B(men_men_n59_), .Y(men_men_n655_));
  OAI210     u0627(.A0(men_men_n655_), .A1(men_men_n654_), .B0(men_men_n244_), .Y(men_men_n656_));
  OAI210     u0628(.A0(men_men_n656_), .A1(men_men_n653_), .B0(j), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n657_), .B(men_men_n649_), .Y(men_men_n658_));
  NO4        u0630(.A(men_men_n658_), .B(men_men_n641_), .C(men_men_n627_), .D(men_men_n621_), .Y(men_men_n659_));
  NA2        u0631(.A(men_men_n379_), .B(men_men_n157_), .Y(men_men_n660_));
  NAi31      u0632(.An(g), .B(h), .C(f), .Y(men_men_n661_));
  OR3        u0633(.A(men_men_n661_), .B(men_men_n271_), .C(n), .Y(men_men_n662_));
  OA210      u0634(.A0(men_men_n530_), .A1(n), .B0(men_men_n586_), .Y(men_men_n663_));
  NA3        u0635(.A(men_men_n415_), .B(men_men_n120_), .C(men_men_n84_), .Y(men_men_n664_));
  OAI210     u0636(.A0(men_men_n663_), .A1(men_men_n91_), .B0(men_men_n664_), .Y(men_men_n665_));
  NOi21      u0637(.An(men_men_n662_), .B(men_men_n665_), .Y(men_men_n666_));
  AOI210     u0638(.A0(men_men_n666_), .A1(men_men_n660_), .B0(men_men_n523_), .Y(men_men_n667_));
  NO3        u0639(.A(g), .B(men_men_n209_), .C(men_men_n54_), .Y(men_men_n668_));
  NO2        u0640(.A(men_men_n510_), .B(men_men_n87_), .Y(men_men_n669_));
  OAI210     u0641(.A0(men_men_n669_), .A1(men_men_n391_), .B0(men_men_n668_), .Y(men_men_n670_));
  OR2        u0642(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n671_));
  NA2        u0643(.A(men_men_n600_), .B(men_men_n339_), .Y(men_men_n672_));
  OA220      u0644(.A0(men_men_n636_), .A1(men_men_n672_), .B0(men_men_n633_), .B1(men_men_n671_), .Y(men_men_n673_));
  AN2        u0645(.A(h), .B(f), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n674_), .B(men_men_n37_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n100_), .B(men_men_n44_), .Y(men_men_n676_));
  OAI220     u0648(.A0(men_men_n676_), .A1(men_men_n330_), .B0(men_men_n675_), .B1(men_men_n463_), .Y(men_men_n677_));
  AOI210     u0649(.A0(men_men_n567_), .A1(men_men_n426_), .B0(men_men_n47_), .Y(men_men_n678_));
  OAI220     u0650(.A0(men_men_n589_), .A1(men_men_n582_), .B0(men_men_n323_), .B1(men_men_n521_), .Y(men_men_n679_));
  AOI210     u0651(.A0(men_men_n679_), .A1(men_men_n678_), .B0(men_men_n677_), .Y(men_men_n680_));
  NA3        u0652(.A(men_men_n680_), .B(men_men_n673_), .C(men_men_n670_), .Y(men_men_n681_));
  NO2        u0653(.A(men_men_n245_), .B(f), .Y(men_men_n682_));
  NO2        u0654(.A(men_men_n624_), .B(men_men_n59_), .Y(men_men_n683_));
  NO3        u0655(.A(men_men_n683_), .B(men_men_n682_), .C(men_men_n34_), .Y(men_men_n684_));
  NA2        u0656(.A(men_men_n326_), .B(men_men_n137_), .Y(men_men_n685_));
  NA2        u0657(.A(men_men_n131_), .B(men_men_n47_), .Y(men_men_n686_));
  AOI220     u0658(.A0(men_men_n686_), .A1(men_men_n526_), .B0(men_men_n360_), .B1(men_men_n113_), .Y(men_men_n687_));
  OA220      u0659(.A0(men_men_n687_), .A1(men_men_n548_), .B0(men_men_n358_), .B1(men_men_n111_), .Y(men_men_n688_));
  OAI210     u0660(.A0(men_men_n685_), .A1(men_men_n684_), .B0(men_men_n688_), .Y(men_men_n689_));
  NO3        u0661(.A(men_men_n402_), .B(men_men_n187_), .C(men_men_n186_), .Y(men_men_n690_));
  NA2        u0662(.A(men_men_n690_), .B(men_men_n225_), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n691_), .B(men_men_n247_), .C(j), .Y(men_men_n692_));
  NA2        u0664(.A(men_men_n462_), .B(men_men_n84_), .Y(men_men_n693_));
  NO4        u0665(.A(men_men_n523_), .B(men_men_n693_), .C(men_men_n130_), .D(men_men_n209_), .Y(men_men_n694_));
  INV        u0666(.A(men_men_n694_), .Y(men_men_n695_));
  NA4        u0667(.A(men_men_n695_), .B(men_men_n692_), .C(men_men_n509_), .D(men_men_n400_), .Y(men_men_n696_));
  NO4        u0668(.A(men_men_n696_), .B(men_men_n689_), .C(men_men_n681_), .D(men_men_n667_), .Y(men_men_n697_));
  NA4        u0669(.A(men_men_n697_), .B(men_men_n659_), .C(men_men_n613_), .D(men_men_n580_), .Y(men08));
  NO2        u0670(.A(k), .B(h), .Y(men_men_n699_));
  AO210      u0671(.A0(men_men_n245_), .A1(men_men_n450_), .B0(men_men_n699_), .Y(men_men_n700_));
  NO2        u0672(.A(men_men_n700_), .B(men_men_n294_), .Y(men_men_n701_));
  NA2        u0673(.A(men_men_n623_), .B(men_men_n84_), .Y(men_men_n702_));
  NA2        u0674(.A(men_men_n702_), .B(men_men_n458_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n703_), .B(men_men_n701_), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n84_), .B(men_men_n110_), .Y(men_men_n705_));
  NO2        u0677(.A(men_men_n705_), .B(men_men_n55_), .Y(men_men_n706_));
  NO4        u0678(.A(men_men_n376_), .B(men_men_n112_), .C(j), .D(men_men_n210_), .Y(men_men_n707_));
  NA2        u0679(.A(men_men_n576_), .B(men_men_n227_), .Y(men_men_n708_));
  AOI220     u0680(.A0(men_men_n708_), .A1(men_men_n345_), .B0(men_men_n707_), .B1(men_men_n706_), .Y(men_men_n709_));
  AOI210     u0681(.A0(men_men_n576_), .A1(men_men_n151_), .B0(men_men_n84_), .Y(men_men_n710_));
  NA4        u0682(.A(men_men_n212_), .B(men_men_n137_), .C(men_men_n43_), .D(h), .Y(men_men_n711_));
  AN2        u0683(.A(l), .B(k), .Y(men_men_n712_));
  NA4        u0684(.A(men_men_n712_), .B(men_men_n109_), .C(men_men_n73_), .D(men_men_n210_), .Y(men_men_n713_));
  OAI210     u0685(.A0(men_men_n711_), .A1(g), .B0(men_men_n713_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n714_), .B(men_men_n710_), .Y(men_men_n715_));
  NA4        u0687(.A(men_men_n715_), .B(men_men_n709_), .C(men_men_n704_), .D(men_men_n347_), .Y(men_men_n716_));
  AN2        u0688(.A(men_men_n531_), .B(men_men_n96_), .Y(men_men_n717_));
  NO4        u0689(.A(men_men_n170_), .B(men_men_n390_), .C(men_men_n112_), .D(g), .Y(men_men_n718_));
  AOI210     u0690(.A0(men_men_n718_), .A1(men_men_n708_), .B0(men_men_n515_), .Y(men_men_n719_));
  NO2        u0691(.A(men_men_n38_), .B(men_men_n209_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n720_), .B(men_men_n564_), .Y(men_men_n721_));
  NAi31      u0693(.An(men_men_n717_), .B(men_men_n721_), .C(men_men_n719_), .Y(men_men_n722_));
  OAI210     u0694(.A0(men_men_n551_), .A1(men_men_n45_), .B0(men_men_n655_), .Y(men_men_n723_));
  NO2        u0695(.A(men_men_n483_), .B(men_men_n131_), .Y(men_men_n724_));
  NA2        u0696(.A(men_men_n724_), .B(men_men_n723_), .Y(men_men_n725_));
  INV        u0697(.A(men_men_n713_), .Y(men_men_n726_));
  NA2        u0698(.A(men_men_n700_), .B(men_men_n134_), .Y(men_men_n727_));
  AOI220     u0699(.A0(men_men_n727_), .A1(men_men_n401_), .B0(men_men_n726_), .B1(men_men_n76_), .Y(men_men_n728_));
  NA2        u0700(.A(men_men_n725_), .B(men_men_n728_), .Y(men_men_n729_));
  NA3        u0701(.A(men_men_n691_), .B(men_men_n332_), .C(men_men_n382_), .Y(men_men_n730_));
  NA2        u0702(.A(men_men_n712_), .B(men_men_n215_), .Y(men_men_n731_));
  NO2        u0703(.A(men_men_n731_), .B(men_men_n325_), .Y(men_men_n732_));
  AOI210     u0704(.A0(men_men_n732_), .A1(men_men_n682_), .B0(men_men_n487_), .Y(men_men_n733_));
  NA3        u0705(.A(m), .B(l), .C(k), .Y(men_men_n734_));
  AOI210     u0706(.A0(men_men_n664_), .A1(men_men_n662_), .B0(men_men_n734_), .Y(men_men_n735_));
  NO2        u0707(.A(men_men_n533_), .B(men_men_n266_), .Y(men_men_n736_));
  NOi21      u0708(.An(men_men_n736_), .B(men_men_n527_), .Y(men_men_n737_));
  NA4        u0709(.A(men_men_n113_), .B(l), .C(k), .D(men_men_n87_), .Y(men_men_n738_));
  NA3        u0710(.A(men_men_n120_), .B(men_men_n410_), .C(i), .Y(men_men_n739_));
  NO2        u0711(.A(men_men_n739_), .B(men_men_n738_), .Y(men_men_n740_));
  NO3        u0712(.A(men_men_n740_), .B(men_men_n737_), .C(men_men_n735_), .Y(men_men_n741_));
  NA3        u0713(.A(men_men_n741_), .B(men_men_n733_), .C(men_men_n730_), .Y(men_men_n742_));
  NO4        u0714(.A(men_men_n742_), .B(men_men_n729_), .C(men_men_n722_), .D(men_men_n716_), .Y(men_men_n743_));
  NA2        u0715(.A(men_men_n625_), .B(men_men_n391_), .Y(men_men_n744_));
  NOi31      u0716(.An(g), .B(h), .C(f), .Y(men_men_n745_));
  NA2        u0717(.A(men_men_n639_), .B(men_men_n745_), .Y(men_men_n746_));
  AO210      u0718(.A0(men_men_n746_), .A1(men_men_n590_), .B0(men_men_n536_), .Y(men_men_n747_));
  INV        u0719(.A(men_men_n495_), .Y(men_men_n748_));
  NA4        u0720(.A(men_men_n748_), .B(men_men_n747_), .C(men_men_n744_), .D(men_men_n244_), .Y(men_men_n749_));
  NA2        u0721(.A(men_men_n712_), .B(men_men_n73_), .Y(men_men_n750_));
  NO4        u0722(.A(men_men_n690_), .B(men_men_n170_), .C(n), .D(i), .Y(men_men_n751_));
  NOi21      u0723(.An(h), .B(j), .Y(men_men_n752_));
  NA2        u0724(.A(men_men_n752_), .B(f), .Y(men_men_n753_));
  INV        u0725(.A(men_men_n751_), .Y(men_men_n754_));
  OAI220     u0726(.A0(men_men_n754_), .A1(men_men_n750_), .B0(men_men_n592_), .B1(men_men_n60_), .Y(men_men_n755_));
  AOI210     u0727(.A0(men_men_n749_), .A1(l), .B0(men_men_n755_), .Y(men_men_n756_));
  NO2        u0728(.A(j), .B(i), .Y(men_men_n757_));
  NA2        u0729(.A(men_men_n757_), .B(men_men_n33_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n420_), .B(men_men_n120_), .Y(men_men_n759_));
  OR2        u0731(.A(men_men_n759_), .B(men_men_n758_), .Y(men_men_n760_));
  NO3        u0732(.A(men_men_n147_), .B(men_men_n47_), .C(men_men_n110_), .Y(men_men_n761_));
  NO3        u0733(.A(men_men_n540_), .B(men_men_n145_), .C(men_men_n73_), .Y(men_men_n762_));
  NO3        u0734(.A(men_men_n483_), .B(men_men_n438_), .C(j), .Y(men_men_n763_));
  OAI210     u0735(.A0(men_men_n762_), .A1(men_men_n761_), .B0(men_men_n763_), .Y(men_men_n764_));
  OAI210     u0736(.A0(men_men_n746_), .A1(men_men_n60_), .B0(men_men_n764_), .Y(men_men_n765_));
  NA2        u0737(.A(k), .B(j), .Y(men_men_n766_));
  NO3        u0738(.A(men_men_n294_), .B(men_men_n766_), .C(men_men_n40_), .Y(men_men_n767_));
  AOI210     u0739(.A0(men_men_n526_), .A1(n), .B0(men_men_n550_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n768_), .B(men_men_n553_), .Y(men_men_n769_));
  AN3        u0741(.A(men_men_n769_), .B(men_men_n767_), .C(men_men_n99_), .Y(men_men_n770_));
  NA2        u0742(.A(men_men_n616_), .B(men_men_n305_), .Y(men_men_n771_));
  NAi31      u0743(.An(men_men_n609_), .B(men_men_n93_), .C(men_men_n84_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n772_), .B(men_men_n771_), .Y(men_men_n773_));
  NO2        u0745(.A(men_men_n294_), .B(men_men_n134_), .Y(men_men_n774_));
  NA2        u0746(.A(men_men_n774_), .B(men_men_n625_), .Y(men_men_n775_));
  NA2        u0747(.A(men_men_n763_), .B(men_men_n678_), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n776_), .B(men_men_n775_), .Y(men_men_n777_));
  OR4        u0749(.A(men_men_n777_), .B(men_men_n773_), .C(men_men_n770_), .D(men_men_n765_), .Y(men_men_n778_));
  NA3        u0750(.A(men_men_n768_), .B(men_men_n553_), .C(men_men_n552_), .Y(men_men_n779_));
  NA4        u0751(.A(men_men_n779_), .B(men_men_n212_), .C(men_men_n450_), .D(men_men_n34_), .Y(men_men_n780_));
  OAI220     u0752(.A0(men_men_n711_), .A1(men_men_n702_), .B0(men_men_n330_), .B1(men_men_n38_), .Y(men_men_n781_));
  INV        u0753(.A(men_men_n781_), .Y(men_men_n782_));
  NA3        u0754(.A(men_men_n543_), .B(men_men_n287_), .C(h), .Y(men_men_n783_));
  NOi21      u0755(.An(men_men_n678_), .B(men_men_n783_), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n92_), .B(men_men_n45_), .Y(men_men_n785_));
  NO2        u0757(.A(men_men_n783_), .B(men_men_n606_), .Y(men_men_n786_));
  AOI210     u0758(.A0(men_men_n785_), .A1(men_men_n644_), .B0(men_men_n786_), .Y(men_men_n787_));
  NAi41      u0759(.An(men_men_n784_), .B(men_men_n787_), .C(men_men_n782_), .D(men_men_n780_), .Y(men_men_n788_));
  AOI220     u0760(.A0(men_men_n96_), .A1(men_men_n233_), .B0(men_men_n763_), .B1(men_men_n637_), .Y(men_men_n789_));
  OAI210     u0761(.A0(men_men_n734_), .A1(men_men_n661_), .B0(men_men_n514_), .Y(men_men_n790_));
  NA3        u0762(.A(men_men_n243_), .B(men_men_n57_), .C(b), .Y(men_men_n791_));
  AOI220     u0763(.A0(men_men_n605_), .A1(men_men_n29_), .B0(men_men_n462_), .B1(men_men_n84_), .Y(men_men_n792_));
  NA2        u0764(.A(men_men_n792_), .B(men_men_n791_), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n783_), .B(men_men_n486_), .Y(men_men_n794_));
  AOI210     u0766(.A0(men_men_n793_), .A1(men_men_n790_), .B0(men_men_n794_), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n795_), .B(men_men_n789_), .Y(men_men_n796_));
  NOi41      u0768(.An(men_men_n760_), .B(men_men_n796_), .C(men_men_n788_), .D(men_men_n778_), .Y(men_men_n797_));
  OR3        u0769(.A(men_men_n711_), .B(men_men_n227_), .C(g), .Y(men_men_n798_));
  NO3        u0770(.A(men_men_n338_), .B(men_men_n296_), .C(men_men_n112_), .Y(men_men_n799_));
  NA2        u0771(.A(men_men_n799_), .B(men_men_n769_), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n44_), .B(men_men_n54_), .Y(men_men_n801_));
  NO3        u0773(.A(men_men_n801_), .B(men_men_n758_), .C(men_men_n271_), .Y(men_men_n802_));
  NO3        u0774(.A(men_men_n521_), .B(men_men_n94_), .C(h), .Y(men_men_n803_));
  AOI210     u0775(.A0(men_men_n803_), .A1(men_men_n706_), .B0(men_men_n802_), .Y(men_men_n804_));
  NA4        u0776(.A(men_men_n804_), .B(men_men_n800_), .C(men_men_n798_), .D(men_men_n403_), .Y(men_men_n805_));
  OR2        u0777(.A(men_men_n661_), .B(men_men_n92_), .Y(men_men_n806_));
  NOi31      u0778(.An(b), .B(d), .C(a), .Y(men_men_n807_));
  NO2        u0779(.A(men_men_n807_), .B(men_men_n603_), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n808_), .B(n), .Y(men_men_n809_));
  NOi21      u0781(.An(men_men_n792_), .B(men_men_n809_), .Y(men_men_n810_));
  OAI220     u0782(.A0(men_men_n810_), .A1(men_men_n806_), .B0(men_men_n783_), .B1(men_men_n604_), .Y(men_men_n811_));
  NO2        u0783(.A(men_men_n551_), .B(men_men_n84_), .Y(men_men_n812_));
  NO3        u0784(.A(men_men_n624_), .B(men_men_n325_), .C(men_men_n116_), .Y(men_men_n813_));
  NOi21      u0785(.An(men_men_n813_), .B(men_men_n155_), .Y(men_men_n814_));
  AOI210     u0786(.A0(men_men_n799_), .A1(men_men_n812_), .B0(men_men_n814_), .Y(men_men_n815_));
  OAI210     u0787(.A0(men_men_n711_), .A1(men_men_n392_), .B0(men_men_n815_), .Y(men_men_n816_));
  NO2        u0788(.A(men_men_n690_), .B(n), .Y(men_men_n817_));
  AOI220     u0789(.A0(men_men_n774_), .A1(men_men_n668_), .B0(men_men_n817_), .B1(men_men_n701_), .Y(men_men_n818_));
  NA2        u0790(.A(men_men_n120_), .B(men_men_n84_), .Y(men_men_n819_));
  AOI210     u0791(.A0(men_men_n424_), .A1(men_men_n416_), .B0(men_men_n819_), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n732_), .B(men_men_n34_), .Y(men_men_n821_));
  NAi21      u0793(.An(men_men_n738_), .B(men_men_n434_), .Y(men_men_n822_));
  NO2        u0794(.A(men_men_n266_), .B(i), .Y(men_men_n823_));
  NA2        u0795(.A(men_men_n718_), .B(men_men_n346_), .Y(men_men_n824_));
  OAI210     u0796(.A0(men_men_n595_), .A1(men_men_n594_), .B0(men_men_n361_), .Y(men_men_n825_));
  AN3        u0797(.A(men_men_n825_), .B(men_men_n824_), .C(men_men_n822_), .Y(men_men_n826_));
  NAi41      u0798(.An(men_men_n820_), .B(men_men_n826_), .C(men_men_n821_), .D(men_men_n818_), .Y(men_men_n827_));
  NO4        u0799(.A(men_men_n827_), .B(men_men_n816_), .C(men_men_n811_), .D(men_men_n805_), .Y(men_men_n828_));
  NA4        u0800(.A(men_men_n828_), .B(men_men_n797_), .C(men_men_n756_), .D(men_men_n743_), .Y(men09));
  INV        u0801(.A(men_men_n121_), .Y(men_men_n830_));
  NA2        u0802(.A(f), .B(e), .Y(men_men_n831_));
  NO2        u0803(.A(men_men_n220_), .B(men_men_n112_), .Y(men_men_n832_));
  NA2        u0804(.A(men_men_n832_), .B(g), .Y(men_men_n833_));
  NA4        u0805(.A(men_men_n307_), .B(men_men_n471_), .C(men_men_n254_), .D(men_men_n118_), .Y(men_men_n834_));
  AOI210     u0806(.A0(men_men_n834_), .A1(g), .B0(men_men_n468_), .Y(men_men_n835_));
  AOI210     u0807(.A0(men_men_n835_), .A1(men_men_n833_), .B0(men_men_n831_), .Y(men_men_n836_));
  NA2        u0808(.A(men_men_n836_), .B(men_men_n830_), .Y(men_men_n837_));
  NA3        u0809(.A(m), .B(l), .C(i), .Y(men_men_n838_));
  OAI220     u0810(.A0(men_men_n589_), .A1(men_men_n838_), .B0(men_men_n351_), .B1(men_men_n522_), .Y(men_men_n839_));
  NA4        u0811(.A(men_men_n88_), .B(men_men_n87_), .C(g), .D(f), .Y(men_men_n840_));
  NAi31      u0812(.An(men_men_n839_), .B(men_men_n840_), .C(men_men_n439_), .Y(men_men_n841_));
  NA3        u0813(.A(men_men_n806_), .B(men_men_n566_), .C(men_men_n514_), .Y(men_men_n842_));
  OA210      u0814(.A0(men_men_n842_), .A1(men_men_n841_), .B0(men_men_n809_), .Y(men_men_n843_));
  INV        u0815(.A(men_men_n335_), .Y(men_men_n844_));
  NO2        u0816(.A(men_men_n126_), .B(men_men_n125_), .Y(men_men_n845_));
  NOi31      u0817(.An(k), .B(m), .C(l), .Y(men_men_n846_));
  NO2        u0818(.A(men_men_n337_), .B(men_men_n846_), .Y(men_men_n847_));
  AOI210     u0819(.A0(men_men_n847_), .A1(men_men_n845_), .B0(men_men_n598_), .Y(men_men_n848_));
  NA2        u0820(.A(men_men_n791_), .B(men_men_n330_), .Y(men_men_n849_));
  NA2        u0821(.A(men_men_n339_), .B(men_men_n341_), .Y(men_men_n850_));
  OAI210     u0822(.A0(men_men_n199_), .A1(men_men_n209_), .B0(men_men_n850_), .Y(men_men_n851_));
  AOI220     u0823(.A0(men_men_n851_), .A1(men_men_n849_), .B0(men_men_n848_), .B1(men_men_n844_), .Y(men_men_n852_));
  NA2        u0824(.A(men_men_n164_), .B(men_men_n114_), .Y(men_men_n853_));
  NA2        u0825(.A(men_men_n853_), .B(men_men_n700_), .Y(men_men_n854_));
  NA3        u0826(.A(men_men_n854_), .B(men_men_n184_), .C(men_men_n31_), .Y(men_men_n855_));
  NA4        u0827(.A(men_men_n855_), .B(men_men_n852_), .C(men_men_n626_), .D(men_men_n82_), .Y(men_men_n856_));
  NO2        u0828(.A(men_men_n585_), .B(men_men_n492_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n857_), .B(men_men_n184_), .Y(men_men_n858_));
  NOi21      u0830(.An(f), .B(d), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n859_), .B(m), .Y(men_men_n860_));
  NO2        u0832(.A(men_men_n860_), .B(men_men_n50_), .Y(men_men_n861_));
  NOi32      u0833(.An(g), .Bn(f), .C(d), .Y(men_men_n862_));
  NA4        u0834(.A(men_men_n862_), .B(men_men_n605_), .C(men_men_n29_), .D(m), .Y(men_men_n863_));
  NOi21      u0835(.An(men_men_n308_), .B(men_men_n863_), .Y(men_men_n864_));
  AOI210     u0836(.A0(men_men_n861_), .A1(men_men_n541_), .B0(men_men_n864_), .Y(men_men_n865_));
  NA3        u0837(.A(men_men_n307_), .B(men_men_n254_), .C(men_men_n118_), .Y(men_men_n866_));
  AN2        u0838(.A(f), .B(d), .Y(men_men_n867_));
  NA3        u0839(.A(men_men_n476_), .B(men_men_n867_), .C(men_men_n84_), .Y(men_men_n868_));
  NO3        u0840(.A(men_men_n868_), .B(men_men_n73_), .C(men_men_n210_), .Y(men_men_n869_));
  NO2        u0841(.A(men_men_n280_), .B(men_men_n54_), .Y(men_men_n870_));
  NA2        u0842(.A(men_men_n866_), .B(men_men_n869_), .Y(men_men_n871_));
  NAi41      u0843(.An(men_men_n485_), .B(men_men_n871_), .C(men_men_n865_), .D(men_men_n858_), .Y(men_men_n872_));
  NO4        u0844(.A(men_men_n624_), .B(men_men_n131_), .C(men_men_n325_), .D(men_men_n148_), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n654_), .B(men_men_n325_), .Y(men_men_n874_));
  AN2        u0846(.A(men_men_n874_), .B(men_men_n682_), .Y(men_men_n875_));
  NO3        u0847(.A(men_men_n875_), .B(men_men_n873_), .C(men_men_n229_), .Y(men_men_n876_));
  NA2        u0848(.A(men_men_n603_), .B(men_men_n84_), .Y(men_men_n877_));
  NO2        u0849(.A(men_men_n850_), .B(men_men_n877_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n868_), .B(men_men_n428_), .Y(men_men_n879_));
  NOi41      u0851(.An(men_men_n218_), .B(men_men_n879_), .C(men_men_n878_), .D(men_men_n303_), .Y(men_men_n880_));
  NA2        u0852(.A(c), .B(men_men_n115_), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n881_), .B(men_men_n407_), .Y(men_men_n882_));
  NA3        u0854(.A(men_men_n882_), .B(men_men_n504_), .C(f), .Y(men_men_n883_));
  OR2        u0855(.A(men_men_n661_), .B(men_men_n537_), .Y(men_men_n884_));
  INV        u0856(.A(men_men_n884_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n808_), .B(men_men_n111_), .Y(men_men_n886_));
  NA2        u0858(.A(men_men_n886_), .B(men_men_n885_), .Y(men_men_n887_));
  NA4        u0859(.A(men_men_n887_), .B(men_men_n883_), .C(men_men_n880_), .D(men_men_n876_), .Y(men_men_n888_));
  NO4        u0860(.A(men_men_n888_), .B(men_men_n872_), .C(men_men_n856_), .D(men_men_n843_), .Y(men_men_n889_));
  OR2        u0861(.A(men_men_n868_), .B(men_men_n73_), .Y(men_men_n890_));
  NA2        u0862(.A(men_men_n832_), .B(g), .Y(men_men_n891_));
  AOI210     u0863(.A0(men_men_n891_), .A1(men_men_n288_), .B0(men_men_n890_), .Y(men_men_n892_));
  NO2        u0864(.A(men_men_n330_), .B(men_men_n840_), .Y(men_men_n893_));
  NO2        u0865(.A(men_men_n134_), .B(men_men_n131_), .Y(men_men_n894_));
  NO2        u0866(.A(men_men_n225_), .B(men_men_n219_), .Y(men_men_n895_));
  AOI220     u0867(.A0(men_men_n895_), .A1(men_men_n222_), .B0(men_men_n301_), .B1(men_men_n894_), .Y(men_men_n896_));
  NO2        u0868(.A(men_men_n428_), .B(men_men_n831_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n897_), .B(men_men_n558_), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n898_), .B(men_men_n896_), .Y(men_men_n899_));
  NA2        u0871(.A(e), .B(d), .Y(men_men_n900_));
  OAI220     u0872(.A0(men_men_n900_), .A1(c), .B0(men_men_n320_), .B1(d), .Y(men_men_n901_));
  NA3        u0873(.A(men_men_n901_), .B(men_men_n453_), .C(men_men_n502_), .Y(men_men_n902_));
  AOI210     u0874(.A0(men_men_n510_), .A1(men_men_n177_), .B0(men_men_n225_), .Y(men_men_n903_));
  INV        u0875(.A(men_men_n903_), .Y(men_men_n904_));
  NA2        u0876(.A(men_men_n280_), .B(men_men_n160_), .Y(men_men_n905_));
  NA2        u0877(.A(men_men_n869_), .B(men_men_n905_), .Y(men_men_n906_));
  NA3        u0878(.A(men_men_n163_), .B(men_men_n85_), .C(men_men_n34_), .Y(men_men_n907_));
  NA4        u0879(.A(men_men_n907_), .B(men_men_n906_), .C(men_men_n904_), .D(men_men_n902_), .Y(men_men_n908_));
  NO4        u0880(.A(men_men_n908_), .B(men_men_n899_), .C(men_men_n893_), .D(men_men_n892_), .Y(men_men_n909_));
  NA2        u0881(.A(men_men_n844_), .B(men_men_n31_), .Y(men_men_n910_));
  AO210      u0882(.A0(men_men_n910_), .A1(men_men_n702_), .B0(men_men_n213_), .Y(men_men_n911_));
  OAI220     u0883(.A0(men_men_n624_), .A1(men_men_n59_), .B0(men_men_n296_), .B1(j), .Y(men_men_n912_));
  AOI220     u0884(.A0(men_men_n912_), .A1(men_men_n874_), .B0(men_men_n614_), .B1(men_men_n623_), .Y(men_men_n913_));
  INV        u0885(.A(men_men_n913_), .Y(men_men_n914_));
  OAI210     u0886(.A0(men_men_n832_), .A1(men_men_n905_), .B0(men_men_n862_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n915_), .B(men_men_n606_), .Y(men_men_n916_));
  AOI210     u0888(.A0(men_men_n117_), .A1(men_men_n116_), .B0(men_men_n253_), .Y(men_men_n917_));
  AN2        u0889(.A(men_men_n849_), .B(men_men_n839_), .Y(men_men_n918_));
  NO3        u0890(.A(men_men_n918_), .B(men_men_n916_), .C(men_men_n914_), .Y(men_men_n919_));
  AO220      u0891(.A0(men_men_n453_), .A1(men_men_n752_), .B0(men_men_n172_), .B1(f), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n920_), .B(men_men_n901_), .Y(men_men_n921_));
  NO2        u0893(.A(men_men_n438_), .B(men_men_n69_), .Y(men_men_n922_));
  OAI210     u0894(.A0(men_men_n842_), .A1(men_men_n922_), .B0(men_men_n706_), .Y(men_men_n923_));
  AN4        u0895(.A(men_men_n923_), .B(men_men_n921_), .C(men_men_n919_), .D(men_men_n911_), .Y(men_men_n924_));
  NA4        u0896(.A(men_men_n924_), .B(men_men_n909_), .C(men_men_n889_), .D(men_men_n837_), .Y(men12));
  NO2        u0897(.A(men_men_n451_), .B(c), .Y(men_men_n926_));
  NO4        u0898(.A(men_men_n443_), .B(men_men_n245_), .C(men_men_n581_), .D(men_men_n210_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n927_), .B(men_men_n926_), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n541_), .B(men_men_n922_), .Y(men_men_n929_));
  NO2        u0901(.A(men_men_n451_), .B(men_men_n115_), .Y(men_men_n930_));
  NO2        u0902(.A(men_men_n845_), .B(men_men_n351_), .Y(men_men_n931_));
  NO2        u0903(.A(men_men_n661_), .B(men_men_n376_), .Y(men_men_n932_));
  AOI220     u0904(.A0(men_men_n932_), .A1(men_men_n539_), .B0(men_men_n931_), .B1(men_men_n930_), .Y(men_men_n933_));
  NA4        u0905(.A(men_men_n933_), .B(men_men_n929_), .C(men_men_n928_), .D(men_men_n442_), .Y(men_men_n934_));
  AOI210     u0906(.A0(men_men_n228_), .A1(men_men_n334_), .B0(men_men_n196_), .Y(men_men_n935_));
  OR2        u0907(.A(men_men_n935_), .B(men_men_n927_), .Y(men_men_n936_));
  NO2        u0908(.A(men_men_n388_), .B(men_men_n210_), .Y(men_men_n937_));
  OAI210     u0909(.A0(men_men_n937_), .A1(men_men_n936_), .B0(men_men_n402_), .Y(men_men_n938_));
  NO2        u0910(.A(men_men_n642_), .B(men_men_n256_), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n589_), .B(men_men_n838_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n940_), .B(men_men_n564_), .Y(men_men_n941_));
  NO2        u0913(.A(men_men_n147_), .B(men_men_n232_), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n942_), .B(men_men_n235_), .C(i), .Y(men_men_n943_));
  NA3        u0915(.A(men_men_n943_), .B(men_men_n941_), .C(men_men_n938_), .Y(men_men_n944_));
  NO3        u0916(.A(men_men_n131_), .B(men_men_n148_), .C(men_men_n210_), .Y(men_men_n945_));
  NA2        u0917(.A(men_men_n945_), .B(men_men_n526_), .Y(men_men_n946_));
  INV        u0918(.A(men_men_n946_), .Y(men_men_n947_));
  NO3        u0919(.A(men_men_n666_), .B(men_men_n92_), .C(men_men_n43_), .Y(men_men_n948_));
  NO4        u0920(.A(men_men_n948_), .B(men_men_n947_), .C(men_men_n944_), .D(men_men_n934_), .Y(men_men_n949_));
  NO2        u0921(.A(men_men_n367_), .B(men_men_n366_), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n586_), .B(men_men_n71_), .Y(men_men_n951_));
  NA2        u0923(.A(men_men_n551_), .B(men_men_n141_), .Y(men_men_n952_));
  NOi21      u0924(.An(men_men_n34_), .B(men_men_n654_), .Y(men_men_n953_));
  AOI220     u0925(.A0(men_men_n953_), .A1(men_men_n952_), .B0(men_men_n951_), .B1(men_men_n950_), .Y(men_men_n954_));
  OAI210     u0926(.A0(men_men_n244_), .A1(men_men_n43_), .B0(men_men_n954_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n434_), .B(men_men_n258_), .Y(men_men_n956_));
  NO3        u0928(.A(men_men_n819_), .B(men_men_n89_), .C(men_men_n407_), .Y(men_men_n957_));
  NAi31      u0929(.An(men_men_n957_), .B(men_men_n956_), .C(men_men_n318_), .Y(men_men_n958_));
  NO2        u0930(.A(men_men_n47_), .B(men_men_n43_), .Y(men_men_n959_));
  NO2        u0931(.A(men_men_n498_), .B(men_men_n296_), .Y(men_men_n960_));
  INV        u0932(.A(men_men_n960_), .Y(men_men_n961_));
  NO2        u0933(.A(men_men_n961_), .B(men_men_n141_), .Y(men_men_n962_));
  NA2        u0934(.A(men_men_n635_), .B(men_men_n361_), .Y(men_men_n963_));
  OAI210     u0935(.A0(men_men_n739_), .A1(men_men_n963_), .B0(men_men_n365_), .Y(men_men_n964_));
  NO4        u0936(.A(men_men_n964_), .B(men_men_n962_), .C(men_men_n958_), .D(men_men_n955_), .Y(men_men_n965_));
  NA2        u0937(.A(men_men_n344_), .B(g), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n157_), .B(i), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n44_), .B(i), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n968_), .B(men_men_n195_), .Y(men_men_n969_));
  AOI210     u0941(.A0(men_men_n418_), .A1(men_men_n37_), .B0(men_men_n969_), .Y(men_men_n970_));
  NO2        u0942(.A(men_men_n141_), .B(men_men_n84_), .Y(men_men_n971_));
  OR2        u0943(.A(men_men_n971_), .B(men_men_n550_), .Y(men_men_n972_));
  NA2        u0944(.A(men_men_n551_), .B(men_men_n380_), .Y(men_men_n973_));
  AOI210     u0945(.A0(men_men_n973_), .A1(n), .B0(men_men_n972_), .Y(men_men_n974_));
  OAI220     u0946(.A0(men_men_n974_), .A1(men_men_n966_), .B0(men_men_n970_), .B1(men_men_n330_), .Y(men_men_n975_));
  NO2        u0947(.A(men_men_n661_), .B(men_men_n492_), .Y(men_men_n976_));
  NA3        u0948(.A(men_men_n339_), .B(men_men_n630_), .C(i), .Y(men_men_n977_));
  OAI210     u0949(.A0(men_men_n438_), .A1(men_men_n307_), .B0(men_men_n977_), .Y(men_men_n978_));
  OAI220     u0950(.A0(men_men_n978_), .A1(men_men_n976_), .B0(men_men_n678_), .B1(men_men_n762_), .Y(men_men_n979_));
  NA2        u0951(.A(men_men_n608_), .B(men_men_n113_), .Y(men_men_n980_));
  OR3        u0952(.A(men_men_n307_), .B(men_men_n433_), .C(f), .Y(men_men_n981_));
  NA3        u0953(.A(men_men_n630_), .B(men_men_n80_), .C(i), .Y(men_men_n982_));
  OA220      u0954(.A0(men_men_n982_), .A1(men_men_n980_), .B0(men_men_n981_), .B1(men_men_n588_), .Y(men_men_n983_));
  NA3        u0955(.A(men_men_n322_), .B(men_men_n117_), .C(g), .Y(men_men_n984_));
  AOI210     u0956(.A0(men_men_n675_), .A1(men_men_n984_), .B0(m), .Y(men_men_n985_));
  OAI210     u0957(.A0(men_men_n985_), .A1(men_men_n931_), .B0(men_men_n321_), .Y(men_men_n986_));
  NA2        u0958(.A(men_men_n693_), .B(men_men_n877_), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n840_), .B(men_men_n439_), .Y(men_men_n988_));
  NA2        u0960(.A(men_men_n216_), .B(men_men_n77_), .Y(men_men_n989_));
  NA3        u0961(.A(men_men_n989_), .B(men_men_n982_), .C(men_men_n981_), .Y(men_men_n990_));
  AOI220     u0962(.A0(men_men_n990_), .A1(men_men_n251_), .B0(men_men_n988_), .B1(men_men_n987_), .Y(men_men_n991_));
  NA4        u0963(.A(men_men_n991_), .B(men_men_n986_), .C(men_men_n983_), .D(men_men_n979_), .Y(men_men_n992_));
  NO2        u0964(.A(men_men_n376_), .B(men_men_n91_), .Y(men_men_n993_));
  OAI210     u0965(.A0(men_men_n993_), .A1(men_men_n939_), .B0(men_men_n233_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n665_), .B(men_men_n88_), .Y(men_men_n995_));
  NO2        u0967(.A(men_men_n457_), .B(men_men_n210_), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n996_), .B(men_men_n381_), .Y(men_men_n997_));
  AOI220     u0969(.A0(men_men_n932_), .A1(men_men_n942_), .B0(men_men_n587_), .B1(men_men_n90_), .Y(men_men_n998_));
  NA4        u0970(.A(men_men_n998_), .B(men_men_n997_), .C(men_men_n995_), .D(men_men_n994_), .Y(men_men_n999_));
  OAI210     u0971(.A0(men_men_n988_), .A1(men_men_n940_), .B0(men_men_n539_), .Y(men_men_n1000_));
  AOI210     u0972(.A0(men_men_n419_), .A1(men_men_n411_), .B0(men_men_n819_), .Y(men_men_n1001_));
  INV        u0973(.A(men_men_n1001_), .Y(men_men_n1002_));
  NA2        u0974(.A(men_men_n985_), .B(men_men_n930_), .Y(men_men_n1003_));
  NA2        u0975(.A(men_men_n645_), .B(men_men_n526_), .Y(men_men_n1004_));
  NA4        u0976(.A(men_men_n1004_), .B(men_men_n1003_), .C(men_men_n1002_), .D(men_men_n1000_), .Y(men_men_n1005_));
  NO4        u0977(.A(men_men_n1005_), .B(men_men_n999_), .C(men_men_n992_), .D(men_men_n975_), .Y(men_men_n1006_));
  NAi31      u0978(.An(men_men_n138_), .B(men_men_n420_), .C(n), .Y(men_men_n1007_));
  NO3        u0979(.A(men_men_n125_), .B(men_men_n337_), .C(men_men_n846_), .Y(men_men_n1008_));
  NO2        u0980(.A(men_men_n1008_), .B(men_men_n1007_), .Y(men_men_n1009_));
  NO3        u0981(.A(men_men_n266_), .B(men_men_n138_), .C(men_men_n407_), .Y(men_men_n1010_));
  AOI210     u0982(.A0(men_men_n1010_), .A1(men_men_n493_), .B0(men_men_n1009_), .Y(men_men_n1011_));
  INV        u0983(.A(men_men_n1011_), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n225_), .B(men_men_n168_), .Y(men_men_n1013_));
  NO3        u0985(.A(men_men_n305_), .B(men_men_n444_), .C(men_men_n172_), .Y(men_men_n1014_));
  NOi31      u0986(.An(men_men_n1013_), .B(men_men_n1014_), .C(men_men_n210_), .Y(men_men_n1015_));
  NAi21      u0987(.An(men_men_n551_), .B(men_men_n996_), .Y(men_men_n1016_));
  NA2        u0988(.A(men_men_n437_), .B(men_men_n877_), .Y(men_men_n1017_));
  NO3        u0989(.A(men_men_n438_), .B(men_men_n307_), .C(men_men_n73_), .Y(men_men_n1018_));
  AOI220     u0990(.A0(men_men_n1018_), .A1(men_men_n1017_), .B0(men_men_n480_), .B1(g), .Y(men_men_n1019_));
  NA2        u0991(.A(men_men_n1019_), .B(men_men_n1016_), .Y(men_men_n1020_));
  OAI220     u0992(.A0(men_men_n1007_), .A1(men_men_n228_), .B0(men_men_n977_), .B1(men_men_n604_), .Y(men_men_n1021_));
  NO2        u0993(.A(men_men_n662_), .B(men_men_n376_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n935_), .B(men_men_n926_), .Y(men_men_n1023_));
  OAI220     u0995(.A0(men_men_n932_), .A1(men_men_n940_), .B0(men_men_n541_), .B1(men_men_n427_), .Y(men_men_n1024_));
  NA3        u0996(.A(men_men_n1024_), .B(men_men_n1023_), .C(men_men_n622_), .Y(men_men_n1025_));
  OAI210     u0997(.A0(men_men_n935_), .A1(men_men_n927_), .B0(men_men_n1013_), .Y(men_men_n1026_));
  NA3        u0998(.A(men_men_n973_), .B(men_men_n484_), .C(men_men_n44_), .Y(men_men_n1027_));
  AOI210     u0999(.A0(men_men_n379_), .A1(men_men_n377_), .B0(men_men_n329_), .Y(men_men_n1028_));
  NA4        u1000(.A(men_men_n1028_), .B(men_men_n1027_), .C(men_men_n1026_), .D(men_men_n267_), .Y(men_men_n1029_));
  OR4        u1001(.A(men_men_n1029_), .B(men_men_n1025_), .C(men_men_n1022_), .D(men_men_n1021_), .Y(men_men_n1030_));
  NO4        u1002(.A(men_men_n1030_), .B(men_men_n1020_), .C(men_men_n1015_), .D(men_men_n1012_), .Y(men_men_n1031_));
  NA4        u1003(.A(men_men_n1031_), .B(men_men_n1006_), .C(men_men_n965_), .D(men_men_n949_), .Y(men13));
  AN2        u1004(.A(c), .B(b), .Y(men_men_n1033_));
  NA3        u1005(.A(men_men_n243_), .B(men_men_n1033_), .C(m), .Y(men_men_n1034_));
  NA2        u1006(.A(d), .B(f), .Y(men_men_n1035_));
  NO4        u1007(.A(men_men_n1035_), .B(men_men_n1034_), .C(j), .D(men_men_n582_), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n258_), .B(men_men_n1033_), .Y(men_men_n1037_));
  NO4        u1009(.A(men_men_n1037_), .B(men_men_n1035_), .C(men_men_n967_), .D(a), .Y(men_men_n1038_));
  NAi32      u1010(.An(d), .Bn(c), .C(e), .Y(men_men_n1039_));
  NA2        u1011(.A(h), .B(men_men_n219_), .Y(men_men_n1040_));
  NA2        u1012(.A(men_men_n410_), .B(men_men_n209_), .Y(men_men_n1041_));
  AN2        u1013(.A(d), .B(c), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n1042_), .B(men_men_n115_), .Y(men_men_n1043_));
  NO4        u1015(.A(men_men_n1043_), .B(men_men_n1041_), .C(men_men_n173_), .D(men_men_n164_), .Y(men_men_n1044_));
  BUFFER     u1016(.A(men_men_n1044_), .Y(men_men_n1045_));
  OR3        u1017(.A(men_men_n1045_), .B(men_men_n1038_), .C(men_men_n1036_), .Y(men_men_n1046_));
  NAi32      u1018(.An(f), .Bn(e), .C(c), .Y(men_men_n1047_));
  NO2        u1019(.A(men_men_n1047_), .B(men_men_n143_), .Y(men_men_n1048_));
  NA2        u1020(.A(men_men_n1048_), .B(g), .Y(men_men_n1049_));
  OR3        u1021(.A(men_men_n219_), .B(men_men_n173_), .C(men_men_n164_), .Y(men_men_n1050_));
  NO2        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .Y(men_men_n1051_));
  NO2        u1023(.A(men_men_n766_), .B(men_men_n112_), .Y(men_men_n1052_));
  NOi41      u1024(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n1053_), .B(men_men_n1052_), .Y(men_men_n1054_));
  NO2        u1026(.A(men_men_n1054_), .B(men_men_n1049_), .Y(men_men_n1055_));
  OR3        u1027(.A(e), .B(d), .C(c), .Y(men_men_n1056_));
  NA3        u1028(.A(k), .B(j), .C(i), .Y(men_men_n1057_));
  NO3        u1029(.A(men_men_n1057_), .B(men_men_n304_), .C(men_men_n91_), .Y(men_men_n1058_));
  NOi21      u1030(.An(men_men_n1058_), .B(men_men_n1056_), .Y(men_men_n1059_));
  OR3        u1031(.A(men_men_n1059_), .B(men_men_n1055_), .C(men_men_n1051_), .Y(men_men_n1060_));
  NO2        u1032(.A(f), .B(c), .Y(men_men_n1061_));
  NOi21      u1033(.An(men_men_n1061_), .B(men_men_n443_), .Y(men_men_n1062_));
  NA2        u1034(.A(men_men_n1062_), .B(men_men_n57_), .Y(men_men_n1063_));
  OR2        u1035(.A(k), .B(i), .Y(men_men_n1064_));
  NO3        u1036(.A(men_men_n1064_), .B(men_men_n239_), .C(l), .Y(men_men_n1065_));
  NOi31      u1037(.An(men_men_n1065_), .B(men_men_n1063_), .C(j), .Y(men_men_n1066_));
  OR3        u1038(.A(men_men_n1066_), .B(men_men_n1060_), .C(men_men_n1046_), .Y(men02));
  OR2        u1039(.A(l), .B(k), .Y(men_men_n1068_));
  OR3        u1040(.A(h), .B(g), .C(f), .Y(men_men_n1069_));
  OR3        u1041(.A(n), .B(m), .C(i), .Y(men_men_n1070_));
  NO4        u1042(.A(men_men_n1070_), .B(men_men_n1069_), .C(men_men_n1068_), .D(men_men_n1056_), .Y(men_men_n1071_));
  NOi31      u1043(.An(e), .B(d), .C(c), .Y(men_men_n1072_));
  NA2        u1044(.A(men_men_n1058_), .B(men_men_n1072_), .Y(men_men_n1073_));
  AN3        u1045(.A(g), .B(f), .C(c), .Y(men_men_n1074_));
  NA2        u1046(.A(men_men_n1074_), .B(men_men_n465_), .Y(men_men_n1075_));
  OR2        u1047(.A(men_men_n1057_), .B(men_men_n304_), .Y(men_men_n1076_));
  OR2        u1048(.A(men_men_n1076_), .B(men_men_n1075_), .Y(men_men_n1077_));
  INV        u1049(.A(men_men_n1051_), .Y(men_men_n1078_));
  NA3        u1050(.A(l), .B(k), .C(j), .Y(men_men_n1079_));
  NA2        u1051(.A(i), .B(h), .Y(men_men_n1080_));
  NO3        u1052(.A(men_men_n1080_), .B(men_men_n1079_), .C(men_men_n131_), .Y(men_men_n1081_));
  NO3        u1053(.A(men_men_n139_), .B(men_men_n278_), .C(men_men_n210_), .Y(men_men_n1082_));
  NA3        u1054(.A(c), .B(b), .C(a), .Y(men_men_n1083_));
  NO3        u1055(.A(men_men_n1083_), .B(men_men_n900_), .C(men_men_n209_), .Y(men_men_n1084_));
  NO3        u1056(.A(men_men_n1057_), .B(men_men_n47_), .C(men_men_n112_), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n1085_), .B(men_men_n1084_), .Y(men_men_n1086_));
  AN3        u1058(.A(men_men_n1086_), .B(men_men_n1078_), .C(men_men_n1077_), .Y(men_men_n1087_));
  NO2        u1059(.A(men_men_n1043_), .B(men_men_n1041_), .Y(men_men_n1088_));
  NA2        u1060(.A(men_men_n1054_), .B(men_men_n1050_), .Y(men_men_n1089_));
  AOI210     u1061(.A0(men_men_n1089_), .A1(men_men_n1088_), .B0(men_men_n1036_), .Y(men_men_n1090_));
  NAi41      u1062(.An(men_men_n1071_), .B(men_men_n1090_), .C(men_men_n1087_), .D(men_men_n1073_), .Y(men03));
  NO2        u1063(.A(men_men_n522_), .B(men_men_n598_), .Y(men_men_n1092_));
  NA4        u1064(.A(men_men_n88_), .B(men_men_n87_), .C(g), .D(men_men_n209_), .Y(men_men_n1093_));
  NA4        u1065(.A(men_men_n573_), .B(m), .C(men_men_n112_), .D(men_men_n209_), .Y(men_men_n1094_));
  NA3        u1066(.A(men_men_n1094_), .B(men_men_n368_), .C(men_men_n1093_), .Y(men_men_n1095_));
  NO2        u1067(.A(men_men_n1095_), .B(men_men_n1092_), .Y(men_men_n1096_));
  NOi41      u1068(.An(men_men_n806_), .B(men_men_n851_), .C(men_men_n841_), .D(men_men_n720_), .Y(men_men_n1097_));
  OAI220     u1069(.A0(men_men_n1097_), .A1(men_men_n693_), .B0(men_men_n1096_), .B1(men_men_n586_), .Y(men_men_n1098_));
  NOi31      u1070(.An(i), .B(k), .C(j), .Y(men_men_n1099_));
  NA4        u1071(.A(men_men_n1099_), .B(men_men_n1072_), .C(men_men_n339_), .D(men_men_n332_), .Y(men_men_n1100_));
  OAI210     u1072(.A0(men_men_n819_), .A1(men_men_n421_), .B0(men_men_n1100_), .Y(men_men_n1101_));
  NOi31      u1073(.An(m), .B(n), .C(f), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n1102_), .B(men_men_n49_), .Y(men_men_n1103_));
  NO2        u1075(.A(men_men_n884_), .B(men_men_n426_), .Y(men_men_n1104_));
  NA2        u1076(.A(men_men_n502_), .B(l), .Y(men_men_n1105_));
  NOi31      u1077(.An(men_men_n862_), .B(men_men_n1034_), .C(men_men_n1105_), .Y(men_men_n1106_));
  NO4        u1078(.A(men_men_n1106_), .B(men_men_n1104_), .C(men_men_n1101_), .D(men_men_n1001_), .Y(men_men_n1107_));
  NO2        u1079(.A(men_men_n278_), .B(a), .Y(men_men_n1108_));
  NO2        u1080(.A(men_men_n1080_), .B(men_men_n483_), .Y(men_men_n1109_));
  NO2        u1081(.A(men_men_n87_), .B(g), .Y(men_men_n1110_));
  AOI210     u1082(.A0(men_men_n1110_), .A1(men_men_n1109_), .B0(men_men_n1065_), .Y(men_men_n1111_));
  OR2        u1083(.A(men_men_n1111_), .B(men_men_n1063_), .Y(men_men_n1112_));
  NA2        u1084(.A(men_men_n1112_), .B(men_men_n1107_), .Y(men_men_n1113_));
  NO4        u1085(.A(men_men_n1113_), .B(men_men_n1098_), .C(men_men_n820_), .D(men_men_n563_), .Y(men_men_n1114_));
  NA2        u1086(.A(c), .B(b), .Y(men_men_n1115_));
  NO2        u1087(.A(men_men_n705_), .B(men_men_n1115_), .Y(men_men_n1116_));
  OAI210     u1088(.A0(men_men_n860_), .A1(men_men_n835_), .B0(men_men_n414_), .Y(men_men_n1117_));
  OAI210     u1089(.A0(men_men_n1117_), .A1(men_men_n861_), .B0(men_men_n1116_), .Y(men_men_n1118_));
  NAi21      u1090(.An(men_men_n422_), .B(men_men_n1116_), .Y(men_men_n1119_));
  OAI210     u1091(.A0(men_men_n545_), .A1(men_men_n39_), .B0(men_men_n1108_), .Y(men_men_n1120_));
  NA2        u1092(.A(men_men_n1120_), .B(men_men_n1119_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n254_), .B(men_men_n118_), .Y(men_men_n1122_));
  OAI210     u1094(.A0(men_men_n1122_), .A1(men_men_n282_), .B0(g), .Y(men_men_n1123_));
  NAi21      u1095(.An(f), .B(d), .Y(men_men_n1124_));
  NO2        u1096(.A(men_men_n1124_), .B(men_men_n1083_), .Y(men_men_n1125_));
  INV        u1097(.A(men_men_n1125_), .Y(men_men_n1126_));
  AOI210     u1098(.A0(men_men_n1123_), .A1(men_men_n288_), .B0(men_men_n1126_), .Y(men_men_n1127_));
  AOI210     u1099(.A0(men_men_n1127_), .A1(men_men_n113_), .B0(men_men_n1121_), .Y(men_men_n1128_));
  NA2        u1100(.A(men_men_n468_), .B(men_men_n467_), .Y(men_men_n1129_));
  NO2        u1101(.A(men_men_n179_), .B(men_men_n232_), .Y(men_men_n1130_));
  NA2        u1102(.A(men_men_n1130_), .B(m), .Y(men_men_n1131_));
  NA3        u1103(.A(men_men_n917_), .B(men_men_n1105_), .C(men_men_n471_), .Y(men_men_n1132_));
  OAI210     u1104(.A0(men_men_n1132_), .A1(men_men_n308_), .B0(men_men_n469_), .Y(men_men_n1133_));
  AOI210     u1105(.A0(men_men_n1133_), .A1(men_men_n1129_), .B0(men_men_n1131_), .Y(men_men_n1134_));
  NA2        u1106(.A(men_men_n558_), .B(men_men_n409_), .Y(men_men_n1135_));
  NO2        u1107(.A(men_men_n963_), .B(men_men_n210_), .Y(men_men_n1136_));
  OAI210     u1108(.A0(men_men_n1136_), .A1(men_men_n447_), .B0(men_men_n1125_), .Y(men_men_n1137_));
  NO2        u1109(.A(men_men_n370_), .B(men_men_n369_), .Y(men_men_n1138_));
  AOI210     u1110(.A0(men_men_n1130_), .A1(men_men_n429_), .B0(men_men_n957_), .Y(men_men_n1139_));
  NAi41      u1111(.An(men_men_n1138_), .B(men_men_n1139_), .C(men_men_n1137_), .D(men_men_n1135_), .Y(men_men_n1140_));
  NO2        u1112(.A(men_men_n1140_), .B(men_men_n1134_), .Y(men_men_n1141_));
  NA4        u1113(.A(men_men_n1141_), .B(men_men_n1128_), .C(men_men_n1118_), .D(men_men_n1114_), .Y(men00));
  AOI210     u1114(.A0(men_men_n295_), .A1(men_men_n210_), .B0(men_men_n270_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n1143_), .B(men_men_n576_), .Y(men_men_n1144_));
  AOI210     u1116(.A0(men_men_n897_), .A1(men_men_n942_), .B0(men_men_n1101_), .Y(men_men_n1145_));
  NO2        u1117(.A(men_men_n957_), .B(men_men_n717_), .Y(men_men_n1146_));
  NA3        u1118(.A(men_men_n1146_), .B(men_men_n1145_), .C(men_men_n1002_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n504_), .B(f), .Y(men_men_n1148_));
  OAI210     u1120(.A0(men_men_n1008_), .A1(men_men_n40_), .B0(men_men_n647_), .Y(men_men_n1149_));
  NA3        u1121(.A(men_men_n1149_), .B(men_men_n250_), .C(n), .Y(men_men_n1150_));
  AOI210     u1122(.A0(men_men_n1150_), .A1(men_men_n1148_), .B0(men_men_n1043_), .Y(men_men_n1151_));
  NO4        u1123(.A(men_men_n1151_), .B(men_men_n1147_), .C(men_men_n1144_), .D(men_men_n1060_), .Y(men_men_n1152_));
  NA3        u1124(.A(men_men_n163_), .B(men_men_n44_), .C(men_men_n43_), .Y(men_men_n1153_));
  NA3        u1125(.A(d), .B(men_men_n54_), .C(b), .Y(men_men_n1154_));
  NOi31      u1126(.An(n), .B(m), .C(i), .Y(men_men_n1155_));
  NA3        u1127(.A(men_men_n1155_), .B(men_men_n650_), .C(men_men_n49_), .Y(men_men_n1156_));
  OAI210     u1128(.A0(men_men_n1154_), .A1(men_men_n1153_), .B0(men_men_n1156_), .Y(men_men_n1157_));
  INV        u1129(.A(men_men_n575_), .Y(men_men_n1158_));
  NO3        u1130(.A(men_men_n1158_), .B(men_men_n1157_), .C(men_men_n1138_), .Y(men_men_n1159_));
  NA3        u1131(.A(men_men_n382_), .B(men_men_n215_), .C(g), .Y(men_men_n1160_));
  NO2        u1132(.A(h), .B(g), .Y(men_men_n1161_));
  NA4        u1133(.A(men_men_n493_), .B(men_men_n465_), .C(men_men_n1161_), .D(men_men_n1033_), .Y(men_men_n1162_));
  NA2        u1134(.A(men_men_n945_), .B(men_men_n574_), .Y(men_men_n1163_));
  NA2        u1135(.A(men_men_n1163_), .B(men_men_n1162_), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n1164_), .B(men_men_n260_), .Y(men_men_n1165_));
  NO2        u1137(.A(men_men_n234_), .B(men_men_n178_), .Y(men_men_n1166_));
  NA2        u1138(.A(men_men_n1166_), .B(men_men_n427_), .Y(men_men_n1167_));
  NA3        u1139(.A(men_men_n176_), .B(men_men_n112_), .C(g), .Y(men_men_n1168_));
  NA3        u1140(.A(men_men_n465_), .B(men_men_n40_), .C(f), .Y(men_men_n1169_));
  NOi31      u1141(.An(men_men_n870_), .B(men_men_n1169_), .C(men_men_n1168_), .Y(men_men_n1170_));
  NAi31      u1142(.An(men_men_n180_), .B(men_men_n857_), .C(men_men_n465_), .Y(men_men_n1171_));
  NAi31      u1143(.An(men_men_n1170_), .B(men_men_n1171_), .C(men_men_n1167_), .Y(men_men_n1172_));
  NO2        u1144(.A(men_men_n269_), .B(men_men_n73_), .Y(men_men_n1173_));
  NO3        u1145(.A(men_men_n426_), .B(men_men_n831_), .C(n), .Y(men_men_n1174_));
  AOI210     u1146(.A0(men_men_n1174_), .A1(men_men_n1173_), .B0(men_men_n1071_), .Y(men_men_n1175_));
  NA2        u1147(.A(men_men_n1175_), .B(men_men_n72_), .Y(men_men_n1176_));
  NO4        u1148(.A(men_men_n1176_), .B(men_men_n1172_), .C(men_men_n577_), .D(men_men_n513_), .Y(men_men_n1177_));
  AN3        u1149(.A(men_men_n1177_), .B(men_men_n1165_), .C(men_men_n1159_), .Y(men_men_n1178_));
  NA2        u1150(.A(men_men_n531_), .B(men_men_n102_), .Y(men_men_n1179_));
  NA3        u1151(.A(men_men_n1102_), .B(men_men_n608_), .C(men_men_n464_), .Y(men_men_n1180_));
  NA4        u1152(.A(men_men_n1180_), .B(men_men_n559_), .C(men_men_n1179_), .D(men_men_n237_), .Y(men_men_n1181_));
  NA2        u1153(.A(men_men_n1095_), .B(men_men_n531_), .Y(men_men_n1182_));
  NA4        u1154(.A(men_men_n650_), .B(men_men_n201_), .C(men_men_n215_), .D(men_men_n157_), .Y(men_men_n1183_));
  NA3        u1155(.A(men_men_n1183_), .B(men_men_n1182_), .C(men_men_n292_), .Y(men_men_n1184_));
  OAI210     u1156(.A0(men_men_n463_), .A1(men_men_n119_), .B0(men_men_n863_), .Y(men_men_n1185_));
  AOI220     u1157(.A0(men_men_n1185_), .A1(men_men_n1132_), .B0(men_men_n558_), .B1(men_men_n409_), .Y(men_men_n1186_));
  OR4        u1158(.A(men_men_n1043_), .B(men_men_n266_), .C(men_men_n217_), .D(e), .Y(men_men_n1187_));
  NO2        u1159(.A(men_men_n213_), .B(men_men_n210_), .Y(men_men_n1188_));
  NA2        u1160(.A(n), .B(e), .Y(men_men_n1189_));
  NO2        u1161(.A(men_men_n1189_), .B(men_men_n143_), .Y(men_men_n1190_));
  AOI220     u1162(.A0(men_men_n1190_), .A1(men_men_n268_), .B0(men_men_n844_), .B1(men_men_n1188_), .Y(men_men_n1191_));
  OAI210     u1163(.A0(men_men_n355_), .A1(men_men_n309_), .B0(men_men_n449_), .Y(men_men_n1192_));
  NA4        u1164(.A(men_men_n1192_), .B(men_men_n1191_), .C(men_men_n1187_), .D(men_men_n1186_), .Y(men_men_n1193_));
  AOI210     u1165(.A0(men_men_n1190_), .A1(men_men_n848_), .B0(men_men_n820_), .Y(men_men_n1194_));
  AOI220     u1166(.A0(men_men_n953_), .A1(men_men_n574_), .B0(men_men_n650_), .B1(men_men_n240_), .Y(men_men_n1195_));
  NO2        u1167(.A(men_men_n66_), .B(h), .Y(men_men_n1196_));
  NO3        u1168(.A(men_men_n1043_), .B(men_men_n1041_), .C(men_men_n731_), .Y(men_men_n1197_));
  INV        u1169(.A(men_men_n131_), .Y(men_men_n1198_));
  AN2        u1170(.A(men_men_n1198_), .B(men_men_n1082_), .Y(men_men_n1199_));
  OAI210     u1171(.A0(men_men_n1199_), .A1(men_men_n1197_), .B0(men_men_n1196_), .Y(men_men_n1200_));
  NA4        u1172(.A(men_men_n1200_), .B(men_men_n1195_), .C(men_men_n1194_), .D(men_men_n865_), .Y(men_men_n1201_));
  NO4        u1173(.A(men_men_n1201_), .B(men_men_n1193_), .C(men_men_n1184_), .D(men_men_n1181_), .Y(men_men_n1202_));
  NA2        u1174(.A(men_men_n836_), .B(men_men_n761_), .Y(men_men_n1203_));
  NA4        u1175(.A(men_men_n1203_), .B(men_men_n1202_), .C(men_men_n1178_), .D(men_men_n1152_), .Y(men01));
  NO3        u1176(.A(men_men_n802_), .B(men_men_n794_), .C(men_men_n276_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n393_), .B(i), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n1206_), .B(men_men_n1205_), .C(men_men_n1023_), .Y(men_men_n1207_));
  NA2        u1179(.A(men_men_n587_), .B(men_men_n90_), .Y(men_men_n1208_));
  NA2        u1180(.A(men_men_n551_), .B(men_men_n265_), .Y(men_men_n1209_));
  NA2        u1181(.A(men_men_n960_), .B(men_men_n1209_), .Y(men_men_n1210_));
  NA4        u1182(.A(men_men_n1210_), .B(men_men_n1208_), .C(men_men_n913_), .D(men_men_n331_), .Y(men_men_n1211_));
  NA2        u1183(.A(men_men_n43_), .B(f), .Y(men_men_n1212_));
  NA2        u1184(.A(men_men_n712_), .B(men_men_n97_), .Y(men_men_n1213_));
  NO2        u1185(.A(men_men_n1213_), .B(men_men_n1212_), .Y(men_men_n1214_));
  OAI210     u1186(.A0(men_men_n783_), .A1(men_men_n604_), .B0(men_men_n1183_), .Y(men_men_n1215_));
  AOI210     u1187(.A0(men_men_n1214_), .A1(men_men_n637_), .B0(men_men_n1215_), .Y(men_men_n1216_));
  INV        u1188(.A(men_men_n117_), .Y(men_men_n1217_));
  OA220      u1189(.A0(men_men_n1217_), .A1(men_men_n584_), .B0(men_men_n663_), .B1(men_men_n368_), .Y(men_men_n1218_));
  NAi41      u1190(.An(men_men_n156_), .B(men_men_n1218_), .C(men_men_n1216_), .D(men_men_n896_), .Y(men_men_n1219_));
  NO3        u1191(.A(men_men_n784_), .B(men_men_n677_), .C(men_men_n507_), .Y(men_men_n1220_));
  NA4        u1192(.A(men_men_n712_), .B(men_men_n97_), .C(men_men_n43_), .D(men_men_n209_), .Y(men_men_n1221_));
  OA220      u1193(.A0(men_men_n1221_), .A1(men_men_n671_), .B0(men_men_n190_), .B1(men_men_n188_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n1222_), .B(men_men_n1220_), .Y(men_men_n1223_));
  NO4        u1195(.A(men_men_n1223_), .B(men_men_n1219_), .C(men_men_n1211_), .D(men_men_n1207_), .Y(men_men_n1224_));
  INV        u1196(.A(men_men_n1160_), .Y(men_men_n1225_));
  OAI210     u1197(.A0(men_men_n1225_), .A1(men_men_n298_), .B0(men_men_n526_), .Y(men_men_n1226_));
  NA2        u1198(.A(men_men_n534_), .B(men_men_n395_), .Y(men_men_n1227_));
  NOi21      u1199(.An(men_men_n560_), .B(men_men_n581_), .Y(men_men_n1228_));
  NA2        u1200(.A(men_men_n1228_), .B(men_men_n1227_), .Y(men_men_n1229_));
  AOI210     u1201(.A0(men_men_n199_), .A1(men_men_n89_), .B0(men_men_n209_), .Y(men_men_n1230_));
  OAI210     u1202(.A0(men_men_n809_), .A1(men_men_n427_), .B0(men_men_n1230_), .Y(men_men_n1231_));
  AN3        u1203(.A(m), .B(l), .C(k), .Y(men_men_n1232_));
  OAI210     u1204(.A0(men_men_n357_), .A1(men_men_n34_), .B0(men_men_n1232_), .Y(men_men_n1233_));
  NA2        u1205(.A(men_men_n198_), .B(men_men_n34_), .Y(men_men_n1234_));
  AO210      u1206(.A0(men_men_n1234_), .A1(men_men_n1233_), .B0(men_men_n330_), .Y(men_men_n1235_));
  NA4        u1207(.A(men_men_n1235_), .B(men_men_n1231_), .C(men_men_n1229_), .D(men_men_n1226_), .Y(men_men_n1236_));
  AOI210     u1208(.A0(men_men_n596_), .A1(men_men_n117_), .B0(men_men_n602_), .Y(men_men_n1237_));
  OAI210     u1209(.A0(men_men_n1217_), .A1(men_men_n593_), .B0(men_men_n1237_), .Y(men_men_n1238_));
  NA2        u1210(.A(men_men_n275_), .B(men_men_n190_), .Y(men_men_n1239_));
  NA2        u1211(.A(men_men_n1239_), .B(men_men_n668_), .Y(men_men_n1240_));
  NO3        u1212(.A(men_men_n819_), .B(men_men_n199_), .C(men_men_n407_), .Y(men_men_n1241_));
  NO2        u1213(.A(men_men_n1241_), .B(men_men_n957_), .Y(men_men_n1242_));
  OAI210     u1214(.A0(men_men_n1214_), .A1(men_men_n324_), .B0(men_men_n678_), .Y(men_men_n1243_));
  NA4        u1215(.A(men_men_n1243_), .B(men_men_n1242_), .C(men_men_n1240_), .D(men_men_n787_), .Y(men_men_n1244_));
  NO3        u1216(.A(men_men_n1244_), .B(men_men_n1238_), .C(men_men_n1236_), .Y(men_men_n1245_));
  NA3        u1217(.A(men_men_n605_), .B(men_men_n29_), .C(f), .Y(men_men_n1246_));
  NO2        u1218(.A(men_men_n1246_), .B(men_men_n199_), .Y(men_men_n1247_));
  AOI210     u1219(.A0(men_men_n499_), .A1(men_men_n56_), .B0(men_men_n1247_), .Y(men_men_n1248_));
  NO2        u1220(.A(men_men_n1221_), .B(men_men_n980_), .Y(men_men_n1249_));
  NO2        u1221(.A(men_men_n202_), .B(men_men_n111_), .Y(men_men_n1250_));
  NO3        u1222(.A(men_men_n1250_), .B(men_men_n1249_), .C(men_men_n1157_), .Y(men_men_n1251_));
  NA3        u1223(.A(men_men_n1251_), .B(men_men_n1248_), .C(men_men_n760_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n967_), .B(men_men_n227_), .Y(men_men_n1253_));
  NO2        u1225(.A(men_men_n968_), .B(men_men_n553_), .Y(men_men_n1254_));
  OAI210     u1226(.A0(men_men_n1254_), .A1(men_men_n1253_), .B0(men_men_n337_), .Y(men_men_n1255_));
  NO3        u1227(.A(men_men_n79_), .B(men_men_n296_), .C(men_men_n43_), .Y(men_men_n1256_));
  NA2        u1228(.A(men_men_n1256_), .B(men_men_n550_), .Y(men_men_n1257_));
  NA2        u1229(.A(men_men_n1257_), .B(men_men_n673_), .Y(men_men_n1258_));
  NO2        u1230(.A(men_men_n368_), .B(men_men_n71_), .Y(men_men_n1259_));
  INV        u1231(.A(men_men_n1259_), .Y(men_men_n1260_));
  NA2        u1232(.A(men_men_n1256_), .B(men_men_n812_), .Y(men_men_n1261_));
  NA3        u1233(.A(men_men_n1261_), .B(men_men_n1260_), .C(men_men_n385_), .Y(men_men_n1262_));
  NOi41      u1234(.An(men_men_n1255_), .B(men_men_n1262_), .C(men_men_n1258_), .D(men_men_n1252_), .Y(men_men_n1263_));
  NO2        u1235(.A(men_men_n130_), .B(men_men_n43_), .Y(men_men_n1264_));
  NO2        u1236(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n1265_));
  AO220      u1237(.A0(men_men_n1265_), .A1(men_men_n625_), .B0(men_men_n1264_), .B1(men_men_n710_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n1266_), .B(men_men_n337_), .Y(men_men_n1267_));
  NO3        u1239(.A(men_men_n1080_), .B(men_men_n173_), .C(men_men_n87_), .Y(men_men_n1268_));
  NA2        u1240(.A(men_men_n1256_), .B(men_men_n971_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n1267_), .Y(men_men_n1270_));
  NO2        u1242(.A(men_men_n616_), .B(men_men_n615_), .Y(men_men_n1271_));
  NO4        u1243(.A(men_men_n1080_), .B(men_men_n1271_), .C(men_men_n171_), .D(men_men_n87_), .Y(men_men_n1272_));
  NO3        u1244(.A(men_men_n1272_), .B(men_men_n1270_), .C(men_men_n641_), .Y(men_men_n1273_));
  NA4        u1245(.A(men_men_n1273_), .B(men_men_n1263_), .C(men_men_n1245_), .D(men_men_n1224_), .Y(men06));
  NO2        u1246(.A(men_men_n408_), .B(men_men_n557_), .Y(men_men_n1275_));
  INV        u1247(.A(men_men_n738_), .Y(men_men_n1276_));
  OAI210     u1248(.A0(men_men_n1276_), .A1(men_men_n261_), .B0(men_men_n1275_), .Y(men_men_n1277_));
  NO2        u1249(.A(men_men_n219_), .B(men_men_n104_), .Y(men_men_n1278_));
  OAI210     u1250(.A0(men_men_n1278_), .A1(men_men_n1268_), .B0(men_men_n381_), .Y(men_men_n1279_));
  NO3        u1251(.A(men_men_n600_), .B(men_men_n807_), .C(men_men_n603_), .Y(men_men_n1280_));
  OR2        u1252(.A(men_men_n1280_), .B(men_men_n884_), .Y(men_men_n1281_));
  NA4        u1253(.A(men_men_n1281_), .B(men_men_n1279_), .C(men_men_n1277_), .D(men_men_n1255_), .Y(men_men_n1282_));
  NO3        u1254(.A(men_men_n1282_), .B(men_men_n1258_), .C(men_men_n249_), .Y(men_men_n1283_));
  NO2        u1255(.A(men_men_n296_), .B(men_men_n43_), .Y(men_men_n1284_));
  AOI210     u1256(.A0(men_men_n1284_), .A1(men_men_n972_), .B0(men_men_n1253_), .Y(men_men_n1285_));
  AOI210     u1257(.A0(men_men_n1284_), .A1(men_men_n554_), .B0(men_men_n1266_), .Y(men_men_n1286_));
  AOI210     u1258(.A0(men_men_n1286_), .A1(men_men_n1285_), .B0(men_men_n334_), .Y(men_men_n1287_));
  OAI210     u1259(.A0(men_men_n89_), .A1(men_men_n40_), .B0(men_men_n676_), .Y(men_men_n1288_));
  NA2        u1260(.A(men_men_n1288_), .B(men_men_n644_), .Y(men_men_n1289_));
  NO2        u1261(.A(men_men_n510_), .B(men_men_n168_), .Y(men_men_n1290_));
  NO2        u1262(.A(men_men_n609_), .B(men_men_n1103_), .Y(men_men_n1291_));
  OAI210     u1263(.A0(men_men_n458_), .A1(men_men_n242_), .B0(men_men_n907_), .Y(men_men_n1292_));
  NO3        u1264(.A(men_men_n1292_), .B(men_men_n1291_), .C(men_men_n1290_), .Y(men_men_n1293_));
  OR2        u1265(.A(men_men_n601_), .B(men_men_n599_), .Y(men_men_n1294_));
  NO2        u1266(.A(men_men_n367_), .B(men_men_n134_), .Y(men_men_n1295_));
  AOI210     u1267(.A0(men_men_n1295_), .A1(men_men_n587_), .B0(men_men_n1294_), .Y(men_men_n1296_));
  NA3        u1268(.A(men_men_n1296_), .B(men_men_n1293_), .C(men_men_n1289_), .Y(men_men_n1297_));
  NO2        u1269(.A(men_men_n753_), .B(men_men_n366_), .Y(men_men_n1298_));
  NO3        u1270(.A(men_men_n678_), .B(men_men_n762_), .C(men_men_n637_), .Y(men_men_n1299_));
  NOi21      u1271(.An(men_men_n1298_), .B(men_men_n1299_), .Y(men_men_n1300_));
  AN2        u1272(.A(men_men_n953_), .B(men_men_n646_), .Y(men_men_n1301_));
  NO4        u1273(.A(men_men_n1301_), .B(men_men_n1300_), .C(men_men_n1297_), .D(men_men_n1287_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n801_), .B(men_men_n271_), .Y(men_men_n1303_));
  OAI220     u1275(.A0(men_men_n738_), .A1(men_men_n45_), .B0(men_men_n219_), .B1(men_men_n618_), .Y(men_men_n1304_));
  OAI210     u1276(.A0(men_men_n271_), .A1(c), .B0(men_men_n643_), .Y(men_men_n1305_));
  AOI220     u1277(.A0(men_men_n1305_), .A1(men_men_n1304_), .B0(men_men_n1303_), .B1(men_men_n261_), .Y(men_men_n1306_));
  NO3        u1278(.A(men_men_n239_), .B(men_men_n104_), .C(men_men_n278_), .Y(men_men_n1307_));
  OAI220     u1279(.A0(men_men_n702_), .A1(men_men_n242_), .B0(men_men_n506_), .B1(men_men_n510_), .Y(men_men_n1308_));
  NO3        u1280(.A(men_men_n1308_), .B(men_men_n1307_), .C(men_men_n1104_), .Y(men_men_n1309_));
  NA4        u1281(.A(men_men_n792_), .B(men_men_n791_), .C(men_men_n437_), .D(men_men_n877_), .Y(men_men_n1310_));
  NAi31      u1282(.An(men_men_n753_), .B(men_men_n1310_), .C(men_men_n198_), .Y(men_men_n1311_));
  NA4        u1283(.A(men_men_n1311_), .B(men_men_n1309_), .C(men_men_n1306_), .D(men_men_n1195_), .Y(men_men_n1312_));
  NOi31      u1284(.An(men_men_n1280_), .B(men_men_n462_), .C(men_men_n394_), .Y(men_men_n1313_));
  OR3        u1285(.A(men_men_n1313_), .B(men_men_n783_), .C(men_men_n537_), .Y(men_men_n1314_));
  OR3        u1286(.A(men_men_n369_), .B(men_men_n219_), .C(men_men_n618_), .Y(men_men_n1315_));
  AOI210     u1287(.A0(men_men_n569_), .A1(men_men_n449_), .B0(men_men_n371_), .Y(men_men_n1316_));
  NA3        u1288(.A(men_men_n1316_), .B(men_men_n1315_), .C(men_men_n1314_), .Y(men_men_n1317_));
  AOI220     u1289(.A0(men_men_n1298_), .A1(men_men_n761_), .B0(men_men_n1295_), .B1(men_men_n233_), .Y(men_men_n1318_));
  AN2        u1290(.A(men_men_n927_), .B(men_men_n926_), .Y(men_men_n1319_));
  NO4        u1291(.A(men_men_n1319_), .B(men_men_n875_), .C(men_men_n495_), .D(men_men_n480_), .Y(men_men_n1320_));
  NA3        u1292(.A(men_men_n1320_), .B(men_men_n1318_), .C(men_men_n1261_), .Y(men_men_n1321_));
  NAi21      u1293(.An(j), .B(i), .Y(men_men_n1322_));
  NO4        u1294(.A(men_men_n1271_), .B(men_men_n1322_), .C(men_men_n443_), .D(men_men_n230_), .Y(men_men_n1323_));
  NO4        u1295(.A(men_men_n1323_), .B(men_men_n1321_), .C(men_men_n1317_), .D(men_men_n1312_), .Y(men_men_n1324_));
  NA4        u1296(.A(men_men_n1324_), .B(men_men_n1302_), .C(men_men_n1283_), .D(men_men_n1273_), .Y(men07));
  NAi32      u1297(.An(m), .Bn(b), .C(n), .Y(men_men_n1326_));
  NO3        u1298(.A(men_men_n1326_), .B(g), .C(f), .Y(men_men_n1327_));
  OAI210     u1299(.A0(men_men_n319_), .A1(men_men_n482_), .B0(men_men_n1327_), .Y(men_men_n1328_));
  NAi21      u1300(.An(f), .B(c), .Y(men_men_n1329_));
  OR2        u1301(.A(e), .B(d), .Y(men_men_n1330_));
  OAI220     u1302(.A0(men_men_n1330_), .A1(men_men_n1329_), .B0(men_men_n631_), .B1(men_men_n320_), .Y(men_men_n1331_));
  NA3        u1303(.A(men_men_n1331_), .B(men_men_n1505_), .C(men_men_n176_), .Y(men_men_n1332_));
  NOi31      u1304(.An(n), .B(m), .C(b), .Y(men_men_n1333_));
  NO3        u1305(.A(men_men_n131_), .B(men_men_n450_), .C(h), .Y(men_men_n1334_));
  NA2        u1306(.A(men_men_n1332_), .B(men_men_n1328_), .Y(men_men_n1335_));
  NOi41      u1307(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1336_));
  NA2        u1308(.A(men_men_n1082_), .B(men_men_n215_), .Y(men_men_n1337_));
  NO2        u1309(.A(men_men_n1337_), .B(men_men_n59_), .Y(men_men_n1338_));
  NO2        u1310(.A(k), .B(i), .Y(men_men_n1339_));
  NO2        u1311(.A(men_men_n1057_), .B(men_men_n304_), .Y(men_men_n1340_));
  NA2        u1312(.A(men_men_n538_), .B(men_men_n80_), .Y(men_men_n1341_));
  NA2        u1313(.A(men_men_n1196_), .B(men_men_n286_), .Y(men_men_n1342_));
  NA2        u1314(.A(men_men_n1342_), .B(men_men_n1341_), .Y(men_men_n1343_));
  NO3        u1315(.A(men_men_n1343_), .B(men_men_n1338_), .C(men_men_n1335_), .Y(men_men_n1344_));
  NO3        u1316(.A(e), .B(d), .C(c), .Y(men_men_n1345_));
  NO2        u1317(.A(men_men_n131_), .B(men_men_n210_), .Y(men_men_n1346_));
  NA2        u1318(.A(men_men_n1346_), .B(men_men_n1345_), .Y(men_men_n1347_));
  NO2        u1319(.A(men_men_n1347_), .B(c), .Y(men_men_n1348_));
  OR2        u1320(.A(h), .B(f), .Y(men_men_n1349_));
  NO3        u1321(.A(n), .B(m), .C(i), .Y(men_men_n1350_));
  NA2        u1322(.A(g), .B(men_men_n1350_), .Y(men_men_n1351_));
  NO2        u1323(.A(i), .B(g), .Y(men_men_n1352_));
  OR3        u1324(.A(men_men_n1352_), .B(men_men_n1326_), .C(men_men_n70_), .Y(men_men_n1353_));
  OAI220     u1325(.A0(men_men_n1353_), .A1(men_men_n482_), .B0(men_men_n1351_), .B1(men_men_n1349_), .Y(men_men_n1354_));
  NA3        u1326(.A(men_men_n699_), .B(men_men_n686_), .C(men_men_n112_), .Y(men_men_n1355_));
  NO2        u1327(.A(men_men_n1355_), .B(men_men_n43_), .Y(men_men_n1356_));
  NO2        u1328(.A(l), .B(k), .Y(men_men_n1357_));
  NOi41      u1329(.An(men_men_n543_), .B(men_men_n1357_), .C(men_men_n477_), .D(men_men_n443_), .Y(men_men_n1358_));
  NO3        u1330(.A(men_men_n443_), .B(d), .C(c), .Y(men_men_n1359_));
  NO4        u1331(.A(men_men_n1358_), .B(men_men_n1356_), .C(men_men_n1354_), .D(men_men_n1348_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n144_), .B(h), .Y(men_men_n1361_));
  NO2        u1333(.A(men_men_n1064_), .B(l), .Y(men_men_n1362_));
  NO2        u1334(.A(g), .B(c), .Y(men_men_n1363_));
  NA3        u1335(.A(men_men_n1363_), .B(men_men_n139_), .C(men_men_n181_), .Y(men_men_n1364_));
  NO2        u1336(.A(men_men_n1364_), .B(men_men_n1362_), .Y(men_men_n1365_));
  NA2        u1337(.A(men_men_n1365_), .B(men_men_n176_), .Y(men_men_n1366_));
  NO2        u1338(.A(men_men_n451_), .B(a), .Y(men_men_n1367_));
  NA3        u1339(.A(men_men_n1367_), .B(k), .C(men_men_n113_), .Y(men_men_n1368_));
  NO2        u1340(.A(i), .B(h), .Y(men_men_n1369_));
  NA2        u1341(.A(men_men_n1124_), .B(h), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n135_), .B(men_men_n215_), .Y(men_men_n1371_));
  NO2        u1343(.A(men_men_n1371_), .B(men_men_n1370_), .Y(men_men_n1372_));
  NO2        u1344(.A(men_men_n758_), .B(men_men_n182_), .Y(men_men_n1373_));
  NOi31      u1345(.An(m), .B(n), .C(b), .Y(men_men_n1374_));
  NOi31      u1346(.An(f), .B(d), .C(c), .Y(men_men_n1375_));
  NA2        u1347(.A(men_men_n1375_), .B(men_men_n1374_), .Y(men_men_n1376_));
  INV        u1348(.A(men_men_n1376_), .Y(men_men_n1377_));
  NO3        u1349(.A(men_men_n1377_), .B(men_men_n1373_), .C(men_men_n1372_), .Y(men_men_n1378_));
  NA2        u1350(.A(men_men_n1074_), .B(men_men_n465_), .Y(men_men_n1379_));
  NO4        u1351(.A(men_men_n1379_), .B(men_men_n1052_), .C(men_men_n443_), .D(men_men_n43_), .Y(men_men_n1380_));
  OAI210     u1352(.A0(men_men_n179_), .A1(men_men_n521_), .B0(men_men_n1053_), .Y(men_men_n1381_));
  NO3        u1353(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1382_));
  INV        u1354(.A(men_men_n1381_), .Y(men_men_n1383_));
  NO2        u1355(.A(men_men_n1383_), .B(men_men_n1380_), .Y(men_men_n1384_));
  AN4        u1356(.A(men_men_n1384_), .B(men_men_n1378_), .C(men_men_n1368_), .D(men_men_n1366_), .Y(men_men_n1385_));
  NA2        u1357(.A(men_men_n1333_), .B(men_men_n378_), .Y(men_men_n1386_));
  NO2        u1358(.A(men_men_n1386_), .B(men_men_n1040_), .Y(men_men_n1387_));
  NA2        u1359(.A(men_men_n1359_), .B(men_men_n211_), .Y(men_men_n1388_));
  NO2        u1360(.A(men_men_n182_), .B(b), .Y(men_men_n1389_));
  AOI210     u1361(.A0(men_men_n1155_), .A1(men_men_n1389_), .B0(men_men_n1081_), .Y(men_men_n1390_));
  NO2        u1362(.A(i), .B(men_men_n209_), .Y(men_men_n1391_));
  NA4        u1363(.A(men_men_n1130_), .B(men_men_n1391_), .C(men_men_n105_), .D(m), .Y(men_men_n1392_));
  NAi41      u1364(.An(men_men_n1387_), .B(men_men_n1392_), .C(men_men_n1390_), .D(men_men_n1388_), .Y(men_men_n1393_));
  NO4        u1365(.A(men_men_n131_), .B(g), .C(f), .D(e), .Y(men_men_n1394_));
  NA3        u1366(.A(men_men_n1339_), .B(men_men_n287_), .C(h), .Y(men_men_n1395_));
  NOi41      u1367(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1396_));
  NA2        u1368(.A(men_men_n1396_), .B(men_men_n113_), .Y(men_men_n1397_));
  NA2        u1369(.A(men_men_n1336_), .B(men_men_n1357_), .Y(men_men_n1398_));
  NA2        u1370(.A(men_men_n1398_), .B(men_men_n1397_), .Y(men_men_n1399_));
  NA2        u1371(.A(men_men_n1102_), .B(men_men_n407_), .Y(men_men_n1400_));
  NO2        u1372(.A(men_men_n1400_), .B(men_men_n436_), .Y(men_men_n1401_));
  AO210      u1373(.A0(men_men_n1401_), .A1(men_men_n115_), .B0(men_men_n1399_), .Y(men_men_n1402_));
  NO2        u1374(.A(men_men_n1402_), .B(men_men_n1393_), .Y(men_men_n1403_));
  NA4        u1375(.A(men_men_n1403_), .B(men_men_n1385_), .C(men_men_n1360_), .D(men_men_n1344_), .Y(men_men_n1404_));
  NO2        u1376(.A(men_men_n390_), .B(j), .Y(men_men_n1405_));
  NA3        u1377(.A(men_men_n1382_), .B(men_men_n1330_), .C(men_men_n1102_), .Y(men_men_n1406_));
  NAi41      u1378(.An(men_men_n1369_), .B(men_men_n1062_), .C(men_men_n164_), .D(men_men_n146_), .Y(men_men_n1407_));
  NA2        u1379(.A(men_men_n1407_), .B(men_men_n1406_), .Y(men_men_n1408_));
  NA3        u1380(.A(g), .B(men_men_n1405_), .C(men_men_n153_), .Y(men_men_n1409_));
  INV        u1381(.A(men_men_n1409_), .Y(men_men_n1410_));
  NO3        u1382(.A(men_men_n753_), .B(men_men_n171_), .C(men_men_n410_), .Y(men_men_n1411_));
  NO3        u1383(.A(men_men_n1411_), .B(men_men_n1410_), .C(men_men_n1408_), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1504_), .B(men_men_n1047_), .Y(men_men_n1413_));
  OR2        u1385(.A(n), .B(i), .Y(men_men_n1414_));
  OAI210     u1386(.A0(men_men_n1414_), .A1(men_men_n1061_), .B0(men_men_n47_), .Y(men_men_n1415_));
  AOI220     u1387(.A0(men_men_n1415_), .A1(men_men_n1161_), .B0(men_men_n823_), .B1(men_men_n189_), .Y(men_men_n1416_));
  INV        u1388(.A(men_men_n1416_), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n219_), .B(k), .Y(men_men_n1418_));
  NO2        u1390(.A(men_men_n1417_), .B(men_men_n1413_), .Y(men_men_n1419_));
  INV        u1391(.A(men_men_n47_), .Y(men_men_n1420_));
  NO3        u1392(.A(men_men_n1083_), .B(men_men_n1330_), .C(men_men_n47_), .Y(men_men_n1421_));
  NA2        u1393(.A(men_men_n1084_), .B(men_men_n1420_), .Y(men_men_n1422_));
  NO2        u1394(.A(men_men_n1070_), .B(h), .Y(men_men_n1423_));
  NA2        u1395(.A(men_men_n1423_), .B(d), .Y(men_men_n1424_));
  OAI220     u1396(.A0(men_men_n1424_), .A1(c), .B0(men_men_n1422_), .B1(j), .Y(men_men_n1425_));
  AOI210     u1397(.A0(men_men_n521_), .A1(h), .B0(men_men_n67_), .Y(men_men_n1426_));
  NA2        u1398(.A(men_men_n1426_), .B(men_men_n1367_), .Y(men_men_n1427_));
  NO2        u1399(.A(men_men_n1322_), .B(men_men_n171_), .Y(men_men_n1428_));
  NOi21      u1400(.An(d), .B(f), .Y(men_men_n1429_));
  NO2        u1401(.A(men_men_n1375_), .B(men_men_n40_), .Y(men_men_n1430_));
  NA2        u1402(.A(men_men_n1430_), .B(men_men_n1428_), .Y(men_men_n1431_));
  NO2        u1403(.A(men_men_n1330_), .B(f), .Y(men_men_n1432_));
  NO2        u1404(.A(men_men_n296_), .B(c), .Y(men_men_n1433_));
  NA2        u1405(.A(men_men_n1433_), .B(men_men_n538_), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1434_), .B(men_men_n1431_), .C(men_men_n1427_), .Y(men_men_n1435_));
  NO2        u1407(.A(men_men_n1435_), .B(men_men_n1425_), .Y(men_men_n1436_));
  NA3        u1408(.A(men_men_n1436_), .B(men_men_n1419_), .C(men_men_n1412_), .Y(men_men_n1437_));
  NO3        u1409(.A(men_men_n1074_), .B(men_men_n1061_), .C(men_men_n40_), .Y(men_men_n1438_));
  NO2        u1410(.A(men_men_n465_), .B(men_men_n296_), .Y(men_men_n1439_));
  OAI210     u1411(.A0(men_men_n1439_), .A1(men_men_n1438_), .B0(men_men_n1340_), .Y(men_men_n1440_));
  OAI210     u1412(.A0(men_men_n1394_), .A1(men_men_n1333_), .B0(men_men_n881_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n1039_), .B(men_men_n131_), .Y(men_men_n1442_));
  NA2        u1414(.A(men_men_n1442_), .B(men_men_n624_), .Y(men_men_n1443_));
  NA3        u1415(.A(men_men_n1443_), .B(men_men_n1441_), .C(men_men_n1440_), .Y(men_men_n1444_));
  NA2        u1416(.A(men_men_n1363_), .B(men_men_n1429_), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n1445_), .B(m), .Y(men_men_n1446_));
  NO2        u1418(.A(men_men_n147_), .B(men_men_n178_), .Y(men_men_n1447_));
  OAI210     u1419(.A0(men_men_n1447_), .A1(men_men_n110_), .B0(men_men_n1374_), .Y(men_men_n1448_));
  INV        u1420(.A(men_men_n1448_), .Y(men_men_n1449_));
  NO3        u1421(.A(men_men_n1449_), .B(men_men_n1446_), .C(men_men_n1444_), .Y(men_men_n1450_));
  NO2        u1422(.A(men_men_n1329_), .B(e), .Y(men_men_n1451_));
  NA2        u1423(.A(men_men_n1451_), .B(men_men_n405_), .Y(men_men_n1452_));
  OAI210     u1424(.A0(men_men_n1432_), .A1(men_men_n1110_), .B0(men_men_n635_), .Y(men_men_n1453_));
  OR3        u1425(.A(men_men_n1418_), .B(men_men_n1196_), .C(men_men_n131_), .Y(men_men_n1454_));
  OAI220     u1426(.A0(men_men_n1454_), .A1(men_men_n1452_), .B0(men_men_n1453_), .B1(men_men_n445_), .Y(men_men_n1455_));
  INV        u1427(.A(men_men_n1455_), .Y(men_men_n1456_));
  NO2        u1428(.A(men_men_n178_), .B(c), .Y(men_men_n1457_));
  NA2        u1429(.A(men_men_n1457_), .B(men_men_n176_), .Y(men_men_n1458_));
  AOI220     u1430(.A0(men_men_n1458_), .A1(men_men_n1063_), .B0(men_men_n528_), .B1(men_men_n366_), .Y(men_men_n1459_));
  AOI210     u1431(.A0(j), .A1(men_men_n1359_), .B0(men_men_n1421_), .Y(men_men_n1460_));
  NA2        u1432(.A(men_men_n1110_), .B(a), .Y(men_men_n1461_));
  OAI220     u1433(.A0(men_men_n1461_), .A1(men_men_n67_), .B0(men_men_n1460_), .B1(men_men_n209_), .Y(men_men_n1462_));
  OR2        u1434(.A(h), .B(men_men_n536_), .Y(men_men_n1463_));
  NO2        u1435(.A(men_men_n1463_), .B(men_men_n171_), .Y(men_men_n1464_));
  NA3        u1436(.A(men_men_n1082_), .B(men_men_n215_), .C(men_men_n66_), .Y(men_men_n1465_));
  NA2        u1437(.A(men_men_n1334_), .B(men_men_n179_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n47_), .B(l), .Y(men_men_n1467_));
  INV        u1439(.A(men_men_n482_), .Y(men_men_n1468_));
  OAI210     u1440(.A0(men_men_n1468_), .A1(men_men_n1084_), .B0(men_men_n1467_), .Y(men_men_n1469_));
  NO2        u1441(.A(men_men_n245_), .B(g), .Y(men_men_n1470_));
  NO2        u1442(.A(m), .B(i), .Y(men_men_n1471_));
  BUFFER     u1443(.A(men_men_n1471_), .Y(men_men_n1472_));
  AOI220     u1444(.A0(men_men_n1472_), .A1(men_men_n1361_), .B0(men_men_n1062_), .B1(men_men_n1470_), .Y(men_men_n1473_));
  NA4        u1445(.A(men_men_n1473_), .B(men_men_n1469_), .C(men_men_n1466_), .D(men_men_n1465_), .Y(men_men_n1474_));
  NO4        u1446(.A(men_men_n1474_), .B(men_men_n1464_), .C(men_men_n1462_), .D(men_men_n1459_), .Y(men_men_n1475_));
  NA3        u1447(.A(men_men_n1475_), .B(men_men_n1456_), .C(men_men_n1450_), .Y(men_men_n1476_));
  NA3        u1448(.A(men_men_n959_), .B(men_men_n135_), .C(men_men_n44_), .Y(men_men_n1477_));
  AOI210     u1449(.A0(d), .A1(c), .B0(men_men_n1477_), .Y(men_men_n1478_));
  NO3        u1450(.A(men_men_n1349_), .B(men_men_n180_), .C(men_men_n450_), .Y(men_men_n1479_));
  NO2        u1451(.A(men_men_n1479_), .B(men_men_n1478_), .Y(men_men_n1480_));
  NO4        u1452(.A(men_men_n219_), .B(men_men_n180_), .C(men_men_n250_), .D(k), .Y(men_men_n1481_));
  NO2        u1453(.A(men_men_n1477_), .B(men_men_n110_), .Y(men_men_n1482_));
  NOi21      u1454(.An(men_men_n1334_), .B(e), .Y(men_men_n1483_));
  NO3        u1455(.A(men_men_n1483_), .B(men_men_n1482_), .C(men_men_n1481_), .Y(men_men_n1484_));
  NA2        u1456(.A(men_men_n1505_), .B(men_men_n154_), .Y(men_men_n1485_));
  NOi31      u1457(.An(men_men_n30_), .B(men_men_n1485_), .C(n), .Y(men_men_n1486_));
  INV        u1458(.A(men_men_n1486_), .Y(men_men_n1487_));
  NA2        u1459(.A(men_men_n57_), .B(a), .Y(men_men_n1488_));
  NO2        u1460(.A(men_men_n1339_), .B(men_men_n117_), .Y(men_men_n1489_));
  OAI220     u1461(.A0(men_men_n1489_), .A1(men_men_n1386_), .B0(men_men_n1400_), .B1(men_men_n1488_), .Y(men_men_n1490_));
  INV        u1462(.A(men_men_n1490_), .Y(men_men_n1491_));
  NA4        u1463(.A(men_men_n1491_), .B(men_men_n1487_), .C(men_men_n1484_), .D(men_men_n1480_), .Y(men_men_n1492_));
  OR4        u1464(.A(men_men_n1492_), .B(men_men_n1476_), .C(men_men_n1437_), .D(men_men_n1404_), .Y(men04));
  NOi31      u1465(.An(men_men_n1394_), .B(men_men_n1395_), .C(men_men_n1043_), .Y(men_men_n1494_));
  NA2        u1466(.A(men_men_n1432_), .B(men_men_n823_), .Y(men_men_n1495_));
  NO4        u1467(.A(men_men_n1495_), .B(men_men_n1034_), .C(men_men_n483_), .D(j), .Y(men_men_n1496_));
  OR3        u1468(.A(men_men_n1496_), .B(men_men_n1494_), .C(men_men_n1055_), .Y(men_men_n1497_));
  INV        u1469(.A(men_men_n1170_), .Y(men_men_n1498_));
  NA2        u1470(.A(men_men_n1498_), .B(men_men_n1200_), .Y(men_men_n1499_));
  NO3        u1471(.A(men_men_n1499_), .B(men_men_n1497_), .C(men_men_n1046_), .Y(men_men_n1500_));
  NA4        u1472(.A(men_men_n1500_), .B(men_men_n1112_), .C(men_men_n1100_), .D(men_men_n1087_), .Y(men05));
  INV        u1473(.A(men_men_n176_), .Y(men_men_n1504_));
  INV        u1474(.A(j), .Y(men_men_n1505_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule