library verilog;
use verilog.vl_types.all;
entity ex_mux_vlg_vec_tst is
end ex_mux_vlg_vec_tst;
