//Benchmark atmr_alu4_1266_0.0313

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n140_, ori_ori_n141_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1111_, men_men_n1112_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  OAI210     o033(.A0(ori_ori_n55_), .A1(ori_ori_n52_), .B0(ori_ori_n45_), .Y(ori_ori_n56_));
  NA3        o034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n57_));
  NO2        o035(.A(i_1_), .B(i_6_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_8_), .B(i_7_), .Y(ori_ori_n59_));
  OAI210     o037(.A0(ori_ori_n59_), .A1(ori_ori_n58_), .B0(ori_ori_n57_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n61_));
  NAi21      o039(.An(i_2_), .B(i_7_), .Y(ori_ori_n62_));
  INV        o040(.A(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NA3        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .C(ori_ori_n31_), .Y(ori_ori_n65_));
  NA2        o043(.A(i_1_), .B(i_10_), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n66_), .B(i_6_), .Y(ori_ori_n67_));
  NAi31      o045(.An(ori_ori_n67_), .B(ori_ori_n65_), .C(ori_ori_n61_), .Y(ori_ori_n68_));
  NA2        o046(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n69_));
  AOI210     o047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_1_), .B(i_6_), .Y(ori_ori_n71_));
  NO2        o049(.A(ori_ori_n71_), .B(ori_ori_n25_), .Y(ori_ori_n72_));
  INV        o050(.A(i_0_), .Y(ori_ori_n73_));
  NAi21      o051(.An(i_5_), .B(i_10_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_5_), .B(i_9_), .Y(ori_ori_n75_));
  AOI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n74_), .B0(ori_ori_n73_), .Y(ori_ori_n76_));
  NO2        o054(.A(ori_ori_n76_), .B(ori_ori_n72_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  OAI210     o056(.A0(ori_ori_n78_), .A1(ori_ori_n68_), .B0(i_0_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_12_), .B(i_5_), .Y(ori_ori_n80_));
  NA2        o058(.A(i_2_), .B(i_8_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n81_), .B(ori_ori_n58_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_9_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_3_), .B(i_7_), .Y(ori_ori_n84_));
  NO2        o062(.A(ori_ori_n83_), .B(ori_ori_n63_), .Y(ori_ori_n85_));
  INV        o063(.A(i_6_), .Y(ori_ori_n86_));
  NO2        o064(.A(i_2_), .B(i_7_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n87_), .Y(ori_ori_n88_));
  OAI210     o066(.A0(ori_ori_n85_), .A1(ori_ori_n82_), .B0(ori_ori_n88_), .Y(ori_ori_n89_));
  NAi21      o067(.An(i_6_), .B(i_10_), .Y(ori_ori_n90_));
  NA2        o068(.A(i_6_), .B(i_9_), .Y(ori_ori_n91_));
  AOI210     o069(.A0(ori_ori_n91_), .A1(ori_ori_n90_), .B0(ori_ori_n63_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_2_), .B(i_6_), .Y(ori_ori_n93_));
  NO3        o071(.A(ori_ori_n93_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n94_), .B(ori_ori_n92_), .Y(ori_ori_n95_));
  AOI210     o073(.A0(ori_ori_n95_), .A1(ori_ori_n89_), .B0(ori_ori_n80_), .Y(ori_ori_n96_));
  AN3        o074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n97_));
  NAi21      o075(.An(i_6_), .B(i_11_), .Y(ori_ori_n98_));
  NO2        o076(.A(i_5_), .B(i_8_), .Y(ori_ori_n99_));
  NOi21      o077(.An(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  AOI220     o078(.A0(ori_ori_n100_), .A1(ori_ori_n62_), .B0(ori_ori_n97_), .B1(ori_ori_n32_), .Y(ori_ori_n101_));
  INV        o079(.A(i_7_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n46_), .B(ori_ori_n102_), .Y(ori_ori_n103_));
  NO2        o081(.A(i_0_), .B(i_5_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(ori_ori_n86_), .Y(ori_ori_n105_));
  NA2        o083(.A(i_12_), .B(i_3_), .Y(ori_ori_n106_));
  INV        o084(.A(ori_ori_n106_), .Y(ori_ori_n107_));
  NA3        o085(.A(ori_ori_n107_), .B(ori_ori_n105_), .C(ori_ori_n103_), .Y(ori_ori_n108_));
  NAi21      o086(.An(i_7_), .B(i_11_), .Y(ori_ori_n109_));
  NO3        o087(.A(ori_ori_n109_), .B(ori_ori_n90_), .C(ori_ori_n53_), .Y(ori_ori_n110_));
  AN2        o088(.A(i_2_), .B(i_10_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(i_7_), .Y(ori_ori_n112_));
  OR2        o090(.A(ori_ori_n80_), .B(ori_ori_n58_), .Y(ori_ori_n113_));
  NO2        o091(.A(i_8_), .B(ori_ori_n102_), .Y(ori_ori_n114_));
  NO3        o092(.A(ori_ori_n114_), .B(ori_ori_n113_), .C(ori_ori_n112_), .Y(ori_ori_n115_));
  NA2        o093(.A(i_12_), .B(i_7_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n63_), .B(ori_ori_n26_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n117_), .B(i_0_), .Y(ori_ori_n118_));
  NA2        o096(.A(i_11_), .B(i_12_), .Y(ori_ori_n119_));
  OAI210     o097(.A0(ori_ori_n118_), .A1(ori_ori_n116_), .B0(ori_ori_n119_), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n120_), .B(ori_ori_n115_), .Y(ori_ori_n121_));
  NAi41      o099(.An(ori_ori_n110_), .B(ori_ori_n121_), .C(ori_ori_n108_), .D(ori_ori_n101_), .Y(ori_ori_n122_));
  NOi21      o100(.An(i_1_), .B(i_5_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(i_11_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n102_), .B(ori_ori_n37_), .Y(ori_ori_n125_));
  NA2        o103(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n126_), .B(ori_ori_n125_), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n127_), .B(ori_ori_n46_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n129_));
  NAi21      o107(.An(i_3_), .B(i_8_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(ori_ori_n62_), .Y(ori_ori_n131_));
  NOi31      o109(.An(ori_ori_n131_), .B(ori_ori_n129_), .C(ori_ori_n128_), .Y(ori_ori_n132_));
  NO2        o110(.A(i_1_), .B(ori_ori_n86_), .Y(ori_ori_n133_));
  NO2        o111(.A(i_6_), .B(i_5_), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n134_), .B(i_3_), .Y(ori_ori_n135_));
  AO210      o113(.A0(ori_ori_n135_), .A1(ori_ori_n47_), .B0(ori_ori_n133_), .Y(ori_ori_n136_));
  OAI220     o114(.A0(ori_ori_n136_), .A1(ori_ori_n109_), .B0(ori_ori_n132_), .B1(ori_ori_n124_), .Y(ori_ori_n137_));
  NO3        o115(.A(ori_ori_n137_), .B(ori_ori_n122_), .C(ori_ori_n96_), .Y(ori_ori_n138_));
  NA3        o116(.A(ori_ori_n138_), .B(ori_ori_n79_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o117(.A(ori_ori_n63_), .B(ori_ori_n37_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n772_), .B(ori_ori_n140_), .Y(ori_ori_n141_));
  NA4        o119(.A(ori_ori_n141_), .B(ori_ori_n77_), .C(ori_ori_n69_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o120(.A(i_8_), .B(i_7_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(i_6_), .Y(ori_ori_n144_));
  NO2        o122(.A(i_12_), .B(i_13_), .Y(ori_ori_n145_));
  NAi21      o123(.An(i_5_), .B(i_11_), .Y(ori_ori_n146_));
  NOi21      o124(.An(ori_ori_n145_), .B(ori_ori_n146_), .Y(ori_ori_n147_));
  NO2        o125(.A(i_0_), .B(i_1_), .Y(ori_ori_n148_));
  NA2        o126(.A(i_2_), .B(i_3_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n149_), .B(i_4_), .Y(ori_ori_n150_));
  AN2        o128(.A(ori_ori_n145_), .B(ori_ori_n83_), .Y(ori_ori_n151_));
  NA2        o129(.A(i_1_), .B(i_5_), .Y(ori_ori_n152_));
  OR2        o130(.A(i_0_), .B(i_1_), .Y(ori_ori_n153_));
  NO3        o131(.A(ori_ori_n153_), .B(ori_ori_n80_), .C(i_13_), .Y(ori_ori_n154_));
  NAi32      o132(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n155_));
  NAi21      o133(.An(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NOi21      o134(.An(i_4_), .B(i_10_), .Y(ori_ori_n157_));
  NA2        o135(.A(ori_ori_n157_), .B(ori_ori_n40_), .Y(ori_ori_n158_));
  NOi21      o136(.An(i_4_), .B(i_9_), .Y(ori_ori_n159_));
  NOi21      o137(.An(i_11_), .B(i_13_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NAi21      o139(.An(i_12_), .B(i_11_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n162_), .B(i_13_), .Y(ori_ori_n163_));
  NO2        o141(.A(ori_ori_n73_), .B(ori_ori_n63_), .Y(ori_ori_n164_));
  NO2        o142(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n165_));
  NO2        o143(.A(i_13_), .B(i_10_), .Y(ori_ori_n166_));
  NA3        o144(.A(ori_ori_n166_), .B(ori_ori_n165_), .C(ori_ori_n44_), .Y(ori_ori_n167_));
  NO2        o145(.A(i_2_), .B(i_1_), .Y(ori_ori_n168_));
  NAi21      o146(.An(i_4_), .B(i_12_), .Y(ori_ori_n169_));
  INV        o147(.A(i_8_), .Y(ori_ori_n170_));
  NO3        o148(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n171_));
  NO2        o149(.A(i_3_), .B(i_8_), .Y(ori_ori_n172_));
  NO3        o150(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n173_));
  NA3        o151(.A(ori_ori_n173_), .B(ori_ori_n172_), .C(ori_ori_n40_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n104_), .B(ori_ori_n58_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n153_), .Y(ori_ori_n176_));
  NO2        o154(.A(i_13_), .B(i_9_), .Y(ori_ori_n177_));
  NAi21      o155(.An(i_12_), .B(i_3_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n176_), .B(ori_ori_n174_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n180_), .B(i_7_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n181_), .B(i_4_), .Y(ori_ori_n182_));
  NAi21      o160(.An(i_12_), .B(i_7_), .Y(ori_ori_n183_));
  NA3        o161(.A(i_13_), .B(ori_ori_n170_), .C(i_10_), .Y(ori_ori_n184_));
  NA2        o162(.A(i_0_), .B(i_5_), .Y(ori_ori_n185_));
  NAi31      o163(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n73_), .B(ori_ori_n26_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n46_), .B(ori_ori_n63_), .Y(ori_ori_n189_));
  INV        o167(.A(i_13_), .Y(ori_ori_n190_));
  NO2        o168(.A(i_12_), .B(ori_ori_n190_), .Y(ori_ori_n191_));
  NO2        o169(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n192_));
  OR2        o170(.A(i_8_), .B(i_7_), .Y(ori_ori_n193_));
  INV        o171(.A(i_12_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n44_), .B(ori_ori_n194_), .Y(ori_ori_n195_));
  NO3        o173(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n196_));
  NA2        o174(.A(i_2_), .B(i_1_), .Y(ori_ori_n197_));
  NO3        o175(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n198_));
  NAi21      o176(.An(i_4_), .B(i_3_), .Y(ori_ori_n199_));
  NO2        o177(.A(i_0_), .B(i_6_), .Y(ori_ori_n200_));
  NOi41      o178(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n201_), .B(ori_ori_n200_), .Y(ori_ori_n202_));
  NO2        o180(.A(i_11_), .B(ori_ori_n190_), .Y(ori_ori_n203_));
  NOi21      o181(.An(i_1_), .B(i_6_), .Y(ori_ori_n204_));
  NAi21      o182(.An(i_3_), .B(i_7_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n194_), .B(i_9_), .Y(ori_ori_n206_));
  OR4        o184(.A(ori_ori_n206_), .B(ori_ori_n205_), .C(ori_ori_n204_), .D(ori_ori_n165_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n73_), .B(i_5_), .Y(ori_ori_n208_));
  NA2        o186(.A(i_3_), .B(i_9_), .Y(ori_ori_n209_));
  NAi21      o187(.An(i_7_), .B(i_10_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n210_), .B(ori_ori_n209_), .Y(ori_ori_n211_));
  NA3        o189(.A(ori_ori_n211_), .B(ori_ori_n208_), .C(ori_ori_n64_), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n212_), .B(ori_ori_n207_), .Y(ori_ori_n213_));
  INV        o191(.A(ori_ori_n144_), .Y(ori_ori_n214_));
  NA2        o192(.A(ori_ori_n194_), .B(i_13_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n215_), .B(ori_ori_n75_), .Y(ori_ori_n216_));
  AOI220     o194(.A0(ori_ori_n216_), .A1(ori_ori_n214_), .B0(ori_ori_n213_), .B1(ori_ori_n203_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n193_), .B(ori_ori_n37_), .Y(ori_ori_n218_));
  NA2        o196(.A(i_12_), .B(i_6_), .Y(ori_ori_n219_));
  OR2        o197(.A(i_13_), .B(i_9_), .Y(ori_ori_n220_));
  NO3        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .C(ori_ori_n48_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n199_), .B(i_2_), .Y(ori_ori_n222_));
  NA3        o200(.A(ori_ori_n222_), .B(ori_ori_n221_), .C(ori_ori_n44_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n203_), .B(i_9_), .Y(ori_ori_n224_));
  NA3        o202(.A(ori_ori_n208_), .B(ori_ori_n153_), .C(ori_ori_n64_), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n225_), .A1(ori_ori_n224_), .B0(ori_ori_n223_), .Y(ori_ori_n226_));
  NO3        o204(.A(i_11_), .B(ori_ori_n190_), .C(ori_ori_n25_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n205_), .B(i_8_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n226_), .B(ori_ori_n218_), .Y(ori_ori_n229_));
  NA2        o207(.A(ori_ori_n229_), .B(ori_ori_n217_), .Y(ori_ori_n230_));
  NO3        o208(.A(i_12_), .B(ori_ori_n190_), .C(ori_ori_n37_), .Y(ori_ori_n231_));
  NO2        o209(.A(i_2_), .B(ori_ori_n102_), .Y(ori_ori_n232_));
  AN2        o210(.A(i_3_), .B(i_10_), .Y(ori_ori_n233_));
  NO2        o211(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n234_));
  NO2        o212(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n230_), .B(ori_ori_n182_), .Y(ori_ori_n236_));
  NO3        o214(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n237_));
  NO2        o215(.A(i_2_), .B(i_3_), .Y(ori_ori_n238_));
  OR2        o216(.A(i_0_), .B(i_5_), .Y(ori_ori_n239_));
  NO2        o217(.A(i_12_), .B(i_10_), .Y(ori_ori_n240_));
  NOi21      o218(.An(i_5_), .B(i_0_), .Y(ori_ori_n241_));
  NA4        o219(.A(ori_ori_n84_), .B(ori_ori_n36_), .C(ori_ori_n86_), .D(i_8_), .Y(ori_ori_n242_));
  NO2        o220(.A(i_1_), .B(i_7_), .Y(ori_ori_n243_));
  NOi21      o221(.An(ori_ori_n152_), .B(ori_ori_n105_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(ori_ori_n126_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n245_), .B(i_3_), .Y(ori_ori_n246_));
  NO2        o224(.A(ori_ori_n170_), .B(i_9_), .Y(ori_ori_n247_));
  NA3        o225(.A(ori_ori_n247_), .B(ori_ori_n175_), .C(ori_ori_n153_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n248_), .B(ori_ori_n46_), .Y(ori_ori_n249_));
  INV        o227(.A(ori_ori_n249_), .Y(ori_ori_n250_));
  AOI210     o228(.A0(ori_ori_n250_), .A1(ori_ori_n246_), .B0(ori_ori_n158_), .Y(ori_ori_n251_));
  INV        o229(.A(ori_ori_n251_), .Y(ori_ori_n252_));
  NOi32      o230(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n253_));
  INV        o231(.A(ori_ori_n253_), .Y(ori_ori_n254_));
  NO2        o232(.A(ori_ori_n186_), .B(ori_ori_n155_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n155_), .B(ori_ori_n153_), .Y(ori_ori_n256_));
  NOi32      o234(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n257_));
  NAi21      o235(.An(i_6_), .B(i_1_), .Y(ori_ori_n258_));
  NA3        o236(.A(ori_ori_n258_), .B(ori_ori_n257_), .C(ori_ori_n46_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n259_), .B(i_0_), .Y(ori_ori_n260_));
  OR3        o238(.A(ori_ori_n260_), .B(ori_ori_n256_), .C(ori_ori_n255_), .Y(ori_ori_n261_));
  NO2        o239(.A(i_1_), .B(ori_ori_n102_), .Y(ori_ori_n262_));
  NAi21      o240(.An(i_3_), .B(i_4_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n263_), .B(i_9_), .Y(ori_ori_n264_));
  AN2        o242(.A(i_6_), .B(i_7_), .Y(ori_ori_n265_));
  OAI210     o243(.A0(ori_ori_n265_), .A1(ori_ori_n262_), .B0(ori_ori_n264_), .Y(ori_ori_n266_));
  NA2        o244(.A(i_2_), .B(i_7_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n263_), .B(i_10_), .Y(ori_ori_n268_));
  NA3        o246(.A(ori_ori_n268_), .B(ori_ori_n267_), .C(ori_ori_n200_), .Y(ori_ori_n269_));
  AOI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n266_), .B0(ori_ori_n165_), .Y(ori_ori_n270_));
  AOI210     o248(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n271_));
  OAI210     o249(.A0(ori_ori_n271_), .A1(ori_ori_n168_), .B0(ori_ori_n268_), .Y(ori_ori_n272_));
  AOI220     o250(.A0(ori_ori_n268_), .A1(ori_ori_n243_), .B0(ori_ori_n196_), .B1(ori_ori_n168_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n273_), .A1(ori_ori_n272_), .B0(i_5_), .Y(ori_ori_n274_));
  NO4        o252(.A(ori_ori_n274_), .B(ori_ori_n270_), .C(ori_ori_n261_), .D(ori_ori_n773_), .Y(ori_ori_n275_));
  NO2        o253(.A(ori_ori_n275_), .B(ori_ori_n254_), .Y(ori_ori_n276_));
  AN2        o254(.A(i_12_), .B(i_5_), .Y(ori_ori_n277_));
  NO2        o255(.A(i_11_), .B(i_6_), .Y(ori_ori_n278_));
  NO2        o256(.A(i_5_), .B(i_10_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n280_));
  NO3        o258(.A(ori_ori_n86_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n281_));
  NO2        o259(.A(i_11_), .B(i_12_), .Y(ori_ori_n282_));
  NAi21      o260(.An(i_13_), .B(i_0_), .Y(ori_ori_n283_));
  NO3        o261(.A(i_1_), .B(i_12_), .C(ori_ori_n86_), .Y(ori_ori_n284_));
  NO2        o262(.A(i_0_), .B(i_11_), .Y(ori_ori_n285_));
  AN2        o263(.A(i_1_), .B(i_6_), .Y(ori_ori_n286_));
  NOi21      o264(.An(i_2_), .B(i_12_), .Y(ori_ori_n287_));
  NAi21      o265(.An(i_9_), .B(i_4_), .Y(ori_ori_n288_));
  OR2        o266(.A(i_13_), .B(i_10_), .Y(ori_ori_n289_));
  NO3        o267(.A(ori_ori_n289_), .B(ori_ori_n119_), .C(ori_ori_n288_), .Y(ori_ori_n290_));
  NO2        o268(.A(ori_ori_n161_), .B(ori_ori_n125_), .Y(ori_ori_n291_));
  NO2        o269(.A(ori_ori_n102_), .B(ori_ori_n25_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n231_), .B(ori_ori_n292_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n293_), .B(ori_ori_n244_), .Y(ori_ori_n294_));
  INV        o272(.A(ori_ori_n294_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n295_), .B(ori_ori_n26_), .Y(ori_ori_n296_));
  NA2        o274(.A(ori_ori_n170_), .B(i_10_), .Y(ori_ori_n297_));
  NA3        o275(.A(ori_ori_n208_), .B(ori_ori_n64_), .C(i_2_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(ori_ori_n297_), .Y(ori_ori_n299_));
  INV        o277(.A(ori_ori_n299_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n300_), .B(ori_ori_n224_), .Y(ori_ori_n301_));
  NO3        o279(.A(ori_ori_n301_), .B(ori_ori_n296_), .C(ori_ori_n276_), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n73_), .B(i_13_), .Y(ori_ori_n303_));
  NO2        o281(.A(i_10_), .B(i_9_), .Y(ori_ori_n304_));
  NAi21      o282(.An(i_12_), .B(i_8_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n305_), .B(i_3_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n235_), .B(i_0_), .Y(ori_ori_n307_));
  NO3        o285(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n219_), .B(ori_ori_n98_), .Y(ori_ori_n309_));
  NA2        o287(.A(ori_ori_n309_), .B(ori_ori_n308_), .Y(ori_ori_n310_));
  NA2        o288(.A(i_8_), .B(i_9_), .Y(ori_ori_n311_));
  AOI210     o289(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n312_));
  OR2        o290(.A(ori_ori_n312_), .B(ori_ori_n311_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n231_), .B(ori_ori_n175_), .Y(ori_ori_n314_));
  OAI220     o292(.A0(ori_ori_n314_), .A1(ori_ori_n313_), .B0(ori_ori_n310_), .B1(ori_ori_n307_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n203_), .B(ori_ori_n234_), .Y(ori_ori_n316_));
  NO3        o294(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n317_));
  INV        o295(.A(ori_ori_n317_), .Y(ori_ori_n318_));
  NA3        o296(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n319_));
  NA4        o297(.A(ori_ori_n146_), .B(ori_ori_n117_), .C(ori_ori_n80_), .D(ori_ori_n23_), .Y(ori_ori_n320_));
  OAI220     o298(.A0(ori_ori_n320_), .A1(ori_ori_n319_), .B0(ori_ori_n318_), .B1(ori_ori_n316_), .Y(ori_ori_n321_));
  NO2        o299(.A(ori_ori_n321_), .B(ori_ori_n315_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n97_), .B(i_13_), .Y(ori_ori_n323_));
  NO2        o301(.A(i_2_), .B(i_13_), .Y(ori_ori_n324_));
  NO3        o302(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n325_));
  NO2        o303(.A(i_6_), .B(i_7_), .Y(ori_ori_n326_));
  NO2        o304(.A(i_11_), .B(i_1_), .Y(ori_ori_n327_));
  NOi21      o305(.An(i_2_), .B(i_7_), .Y(ori_ori_n328_));
  NO2        o306(.A(i_3_), .B(ori_ori_n170_), .Y(ori_ori_n329_));
  NO2        o307(.A(i_6_), .B(i_10_), .Y(ori_ori_n330_));
  NA3        o308(.A(ori_ori_n201_), .B(ori_ori_n160_), .C(ori_ori_n134_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n153_), .B(i_3_), .Y(ori_ori_n333_));
  NAi31      o311(.An(ori_ori_n332_), .B(ori_ori_n333_), .C(ori_ori_n191_), .Y(ori_ori_n334_));
  NA3        o312(.A(ori_ori_n280_), .B(ori_ori_n164_), .C(ori_ori_n150_), .Y(ori_ori_n335_));
  NA3        o313(.A(ori_ori_n335_), .B(ori_ori_n334_), .C(ori_ori_n331_), .Y(ori_ori_n336_));
  INV        o314(.A(ori_ori_n336_), .Y(ori_ori_n337_));
  NA2        o315(.A(ori_ori_n308_), .B(ori_ori_n277_), .Y(ori_ori_n338_));
  NA2        o316(.A(ori_ori_n317_), .B(ori_ori_n279_), .Y(ori_ori_n339_));
  NAi21      o317(.An(ori_ori_n184_), .B(ori_ori_n282_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n243_), .B(ori_ori_n185_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n340_), .Y(ori_ori_n342_));
  NA2        o320(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n237_), .B(ori_ori_n196_), .Y(ori_ori_n344_));
  OAI220     o322(.A0(ori_ori_n344_), .A1(ori_ori_n298_), .B0(ori_ori_n343_), .B1(ori_ori_n323_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n345_), .B(ori_ori_n342_), .Y(ori_ori_n346_));
  NA3        o324(.A(ori_ori_n346_), .B(ori_ori_n337_), .C(ori_ori_n322_), .Y(ori_ori_n347_));
  NA2        o325(.A(ori_ori_n277_), .B(ori_ori_n190_), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n265_), .B(ori_ori_n257_), .Y(ori_ori_n349_));
  OR2        o327(.A(ori_ori_n348_), .B(ori_ori_n349_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n351_));
  AOI210     o329(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n290_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n352_), .B(ori_ori_n350_), .Y(ori_ori_n353_));
  INV        o331(.A(ori_ori_n353_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n208_), .B(ori_ori_n64_), .Y(ori_ori_n355_));
  OAI210     o333(.A0(i_8_), .A1(ori_ori_n355_), .B0(ori_ori_n136_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(ori_ori_n291_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n357_), .B(ori_ori_n354_), .Y(ori_ori_n358_));
  NO2        o336(.A(i_12_), .B(ori_ori_n170_), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n360_));
  NO2        o338(.A(ori_ori_n360_), .B(i_6_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n153_), .B(i_5_), .Y(ori_ori_n362_));
  NA3        o340(.A(ori_ori_n185_), .B(ori_ori_n71_), .C(ori_ori_n44_), .Y(ori_ori_n363_));
  NA2        o341(.A(ori_ori_n231_), .B(ori_ori_n84_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n363_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  NA2        o343(.A(ori_ori_n189_), .B(ori_ori_n188_), .Y(ori_ori_n366_));
  NA2        o344(.A(ori_ori_n304_), .B(ori_ori_n187_), .Y(ori_ori_n367_));
  NO2        o345(.A(ori_ori_n366_), .B(ori_ori_n367_), .Y(ori_ori_n368_));
  AOI210     o346(.A0(ori_ori_n258_), .A1(ori_ori_n46_), .B0(ori_ori_n262_), .Y(ori_ori_n369_));
  NA2        o347(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n370_));
  NA3        o348(.A(ori_ori_n359_), .B(ori_ori_n227_), .C(ori_ori_n370_), .Y(ori_ori_n371_));
  NO2        o349(.A(ori_ori_n369_), .B(ori_ori_n371_), .Y(ori_ori_n372_));
  NO3        o350(.A(ori_ori_n372_), .B(ori_ori_n368_), .C(ori_ori_n365_), .Y(ori_ori_n373_));
  NO4        o351(.A(ori_ori_n204_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n374_));
  NO3        o352(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n289_), .B(i_1_), .Y(ori_ori_n376_));
  NOi31      o354(.An(ori_ori_n376_), .B(ori_ori_n309_), .C(ori_ori_n73_), .Y(ori_ori_n377_));
  NOi21      o355(.An(i_10_), .B(i_6_), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n379_));
  AOI220     o357(.A0(ori_ori_n231_), .A1(ori_ori_n379_), .B0(ori_ori_n227_), .B1(ori_ori_n378_), .Y(ori_ori_n380_));
  NO2        o358(.A(ori_ori_n380_), .B(ori_ori_n307_), .Y(ori_ori_n381_));
  NO2        o359(.A(ori_ori_n116_), .B(ori_ori_n23_), .Y(ori_ori_n382_));
  NOi31      o360(.An(ori_ori_n147_), .B(i_10_), .C(ori_ori_n242_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n383_), .B(ori_ori_n381_), .Y(ori_ori_n384_));
  INV        o362(.A(ori_ori_n238_), .Y(ori_ori_n385_));
  NO2        o363(.A(i_12_), .B(ori_ori_n86_), .Y(ori_ori_n386_));
  NA3        o364(.A(ori_ori_n386_), .B(ori_ori_n227_), .C(ori_ori_n370_), .Y(ori_ori_n387_));
  NA3        o365(.A(ori_ori_n278_), .B(ori_ori_n231_), .C(ori_ori_n185_), .Y(ori_ori_n388_));
  AOI210     o366(.A0(ori_ori_n388_), .A1(ori_ori_n387_), .B0(ori_ori_n385_), .Y(ori_ori_n389_));
  OR2        o367(.A(i_2_), .B(i_5_), .Y(ori_ori_n390_));
  OR2        o368(.A(ori_ori_n390_), .B(ori_ori_n286_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n267_), .B(ori_ori_n200_), .Y(ori_ori_n392_));
  AOI210     o370(.A0(ori_ori_n392_), .A1(ori_ori_n391_), .B0(ori_ori_n340_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n393_), .B(ori_ori_n389_), .Y(ori_ori_n394_));
  NA3        o372(.A(ori_ori_n394_), .B(ori_ori_n384_), .C(ori_ori_n373_), .Y(ori_ori_n395_));
  NO3        o373(.A(ori_ori_n395_), .B(ori_ori_n358_), .C(ori_ori_n347_), .Y(ori_ori_n396_));
  NA4        o374(.A(ori_ori_n396_), .B(ori_ori_n302_), .C(ori_ori_n252_), .D(ori_ori_n236_), .Y(ori7));
  NO2        o375(.A(ori_ori_n93_), .B(ori_ori_n54_), .Y(ori_ori_n398_));
  NA2        o376(.A(ori_ori_n330_), .B(ori_ori_n84_), .Y(ori_ori_n399_));
  NA2        o377(.A(i_11_), .B(ori_ori_n170_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n145_), .B(ori_ori_n400_), .Y(ori_ori_n401_));
  NO2        o379(.A(ori_ori_n401_), .B(ori_ori_n399_), .Y(ori_ori_n402_));
  NA3        o380(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n403_));
  NO2        o381(.A(ori_ori_n194_), .B(i_4_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n404_), .B(i_8_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n106_), .B(ori_ori_n403_), .Y(ori_ori_n406_));
  NA2        o384(.A(i_2_), .B(ori_ori_n86_), .Y(ori_ori_n407_));
  OAI210     o385(.A0(ori_ori_n87_), .A1(ori_ori_n172_), .B0(ori_ori_n173_), .Y(ori_ori_n408_));
  NO2        o386(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n409_));
  NA2        o387(.A(i_4_), .B(i_8_), .Y(ori_ori_n410_));
  AOI210     o388(.A0(ori_ori_n410_), .A1(ori_ori_n233_), .B0(ori_ori_n409_), .Y(ori_ori_n411_));
  OAI220     o389(.A0(ori_ori_n411_), .A1(ori_ori_n407_), .B0(ori_ori_n408_), .B1(i_13_), .Y(ori_ori_n412_));
  NO4        o390(.A(ori_ori_n412_), .B(ori_ori_n406_), .C(ori_ori_n402_), .D(ori_ori_n398_), .Y(ori_ori_n413_));
  AOI210     o391(.A0(ori_ori_n130_), .A1(ori_ori_n62_), .B0(i_10_), .Y(ori_ori_n414_));
  AOI210     o392(.A0(ori_ori_n414_), .A1(ori_ori_n194_), .B0(ori_ori_n157_), .Y(ori_ori_n415_));
  OR2        o393(.A(i_6_), .B(i_10_), .Y(ori_ori_n416_));
  NO2        o394(.A(ori_ori_n416_), .B(ori_ori_n23_), .Y(ori_ori_n417_));
  OR3        o395(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n418_));
  INV        o396(.A(ori_ori_n171_), .Y(ori_ori_n419_));
  INV        o397(.A(ori_ori_n417_), .Y(ori_ori_n420_));
  OA220      o398(.A0(ori_ori_n420_), .A1(ori_ori_n385_), .B0(ori_ori_n415_), .B1(ori_ori_n220_), .Y(ori_ori_n421_));
  AOI210     o399(.A0(ori_ori_n421_), .A1(ori_ori_n413_), .B0(ori_ori_n63_), .Y(ori_ori_n422_));
  NOi21      o400(.An(i_11_), .B(i_7_), .Y(ori_ori_n423_));
  AO210      o401(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n424_));
  NO2        o402(.A(ori_ori_n424_), .B(ori_ori_n423_), .Y(ori_ori_n425_));
  NA2        o403(.A(ori_ori_n425_), .B(ori_ori_n177_), .Y(ori_ori_n426_));
  NA3        o404(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n427_));
  NO2        o405(.A(ori_ori_n426_), .B(ori_ori_n63_), .Y(ori_ori_n428_));
  OR2        o406(.A(ori_ori_n273_), .B(ori_ori_n41_), .Y(ori_ori_n429_));
  NO3        o407(.A(ori_ori_n210_), .B(ori_ori_n178_), .C(ori_ori_n400_), .Y(ori_ori_n430_));
  OAI210     o408(.A0(ori_ori_n430_), .A1(ori_ori_n191_), .B0(ori_ori_n63_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n287_), .B(ori_ori_n31_), .Y(ori_ori_n432_));
  OR2        o410(.A(ori_ori_n178_), .B(ori_ori_n109_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n433_), .B(ori_ori_n432_), .Y(ori_ori_n434_));
  NO2        o412(.A(i_1_), .B(i_4_), .Y(ori_ori_n435_));
  NA2        o413(.A(ori_ori_n435_), .B(ori_ori_n434_), .Y(ori_ori_n436_));
  NO2        o414(.A(i_1_), .B(i_12_), .Y(ori_ori_n437_));
  NA3        o415(.A(ori_ori_n437_), .B(ori_ori_n111_), .C(ori_ori_n24_), .Y(ori_ori_n438_));
  BUFFER     o416(.A(ori_ori_n438_), .Y(ori_ori_n439_));
  NA4        o417(.A(ori_ori_n439_), .B(ori_ori_n436_), .C(ori_ori_n431_), .D(ori_ori_n429_), .Y(ori_ori_n440_));
  OAI210     o418(.A0(ori_ori_n440_), .A1(ori_ori_n428_), .B0(i_6_), .Y(ori_ori_n441_));
  NO2        o419(.A(ori_ori_n427_), .B(ori_ori_n109_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n442_), .B(ori_ori_n386_), .Y(ori_ori_n443_));
  NO2        o421(.A(i_6_), .B(i_11_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n443_), .B(ori_ori_n310_), .Y(ori_ori_n445_));
  NO3        o423(.A(ori_ori_n416_), .B(ori_ori_n193_), .C(ori_ori_n23_), .Y(ori_ori_n446_));
  AOI210     o424(.A0(i_1_), .A1(ori_ori_n211_), .B0(ori_ori_n446_), .Y(ori_ori_n447_));
  NO2        o425(.A(ori_ori_n447_), .B(ori_ori_n44_), .Y(ori_ori_n448_));
  INV        o426(.A(i_2_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n140_), .B(i_9_), .Y(ori_ori_n450_));
  NA3        o428(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n451_));
  NO2        o429(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n452_));
  NA3        o430(.A(ori_ori_n452_), .B(ori_ori_n219_), .C(ori_ori_n44_), .Y(ori_ori_n453_));
  OAI220     o431(.A0(ori_ori_n453_), .A1(ori_ori_n451_), .B0(ori_ori_n450_), .B1(ori_ori_n449_), .Y(ori_ori_n454_));
  AOI210     o432(.A0(ori_ori_n327_), .A1(ori_ori_n292_), .B0(ori_ori_n198_), .Y(ori_ori_n455_));
  NO2        o433(.A(ori_ori_n455_), .B(ori_ori_n407_), .Y(ori_ori_n456_));
  NO2        o434(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n457_));
  OR2        o435(.A(ori_ori_n456_), .B(ori_ori_n454_), .Y(ori_ori_n458_));
  NO3        o436(.A(ori_ori_n458_), .B(ori_ori_n448_), .C(ori_ori_n445_), .Y(ori_ori_n459_));
  NO2        o437(.A(ori_ori_n194_), .B(ori_ori_n102_), .Y(ori_ori_n460_));
  NO2        o438(.A(ori_ori_n460_), .B(ori_ori_n423_), .Y(ori_ori_n461_));
  NA2        o439(.A(ori_ori_n461_), .B(i_1_), .Y(ori_ori_n462_));
  NO2        o440(.A(ori_ori_n462_), .B(ori_ori_n418_), .Y(ori_ori_n463_));
  NO2        o441(.A(ori_ori_n288_), .B(ori_ori_n86_), .Y(ori_ori_n464_));
  NA2        o442(.A(ori_ori_n463_), .B(ori_ori_n46_), .Y(ori_ori_n465_));
  NA2        o443(.A(i_3_), .B(ori_ori_n170_), .Y(ori_ori_n466_));
  NO2        o444(.A(ori_ori_n466_), .B(ori_ori_n116_), .Y(ori_ori_n467_));
  AN2        o445(.A(ori_ori_n467_), .B(ori_ori_n361_), .Y(ori_ori_n468_));
  NO2        o446(.A(ori_ori_n193_), .B(ori_ori_n44_), .Y(ori_ori_n469_));
  NO3        o447(.A(ori_ori_n469_), .B(ori_ori_n235_), .C(ori_ori_n195_), .Y(ori_ori_n470_));
  NO2        o448(.A(ori_ori_n119_), .B(ori_ori_n37_), .Y(ori_ori_n471_));
  NO2        o449(.A(ori_ori_n471_), .B(i_6_), .Y(ori_ori_n472_));
  NO2        o450(.A(ori_ori_n86_), .B(i_9_), .Y(ori_ori_n473_));
  NO2        o451(.A(ori_ori_n473_), .B(ori_ori_n63_), .Y(ori_ori_n474_));
  NO2        o452(.A(ori_ori_n474_), .B(ori_ori_n437_), .Y(ori_ori_n475_));
  NO4        o453(.A(ori_ori_n475_), .B(ori_ori_n472_), .C(ori_ori_n470_), .D(i_4_), .Y(ori_ori_n476_));
  NA2        o454(.A(i_1_), .B(i_3_), .Y(ori_ori_n477_));
  NO2        o455(.A(ori_ori_n311_), .B(ori_ori_n93_), .Y(ori_ori_n478_));
  AOI210     o456(.A0(ori_ori_n469_), .A1(ori_ori_n378_), .B0(ori_ori_n478_), .Y(ori_ori_n479_));
  NO2        o457(.A(ori_ori_n479_), .B(ori_ori_n477_), .Y(ori_ori_n480_));
  NO3        o458(.A(ori_ori_n480_), .B(ori_ori_n476_), .C(ori_ori_n468_), .Y(ori_ori_n481_));
  NA4        o459(.A(ori_ori_n481_), .B(ori_ori_n465_), .C(ori_ori_n459_), .D(ori_ori_n441_), .Y(ori_ori_n482_));
  AN2        o460(.A(ori_ori_n201_), .B(ori_ori_n86_), .Y(ori_ori_n483_));
  NA2        o461(.A(ori_ori_n265_), .B(ori_ori_n264_), .Y(ori_ori_n484_));
  NO3        o462(.A(ori_ori_n328_), .B(ori_ori_n410_), .C(ori_ori_n86_), .Y(ori_ori_n485_));
  NA2        o463(.A(ori_ori_n485_), .B(ori_ori_n25_), .Y(ori_ori_n486_));
  NA2        o464(.A(ori_ori_n486_), .B(ori_ori_n484_), .Y(ori_ori_n487_));
  OAI210     o465(.A0(ori_ori_n487_), .A1(ori_ori_n483_), .B0(i_1_), .Y(ori_ori_n488_));
  AOI210     o466(.A0(ori_ori_n219_), .A1(ori_ori_n98_), .B0(i_1_), .Y(ori_ori_n489_));
  NO2        o467(.A(ori_ori_n263_), .B(i_2_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n490_), .B(ori_ori_n489_), .Y(ori_ori_n491_));
  AOI210     o469(.A0(ori_ori_n491_), .A1(ori_ori_n488_), .B0(i_13_), .Y(ori_ori_n492_));
  OR2        o470(.A(i_11_), .B(i_7_), .Y(ori_ori_n493_));
  NO2        o471(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n494_));
  NO2        o472(.A(ori_ori_n328_), .B(ori_ori_n24_), .Y(ori_ori_n495_));
  AOI220     o473(.A0(ori_ori_n495_), .A1(ori_ori_n464_), .B0(ori_ori_n201_), .B1(ori_ori_n133_), .Y(ori_ori_n496_));
  OAI220     o474(.A0(ori_ori_n496_), .A1(ori_ori_n41_), .B0(ori_ori_n771_), .B1(ori_ori_n93_), .Y(ori_ori_n497_));
  INV        o475(.A(ori_ori_n497_), .Y(ori_ori_n498_));
  INV        o476(.A(ori_ori_n116_), .Y(ori_ori_n499_));
  AOI220     o477(.A0(ori_ori_n499_), .A1(ori_ori_n72_), .B0(ori_ori_n278_), .B1(ori_ori_n452_), .Y(ori_ori_n500_));
  NO2        o478(.A(ori_ori_n500_), .B(ori_ori_n199_), .Y(ori_ori_n501_));
  AOI210     o479(.A0(ori_ori_n305_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n502_));
  NOi31      o480(.An(ori_ori_n502_), .B(ori_ori_n399_), .C(ori_ori_n44_), .Y(ori_ori_n503_));
  NA2        o481(.A(ori_ori_n129_), .B(i_13_), .Y(ori_ori_n504_));
  NO2        o482(.A(ori_ori_n451_), .B(ori_ori_n116_), .Y(ori_ori_n505_));
  INV        o483(.A(ori_ori_n505_), .Y(ori_ori_n506_));
  OAI220     o484(.A0(ori_ori_n506_), .A1(ori_ori_n71_), .B0(ori_ori_n504_), .B1(ori_ori_n489_), .Y(ori_ori_n507_));
  NO3        o485(.A(ori_ori_n71_), .B(ori_ori_n32_), .C(ori_ori_n102_), .Y(ori_ori_n508_));
  NA2        o486(.A(ori_ori_n26_), .B(ori_ori_n170_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n509_), .B(i_7_), .Y(ori_ori_n510_));
  NO3        o488(.A(ori_ori_n328_), .B(ori_ori_n194_), .C(ori_ori_n86_), .Y(ori_ori_n511_));
  AOI210     o489(.A0(ori_ori_n511_), .A1(ori_ori_n510_), .B0(ori_ori_n508_), .Y(ori_ori_n512_));
  AOI220     o490(.A0(ori_ori_n278_), .A1(ori_ori_n452_), .B0(ori_ori_n92_), .B1(ori_ori_n103_), .Y(ori_ori_n513_));
  OAI220     o491(.A0(ori_ori_n513_), .A1(ori_ori_n405_), .B0(ori_ori_n512_), .B1(ori_ori_n419_), .Y(ori_ori_n514_));
  NO4        o492(.A(ori_ori_n514_), .B(ori_ori_n507_), .C(ori_ori_n503_), .D(ori_ori_n501_), .Y(ori_ori_n515_));
  OR2        o493(.A(i_11_), .B(i_6_), .Y(ori_ori_n516_));
  NA3        o494(.A(ori_ori_n404_), .B(ori_ori_n509_), .C(i_7_), .Y(ori_ori_n517_));
  AOI210     o495(.A0(ori_ori_n517_), .A1(ori_ori_n506_), .B0(ori_ori_n516_), .Y(ori_ori_n518_));
  NA3        o496(.A(ori_ori_n287_), .B(ori_ori_n409_), .C(ori_ori_n98_), .Y(ori_ori_n519_));
  NA2        o497(.A(ori_ori_n444_), .B(i_13_), .Y(ori_ori_n520_));
  NA2        o498(.A(ori_ori_n103_), .B(ori_ori_n509_), .Y(ori_ori_n521_));
  NAi21      o499(.An(i_11_), .B(i_12_), .Y(ori_ori_n522_));
  NOi41      o500(.An(ori_ori_n112_), .B(ori_ori_n522_), .C(i_13_), .D(ori_ori_n86_), .Y(ori_ori_n523_));
  NO3        o501(.A(ori_ori_n328_), .B(ori_ori_n386_), .C(ori_ori_n410_), .Y(ori_ori_n524_));
  AOI220     o502(.A0(ori_ori_n524_), .A1(ori_ori_n237_), .B0(ori_ori_n523_), .B1(ori_ori_n521_), .Y(ori_ori_n525_));
  NA3        o503(.A(ori_ori_n525_), .B(ori_ori_n520_), .C(ori_ori_n519_), .Y(ori_ori_n526_));
  OAI210     o504(.A0(ori_ori_n526_), .A1(ori_ori_n518_), .B0(ori_ori_n63_), .Y(ori_ori_n527_));
  NO2        o505(.A(i_2_), .B(i_12_), .Y(ori_ori_n528_));
  NA2        o506(.A(ori_ori_n262_), .B(ori_ori_n528_), .Y(ori_ori_n529_));
  NA2        o507(.A(ori_ori_n264_), .B(ori_ori_n262_), .Y(ori_ori_n530_));
  NO2        o508(.A(ori_ori_n130_), .B(i_2_), .Y(ori_ori_n531_));
  NA2        o509(.A(ori_ori_n531_), .B(ori_ori_n437_), .Y(ori_ori_n532_));
  NA3        o510(.A(ori_ori_n532_), .B(ori_ori_n530_), .C(ori_ori_n529_), .Y(ori_ori_n533_));
  NA3        o511(.A(ori_ori_n533_), .B(ori_ori_n45_), .C(ori_ori_n190_), .Y(ori_ori_n534_));
  NA4        o512(.A(ori_ori_n534_), .B(ori_ori_n527_), .C(ori_ori_n515_), .D(ori_ori_n498_), .Y(ori_ori_n535_));
  OR4        o513(.A(ori_ori_n535_), .B(ori_ori_n492_), .C(ori_ori_n482_), .D(ori_ori_n422_), .Y(ori5));
  NA2        o514(.A(ori_ori_n461_), .B(ori_ori_n222_), .Y(ori_ori_n537_));
  AN2        o515(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n538_));
  NA3        o516(.A(ori_ori_n538_), .B(ori_ori_n528_), .C(ori_ori_n109_), .Y(ori_ori_n539_));
  NO2        o517(.A(ori_ori_n405_), .B(i_11_), .Y(ori_ori_n540_));
  NA2        o518(.A(ori_ori_n87_), .B(ori_ori_n540_), .Y(ori_ori_n541_));
  NA3        o519(.A(ori_ori_n541_), .B(ori_ori_n539_), .C(ori_ori_n537_), .Y(ori_ori_n542_));
  NO3        o520(.A(i_11_), .B(ori_ori_n194_), .C(i_13_), .Y(ori_ori_n543_));
  NO2        o521(.A(ori_ori_n126_), .B(ori_ori_n23_), .Y(ori_ori_n544_));
  NA2        o522(.A(i_12_), .B(i_8_), .Y(ori_ori_n545_));
  OAI210     o523(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n545_), .Y(ori_ori_n546_));
  INV        o524(.A(ori_ori_n304_), .Y(ori_ori_n547_));
  AOI220     o525(.A0(ori_ori_n238_), .A1(ori_ori_n382_), .B0(ori_ori_n546_), .B1(ori_ori_n544_), .Y(ori_ori_n548_));
  INV        o526(.A(ori_ori_n548_), .Y(ori_ori_n549_));
  NO2        o527(.A(ori_ori_n549_), .B(ori_ori_n542_), .Y(ori_ori_n550_));
  INV        o528(.A(ori_ori_n160_), .Y(ori_ori_n551_));
  INV        o529(.A(ori_ori_n201_), .Y(ori_ori_n552_));
  OAI210     o530(.A0(ori_ori_n490_), .A1(ori_ori_n306_), .B0(ori_ori_n112_), .Y(ori_ori_n553_));
  AOI210     o531(.A0(ori_ori_n553_), .A1(ori_ori_n552_), .B0(ori_ori_n551_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n311_), .B(ori_ori_n26_), .Y(ori_ori_n555_));
  NO2        o533(.A(ori_ori_n555_), .B(ori_ori_n292_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n556_), .B(i_2_), .Y(ori_ori_n557_));
  INV        o535(.A(ori_ori_n557_), .Y(ori_ori_n558_));
  AOI210     o536(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n289_), .Y(ori_ori_n559_));
  AOI210     o537(.A0(ori_ori_n559_), .A1(ori_ori_n558_), .B0(ori_ori_n554_), .Y(ori_ori_n560_));
  NO2        o538(.A(ori_ori_n169_), .B(ori_ori_n127_), .Y(ori_ori_n561_));
  OAI210     o539(.A0(ori_ori_n561_), .A1(ori_ori_n544_), .B0(i_2_), .Y(ori_ori_n562_));
  INV        o540(.A(ori_ori_n161_), .Y(ori_ori_n563_));
  NO3        o541(.A(ori_ori_n424_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n564_));
  AOI210     o542(.A0(ori_ori_n563_), .A1(ori_ori_n87_), .B0(ori_ori_n564_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n565_), .A1(ori_ori_n562_), .B0(ori_ori_n170_), .Y(ori_ori_n566_));
  OA210      o544(.A0(ori_ori_n425_), .A1(ori_ori_n128_), .B0(i_13_), .Y(ori_ori_n567_));
  NA2        o545(.A(ori_ori_n171_), .B(ori_ori_n172_), .Y(ori_ori_n568_));
  NA2        o546(.A(ori_ori_n151_), .B(ori_ori_n400_), .Y(ori_ori_n569_));
  AOI210     o547(.A0(ori_ori_n569_), .A1(ori_ori_n568_), .B0(ori_ori_n267_), .Y(ori_ori_n570_));
  AOI210     o548(.A0(ori_ori_n178_), .A1(ori_ori_n149_), .B0(ori_ori_n351_), .Y(ori_ori_n571_));
  OAI210     o549(.A0(ori_ori_n571_), .A1(ori_ori_n191_), .B0(ori_ori_n292_), .Y(ori_ori_n572_));
  NO2        o550(.A(ori_ori_n103_), .B(ori_ori_n44_), .Y(ori_ori_n573_));
  INV        o551(.A(ori_ori_n232_), .Y(ori_ori_n574_));
  NA4        o552(.A(ori_ori_n574_), .B(ori_ori_n233_), .C(ori_ori_n126_), .D(ori_ori_n42_), .Y(ori_ori_n575_));
  OAI210     o553(.A0(ori_ori_n575_), .A1(ori_ori_n573_), .B0(ori_ori_n572_), .Y(ori_ori_n576_));
  NO4        o554(.A(ori_ori_n576_), .B(ori_ori_n570_), .C(ori_ori_n567_), .D(ori_ori_n566_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n382_), .B(ori_ori_n28_), .Y(ori_ori_n578_));
  NA2        o556(.A(ori_ori_n543_), .B(ori_ori_n228_), .Y(ori_ori_n579_));
  NA2        o557(.A(ori_ori_n579_), .B(ori_ori_n578_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n62_), .B(i_12_), .Y(ori_ori_n581_));
  NO2        o559(.A(ori_ori_n581_), .B(ori_ori_n128_), .Y(ori_ori_n582_));
  NO2        o560(.A(ori_ori_n582_), .B(ori_ori_n400_), .Y(ori_ori_n583_));
  AOI220     o561(.A0(ori_ori_n583_), .A1(ori_ori_n36_), .B0(ori_ori_n580_), .B1(ori_ori_n46_), .Y(ori_ori_n584_));
  NA4        o562(.A(ori_ori_n584_), .B(ori_ori_n577_), .C(ori_ori_n560_), .D(ori_ori_n550_), .Y(ori6));
  NA4        o563(.A(ori_ori_n279_), .B(ori_ori_n329_), .C(ori_ori_n71_), .D(ori_ori_n102_), .Y(ori_ori_n586_));
  INV        o564(.A(ori_ori_n586_), .Y(ori_ori_n587_));
  NO2        o565(.A(ori_ori_n186_), .B(ori_ori_n332_), .Y(ori_ori_n588_));
  NO2        o566(.A(ori_ori_n587_), .B(ori_ori_n241_), .Y(ori_ori_n589_));
  OR2        o567(.A(ori_ori_n589_), .B(i_12_), .Y(ori_ori_n590_));
  NA2        o568(.A(ori_ori_n386_), .B(ori_ori_n63_), .Y(ori_ori_n591_));
  INV        o569(.A(ori_ori_n591_), .Y(ori_ori_n592_));
  NA2        o570(.A(ori_ori_n592_), .B(ori_ori_n73_), .Y(ori_ori_n593_));
  INV        o571(.A(ori_ori_n240_), .Y(ori_ori_n594_));
  NA2        o572(.A(ori_ori_n75_), .B(ori_ori_n133_), .Y(ori_ori_n595_));
  INV        o573(.A(ori_ori_n126_), .Y(ori_ori_n596_));
  NA2        o574(.A(ori_ori_n596_), .B(ori_ori_n46_), .Y(ori_ori_n597_));
  AOI210     o575(.A0(ori_ori_n597_), .A1(ori_ori_n595_), .B0(ori_ori_n594_), .Y(ori_ori_n598_));
  NO2        o576(.A(ori_ori_n204_), .B(i_9_), .Y(ori_ori_n599_));
  NA2        o577(.A(ori_ori_n599_), .B(ori_ori_n581_), .Y(ori_ori_n600_));
  AOI210     o578(.A0(ori_ori_n600_), .A1(ori_ori_n349_), .B0(ori_ori_n165_), .Y(ori_ori_n601_));
  NO2        o579(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n602_));
  NAi32      o580(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n603_));
  NO2        o581(.A(ori_ori_n516_), .B(ori_ori_n603_), .Y(ori_ori_n604_));
  OR3        o582(.A(ori_ori_n604_), .B(ori_ori_n601_), .C(ori_ori_n598_), .Y(ori_ori_n605_));
  NO2        o583(.A(ori_ori_n493_), .B(i_2_), .Y(ori_ori_n606_));
  NA2        o584(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n607_));
  NO2        o585(.A(ori_ori_n607_), .B(ori_ori_n286_), .Y(ori_ori_n608_));
  NA2        o586(.A(ori_ori_n608_), .B(ori_ori_n606_), .Y(ori_ori_n609_));
  OR2        o587(.A(ori_ori_n425_), .B(ori_ori_n306_), .Y(ori_ori_n610_));
  NA3        o588(.A(ori_ori_n610_), .B(ori_ori_n148_), .C(ori_ori_n69_), .Y(ori_ori_n611_));
  AO210      o589(.A0(ori_ori_n339_), .A1(ori_ori_n547_), .B0(ori_ori_n36_), .Y(ori_ori_n612_));
  NA3        o590(.A(ori_ori_n612_), .B(ori_ori_n611_), .C(ori_ori_n609_), .Y(ori_ori_n613_));
  NO2        o591(.A(i_6_), .B(i_11_), .Y(ori_ori_n614_));
  AOI220     o592(.A0(ori_ori_n614_), .A1(ori_ori_n375_), .B0(ori_ori_n588_), .B1(ori_ori_n510_), .Y(ori_ori_n615_));
  NA3        o593(.A(ori_ori_n267_), .B(ori_ori_n196_), .C(ori_ori_n148_), .Y(ori_ori_n616_));
  NA2        o594(.A(ori_ori_n281_), .B(ori_ori_n70_), .Y(ori_ori_n617_));
  NA4        o595(.A(ori_ori_n617_), .B(ori_ori_n616_), .C(ori_ori_n615_), .D(ori_ori_n408_), .Y(ori_ori_n618_));
  AOI210     o596(.A0(ori_ori_n306_), .A1(ori_ori_n304_), .B0(ori_ori_n374_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n416_), .B(ori_ori_n103_), .Y(ori_ori_n620_));
  OAI210     o598(.A0(ori_ori_n620_), .A1(ori_ori_n113_), .B0(ori_ori_n285_), .Y(ori_ori_n621_));
  INV        o599(.A(ori_ori_n391_), .Y(ori_ori_n622_));
  NA3        o600(.A(ori_ori_n622_), .B(ori_ori_n240_), .C(i_7_), .Y(ori_ori_n623_));
  NA3        o601(.A(ori_ori_n623_), .B(ori_ori_n621_), .C(ori_ori_n619_), .Y(ori_ori_n624_));
  NO4        o602(.A(ori_ori_n624_), .B(ori_ori_n618_), .C(ori_ori_n613_), .D(ori_ori_n605_), .Y(ori_ori_n625_));
  NA4        o603(.A(ori_ori_n625_), .B(ori_ori_n593_), .C(ori_ori_n590_), .D(ori_ori_n275_), .Y(ori3));
  NA2        o604(.A(i_12_), .B(i_10_), .Y(ori_ori_n627_));
  NO2        o605(.A(i_11_), .B(ori_ori_n194_), .Y(ori_ori_n628_));
  NA3        o606(.A(ori_ori_n616_), .B(ori_ori_n408_), .C(ori_ori_n266_), .Y(ori_ori_n629_));
  NA2        o607(.A(ori_ori_n629_), .B(ori_ori_n40_), .Y(ori_ori_n630_));
  NOi21      o608(.An(ori_ori_n97_), .B(ori_ori_n556_), .Y(ori_ori_n631_));
  NO3        o609(.A(ori_ori_n433_), .B(ori_ori_n311_), .C(ori_ori_n133_), .Y(ori_ori_n632_));
  NA2        o610(.A(ori_ori_n287_), .B(ori_ori_n45_), .Y(ori_ori_n633_));
  AN2        o611(.A(ori_ori_n309_), .B(ori_ori_n55_), .Y(ori_ori_n634_));
  NO3        o612(.A(ori_ori_n634_), .B(ori_ori_n632_), .C(ori_ori_n631_), .Y(ori_ori_n635_));
  AOI210     o613(.A0(ori_ori_n635_), .A1(ori_ori_n630_), .B0(ori_ori_n48_), .Y(ori_ori_n636_));
  NO4        o614(.A(ori_ori_n271_), .B(ori_ori_n277_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n637_));
  NA2        o615(.A(ori_ori_n165_), .B(ori_ori_n378_), .Y(ori_ori_n638_));
  NOi31      o616(.An(ori_ori_n638_), .B(ori_ori_n637_), .C(ori_ori_n39_), .Y(ori_ori_n639_));
  NO2        o617(.A(ori_ori_n639_), .B(ori_ori_n63_), .Y(ori_ori_n640_));
  NOi21      o618(.An(i_5_), .B(i_9_), .Y(ori_ori_n641_));
  NA2        o619(.A(ori_ori_n641_), .B(ori_ori_n303_), .Y(ori_ori_n642_));
  BUFFER     o620(.A(ori_ori_n219_), .Y(ori_ori_n643_));
  AOI210     o621(.A0(ori_ori_n643_), .A1(ori_ori_n327_), .B0(ori_ori_n485_), .Y(ori_ori_n644_));
  NO2        o622(.A(ori_ori_n644_), .B(ori_ori_n642_), .Y(ori_ori_n645_));
  NO3        o623(.A(ori_ori_n645_), .B(ori_ori_n640_), .C(ori_ori_n636_), .Y(ori_ori_n646_));
  NA2        o624(.A(ori_ori_n165_), .B(ori_ori_n24_), .Y(ori_ori_n647_));
  INV        o625(.A(ori_ori_n471_), .Y(ori_ori_n648_));
  NO2        o626(.A(ori_ori_n648_), .B(ori_ori_n647_), .Y(ori_ori_n649_));
  INV        o627(.A(ori_ori_n649_), .Y(ori_ori_n650_));
  NA2        o628(.A(ori_ori_n379_), .B(i_0_), .Y(ori_ori_n651_));
  NO4        o629(.A(ori_ori_n390_), .B(ori_ori_n183_), .C(ori_ori_n289_), .D(ori_ori_n286_), .Y(ori_ori_n652_));
  NA2        o630(.A(ori_ori_n652_), .B(i_11_), .Y(ori_ori_n653_));
  NA2        o631(.A(ori_ori_n543_), .B(ori_ori_n241_), .Y(ori_ori_n654_));
  AOI210     o632(.A0(ori_ori_n330_), .A1(ori_ori_n87_), .B0(ori_ori_n58_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n655_), .B(ori_ori_n654_), .Y(ori_ori_n656_));
  NO2        o634(.A(ori_ori_n206_), .B(ori_ori_n152_), .Y(ori_ori_n657_));
  NA2        o635(.A(i_0_), .B(i_10_), .Y(ori_ori_n658_));
  INV        o636(.A(ori_ori_n360_), .Y(ori_ori_n659_));
  NO4        o637(.A(ori_ori_n116_), .B(ori_ori_n58_), .C(ori_ori_n466_), .D(i_5_), .Y(ori_ori_n660_));
  AO220      o638(.A0(ori_ori_n660_), .A1(ori_ori_n659_), .B0(ori_ori_n657_), .B1(i_6_), .Y(ori_ori_n661_));
  NO2        o639(.A(ori_ori_n661_), .B(ori_ori_n656_), .Y(ori_ori_n662_));
  NA3        o640(.A(ori_ori_n662_), .B(ori_ori_n653_), .C(ori_ori_n650_), .Y(ori_ori_n663_));
  NO2        o641(.A(ori_ori_n104_), .B(ori_ori_n37_), .Y(ori_ori_n664_));
  NA2        o642(.A(i_11_), .B(i_9_), .Y(ori_ori_n665_));
  NO3        o643(.A(i_12_), .B(ori_ori_n665_), .C(ori_ori_n407_), .Y(ori_ori_n666_));
  AN2        o644(.A(ori_ori_n666_), .B(ori_ori_n664_), .Y(ori_ori_n667_));
  NA2        o645(.A(ori_ori_n280_), .B(ori_ori_n164_), .Y(ori_ori_n668_));
  NA2        o646(.A(ori_ori_n668_), .B(ori_ori_n156_), .Y(ori_ori_n669_));
  NO2        o647(.A(ori_ori_n665_), .B(ori_ori_n73_), .Y(ori_ori_n670_));
  NO2        o648(.A(ori_ori_n162_), .B(i_0_), .Y(ori_ori_n671_));
  INV        o649(.A(ori_ori_n284_), .Y(ori_ori_n672_));
  NO2        o650(.A(ori_ori_n672_), .B(ori_ori_n642_), .Y(ori_ori_n673_));
  NO3        o651(.A(ori_ori_n673_), .B(ori_ori_n669_), .C(ori_ori_n667_), .Y(ori_ori_n674_));
  NA2        o652(.A(ori_ori_n457_), .B(ori_ori_n123_), .Y(ori_ori_n675_));
  NO2        o653(.A(i_6_), .B(ori_ori_n675_), .Y(ori_ori_n676_));
  AOI210     o654(.A0(ori_ori_n305_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n677_));
  NA2        o655(.A(ori_ori_n160_), .B(ori_ori_n104_), .Y(ori_ori_n678_));
  NOi32      o656(.An(ori_ori_n677_), .Bn(ori_ori_n168_), .C(ori_ori_n678_), .Y(ori_ori_n679_));
  NA2        o657(.A(ori_ori_n409_), .B(ori_ori_n241_), .Y(ori_ori_n680_));
  NO2        o658(.A(ori_ori_n680_), .B(ori_ori_n633_), .Y(ori_ori_n681_));
  NO3        o659(.A(ori_ori_n681_), .B(ori_ori_n679_), .C(ori_ori_n676_), .Y(ori_ori_n682_));
  NOi21      o660(.An(i_7_), .B(i_5_), .Y(ori_ori_n683_));
  INV        o661(.A(ori_ori_n239_), .Y(ori_ori_n684_));
  NA2        o662(.A(ori_ori_n682_), .B(ori_ori_n674_), .Y(ori_ori_n685_));
  NO2        o663(.A(ori_ori_n627_), .B(ori_ori_n238_), .Y(ori_ori_n686_));
  OA210      o664(.A0(ori_ori_n326_), .A1(ori_ori_n189_), .B0(ori_ori_n325_), .Y(ori_ori_n687_));
  NA2        o665(.A(ori_ori_n686_), .B(ori_ori_n670_), .Y(ori_ori_n688_));
  NA2        o666(.A(ori_ori_n670_), .B(ori_ori_n233_), .Y(ori_ori_n689_));
  OAI210     o667(.A0(i_2_), .A1(ori_ori_n167_), .B0(ori_ori_n689_), .Y(ori_ori_n690_));
  NA2        o668(.A(ori_ori_n690_), .B(ori_ori_n326_), .Y(ori_ori_n691_));
  NO2        o669(.A(ori_ori_n75_), .B(ori_ori_n545_), .Y(ori_ori_n692_));
  NA2        o670(.A(ori_ori_n692_), .B(i_11_), .Y(ori_ori_n693_));
  NO2        o671(.A(ori_ori_n693_), .B(ori_ori_n47_), .Y(ori_ori_n694_));
  NA2        o672(.A(ori_ori_n495_), .B(ori_ori_n362_), .Y(ori_ori_n695_));
  NAi21      o673(.An(i_9_), .B(i_5_), .Y(ori_ori_n696_));
  NO2        o674(.A(ori_ori_n696_), .B(ori_ori_n283_), .Y(ori_ori_n697_));
  NO2        o675(.A(ori_ori_n403_), .B(ori_ori_n106_), .Y(ori_ori_n698_));
  AOI220     o676(.A0(ori_ori_n698_), .A1(i_0_), .B0(ori_ori_n697_), .B1(ori_ori_n425_), .Y(ori_ori_n699_));
  OAI220     o677(.A0(ori_ori_n699_), .A1(ori_ori_n86_), .B0(ori_ori_n695_), .B1(ori_ori_n161_), .Y(ori_ori_n700_));
  NO3        o678(.A(ori_ori_n700_), .B(ori_ori_n694_), .C(ori_ori_n353_), .Y(ori_ori_n701_));
  NA3        o679(.A(ori_ori_n701_), .B(ori_ori_n691_), .C(ori_ori_n688_), .Y(ori_ori_n702_));
  NO3        o680(.A(ori_ori_n702_), .B(ori_ori_n685_), .C(ori_ori_n663_), .Y(ori_ori_n703_));
  NO2        o681(.A(i_0_), .B(ori_ori_n522_), .Y(ori_ori_n704_));
  AOI210     o682(.A0(ori_ori_n591_), .A1(ori_ori_n484_), .B0(ori_ori_n678_), .Y(ori_ori_n705_));
  INV        o683(.A(ori_ori_n705_), .Y(ori_ori_n706_));
  OAI210     o684(.A0(ori_ori_n200_), .A1(i_9_), .B0(ori_ori_n192_), .Y(ori_ori_n707_));
  AOI210     o685(.A0(ori_ori_n707_), .A1(ori_ori_n651_), .B0(ori_ori_n152_), .Y(ori_ori_n708_));
  INV        o686(.A(ori_ori_n708_), .Y(ori_ori_n709_));
  NA2        o687(.A(ori_ori_n709_), .B(ori_ori_n706_), .Y(ori_ori_n710_));
  NO3        o688(.A(ori_ori_n658_), .B(ori_ori_n641_), .C(ori_ori_n169_), .Y(ori_ori_n711_));
  AOI220     o689(.A0(ori_ori_n711_), .A1(i_11_), .B0(ori_ori_n377_), .B1(ori_ori_n75_), .Y(ori_ori_n712_));
  NO3        o690(.A(ori_ori_n179_), .B(ori_ori_n277_), .C(i_0_), .Y(ori_ori_n713_));
  OAI210     o691(.A0(ori_ori_n713_), .A1(ori_ori_n76_), .B0(i_13_), .Y(ori_ori_n714_));
  NA2        o692(.A(ori_ori_n714_), .B(ori_ori_n712_), .Y(ori_ori_n715_));
  NO2        o693(.A(ori_ori_n199_), .B(ori_ori_n93_), .Y(ori_ori_n716_));
  AOI210     o694(.A0(ori_ori_n716_), .A1(ori_ori_n704_), .B0(ori_ori_n110_), .Y(ori_ori_n717_));
  OR2        o695(.A(ori_ori_n717_), .B(i_5_), .Y(ori_ori_n718_));
  AOI210     o696(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n162_), .Y(ori_ori_n719_));
  NA2        o697(.A(ori_ori_n719_), .B(ori_ori_n687_), .Y(ori_ori_n720_));
  NO3        o698(.A(ori_ori_n633_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n721_));
  NA2        o699(.A(ori_ori_n338_), .B(ori_ori_n331_), .Y(ori_ori_n722_));
  NO2        o700(.A(ori_ori_n722_), .B(ori_ori_n721_), .Y(ori_ori_n723_));
  NA3        o701(.A(ori_ori_n279_), .B(ori_ori_n160_), .C(ori_ori_n159_), .Y(ori_ori_n724_));
  INV        o702(.A(ori_ori_n724_), .Y(ori_ori_n725_));
  NO3        o703(.A(ori_ori_n665_), .B(ori_ori_n185_), .C(ori_ori_n169_), .Y(ori_ori_n726_));
  NO2        o704(.A(ori_ori_n726_), .B(ori_ori_n725_), .Y(ori_ori_n727_));
  NA4        o705(.A(ori_ori_n727_), .B(ori_ori_n723_), .C(ori_ori_n720_), .D(ori_ori_n718_), .Y(ori_ori_n728_));
  NO2        o706(.A(ori_ori_n86_), .B(i_5_), .Y(ori_ori_n729_));
  NA3        o707(.A(ori_ori_n628_), .B(ori_ori_n111_), .C(ori_ori_n126_), .Y(ori_ori_n730_));
  INV        o708(.A(ori_ori_n730_), .Y(ori_ori_n731_));
  NA2        o709(.A(ori_ori_n731_), .B(ori_ori_n729_), .Y(ori_ori_n732_));
  NAi21      o710(.An(ori_ori_n198_), .B(ori_ori_n199_), .Y(ori_ori_n733_));
  NO4        o711(.A(ori_ori_n197_), .B(ori_ori_n179_), .C(i_0_), .D(i_12_), .Y(ori_ori_n734_));
  AOI220     o712(.A0(ori_ori_n734_), .A1(ori_ori_n733_), .B0(ori_ori_n587_), .B1(ori_ori_n163_), .Y(ori_ori_n735_));
  NA2        o713(.A(ori_ori_n683_), .B(ori_ori_n324_), .Y(ori_ori_n736_));
  NO2        o714(.A(ori_ori_n736_), .B(ori_ori_n474_), .Y(ori_ori_n737_));
  NA2        o715(.A(ori_ori_n737_), .B(ori_ori_n671_), .Y(ori_ori_n738_));
  NA3        o716(.A(ori_ori_n738_), .B(ori_ori_n735_), .C(ori_ori_n732_), .Y(ori_ori_n739_));
  NO4        o717(.A(ori_ori_n739_), .B(ori_ori_n728_), .C(ori_ori_n715_), .D(ori_ori_n710_), .Y(ori_ori_n740_));
  OAI210     o718(.A0(ori_ori_n606_), .A1(ori_ori_n602_), .B0(ori_ori_n37_), .Y(ori_ori_n741_));
  NA2        o719(.A(ori_ori_n741_), .B(ori_ori_n415_), .Y(ori_ori_n742_));
  NA2        o720(.A(ori_ori_n742_), .B(ori_ori_n177_), .Y(ori_ori_n743_));
  NA2        o721(.A(ori_ori_n166_), .B(ori_ori_n168_), .Y(ori_ori_n744_));
  AO210      o722(.A0(ori_ori_n493_), .A1(ori_ori_n33_), .B0(ori_ori_n744_), .Y(ori_ori_n745_));
  NAi31      o723(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n746_));
  AOI210     o724(.A0(ori_ori_n119_), .A1(ori_ori_n70_), .B0(ori_ori_n746_), .Y(ori_ori_n747_));
  NO2        o725(.A(ori_ori_n747_), .B(ori_ori_n446_), .Y(ori_ori_n748_));
  NA2        o726(.A(ori_ori_n748_), .B(ori_ori_n745_), .Y(ori_ori_n749_));
  NO2        o727(.A(ori_ori_n319_), .B(ori_ori_n219_), .Y(ori_ori_n750_));
  NO2        o728(.A(ori_ori_n750_), .B(ori_ori_n652_), .Y(ori_ori_n751_));
  INV        o729(.A(ori_ori_n751_), .Y(ori_ori_n752_));
  AOI210     o730(.A0(ori_ori_n749_), .A1(ori_ori_n48_), .B0(ori_ori_n752_), .Y(ori_ori_n753_));
  AOI210     o731(.A0(ori_ori_n753_), .A1(ori_ori_n743_), .B0(ori_ori_n73_), .Y(ori_ori_n754_));
  INV        o732(.A(ori_ori_n274_), .Y(ori_ori_n755_));
  NO2        o733(.A(ori_ori_n755_), .B(ori_ori_n551_), .Y(ori_ori_n756_));
  OAI210     o734(.A0(ori_ori_n221_), .A1(ori_ori_n154_), .B0(ori_ori_n87_), .Y(ori_ori_n757_));
  NO2        o735(.A(ori_ori_n757_), .B(i_11_), .Y(ori_ori_n758_));
  NO3        o736(.A(ori_ori_n59_), .B(ori_ori_n58_), .C(i_4_), .Y(ori_ori_n759_));
  OAI210     o737(.A0(ori_ori_n684_), .A1(ori_ori_n234_), .B0(ori_ori_n759_), .Y(ori_ori_n760_));
  NO2        o738(.A(ori_ori_n760_), .B(ori_ori_n522_), .Y(ori_ori_n761_));
  INV        o739(.A(ori_ori_n374_), .Y(ori_ori_n762_));
  NO2        o740(.A(ori_ori_n604_), .B(ori_ori_n255_), .Y(ori_ori_n763_));
  AOI210     o741(.A0(ori_ori_n763_), .A1(ori_ori_n762_), .B0(ori_ori_n41_), .Y(ori_ori_n764_));
  NO3        o742(.A(ori_ori_n764_), .B(ori_ori_n761_), .C(ori_ori_n758_), .Y(ori_ori_n765_));
  INV        o743(.A(ori_ori_n765_), .Y(ori_ori_n766_));
  NO3        o744(.A(ori_ori_n766_), .B(ori_ori_n756_), .C(ori_ori_n754_), .Y(ori_ori_n767_));
  NA4        o745(.A(ori_ori_n767_), .B(ori_ori_n740_), .C(ori_ori_n703_), .D(ori_ori_n646_), .Y(ori4));
  INV        o746(.A(ori_ori_n494_), .Y(ori_ori_n771_));
  INV        o747(.A(i_6_), .Y(ori_ori_n772_));
  INV        o748(.A(ori_ori_n202_), .Y(ori_ori_n773_));
  NAi21      m0000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m0001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m0002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m0003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m0004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m0005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m0006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m0007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m0008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m0010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m0011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m0012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m0013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m0014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m0015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m0016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m0017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m0018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m0019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m0021(.A(mai_mai_n35_), .Y(mai1));
  INV        m0022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m0023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m0024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m0025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m0026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m0027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m0028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m0029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m0030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m0031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m0032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NA2        m0033(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n56_));
  NA3        m0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n57_));
  NO2        m0035(.A(i_1_), .B(i_6_), .Y(mai_mai_n58_));
  NA2        m0036(.A(i_8_), .B(i_7_), .Y(mai_mai_n59_));
  OAI210     m0037(.A0(mai_mai_n59_), .A1(mai_mai_n58_), .B0(mai_mai_n57_), .Y(mai_mai_n60_));
  NA2        m0038(.A(mai_mai_n60_), .B(i_12_), .Y(mai_mai_n61_));
  NAi21      m0039(.An(i_2_), .B(i_7_), .Y(mai_mai_n62_));
  INV        m0040(.A(i_1_), .Y(mai_mai_n63_));
  NA2        m0041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NA3        m0042(.A(mai_mai_n64_), .B(mai_mai_n62_), .C(mai_mai_n31_), .Y(mai_mai_n65_));
  NA2        m0043(.A(i_1_), .B(i_10_), .Y(mai_mai_n66_));
  NO2        m0044(.A(mai_mai_n66_), .B(i_6_), .Y(mai_mai_n67_));
  NAi31      m0045(.An(mai_mai_n67_), .B(mai_mai_n65_), .C(mai_mai_n61_), .Y(mai_mai_n68_));
  NA2        m0046(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n69_));
  AOI210     m0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n70_));
  NA2        m0048(.A(i_1_), .B(i_6_), .Y(mai_mai_n71_));
  NO2        m0049(.A(mai_mai_n71_), .B(mai_mai_n25_), .Y(mai_mai_n72_));
  INV        m0050(.A(i_0_), .Y(mai_mai_n73_));
  NAi21      m0051(.An(i_5_), .B(i_10_), .Y(mai_mai_n74_));
  NA2        m0052(.A(i_5_), .B(i_9_), .Y(mai_mai_n75_));
  AOI210     m0053(.A0(mai_mai_n75_), .A1(mai_mai_n74_), .B0(mai_mai_n73_), .Y(mai_mai_n76_));
  NO2        m0054(.A(mai_mai_n76_), .B(mai_mai_n72_), .Y(mai_mai_n77_));
  OAI210     m0055(.A0(mai_mai_n70_), .A1(mai_mai_n69_), .B0(mai_mai_n77_), .Y(mai_mai_n78_));
  OAI210     m0056(.A0(mai_mai_n78_), .A1(mai_mai_n68_), .B0(i_0_), .Y(mai_mai_n79_));
  NA2        m0057(.A(i_12_), .B(i_5_), .Y(mai_mai_n80_));
  NA2        m0058(.A(i_2_), .B(i_8_), .Y(mai_mai_n81_));
  NO2        m0059(.A(mai_mai_n81_), .B(mai_mai_n58_), .Y(mai_mai_n82_));
  NO2        m0060(.A(i_3_), .B(i_9_), .Y(mai_mai_n83_));
  NO2        m0061(.A(i_3_), .B(i_7_), .Y(mai_mai_n84_));
  NO3        m0062(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(mai_mai_n63_), .Y(mai_mai_n85_));
  INV        m0063(.A(i_6_), .Y(mai_mai_n86_));
  OR4        m0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n87_));
  INV        m0065(.A(mai_mai_n87_), .Y(mai_mai_n88_));
  NO2        m0066(.A(i_2_), .B(i_7_), .Y(mai_mai_n89_));
  AOI210     m0067(.A0(mai_mai_n88_), .A1(mai_mai_n86_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  OAI210     m0068(.A0(mai_mai_n85_), .A1(mai_mai_n82_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  NAi21      m0069(.An(i_6_), .B(i_10_), .Y(mai_mai_n92_));
  NA2        m0070(.A(i_6_), .B(i_9_), .Y(mai_mai_n93_));
  AOI210     m0071(.A0(mai_mai_n93_), .A1(mai_mai_n92_), .B0(mai_mai_n63_), .Y(mai_mai_n94_));
  NA2        m0072(.A(i_2_), .B(i_6_), .Y(mai_mai_n95_));
  INV        m0073(.A(mai_mai_n94_), .Y(mai_mai_n96_));
  AOI210     m0074(.A0(mai_mai_n96_), .A1(mai_mai_n91_), .B0(mai_mai_n80_), .Y(mai_mai_n97_));
  AN3        m0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n98_));
  NAi21      m0076(.An(i_6_), .B(i_11_), .Y(mai_mai_n99_));
  NO2        m0077(.A(i_5_), .B(i_8_), .Y(mai_mai_n100_));
  NOi21      m0078(.An(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  AOI220     m0079(.A0(mai_mai_n101_), .A1(mai_mai_n62_), .B0(mai_mai_n98_), .B1(mai_mai_n32_), .Y(mai_mai_n102_));
  INV        m0080(.A(i_7_), .Y(mai_mai_n103_));
  NA2        m0081(.A(mai_mai_n47_), .B(mai_mai_n103_), .Y(mai_mai_n104_));
  NO2        m0082(.A(i_0_), .B(i_5_), .Y(mai_mai_n105_));
  NO2        m0083(.A(mai_mai_n105_), .B(mai_mai_n86_), .Y(mai_mai_n106_));
  NA2        m0084(.A(i_12_), .B(i_3_), .Y(mai_mai_n107_));
  INV        m0085(.A(mai_mai_n107_), .Y(mai_mai_n108_));
  NA3        m0086(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n104_), .Y(mai_mai_n109_));
  NAi21      m0087(.An(i_7_), .B(i_11_), .Y(mai_mai_n110_));
  AN2        m0088(.A(i_2_), .B(i_10_), .Y(mai_mai_n111_));
  NO2        m0089(.A(mai_mai_n111_), .B(i_7_), .Y(mai_mai_n112_));
  OR2        m0090(.A(mai_mai_n80_), .B(mai_mai_n58_), .Y(mai_mai_n113_));
  NO2        m0091(.A(i_8_), .B(mai_mai_n103_), .Y(mai_mai_n114_));
  NO3        m0092(.A(mai_mai_n114_), .B(mai_mai_n113_), .C(mai_mai_n112_), .Y(mai_mai_n115_));
  NA2        m0093(.A(i_12_), .B(i_7_), .Y(mai_mai_n116_));
  NA2        m0094(.A(i_11_), .B(i_12_), .Y(mai_mai_n117_));
  INV        m0095(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NO2        m0096(.A(mai_mai_n118_), .B(mai_mai_n115_), .Y(mai_mai_n119_));
  NA3        m0097(.A(mai_mai_n119_), .B(mai_mai_n109_), .C(mai_mai_n102_), .Y(mai_mai_n120_));
  NOi21      m0098(.An(i_1_), .B(i_5_), .Y(mai_mai_n121_));
  NA2        m0099(.A(mai_mai_n121_), .B(i_11_), .Y(mai_mai_n122_));
  NA2        m0100(.A(mai_mai_n103_), .B(mai_mai_n37_), .Y(mai_mai_n123_));
  NA2        m0101(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n124_));
  NA2        m0102(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n125_));
  NO2        m0103(.A(mai_mai_n125_), .B(mai_mai_n47_), .Y(mai_mai_n126_));
  NA2        m0104(.A(mai_mai_n93_), .B(mai_mai_n92_), .Y(mai_mai_n127_));
  NAi21      m0105(.An(i_3_), .B(i_8_), .Y(mai_mai_n128_));
  NA2        m0106(.A(mai_mai_n128_), .B(mai_mai_n62_), .Y(mai_mai_n129_));
  NOi31      m0107(.An(mai_mai_n129_), .B(mai_mai_n127_), .C(mai_mai_n126_), .Y(mai_mai_n130_));
  NO2        m0108(.A(i_1_), .B(mai_mai_n86_), .Y(mai_mai_n131_));
  NO2        m0109(.A(i_6_), .B(i_5_), .Y(mai_mai_n132_));
  NA2        m0110(.A(mai_mai_n132_), .B(i_3_), .Y(mai_mai_n133_));
  AO210      m0111(.A0(mai_mai_n133_), .A1(mai_mai_n48_), .B0(mai_mai_n131_), .Y(mai_mai_n134_));
  OAI220     m0112(.A0(mai_mai_n134_), .A1(mai_mai_n110_), .B0(mai_mai_n130_), .B1(mai_mai_n122_), .Y(mai_mai_n135_));
  NO3        m0113(.A(mai_mai_n135_), .B(mai_mai_n120_), .C(mai_mai_n97_), .Y(mai_mai_n136_));
  NA3        m0114(.A(mai_mai_n136_), .B(mai_mai_n79_), .C(mai_mai_n56_), .Y(mai2));
  NO2        m0115(.A(mai_mai_n63_), .B(mai_mai_n37_), .Y(mai_mai_n138_));
  NA2        m0116(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n139_));
  NA2        m0117(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NA4        m0118(.A(mai_mai_n140_), .B(mai_mai_n77_), .C(mai_mai_n69_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m0119(.A(i_8_), .B(i_7_), .Y(mai_mai_n142_));
  NA2        m0120(.A(mai_mai_n142_), .B(i_6_), .Y(mai_mai_n143_));
  NO2        m0121(.A(i_12_), .B(i_13_), .Y(mai_mai_n144_));
  NAi21      m0122(.An(i_5_), .B(i_11_), .Y(mai_mai_n145_));
  NOi21      m0123(.An(mai_mai_n144_), .B(mai_mai_n145_), .Y(mai_mai_n146_));
  NO2        m0124(.A(i_0_), .B(i_1_), .Y(mai_mai_n147_));
  NA2        m0125(.A(i_2_), .B(i_3_), .Y(mai_mai_n148_));
  NO2        m0126(.A(mai_mai_n148_), .B(i_4_), .Y(mai_mai_n149_));
  NA3        m0127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n150_));
  AN2        m0128(.A(mai_mai_n144_), .B(mai_mai_n83_), .Y(mai_mai_n151_));
  NO2        m0129(.A(mai_mai_n151_), .B(mai_mai_n27_), .Y(mai_mai_n152_));
  NA2        m0130(.A(i_1_), .B(i_5_), .Y(mai_mai_n153_));
  NO2        m0131(.A(mai_mai_n73_), .B(mai_mai_n47_), .Y(mai_mai_n154_));
  NA2        m0132(.A(mai_mai_n154_), .B(mai_mai_n36_), .Y(mai_mai_n155_));
  NO3        m0133(.A(mai_mai_n155_), .B(mai_mai_n153_), .C(mai_mai_n152_), .Y(mai_mai_n156_));
  OR2        m0134(.A(i_0_), .B(i_1_), .Y(mai_mai_n157_));
  NO3        m0135(.A(mai_mai_n157_), .B(mai_mai_n80_), .C(i_13_), .Y(mai_mai_n158_));
  NAi32      m0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n159_));
  NAi21      m0137(.An(mai_mai_n159_), .B(mai_mai_n158_), .Y(mai_mai_n160_));
  NOi21      m0138(.An(i_4_), .B(i_10_), .Y(mai_mai_n161_));
  NA2        m0139(.A(mai_mai_n161_), .B(mai_mai_n40_), .Y(mai_mai_n162_));
  NO2        m0140(.A(i_3_), .B(i_5_), .Y(mai_mai_n163_));
  NO3        m0141(.A(mai_mai_n73_), .B(i_2_), .C(i_1_), .Y(mai_mai_n164_));
  NA2        m0142(.A(mai_mai_n164_), .B(mai_mai_n163_), .Y(mai_mai_n165_));
  OAI210     m0143(.A0(mai_mai_n165_), .A1(mai_mai_n162_), .B0(mai_mai_n160_), .Y(mai_mai_n166_));
  NO2        m0144(.A(mai_mai_n166_), .B(mai_mai_n156_), .Y(mai_mai_n167_));
  AOI210     m0145(.A0(mai_mai_n167_), .A1(mai_mai_n150_), .B0(mai_mai_n143_), .Y(mai_mai_n168_));
  NA3        m0146(.A(mai_mai_n73_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n169_));
  NA2        m0147(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n170_));
  NOi21      m0148(.An(i_4_), .B(i_9_), .Y(mai_mai_n171_));
  NOi21      m0149(.An(i_11_), .B(i_13_), .Y(mai_mai_n172_));
  NA2        m0150(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  OR2        m0151(.A(mai_mai_n173_), .B(mai_mai_n170_), .Y(mai_mai_n174_));
  NO2        m0152(.A(i_4_), .B(i_5_), .Y(mai_mai_n175_));
  NAi21      m0153(.An(i_12_), .B(i_11_), .Y(mai_mai_n176_));
  NO2        m0154(.A(mai_mai_n176_), .B(i_13_), .Y(mai_mai_n177_));
  NA3        m0155(.A(mai_mai_n177_), .B(mai_mai_n175_), .C(mai_mai_n83_), .Y(mai_mai_n178_));
  AOI210     m0156(.A0(mai_mai_n178_), .A1(mai_mai_n174_), .B0(mai_mai_n169_), .Y(mai_mai_n179_));
  NO2        m0157(.A(mai_mai_n73_), .B(mai_mai_n63_), .Y(mai_mai_n180_));
  NA2        m0158(.A(mai_mai_n180_), .B(mai_mai_n47_), .Y(mai_mai_n181_));
  NA2        m0159(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n182_));
  NAi31      m0160(.An(mai_mai_n182_), .B(mai_mai_n151_), .C(i_11_), .Y(mai_mai_n183_));
  NA2        m0161(.A(i_3_), .B(i_5_), .Y(mai_mai_n184_));
  OR2        m0162(.A(mai_mai_n184_), .B(mai_mai_n173_), .Y(mai_mai_n185_));
  AOI210     m0163(.A0(mai_mai_n185_), .A1(mai_mai_n183_), .B0(mai_mai_n181_), .Y(mai_mai_n186_));
  NO2        m0164(.A(mai_mai_n73_), .B(i_5_), .Y(mai_mai_n187_));
  NO2        m0165(.A(i_13_), .B(i_10_), .Y(mai_mai_n188_));
  NA3        m0166(.A(mai_mai_n188_), .B(mai_mai_n187_), .C(mai_mai_n45_), .Y(mai_mai_n189_));
  NO2        m0167(.A(i_2_), .B(i_1_), .Y(mai_mai_n190_));
  NA2        m0168(.A(mai_mai_n190_), .B(i_3_), .Y(mai_mai_n191_));
  NAi21      m0169(.An(i_4_), .B(i_12_), .Y(mai_mai_n192_));
  NO4        m0170(.A(mai_mai_n192_), .B(mai_mai_n191_), .C(mai_mai_n189_), .D(mai_mai_n25_), .Y(mai_mai_n193_));
  NO3        m0171(.A(mai_mai_n193_), .B(mai_mai_n186_), .C(mai_mai_n179_), .Y(mai_mai_n194_));
  INV        m0172(.A(i_8_), .Y(mai_mai_n195_));
  NO2        m0173(.A(mai_mai_n195_), .B(i_7_), .Y(mai_mai_n196_));
  NA2        m0174(.A(mai_mai_n196_), .B(i_6_), .Y(mai_mai_n197_));
  NO3        m0175(.A(i_3_), .B(mai_mai_n86_), .C(mai_mai_n49_), .Y(mai_mai_n198_));
  NA2        m0176(.A(mai_mai_n198_), .B(mai_mai_n114_), .Y(mai_mai_n199_));
  NO3        m0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n200_));
  NA3        m0178(.A(mai_mai_n200_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n201_));
  NO3        m0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n202_));
  OAI210     m0180(.A0(mai_mai_n98_), .A1(i_12_), .B0(mai_mai_n202_), .Y(mai_mai_n203_));
  AOI210     m0181(.A0(mai_mai_n203_), .A1(mai_mai_n201_), .B0(mai_mai_n199_), .Y(mai_mai_n204_));
  NO2        m0182(.A(i_3_), .B(i_8_), .Y(mai_mai_n205_));
  NO3        m0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n206_));
  NA3        m0184(.A(mai_mai_n206_), .B(mai_mai_n205_), .C(mai_mai_n40_), .Y(mai_mai_n207_));
  NO2        m0185(.A(mai_mai_n105_), .B(mai_mai_n58_), .Y(mai_mai_n208_));
  NO2        m0186(.A(i_13_), .B(i_9_), .Y(mai_mai_n209_));
  NA3        m0187(.A(mai_mai_n209_), .B(i_6_), .C(mai_mai_n195_), .Y(mai_mai_n210_));
  NAi21      m0188(.An(i_12_), .B(i_3_), .Y(mai_mai_n211_));
  NO2        m0189(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n212_));
  NO3        m0190(.A(i_0_), .B(i_2_), .C(mai_mai_n63_), .Y(mai_mai_n213_));
  NA3        m0191(.A(mai_mai_n213_), .B(mai_mai_n212_), .C(i_10_), .Y(mai_mai_n214_));
  NO2        m0192(.A(mai_mai_n214_), .B(mai_mai_n210_), .Y(mai_mai_n215_));
  AOI210     m0193(.A0(mai_mai_n215_), .A1(i_7_), .B0(mai_mai_n204_), .Y(mai_mai_n216_));
  OAI220     m0194(.A0(mai_mai_n216_), .A1(i_4_), .B0(mai_mai_n197_), .B1(mai_mai_n194_), .Y(mai_mai_n217_));
  NAi21      m0195(.An(i_12_), .B(i_7_), .Y(mai_mai_n218_));
  NA3        m0196(.A(i_13_), .B(mai_mai_n195_), .C(i_10_), .Y(mai_mai_n219_));
  NO2        m0197(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n220_));
  NA2        m0198(.A(i_0_), .B(i_5_), .Y(mai_mai_n221_));
  NA2        m0199(.A(mai_mai_n221_), .B(mai_mai_n106_), .Y(mai_mai_n222_));
  OAI220     m0200(.A0(mai_mai_n222_), .A1(mai_mai_n191_), .B0(mai_mai_n181_), .B1(mai_mai_n133_), .Y(mai_mai_n223_));
  NAi31      m0201(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n224_));
  NO2        m0202(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n225_));
  NO2        m0203(.A(mai_mai_n73_), .B(mai_mai_n26_), .Y(mai_mai_n226_));
  NO2        m0204(.A(mai_mai_n47_), .B(mai_mai_n63_), .Y(mai_mai_n227_));
  NA3        m0205(.A(mai_mai_n227_), .B(mai_mai_n226_), .C(mai_mai_n225_), .Y(mai_mai_n228_));
  INV        m0206(.A(i_13_), .Y(mai_mai_n229_));
  NO2        m0207(.A(i_12_), .B(mai_mai_n229_), .Y(mai_mai_n230_));
  NA3        m0208(.A(mai_mai_n230_), .B(mai_mai_n200_), .C(mai_mai_n198_), .Y(mai_mai_n231_));
  OAI210     m0209(.A0(mai_mai_n228_), .A1(mai_mai_n224_), .B0(mai_mai_n231_), .Y(mai_mai_n232_));
  AOI220     m0210(.A0(mai_mai_n232_), .A1(mai_mai_n142_), .B0(mai_mai_n223_), .B1(mai_mai_n220_), .Y(mai_mai_n233_));
  NO2        m0211(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n234_));
  NO2        m0212(.A(mai_mai_n184_), .B(i_4_), .Y(mai_mai_n235_));
  NA2        m0213(.A(mai_mai_n235_), .B(mai_mai_n234_), .Y(mai_mai_n236_));
  OR2        m0214(.A(i_8_), .B(i_7_), .Y(mai_mai_n237_));
  NO2        m0215(.A(mai_mai_n237_), .B(mai_mai_n86_), .Y(mai_mai_n238_));
  NO2        m0216(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n239_));
  NA2        m0217(.A(mai_mai_n239_), .B(mai_mai_n238_), .Y(mai_mai_n240_));
  INV        m0218(.A(i_12_), .Y(mai_mai_n241_));
  NO2        m0219(.A(mai_mai_n45_), .B(mai_mai_n241_), .Y(mai_mai_n242_));
  NO3        m0220(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n243_));
  NA2        m0221(.A(i_2_), .B(i_1_), .Y(mai_mai_n244_));
  NO2        m0222(.A(mai_mai_n240_), .B(mai_mai_n236_), .Y(mai_mai_n245_));
  NO3        m0223(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n246_));
  NAi21      m0224(.An(i_4_), .B(i_3_), .Y(mai_mai_n247_));
  NO2        m0225(.A(mai_mai_n247_), .B(mai_mai_n75_), .Y(mai_mai_n248_));
  NO2        m0226(.A(i_0_), .B(i_6_), .Y(mai_mai_n249_));
  NOi41      m0227(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n250_));
  NA2        m0228(.A(mai_mai_n250_), .B(mai_mai_n249_), .Y(mai_mai_n251_));
  NO2        m0229(.A(mai_mai_n244_), .B(mai_mai_n184_), .Y(mai_mai_n252_));
  NAi21      m0230(.An(mai_mai_n251_), .B(mai_mai_n252_), .Y(mai_mai_n253_));
  INV        m0231(.A(mai_mai_n253_), .Y(mai_mai_n254_));
  AOI220     m0232(.A0(mai_mai_n254_), .A1(mai_mai_n40_), .B0(mai_mai_n245_), .B1(mai_mai_n209_), .Y(mai_mai_n255_));
  NO2        m0233(.A(i_11_), .B(mai_mai_n229_), .Y(mai_mai_n256_));
  NOi21      m0234(.An(i_1_), .B(i_6_), .Y(mai_mai_n257_));
  NAi21      m0235(.An(i_3_), .B(i_7_), .Y(mai_mai_n258_));
  NA2        m0236(.A(mai_mai_n241_), .B(i_9_), .Y(mai_mai_n259_));
  OR4        m0237(.A(mai_mai_n259_), .B(mai_mai_n258_), .C(mai_mai_n257_), .D(mai_mai_n187_), .Y(mai_mai_n260_));
  NO2        m0238(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n261_));
  NO2        m0239(.A(i_12_), .B(i_3_), .Y(mai_mai_n262_));
  NA2        m0240(.A(mai_mai_n73_), .B(i_5_), .Y(mai_mai_n263_));
  NA2        m0241(.A(i_3_), .B(i_9_), .Y(mai_mai_n264_));
  NAi21      m0242(.An(i_7_), .B(i_10_), .Y(mai_mai_n265_));
  NO2        m0243(.A(mai_mai_n265_), .B(mai_mai_n264_), .Y(mai_mai_n266_));
  NA3        m0244(.A(mai_mai_n266_), .B(mai_mai_n263_), .C(mai_mai_n64_), .Y(mai_mai_n267_));
  NA2        m0245(.A(mai_mai_n267_), .B(mai_mai_n260_), .Y(mai_mai_n268_));
  NA3        m0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n269_));
  INV        m0247(.A(mai_mai_n143_), .Y(mai_mai_n270_));
  NA2        m0248(.A(mai_mai_n241_), .B(i_13_), .Y(mai_mai_n271_));
  NO2        m0249(.A(mai_mai_n271_), .B(mai_mai_n75_), .Y(mai_mai_n272_));
  AOI220     m0250(.A0(mai_mai_n272_), .A1(mai_mai_n270_), .B0(mai_mai_n268_), .B1(mai_mai_n256_), .Y(mai_mai_n273_));
  NO2        m0251(.A(mai_mai_n237_), .B(mai_mai_n37_), .Y(mai_mai_n274_));
  NA2        m0252(.A(i_12_), .B(i_6_), .Y(mai_mai_n275_));
  OR2        m0253(.A(i_13_), .B(i_9_), .Y(mai_mai_n276_));
  NO2        m0254(.A(mai_mai_n247_), .B(i_2_), .Y(mai_mai_n277_));
  NA2        m0255(.A(mai_mai_n256_), .B(i_9_), .Y(mai_mai_n278_));
  NA2        m0256(.A(mai_mai_n154_), .B(mai_mai_n63_), .Y(mai_mai_n279_));
  NO3        m0257(.A(i_11_), .B(mai_mai_n229_), .C(mai_mai_n25_), .Y(mai_mai_n280_));
  NO2        m0258(.A(mai_mai_n258_), .B(i_8_), .Y(mai_mai_n281_));
  NO2        m0259(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n282_));
  NA3        m0260(.A(mai_mai_n282_), .B(mai_mai_n281_), .C(mai_mai_n280_), .Y(mai_mai_n283_));
  NO3        m0261(.A(mai_mai_n26_), .B(mai_mai_n86_), .C(i_5_), .Y(mai_mai_n284_));
  NA3        m0262(.A(mai_mai_n284_), .B(mai_mai_n274_), .C(mai_mai_n230_), .Y(mai_mai_n285_));
  AOI210     m0263(.A0(mai_mai_n285_), .A1(mai_mai_n283_), .B0(mai_mai_n279_), .Y(mai_mai_n286_));
  INV        m0264(.A(mai_mai_n286_), .Y(mai_mai_n287_));
  NA4        m0265(.A(mai_mai_n287_), .B(mai_mai_n273_), .C(mai_mai_n255_), .D(mai_mai_n233_), .Y(mai_mai_n288_));
  NO3        m0266(.A(i_12_), .B(mai_mai_n229_), .C(mai_mai_n37_), .Y(mai_mai_n289_));
  INV        m0267(.A(mai_mai_n289_), .Y(mai_mai_n290_));
  NA2        m0268(.A(i_8_), .B(mai_mai_n103_), .Y(mai_mai_n291_));
  NOi21      m0269(.An(mai_mai_n163_), .B(mai_mai_n86_), .Y(mai_mai_n292_));
  NO3        m0270(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n293_));
  AOI220     m0271(.A0(mai_mai_n293_), .A1(mai_mai_n198_), .B0(mai_mai_n292_), .B1(mai_mai_n239_), .Y(mai_mai_n294_));
  NO2        m0272(.A(mai_mai_n294_), .B(mai_mai_n291_), .Y(mai_mai_n295_));
  NO3        m0273(.A(i_0_), .B(i_2_), .C(mai_mai_n63_), .Y(mai_mai_n296_));
  NO2        m0274(.A(mai_mai_n244_), .B(i_0_), .Y(mai_mai_n297_));
  AOI220     m0275(.A0(mai_mai_n297_), .A1(mai_mai_n196_), .B0(mai_mai_n296_), .B1(mai_mai_n142_), .Y(mai_mai_n298_));
  NA2        m0276(.A(mai_mai_n282_), .B(mai_mai_n26_), .Y(mai_mai_n299_));
  NO2        m0277(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n300_));
  NA2        m0278(.A(i_0_), .B(i_1_), .Y(mai_mai_n301_));
  NO2        m0279(.A(mai_mai_n301_), .B(i_2_), .Y(mai_mai_n302_));
  NO2        m0280(.A(mai_mai_n59_), .B(i_6_), .Y(mai_mai_n303_));
  NA3        m0281(.A(mai_mai_n303_), .B(mai_mai_n302_), .C(mai_mai_n163_), .Y(mai_mai_n304_));
  OAI210     m0282(.A0(mai_mai_n165_), .A1(mai_mai_n143_), .B0(mai_mai_n304_), .Y(mai_mai_n305_));
  NO3        m0283(.A(mai_mai_n305_), .B(mai_mai_n300_), .C(mai_mai_n295_), .Y(mai_mai_n306_));
  NO2        m0284(.A(i_3_), .B(i_10_), .Y(mai_mai_n307_));
  NA3        m0285(.A(mai_mai_n307_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n308_));
  NO2        m0286(.A(i_2_), .B(mai_mai_n103_), .Y(mai_mai_n309_));
  NA2        m0287(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n310_));
  NO2        m0288(.A(mai_mai_n310_), .B(i_8_), .Y(mai_mai_n311_));
  NA2        m0289(.A(mai_mai_n311_), .B(mai_mai_n309_), .Y(mai_mai_n312_));
  AN2        m0290(.A(i_3_), .B(i_10_), .Y(mai_mai_n313_));
  NA4        m0291(.A(mai_mai_n313_), .B(mai_mai_n200_), .C(mai_mai_n177_), .D(mai_mai_n175_), .Y(mai_mai_n314_));
  NO2        m0292(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n315_));
  NO2        m0293(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n316_));
  OR2        m0294(.A(mai_mai_n312_), .B(mai_mai_n308_), .Y(mai_mai_n317_));
  OAI220     m0295(.A0(mai_mai_n317_), .A1(i_6_), .B0(mai_mai_n306_), .B1(mai_mai_n290_), .Y(mai_mai_n318_));
  NO4        m0296(.A(mai_mai_n318_), .B(mai_mai_n288_), .C(mai_mai_n217_), .D(mai_mai_n168_), .Y(mai_mai_n319_));
  NO3        m0297(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n320_));
  NO2        m0298(.A(mai_mai_n59_), .B(mai_mai_n86_), .Y(mai_mai_n321_));
  NA2        m0299(.A(mai_mai_n297_), .B(mai_mai_n321_), .Y(mai_mai_n322_));
  NO3        m0300(.A(i_6_), .B(mai_mai_n195_), .C(i_7_), .Y(mai_mai_n323_));
  NA2        m0301(.A(mai_mai_n323_), .B(mai_mai_n200_), .Y(mai_mai_n324_));
  AOI210     m0302(.A0(mai_mai_n324_), .A1(mai_mai_n322_), .B0(mai_mai_n170_), .Y(mai_mai_n325_));
  NO2        m0303(.A(i_2_), .B(i_3_), .Y(mai_mai_n326_));
  OR2        m0304(.A(i_0_), .B(i_5_), .Y(mai_mai_n327_));
  NA2        m0305(.A(mai_mai_n221_), .B(mai_mai_n327_), .Y(mai_mai_n328_));
  NA4        m0306(.A(mai_mai_n328_), .B(mai_mai_n238_), .C(mai_mai_n326_), .D(i_1_), .Y(mai_mai_n329_));
  NA3        m0307(.A(mai_mai_n297_), .B(mai_mai_n292_), .C(mai_mai_n114_), .Y(mai_mai_n330_));
  NAi21      m0308(.An(i_8_), .B(i_7_), .Y(mai_mai_n331_));
  NO2        m0309(.A(mai_mai_n331_), .B(i_6_), .Y(mai_mai_n332_));
  NO2        m0310(.A(mai_mai_n157_), .B(mai_mai_n47_), .Y(mai_mai_n333_));
  NA3        m0311(.A(mai_mai_n333_), .B(mai_mai_n332_), .C(mai_mai_n163_), .Y(mai_mai_n334_));
  NA3        m0312(.A(mai_mai_n334_), .B(mai_mai_n330_), .C(mai_mai_n329_), .Y(mai_mai_n335_));
  OAI210     m0313(.A0(mai_mai_n335_), .A1(mai_mai_n325_), .B0(i_4_), .Y(mai_mai_n336_));
  NO2        m0314(.A(i_12_), .B(i_10_), .Y(mai_mai_n337_));
  NOi21      m0315(.An(i_5_), .B(i_0_), .Y(mai_mai_n338_));
  NO3        m0316(.A(mai_mai_n310_), .B(mai_mai_n338_), .C(mai_mai_n128_), .Y(mai_mai_n339_));
  NA4        m0317(.A(mai_mai_n84_), .B(mai_mai_n36_), .C(mai_mai_n86_), .D(i_8_), .Y(mai_mai_n340_));
  NA2        m0318(.A(mai_mai_n339_), .B(mai_mai_n337_), .Y(mai_mai_n341_));
  NO2        m0319(.A(i_6_), .B(i_8_), .Y(mai_mai_n342_));
  NOi21      m0320(.An(i_0_), .B(i_2_), .Y(mai_mai_n343_));
  AN2        m0321(.A(mai_mai_n343_), .B(mai_mai_n342_), .Y(mai_mai_n344_));
  NO2        m0322(.A(i_1_), .B(i_7_), .Y(mai_mai_n345_));
  AO220      m0323(.A0(mai_mai_n345_), .A1(mai_mai_n344_), .B0(mai_mai_n332_), .B1(mai_mai_n239_), .Y(mai_mai_n346_));
  NA3        m0324(.A(mai_mai_n346_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n347_));
  NA3        m0325(.A(mai_mai_n347_), .B(mai_mai_n341_), .C(mai_mai_n336_), .Y(mai_mai_n348_));
  NO3        m0326(.A(mai_mai_n237_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n349_));
  NO3        m0327(.A(mai_mai_n331_), .B(i_2_), .C(i_1_), .Y(mai_mai_n350_));
  OAI210     m0328(.A0(mai_mai_n350_), .A1(mai_mai_n349_), .B0(i_6_), .Y(mai_mai_n351_));
  NA3        m0329(.A(mai_mai_n257_), .B(mai_mai_n309_), .C(mai_mai_n195_), .Y(mai_mai_n352_));
  AOI210     m0330(.A0(mai_mai_n352_), .A1(mai_mai_n351_), .B0(mai_mai_n328_), .Y(mai_mai_n353_));
  NOi21      m0331(.An(mai_mai_n153_), .B(mai_mai_n106_), .Y(mai_mai_n354_));
  NA2        m0332(.A(mai_mai_n353_), .B(i_3_), .Y(mai_mai_n355_));
  INV        m0333(.A(mai_mai_n84_), .Y(mai_mai_n356_));
  NO2        m0334(.A(mai_mai_n301_), .B(mai_mai_n81_), .Y(mai_mai_n357_));
  NA2        m0335(.A(mai_mai_n357_), .B(mai_mai_n132_), .Y(mai_mai_n358_));
  NO2        m0336(.A(mai_mai_n95_), .B(mai_mai_n195_), .Y(mai_mai_n359_));
  NA2        m0337(.A(mai_mai_n359_), .B(mai_mai_n63_), .Y(mai_mai_n360_));
  AOI210     m0338(.A0(mai_mai_n360_), .A1(mai_mai_n358_), .B0(mai_mai_n356_), .Y(mai_mai_n361_));
  NO2        m0339(.A(mai_mai_n195_), .B(i_9_), .Y(mai_mai_n362_));
  NA3        m0340(.A(mai_mai_n362_), .B(mai_mai_n208_), .C(mai_mai_n157_), .Y(mai_mai_n363_));
  NO2        m0341(.A(mai_mai_n361_), .B(mai_mai_n300_), .Y(mai_mai_n364_));
  AOI210     m0342(.A0(mai_mai_n364_), .A1(mai_mai_n355_), .B0(mai_mai_n162_), .Y(mai_mai_n365_));
  AOI210     m0343(.A0(mai_mai_n348_), .A1(mai_mai_n320_), .B0(mai_mai_n365_), .Y(mai_mai_n366_));
  NOi32      m0344(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n367_));
  INV        m0345(.A(mai_mai_n367_), .Y(mai_mai_n368_));
  NAi21      m0346(.An(i_0_), .B(i_6_), .Y(mai_mai_n369_));
  NAi21      m0347(.An(i_1_), .B(i_5_), .Y(mai_mai_n370_));
  NA2        m0348(.A(mai_mai_n370_), .B(mai_mai_n369_), .Y(mai_mai_n371_));
  NA2        m0349(.A(mai_mai_n371_), .B(mai_mai_n25_), .Y(mai_mai_n372_));
  OAI210     m0350(.A0(mai_mai_n372_), .A1(mai_mai_n159_), .B0(mai_mai_n251_), .Y(mai_mai_n373_));
  NAi41      m0351(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n374_));
  OAI220     m0352(.A0(mai_mai_n374_), .A1(mai_mai_n370_), .B0(mai_mai_n224_), .B1(mai_mai_n159_), .Y(mai_mai_n375_));
  AOI210     m0353(.A0(mai_mai_n374_), .A1(mai_mai_n159_), .B0(mai_mai_n157_), .Y(mai_mai_n376_));
  NOi32      m0354(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n377_));
  OR2        m0355(.A(mai_mai_n376_), .B(mai_mai_n375_), .Y(mai_mai_n378_));
  NO2        m0356(.A(i_1_), .B(mai_mai_n103_), .Y(mai_mai_n379_));
  NAi21      m0357(.An(i_3_), .B(i_4_), .Y(mai_mai_n380_));
  NO2        m0358(.A(mai_mai_n380_), .B(i_9_), .Y(mai_mai_n381_));
  AN2        m0359(.A(i_6_), .B(i_7_), .Y(mai_mai_n382_));
  OAI210     m0360(.A0(mai_mai_n382_), .A1(mai_mai_n379_), .B0(mai_mai_n381_), .Y(mai_mai_n383_));
  NA2        m0361(.A(i_2_), .B(i_7_), .Y(mai_mai_n384_));
  NO2        m0362(.A(mai_mai_n380_), .B(i_10_), .Y(mai_mai_n385_));
  NA3        m0363(.A(mai_mai_n385_), .B(mai_mai_n384_), .C(mai_mai_n249_), .Y(mai_mai_n386_));
  AOI210     m0364(.A0(mai_mai_n386_), .A1(mai_mai_n383_), .B0(mai_mai_n187_), .Y(mai_mai_n387_));
  AOI210     m0365(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n388_));
  OAI210     m0366(.A0(mai_mai_n388_), .A1(mai_mai_n190_), .B0(mai_mai_n385_), .Y(mai_mai_n389_));
  AOI220     m0367(.A0(mai_mai_n385_), .A1(mai_mai_n345_), .B0(mai_mai_n243_), .B1(mai_mai_n190_), .Y(mai_mai_n390_));
  AOI210     m0368(.A0(mai_mai_n390_), .A1(mai_mai_n389_), .B0(i_5_), .Y(mai_mai_n391_));
  NO4        m0369(.A(mai_mai_n391_), .B(mai_mai_n387_), .C(mai_mai_n378_), .D(mai_mai_n373_), .Y(mai_mai_n392_));
  NO2        m0370(.A(mai_mai_n392_), .B(mai_mai_n368_), .Y(mai_mai_n393_));
  NO2        m0371(.A(mai_mai_n59_), .B(mai_mai_n25_), .Y(mai_mai_n394_));
  AN2        m0372(.A(i_12_), .B(i_5_), .Y(mai_mai_n395_));
  NO2        m0373(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n396_));
  NA2        m0374(.A(mai_mai_n396_), .B(mai_mai_n395_), .Y(mai_mai_n397_));
  NO2        m0375(.A(i_11_), .B(i_6_), .Y(mai_mai_n398_));
  NA3        m0376(.A(mai_mai_n398_), .B(mai_mai_n333_), .C(mai_mai_n229_), .Y(mai_mai_n399_));
  NO2        m0377(.A(mai_mai_n399_), .B(mai_mai_n397_), .Y(mai_mai_n400_));
  NO2        m0378(.A(mai_mai_n247_), .B(i_5_), .Y(mai_mai_n401_));
  NO2        m0379(.A(i_5_), .B(i_10_), .Y(mai_mai_n402_));
  AOI220     m0380(.A0(mai_mai_n402_), .A1(mai_mai_n277_), .B0(mai_mai_n401_), .B1(mai_mai_n200_), .Y(mai_mai_n403_));
  NA2        m0381(.A(mai_mai_n144_), .B(mai_mai_n46_), .Y(mai_mai_n404_));
  NO2        m0382(.A(mai_mai_n404_), .B(mai_mai_n403_), .Y(mai_mai_n405_));
  OAI210     m0383(.A0(mai_mai_n405_), .A1(mai_mai_n400_), .B0(mai_mai_n394_), .Y(mai_mai_n406_));
  NO2        m0384(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n407_));
  NO2        m0385(.A(mai_mai_n150_), .B(mai_mai_n86_), .Y(mai_mai_n408_));
  OAI210     m0386(.A0(mai_mai_n408_), .A1(mai_mai_n400_), .B0(mai_mai_n407_), .Y(mai_mai_n409_));
  NO3        m0387(.A(mai_mai_n86_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n410_));
  NO2        m0388(.A(i_3_), .B(mai_mai_n103_), .Y(mai_mai_n411_));
  NA4        m0389(.A(mai_mai_n307_), .B(mai_mai_n93_), .C(mai_mai_n75_), .D(mai_mai_n55_), .Y(mai_mai_n412_));
  NO2        m0390(.A(i_11_), .B(i_12_), .Y(mai_mai_n413_));
  NA2        m0391(.A(mai_mai_n413_), .B(mai_mai_n36_), .Y(mai_mai_n414_));
  NO2        m0392(.A(mai_mai_n412_), .B(mai_mai_n414_), .Y(mai_mai_n415_));
  NA2        m0393(.A(mai_mai_n402_), .B(mai_mai_n241_), .Y(mai_mai_n416_));
  NA3        m0394(.A(mai_mai_n114_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n417_));
  NO2        m0395(.A(mai_mai_n417_), .B(mai_mai_n224_), .Y(mai_mai_n418_));
  NAi21      m0396(.An(i_13_), .B(i_0_), .Y(mai_mai_n419_));
  NO2        m0397(.A(mai_mai_n419_), .B(mai_mai_n244_), .Y(mai_mai_n420_));
  OAI210     m0398(.A0(mai_mai_n418_), .A1(mai_mai_n415_), .B0(mai_mai_n420_), .Y(mai_mai_n421_));
  NA3        m0399(.A(mai_mai_n421_), .B(mai_mai_n409_), .C(mai_mai_n406_), .Y(mai_mai_n422_));
  NA2        m0400(.A(mai_mai_n45_), .B(mai_mai_n229_), .Y(mai_mai_n423_));
  NO3        m0401(.A(i_1_), .B(i_12_), .C(mai_mai_n86_), .Y(mai_mai_n424_));
  NO2        m0402(.A(i_0_), .B(i_11_), .Y(mai_mai_n425_));
  INV        m0403(.A(i_5_), .Y(mai_mai_n426_));
  AN2        m0404(.A(i_1_), .B(i_6_), .Y(mai_mai_n427_));
  NOi21      m0405(.An(i_2_), .B(i_12_), .Y(mai_mai_n428_));
  NA2        m0406(.A(mai_mai_n428_), .B(mai_mai_n427_), .Y(mai_mai_n429_));
  NO2        m0407(.A(mai_mai_n429_), .B(mai_mai_n426_), .Y(mai_mai_n430_));
  NA2        m0408(.A(mai_mai_n142_), .B(i_9_), .Y(mai_mai_n431_));
  NO2        m0409(.A(mai_mai_n431_), .B(i_4_), .Y(mai_mai_n432_));
  NA2        m0410(.A(mai_mai_n430_), .B(mai_mai_n432_), .Y(mai_mai_n433_));
  NAi21      m0411(.An(i_9_), .B(i_4_), .Y(mai_mai_n434_));
  OR2        m0412(.A(i_13_), .B(i_10_), .Y(mai_mai_n435_));
  NO3        m0413(.A(mai_mai_n435_), .B(mai_mai_n117_), .C(mai_mai_n434_), .Y(mai_mai_n436_));
  OR2        m0414(.A(mai_mai_n219_), .B(mai_mai_n218_), .Y(mai_mai_n437_));
  NO2        m0415(.A(mai_mai_n103_), .B(mai_mai_n25_), .Y(mai_mai_n438_));
  NA2        m0416(.A(mai_mai_n289_), .B(mai_mai_n438_), .Y(mai_mai_n439_));
  NA2        m0417(.A(mai_mai_n282_), .B(mai_mai_n213_), .Y(mai_mai_n440_));
  OAI220     m0418(.A0(mai_mai_n440_), .A1(mai_mai_n437_), .B0(mai_mai_n439_), .B1(mai_mai_n354_), .Y(mai_mai_n441_));
  INV        m0419(.A(mai_mai_n441_), .Y(mai_mai_n442_));
  AOI210     m0420(.A0(mai_mai_n442_), .A1(mai_mai_n433_), .B0(mai_mai_n26_), .Y(mai_mai_n443_));
  NA2        m0421(.A(mai_mai_n330_), .B(mai_mai_n329_), .Y(mai_mai_n444_));
  AOI220     m0422(.A0(mai_mai_n303_), .A1(mai_mai_n293_), .B0(mai_mai_n297_), .B1(mai_mai_n321_), .Y(mai_mai_n445_));
  NO2        m0423(.A(mai_mai_n445_), .B(mai_mai_n170_), .Y(mai_mai_n446_));
  NO2        m0424(.A(mai_mai_n184_), .B(mai_mai_n86_), .Y(mai_mai_n447_));
  AOI220     m0425(.A0(mai_mai_n447_), .A1(mai_mai_n302_), .B0(mai_mai_n284_), .B1(mai_mai_n213_), .Y(mai_mai_n448_));
  NO2        m0426(.A(mai_mai_n448_), .B(mai_mai_n291_), .Y(mai_mai_n449_));
  NO3        m0427(.A(mai_mai_n449_), .B(mai_mai_n446_), .C(mai_mai_n444_), .Y(mai_mai_n450_));
  NA2        m0428(.A(mai_mai_n198_), .B(mai_mai_n98_), .Y(mai_mai_n451_));
  NA3        m0429(.A(mai_mai_n333_), .B(mai_mai_n163_), .C(mai_mai_n86_), .Y(mai_mai_n452_));
  AOI210     m0430(.A0(mai_mai_n452_), .A1(mai_mai_n451_), .B0(mai_mai_n331_), .Y(mai_mai_n453_));
  NA2        m0431(.A(mai_mai_n195_), .B(i_10_), .Y(mai_mai_n454_));
  NA3        m0432(.A(mai_mai_n263_), .B(mai_mai_n64_), .C(i_2_), .Y(mai_mai_n455_));
  NA2        m0433(.A(mai_mai_n303_), .B(mai_mai_n239_), .Y(mai_mai_n456_));
  OAI220     m0434(.A0(mai_mai_n456_), .A1(mai_mai_n184_), .B0(mai_mai_n455_), .B1(mai_mai_n454_), .Y(mai_mai_n457_));
  NO2        m0435(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n458_));
  NA3        m0436(.A(mai_mai_n345_), .B(mai_mai_n344_), .C(mai_mai_n458_), .Y(mai_mai_n459_));
  NA2        m0437(.A(mai_mai_n323_), .B(mai_mai_n328_), .Y(mai_mai_n460_));
  OAI210     m0438(.A0(mai_mai_n460_), .A1(mai_mai_n191_), .B0(mai_mai_n459_), .Y(mai_mai_n461_));
  NO3        m0439(.A(mai_mai_n461_), .B(mai_mai_n457_), .C(mai_mai_n453_), .Y(mai_mai_n462_));
  AOI210     m0440(.A0(mai_mai_n462_), .A1(mai_mai_n450_), .B0(mai_mai_n278_), .Y(mai_mai_n463_));
  NO4        m0441(.A(mai_mai_n463_), .B(mai_mai_n443_), .C(mai_mai_n422_), .D(mai_mai_n393_), .Y(mai_mai_n464_));
  NO2        m0442(.A(mai_mai_n63_), .B(i_4_), .Y(mai_mai_n465_));
  NO2        m0443(.A(mai_mai_n73_), .B(i_13_), .Y(mai_mai_n466_));
  NO2        m0444(.A(i_10_), .B(i_9_), .Y(mai_mai_n467_));
  NAi21      m0445(.An(i_12_), .B(i_8_), .Y(mai_mai_n468_));
  NO2        m0446(.A(mai_mai_n468_), .B(i_3_), .Y(mai_mai_n469_));
  NO2        m0447(.A(mai_mai_n47_), .B(i_4_), .Y(mai_mai_n470_));
  NA2        m0448(.A(mai_mai_n470_), .B(mai_mai_n106_), .Y(mai_mai_n471_));
  NO2        m0449(.A(mai_mai_n471_), .B(mai_mai_n207_), .Y(mai_mai_n472_));
  NA2        m0450(.A(mai_mai_n316_), .B(i_0_), .Y(mai_mai_n473_));
  NO3        m0451(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n474_));
  NA2        m0452(.A(mai_mai_n275_), .B(mai_mai_n99_), .Y(mai_mai_n475_));
  NA2        m0453(.A(mai_mai_n475_), .B(mai_mai_n474_), .Y(mai_mai_n476_));
  NA2        m0454(.A(i_8_), .B(i_9_), .Y(mai_mai_n477_));
  AOI210     m0455(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n478_));
  OR2        m0456(.A(mai_mai_n478_), .B(mai_mai_n477_), .Y(mai_mai_n479_));
  NA2        m0457(.A(mai_mai_n289_), .B(mai_mai_n208_), .Y(mai_mai_n480_));
  NO2        m0458(.A(mai_mai_n480_), .B(mai_mai_n479_), .Y(mai_mai_n481_));
  NA2        m0459(.A(mai_mai_n256_), .B(mai_mai_n315_), .Y(mai_mai_n482_));
  NO3        m0460(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n483_));
  AOI210     m0461(.A0(mai_mai_n262_), .A1(mai_mai_n190_), .B0(mai_mai_n483_), .Y(mai_mai_n484_));
  NO2        m0462(.A(mai_mai_n484_), .B(mai_mai_n482_), .Y(mai_mai_n485_));
  NO3        m0463(.A(mai_mai_n485_), .B(mai_mai_n481_), .C(mai_mai_n472_), .Y(mai_mai_n486_));
  OR2        m0464(.A(mai_mai_n301_), .B(mai_mai_n210_), .Y(mai_mai_n487_));
  OA210      m0465(.A0(mai_mai_n363_), .A1(mai_mai_n103_), .B0(mai_mai_n304_), .Y(mai_mai_n488_));
  OA220      m0466(.A0(mai_mai_n488_), .A1(mai_mai_n162_), .B0(mai_mai_n487_), .B1(mai_mai_n236_), .Y(mai_mai_n489_));
  NA2        m0467(.A(mai_mai_n98_), .B(i_13_), .Y(mai_mai_n490_));
  NA2        m0468(.A(mai_mai_n447_), .B(mai_mai_n394_), .Y(mai_mai_n491_));
  NO2        m0469(.A(i_2_), .B(i_13_), .Y(mai_mai_n492_));
  NA3        m0470(.A(mai_mai_n492_), .B(mai_mai_n161_), .C(mai_mai_n101_), .Y(mai_mai_n493_));
  OAI220     m0471(.A0(mai_mai_n493_), .A1(mai_mai_n241_), .B0(mai_mai_n491_), .B1(mai_mai_n490_), .Y(mai_mai_n494_));
  NO3        m0472(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n495_));
  NO2        m0473(.A(i_6_), .B(i_7_), .Y(mai_mai_n496_));
  NA2        m0474(.A(mai_mai_n496_), .B(mai_mai_n495_), .Y(mai_mai_n497_));
  NO2        m0475(.A(i_11_), .B(i_1_), .Y(mai_mai_n498_));
  NO2        m0476(.A(mai_mai_n73_), .B(i_3_), .Y(mai_mai_n499_));
  OR2        m0477(.A(i_11_), .B(i_8_), .Y(mai_mai_n500_));
  NOi21      m0478(.An(i_2_), .B(i_7_), .Y(mai_mai_n501_));
  NAi31      m0479(.An(mai_mai_n500_), .B(mai_mai_n501_), .C(mai_mai_n499_), .Y(mai_mai_n502_));
  NO2        m0480(.A(mai_mai_n435_), .B(i_6_), .Y(mai_mai_n503_));
  NA3        m0481(.A(mai_mai_n503_), .B(mai_mai_n465_), .C(mai_mai_n75_), .Y(mai_mai_n504_));
  NO2        m0482(.A(mai_mai_n504_), .B(mai_mai_n502_), .Y(mai_mai_n505_));
  NO2        m0483(.A(i_3_), .B(mai_mai_n195_), .Y(mai_mai_n506_));
  NO2        m0484(.A(i_6_), .B(i_10_), .Y(mai_mai_n507_));
  NA4        m0485(.A(mai_mai_n507_), .B(mai_mai_n320_), .C(mai_mai_n506_), .D(mai_mai_n241_), .Y(mai_mai_n508_));
  NO2        m0486(.A(mai_mai_n508_), .B(mai_mai_n155_), .Y(mai_mai_n509_));
  NA3        m0487(.A(mai_mai_n250_), .B(mai_mai_n172_), .C(mai_mai_n132_), .Y(mai_mai_n510_));
  NA2        m0488(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n511_));
  NO2        m0489(.A(mai_mai_n157_), .B(i_3_), .Y(mai_mai_n512_));
  NAi31      m0490(.An(mai_mai_n511_), .B(mai_mai_n512_), .C(mai_mai_n230_), .Y(mai_mai_n513_));
  NA3        m0491(.A(mai_mai_n407_), .B(mai_mai_n180_), .C(mai_mai_n149_), .Y(mai_mai_n514_));
  NA3        m0492(.A(mai_mai_n514_), .B(mai_mai_n513_), .C(mai_mai_n510_), .Y(mai_mai_n515_));
  NO4        m0493(.A(mai_mai_n515_), .B(mai_mai_n509_), .C(mai_mai_n505_), .D(mai_mai_n494_), .Y(mai_mai_n516_));
  NA2        m0494(.A(mai_mai_n474_), .B(mai_mai_n395_), .Y(mai_mai_n517_));
  NA2        m0495(.A(mai_mai_n483_), .B(mai_mai_n402_), .Y(mai_mai_n518_));
  NO2        m0496(.A(mai_mai_n518_), .B(mai_mai_n228_), .Y(mai_mai_n519_));
  NAi21      m0497(.An(mai_mai_n219_), .B(mai_mai_n413_), .Y(mai_mai_n520_));
  NO2        m0498(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n521_));
  NO2        m0499(.A(i_0_), .B(mai_mai_n86_), .Y(mai_mai_n522_));
  NA3        m0500(.A(mai_mai_n522_), .B(mai_mai_n521_), .C(mai_mai_n142_), .Y(mai_mai_n523_));
  OR3        m0501(.A(mai_mai_n310_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n524_));
  NO2        m0502(.A(mai_mai_n524_), .B(mai_mai_n523_), .Y(mai_mai_n525_));
  NA2        m0503(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n526_));
  NA2        m0504(.A(mai_mai_n320_), .B(mai_mai_n243_), .Y(mai_mai_n527_));
  OAI220     m0505(.A0(mai_mai_n527_), .A1(mai_mai_n455_), .B0(mai_mai_n526_), .B1(mai_mai_n490_), .Y(mai_mai_n528_));
  NA4        m0506(.A(mai_mai_n313_), .B(mai_mai_n227_), .C(mai_mai_n73_), .D(mai_mai_n241_), .Y(mai_mai_n529_));
  NO2        m0507(.A(mai_mai_n529_), .B(mai_mai_n497_), .Y(mai_mai_n530_));
  NO4        m0508(.A(mai_mai_n530_), .B(mai_mai_n528_), .C(mai_mai_n525_), .D(mai_mai_n519_), .Y(mai_mai_n531_));
  NA4        m0509(.A(mai_mai_n531_), .B(mai_mai_n516_), .C(mai_mai_n489_), .D(mai_mai_n486_), .Y(mai_mai_n532_));
  NA3        m0510(.A(mai_mai_n313_), .B(mai_mai_n177_), .C(mai_mai_n175_), .Y(mai_mai_n533_));
  OAI210     m0511(.A0(mai_mai_n308_), .A1(mai_mai_n182_), .B0(mai_mai_n533_), .Y(mai_mai_n534_));
  AN2        m0512(.A(mai_mai_n293_), .B(mai_mai_n238_), .Y(mai_mai_n535_));
  NA2        m0513(.A(mai_mai_n535_), .B(mai_mai_n534_), .Y(mai_mai_n536_));
  NA2        m0514(.A(mai_mai_n122_), .B(mai_mai_n113_), .Y(mai_mai_n537_));
  AN2        m0515(.A(mai_mai_n537_), .B(mai_mai_n474_), .Y(mai_mai_n538_));
  NA2        m0516(.A(mai_mai_n320_), .B(mai_mai_n164_), .Y(mai_mai_n539_));
  OAI210     m0517(.A0(mai_mai_n539_), .A1(mai_mai_n236_), .B0(mai_mai_n314_), .Y(mai_mai_n540_));
  AOI220     m0518(.A0(mai_mai_n540_), .A1(mai_mai_n332_), .B0(mai_mai_n538_), .B1(mai_mai_n316_), .Y(mai_mai_n541_));
  NA2        m0519(.A(mai_mai_n395_), .B(mai_mai_n229_), .Y(mai_mai_n542_));
  NA2        m0520(.A(mai_mai_n367_), .B(mai_mai_n73_), .Y(mai_mai_n543_));
  NA2        m0521(.A(mai_mai_n382_), .B(mai_mai_n377_), .Y(mai_mai_n544_));
  AO210      m0522(.A0(mai_mai_n543_), .A1(mai_mai_n542_), .B0(mai_mai_n544_), .Y(mai_mai_n545_));
  NO2        m0523(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n546_));
  AOI210     m0524(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n436_), .Y(mai_mai_n547_));
  NA2        m0525(.A(mai_mai_n547_), .B(mai_mai_n545_), .Y(mai_mai_n548_));
  INV        m0526(.A(mai_mai_n548_), .Y(mai_mai_n549_));
  NO2        m0527(.A(i_7_), .B(mai_mai_n201_), .Y(mai_mai_n550_));
  OR2        m0528(.A(mai_mai_n184_), .B(i_4_), .Y(mai_mai_n551_));
  NO2        m0529(.A(mai_mai_n551_), .B(mai_mai_n86_), .Y(mai_mai_n552_));
  NA2        m0530(.A(mai_mai_n552_), .B(mai_mai_n550_), .Y(mai_mai_n553_));
  NA4        m0531(.A(mai_mai_n553_), .B(mai_mai_n549_), .C(mai_mai_n541_), .D(mai_mai_n536_), .Y(mai_mai_n554_));
  NA2        m0532(.A(mai_mai_n401_), .B(mai_mai_n302_), .Y(mai_mai_n555_));
  OAI210     m0533(.A0(mai_mai_n397_), .A1(mai_mai_n169_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  NO2        m0534(.A(i_12_), .B(mai_mai_n195_), .Y(mai_mai_n557_));
  NA2        m0535(.A(mai_mai_n557_), .B(mai_mai_n229_), .Y(mai_mai_n558_));
  NO2        m0536(.A(mai_mai_n1080_), .B(mai_mai_n558_), .Y(mai_mai_n559_));
  NOi31      m0537(.An(mai_mai_n323_), .B(mai_mai_n435_), .C(mai_mai_n38_), .Y(mai_mai_n560_));
  OAI210     m0538(.A0(mai_mai_n560_), .A1(mai_mai_n559_), .B0(mai_mai_n556_), .Y(mai_mai_n561_));
  NO2        m0539(.A(i_8_), .B(i_7_), .Y(mai_mai_n562_));
  OAI210     m0540(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n563_));
  NA2        m0541(.A(mai_mai_n563_), .B(mai_mai_n227_), .Y(mai_mai_n564_));
  AOI220     m0542(.A0(mai_mai_n333_), .A1(mai_mai_n40_), .B0(mai_mai_n239_), .B1(mai_mai_n209_), .Y(mai_mai_n565_));
  OAI220     m0543(.A0(mai_mai_n565_), .A1(mai_mai_n551_), .B0(mai_mai_n564_), .B1(mai_mai_n247_), .Y(mai_mai_n566_));
  NA2        m0544(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n567_));
  NO2        m0545(.A(mai_mai_n567_), .B(i_6_), .Y(mai_mai_n568_));
  NA3        m0546(.A(mai_mai_n568_), .B(mai_mai_n566_), .C(mai_mai_n562_), .Y(mai_mai_n569_));
  AOI220     m0547(.A0(mai_mai_n447_), .A1(mai_mai_n333_), .B0(mai_mai_n252_), .B1(mai_mai_n249_), .Y(mai_mai_n570_));
  OAI220     m0548(.A0(mai_mai_n570_), .A1(mai_mai_n271_), .B0(mai_mai_n490_), .B1(mai_mai_n133_), .Y(mai_mai_n571_));
  NA2        m0549(.A(mai_mai_n571_), .B(mai_mai_n274_), .Y(mai_mai_n572_));
  NOi31      m0550(.An(mai_mai_n297_), .B(mai_mai_n308_), .C(mai_mai_n182_), .Y(mai_mai_n573_));
  NA3        m0551(.A(mai_mai_n313_), .B(mai_mai_n175_), .C(mai_mai_n98_), .Y(mai_mai_n574_));
  NO2        m0552(.A(mai_mai_n225_), .B(mai_mai_n45_), .Y(mai_mai_n575_));
  NO2        m0553(.A(mai_mai_n157_), .B(i_5_), .Y(mai_mai_n576_));
  NA3        m0554(.A(mai_mai_n576_), .B(mai_mai_n423_), .C(mai_mai_n326_), .Y(mai_mai_n577_));
  OAI210     m0555(.A0(mai_mai_n577_), .A1(mai_mai_n575_), .B0(mai_mai_n574_), .Y(mai_mai_n578_));
  OAI210     m0556(.A0(mai_mai_n578_), .A1(mai_mai_n573_), .B0(mai_mai_n483_), .Y(mai_mai_n579_));
  NA4        m0557(.A(mai_mai_n579_), .B(mai_mai_n572_), .C(mai_mai_n569_), .D(mai_mai_n561_), .Y(mai_mai_n580_));
  NA3        m0558(.A(mai_mai_n221_), .B(mai_mai_n71_), .C(mai_mai_n45_), .Y(mai_mai_n581_));
  NA2        m0559(.A(mai_mai_n289_), .B(mai_mai_n84_), .Y(mai_mai_n582_));
  AOI210     m0560(.A0(mai_mai_n581_), .A1(mai_mai_n358_), .B0(mai_mai_n582_), .Y(mai_mai_n583_));
  NA2        m0561(.A(mai_mai_n303_), .B(mai_mai_n293_), .Y(mai_mai_n584_));
  NO2        m0562(.A(mai_mai_n584_), .B(mai_mai_n174_), .Y(mai_mai_n585_));
  NA2        m0563(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n586_));
  NA2        m0564(.A(mai_mai_n467_), .B(mai_mai_n225_), .Y(mai_mai_n587_));
  NO2        m0565(.A(mai_mai_n586_), .B(mai_mai_n587_), .Y(mai_mai_n588_));
  AOI210     m0566(.A0(i_6_), .A1(mai_mai_n47_), .B0(mai_mai_n379_), .Y(mai_mai_n589_));
  NA2        m0567(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n590_));
  NA3        m0568(.A(mai_mai_n557_), .B(mai_mai_n280_), .C(mai_mai_n590_), .Y(mai_mai_n591_));
  NO2        m0569(.A(mai_mai_n589_), .B(mai_mai_n591_), .Y(mai_mai_n592_));
  NO4        m0570(.A(mai_mai_n592_), .B(mai_mai_n588_), .C(mai_mai_n585_), .D(mai_mai_n583_), .Y(mai_mai_n593_));
  NO4        m0571(.A(mai_mai_n257_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n594_));
  NO3        m0572(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n595_));
  NO2        m0573(.A(mai_mai_n237_), .B(mai_mai_n36_), .Y(mai_mai_n596_));
  AN2        m0574(.A(mai_mai_n596_), .B(mai_mai_n595_), .Y(mai_mai_n597_));
  OA210      m0575(.A0(mai_mai_n597_), .A1(mai_mai_n594_), .B0(mai_mai_n367_), .Y(mai_mai_n598_));
  NO2        m0576(.A(mai_mai_n435_), .B(i_1_), .Y(mai_mai_n599_));
  NOi31      m0577(.An(mai_mai_n599_), .B(mai_mai_n475_), .C(mai_mai_n73_), .Y(mai_mai_n600_));
  AN4        m0578(.A(mai_mai_n600_), .B(mai_mai_n432_), .C(mai_mai_n521_), .D(i_2_), .Y(mai_mai_n601_));
  NO2        m0579(.A(mai_mai_n445_), .B(mai_mai_n178_), .Y(mai_mai_n602_));
  NO3        m0580(.A(mai_mai_n602_), .B(mai_mai_n601_), .C(mai_mai_n598_), .Y(mai_mai_n603_));
  NOi21      m0581(.An(i_10_), .B(i_6_), .Y(mai_mai_n604_));
  NO2        m0582(.A(mai_mai_n86_), .B(mai_mai_n25_), .Y(mai_mai_n605_));
  NO2        m0583(.A(mai_mai_n116_), .B(mai_mai_n23_), .Y(mai_mai_n606_));
  NA2        m0584(.A(mai_mai_n323_), .B(mai_mai_n164_), .Y(mai_mai_n607_));
  AOI220     m0585(.A0(mai_mai_n607_), .A1(mai_mai_n456_), .B0(mai_mai_n185_), .B1(mai_mai_n183_), .Y(mai_mai_n608_));
  NOi31      m0586(.An(mai_mai_n146_), .B(i_1_), .C(mai_mai_n340_), .Y(mai_mai_n609_));
  NO2        m0587(.A(mai_mai_n609_), .B(mai_mai_n608_), .Y(mai_mai_n610_));
  NO2        m0588(.A(mai_mai_n543_), .B(mai_mai_n390_), .Y(mai_mai_n611_));
  INV        m0589(.A(mai_mai_n326_), .Y(mai_mai_n612_));
  NO2        m0590(.A(i_12_), .B(mai_mai_n86_), .Y(mai_mai_n613_));
  NA2        m0591(.A(mai_mai_n175_), .B(i_0_), .Y(mai_mai_n614_));
  NO3        m0592(.A(mai_mai_n614_), .B(mai_mai_n351_), .C(mai_mai_n308_), .Y(mai_mai_n615_));
  OR2        m0593(.A(i_2_), .B(i_5_), .Y(mai_mai_n616_));
  OR2        m0594(.A(mai_mai_n616_), .B(mai_mai_n427_), .Y(mai_mai_n617_));
  AOI210     m0595(.A0(mai_mai_n384_), .A1(mai_mai_n249_), .B0(mai_mai_n200_), .Y(mai_mai_n618_));
  AOI210     m0596(.A0(mai_mai_n618_), .A1(mai_mai_n617_), .B0(mai_mai_n520_), .Y(mai_mai_n619_));
  NO3        m0597(.A(mai_mai_n619_), .B(mai_mai_n615_), .C(mai_mai_n611_), .Y(mai_mai_n620_));
  NA4        m0598(.A(mai_mai_n620_), .B(mai_mai_n610_), .C(mai_mai_n603_), .D(mai_mai_n593_), .Y(mai_mai_n621_));
  NO4        m0599(.A(mai_mai_n621_), .B(mai_mai_n580_), .C(mai_mai_n554_), .D(mai_mai_n532_), .Y(mai_mai_n622_));
  NA4        m0600(.A(mai_mai_n622_), .B(mai_mai_n464_), .C(mai_mai_n366_), .D(mai_mai_n319_), .Y(mai7));
  NO2        m0601(.A(mai_mai_n95_), .B(mai_mai_n55_), .Y(mai_mai_n624_));
  NO2        m0602(.A(mai_mai_n110_), .B(mai_mai_n92_), .Y(mai_mai_n625_));
  NA2        m0603(.A(mai_mai_n396_), .B(mai_mai_n625_), .Y(mai_mai_n626_));
  NA2        m0604(.A(mai_mai_n507_), .B(mai_mai_n84_), .Y(mai_mai_n627_));
  NA2        m0605(.A(i_11_), .B(mai_mai_n195_), .Y(mai_mai_n628_));
  INV        m0606(.A(mai_mai_n626_), .Y(mai_mai_n629_));
  NA3        m0607(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n630_));
  NO2        m0608(.A(mai_mai_n241_), .B(i_4_), .Y(mai_mai_n631_));
  NA2        m0609(.A(mai_mai_n631_), .B(i_8_), .Y(mai_mai_n632_));
  NO2        m0610(.A(mai_mai_n107_), .B(mai_mai_n630_), .Y(mai_mai_n633_));
  NA2        m0611(.A(i_2_), .B(mai_mai_n86_), .Y(mai_mai_n634_));
  OAI210     m0612(.A0(mai_mai_n89_), .A1(mai_mai_n205_), .B0(mai_mai_n206_), .Y(mai_mai_n635_));
  NO2        m0613(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n636_));
  NA2        m0614(.A(i_4_), .B(i_8_), .Y(mai_mai_n637_));
  AOI210     m0615(.A0(mai_mai_n637_), .A1(mai_mai_n313_), .B0(mai_mai_n636_), .Y(mai_mai_n638_));
  OAI220     m0616(.A0(mai_mai_n638_), .A1(mai_mai_n634_), .B0(mai_mai_n635_), .B1(i_13_), .Y(mai_mai_n639_));
  NO4        m0617(.A(mai_mai_n639_), .B(mai_mai_n633_), .C(mai_mai_n629_), .D(mai_mai_n624_), .Y(mai_mai_n640_));
  AOI210     m0618(.A0(mai_mai_n128_), .A1(mai_mai_n62_), .B0(i_10_), .Y(mai_mai_n641_));
  AOI210     m0619(.A0(mai_mai_n641_), .A1(mai_mai_n241_), .B0(mai_mai_n161_), .Y(mai_mai_n642_));
  OR2        m0620(.A(i_6_), .B(i_10_), .Y(mai_mai_n643_));
  NO2        m0621(.A(mai_mai_n643_), .B(mai_mai_n23_), .Y(mai_mai_n644_));
  OR3        m0622(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n645_));
  NO3        m0623(.A(mai_mai_n645_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n646_));
  INV        m0624(.A(mai_mai_n202_), .Y(mai_mai_n647_));
  NO2        m0625(.A(mai_mai_n646_), .B(mai_mai_n644_), .Y(mai_mai_n648_));
  OA220      m0626(.A0(mai_mai_n648_), .A1(mai_mai_n612_), .B0(mai_mai_n642_), .B1(mai_mai_n276_), .Y(mai_mai_n649_));
  AOI210     m0627(.A0(mai_mai_n649_), .A1(mai_mai_n640_), .B0(mai_mai_n63_), .Y(mai_mai_n650_));
  NOi21      m0628(.An(i_11_), .B(i_7_), .Y(mai_mai_n651_));
  AO210      m0629(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n652_));
  NO2        m0630(.A(mai_mai_n652_), .B(mai_mai_n651_), .Y(mai_mai_n653_));
  NA2        m0631(.A(mai_mai_n653_), .B(mai_mai_n209_), .Y(mai_mai_n654_));
  NA3        m0632(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n655_));
  NAi31      m0633(.An(mai_mai_n655_), .B(mai_mai_n218_), .C(i_11_), .Y(mai_mai_n656_));
  AOI210     m0634(.A0(mai_mai_n656_), .A1(mai_mai_n654_), .B0(mai_mai_n63_), .Y(mai_mai_n657_));
  NA2        m0635(.A(mai_mai_n88_), .B(mai_mai_n63_), .Y(mai_mai_n658_));
  AO210      m0636(.A0(mai_mai_n658_), .A1(mai_mai_n390_), .B0(mai_mai_n41_), .Y(mai_mai_n659_));
  NA2        m0637(.A(mai_mai_n230_), .B(mai_mai_n63_), .Y(mai_mai_n660_));
  NO2        m0638(.A(mai_mai_n63_), .B(i_9_), .Y(mai_mai_n661_));
  NO2        m0639(.A(i_1_), .B(i_12_), .Y(mai_mai_n662_));
  NA2        m0640(.A(mai_mai_n660_), .B(mai_mai_n659_), .Y(mai_mai_n663_));
  OAI210     m0641(.A0(mai_mai_n663_), .A1(mai_mai_n657_), .B0(i_6_), .Y(mai_mai_n664_));
  NO2        m0642(.A(mai_mai_n655_), .B(mai_mai_n110_), .Y(mai_mai_n665_));
  NA2        m0643(.A(mai_mai_n665_), .B(mai_mai_n613_), .Y(mai_mai_n666_));
  NO2        m0644(.A(mai_mai_n241_), .B(mai_mai_n86_), .Y(mai_mai_n667_));
  NO2        m0645(.A(mai_mai_n667_), .B(i_11_), .Y(mai_mai_n668_));
  NA2        m0646(.A(mai_mai_n666_), .B(mai_mai_n476_), .Y(mai_mai_n669_));
  NO4        m0647(.A(mai_mai_n218_), .B(mai_mai_n128_), .C(i_13_), .D(mai_mai_n86_), .Y(mai_mai_n670_));
  NA2        m0648(.A(mai_mai_n670_), .B(mai_mai_n661_), .Y(mai_mai_n671_));
  NA2        m0649(.A(mai_mai_n241_), .B(i_6_), .Y(mai_mai_n672_));
  NA2        m0650(.A(i_1_), .B(mai_mai_n266_), .Y(mai_mai_n673_));
  OAI210     m0651(.A0(mai_mai_n673_), .A1(mai_mai_n45_), .B0(mai_mai_n671_), .Y(mai_mai_n674_));
  NA3        m0652(.A(mai_mai_n562_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n675_));
  NA2        m0653(.A(mai_mai_n138_), .B(i_9_), .Y(mai_mai_n676_));
  NA3        m0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n677_));
  NO2        m0655(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n678_));
  NO2        m0656(.A(mai_mai_n676_), .B(mai_mai_n1078_), .Y(mai_mai_n679_));
  NA3        m0657(.A(mai_mai_n661_), .B(mai_mai_n326_), .C(i_6_), .Y(mai_mai_n680_));
  NO2        m0658(.A(mai_mai_n680_), .B(mai_mai_n23_), .Y(mai_mai_n681_));
  AOI210     m0659(.A0(mai_mai_n498_), .A1(mai_mai_n438_), .B0(mai_mai_n246_), .Y(mai_mai_n682_));
  NO2        m0660(.A(mai_mai_n682_), .B(mai_mai_n634_), .Y(mai_mai_n683_));
  NAi21      m0661(.An(mai_mai_n675_), .B(mai_mai_n94_), .Y(mai_mai_n684_));
  NA2        m0662(.A(mai_mai_n678_), .B(mai_mai_n275_), .Y(mai_mai_n685_));
  NO2        m0663(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n686_));
  NA2        m0664(.A(mai_mai_n686_), .B(mai_mai_n24_), .Y(mai_mai_n687_));
  OAI210     m0665(.A0(mai_mai_n687_), .A1(mai_mai_n685_), .B0(mai_mai_n684_), .Y(mai_mai_n688_));
  OR4        m0666(.A(mai_mai_n688_), .B(mai_mai_n683_), .C(mai_mai_n681_), .D(mai_mai_n679_), .Y(mai_mai_n689_));
  NO3        m0667(.A(mai_mai_n689_), .B(mai_mai_n674_), .C(mai_mai_n669_), .Y(mai_mai_n690_));
  NO2        m0668(.A(mai_mai_n241_), .B(mai_mai_n103_), .Y(mai_mai_n691_));
  NO2        m0669(.A(mai_mai_n691_), .B(mai_mai_n651_), .Y(mai_mai_n692_));
  NA2        m0670(.A(mai_mai_n692_), .B(i_1_), .Y(mai_mai_n693_));
  NO2        m0671(.A(mai_mai_n693_), .B(mai_mai_n645_), .Y(mai_mai_n694_));
  NO2        m0672(.A(mai_mai_n434_), .B(mai_mai_n86_), .Y(mai_mai_n695_));
  NA2        m0673(.A(mai_mai_n694_), .B(mai_mai_n47_), .Y(mai_mai_n696_));
  NO2        m0674(.A(mai_mai_n237_), .B(mai_mai_n45_), .Y(mai_mai_n697_));
  NO3        m0675(.A(mai_mai_n697_), .B(mai_mai_n316_), .C(mai_mai_n242_), .Y(mai_mai_n698_));
  NO2        m0676(.A(mai_mai_n117_), .B(mai_mai_n37_), .Y(mai_mai_n699_));
  NO2        m0677(.A(mai_mai_n699_), .B(i_6_), .Y(mai_mai_n700_));
  NO2        m0678(.A(mai_mai_n86_), .B(i_9_), .Y(mai_mai_n701_));
  NO2        m0679(.A(mai_mai_n701_), .B(mai_mai_n63_), .Y(mai_mai_n702_));
  NO2        m0680(.A(mai_mai_n702_), .B(mai_mai_n662_), .Y(mai_mai_n703_));
  NO4        m0681(.A(mai_mai_n703_), .B(mai_mai_n700_), .C(mai_mai_n698_), .D(i_4_), .Y(mai_mai_n704_));
  NA2        m0682(.A(i_1_), .B(i_3_), .Y(mai_mai_n705_));
  INV        m0683(.A(mai_mai_n704_), .Y(mai_mai_n706_));
  NA4        m0684(.A(mai_mai_n706_), .B(mai_mai_n696_), .C(mai_mai_n690_), .D(mai_mai_n664_), .Y(mai_mai_n707_));
  NO3        m0685(.A(mai_mai_n500_), .B(i_3_), .C(i_7_), .Y(mai_mai_n708_));
  NOi21      m0686(.An(mai_mai_n708_), .B(i_10_), .Y(mai_mai_n709_));
  OA210      m0687(.A0(mai_mai_n709_), .A1(mai_mai_n250_), .B0(mai_mai_n86_), .Y(mai_mai_n710_));
  NA3        m0688(.A(mai_mai_n507_), .B(mai_mai_n546_), .C(mai_mai_n47_), .Y(mai_mai_n711_));
  NA3        m0689(.A(mai_mai_n161_), .B(mai_mai_n84_), .C(mai_mai_n86_), .Y(mai_mai_n712_));
  NA2        m0690(.A(mai_mai_n712_), .B(mai_mai_n711_), .Y(mai_mai_n713_));
  OAI210     m0691(.A0(mai_mai_n713_), .A1(mai_mai_n710_), .B0(i_1_), .Y(mai_mai_n714_));
  AOI210     m0692(.A0(mai_mai_n275_), .A1(mai_mai_n99_), .B0(i_1_), .Y(mai_mai_n715_));
  NO2        m0693(.A(mai_mai_n380_), .B(i_2_), .Y(mai_mai_n716_));
  NA2        m0694(.A(mai_mai_n716_), .B(mai_mai_n715_), .Y(mai_mai_n717_));
  OAI210     m0695(.A0(mai_mai_n680_), .A1(mai_mai_n468_), .B0(mai_mai_n717_), .Y(mai_mai_n718_));
  INV        m0696(.A(mai_mai_n718_), .Y(mai_mai_n719_));
  AOI210     m0697(.A0(mai_mai_n719_), .A1(mai_mai_n714_), .B0(i_13_), .Y(mai_mai_n720_));
  OR2        m0698(.A(i_11_), .B(i_7_), .Y(mai_mai_n721_));
  NA3        m0699(.A(mai_mai_n721_), .B(mai_mai_n108_), .C(mai_mai_n138_), .Y(mai_mai_n722_));
  AOI220     m0700(.A0(mai_mai_n492_), .A1(mai_mai_n161_), .B0(mai_mai_n470_), .B1(mai_mai_n138_), .Y(mai_mai_n723_));
  OAI210     m0701(.A0(mai_mai_n723_), .A1(mai_mai_n45_), .B0(mai_mai_n722_), .Y(mai_mai_n724_));
  NO2        m0702(.A(mai_mai_n55_), .B(i_12_), .Y(mai_mai_n725_));
  INV        m0703(.A(mai_mai_n725_), .Y(mai_mai_n726_));
  NO2        m0704(.A(mai_mai_n501_), .B(mai_mai_n24_), .Y(mai_mai_n727_));
  AOI220     m0705(.A0(mai_mai_n727_), .A1(mai_mai_n695_), .B0(mai_mai_n250_), .B1(mai_mai_n131_), .Y(mai_mai_n728_));
  OAI220     m0706(.A0(mai_mai_n728_), .A1(mai_mai_n41_), .B0(mai_mai_n726_), .B1(mai_mai_n95_), .Y(mai_mai_n729_));
  AOI210     m0707(.A0(mai_mai_n724_), .A1(mai_mai_n342_), .B0(mai_mai_n729_), .Y(mai_mai_n730_));
  NA2        m0708(.A(mai_mai_n398_), .B(mai_mai_n678_), .Y(mai_mai_n731_));
  NO2        m0709(.A(mai_mai_n731_), .B(mai_mai_n247_), .Y(mai_mai_n732_));
  AOI210     m0710(.A0(mai_mai_n468_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n733_));
  NOi31      m0711(.An(mai_mai_n733_), .B(mai_mai_n627_), .C(mai_mai_n45_), .Y(mai_mai_n734_));
  NA2        m0712(.A(mai_mai_n127_), .B(i_13_), .Y(mai_mai_n735_));
  NO2        m0713(.A(mai_mai_n677_), .B(mai_mai_n116_), .Y(mai_mai_n736_));
  INV        m0714(.A(mai_mai_n736_), .Y(mai_mai_n737_));
  OAI220     m0715(.A0(mai_mai_n737_), .A1(mai_mai_n71_), .B0(mai_mai_n735_), .B1(mai_mai_n715_), .Y(mai_mai_n738_));
  NA2        m0716(.A(mai_mai_n26_), .B(mai_mai_n195_), .Y(mai_mai_n739_));
  INV        m0717(.A(i_7_), .Y(mai_mai_n740_));
  AOI220     m0718(.A0(mai_mai_n398_), .A1(mai_mai_n678_), .B0(mai_mai_n94_), .B1(mai_mai_n104_), .Y(mai_mai_n741_));
  NO2        m0719(.A(mai_mai_n741_), .B(mai_mai_n632_), .Y(mai_mai_n742_));
  NO4        m0720(.A(mai_mai_n742_), .B(mai_mai_n738_), .C(mai_mai_n734_), .D(mai_mai_n732_), .Y(mai_mai_n743_));
  OR2        m0721(.A(i_11_), .B(i_6_), .Y(mai_mai_n744_));
  NA3        m0722(.A(mai_mai_n631_), .B(mai_mai_n739_), .C(i_7_), .Y(mai_mai_n745_));
  AOI210     m0723(.A0(mai_mai_n745_), .A1(mai_mai_n737_), .B0(mai_mai_n744_), .Y(mai_mai_n746_));
  NA3        m0724(.A(mai_mai_n428_), .B(mai_mai_n636_), .C(mai_mai_n99_), .Y(mai_mai_n747_));
  NA2        m0725(.A(mai_mai_n668_), .B(i_13_), .Y(mai_mai_n748_));
  NA2        m0726(.A(mai_mai_n104_), .B(mai_mai_n739_), .Y(mai_mai_n749_));
  NAi21      m0727(.An(i_11_), .B(i_12_), .Y(mai_mai_n750_));
  NOi41      m0728(.An(mai_mai_n112_), .B(mai_mai_n750_), .C(i_13_), .D(mai_mai_n86_), .Y(mai_mai_n751_));
  NA2        m0729(.A(mai_mai_n751_), .B(mai_mai_n749_), .Y(mai_mai_n752_));
  NA3        m0730(.A(mai_mai_n752_), .B(mai_mai_n748_), .C(mai_mai_n747_), .Y(mai_mai_n753_));
  OAI210     m0731(.A0(mai_mai_n753_), .A1(mai_mai_n746_), .B0(mai_mai_n63_), .Y(mai_mai_n754_));
  NO2        m0732(.A(i_2_), .B(i_12_), .Y(mai_mai_n755_));
  NA2        m0733(.A(mai_mai_n379_), .B(mai_mai_n755_), .Y(mai_mai_n756_));
  NA2        m0734(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n757_));
  NO3        m0735(.A(mai_mai_n757_), .B(mai_mai_n396_), .C(mai_mai_n631_), .Y(mai_mai_n758_));
  OAI210     m0736(.A0(mai_mai_n758_), .A1(mai_mai_n381_), .B0(mai_mai_n379_), .Y(mai_mai_n759_));
  NO2        m0737(.A(mai_mai_n128_), .B(i_2_), .Y(mai_mai_n760_));
  NA2        m0738(.A(mai_mai_n759_), .B(mai_mai_n756_), .Y(mai_mai_n761_));
  NA3        m0739(.A(mai_mai_n761_), .B(mai_mai_n46_), .C(mai_mai_n229_), .Y(mai_mai_n762_));
  NA4        m0740(.A(mai_mai_n762_), .B(mai_mai_n754_), .C(mai_mai_n743_), .D(mai_mai_n730_), .Y(mai_mai_n763_));
  OR4        m0741(.A(mai_mai_n763_), .B(mai_mai_n720_), .C(mai_mai_n707_), .D(mai_mai_n650_), .Y(mai5));
  NA2        m0742(.A(mai_mai_n692_), .B(mai_mai_n277_), .Y(mai_mai_n765_));
  AN2        m0743(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n766_));
  NA3        m0744(.A(mai_mai_n766_), .B(mai_mai_n755_), .C(mai_mai_n110_), .Y(mai_mai_n767_));
  NO2        m0745(.A(mai_mai_n632_), .B(i_11_), .Y(mai_mai_n768_));
  NA2        m0746(.A(mai_mai_n89_), .B(mai_mai_n768_), .Y(mai_mai_n769_));
  NA3        m0747(.A(mai_mai_n769_), .B(mai_mai_n767_), .C(mai_mai_n765_), .Y(mai_mai_n770_));
  NO3        m0748(.A(i_11_), .B(mai_mai_n241_), .C(i_13_), .Y(mai_mai_n771_));
  NO2        m0749(.A(mai_mai_n124_), .B(mai_mai_n23_), .Y(mai_mai_n772_));
  NA2        m0750(.A(i_12_), .B(i_8_), .Y(mai_mai_n773_));
  OAI210     m0751(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n773_), .Y(mai_mai_n774_));
  INV        m0752(.A(mai_mai_n467_), .Y(mai_mai_n775_));
  AOI220     m0753(.A0(mai_mai_n326_), .A1(mai_mai_n606_), .B0(mai_mai_n774_), .B1(mai_mai_n772_), .Y(mai_mai_n776_));
  INV        m0754(.A(mai_mai_n776_), .Y(mai_mai_n777_));
  NO2        m0755(.A(mai_mai_n777_), .B(mai_mai_n770_), .Y(mai_mai_n778_));
  INV        m0756(.A(mai_mai_n172_), .Y(mai_mai_n779_));
  INV        m0757(.A(mai_mai_n250_), .Y(mai_mai_n780_));
  OAI210     m0758(.A0(mai_mai_n716_), .A1(mai_mai_n469_), .B0(mai_mai_n112_), .Y(mai_mai_n781_));
  AOI210     m0759(.A0(mai_mai_n781_), .A1(mai_mai_n780_), .B0(mai_mai_n779_), .Y(mai_mai_n782_));
  NO2        m0760(.A(mai_mai_n477_), .B(mai_mai_n26_), .Y(mai_mai_n783_));
  NO2        m0761(.A(mai_mai_n783_), .B(mai_mai_n438_), .Y(mai_mai_n784_));
  NA2        m0762(.A(mai_mai_n784_), .B(i_2_), .Y(mai_mai_n785_));
  INV        m0763(.A(mai_mai_n785_), .Y(mai_mai_n786_));
  AOI210     m0764(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n435_), .Y(mai_mai_n787_));
  AOI210     m0765(.A0(mai_mai_n787_), .A1(mai_mai_n786_), .B0(mai_mai_n782_), .Y(mai_mai_n788_));
  NO2        m0766(.A(mai_mai_n192_), .B(mai_mai_n125_), .Y(mai_mai_n789_));
  OAI210     m0767(.A0(mai_mai_n789_), .A1(mai_mai_n772_), .B0(i_2_), .Y(mai_mai_n790_));
  INV        m0768(.A(mai_mai_n173_), .Y(mai_mai_n791_));
  NO3        m0769(.A(mai_mai_n652_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n792_));
  AOI210     m0770(.A0(mai_mai_n791_), .A1(mai_mai_n89_), .B0(mai_mai_n792_), .Y(mai_mai_n793_));
  AOI210     m0771(.A0(mai_mai_n793_), .A1(mai_mai_n790_), .B0(mai_mai_n195_), .Y(mai_mai_n794_));
  OA210      m0772(.A0(mai_mai_n653_), .A1(mai_mai_n126_), .B0(i_13_), .Y(mai_mai_n795_));
  NA2        m0773(.A(mai_mai_n151_), .B(mai_mai_n628_), .Y(mai_mai_n796_));
  NO2        m0774(.A(mai_mai_n796_), .B(mai_mai_n384_), .Y(mai_mai_n797_));
  AOI210     m0775(.A0(mai_mai_n211_), .A1(mai_mai_n148_), .B0(mai_mai_n546_), .Y(mai_mai_n798_));
  OAI210     m0776(.A0(mai_mai_n798_), .A1(mai_mai_n230_), .B0(mai_mai_n438_), .Y(mai_mai_n799_));
  NO2        m0777(.A(mai_mai_n104_), .B(mai_mai_n45_), .Y(mai_mai_n800_));
  INV        m0778(.A(mai_mai_n309_), .Y(mai_mai_n801_));
  NA4        m0779(.A(mai_mai_n801_), .B(mai_mai_n313_), .C(mai_mai_n124_), .D(mai_mai_n43_), .Y(mai_mai_n802_));
  OAI210     m0780(.A0(mai_mai_n802_), .A1(mai_mai_n800_), .B0(mai_mai_n799_), .Y(mai_mai_n803_));
  NO4        m0781(.A(mai_mai_n803_), .B(mai_mai_n797_), .C(mai_mai_n795_), .D(mai_mai_n794_), .Y(mai_mai_n804_));
  NA2        m0782(.A(mai_mai_n606_), .B(mai_mai_n28_), .Y(mai_mai_n805_));
  NA2        m0783(.A(mai_mai_n771_), .B(mai_mai_n281_), .Y(mai_mai_n806_));
  NA2        m0784(.A(mai_mai_n806_), .B(mai_mai_n805_), .Y(mai_mai_n807_));
  NO2        m0785(.A(mai_mai_n62_), .B(i_12_), .Y(mai_mai_n808_));
  NO2        m0786(.A(mai_mai_n808_), .B(mai_mai_n126_), .Y(mai_mai_n809_));
  NO2        m0787(.A(mai_mai_n809_), .B(mai_mai_n628_), .Y(mai_mai_n810_));
  AOI220     m0788(.A0(mai_mai_n810_), .A1(mai_mai_n36_), .B0(mai_mai_n807_), .B1(mai_mai_n47_), .Y(mai_mai_n811_));
  NA4        m0789(.A(mai_mai_n811_), .B(mai_mai_n804_), .C(mai_mai_n788_), .D(mai_mai_n778_), .Y(mai6));
  NO3        m0790(.A(mai_mai_n261_), .B(mai_mai_n315_), .C(i_1_), .Y(mai_mai_n813_));
  NO2        m0791(.A(mai_mai_n187_), .B(mai_mai_n139_), .Y(mai_mai_n814_));
  OAI210     m0792(.A0(mai_mai_n814_), .A1(mai_mai_n813_), .B0(mai_mai_n760_), .Y(mai_mai_n815_));
  NO2        m0793(.A(mai_mai_n224_), .B(mai_mai_n511_), .Y(mai_mai_n816_));
  NO2        m0794(.A(i_11_), .B(i_9_), .Y(mai_mai_n817_));
  AO210      m0795(.A0(mai_mai_n1079_), .A1(mai_mai_n815_), .B0(i_12_), .Y(mai_mai_n818_));
  NA2        m0796(.A(mai_mai_n385_), .B(mai_mai_n345_), .Y(mai_mai_n819_));
  NA2        m0797(.A(mai_mai_n613_), .B(mai_mai_n63_), .Y(mai_mai_n820_));
  NA2        m0798(.A(mai_mai_n709_), .B(mai_mai_n71_), .Y(mai_mai_n821_));
  BUFFER     m0799(.A(mai_mai_n658_), .Y(mai_mai_n822_));
  NA4        m0800(.A(mai_mai_n822_), .B(mai_mai_n821_), .C(mai_mai_n820_), .D(mai_mai_n819_), .Y(mai_mai_n823_));
  INV        m0801(.A(mai_mai_n199_), .Y(mai_mai_n824_));
  AOI220     m0802(.A0(mai_mai_n824_), .A1(mai_mai_n817_), .B0(mai_mai_n823_), .B1(mai_mai_n73_), .Y(mai_mai_n825_));
  INV        m0803(.A(mai_mai_n337_), .Y(mai_mai_n826_));
  NA2        m0804(.A(mai_mai_n75_), .B(mai_mai_n131_), .Y(mai_mai_n827_));
  INV        m0805(.A(mai_mai_n124_), .Y(mai_mai_n828_));
  NA2        m0806(.A(mai_mai_n828_), .B(mai_mai_n47_), .Y(mai_mai_n829_));
  AOI210     m0807(.A0(mai_mai_n829_), .A1(mai_mai_n827_), .B0(mai_mai_n826_), .Y(mai_mai_n830_));
  NO2        m0808(.A(mai_mai_n257_), .B(i_9_), .Y(mai_mai_n831_));
  NA2        m0809(.A(mai_mai_n831_), .B(mai_mai_n808_), .Y(mai_mai_n832_));
  AOI210     m0810(.A0(mai_mai_n832_), .A1(mai_mai_n544_), .B0(mai_mai_n187_), .Y(mai_mai_n833_));
  NO2        m0811(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n834_));
  NA3        m0812(.A(mai_mai_n834_), .B(mai_mai_n496_), .C(mai_mai_n402_), .Y(mai_mai_n835_));
  NAi32      m0813(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n836_));
  AOI210     m0814(.A0(mai_mai_n744_), .A1(mai_mai_n87_), .B0(mai_mai_n836_), .Y(mai_mai_n837_));
  OAI210     m0815(.A0(mai_mai_n708_), .A1(mai_mai_n596_), .B0(mai_mai_n595_), .Y(mai_mai_n838_));
  NAi31      m0816(.An(mai_mai_n837_), .B(mai_mai_n838_), .C(mai_mai_n835_), .Y(mai_mai_n839_));
  OR3        m0817(.A(mai_mai_n839_), .B(mai_mai_n833_), .C(mai_mai_n830_), .Y(mai_mai_n840_));
  NO2        m0818(.A(mai_mai_n721_), .B(i_2_), .Y(mai_mai_n841_));
  NA2        m0819(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n842_));
  OAI210     m0820(.A0(mai_mai_n842_), .A1(mai_mai_n427_), .B0(mai_mai_n372_), .Y(mai_mai_n843_));
  NA2        m0821(.A(mai_mai_n843_), .B(mai_mai_n841_), .Y(mai_mai_n844_));
  AO220      m0822(.A0(mai_mai_n371_), .A1(mai_mai_n362_), .B0(mai_mai_n410_), .B1(mai_mai_n628_), .Y(mai_mai_n845_));
  NA3        m0823(.A(mai_mai_n845_), .B(mai_mai_n262_), .C(i_7_), .Y(mai_mai_n846_));
  BUFFER     m0824(.A(mai_mai_n653_), .Y(mai_mai_n847_));
  NA3        m0825(.A(mai_mai_n847_), .B(mai_mai_n147_), .C(mai_mai_n69_), .Y(mai_mai_n848_));
  AO210      m0826(.A0(mai_mai_n518_), .A1(mai_mai_n775_), .B0(mai_mai_n36_), .Y(mai_mai_n849_));
  NA4        m0827(.A(mai_mai_n849_), .B(mai_mai_n848_), .C(mai_mai_n846_), .D(mai_mai_n844_), .Y(mai_mai_n850_));
  OAI210     m0828(.A0(mai_mai_n667_), .A1(i_11_), .B0(mai_mai_n87_), .Y(mai_mai_n851_));
  AOI220     m0829(.A0(mai_mai_n851_), .A1(mai_mai_n595_), .B0(mai_mai_n816_), .B1(mai_mai_n740_), .Y(mai_mai_n852_));
  NA2        m0830(.A(mai_mai_n410_), .B(mai_mai_n70_), .Y(mai_mai_n853_));
  NA3        m0831(.A(mai_mai_n853_), .B(mai_mai_n852_), .C(mai_mai_n635_), .Y(mai_mai_n854_));
  AO210      m0832(.A0(mai_mai_n546_), .A1(mai_mai_n47_), .B0(mai_mai_n88_), .Y(mai_mai_n855_));
  NA3        m0833(.A(mai_mai_n855_), .B(mai_mai_n507_), .C(mai_mai_n221_), .Y(mai_mai_n856_));
  AOI210     m0834(.A0(mai_mai_n469_), .A1(mai_mai_n467_), .B0(mai_mai_n594_), .Y(mai_mai_n857_));
  NA2        m0835(.A(mai_mai_n113_), .B(mai_mai_n425_), .Y(mai_mai_n858_));
  NA2        m0836(.A(mai_mai_n249_), .B(mai_mai_n47_), .Y(mai_mai_n859_));
  NA2        m0837(.A(mai_mai_n859_), .B(mai_mai_n617_), .Y(mai_mai_n860_));
  NA3        m0838(.A(mai_mai_n860_), .B(mai_mai_n337_), .C(i_7_), .Y(mai_mai_n861_));
  NA4        m0839(.A(mai_mai_n861_), .B(mai_mai_n858_), .C(mai_mai_n857_), .D(mai_mai_n856_), .Y(mai_mai_n862_));
  NO4        m0840(.A(mai_mai_n862_), .B(mai_mai_n854_), .C(mai_mai_n850_), .D(mai_mai_n840_), .Y(mai_mai_n863_));
  NA4        m0841(.A(mai_mai_n863_), .B(mai_mai_n825_), .C(mai_mai_n818_), .D(mai_mai_n392_), .Y(mai3));
  NA2        m0842(.A(i_12_), .B(i_10_), .Y(mai_mai_n865_));
  NA2        m0843(.A(i_6_), .B(i_7_), .Y(mai_mai_n866_));
  NO2        m0844(.A(mai_mai_n866_), .B(i_0_), .Y(mai_mai_n867_));
  NO2        m0845(.A(i_11_), .B(mai_mai_n241_), .Y(mai_mai_n868_));
  OAI210     m0846(.A0(mai_mai_n867_), .A1(mai_mai_n297_), .B0(mai_mai_n868_), .Y(mai_mai_n869_));
  NO2        m0847(.A(mai_mai_n869_), .B(mai_mai_n195_), .Y(mai_mai_n870_));
  NO3        m0848(.A(mai_mai_n473_), .B(mai_mai_n92_), .C(mai_mai_n45_), .Y(mai_mai_n871_));
  OA210      m0849(.A0(mai_mai_n871_), .A1(mai_mai_n870_), .B0(mai_mai_n175_), .Y(mai_mai_n872_));
  NA2        m0850(.A(mai_mai_n428_), .B(mai_mai_n46_), .Y(mai_mai_n873_));
  NO4        m0851(.A(mai_mai_n388_), .B(mai_mai_n395_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n874_));
  NA2        m0852(.A(mai_mai_n187_), .B(mai_mai_n604_), .Y(mai_mai_n875_));
  NOi31      m0853(.An(mai_mai_n875_), .B(mai_mai_n874_), .C(mai_mai_n39_), .Y(mai_mai_n876_));
  NA2        m0854(.A(mai_mai_n733_), .B(mai_mai_n701_), .Y(mai_mai_n877_));
  NA2        m0855(.A(mai_mai_n343_), .B(mai_mai_n458_), .Y(mai_mai_n878_));
  OAI220     m0856(.A0(mai_mai_n878_), .A1(mai_mai_n877_), .B0(mai_mai_n876_), .B1(mai_mai_n63_), .Y(mai_mai_n879_));
  NOi21      m0857(.An(i_5_), .B(i_9_), .Y(mai_mai_n880_));
  NA2        m0858(.A(mai_mai_n880_), .B(mai_mai_n466_), .Y(mai_mai_n881_));
  BUFFER     m0859(.A(mai_mai_n275_), .Y(mai_mai_n882_));
  NA2        m0860(.A(mai_mai_n882_), .B(mai_mai_n498_), .Y(mai_mai_n883_));
  NO3        m0861(.A(mai_mai_n431_), .B(mai_mai_n275_), .C(mai_mai_n73_), .Y(mai_mai_n884_));
  NO2        m0862(.A(mai_mai_n176_), .B(mai_mai_n148_), .Y(mai_mai_n885_));
  AOI210     m0863(.A0(mai_mai_n885_), .A1(mai_mai_n249_), .B0(mai_mai_n884_), .Y(mai_mai_n886_));
  OAI220     m0864(.A0(mai_mai_n886_), .A1(mai_mai_n182_), .B0(mai_mai_n883_), .B1(mai_mai_n881_), .Y(mai_mai_n887_));
  NO3        m0865(.A(mai_mai_n887_), .B(mai_mai_n879_), .C(mai_mai_n872_), .Y(mai_mai_n888_));
  NA2        m0866(.A(mai_mai_n187_), .B(mai_mai_n24_), .Y(mai_mai_n889_));
  NO2        m0867(.A(mai_mai_n699_), .B(mai_mai_n625_), .Y(mai_mai_n890_));
  NO2        m0868(.A(mai_mai_n890_), .B(mai_mai_n889_), .Y(mai_mai_n891_));
  NA2        m0869(.A(mai_mai_n320_), .B(mai_mai_n129_), .Y(mai_mai_n892_));
  NAi21      m0870(.An(mai_mai_n162_), .B(mai_mai_n458_), .Y(mai_mai_n893_));
  OAI220     m0871(.A0(mai_mai_n893_), .A1(mai_mai_n859_), .B0(mai_mai_n892_), .B1(mai_mai_n416_), .Y(mai_mai_n894_));
  NO2        m0872(.A(mai_mai_n894_), .B(mai_mai_n891_), .Y(mai_mai_n895_));
  NO2        m0873(.A(mai_mai_n402_), .B(mai_mai_n301_), .Y(mai_mai_n896_));
  NA2        m0874(.A(mai_mai_n896_), .B(mai_mai_n736_), .Y(mai_mai_n897_));
  NA2        m0875(.A(mai_mai_n605_), .B(i_0_), .Y(mai_mai_n898_));
  NO3        m0876(.A(mai_mai_n898_), .B(mai_mai_n397_), .C(mai_mai_n89_), .Y(mai_mai_n899_));
  INV        m0877(.A(mai_mai_n899_), .Y(mai_mai_n900_));
  INV        m0878(.A(mai_mai_n496_), .Y(mai_mai_n901_));
  AN2        m0879(.A(mai_mai_n98_), .B(mai_mai_n248_), .Y(mai_mai_n902_));
  NA2        m0880(.A(mai_mai_n771_), .B(mai_mai_n338_), .Y(mai_mai_n903_));
  INV        m0881(.A(mai_mai_n58_), .Y(mai_mai_n904_));
  OAI220     m0882(.A0(mai_mai_n904_), .A1(mai_mai_n903_), .B0(mai_mai_n687_), .B1(mai_mai_n564_), .Y(mai_mai_n905_));
  NO2        m0883(.A(mai_mai_n259_), .B(mai_mai_n153_), .Y(mai_mai_n906_));
  NA2        m0884(.A(i_0_), .B(i_10_), .Y(mai_mai_n907_));
  AN2        m0885(.A(mai_mai_n906_), .B(i_6_), .Y(mai_mai_n908_));
  AOI220     m0886(.A0(mai_mai_n343_), .A1(mai_mai_n100_), .B0(mai_mai_n187_), .B1(mai_mai_n84_), .Y(mai_mai_n909_));
  NA2        m0887(.A(mai_mai_n599_), .B(i_4_), .Y(mai_mai_n910_));
  NA2        m0888(.A(mai_mai_n190_), .B(mai_mai_n205_), .Y(mai_mai_n911_));
  OAI220     m0889(.A0(mai_mai_n911_), .A1(mai_mai_n903_), .B0(mai_mai_n910_), .B1(mai_mai_n909_), .Y(mai_mai_n912_));
  NO4        m0890(.A(mai_mai_n912_), .B(mai_mai_n908_), .C(mai_mai_n905_), .D(mai_mai_n902_), .Y(mai_mai_n913_));
  NA4        m0891(.A(mai_mai_n913_), .B(mai_mai_n900_), .C(mai_mai_n897_), .D(mai_mai_n895_), .Y(mai_mai_n914_));
  NA2        m0892(.A(i_11_), .B(i_9_), .Y(mai_mai_n915_));
  NO2        m0893(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n916_));
  NA2        m0894(.A(mai_mai_n407_), .B(mai_mai_n180_), .Y(mai_mai_n917_));
  NA2        m0895(.A(mai_mai_n917_), .B(mai_mai_n160_), .Y(mai_mai_n918_));
  NO2        m0896(.A(mai_mai_n915_), .B(mai_mai_n73_), .Y(mai_mai_n919_));
  NO2        m0897(.A(mai_mai_n176_), .B(i_0_), .Y(mai_mai_n920_));
  INV        m0898(.A(mai_mai_n920_), .Y(mai_mai_n921_));
  NA2        m0899(.A(mai_mai_n496_), .B(mai_mai_n235_), .Y(mai_mai_n922_));
  AOI210     m0900(.A0(mai_mai_n382_), .A1(mai_mai_n42_), .B0(mai_mai_n424_), .Y(mai_mai_n923_));
  OAI220     m0901(.A0(mai_mai_n923_), .A1(mai_mai_n881_), .B0(mai_mai_n922_), .B1(mai_mai_n921_), .Y(mai_mai_n924_));
  NO2        m0902(.A(mai_mai_n924_), .B(mai_mai_n918_), .Y(mai_mai_n925_));
  NA2        m0903(.A(mai_mai_n686_), .B(mai_mai_n121_), .Y(mai_mai_n926_));
  NO2        m0904(.A(i_6_), .B(mai_mai_n926_), .Y(mai_mai_n927_));
  AOI210     m0905(.A0(mai_mai_n468_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n928_));
  NA2        m0906(.A(mai_mai_n172_), .B(mai_mai_n105_), .Y(mai_mai_n929_));
  INV        m0907(.A(mai_mai_n927_), .Y(mai_mai_n930_));
  NOi21      m0908(.An(i_7_), .B(i_5_), .Y(mai_mai_n931_));
  NOi31      m0909(.An(mai_mai_n931_), .B(i_0_), .C(mai_mai_n750_), .Y(mai_mai_n932_));
  NA3        m0910(.A(mai_mai_n932_), .B(mai_mai_n396_), .C(i_6_), .Y(mai_mai_n933_));
  OA210      m0911(.A0(mai_mai_n929_), .A1(mai_mai_n544_), .B0(mai_mai_n933_), .Y(mai_mai_n934_));
  NO3        m0912(.A(mai_mai_n419_), .B(mai_mai_n374_), .C(mai_mai_n370_), .Y(mai_mai_n935_));
  NO2        m0913(.A(mai_mai_n269_), .B(mai_mai_n327_), .Y(mai_mai_n936_));
  NO2        m0914(.A(mai_mai_n750_), .B(mai_mai_n264_), .Y(mai_mai_n937_));
  AOI210     m0915(.A0(mai_mai_n937_), .A1(mai_mai_n936_), .B0(mai_mai_n935_), .Y(mai_mai_n938_));
  NA4        m0916(.A(mai_mai_n938_), .B(mai_mai_n934_), .C(mai_mai_n930_), .D(mai_mai_n925_), .Y(mai_mai_n939_));
  NO2        m0917(.A(mai_mai_n889_), .B(mai_mai_n244_), .Y(mai_mai_n940_));
  AN2        m0918(.A(mai_mai_n342_), .B(mai_mai_n338_), .Y(mai_mai_n941_));
  AO220      m0919(.A0(mai_mai_n941_), .A1(mai_mai_n885_), .B0(mai_mai_n357_), .B1(mai_mai_n27_), .Y(mai_mai_n942_));
  OAI210     m0920(.A0(mai_mai_n942_), .A1(mai_mai_n940_), .B0(i_10_), .Y(mai_mai_n943_));
  NO2        m0921(.A(mai_mai_n865_), .B(mai_mai_n326_), .Y(mai_mai_n944_));
  NA2        m0922(.A(mai_mai_n944_), .B(mai_mai_n919_), .Y(mai_mai_n945_));
  NA3        m0923(.A(mai_mai_n495_), .B(mai_mai_n428_), .C(mai_mai_n46_), .Y(mai_mai_n946_));
  OAI210     m0924(.A0(mai_mai_n893_), .A1(mai_mai_n901_), .B0(mai_mai_n946_), .Y(mai_mai_n947_));
  NO2        m0925(.A(mai_mai_n262_), .B(mai_mai_n47_), .Y(mai_mai_n948_));
  NO2        m0926(.A(mai_mai_n948_), .B(mai_mai_n189_), .Y(mai_mai_n949_));
  AOI220     m0927(.A0(mai_mai_n949_), .A1(mai_mai_n496_), .B0(mai_mai_n947_), .B1(mai_mai_n73_), .Y(mai_mai_n950_));
  NA3        m0928(.A(mai_mai_n842_), .B(mai_mai_n394_), .C(mai_mai_n667_), .Y(mai_mai_n951_));
  NA2        m0929(.A(mai_mai_n95_), .B(mai_mai_n45_), .Y(mai_mai_n952_));
  NO2        m0930(.A(mai_mai_n75_), .B(mai_mai_n773_), .Y(mai_mai_n953_));
  AOI220     m0931(.A0(mai_mai_n953_), .A1(mai_mai_n952_), .B0(mai_mai_n175_), .B1(mai_mai_n625_), .Y(mai_mai_n954_));
  AOI210     m0932(.A0(mai_mai_n954_), .A1(mai_mai_n951_), .B0(mai_mai_n48_), .Y(mai_mai_n955_));
  NO3        m0933(.A(mai_mai_n616_), .B(mai_mai_n369_), .C(mai_mai_n24_), .Y(mai_mai_n956_));
  AOI210     m0934(.A0(mai_mai_n727_), .A1(mai_mai_n576_), .B0(mai_mai_n956_), .Y(mai_mai_n957_));
  NAi21      m0935(.An(i_9_), .B(i_5_), .Y(mai_mai_n958_));
  NO2        m0936(.A(mai_mai_n958_), .B(mai_mai_n419_), .Y(mai_mai_n959_));
  NA2        m0937(.A(mai_mai_n959_), .B(mai_mai_n653_), .Y(mai_mai_n960_));
  OAI220     m0938(.A0(mai_mai_n960_), .A1(mai_mai_n86_), .B0(mai_mai_n957_), .B1(mai_mai_n173_), .Y(mai_mai_n961_));
  NO3        m0939(.A(mai_mai_n961_), .B(mai_mai_n955_), .C(mai_mai_n548_), .Y(mai_mai_n962_));
  NA4        m0940(.A(mai_mai_n962_), .B(mai_mai_n950_), .C(mai_mai_n945_), .D(mai_mai_n943_), .Y(mai_mai_n963_));
  NO3        m0941(.A(mai_mai_n963_), .B(mai_mai_n939_), .C(mai_mai_n914_), .Y(mai_mai_n964_));
  NO2        m0942(.A(i_0_), .B(mai_mai_n750_), .Y(mai_mai_n965_));
  NA2        m0943(.A(mai_mai_n73_), .B(mai_mai_n45_), .Y(mai_mai_n966_));
  NA2        m0944(.A(mai_mai_n907_), .B(mai_mai_n966_), .Y(mai_mai_n967_));
  NO3        m0945(.A(mai_mai_n107_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n968_));
  AO220      m0946(.A0(mai_mai_n968_), .A1(mai_mai_n967_), .B0(mai_mai_n965_), .B1(mai_mai_n175_), .Y(mai_mai_n969_));
  NO2        m0947(.A(mai_mai_n820_), .B(mai_mai_n929_), .Y(mai_mai_n970_));
  AOI210     m0948(.A0(mai_mai_n969_), .A1(mai_mai_n359_), .B0(mai_mai_n970_), .Y(mai_mai_n971_));
  NA2        m0949(.A(mai_mai_n760_), .B(mai_mai_n146_), .Y(mai_mai_n972_));
  INV        m0950(.A(mai_mai_n972_), .Y(mai_mai_n973_));
  NA3        m0951(.A(mai_mai_n973_), .B(mai_mai_n701_), .C(mai_mai_n73_), .Y(mai_mai_n974_));
  NO2        m0952(.A(mai_mai_n838_), .B(mai_mai_n419_), .Y(mai_mai_n975_));
  NA3        m0953(.A(mai_mai_n867_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n976_));
  NA2        m0954(.A(mai_mai_n868_), .B(i_9_), .Y(mai_mai_n977_));
  AOI210     m0955(.A0(mai_mai_n976_), .A1(mai_mai_n523_), .B0(mai_mai_n977_), .Y(mai_mai_n978_));
  OAI210     m0956(.A0(mai_mai_n249_), .A1(i_9_), .B0(mai_mai_n234_), .Y(mai_mai_n979_));
  AOI210     m0957(.A0(mai_mai_n979_), .A1(mai_mai_n898_), .B0(mai_mai_n153_), .Y(mai_mai_n980_));
  NO3        m0958(.A(mai_mai_n980_), .B(mai_mai_n978_), .C(mai_mai_n975_), .Y(mai_mai_n981_));
  NA3        m0959(.A(mai_mai_n981_), .B(mai_mai_n974_), .C(mai_mai_n971_), .Y(mai_mai_n982_));
  NA2        m0960(.A(mai_mai_n941_), .B(mai_mai_n384_), .Y(mai_mai_n983_));
  AOI210     m0961(.A0(mai_mai_n308_), .A1(mai_mai_n162_), .B0(mai_mai_n983_), .Y(mai_mai_n984_));
  NA3        m0962(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n985_));
  NA2        m0963(.A(mai_mai_n916_), .B(mai_mai_n512_), .Y(mai_mai_n986_));
  AOI210     m0964(.A0(mai_mai_n985_), .A1(mai_mai_n162_), .B0(mai_mai_n986_), .Y(mai_mai_n987_));
  NO2        m0965(.A(mai_mai_n987_), .B(mai_mai_n984_), .Y(mai_mai_n988_));
  NO3        m0966(.A(mai_mai_n907_), .B(mai_mai_n880_), .C(mai_mai_n192_), .Y(mai_mai_n989_));
  AOI220     m0967(.A0(mai_mai_n989_), .A1(i_11_), .B0(mai_mai_n600_), .B1(mai_mai_n75_), .Y(mai_mai_n990_));
  NO3        m0968(.A(mai_mai_n212_), .B(mai_mai_n395_), .C(i_0_), .Y(mai_mai_n991_));
  OAI210     m0969(.A0(mai_mai_n991_), .A1(mai_mai_n76_), .B0(i_13_), .Y(mai_mai_n992_));
  INV        m0970(.A(mai_mai_n221_), .Y(mai_mai_n993_));
  OAI220     m0971(.A0(mai_mai_n558_), .A1(mai_mai_n139_), .B0(mai_mai_n672_), .B1(mai_mai_n647_), .Y(mai_mai_n994_));
  NA3        m0972(.A(mai_mai_n994_), .B(mai_mai_n411_), .C(mai_mai_n993_), .Y(mai_mai_n995_));
  NA4        m0973(.A(mai_mai_n995_), .B(mai_mai_n992_), .C(mai_mai_n990_), .D(mai_mai_n988_), .Y(mai_mai_n996_));
  AOI220     m0974(.A0(mai_mai_n931_), .A1(mai_mai_n512_), .B0(mai_mai_n867_), .B1(mai_mai_n163_), .Y(mai_mai_n997_));
  NA2        m0975(.A(mai_mai_n362_), .B(mai_mai_n177_), .Y(mai_mai_n998_));
  OR2        m0976(.A(mai_mai_n998_), .B(mai_mai_n997_), .Y(mai_mai_n999_));
  AOI210     m0977(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n176_), .Y(mai_mai_n1000_));
  NA3        m0978(.A(mai_mai_n644_), .B(mai_mai_n187_), .C(mai_mai_n84_), .Y(mai_mai_n1001_));
  NA2        m0979(.A(mai_mai_n1001_), .B(mai_mai_n574_), .Y(mai_mai_n1002_));
  NO3        m0980(.A(mai_mai_n873_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n1003_));
  NA3        m0981(.A(mai_mai_n517_), .B(mai_mai_n510_), .C(mai_mai_n493_), .Y(mai_mai_n1004_));
  NO3        m0982(.A(mai_mai_n1004_), .B(mai_mai_n1003_), .C(mai_mai_n1002_), .Y(mai_mai_n1005_));
  NA3        m0983(.A(mai_mai_n916_), .B(mai_mai_n297_), .C(mai_mai_n234_), .Y(mai_mai_n1006_));
  INV        m0984(.A(mai_mai_n1006_), .Y(mai_mai_n1007_));
  NA3        m0985(.A(mai_mai_n402_), .B(mai_mai_n344_), .C(mai_mai_n225_), .Y(mai_mai_n1008_));
  OAI210     m0986(.A0(mai_mai_n875_), .A1(mai_mai_n675_), .B0(mai_mai_n1008_), .Y(mai_mai_n1009_));
  NOi31      m0987(.An(mai_mai_n401_), .B(mai_mai_n966_), .C(mai_mai_n244_), .Y(mai_mai_n1010_));
  NO3        m0988(.A(mai_mai_n915_), .B(mai_mai_n221_), .C(mai_mai_n192_), .Y(mai_mai_n1011_));
  NO4        m0989(.A(mai_mai_n1011_), .B(mai_mai_n1010_), .C(mai_mai_n1009_), .D(mai_mai_n1007_), .Y(mai_mai_n1012_));
  NA3        m0990(.A(mai_mai_n1012_), .B(mai_mai_n1005_), .C(mai_mai_n999_), .Y(mai_mai_n1013_));
  INV        m0991(.A(mai_mai_n646_), .Y(mai_mai_n1014_));
  NO3        m0992(.A(mai_mai_n1014_), .B(mai_mai_n590_), .C(mai_mai_n356_), .Y(mai_mai_n1015_));
  NO2        m0993(.A(mai_mai_n86_), .B(i_5_), .Y(mai_mai_n1016_));
  NA3        m0994(.A(mai_mai_n868_), .B(mai_mai_n111_), .C(mai_mai_n124_), .Y(mai_mai_n1017_));
  INV        m0995(.A(mai_mai_n1017_), .Y(mai_mai_n1018_));
  AOI210     m0996(.A0(mai_mai_n1018_), .A1(mai_mai_n1016_), .B0(mai_mai_n1015_), .Y(mai_mai_n1019_));
  NA3        m0997(.A(mai_mai_n313_), .B(i_5_), .C(mai_mai_n195_), .Y(mai_mai_n1020_));
  NA2        m0998(.A(mai_mai_n1020_), .B(mai_mai_n247_), .Y(mai_mai_n1021_));
  NO4        m0999(.A(mai_mai_n244_), .B(mai_mai_n212_), .C(i_0_), .D(i_12_), .Y(mai_mai_n1022_));
  NA2        m1000(.A(mai_mai_n1022_), .B(mai_mai_n1021_), .Y(mai_mai_n1023_));
  AN2        m1001(.A(mai_mai_n907_), .B(mai_mai_n153_), .Y(mai_mai_n1024_));
  NO4        m1002(.A(mai_mai_n1024_), .B(i_12_), .C(mai_mai_n675_), .D(mai_mai_n131_), .Y(mai_mai_n1025_));
  NA2        m1003(.A(mai_mai_n1025_), .B(mai_mai_n221_), .Y(mai_mai_n1026_));
  NA3        m1004(.A(mai_mai_n100_), .B(mai_mai_n604_), .C(i_11_), .Y(mai_mai_n1027_));
  NO2        m1005(.A(mai_mai_n1027_), .B(mai_mai_n155_), .Y(mai_mai_n1028_));
  NA2        m1006(.A(mai_mai_n931_), .B(mai_mai_n492_), .Y(mai_mai_n1029_));
  NA2        m1007(.A(mai_mai_n64_), .B(mai_mai_n103_), .Y(mai_mai_n1030_));
  OAI220     m1008(.A0(mai_mai_n1030_), .A1(mai_mai_n1020_), .B0(mai_mai_n1029_), .B1(mai_mai_n702_), .Y(mai_mai_n1031_));
  AOI210     m1009(.A0(mai_mai_n1031_), .A1(mai_mai_n920_), .B0(mai_mai_n1028_), .Y(mai_mai_n1032_));
  NA4        m1010(.A(mai_mai_n1032_), .B(mai_mai_n1026_), .C(mai_mai_n1023_), .D(mai_mai_n1019_), .Y(mai_mai_n1033_));
  NO4        m1011(.A(mai_mai_n1033_), .B(mai_mai_n1013_), .C(mai_mai_n996_), .D(mai_mai_n982_), .Y(mai_mai_n1034_));
  OAI210     m1012(.A0(mai_mai_n841_), .A1(mai_mai_n834_), .B0(mai_mai_n37_), .Y(mai_mai_n1035_));
  NA3        m1013(.A(mai_mai_n928_), .B(mai_mai_n379_), .C(i_5_), .Y(mai_mai_n1036_));
  NA3        m1014(.A(mai_mai_n1036_), .B(mai_mai_n1035_), .C(mai_mai_n642_), .Y(mai_mai_n1037_));
  NA2        m1015(.A(mai_mai_n1037_), .B(mai_mai_n209_), .Y(mai_mai_n1038_));
  BUFFER     m1016(.A(mai_mai_n380_), .Y(mai_mai_n1039_));
  NA2        m1017(.A(mai_mai_n188_), .B(mai_mai_n190_), .Y(mai_mai_n1040_));
  AO210      m1018(.A0(mai_mai_n1039_), .A1(mai_mai_n33_), .B0(mai_mai_n1040_), .Y(mai_mai_n1041_));
  OAI210     m1019(.A0(mai_mai_n646_), .A1(mai_mai_n644_), .B0(mai_mai_n326_), .Y(mai_mai_n1042_));
  NA2        m1020(.A(mai_mai_n1042_), .B(mai_mai_n1041_), .Y(mai_mai_n1043_));
  NO4        m1021(.A(mai_mai_n237_), .B(mai_mai_n145_), .C(mai_mai_n705_), .D(mai_mai_n37_), .Y(mai_mai_n1044_));
  INV        m1022(.A(mai_mai_n1044_), .Y(mai_mai_n1045_));
  OAI210     m1023(.A0(mai_mai_n1027_), .A1(mai_mai_n148_), .B0(mai_mai_n1045_), .Y(mai_mai_n1046_));
  AOI210     m1024(.A0(mai_mai_n1043_), .A1(mai_mai_n49_), .B0(mai_mai_n1046_), .Y(mai_mai_n1047_));
  AOI210     m1025(.A0(mai_mai_n1047_), .A1(mai_mai_n1038_), .B0(mai_mai_n73_), .Y(mai_mai_n1048_));
  NO2        m1026(.A(mai_mai_n597_), .B(mai_mai_n391_), .Y(mai_mai_n1049_));
  NO2        m1027(.A(mai_mai_n1049_), .B(mai_mai_n779_), .Y(mai_mai_n1050_));
  OAI210     m1028(.A0(mai_mai_n80_), .A1(mai_mai_n55_), .B0(mai_mai_n110_), .Y(mai_mai_n1051_));
  NA2        m1029(.A(mai_mai_n1051_), .B(mai_mai_n76_), .Y(mai_mai_n1052_));
  AOI210     m1030(.A0(mai_mai_n1000_), .A1(mai_mai_n916_), .B0(mai_mai_n932_), .Y(mai_mai_n1053_));
  AOI210     m1031(.A0(mai_mai_n1053_), .A1(mai_mai_n1052_), .B0(mai_mai_n705_), .Y(mai_mai_n1054_));
  NA2        m1032(.A(mai_mai_n269_), .B(mai_mai_n57_), .Y(mai_mai_n1055_));
  AOI220     m1033(.A0(mai_mai_n1055_), .A1(mai_mai_n76_), .B0(mai_mai_n357_), .B1(mai_mai_n261_), .Y(mai_mai_n1056_));
  NO2        m1034(.A(mai_mai_n1056_), .B(mai_mai_n241_), .Y(mai_mai_n1057_));
  NA3        m1035(.A(mai_mai_n98_), .B(mai_mai_n315_), .C(mai_mai_n31_), .Y(mai_mai_n1058_));
  INV        m1036(.A(mai_mai_n1058_), .Y(mai_mai_n1059_));
  NO3        m1037(.A(mai_mai_n1059_), .B(mai_mai_n1057_), .C(mai_mai_n1054_), .Y(mai_mai_n1060_));
  NA2        m1038(.A(mai_mai_n158_), .B(mai_mai_n89_), .Y(mai_mai_n1061_));
  NA3        m1039(.A(mai_mai_n783_), .B(mai_mai_n297_), .C(mai_mai_n80_), .Y(mai_mai_n1062_));
  AOI210     m1040(.A0(mai_mai_n1062_), .A1(mai_mai_n1061_), .B0(i_11_), .Y(mai_mai_n1063_));
  NA2        m1041(.A(mai_mai_n637_), .B(mai_mai_n218_), .Y(mai_mai_n1064_));
  OAI210     m1042(.A0(mai_mai_n1064_), .A1(mai_mai_n928_), .B0(mai_mai_n209_), .Y(mai_mai_n1065_));
  NA2        m1043(.A(mai_mai_n164_), .B(i_5_), .Y(mai_mai_n1066_));
  NO2        m1044(.A(mai_mai_n1065_), .B(mai_mai_n1066_), .Y(mai_mai_n1067_));
  NO4        m1045(.A(mai_mai_n958_), .B(mai_mai_n500_), .C(mai_mai_n258_), .D(mai_mai_n257_), .Y(mai_mai_n1068_));
  NO2        m1046(.A(mai_mai_n1068_), .B(mai_mai_n594_), .Y(mai_mai_n1069_));
  NO2        m1047(.A(mai_mai_n837_), .B(mai_mai_n375_), .Y(mai_mai_n1070_));
  AOI210     m1048(.A0(mai_mai_n1070_), .A1(mai_mai_n1069_), .B0(mai_mai_n41_), .Y(mai_mai_n1071_));
  NO3        m1049(.A(mai_mai_n1071_), .B(mai_mai_n1067_), .C(mai_mai_n1063_), .Y(mai_mai_n1072_));
  OAI210     m1050(.A0(mai_mai_n1060_), .A1(i_4_), .B0(mai_mai_n1072_), .Y(mai_mai_n1073_));
  NO3        m1051(.A(mai_mai_n1073_), .B(mai_mai_n1050_), .C(mai_mai_n1048_), .Y(mai_mai_n1074_));
  NA4        m1052(.A(mai_mai_n1074_), .B(mai_mai_n1034_), .C(mai_mai_n964_), .D(mai_mai_n888_), .Y(mai4));
  INV        m1053(.A(i_2_), .Y(mai_mai_n1078_));
  INV        m1054(.A(mai_mai_n338_), .Y(mai_mai_n1079_));
  INV        m1055(.A(mai_mai_n507_), .Y(mai_mai_n1080_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u0033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  OAI210     u0034(.A0(men_men_n56_), .A1(men_men_n53_), .B0(men_men_n46_), .Y(men_men_n57_));
  NA3        u0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n58_));
  NO2        u0036(.A(i_1_), .B(i_6_), .Y(men_men_n59_));
  NA2        u0037(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  OAI210     u0038(.A0(men_men_n60_), .A1(men_men_n59_), .B0(men_men_n58_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_12_), .Y(men_men_n62_));
  NAi21      u0040(.An(i_2_), .B(i_7_), .Y(men_men_n63_));
  INV        u0041(.A(i_1_), .Y(men_men_n64_));
  NA2        u0042(.A(men_men_n64_), .B(i_6_), .Y(men_men_n65_));
  NA3        u0043(.A(men_men_n65_), .B(men_men_n63_), .C(men_men_n31_), .Y(men_men_n66_));
  NA2        u0044(.A(i_1_), .B(i_10_), .Y(men_men_n67_));
  NO2        u0045(.A(men_men_n67_), .B(i_6_), .Y(men_men_n68_));
  NAi31      u0046(.An(men_men_n68_), .B(men_men_n66_), .C(men_men_n62_), .Y(men_men_n69_));
  NA2        u0047(.A(men_men_n51_), .B(i_2_), .Y(men_men_n70_));
  AOI210     u0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n71_));
  NA2        u0049(.A(i_1_), .B(i_6_), .Y(men_men_n72_));
  NO2        u0050(.A(men_men_n72_), .B(men_men_n25_), .Y(men_men_n73_));
  INV        u0051(.A(i_0_), .Y(men_men_n74_));
  NAi21      u0052(.An(i_5_), .B(i_10_), .Y(men_men_n75_));
  NA2        u0053(.A(i_5_), .B(i_9_), .Y(men_men_n76_));
  AOI210     u0054(.A0(men_men_n76_), .A1(men_men_n75_), .B0(men_men_n74_), .Y(men_men_n77_));
  NO2        u0055(.A(men_men_n77_), .B(men_men_n73_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n78_), .Y(men_men_n79_));
  OAI210     u0057(.A0(men_men_n79_), .A1(men_men_n69_), .B0(i_0_), .Y(men_men_n80_));
  NA2        u0058(.A(i_12_), .B(i_5_), .Y(men_men_n81_));
  NA2        u0059(.A(i_2_), .B(i_8_), .Y(men_men_n82_));
  NO2        u0060(.A(men_men_n82_), .B(men_men_n59_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_9_), .Y(men_men_n84_));
  NO2        u0062(.A(i_3_), .B(i_7_), .Y(men_men_n85_));
  NO3        u0063(.A(men_men_n85_), .B(men_men_n84_), .C(men_men_n64_), .Y(men_men_n86_));
  INV        u0064(.A(i_6_), .Y(men_men_n87_));
  OR4        u0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n88_));
  INV        u0066(.A(men_men_n88_), .Y(men_men_n89_));
  NO2        u0067(.A(i_2_), .B(i_7_), .Y(men_men_n90_));
  OAI210     u0068(.A0(men_men_n86_), .A1(men_men_n83_), .B0(i_2_), .Y(men_men_n91_));
  NAi21      u0069(.An(i_6_), .B(i_10_), .Y(men_men_n92_));
  NA2        u0070(.A(i_6_), .B(i_9_), .Y(men_men_n93_));
  AOI210     u0071(.A0(men_men_n93_), .A1(men_men_n92_), .B0(men_men_n64_), .Y(men_men_n94_));
  NA2        u0072(.A(i_2_), .B(i_6_), .Y(men_men_n95_));
  NO3        u0073(.A(men_men_n95_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n96_));
  NO2        u0074(.A(men_men_n96_), .B(men_men_n94_), .Y(men_men_n97_));
  AOI210     u0075(.A0(men_men_n97_), .A1(men_men_n91_), .B0(men_men_n81_), .Y(men_men_n98_));
  AN3        u0076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n99_));
  NAi21      u0077(.An(i_6_), .B(i_11_), .Y(men_men_n100_));
  NO2        u0078(.A(i_5_), .B(i_8_), .Y(men_men_n101_));
  NOi21      u0079(.An(men_men_n101_), .B(men_men_n100_), .Y(men_men_n102_));
  AOI220     u0080(.A0(men_men_n102_), .A1(men_men_n63_), .B0(men_men_n99_), .B1(men_men_n32_), .Y(men_men_n103_));
  INV        u0081(.A(i_7_), .Y(men_men_n104_));
  NA2        u0082(.A(men_men_n47_), .B(men_men_n104_), .Y(men_men_n105_));
  NO2        u0083(.A(i_0_), .B(i_5_), .Y(men_men_n106_));
  NO2        u0084(.A(men_men_n106_), .B(men_men_n87_), .Y(men_men_n107_));
  NA2        u0085(.A(i_12_), .B(i_3_), .Y(men_men_n108_));
  INV        u0086(.A(men_men_n108_), .Y(men_men_n109_));
  NA3        u0087(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n105_), .Y(men_men_n110_));
  NAi21      u0088(.An(i_7_), .B(i_11_), .Y(men_men_n111_));
  NO3        u0089(.A(men_men_n111_), .B(men_men_n92_), .C(men_men_n54_), .Y(men_men_n112_));
  AN2        u0090(.A(i_2_), .B(i_10_), .Y(men_men_n113_));
  NO2        u0091(.A(men_men_n113_), .B(i_7_), .Y(men_men_n114_));
  OR2        u0092(.A(men_men_n81_), .B(men_men_n59_), .Y(men_men_n115_));
  NO2        u0093(.A(i_8_), .B(men_men_n104_), .Y(men_men_n116_));
  NO3        u0094(.A(men_men_n116_), .B(men_men_n115_), .C(men_men_n114_), .Y(men_men_n117_));
  NA2        u0095(.A(i_12_), .B(i_7_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n64_), .B(men_men_n26_), .Y(men_men_n119_));
  NA2        u0097(.A(men_men_n119_), .B(i_0_), .Y(men_men_n120_));
  NA2        u0098(.A(i_11_), .B(i_12_), .Y(men_men_n121_));
  OAI210     u0099(.A0(men_men_n120_), .A1(men_men_n118_), .B0(men_men_n121_), .Y(men_men_n122_));
  NO2        u0100(.A(men_men_n122_), .B(men_men_n117_), .Y(men_men_n123_));
  NAi41      u0101(.An(men_men_n112_), .B(men_men_n123_), .C(men_men_n110_), .D(men_men_n103_), .Y(men_men_n124_));
  NOi21      u0102(.An(i_1_), .B(i_5_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n125_), .B(i_11_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n104_), .B(men_men_n37_), .Y(men_men_n127_));
  NA2        u0105(.A(i_7_), .B(men_men_n25_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n129_));
  NO2        u0107(.A(men_men_n129_), .B(men_men_n47_), .Y(men_men_n130_));
  NA2        u0108(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n131_));
  NAi21      u0109(.An(i_3_), .B(i_8_), .Y(men_men_n132_));
  NA2        u0110(.A(men_men_n132_), .B(men_men_n63_), .Y(men_men_n133_));
  NOi31      u0111(.An(men_men_n133_), .B(men_men_n131_), .C(men_men_n130_), .Y(men_men_n134_));
  NO2        u0112(.A(i_1_), .B(men_men_n87_), .Y(men_men_n135_));
  NO2        u0113(.A(i_6_), .B(i_5_), .Y(men_men_n136_));
  NA2        u0114(.A(men_men_n136_), .B(i_3_), .Y(men_men_n137_));
  AO210      u0115(.A0(men_men_n137_), .A1(men_men_n48_), .B0(men_men_n135_), .Y(men_men_n138_));
  OAI220     u0116(.A0(men_men_n138_), .A1(men_men_n111_), .B0(men_men_n134_), .B1(men_men_n126_), .Y(men_men_n139_));
  NO3        u0117(.A(men_men_n139_), .B(men_men_n124_), .C(men_men_n98_), .Y(men_men_n140_));
  NA3        u0118(.A(men_men_n140_), .B(men_men_n80_), .C(men_men_n57_), .Y(men2));
  NO2        u0119(.A(men_men_n64_), .B(men_men_n37_), .Y(men_men_n142_));
  NA2        u0120(.A(i_6_), .B(men_men_n25_), .Y(men_men_n143_));
  NA2        u0121(.A(men_men_n143_), .B(men_men_n142_), .Y(men_men_n144_));
  NA4        u0122(.A(men_men_n144_), .B(men_men_n78_), .C(men_men_n70_), .D(men_men_n30_), .Y(men0));
  AN2        u0123(.A(i_8_), .B(i_7_), .Y(men_men_n146_));
  NA2        u0124(.A(men_men_n146_), .B(i_6_), .Y(men_men_n147_));
  NO2        u0125(.A(i_12_), .B(i_13_), .Y(men_men_n148_));
  NAi21      u0126(.An(i_5_), .B(i_11_), .Y(men_men_n149_));
  NOi21      u0127(.An(men_men_n148_), .B(men_men_n149_), .Y(men_men_n150_));
  NO2        u0128(.A(i_0_), .B(i_1_), .Y(men_men_n151_));
  NA2        u0129(.A(i_2_), .B(i_3_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n152_), .B(i_4_), .Y(men_men_n153_));
  NA3        u0131(.A(men_men_n153_), .B(men_men_n151_), .C(men_men_n150_), .Y(men_men_n154_));
  OR2        u0132(.A(men_men_n154_), .B(men_men_n25_), .Y(men_men_n155_));
  AN2        u0133(.A(men_men_n148_), .B(men_men_n84_), .Y(men_men_n156_));
  NO2        u0134(.A(men_men_n156_), .B(men_men_n27_), .Y(men_men_n157_));
  NA2        u0135(.A(i_1_), .B(i_5_), .Y(men_men_n158_));
  NO2        u0136(.A(men_men_n74_), .B(men_men_n47_), .Y(men_men_n159_));
  NA2        u0137(.A(men_men_n159_), .B(men_men_n36_), .Y(men_men_n160_));
  NO3        u0138(.A(men_men_n160_), .B(men_men_n158_), .C(men_men_n157_), .Y(men_men_n161_));
  OR2        u0139(.A(i_0_), .B(i_1_), .Y(men_men_n162_));
  NO3        u0140(.A(men_men_n162_), .B(men_men_n81_), .C(i_13_), .Y(men_men_n163_));
  NAi32      u0141(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n164_));
  NAi21      u0142(.An(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NOi21      u0143(.An(i_4_), .B(i_10_), .Y(men_men_n166_));
  NA2        u0144(.A(men_men_n166_), .B(men_men_n40_), .Y(men_men_n167_));
  NO2        u0145(.A(i_3_), .B(i_5_), .Y(men_men_n168_));
  NO3        u0146(.A(men_men_n74_), .B(i_2_), .C(i_1_), .Y(men_men_n169_));
  NA2        u0147(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  OAI210     u0148(.A0(men_men_n170_), .A1(men_men_n167_), .B0(men_men_n165_), .Y(men_men_n171_));
  NO2        u0149(.A(men_men_n171_), .B(men_men_n161_), .Y(men_men_n172_));
  AOI210     u0150(.A0(men_men_n172_), .A1(men_men_n155_), .B0(men_men_n147_), .Y(men_men_n173_));
  NA3        u0151(.A(men_men_n74_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n174_));
  NA2        u0152(.A(i_3_), .B(men_men_n49_), .Y(men_men_n175_));
  NOi21      u0153(.An(i_4_), .B(i_9_), .Y(men_men_n176_));
  NOi21      u0154(.An(i_11_), .B(i_13_), .Y(men_men_n177_));
  NA2        u0155(.A(men_men_n177_), .B(men_men_n176_), .Y(men_men_n178_));
  OR2        u0156(.A(men_men_n178_), .B(men_men_n175_), .Y(men_men_n179_));
  NO2        u0157(.A(i_4_), .B(i_5_), .Y(men_men_n180_));
  NAi21      u0158(.An(i_12_), .B(i_11_), .Y(men_men_n181_));
  NO2        u0159(.A(men_men_n181_), .B(i_13_), .Y(men_men_n182_));
  NA3        u0160(.A(men_men_n182_), .B(men_men_n180_), .C(men_men_n84_), .Y(men_men_n183_));
  AOI210     u0161(.A0(men_men_n183_), .A1(men_men_n179_), .B0(men_men_n174_), .Y(men_men_n184_));
  NO2        u0162(.A(men_men_n74_), .B(men_men_n64_), .Y(men_men_n185_));
  NA2        u0163(.A(men_men_n185_), .B(men_men_n47_), .Y(men_men_n186_));
  NA2        u0164(.A(men_men_n36_), .B(i_5_), .Y(men_men_n187_));
  NAi31      u0165(.An(men_men_n187_), .B(men_men_n156_), .C(i_11_), .Y(men_men_n188_));
  NA2        u0166(.A(i_3_), .B(i_5_), .Y(men_men_n189_));
  OR2        u0167(.A(men_men_n189_), .B(men_men_n178_), .Y(men_men_n190_));
  AOI210     u0168(.A0(men_men_n190_), .A1(men_men_n188_), .B0(men_men_n186_), .Y(men_men_n191_));
  NO2        u0169(.A(men_men_n74_), .B(i_5_), .Y(men_men_n192_));
  NO2        u0170(.A(i_13_), .B(i_10_), .Y(men_men_n193_));
  NA3        u0171(.A(men_men_n193_), .B(men_men_n192_), .C(men_men_n45_), .Y(men_men_n194_));
  NO2        u0172(.A(i_2_), .B(i_1_), .Y(men_men_n195_));
  NA2        u0173(.A(men_men_n195_), .B(i_3_), .Y(men_men_n196_));
  NAi21      u0174(.An(i_4_), .B(i_12_), .Y(men_men_n197_));
  NO4        u0175(.A(men_men_n197_), .B(men_men_n196_), .C(men_men_n194_), .D(men_men_n25_), .Y(men_men_n198_));
  NO3        u0176(.A(men_men_n198_), .B(men_men_n191_), .C(men_men_n184_), .Y(men_men_n199_));
  INV        u0177(.A(i_8_), .Y(men_men_n200_));
  NO2        u0178(.A(men_men_n200_), .B(i_7_), .Y(men_men_n201_));
  NA2        u0179(.A(men_men_n201_), .B(i_6_), .Y(men_men_n202_));
  NO3        u0180(.A(i_3_), .B(men_men_n87_), .C(men_men_n49_), .Y(men_men_n203_));
  NA2        u0181(.A(men_men_n203_), .B(men_men_n116_), .Y(men_men_n204_));
  NO3        u0182(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n205_));
  NA3        u0183(.A(men_men_n205_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n206_));
  NO3        u0184(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n207_));
  OAI210     u0185(.A0(men_men_n99_), .A1(i_12_), .B0(men_men_n207_), .Y(men_men_n208_));
  AOI210     u0186(.A0(men_men_n208_), .A1(men_men_n206_), .B0(men_men_n204_), .Y(men_men_n209_));
  NO2        u0187(.A(i_3_), .B(i_8_), .Y(men_men_n210_));
  NO3        u0188(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n211_));
  NA3        u0189(.A(men_men_n211_), .B(men_men_n210_), .C(men_men_n40_), .Y(men_men_n212_));
  NO2        u0190(.A(men_men_n106_), .B(men_men_n59_), .Y(men_men_n213_));
  NO2        u0191(.A(i_13_), .B(i_9_), .Y(men_men_n214_));
  NA3        u0192(.A(men_men_n214_), .B(i_6_), .C(men_men_n200_), .Y(men_men_n215_));
  NAi21      u0193(.An(i_12_), .B(i_3_), .Y(men_men_n216_));
  OR2        u0194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n45_), .B(i_5_), .Y(men_men_n218_));
  NO3        u0196(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n219_));
  NA2        u0197(.A(men_men_n219_), .B(i_10_), .Y(men_men_n220_));
  OAI220     u0198(.A0(men_men_n220_), .A1(men_men_n217_), .B0(men_men_n106_), .B1(men_men_n212_), .Y(men_men_n221_));
  AOI210     u0199(.A0(men_men_n221_), .A1(i_7_), .B0(men_men_n209_), .Y(men_men_n222_));
  OAI220     u0200(.A0(men_men_n222_), .A1(i_4_), .B0(men_men_n202_), .B1(men_men_n199_), .Y(men_men_n223_));
  NAi21      u0201(.An(i_12_), .B(i_7_), .Y(men_men_n224_));
  NA3        u0202(.A(i_13_), .B(men_men_n200_), .C(i_10_), .Y(men_men_n225_));
  NO2        u0203(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  NA2        u0204(.A(i_0_), .B(i_5_), .Y(men_men_n227_));
  OAI220     u0205(.A0(men_men_n87_), .A1(men_men_n196_), .B0(men_men_n186_), .B1(men_men_n137_), .Y(men_men_n228_));
  NAi31      u0206(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n229_));
  NO2        u0207(.A(men_men_n36_), .B(i_13_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n47_), .B(men_men_n64_), .Y(men_men_n231_));
  NA3        u0209(.A(men_men_n231_), .B(i_0_), .C(men_men_n230_), .Y(men_men_n232_));
  INV        u0210(.A(i_13_), .Y(men_men_n233_));
  NO2        u0211(.A(i_12_), .B(men_men_n233_), .Y(men_men_n234_));
  NA3        u0212(.A(men_men_n234_), .B(men_men_n205_), .C(men_men_n203_), .Y(men_men_n235_));
  OAI210     u0213(.A0(men_men_n232_), .A1(men_men_n229_), .B0(men_men_n235_), .Y(men_men_n236_));
  AOI220     u0214(.A0(men_men_n236_), .A1(men_men_n146_), .B0(men_men_n228_), .B1(men_men_n226_), .Y(men_men_n237_));
  NO2        u0215(.A(i_12_), .B(men_men_n37_), .Y(men_men_n238_));
  NO2        u0216(.A(men_men_n189_), .B(i_4_), .Y(men_men_n239_));
  NA2        u0217(.A(men_men_n239_), .B(men_men_n238_), .Y(men_men_n240_));
  OR2        u0218(.A(i_8_), .B(i_7_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n241_), .B(men_men_n87_), .Y(men_men_n242_));
  NO2        u0220(.A(men_men_n54_), .B(i_1_), .Y(men_men_n243_));
  NA2        u0221(.A(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  INV        u0222(.A(i_12_), .Y(men_men_n245_));
  NO2        u0223(.A(men_men_n45_), .B(men_men_n245_), .Y(men_men_n246_));
  NO3        u0224(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n247_));
  NA2        u0225(.A(i_2_), .B(i_1_), .Y(men_men_n248_));
  NO2        u0226(.A(men_men_n244_), .B(men_men_n240_), .Y(men_men_n249_));
  NO3        u0227(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n250_));
  NAi21      u0228(.An(i_4_), .B(i_3_), .Y(men_men_n251_));
  NO2        u0229(.A(men_men_n251_), .B(men_men_n76_), .Y(men_men_n252_));
  NO2        u0230(.A(i_0_), .B(i_6_), .Y(men_men_n253_));
  NOi41      u0231(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n254_));
  NA2        u0232(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NO2        u0233(.A(men_men_n248_), .B(men_men_n189_), .Y(men_men_n256_));
  NAi21      u0234(.An(men_men_n255_), .B(men_men_n256_), .Y(men_men_n257_));
  INV        u0235(.A(men_men_n257_), .Y(men_men_n258_));
  AOI220     u0236(.A0(men_men_n258_), .A1(men_men_n40_), .B0(men_men_n249_), .B1(men_men_n214_), .Y(men_men_n259_));
  NO2        u0237(.A(i_11_), .B(men_men_n233_), .Y(men_men_n260_));
  NOi21      u0238(.An(i_1_), .B(i_6_), .Y(men_men_n261_));
  NAi21      u0239(.An(i_3_), .B(i_7_), .Y(men_men_n262_));
  NO2        u0240(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n263_));
  NO2        u0241(.A(i_12_), .B(i_3_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n74_), .B(i_5_), .Y(men_men_n265_));
  NA2        u0243(.A(i_3_), .B(i_9_), .Y(men_men_n266_));
  NAi21      u0244(.An(i_7_), .B(i_10_), .Y(men_men_n267_));
  NO2        u0245(.A(men_men_n267_), .B(men_men_n266_), .Y(men_men_n268_));
  NA3        u0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n269_));
  INV        u0247(.A(men_men_n147_), .Y(men_men_n270_));
  NA2        u0248(.A(men_men_n245_), .B(i_13_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n271_), .B(men_men_n76_), .Y(men_men_n272_));
  NA2        u0250(.A(men_men_n272_), .B(men_men_n270_), .Y(men_men_n273_));
  NO2        u0251(.A(men_men_n241_), .B(men_men_n37_), .Y(men_men_n274_));
  NA2        u0252(.A(i_12_), .B(i_6_), .Y(men_men_n275_));
  OR2        u0253(.A(i_13_), .B(i_9_), .Y(men_men_n276_));
  NO3        u0254(.A(men_men_n276_), .B(men_men_n275_), .C(men_men_n49_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n251_), .B(i_2_), .Y(men_men_n278_));
  NA3        u0256(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n45_), .Y(men_men_n279_));
  NA2        u0257(.A(men_men_n260_), .B(i_9_), .Y(men_men_n280_));
  NA3        u0258(.A(men_men_n265_), .B(men_men_n162_), .C(men_men_n65_), .Y(men_men_n281_));
  OAI210     u0259(.A0(men_men_n281_), .A1(men_men_n280_), .B0(men_men_n279_), .Y(men_men_n282_));
  NA2        u0260(.A(men_men_n159_), .B(men_men_n64_), .Y(men_men_n283_));
  NO3        u0261(.A(i_11_), .B(men_men_n233_), .C(men_men_n25_), .Y(men_men_n284_));
  NO2        u0262(.A(men_men_n262_), .B(i_8_), .Y(men_men_n285_));
  NO2        u0263(.A(i_6_), .B(men_men_n49_), .Y(men_men_n286_));
  NA3        u0264(.A(men_men_n286_), .B(men_men_n285_), .C(men_men_n284_), .Y(men_men_n287_));
  NO3        u0265(.A(men_men_n26_), .B(men_men_n87_), .C(i_5_), .Y(men_men_n288_));
  NA3        u0266(.A(men_men_n288_), .B(men_men_n274_), .C(men_men_n234_), .Y(men_men_n289_));
  AOI210     u0267(.A0(men_men_n289_), .A1(men_men_n287_), .B0(men_men_n283_), .Y(men_men_n290_));
  AOI210     u0268(.A0(men_men_n282_), .A1(men_men_n274_), .B0(men_men_n290_), .Y(men_men_n291_));
  NA4        u0269(.A(men_men_n291_), .B(men_men_n273_), .C(men_men_n259_), .D(men_men_n237_), .Y(men_men_n292_));
  NO3        u0270(.A(i_12_), .B(men_men_n233_), .C(men_men_n37_), .Y(men_men_n293_));
  INV        u0271(.A(men_men_n293_), .Y(men_men_n294_));
  NA2        u0272(.A(i_8_), .B(men_men_n104_), .Y(men_men_n295_));
  NO3        u0273(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n296_));
  AOI220     u0274(.A0(men_men_n296_), .A1(men_men_n203_), .B0(men_men_n168_), .B1(men_men_n243_), .Y(men_men_n297_));
  NO2        u0275(.A(men_men_n297_), .B(men_men_n295_), .Y(men_men_n298_));
  NO3        u0276(.A(i_0_), .B(i_2_), .C(men_men_n64_), .Y(men_men_n299_));
  NO2        u0277(.A(men_men_n248_), .B(i_0_), .Y(men_men_n300_));
  AOI220     u0278(.A0(men_men_n300_), .A1(men_men_n201_), .B0(men_men_n299_), .B1(men_men_n146_), .Y(men_men_n301_));
  NA2        u0279(.A(men_men_n286_), .B(men_men_n26_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n302_), .B(men_men_n301_), .Y(men_men_n303_));
  NA2        u0281(.A(i_0_), .B(i_1_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n304_), .B(i_2_), .Y(men_men_n305_));
  NO2        u0283(.A(men_men_n60_), .B(i_6_), .Y(men_men_n306_));
  NA3        u0284(.A(men_men_n306_), .B(men_men_n305_), .C(men_men_n168_), .Y(men_men_n307_));
  OAI210     u0285(.A0(men_men_n170_), .A1(men_men_n147_), .B0(men_men_n307_), .Y(men_men_n308_));
  NO3        u0286(.A(men_men_n308_), .B(men_men_n303_), .C(men_men_n298_), .Y(men_men_n309_));
  NO2        u0287(.A(i_3_), .B(i_10_), .Y(men_men_n310_));
  NA3        u0288(.A(men_men_n310_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n311_));
  NO2        u0289(.A(i_2_), .B(men_men_n104_), .Y(men_men_n312_));
  NA2        u0290(.A(i_1_), .B(men_men_n36_), .Y(men_men_n313_));
  NOi21      u0291(.An(men_men_n227_), .B(men_men_n106_), .Y(men_men_n314_));
  NA3        u0292(.A(men_men_n314_), .B(i_1_), .C(men_men_n312_), .Y(men_men_n315_));
  AN2        u0293(.A(i_3_), .B(i_10_), .Y(men_men_n316_));
  NA4        u0294(.A(men_men_n316_), .B(men_men_n205_), .C(men_men_n182_), .D(men_men_n180_), .Y(men_men_n317_));
  NO2        u0295(.A(i_5_), .B(men_men_n37_), .Y(men_men_n318_));
  NO2        u0296(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n319_));
  OR2        u0297(.A(men_men_n315_), .B(men_men_n311_), .Y(men_men_n320_));
  OAI220     u0298(.A0(men_men_n320_), .A1(i_6_), .B0(men_men_n309_), .B1(men_men_n294_), .Y(men_men_n321_));
  NO4        u0299(.A(men_men_n321_), .B(men_men_n292_), .C(men_men_n223_), .D(men_men_n173_), .Y(men_men_n322_));
  NO3        u0300(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n323_));
  NO2        u0301(.A(men_men_n60_), .B(men_men_n87_), .Y(men_men_n324_));
  NA2        u0302(.A(men_men_n300_), .B(men_men_n324_), .Y(men_men_n325_));
  NO3        u0303(.A(i_6_), .B(men_men_n200_), .C(i_7_), .Y(men_men_n326_));
  NA2        u0304(.A(men_men_n326_), .B(men_men_n205_), .Y(men_men_n327_));
  AOI210     u0305(.A0(men_men_n327_), .A1(men_men_n325_), .B0(men_men_n175_), .Y(men_men_n328_));
  NO2        u0306(.A(i_2_), .B(i_3_), .Y(men_men_n329_));
  OR2        u0307(.A(i_0_), .B(i_5_), .Y(men_men_n330_));
  NA2        u0308(.A(men_men_n227_), .B(men_men_n330_), .Y(men_men_n331_));
  NA4        u0309(.A(men_men_n331_), .B(men_men_n242_), .C(men_men_n329_), .D(i_1_), .Y(men_men_n332_));
  NA3        u0310(.A(men_men_n300_), .B(men_men_n168_), .C(men_men_n116_), .Y(men_men_n333_));
  NAi21      u0311(.An(i_8_), .B(i_7_), .Y(men_men_n334_));
  NO2        u0312(.A(men_men_n334_), .B(i_6_), .Y(men_men_n335_));
  NO2        u0313(.A(men_men_n162_), .B(men_men_n47_), .Y(men_men_n336_));
  NA3        u0314(.A(men_men_n336_), .B(men_men_n335_), .C(men_men_n168_), .Y(men_men_n337_));
  NA3        u0315(.A(men_men_n337_), .B(men_men_n333_), .C(men_men_n332_), .Y(men_men_n338_));
  OAI210     u0316(.A0(men_men_n338_), .A1(men_men_n328_), .B0(i_4_), .Y(men_men_n339_));
  NO2        u0317(.A(i_12_), .B(i_10_), .Y(men_men_n340_));
  NOi21      u0318(.An(i_5_), .B(i_0_), .Y(men_men_n341_));
  AOI210     u0319(.A0(i_2_), .A1(men_men_n49_), .B0(men_men_n104_), .Y(men_men_n342_));
  NO4        u0320(.A(men_men_n342_), .B(men_men_n313_), .C(men_men_n341_), .D(men_men_n132_), .Y(men_men_n343_));
  NA4        u0321(.A(men_men_n85_), .B(men_men_n36_), .C(men_men_n87_), .D(i_8_), .Y(men_men_n344_));
  NA2        u0322(.A(men_men_n343_), .B(men_men_n340_), .Y(men_men_n345_));
  NO2        u0323(.A(i_6_), .B(i_8_), .Y(men_men_n346_));
  NOi21      u0324(.An(i_0_), .B(i_2_), .Y(men_men_n347_));
  AN2        u0325(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NO2        u0326(.A(i_1_), .B(i_7_), .Y(men_men_n349_));
  AO220      u0327(.A0(men_men_n349_), .A1(men_men_n348_), .B0(men_men_n335_), .B1(men_men_n243_), .Y(men_men_n350_));
  NA3        u0328(.A(men_men_n350_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n351_));
  NA3        u0329(.A(men_men_n351_), .B(men_men_n345_), .C(men_men_n339_), .Y(men_men_n352_));
  NO3        u0330(.A(men_men_n241_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n353_));
  NO3        u0331(.A(men_men_n334_), .B(i_2_), .C(i_1_), .Y(men_men_n354_));
  OAI210     u0332(.A0(men_men_n354_), .A1(men_men_n353_), .B0(i_6_), .Y(men_men_n355_));
  NA3        u0333(.A(men_men_n261_), .B(men_men_n312_), .C(men_men_n200_), .Y(men_men_n356_));
  AOI210     u0334(.A0(men_men_n356_), .A1(men_men_n355_), .B0(men_men_n331_), .Y(men_men_n357_));
  NOi21      u0335(.An(men_men_n158_), .B(men_men_n107_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n358_), .B(men_men_n128_), .Y(men_men_n359_));
  OAI210     u0337(.A0(men_men_n359_), .A1(men_men_n357_), .B0(i_3_), .Y(men_men_n360_));
  INV        u0338(.A(men_men_n85_), .Y(men_men_n361_));
  NO2        u0339(.A(men_men_n304_), .B(men_men_n82_), .Y(men_men_n362_));
  NA2        u0340(.A(men_men_n362_), .B(men_men_n136_), .Y(men_men_n363_));
  NO2        u0341(.A(men_men_n95_), .B(men_men_n200_), .Y(men_men_n364_));
  NA3        u0342(.A(men_men_n314_), .B(men_men_n364_), .C(men_men_n64_), .Y(men_men_n365_));
  AOI210     u0343(.A0(men_men_n365_), .A1(men_men_n363_), .B0(men_men_n361_), .Y(men_men_n366_));
  NO2        u0344(.A(men_men_n200_), .B(i_9_), .Y(men_men_n367_));
  NA3        u0345(.A(men_men_n367_), .B(men_men_n213_), .C(men_men_n162_), .Y(men_men_n368_));
  NO2        u0346(.A(men_men_n368_), .B(men_men_n47_), .Y(men_men_n369_));
  NO3        u0347(.A(men_men_n369_), .B(men_men_n366_), .C(men_men_n303_), .Y(men_men_n370_));
  AOI210     u0348(.A0(men_men_n370_), .A1(men_men_n360_), .B0(men_men_n167_), .Y(men_men_n371_));
  AOI210     u0349(.A0(men_men_n352_), .A1(men_men_n323_), .B0(men_men_n371_), .Y(men_men_n372_));
  NOi32      u0350(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n373_));
  INV        u0351(.A(men_men_n373_), .Y(men_men_n374_));
  NAi21      u0352(.An(i_0_), .B(i_6_), .Y(men_men_n375_));
  NAi21      u0353(.An(i_1_), .B(i_5_), .Y(men_men_n376_));
  NA2        u0354(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n377_));
  NA2        u0355(.A(men_men_n377_), .B(men_men_n25_), .Y(men_men_n378_));
  OAI210     u0356(.A0(men_men_n378_), .A1(men_men_n164_), .B0(men_men_n255_), .Y(men_men_n379_));
  NAi41      u0357(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n380_));
  OAI220     u0358(.A0(men_men_n380_), .A1(men_men_n376_), .B0(men_men_n229_), .B1(men_men_n164_), .Y(men_men_n381_));
  AOI210     u0359(.A0(men_men_n380_), .A1(men_men_n164_), .B0(men_men_n162_), .Y(men_men_n382_));
  NOi32      u0360(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n383_));
  NAi21      u0361(.An(i_6_), .B(i_1_), .Y(men_men_n384_));
  NA3        u0362(.A(men_men_n384_), .B(men_men_n383_), .C(men_men_n47_), .Y(men_men_n385_));
  NO2        u0363(.A(men_men_n385_), .B(i_0_), .Y(men_men_n386_));
  OR3        u0364(.A(men_men_n386_), .B(men_men_n382_), .C(men_men_n381_), .Y(men_men_n387_));
  NO2        u0365(.A(i_1_), .B(men_men_n104_), .Y(men_men_n388_));
  NAi21      u0366(.An(i_3_), .B(i_4_), .Y(men_men_n389_));
  NO2        u0367(.A(men_men_n389_), .B(i_9_), .Y(men_men_n390_));
  AN2        u0368(.A(i_6_), .B(i_7_), .Y(men_men_n391_));
  OAI210     u0369(.A0(men_men_n391_), .A1(men_men_n388_), .B0(men_men_n390_), .Y(men_men_n392_));
  NA2        u0370(.A(i_2_), .B(i_7_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n389_), .B(i_10_), .Y(men_men_n394_));
  NO2        u0372(.A(men_men_n392_), .B(men_men_n192_), .Y(men_men_n395_));
  AOI210     u0373(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n396_));
  OAI210     u0374(.A0(men_men_n396_), .A1(men_men_n195_), .B0(men_men_n394_), .Y(men_men_n397_));
  AOI220     u0375(.A0(men_men_n394_), .A1(men_men_n349_), .B0(men_men_n247_), .B1(men_men_n195_), .Y(men_men_n398_));
  AOI210     u0376(.A0(men_men_n398_), .A1(men_men_n397_), .B0(i_5_), .Y(men_men_n399_));
  NO4        u0377(.A(men_men_n399_), .B(men_men_n395_), .C(men_men_n387_), .D(men_men_n379_), .Y(men_men_n400_));
  NO2        u0378(.A(men_men_n400_), .B(men_men_n374_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n60_), .B(men_men_n25_), .Y(men_men_n402_));
  AN2        u0380(.A(i_12_), .B(i_5_), .Y(men_men_n403_));
  NO2        u0381(.A(i_4_), .B(men_men_n26_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n404_), .B(men_men_n403_), .Y(men_men_n405_));
  NO2        u0383(.A(i_11_), .B(i_6_), .Y(men_men_n406_));
  NA3        u0384(.A(men_men_n406_), .B(men_men_n336_), .C(men_men_n233_), .Y(men_men_n407_));
  NO2        u0385(.A(men_men_n407_), .B(men_men_n405_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n251_), .B(i_5_), .Y(men_men_n409_));
  NO2        u0387(.A(i_5_), .B(i_10_), .Y(men_men_n410_));
  AOI220     u0388(.A0(men_men_n410_), .A1(men_men_n278_), .B0(men_men_n409_), .B1(men_men_n205_), .Y(men_men_n411_));
  NA2        u0389(.A(men_men_n148_), .B(men_men_n46_), .Y(men_men_n412_));
  NO2        u0390(.A(men_men_n412_), .B(men_men_n411_), .Y(men_men_n413_));
  OAI210     u0391(.A0(men_men_n413_), .A1(men_men_n408_), .B0(men_men_n402_), .Y(men_men_n414_));
  NO2        u0392(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n154_), .B(men_men_n87_), .Y(men_men_n416_));
  OAI210     u0394(.A0(men_men_n416_), .A1(men_men_n408_), .B0(men_men_n415_), .Y(men_men_n417_));
  NO3        u0395(.A(men_men_n87_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n418_));
  NO2        u0396(.A(i_3_), .B(men_men_n104_), .Y(men_men_n419_));
  NO2        u0397(.A(i_11_), .B(i_12_), .Y(men_men_n420_));
  NA2        u0398(.A(men_men_n410_), .B(men_men_n245_), .Y(men_men_n421_));
  NA3        u0399(.A(men_men_n116_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n422_));
  OAI220     u0400(.A0(men_men_n422_), .A1(men_men_n229_), .B0(men_men_n421_), .B1(men_men_n344_), .Y(men_men_n423_));
  NAi21      u0401(.An(i_13_), .B(i_0_), .Y(men_men_n424_));
  NO2        u0402(.A(men_men_n424_), .B(men_men_n248_), .Y(men_men_n425_));
  NA2        u0403(.A(men_men_n423_), .B(men_men_n425_), .Y(men_men_n426_));
  NA3        u0404(.A(men_men_n426_), .B(men_men_n417_), .C(men_men_n414_), .Y(men_men_n427_));
  NA2        u0405(.A(men_men_n45_), .B(men_men_n233_), .Y(men_men_n428_));
  NO3        u0406(.A(i_1_), .B(i_12_), .C(men_men_n87_), .Y(men_men_n429_));
  NO2        u0407(.A(i_0_), .B(i_11_), .Y(men_men_n430_));
  INV        u0408(.A(i_5_), .Y(men_men_n431_));
  AN2        u0409(.A(i_1_), .B(i_6_), .Y(men_men_n432_));
  NOi21      u0410(.An(i_2_), .B(i_12_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n433_), .B(men_men_n432_), .Y(men_men_n434_));
  NO2        u0412(.A(men_men_n434_), .B(men_men_n431_), .Y(men_men_n435_));
  NA2        u0413(.A(men_men_n146_), .B(i_9_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(i_4_), .Y(men_men_n437_));
  NA2        u0415(.A(men_men_n435_), .B(men_men_n437_), .Y(men_men_n438_));
  OR2        u0416(.A(i_13_), .B(i_10_), .Y(men_men_n439_));
  NO2        u0417(.A(men_men_n178_), .B(men_men_n127_), .Y(men_men_n440_));
  OR2        u0418(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n104_), .B(men_men_n25_), .Y(men_men_n442_));
  NA2        u0420(.A(men_men_n293_), .B(men_men_n442_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n286_), .B(men_men_n219_), .Y(men_men_n444_));
  OAI220     u0422(.A0(men_men_n444_), .A1(men_men_n441_), .B0(men_men_n443_), .B1(men_men_n358_), .Y(men_men_n445_));
  INV        u0423(.A(men_men_n445_), .Y(men_men_n446_));
  AOI210     u0424(.A0(men_men_n446_), .A1(men_men_n438_), .B0(men_men_n26_), .Y(men_men_n447_));
  NA2        u0425(.A(men_men_n333_), .B(men_men_n332_), .Y(men_men_n448_));
  AOI220     u0426(.A0(men_men_n306_), .A1(men_men_n296_), .B0(men_men_n300_), .B1(men_men_n324_), .Y(men_men_n449_));
  NO2        u0427(.A(men_men_n449_), .B(men_men_n175_), .Y(men_men_n450_));
  NO2        u0428(.A(men_men_n189_), .B(men_men_n87_), .Y(men_men_n451_));
  AOI220     u0429(.A0(men_men_n451_), .A1(men_men_n305_), .B0(men_men_n288_), .B1(men_men_n219_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n452_), .B(men_men_n295_), .Y(men_men_n453_));
  NO3        u0431(.A(men_men_n453_), .B(men_men_n450_), .C(men_men_n448_), .Y(men_men_n454_));
  NA2        u0432(.A(men_men_n203_), .B(men_men_n99_), .Y(men_men_n455_));
  NA3        u0433(.A(men_men_n336_), .B(men_men_n168_), .C(men_men_n87_), .Y(men_men_n456_));
  AOI210     u0434(.A0(men_men_n456_), .A1(men_men_n455_), .B0(men_men_n334_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n306_), .B(men_men_n243_), .Y(men_men_n458_));
  NO2        u0436(.A(men_men_n458_), .B(men_men_n189_), .Y(men_men_n459_));
  NO2        u0437(.A(i_3_), .B(men_men_n49_), .Y(men_men_n460_));
  NA3        u0438(.A(men_men_n349_), .B(men_men_n348_), .C(men_men_n460_), .Y(men_men_n461_));
  NA2        u0439(.A(men_men_n326_), .B(men_men_n331_), .Y(men_men_n462_));
  OAI210     u0440(.A0(men_men_n462_), .A1(men_men_n196_), .B0(men_men_n461_), .Y(men_men_n463_));
  NO3        u0441(.A(men_men_n463_), .B(men_men_n459_), .C(men_men_n457_), .Y(men_men_n464_));
  AOI210     u0442(.A0(men_men_n464_), .A1(men_men_n454_), .B0(men_men_n280_), .Y(men_men_n465_));
  NO4        u0443(.A(men_men_n465_), .B(men_men_n447_), .C(men_men_n427_), .D(men_men_n401_), .Y(men_men_n466_));
  NO2        u0444(.A(men_men_n64_), .B(i_4_), .Y(men_men_n467_));
  NO2        u0445(.A(men_men_n74_), .B(i_13_), .Y(men_men_n468_));
  NA3        u0446(.A(men_men_n468_), .B(men_men_n467_), .C(i_2_), .Y(men_men_n469_));
  NO2        u0447(.A(i_10_), .B(i_9_), .Y(men_men_n470_));
  NAi21      u0448(.An(i_12_), .B(i_8_), .Y(men_men_n471_));
  NO2        u0449(.A(men_men_n471_), .B(i_3_), .Y(men_men_n472_));
  NA2        u0450(.A(men_men_n472_), .B(men_men_n470_), .Y(men_men_n473_));
  NO2        u0451(.A(men_men_n47_), .B(i_4_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n474_), .B(men_men_n107_), .Y(men_men_n475_));
  OAI220     u0453(.A0(men_men_n475_), .A1(men_men_n212_), .B0(men_men_n473_), .B1(men_men_n469_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n319_), .B(i_0_), .Y(men_men_n477_));
  NO3        u0455(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n275_), .B(men_men_n100_), .Y(men_men_n479_));
  NA2        u0457(.A(men_men_n479_), .B(men_men_n478_), .Y(men_men_n480_));
  NA2        u0458(.A(i_8_), .B(i_9_), .Y(men_men_n481_));
  NO2        u0459(.A(men_men_n480_), .B(men_men_n477_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n260_), .B(men_men_n318_), .Y(men_men_n483_));
  NO3        u0461(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n484_));
  AOI210     u0462(.A0(men_men_n264_), .A1(men_men_n195_), .B0(men_men_n484_), .Y(men_men_n485_));
  NA3        u0463(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n486_));
  NA4        u0464(.A(men_men_n149_), .B(men_men_n119_), .C(men_men_n81_), .D(men_men_n23_), .Y(men_men_n487_));
  OAI220     u0465(.A0(men_men_n487_), .A1(men_men_n486_), .B0(men_men_n485_), .B1(men_men_n483_), .Y(men_men_n488_));
  NO3        u0466(.A(men_men_n488_), .B(men_men_n482_), .C(men_men_n476_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n305_), .B(men_men_n111_), .Y(men_men_n490_));
  OR2        u0468(.A(men_men_n490_), .B(men_men_n215_), .Y(men_men_n491_));
  OA210      u0469(.A0(men_men_n368_), .A1(men_men_n104_), .B0(men_men_n307_), .Y(men_men_n492_));
  OA220      u0470(.A0(men_men_n492_), .A1(men_men_n167_), .B0(men_men_n491_), .B1(men_men_n240_), .Y(men_men_n493_));
  NA2        u0471(.A(men_men_n99_), .B(i_13_), .Y(men_men_n494_));
  NA2        u0472(.A(men_men_n451_), .B(men_men_n402_), .Y(men_men_n495_));
  NO2        u0473(.A(i_2_), .B(i_13_), .Y(men_men_n496_));
  NA3        u0474(.A(men_men_n496_), .B(men_men_n166_), .C(men_men_n102_), .Y(men_men_n497_));
  OAI220     u0475(.A0(men_men_n497_), .A1(men_men_n245_), .B0(men_men_n495_), .B1(men_men_n494_), .Y(men_men_n498_));
  NO3        u0476(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n499_));
  NO2        u0477(.A(i_6_), .B(i_7_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n500_), .B(men_men_n499_), .Y(men_men_n501_));
  NO2        u0479(.A(i_11_), .B(i_1_), .Y(men_men_n502_));
  OR2        u0480(.A(i_11_), .B(i_8_), .Y(men_men_n503_));
  NOi21      u0481(.An(i_2_), .B(i_7_), .Y(men_men_n504_));
  NAi31      u0482(.An(men_men_n503_), .B(men_men_n504_), .C(i_0_), .Y(men_men_n505_));
  NO2        u0483(.A(men_men_n439_), .B(i_6_), .Y(men_men_n506_));
  NA3        u0484(.A(men_men_n506_), .B(men_men_n467_), .C(men_men_n76_), .Y(men_men_n507_));
  NO2        u0485(.A(men_men_n507_), .B(men_men_n505_), .Y(men_men_n508_));
  NO2        u0486(.A(i_3_), .B(men_men_n200_), .Y(men_men_n509_));
  NO2        u0487(.A(i_6_), .B(i_10_), .Y(men_men_n510_));
  NA4        u0488(.A(men_men_n510_), .B(men_men_n323_), .C(men_men_n509_), .D(men_men_n245_), .Y(men_men_n511_));
  NO2        u0489(.A(men_men_n511_), .B(men_men_n160_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n513_));
  NO2        u0491(.A(men_men_n162_), .B(i_3_), .Y(men_men_n514_));
  NAi31      u0492(.An(men_men_n513_), .B(men_men_n514_), .C(men_men_n234_), .Y(men_men_n515_));
  NA3        u0493(.A(men_men_n415_), .B(men_men_n185_), .C(men_men_n153_), .Y(men_men_n516_));
  NA2        u0494(.A(men_men_n516_), .B(men_men_n515_), .Y(men_men_n517_));
  NO4        u0495(.A(men_men_n517_), .B(men_men_n512_), .C(men_men_n508_), .D(men_men_n498_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n478_), .B(men_men_n403_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n484_), .B(men_men_n410_), .Y(men_men_n520_));
  NO2        u0498(.A(men_men_n520_), .B(men_men_n232_), .Y(men_men_n521_));
  NAi21      u0499(.An(men_men_n225_), .B(men_men_n420_), .Y(men_men_n522_));
  NA2        u0500(.A(men_men_n349_), .B(men_men_n227_), .Y(men_men_n523_));
  NO2        u0501(.A(men_men_n26_), .B(i_5_), .Y(men_men_n524_));
  NO2        u0502(.A(i_0_), .B(men_men_n87_), .Y(men_men_n525_));
  NA3        u0503(.A(men_men_n525_), .B(men_men_n524_), .C(men_men_n146_), .Y(men_men_n526_));
  OR3        u0504(.A(men_men_n313_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n527_));
  OAI220     u0505(.A0(men_men_n527_), .A1(men_men_n526_), .B0(men_men_n523_), .B1(men_men_n522_), .Y(men_men_n528_));
  NA4        u0506(.A(men_men_n316_), .B(men_men_n231_), .C(men_men_n74_), .D(men_men_n245_), .Y(men_men_n529_));
  NO2        u0507(.A(men_men_n529_), .B(men_men_n501_), .Y(men_men_n530_));
  NO3        u0508(.A(men_men_n530_), .B(men_men_n528_), .C(men_men_n521_), .Y(men_men_n531_));
  NA4        u0509(.A(men_men_n531_), .B(men_men_n518_), .C(men_men_n493_), .D(men_men_n489_), .Y(men_men_n532_));
  NA3        u0510(.A(men_men_n316_), .B(men_men_n182_), .C(men_men_n180_), .Y(men_men_n533_));
  OAI210     u0511(.A0(men_men_n311_), .A1(men_men_n187_), .B0(men_men_n533_), .Y(men_men_n534_));
  AN2        u0512(.A(men_men_n296_), .B(men_men_n242_), .Y(men_men_n535_));
  NA2        u0513(.A(men_men_n535_), .B(men_men_n534_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n126_), .B(men_men_n115_), .Y(men_men_n537_));
  AN2        u0515(.A(men_men_n537_), .B(men_men_n478_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n323_), .B(men_men_n169_), .Y(men_men_n539_));
  OAI210     u0517(.A0(men_men_n539_), .A1(men_men_n240_), .B0(men_men_n317_), .Y(men_men_n540_));
  AOI220     u0518(.A0(men_men_n540_), .A1(men_men_n335_), .B0(men_men_n538_), .B1(men_men_n319_), .Y(men_men_n541_));
  NA4        u0519(.A(men_men_n468_), .B(men_men_n467_), .C(men_men_n210_), .D(i_2_), .Y(men_men_n542_));
  INV        u0520(.A(men_men_n542_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n373_), .B(men_men_n74_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n391_), .B(men_men_n383_), .Y(men_men_n545_));
  NO2        u0523(.A(men_men_n36_), .B(i_8_), .Y(men_men_n546_));
  NA2        u0524(.A(men_men_n39_), .B(i_13_), .Y(men_men_n547_));
  INV        u0525(.A(men_men_n547_), .Y(men_men_n548_));
  AOI210     u0526(.A0(men_men_n543_), .A1(men_men_n211_), .B0(men_men_n548_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n265_), .B(men_men_n65_), .Y(men_men_n550_));
  OAI210     u0528(.A0(i_8_), .A1(men_men_n550_), .B0(men_men_n138_), .Y(men_men_n551_));
  AOI210     u0529(.A0(men_men_n201_), .A1(i_9_), .B0(men_men_n274_), .Y(men_men_n552_));
  NO2        u0530(.A(men_men_n552_), .B(men_men_n206_), .Y(men_men_n553_));
  NO2        u0531(.A(men_men_n189_), .B(men_men_n87_), .Y(men_men_n554_));
  AOI220     u0532(.A0(men_men_n554_), .A1(men_men_n553_), .B0(men_men_n551_), .B1(men_men_n440_), .Y(men_men_n555_));
  NA4        u0533(.A(men_men_n555_), .B(men_men_n549_), .C(men_men_n541_), .D(men_men_n536_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n409_), .B(men_men_n305_), .Y(men_men_n557_));
  OAI210     u0535(.A0(men_men_n405_), .A1(men_men_n174_), .B0(men_men_n557_), .Y(men_men_n558_));
  NO2        u0536(.A(i_12_), .B(men_men_n200_), .Y(men_men_n559_));
  NA2        u0537(.A(men_men_n559_), .B(men_men_n233_), .Y(men_men_n560_));
  NA2        u0538(.A(men_men_n510_), .B(men_men_n27_), .Y(men_men_n561_));
  NO3        u0539(.A(men_men_n561_), .B(men_men_n560_), .C(men_men_n490_), .Y(men_men_n562_));
  NOi31      u0540(.An(men_men_n326_), .B(men_men_n439_), .C(men_men_n38_), .Y(men_men_n563_));
  OAI210     u0541(.A0(men_men_n563_), .A1(men_men_n562_), .B0(men_men_n558_), .Y(men_men_n564_));
  NO2        u0542(.A(i_8_), .B(i_7_), .Y(men_men_n565_));
  OAI210     u0543(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n566_));
  NA2        u0544(.A(men_men_n566_), .B(men_men_n231_), .Y(men_men_n567_));
  AOI220     u0545(.A0(men_men_n336_), .A1(men_men_n40_), .B0(men_men_n243_), .B1(men_men_n214_), .Y(men_men_n568_));
  OAI220     u0546(.A0(men_men_n568_), .A1(men_men_n189_), .B0(men_men_n567_), .B1(men_men_n251_), .Y(men_men_n569_));
  NA2        u0547(.A(men_men_n45_), .B(i_10_), .Y(men_men_n570_));
  NO2        u0548(.A(men_men_n570_), .B(i_6_), .Y(men_men_n571_));
  NA3        u0549(.A(men_men_n571_), .B(men_men_n569_), .C(men_men_n565_), .Y(men_men_n572_));
  AOI220     u0550(.A0(men_men_n451_), .A1(men_men_n336_), .B0(men_men_n256_), .B1(men_men_n253_), .Y(men_men_n573_));
  OAI220     u0551(.A0(men_men_n573_), .A1(men_men_n271_), .B0(men_men_n494_), .B1(men_men_n137_), .Y(men_men_n574_));
  NA2        u0552(.A(men_men_n574_), .B(men_men_n274_), .Y(men_men_n575_));
  NOi31      u0553(.An(men_men_n300_), .B(men_men_n311_), .C(men_men_n187_), .Y(men_men_n576_));
  NA3        u0554(.A(men_men_n316_), .B(men_men_n180_), .C(men_men_n99_), .Y(men_men_n577_));
  NO2        u0555(.A(men_men_n230_), .B(men_men_n45_), .Y(men_men_n578_));
  NO2        u0556(.A(men_men_n162_), .B(i_5_), .Y(men_men_n579_));
  NA3        u0557(.A(men_men_n579_), .B(men_men_n428_), .C(men_men_n329_), .Y(men_men_n580_));
  OAI210     u0558(.A0(men_men_n580_), .A1(men_men_n578_), .B0(men_men_n577_), .Y(men_men_n581_));
  OAI210     u0559(.A0(men_men_n581_), .A1(men_men_n576_), .B0(men_men_n484_), .Y(men_men_n582_));
  NA4        u0560(.A(men_men_n582_), .B(men_men_n575_), .C(men_men_n572_), .D(men_men_n564_), .Y(men_men_n583_));
  NA2        u0561(.A(men_men_n293_), .B(men_men_n85_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n363_), .B(men_men_n584_), .Y(men_men_n585_));
  NA2        u0563(.A(men_men_n306_), .B(men_men_n296_), .Y(men_men_n586_));
  NO2        u0564(.A(men_men_n586_), .B(men_men_n179_), .Y(men_men_n587_));
  AOI210     u0565(.A0(men_men_n384_), .A1(men_men_n47_), .B0(men_men_n388_), .Y(men_men_n588_));
  NA2        u0566(.A(i_0_), .B(men_men_n49_), .Y(men_men_n589_));
  NA3        u0567(.A(men_men_n559_), .B(men_men_n284_), .C(men_men_n589_), .Y(men_men_n590_));
  NO2        u0568(.A(men_men_n588_), .B(men_men_n590_), .Y(men_men_n591_));
  NO3        u0569(.A(men_men_n591_), .B(men_men_n587_), .C(men_men_n585_), .Y(men_men_n592_));
  NO4        u0570(.A(men_men_n261_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n593_));
  NO3        u0571(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n594_));
  NO2        u0572(.A(men_men_n241_), .B(men_men_n36_), .Y(men_men_n595_));
  AN2        u0573(.A(men_men_n595_), .B(men_men_n594_), .Y(men_men_n596_));
  OA210      u0574(.A0(men_men_n596_), .A1(men_men_n593_), .B0(men_men_n373_), .Y(men_men_n597_));
  NO2        u0575(.A(men_men_n439_), .B(i_1_), .Y(men_men_n598_));
  NOi31      u0576(.An(men_men_n598_), .B(men_men_n479_), .C(men_men_n74_), .Y(men_men_n599_));
  AN4        u0577(.A(men_men_n599_), .B(men_men_n437_), .C(men_men_n524_), .D(i_2_), .Y(men_men_n600_));
  NO2        u0578(.A(men_men_n449_), .B(men_men_n183_), .Y(men_men_n601_));
  NO3        u0579(.A(men_men_n601_), .B(men_men_n600_), .C(men_men_n597_), .Y(men_men_n602_));
  NOi21      u0580(.An(i_10_), .B(i_6_), .Y(men_men_n603_));
  NO2        u0581(.A(men_men_n87_), .B(men_men_n25_), .Y(men_men_n604_));
  AOI220     u0582(.A0(men_men_n293_), .A1(men_men_n604_), .B0(men_men_n284_), .B1(men_men_n603_), .Y(men_men_n605_));
  NO2        u0583(.A(men_men_n605_), .B(men_men_n477_), .Y(men_men_n606_));
  NO2        u0584(.A(men_men_n118_), .B(men_men_n23_), .Y(men_men_n607_));
  NA2        u0585(.A(men_men_n326_), .B(men_men_n169_), .Y(men_men_n608_));
  AOI220     u0586(.A0(men_men_n608_), .A1(men_men_n458_), .B0(men_men_n190_), .B1(men_men_n188_), .Y(men_men_n609_));
  NO2        u0587(.A(men_men_n205_), .B(men_men_n37_), .Y(men_men_n610_));
  NOi31      u0588(.An(men_men_n150_), .B(men_men_n610_), .C(men_men_n344_), .Y(men_men_n611_));
  NO3        u0589(.A(men_men_n611_), .B(men_men_n609_), .C(men_men_n606_), .Y(men_men_n612_));
  NO2        u0590(.A(men_men_n544_), .B(men_men_n398_), .Y(men_men_n613_));
  INV        u0591(.A(men_men_n329_), .Y(men_men_n614_));
  NO2        u0592(.A(i_12_), .B(men_men_n87_), .Y(men_men_n615_));
  NA3        u0593(.A(men_men_n615_), .B(men_men_n284_), .C(men_men_n589_), .Y(men_men_n616_));
  NA3        u0594(.A(men_men_n406_), .B(men_men_n293_), .C(men_men_n227_), .Y(men_men_n617_));
  AOI210     u0595(.A0(men_men_n617_), .A1(men_men_n616_), .B0(men_men_n614_), .Y(men_men_n618_));
  NO3        u0596(.A(i_4_), .B(men_men_n355_), .C(men_men_n311_), .Y(men_men_n619_));
  OR2        u0597(.A(i_2_), .B(i_5_), .Y(men_men_n620_));
  NO3        u0598(.A(men_men_n619_), .B(men_men_n618_), .C(men_men_n613_), .Y(men_men_n621_));
  NA4        u0599(.A(men_men_n621_), .B(men_men_n612_), .C(men_men_n602_), .D(men_men_n592_), .Y(men_men_n622_));
  NO4        u0600(.A(men_men_n622_), .B(men_men_n583_), .C(men_men_n556_), .D(men_men_n532_), .Y(men_men_n623_));
  NA4        u0601(.A(men_men_n623_), .B(men_men_n466_), .C(men_men_n372_), .D(men_men_n322_), .Y(men7));
  NO2        u0602(.A(men_men_n95_), .B(men_men_n55_), .Y(men_men_n625_));
  NO2        u0603(.A(men_men_n111_), .B(men_men_n92_), .Y(men_men_n626_));
  NA2        u0604(.A(men_men_n404_), .B(men_men_n626_), .Y(men_men_n627_));
  NA2        u0605(.A(men_men_n510_), .B(men_men_n85_), .Y(men_men_n628_));
  NA2        u0606(.A(i_11_), .B(men_men_n200_), .Y(men_men_n629_));
  NA2        u0607(.A(men_men_n148_), .B(men_men_n629_), .Y(men_men_n630_));
  OAI210     u0608(.A0(men_men_n630_), .A1(men_men_n628_), .B0(men_men_n627_), .Y(men_men_n631_));
  NA3        u0609(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n632_));
  NO2        u0610(.A(men_men_n245_), .B(i_4_), .Y(men_men_n633_));
  NA2        u0611(.A(men_men_n633_), .B(i_8_), .Y(men_men_n634_));
  NO2        u0612(.A(men_men_n108_), .B(men_men_n632_), .Y(men_men_n635_));
  NA2        u0613(.A(i_2_), .B(men_men_n87_), .Y(men_men_n636_));
  OAI210     u0614(.A0(men_men_n90_), .A1(men_men_n210_), .B0(men_men_n211_), .Y(men_men_n637_));
  NO2        u0615(.A(i_7_), .B(men_men_n37_), .Y(men_men_n638_));
  NA2        u0616(.A(i_4_), .B(i_8_), .Y(men_men_n639_));
  AOI210     u0617(.A0(men_men_n639_), .A1(men_men_n316_), .B0(men_men_n638_), .Y(men_men_n640_));
  OAI220     u0618(.A0(men_men_n640_), .A1(men_men_n636_), .B0(men_men_n637_), .B1(i_13_), .Y(men_men_n641_));
  NO4        u0619(.A(men_men_n641_), .B(men_men_n635_), .C(men_men_n631_), .D(men_men_n625_), .Y(men_men_n642_));
  AOI210     u0620(.A0(men_men_n132_), .A1(men_men_n63_), .B0(i_10_), .Y(men_men_n643_));
  AOI210     u0621(.A0(men_men_n643_), .A1(men_men_n245_), .B0(men_men_n166_), .Y(men_men_n644_));
  OR2        u0622(.A(i_6_), .B(i_10_), .Y(men_men_n645_));
  NO2        u0623(.A(men_men_n645_), .B(men_men_n23_), .Y(men_men_n646_));
  OR3        u0624(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n647_));
  NO3        u0625(.A(men_men_n647_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n648_));
  INV        u0626(.A(men_men_n207_), .Y(men_men_n649_));
  NO2        u0627(.A(men_men_n648_), .B(men_men_n646_), .Y(men_men_n650_));
  OA220      u0628(.A0(men_men_n650_), .A1(men_men_n614_), .B0(men_men_n644_), .B1(men_men_n276_), .Y(men_men_n651_));
  AOI210     u0629(.A0(men_men_n651_), .A1(men_men_n642_), .B0(men_men_n64_), .Y(men_men_n652_));
  NOi21      u0630(.An(i_11_), .B(i_7_), .Y(men_men_n653_));
  AO210      u0631(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n654_));
  NO2        u0632(.A(men_men_n654_), .B(men_men_n653_), .Y(men_men_n655_));
  NA2        u0633(.A(men_men_n655_), .B(men_men_n214_), .Y(men_men_n656_));
  NA3        u0634(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n657_));
  NAi31      u0635(.An(men_men_n657_), .B(men_men_n224_), .C(i_11_), .Y(men_men_n658_));
  AOI210     u0636(.A0(men_men_n658_), .A1(men_men_n656_), .B0(men_men_n64_), .Y(men_men_n659_));
  NA2        u0637(.A(men_men_n89_), .B(men_men_n64_), .Y(men_men_n660_));
  AO210      u0638(.A0(men_men_n660_), .A1(men_men_n398_), .B0(men_men_n41_), .Y(men_men_n661_));
  NO3        u0639(.A(men_men_n267_), .B(men_men_n216_), .C(men_men_n629_), .Y(men_men_n662_));
  OAI210     u0640(.A0(men_men_n662_), .A1(men_men_n234_), .B0(men_men_n64_), .Y(men_men_n663_));
  NA2        u0641(.A(men_men_n433_), .B(men_men_n31_), .Y(men_men_n664_));
  OR2        u0642(.A(men_men_n216_), .B(men_men_n111_), .Y(men_men_n665_));
  NA2        u0643(.A(men_men_n665_), .B(men_men_n664_), .Y(men_men_n666_));
  NO2        u0644(.A(men_men_n64_), .B(i_9_), .Y(men_men_n667_));
  NO2        u0645(.A(men_men_n667_), .B(i_4_), .Y(men_men_n668_));
  NA2        u0646(.A(men_men_n668_), .B(men_men_n666_), .Y(men_men_n669_));
  NO2        u0647(.A(i_1_), .B(i_12_), .Y(men_men_n670_));
  NA3        u0648(.A(men_men_n670_), .B(men_men_n113_), .C(men_men_n24_), .Y(men_men_n671_));
  NA4        u0649(.A(men_men_n671_), .B(men_men_n669_), .C(men_men_n663_), .D(men_men_n661_), .Y(men_men_n672_));
  OAI210     u0650(.A0(men_men_n672_), .A1(men_men_n659_), .B0(i_6_), .Y(men_men_n673_));
  NO2        u0651(.A(men_men_n245_), .B(men_men_n87_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(i_11_), .Y(men_men_n675_));
  INV        u0653(.A(men_men_n480_), .Y(men_men_n676_));
  NO4        u0654(.A(men_men_n224_), .B(men_men_n132_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n677_));
  NA2        u0655(.A(men_men_n677_), .B(men_men_n667_), .Y(men_men_n678_));
  NA2        u0656(.A(men_men_n245_), .B(i_6_), .Y(men_men_n679_));
  NO3        u0657(.A(men_men_n645_), .B(men_men_n241_), .C(men_men_n23_), .Y(men_men_n680_));
  AOI210     u0658(.A0(i_1_), .A1(men_men_n268_), .B0(men_men_n680_), .Y(men_men_n681_));
  OAI210     u0659(.A0(men_men_n681_), .A1(men_men_n45_), .B0(men_men_n678_), .Y(men_men_n682_));
  NA3        u0660(.A(men_men_n565_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n683_));
  NA2        u0661(.A(men_men_n142_), .B(i_9_), .Y(men_men_n684_));
  NA3        u0662(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n47_), .B(i_1_), .Y(men_men_n686_));
  NA3        u0664(.A(men_men_n686_), .B(men_men_n275_), .C(men_men_n45_), .Y(men_men_n687_));
  OAI220     u0665(.A0(men_men_n687_), .A1(men_men_n685_), .B0(men_men_n684_), .B1(men_men_n1112_), .Y(men_men_n688_));
  NA3        u0666(.A(men_men_n667_), .B(men_men_n329_), .C(i_6_), .Y(men_men_n689_));
  NO2        u0667(.A(men_men_n689_), .B(men_men_n23_), .Y(men_men_n690_));
  AOI210     u0668(.A0(men_men_n502_), .A1(men_men_n442_), .B0(men_men_n250_), .Y(men_men_n691_));
  NO2        u0669(.A(men_men_n691_), .B(men_men_n636_), .Y(men_men_n692_));
  NAi21      u0670(.An(men_men_n683_), .B(men_men_n94_), .Y(men_men_n693_));
  NA2        u0671(.A(men_men_n686_), .B(men_men_n275_), .Y(men_men_n694_));
  NO2        u0672(.A(i_11_), .B(men_men_n37_), .Y(men_men_n695_));
  NA2        u0673(.A(men_men_n695_), .B(men_men_n24_), .Y(men_men_n696_));
  OAI210     u0674(.A0(men_men_n696_), .A1(men_men_n694_), .B0(men_men_n693_), .Y(men_men_n697_));
  OR4        u0675(.A(men_men_n697_), .B(men_men_n692_), .C(men_men_n690_), .D(men_men_n688_), .Y(men_men_n698_));
  NO3        u0676(.A(men_men_n698_), .B(men_men_n682_), .C(men_men_n676_), .Y(men_men_n699_));
  NO2        u0677(.A(men_men_n245_), .B(men_men_n104_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n700_), .B(men_men_n653_), .Y(men_men_n701_));
  NA2        u0679(.A(men_men_n701_), .B(i_1_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n702_), .B(men_men_n647_), .Y(men_men_n703_));
  NA2        u0681(.A(men_men_n703_), .B(men_men_n47_), .Y(men_men_n704_));
  NA2        u0682(.A(i_3_), .B(men_men_n200_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(men_men_n118_), .Y(men_men_n706_));
  AN2        u0684(.A(men_men_n706_), .B(men_men_n571_), .Y(men_men_n707_));
  NO2        u0685(.A(men_men_n241_), .B(men_men_n45_), .Y(men_men_n708_));
  NO3        u0686(.A(men_men_n708_), .B(men_men_n319_), .C(men_men_n246_), .Y(men_men_n709_));
  NO2        u0687(.A(men_men_n121_), .B(men_men_n37_), .Y(men_men_n710_));
  NO2        u0688(.A(men_men_n710_), .B(i_6_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n87_), .B(i_9_), .Y(men_men_n712_));
  NO2        u0690(.A(men_men_n712_), .B(men_men_n64_), .Y(men_men_n713_));
  NO2        u0691(.A(men_men_n713_), .B(men_men_n670_), .Y(men_men_n714_));
  NO4        u0692(.A(men_men_n714_), .B(men_men_n711_), .C(men_men_n709_), .D(i_4_), .Y(men_men_n715_));
  NA2        u0693(.A(i_1_), .B(i_3_), .Y(men_men_n716_));
  NO2        u0694(.A(men_men_n481_), .B(men_men_n95_), .Y(men_men_n717_));
  AOI210     u0695(.A0(men_men_n708_), .A1(men_men_n603_), .B0(men_men_n717_), .Y(men_men_n718_));
  NO2        u0696(.A(men_men_n718_), .B(men_men_n716_), .Y(men_men_n719_));
  NO3        u0697(.A(men_men_n719_), .B(men_men_n715_), .C(men_men_n707_), .Y(men_men_n720_));
  NA4        u0698(.A(men_men_n720_), .B(men_men_n704_), .C(men_men_n699_), .D(men_men_n673_), .Y(men_men_n721_));
  NO3        u0699(.A(men_men_n503_), .B(i_3_), .C(i_7_), .Y(men_men_n722_));
  NOi21      u0700(.An(men_men_n722_), .B(i_10_), .Y(men_men_n723_));
  OA210      u0701(.A0(men_men_n723_), .A1(men_men_n254_), .B0(men_men_n87_), .Y(men_men_n724_));
  NA2        u0702(.A(men_men_n391_), .B(men_men_n390_), .Y(men_men_n725_));
  NA3        u0703(.A(men_men_n510_), .B(men_men_n546_), .C(men_men_n47_), .Y(men_men_n726_));
  NO3        u0704(.A(men_men_n504_), .B(men_men_n639_), .C(men_men_n87_), .Y(men_men_n727_));
  NA2        u0705(.A(men_men_n727_), .B(men_men_n25_), .Y(men_men_n728_));
  NA3        u0706(.A(men_men_n166_), .B(men_men_n85_), .C(men_men_n87_), .Y(men_men_n729_));
  NA4        u0707(.A(men_men_n729_), .B(men_men_n728_), .C(men_men_n726_), .D(men_men_n725_), .Y(men_men_n730_));
  OAI210     u0708(.A0(men_men_n730_), .A1(men_men_n724_), .B0(i_1_), .Y(men_men_n731_));
  AOI210     u0709(.A0(men_men_n275_), .A1(men_men_n100_), .B0(i_1_), .Y(men_men_n732_));
  NO2        u0710(.A(men_men_n389_), .B(i_2_), .Y(men_men_n733_));
  NA2        u0711(.A(men_men_n733_), .B(men_men_n732_), .Y(men_men_n734_));
  OAI210     u0712(.A0(men_men_n689_), .A1(men_men_n471_), .B0(men_men_n734_), .Y(men_men_n735_));
  INV        u0713(.A(men_men_n735_), .Y(men_men_n736_));
  AOI210     u0714(.A0(men_men_n736_), .A1(men_men_n731_), .B0(i_13_), .Y(men_men_n737_));
  OR2        u0715(.A(i_11_), .B(i_7_), .Y(men_men_n738_));
  NA3        u0716(.A(men_men_n738_), .B(men_men_n109_), .C(men_men_n142_), .Y(men_men_n739_));
  AOI220     u0717(.A0(men_men_n496_), .A1(men_men_n166_), .B0(men_men_n474_), .B1(men_men_n142_), .Y(men_men_n740_));
  OAI210     u0718(.A0(men_men_n740_), .A1(men_men_n45_), .B0(men_men_n739_), .Y(men_men_n741_));
  AOI210     u0719(.A0(men_men_n685_), .A1(men_men_n55_), .B0(i_12_), .Y(men_men_n742_));
  NO2        u0720(.A(men_men_n1111_), .B(men_men_n95_), .Y(men_men_n743_));
  AOI210     u0721(.A0(men_men_n741_), .A1(men_men_n346_), .B0(men_men_n743_), .Y(men_men_n744_));
  NA2        u0722(.A(men_men_n118_), .B(men_men_n111_), .Y(men_men_n745_));
  AOI220     u0723(.A0(men_men_n745_), .A1(men_men_n73_), .B0(men_men_n406_), .B1(men_men_n686_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n746_), .B(men_men_n251_), .Y(men_men_n747_));
  AOI210     u0725(.A0(men_men_n471_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n748_));
  NA2        u0726(.A(men_men_n131_), .B(i_13_), .Y(men_men_n749_));
  NO2        u0727(.A(men_men_n685_), .B(men_men_n118_), .Y(men_men_n750_));
  NO2        u0728(.A(men_men_n749_), .B(men_men_n732_), .Y(men_men_n751_));
  NO3        u0729(.A(men_men_n72_), .B(men_men_n32_), .C(men_men_n104_), .Y(men_men_n752_));
  NA2        u0730(.A(men_men_n26_), .B(men_men_n200_), .Y(men_men_n753_));
  NA2        u0731(.A(men_men_n753_), .B(i_7_), .Y(men_men_n754_));
  NO3        u0732(.A(men_men_n504_), .B(men_men_n245_), .C(men_men_n87_), .Y(men_men_n755_));
  AOI210     u0733(.A0(men_men_n755_), .A1(men_men_n754_), .B0(men_men_n752_), .Y(men_men_n756_));
  AOI220     u0734(.A0(men_men_n406_), .A1(men_men_n686_), .B0(men_men_n94_), .B1(men_men_n105_), .Y(men_men_n757_));
  OAI220     u0735(.A0(men_men_n757_), .A1(men_men_n634_), .B0(men_men_n756_), .B1(men_men_n649_), .Y(men_men_n758_));
  NO3        u0736(.A(men_men_n758_), .B(men_men_n751_), .C(men_men_n747_), .Y(men_men_n759_));
  OR2        u0737(.A(i_11_), .B(i_6_), .Y(men_men_n760_));
  NA3        u0738(.A(men_men_n633_), .B(men_men_n753_), .C(i_7_), .Y(men_men_n761_));
  NO2        u0739(.A(men_men_n761_), .B(men_men_n760_), .Y(men_men_n762_));
  NA3        u0740(.A(men_men_n433_), .B(men_men_n638_), .C(men_men_n100_), .Y(men_men_n763_));
  NA2        u0741(.A(men_men_n675_), .B(i_13_), .Y(men_men_n764_));
  NAi21      u0742(.An(i_11_), .B(i_12_), .Y(men_men_n765_));
  NOi41      u0743(.An(men_men_n114_), .B(men_men_n765_), .C(i_13_), .D(men_men_n87_), .Y(men_men_n766_));
  NO3        u0744(.A(men_men_n504_), .B(men_men_n615_), .C(men_men_n639_), .Y(men_men_n767_));
  AOI220     u0745(.A0(men_men_n767_), .A1(men_men_n323_), .B0(men_men_n766_), .B1(men_men_n47_), .Y(men_men_n768_));
  NA3        u0746(.A(men_men_n768_), .B(men_men_n764_), .C(men_men_n763_), .Y(men_men_n769_));
  OAI210     u0747(.A0(men_men_n769_), .A1(men_men_n762_), .B0(men_men_n64_), .Y(men_men_n770_));
  NO2        u0748(.A(i_2_), .B(i_12_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n388_), .B(men_men_n771_), .Y(men_men_n772_));
  NA2        u0750(.A(i_8_), .B(men_men_n25_), .Y(men_men_n773_));
  NO3        u0751(.A(men_men_n773_), .B(men_men_n404_), .C(men_men_n633_), .Y(men_men_n774_));
  OAI210     u0752(.A0(men_men_n774_), .A1(men_men_n390_), .B0(men_men_n388_), .Y(men_men_n775_));
  NO2        u0753(.A(men_men_n132_), .B(i_2_), .Y(men_men_n776_));
  NA2        u0754(.A(men_men_n776_), .B(men_men_n670_), .Y(men_men_n777_));
  NA3        u0755(.A(men_men_n777_), .B(men_men_n775_), .C(men_men_n772_), .Y(men_men_n778_));
  NA3        u0756(.A(men_men_n778_), .B(men_men_n46_), .C(men_men_n233_), .Y(men_men_n779_));
  NA4        u0757(.A(men_men_n779_), .B(men_men_n770_), .C(men_men_n759_), .D(men_men_n744_), .Y(men_men_n780_));
  OR4        u0758(.A(men_men_n780_), .B(men_men_n737_), .C(men_men_n721_), .D(men_men_n652_), .Y(men5));
  AOI210     u0759(.A0(men_men_n701_), .A1(men_men_n278_), .B0(men_men_n440_), .Y(men_men_n782_));
  AN2        u0760(.A(men_men_n24_), .B(i_10_), .Y(men_men_n783_));
  NA3        u0761(.A(men_men_n783_), .B(men_men_n771_), .C(men_men_n111_), .Y(men_men_n784_));
  NO2        u0762(.A(men_men_n634_), .B(i_11_), .Y(men_men_n785_));
  OAI210     u0763(.A0(men_men_n638_), .A1(men_men_n90_), .B0(men_men_n785_), .Y(men_men_n786_));
  NA3        u0764(.A(men_men_n786_), .B(men_men_n784_), .C(men_men_n782_), .Y(men_men_n787_));
  NO3        u0765(.A(i_11_), .B(men_men_n245_), .C(i_13_), .Y(men_men_n788_));
  NO2        u0766(.A(men_men_n128_), .B(men_men_n23_), .Y(men_men_n789_));
  NA2        u0767(.A(i_12_), .B(i_8_), .Y(men_men_n790_));
  OAI210     u0768(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n790_), .Y(men_men_n791_));
  INV        u0769(.A(men_men_n470_), .Y(men_men_n792_));
  AOI220     u0770(.A0(men_men_n329_), .A1(men_men_n607_), .B0(men_men_n791_), .B1(men_men_n789_), .Y(men_men_n793_));
  INV        u0771(.A(men_men_n793_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n794_), .B(men_men_n787_), .Y(men_men_n795_));
  INV        u0773(.A(men_men_n177_), .Y(men_men_n796_));
  INV        u0774(.A(men_men_n254_), .Y(men_men_n797_));
  OAI210     u0775(.A0(men_men_n733_), .A1(men_men_n472_), .B0(men_men_n114_), .Y(men_men_n798_));
  AOI210     u0776(.A0(men_men_n798_), .A1(men_men_n797_), .B0(men_men_n796_), .Y(men_men_n799_));
  NO2        u0777(.A(men_men_n481_), .B(men_men_n26_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n800_), .B(men_men_n442_), .Y(men_men_n801_));
  NA2        u0779(.A(men_men_n801_), .B(i_2_), .Y(men_men_n802_));
  INV        u0780(.A(men_men_n802_), .Y(men_men_n803_));
  AOI210     u0781(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n439_), .Y(men_men_n804_));
  AOI210     u0782(.A0(men_men_n804_), .A1(men_men_n803_), .B0(men_men_n799_), .Y(men_men_n805_));
  NO2        u0783(.A(men_men_n197_), .B(men_men_n129_), .Y(men_men_n806_));
  OAI210     u0784(.A0(men_men_n806_), .A1(men_men_n789_), .B0(i_2_), .Y(men_men_n807_));
  INV        u0785(.A(men_men_n178_), .Y(men_men_n808_));
  NO3        u0786(.A(men_men_n654_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n809_));
  AOI210     u0787(.A0(men_men_n808_), .A1(men_men_n90_), .B0(men_men_n809_), .Y(men_men_n810_));
  AOI210     u0788(.A0(men_men_n810_), .A1(men_men_n807_), .B0(men_men_n200_), .Y(men_men_n811_));
  OA210      u0789(.A0(men_men_n655_), .A1(men_men_n130_), .B0(i_13_), .Y(men_men_n812_));
  NA2        u0790(.A(men_men_n207_), .B(men_men_n210_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n156_), .B(men_men_n629_), .Y(men_men_n814_));
  AOI210     u0792(.A0(men_men_n814_), .A1(men_men_n813_), .B0(men_men_n393_), .Y(men_men_n815_));
  AOI210     u0793(.A0(men_men_n216_), .A1(men_men_n152_), .B0(men_men_n546_), .Y(men_men_n816_));
  OAI210     u0794(.A0(men_men_n816_), .A1(men_men_n234_), .B0(men_men_n442_), .Y(men_men_n817_));
  NO2        u0795(.A(men_men_n105_), .B(men_men_n45_), .Y(men_men_n818_));
  INV        u0796(.A(men_men_n312_), .Y(men_men_n819_));
  NA4        u0797(.A(men_men_n819_), .B(men_men_n316_), .C(men_men_n128_), .D(men_men_n43_), .Y(men_men_n820_));
  OAI210     u0798(.A0(men_men_n820_), .A1(men_men_n818_), .B0(men_men_n817_), .Y(men_men_n821_));
  NO4        u0799(.A(men_men_n821_), .B(men_men_n815_), .C(men_men_n812_), .D(men_men_n811_), .Y(men_men_n822_));
  NA2        u0800(.A(men_men_n607_), .B(men_men_n28_), .Y(men_men_n823_));
  NA2        u0801(.A(men_men_n788_), .B(men_men_n285_), .Y(men_men_n824_));
  NA2        u0802(.A(men_men_n824_), .B(men_men_n823_), .Y(men_men_n825_));
  NO2        u0803(.A(men_men_n63_), .B(i_12_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n826_), .B(men_men_n130_), .Y(men_men_n827_));
  NO2        u0805(.A(men_men_n827_), .B(men_men_n629_), .Y(men_men_n828_));
  AOI220     u0806(.A0(men_men_n828_), .A1(men_men_n36_), .B0(men_men_n825_), .B1(men_men_n47_), .Y(men_men_n829_));
  NA4        u0807(.A(men_men_n829_), .B(men_men_n822_), .C(men_men_n805_), .D(men_men_n795_), .Y(men6));
  NO3        u0808(.A(men_men_n263_), .B(men_men_n318_), .C(i_1_), .Y(men_men_n831_));
  NO2        u0809(.A(men_men_n192_), .B(men_men_n143_), .Y(men_men_n832_));
  OAI210     u0810(.A0(men_men_n832_), .A1(men_men_n831_), .B0(men_men_n776_), .Y(men_men_n833_));
  NA4        u0811(.A(men_men_n410_), .B(men_men_n509_), .C(men_men_n72_), .D(men_men_n104_), .Y(men_men_n834_));
  INV        u0812(.A(men_men_n834_), .Y(men_men_n835_));
  NO2        u0813(.A(i_11_), .B(i_9_), .Y(men_men_n836_));
  NO2        u0814(.A(men_men_n835_), .B(men_men_n341_), .Y(men_men_n837_));
  AO210      u0815(.A0(men_men_n837_), .A1(men_men_n833_), .B0(i_12_), .Y(men_men_n838_));
  NA2        u0816(.A(men_men_n394_), .B(men_men_n349_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n615_), .B(men_men_n64_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n723_), .B(men_men_n72_), .Y(men_men_n841_));
  NA4        u0819(.A(men_men_n660_), .B(men_men_n841_), .C(men_men_n840_), .D(men_men_n839_), .Y(men_men_n842_));
  INV        u0820(.A(men_men_n204_), .Y(men_men_n843_));
  AOI220     u0821(.A0(men_men_n843_), .A1(men_men_n836_), .B0(men_men_n842_), .B1(men_men_n74_), .Y(men_men_n844_));
  INV        u0822(.A(men_men_n340_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n76_), .B(men_men_n135_), .Y(men_men_n846_));
  INV        u0824(.A(men_men_n128_), .Y(men_men_n847_));
  NA2        u0825(.A(men_men_n847_), .B(men_men_n47_), .Y(men_men_n848_));
  AOI210     u0826(.A0(men_men_n848_), .A1(men_men_n846_), .B0(men_men_n845_), .Y(men_men_n849_));
  NO2        u0827(.A(men_men_n545_), .B(men_men_n192_), .Y(men_men_n850_));
  NO2        u0828(.A(men_men_n32_), .B(i_11_), .Y(men_men_n851_));
  NA3        u0829(.A(men_men_n851_), .B(men_men_n500_), .C(men_men_n410_), .Y(men_men_n852_));
  NAi32      u0830(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n853_));
  AOI210     u0831(.A0(men_men_n760_), .A1(men_men_n88_), .B0(men_men_n853_), .Y(men_men_n854_));
  OAI210     u0832(.A0(men_men_n722_), .A1(men_men_n595_), .B0(men_men_n594_), .Y(men_men_n855_));
  NAi31      u0833(.An(men_men_n854_), .B(men_men_n855_), .C(men_men_n852_), .Y(men_men_n856_));
  OR3        u0834(.A(men_men_n856_), .B(men_men_n850_), .C(men_men_n849_), .Y(men_men_n857_));
  NO2        u0835(.A(men_men_n738_), .B(i_2_), .Y(men_men_n858_));
  NA2        u0836(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n859_));
  OAI210     u0837(.A0(men_men_n859_), .A1(men_men_n432_), .B0(men_men_n378_), .Y(men_men_n860_));
  NA2        u0838(.A(men_men_n860_), .B(men_men_n858_), .Y(men_men_n861_));
  AO220      u0839(.A0(men_men_n377_), .A1(men_men_n367_), .B0(men_men_n418_), .B1(men_men_n629_), .Y(men_men_n862_));
  NA3        u0840(.A(men_men_n862_), .B(men_men_n264_), .C(i_7_), .Y(men_men_n863_));
  OR2        u0841(.A(men_men_n655_), .B(men_men_n472_), .Y(men_men_n864_));
  NA3        u0842(.A(men_men_n864_), .B(men_men_n151_), .C(men_men_n70_), .Y(men_men_n865_));
  AO210      u0843(.A0(men_men_n520_), .A1(men_men_n792_), .B0(men_men_n36_), .Y(men_men_n866_));
  NA4        u0844(.A(men_men_n866_), .B(men_men_n865_), .C(men_men_n863_), .D(men_men_n861_), .Y(men_men_n867_));
  OAI210     u0845(.A0(men_men_n674_), .A1(i_11_), .B0(men_men_n88_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n868_), .B(men_men_n594_), .Y(men_men_n869_));
  NA3        u0847(.A(men_men_n393_), .B(men_men_n247_), .C(men_men_n151_), .Y(men_men_n870_));
  OAI210     u0848(.A0(men_men_n418_), .A1(men_men_n211_), .B0(men_men_n71_), .Y(men_men_n871_));
  NA4        u0849(.A(men_men_n871_), .B(men_men_n870_), .C(men_men_n869_), .D(men_men_n637_), .Y(men_men_n872_));
  AO210      u0850(.A0(men_men_n546_), .A1(men_men_n47_), .B0(men_men_n89_), .Y(men_men_n873_));
  NA3        u0851(.A(men_men_n873_), .B(men_men_n510_), .C(men_men_n227_), .Y(men_men_n874_));
  AOI210     u0852(.A0(men_men_n472_), .A1(men_men_n470_), .B0(men_men_n593_), .Y(men_men_n875_));
  NO2        u0853(.A(men_men_n645_), .B(men_men_n105_), .Y(men_men_n876_));
  OAI210     u0854(.A0(men_men_n876_), .A1(men_men_n115_), .B0(men_men_n430_), .Y(men_men_n877_));
  NA2        u0855(.A(men_men_n253_), .B(men_men_n47_), .Y(men_men_n878_));
  NA3        u0856(.A(men_men_n877_), .B(men_men_n875_), .C(men_men_n874_), .Y(men_men_n879_));
  NO4        u0857(.A(men_men_n879_), .B(men_men_n872_), .C(men_men_n867_), .D(men_men_n857_), .Y(men_men_n880_));
  NA4        u0858(.A(men_men_n880_), .B(men_men_n844_), .C(men_men_n838_), .D(men_men_n400_), .Y(men3));
  NA2        u0859(.A(i_6_), .B(i_7_), .Y(men_men_n882_));
  NO2        u0860(.A(men_men_n882_), .B(i_0_), .Y(men_men_n883_));
  NO2        u0861(.A(i_11_), .B(men_men_n245_), .Y(men_men_n884_));
  OAI210     u0862(.A0(men_men_n883_), .A1(men_men_n300_), .B0(men_men_n884_), .Y(men_men_n885_));
  NO2        u0863(.A(men_men_n885_), .B(men_men_n200_), .Y(men_men_n886_));
  NO3        u0864(.A(men_men_n477_), .B(men_men_n92_), .C(men_men_n45_), .Y(men_men_n887_));
  OA210      u0865(.A0(men_men_n887_), .A1(men_men_n886_), .B0(men_men_n180_), .Y(men_men_n888_));
  NA3        u0866(.A(men_men_n870_), .B(men_men_n637_), .C(men_men_n392_), .Y(men_men_n889_));
  NA2        u0867(.A(men_men_n889_), .B(men_men_n40_), .Y(men_men_n890_));
  NOi21      u0868(.An(men_men_n99_), .B(men_men_n801_), .Y(men_men_n891_));
  NO3        u0869(.A(men_men_n665_), .B(men_men_n481_), .C(men_men_n135_), .Y(men_men_n892_));
  NA2        u0870(.A(men_men_n433_), .B(men_men_n46_), .Y(men_men_n893_));
  AN2        u0871(.A(men_men_n479_), .B(men_men_n56_), .Y(men_men_n894_));
  NO3        u0872(.A(men_men_n894_), .B(men_men_n892_), .C(men_men_n891_), .Y(men_men_n895_));
  AOI210     u0873(.A0(men_men_n895_), .A1(men_men_n890_), .B0(men_men_n49_), .Y(men_men_n896_));
  NO4        u0874(.A(men_men_n396_), .B(men_men_n403_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n897_));
  NA2        u0875(.A(men_men_n192_), .B(men_men_n603_), .Y(men_men_n898_));
  NOi31      u0876(.An(men_men_n898_), .B(men_men_n897_), .C(men_men_n39_), .Y(men_men_n899_));
  NA2        u0877(.A(men_men_n748_), .B(men_men_n712_), .Y(men_men_n900_));
  NA2        u0878(.A(men_men_n347_), .B(men_men_n460_), .Y(men_men_n901_));
  OAI220     u0879(.A0(men_men_n901_), .A1(men_men_n900_), .B0(men_men_n899_), .B1(men_men_n64_), .Y(men_men_n902_));
  NOi21      u0880(.An(i_5_), .B(i_9_), .Y(men_men_n903_));
  NA2        u0881(.A(men_men_n903_), .B(men_men_n468_), .Y(men_men_n904_));
  AOI210     u0882(.A0(men_men_n275_), .A1(men_men_n502_), .B0(men_men_n727_), .Y(men_men_n905_));
  NO3        u0883(.A(men_men_n436_), .B(men_men_n275_), .C(men_men_n74_), .Y(men_men_n906_));
  NO2        u0884(.A(men_men_n181_), .B(men_men_n152_), .Y(men_men_n907_));
  AOI210     u0885(.A0(men_men_n907_), .A1(men_men_n253_), .B0(men_men_n906_), .Y(men_men_n908_));
  OAI220     u0886(.A0(men_men_n908_), .A1(men_men_n187_), .B0(men_men_n905_), .B1(men_men_n904_), .Y(men_men_n909_));
  NO4        u0887(.A(men_men_n909_), .B(men_men_n902_), .C(men_men_n896_), .D(men_men_n888_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n192_), .B(men_men_n24_), .Y(men_men_n911_));
  NO2        u0889(.A(men_men_n710_), .B(men_men_n626_), .Y(men_men_n912_));
  NO2        u0890(.A(men_men_n912_), .B(men_men_n911_), .Y(men_men_n913_));
  NA2        u0891(.A(men_men_n323_), .B(men_men_n133_), .Y(men_men_n914_));
  NAi21      u0892(.An(men_men_n167_), .B(men_men_n460_), .Y(men_men_n915_));
  OAI220     u0893(.A0(men_men_n915_), .A1(men_men_n878_), .B0(men_men_n914_), .B1(men_men_n421_), .Y(men_men_n916_));
  NO2        u0894(.A(men_men_n916_), .B(men_men_n913_), .Y(men_men_n917_));
  NO2        u0895(.A(men_men_n410_), .B(men_men_n304_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n918_), .B(men_men_n750_), .Y(men_men_n919_));
  NA2        u0897(.A(men_men_n604_), .B(i_0_), .Y(men_men_n920_));
  NO3        u0898(.A(men_men_n920_), .B(men_men_n405_), .C(men_men_n90_), .Y(men_men_n921_));
  NO4        u0899(.A(men_men_n620_), .B(men_men_n224_), .C(men_men_n439_), .D(men_men_n432_), .Y(men_men_n922_));
  AOI210     u0900(.A0(men_men_n922_), .A1(i_11_), .B0(men_men_n921_), .Y(men_men_n923_));
  INV        u0901(.A(men_men_n500_), .Y(men_men_n924_));
  AN2        u0902(.A(men_men_n99_), .B(men_men_n252_), .Y(men_men_n925_));
  NA2        u0903(.A(men_men_n788_), .B(men_men_n341_), .Y(men_men_n926_));
  AOI210     u0904(.A0(men_men_n510_), .A1(men_men_n90_), .B0(men_men_n59_), .Y(men_men_n927_));
  OAI220     u0905(.A0(men_men_n927_), .A1(men_men_n926_), .B0(men_men_n696_), .B1(men_men_n567_), .Y(men_men_n928_));
  NA2        u0906(.A(i_0_), .B(i_10_), .Y(men_men_n929_));
  OAI210     u0907(.A0(men_men_n929_), .A1(men_men_n87_), .B0(men_men_n570_), .Y(men_men_n930_));
  NO4        u0908(.A(men_men_n118_), .B(men_men_n59_), .C(men_men_n705_), .D(i_5_), .Y(men_men_n931_));
  AN2        u0909(.A(men_men_n931_), .B(men_men_n930_), .Y(men_men_n932_));
  AOI220     u0910(.A0(men_men_n347_), .A1(men_men_n101_), .B0(men_men_n192_), .B1(men_men_n85_), .Y(men_men_n933_));
  NA2        u0911(.A(men_men_n598_), .B(i_4_), .Y(men_men_n934_));
  NA2        u0912(.A(men_men_n195_), .B(men_men_n210_), .Y(men_men_n935_));
  OAI220     u0913(.A0(men_men_n935_), .A1(men_men_n926_), .B0(men_men_n934_), .B1(men_men_n933_), .Y(men_men_n936_));
  NO4        u0914(.A(men_men_n936_), .B(men_men_n932_), .C(men_men_n928_), .D(men_men_n925_), .Y(men_men_n937_));
  NA4        u0915(.A(men_men_n937_), .B(men_men_n923_), .C(men_men_n919_), .D(men_men_n917_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n106_), .B(men_men_n37_), .Y(men_men_n939_));
  NA2        u0917(.A(i_11_), .B(i_9_), .Y(men_men_n940_));
  NO3        u0918(.A(i_12_), .B(men_men_n940_), .C(men_men_n636_), .Y(men_men_n941_));
  AO220      u0919(.A0(men_men_n941_), .A1(men_men_n939_), .B0(men_men_n277_), .B1(men_men_n89_), .Y(men_men_n942_));
  NO2        u0920(.A(men_men_n49_), .B(i_7_), .Y(men_men_n943_));
  NA2        u0921(.A(men_men_n415_), .B(men_men_n185_), .Y(men_men_n944_));
  NA2        u0922(.A(men_men_n944_), .B(men_men_n165_), .Y(men_men_n945_));
  NO2        u0923(.A(men_men_n940_), .B(men_men_n74_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n181_), .B(i_0_), .Y(men_men_n947_));
  INV        u0925(.A(men_men_n947_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n500_), .B(men_men_n239_), .Y(men_men_n949_));
  AOI210     u0927(.A0(men_men_n391_), .A1(men_men_n42_), .B0(men_men_n429_), .Y(men_men_n950_));
  OAI220     u0928(.A0(men_men_n950_), .A1(men_men_n904_), .B0(men_men_n949_), .B1(men_men_n948_), .Y(men_men_n951_));
  NO3        u0929(.A(men_men_n951_), .B(men_men_n945_), .C(men_men_n942_), .Y(men_men_n952_));
  NA2        u0930(.A(men_men_n695_), .B(men_men_n125_), .Y(men_men_n953_));
  NO2        u0931(.A(i_6_), .B(men_men_n953_), .Y(men_men_n954_));
  AOI210     u0932(.A0(men_men_n471_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n955_));
  NA2        u0933(.A(men_men_n177_), .B(men_men_n106_), .Y(men_men_n956_));
  NOi32      u0934(.An(men_men_n955_), .Bn(men_men_n195_), .C(men_men_n956_), .Y(men_men_n957_));
  AOI210     u0935(.A0(men_men_n638_), .A1(men_men_n341_), .B0(men_men_n252_), .Y(men_men_n958_));
  NO2        u0936(.A(men_men_n958_), .B(men_men_n893_), .Y(men_men_n959_));
  NO3        u0937(.A(men_men_n959_), .B(men_men_n957_), .C(men_men_n954_), .Y(men_men_n960_));
  NOi21      u0938(.An(i_7_), .B(i_5_), .Y(men_men_n961_));
  NOi31      u0939(.An(men_men_n961_), .B(i_0_), .C(men_men_n765_), .Y(men_men_n962_));
  NA3        u0940(.A(men_men_n962_), .B(men_men_n404_), .C(i_6_), .Y(men_men_n963_));
  OA210      u0941(.A0(men_men_n956_), .A1(men_men_n545_), .B0(men_men_n963_), .Y(men_men_n964_));
  NO3        u0942(.A(men_men_n424_), .B(men_men_n380_), .C(men_men_n376_), .Y(men_men_n965_));
  NO2        u0943(.A(men_men_n269_), .B(men_men_n330_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n765_), .B(men_men_n266_), .Y(men_men_n967_));
  AOI210     u0945(.A0(men_men_n967_), .A1(men_men_n966_), .B0(men_men_n965_), .Y(men_men_n968_));
  NA4        u0946(.A(men_men_n968_), .B(men_men_n964_), .C(men_men_n960_), .D(men_men_n952_), .Y(men_men_n969_));
  NO2        u0947(.A(men_men_n911_), .B(men_men_n248_), .Y(men_men_n970_));
  AN2        u0948(.A(men_men_n346_), .B(men_men_n341_), .Y(men_men_n971_));
  AO220      u0949(.A0(men_men_n971_), .A1(men_men_n907_), .B0(men_men_n362_), .B1(men_men_n27_), .Y(men_men_n972_));
  OAI210     u0950(.A0(men_men_n972_), .A1(men_men_n970_), .B0(i_10_), .Y(men_men_n973_));
  OA210      u0951(.A0(men_men_n500_), .A1(men_men_n231_), .B0(men_men_n499_), .Y(men_men_n974_));
  NA3        u0952(.A(men_men_n499_), .B(men_men_n433_), .C(men_men_n46_), .Y(men_men_n975_));
  OAI210     u0953(.A0(men_men_n915_), .A1(men_men_n924_), .B0(men_men_n975_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n946_), .B(men_men_n316_), .Y(men_men_n977_));
  NA2        u0955(.A(men_men_n194_), .B(men_men_n977_), .Y(men_men_n978_));
  AOI220     u0956(.A0(men_men_n978_), .A1(men_men_n500_), .B0(men_men_n976_), .B1(men_men_n74_), .Y(men_men_n979_));
  NA3        u0957(.A(men_men_n859_), .B(men_men_n402_), .C(men_men_n674_), .Y(men_men_n980_));
  NA2        u0958(.A(men_men_n95_), .B(men_men_n45_), .Y(men_men_n981_));
  NO2        u0959(.A(men_men_n76_), .B(men_men_n790_), .Y(men_men_n982_));
  AOI220     u0960(.A0(men_men_n982_), .A1(men_men_n981_), .B0(men_men_n180_), .B1(men_men_n626_), .Y(men_men_n983_));
  AOI210     u0961(.A0(men_men_n983_), .A1(men_men_n980_), .B0(men_men_n48_), .Y(men_men_n984_));
  NO3        u0962(.A(men_men_n620_), .B(men_men_n375_), .C(men_men_n24_), .Y(men_men_n985_));
  INV        u0963(.A(men_men_n985_), .Y(men_men_n986_));
  NAi21      u0964(.An(i_9_), .B(i_5_), .Y(men_men_n987_));
  NO2        u0965(.A(men_men_n632_), .B(men_men_n108_), .Y(men_men_n988_));
  NA2        u0966(.A(men_men_n988_), .B(i_0_), .Y(men_men_n989_));
  OAI220     u0967(.A0(men_men_n989_), .A1(men_men_n87_), .B0(men_men_n986_), .B1(men_men_n178_), .Y(men_men_n990_));
  NO2        u0968(.A(men_men_n990_), .B(men_men_n984_), .Y(men_men_n991_));
  NA3        u0969(.A(men_men_n991_), .B(men_men_n979_), .C(men_men_n973_), .Y(men_men_n992_));
  NO3        u0970(.A(men_men_n992_), .B(men_men_n969_), .C(men_men_n938_), .Y(men_men_n993_));
  NO2        u0971(.A(i_0_), .B(men_men_n765_), .Y(men_men_n994_));
  NA2        u0972(.A(men_men_n74_), .B(men_men_n45_), .Y(men_men_n995_));
  NA2        u0973(.A(men_men_n929_), .B(men_men_n995_), .Y(men_men_n996_));
  NO3        u0974(.A(men_men_n108_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n997_));
  AO220      u0975(.A0(men_men_n997_), .A1(men_men_n996_), .B0(men_men_n994_), .B1(men_men_n180_), .Y(men_men_n998_));
  AOI210     u0976(.A0(men_men_n840_), .A1(men_men_n725_), .B0(men_men_n956_), .Y(men_men_n999_));
  AOI210     u0977(.A0(men_men_n998_), .A1(men_men_n364_), .B0(men_men_n999_), .Y(men_men_n1000_));
  NA2        u0978(.A(men_men_n776_), .B(men_men_n150_), .Y(men_men_n1001_));
  INV        u0979(.A(men_men_n1001_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n1002_), .B(men_men_n712_), .C(men_men_n74_), .Y(men_men_n1003_));
  NO2        u0981(.A(men_men_n855_), .B(men_men_n424_), .Y(men_men_n1004_));
  NA3        u0982(.A(men_men_n883_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n884_), .B(i_9_), .Y(men_men_n1006_));
  AOI210     u0984(.A0(men_men_n1005_), .A1(men_men_n526_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  OAI210     u0985(.A0(men_men_n253_), .A1(i_9_), .B0(men_men_n238_), .Y(men_men_n1008_));
  AOI210     u0986(.A0(men_men_n1008_), .A1(men_men_n920_), .B0(men_men_n158_), .Y(men_men_n1009_));
  NO3        u0987(.A(men_men_n1009_), .B(men_men_n1007_), .C(men_men_n1004_), .Y(men_men_n1010_));
  NA3        u0988(.A(men_men_n1010_), .B(men_men_n1003_), .C(men_men_n1000_), .Y(men_men_n1011_));
  NA2        u0989(.A(men_men_n971_), .B(men_men_n393_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n311_), .A1(men_men_n167_), .B0(men_men_n1012_), .Y(men_men_n1013_));
  NA3        u0991(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n1014_));
  NA2        u0992(.A(men_men_n943_), .B(men_men_n514_), .Y(men_men_n1015_));
  AOI210     u0993(.A0(men_men_n1014_), .A1(men_men_n167_), .B0(men_men_n1015_), .Y(men_men_n1016_));
  NO2        u0994(.A(men_men_n1016_), .B(men_men_n1013_), .Y(men_men_n1017_));
  NO3        u0995(.A(men_men_n929_), .B(men_men_n903_), .C(men_men_n197_), .Y(men_men_n1018_));
  AOI220     u0996(.A0(men_men_n1018_), .A1(i_11_), .B0(men_men_n599_), .B1(men_men_n76_), .Y(men_men_n1019_));
  NO3        u0997(.A(men_men_n218_), .B(men_men_n403_), .C(i_0_), .Y(men_men_n1020_));
  OAI210     u0998(.A0(men_men_n1020_), .A1(men_men_n77_), .B0(i_13_), .Y(men_men_n1021_));
  INV        u0999(.A(men_men_n227_), .Y(men_men_n1022_));
  OAI220     u1000(.A0(men_men_n560_), .A1(men_men_n143_), .B0(men_men_n679_), .B1(men_men_n649_), .Y(men_men_n1023_));
  NA3        u1001(.A(men_men_n1023_), .B(men_men_n419_), .C(men_men_n1022_), .Y(men_men_n1024_));
  NA4        u1002(.A(men_men_n1024_), .B(men_men_n1021_), .C(men_men_n1019_), .D(men_men_n1017_), .Y(men_men_n1025_));
  NO2        u1003(.A(men_men_n251_), .B(men_men_n95_), .Y(men_men_n1026_));
  AOI210     u1004(.A0(men_men_n1026_), .A1(men_men_n994_), .B0(men_men_n112_), .Y(men_men_n1027_));
  AOI220     u1005(.A0(men_men_n961_), .A1(men_men_n514_), .B0(men_men_n883_), .B1(men_men_n168_), .Y(men_men_n1028_));
  NA2        u1006(.A(men_men_n367_), .B(men_men_n182_), .Y(men_men_n1029_));
  OA220      u1007(.A0(men_men_n1029_), .A1(men_men_n1028_), .B0(men_men_n1027_), .B1(i_5_), .Y(men_men_n1030_));
  AOI210     u1008(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n181_), .Y(men_men_n1031_));
  NA2        u1009(.A(men_men_n1031_), .B(men_men_n974_), .Y(men_men_n1032_));
  NA3        u1010(.A(men_men_n646_), .B(men_men_n192_), .C(men_men_n85_), .Y(men_men_n1033_));
  NA2        u1011(.A(men_men_n1033_), .B(men_men_n577_), .Y(men_men_n1034_));
  NA2        u1012(.A(men_men_n519_), .B(men_men_n497_), .Y(men_men_n1035_));
  NO2        u1013(.A(men_men_n1035_), .B(men_men_n1034_), .Y(men_men_n1036_));
  NA3        u1014(.A(men_men_n410_), .B(men_men_n177_), .C(men_men_n176_), .Y(men_men_n1037_));
  NA3        u1015(.A(men_men_n943_), .B(men_men_n300_), .C(men_men_n238_), .Y(men_men_n1038_));
  NA2        u1016(.A(men_men_n1038_), .B(men_men_n1037_), .Y(men_men_n1039_));
  NA3        u1017(.A(men_men_n410_), .B(men_men_n348_), .C(men_men_n230_), .Y(men_men_n1040_));
  OAI210     u1018(.A0(men_men_n898_), .A1(men_men_n683_), .B0(men_men_n1040_), .Y(men_men_n1041_));
  NOi31      u1019(.An(men_men_n409_), .B(men_men_n995_), .C(men_men_n248_), .Y(men_men_n1042_));
  NO3        u1020(.A(men_men_n940_), .B(men_men_n227_), .C(men_men_n197_), .Y(men_men_n1043_));
  NO4        u1021(.A(men_men_n1043_), .B(men_men_n1042_), .C(men_men_n1041_), .D(men_men_n1039_), .Y(men_men_n1044_));
  NA4        u1022(.A(men_men_n1044_), .B(men_men_n1036_), .C(men_men_n1032_), .D(men_men_n1030_), .Y(men_men_n1045_));
  INV        u1023(.A(men_men_n648_), .Y(men_men_n1046_));
  NO3        u1024(.A(men_men_n1046_), .B(men_men_n589_), .C(men_men_n361_), .Y(men_men_n1047_));
  INV        u1025(.A(men_men_n1047_), .Y(men_men_n1048_));
  NA3        u1026(.A(men_men_n316_), .B(i_5_), .C(men_men_n200_), .Y(men_men_n1049_));
  NAi31      u1027(.An(men_men_n250_), .B(men_men_n1049_), .C(men_men_n251_), .Y(men_men_n1050_));
  NO4        u1028(.A(men_men_n248_), .B(men_men_n218_), .C(i_0_), .D(i_12_), .Y(men_men_n1051_));
  AOI220     u1029(.A0(men_men_n1051_), .A1(men_men_n1050_), .B0(men_men_n835_), .B1(men_men_n182_), .Y(men_men_n1052_));
  AN2        u1030(.A(men_men_n929_), .B(men_men_n158_), .Y(men_men_n1053_));
  NO4        u1031(.A(men_men_n1053_), .B(i_12_), .C(men_men_n683_), .D(men_men_n135_), .Y(men_men_n1054_));
  NA2        u1032(.A(men_men_n1054_), .B(men_men_n227_), .Y(men_men_n1055_));
  NA3        u1033(.A(men_men_n101_), .B(men_men_n603_), .C(i_11_), .Y(men_men_n1056_));
  NO2        u1034(.A(men_men_n1056_), .B(men_men_n160_), .Y(men_men_n1057_));
  NA2        u1035(.A(men_men_n65_), .B(men_men_n104_), .Y(men_men_n1058_));
  NO2        u1036(.A(men_men_n1058_), .B(men_men_n1049_), .Y(men_men_n1059_));
  AOI210     u1037(.A0(men_men_n1059_), .A1(men_men_n947_), .B0(men_men_n1057_), .Y(men_men_n1060_));
  NA4        u1038(.A(men_men_n1060_), .B(men_men_n1055_), .C(men_men_n1052_), .D(men_men_n1048_), .Y(men_men_n1061_));
  NO4        u1039(.A(men_men_n1061_), .B(men_men_n1045_), .C(men_men_n1025_), .D(men_men_n1011_), .Y(men_men_n1062_));
  OAI210     u1040(.A0(men_men_n858_), .A1(men_men_n851_), .B0(men_men_n37_), .Y(men_men_n1063_));
  NA3        u1041(.A(men_men_n955_), .B(men_men_n388_), .C(i_5_), .Y(men_men_n1064_));
  NA3        u1042(.A(men_men_n1064_), .B(men_men_n1063_), .C(men_men_n644_), .Y(men_men_n1065_));
  NA2        u1043(.A(men_men_n1065_), .B(men_men_n214_), .Y(men_men_n1066_));
  NA2        u1044(.A(men_men_n193_), .B(men_men_n195_), .Y(men_men_n1067_));
  AO210      u1045(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n1067_), .Y(men_men_n1068_));
  OAI210     u1046(.A0(men_men_n648_), .A1(men_men_n646_), .B0(men_men_n329_), .Y(men_men_n1069_));
  NAi31      u1047(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1070_));
  AOI210     u1048(.A0(men_men_n121_), .A1(men_men_n71_), .B0(men_men_n1070_), .Y(men_men_n1071_));
  NO2        u1049(.A(men_men_n1071_), .B(men_men_n680_), .Y(men_men_n1072_));
  NA3        u1050(.A(men_men_n1072_), .B(men_men_n1069_), .C(men_men_n1068_), .Y(men_men_n1073_));
  NO2        u1051(.A(men_men_n486_), .B(men_men_n275_), .Y(men_men_n1074_));
  NO4        u1052(.A(men_men_n241_), .B(men_men_n149_), .C(men_men_n716_), .D(men_men_n37_), .Y(men_men_n1075_));
  NO3        u1053(.A(men_men_n1075_), .B(men_men_n1074_), .C(men_men_n922_), .Y(men_men_n1076_));
  OAI210     u1054(.A0(men_men_n1056_), .A1(men_men_n152_), .B0(men_men_n1076_), .Y(men_men_n1077_));
  AOI210     u1055(.A0(men_men_n1073_), .A1(men_men_n49_), .B0(men_men_n1077_), .Y(men_men_n1078_));
  AOI210     u1056(.A0(men_men_n1078_), .A1(men_men_n1066_), .B0(men_men_n74_), .Y(men_men_n1079_));
  NO2        u1057(.A(men_men_n596_), .B(men_men_n399_), .Y(men_men_n1080_));
  NO2        u1058(.A(men_men_n1080_), .B(men_men_n796_), .Y(men_men_n1081_));
  INV        u1059(.A(men_men_n77_), .Y(men_men_n1082_));
  AOI210     u1060(.A0(men_men_n1031_), .A1(men_men_n943_), .B0(men_men_n962_), .Y(men_men_n1083_));
  AOI210     u1061(.A0(men_men_n1083_), .A1(men_men_n1082_), .B0(men_men_n716_), .Y(men_men_n1084_));
  NA2        u1062(.A(men_men_n269_), .B(men_men_n58_), .Y(men_men_n1085_));
  AOI220     u1063(.A0(men_men_n1085_), .A1(men_men_n77_), .B0(men_men_n362_), .B1(men_men_n263_), .Y(men_men_n1086_));
  NO2        u1064(.A(men_men_n1086_), .B(men_men_n245_), .Y(men_men_n1087_));
  NA3        u1065(.A(men_men_n99_), .B(men_men_n318_), .C(men_men_n31_), .Y(men_men_n1088_));
  INV        u1066(.A(men_men_n1088_), .Y(men_men_n1089_));
  NO3        u1067(.A(men_men_n1089_), .B(men_men_n1087_), .C(men_men_n1084_), .Y(men_men_n1090_));
  OAI210     u1068(.A0(men_men_n277_), .A1(men_men_n163_), .B0(men_men_n90_), .Y(men_men_n1091_));
  NA3        u1069(.A(men_men_n800_), .B(men_men_n300_), .C(men_men_n81_), .Y(men_men_n1092_));
  AOI210     u1070(.A0(men_men_n1092_), .A1(men_men_n1091_), .B0(i_11_), .Y(men_men_n1093_));
  NA2        u1071(.A(men_men_n639_), .B(men_men_n224_), .Y(men_men_n1094_));
  OAI210     u1072(.A0(men_men_n1094_), .A1(men_men_n955_), .B0(men_men_n214_), .Y(men_men_n1095_));
  NA2        u1073(.A(men_men_n169_), .B(i_5_), .Y(men_men_n1096_));
  AOI210     u1074(.A0(men_men_n1095_), .A1(men_men_n813_), .B0(men_men_n1096_), .Y(men_men_n1097_));
  NO3        u1075(.A(men_men_n60_), .B(men_men_n59_), .C(i_4_), .Y(men_men_n1098_));
  OAI210     u1076(.A0(men_men_n966_), .A1(men_men_n318_), .B0(men_men_n1098_), .Y(men_men_n1099_));
  NO2        u1077(.A(men_men_n1099_), .B(men_men_n765_), .Y(men_men_n1100_));
  NO4        u1078(.A(men_men_n987_), .B(men_men_n503_), .C(men_men_n262_), .D(men_men_n261_), .Y(men_men_n1101_));
  NO2        u1079(.A(men_men_n1101_), .B(men_men_n593_), .Y(men_men_n1102_));
  NO2        u1080(.A(men_men_n854_), .B(men_men_n381_), .Y(men_men_n1103_));
  AOI210     u1081(.A0(men_men_n1103_), .A1(men_men_n1102_), .B0(men_men_n41_), .Y(men_men_n1104_));
  NO4        u1082(.A(men_men_n1104_), .B(men_men_n1100_), .C(men_men_n1097_), .D(men_men_n1093_), .Y(men_men_n1105_));
  OAI210     u1083(.A0(men_men_n1090_), .A1(i_4_), .B0(men_men_n1105_), .Y(men_men_n1106_));
  NO3        u1084(.A(men_men_n1106_), .B(men_men_n1081_), .C(men_men_n1079_), .Y(men_men_n1107_));
  NA4        u1085(.A(men_men_n1107_), .B(men_men_n1062_), .C(men_men_n993_), .D(men_men_n910_), .Y(men4));
  INV        u1086(.A(men_men_n742_), .Y(men_men_n1111_));
  INV        u1087(.A(i_2_), .Y(men_men_n1112_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule