//Benchmark atmr_misex3_1774_0.0625

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  INV        o0001(.A(d), .Y(ori_ori_n30_));
  NA3        o0002(.A(e), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n31_));
  NOi32      o0003(.An(m), .Bn(l), .C(n), .Y(ori_ori_n32_));
  NOi32      o0004(.An(i), .Bn(o), .C(h), .Y(ori_ori_n33_));
  NA2        o0005(.A(ori_ori_n33_), .B(ori_ori_n32_), .Y(ori_ori_n34_));
  AN2        o0006(.A(m), .B(l), .Y(ori_ori_n35_));
  NOi32      o0007(.An(j), .Bn(o), .C(k), .Y(ori_ori_n36_));
  NA2        o0008(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n37_));
  NO2        o0009(.A(ori_ori_n37_), .B(n), .Y(ori_ori_n38_));
  INV        o0010(.A(h), .Y(ori_ori_n39_));
  NAi21      o0011(.An(j), .B(l), .Y(ori_ori_n40_));
  NAi32      o0012(.An(n), .Bn(o), .C(m), .Y(ori_ori_n41_));
  NO3        o0013(.A(ori_ori_n41_), .B(ori_ori_n40_), .C(ori_ori_n39_), .Y(ori_ori_n42_));
  NAi31      o0014(.An(n), .B(m), .C(l), .Y(ori_ori_n43_));
  INV        o0015(.A(i), .Y(ori_ori_n44_));
  AN2        o0016(.A(h), .B(o), .Y(ori_ori_n45_));
  NA2        o0017(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori_ori_n46_));
  NO2        o0018(.A(ori_ori_n46_), .B(ori_ori_n43_), .Y(ori_ori_n47_));
  NAi21      o0019(.An(n), .B(m), .Y(ori_ori_n48_));
  NOi32      o0020(.An(k), .Bn(h), .C(l), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(o), .Y(ori_ori_n50_));
  INV        o0022(.A(ori_ori_n50_), .Y(ori_ori_n51_));
  NO2        o0023(.A(ori_ori_n51_), .B(ori_ori_n48_), .Y(ori_ori_n52_));
  NO3        o0024(.A(ori_ori_n52_), .B(ori_ori_n47_), .C(ori_ori_n42_), .Y(ori_ori_n53_));
  AOI210     o0025(.A0(ori_ori_n53_), .A1(ori_ori_n34_), .B0(ori_ori_n31_), .Y(ori_ori_n54_));
  INV        o0026(.A(c), .Y(ori_ori_n55_));
  NA2        o0027(.A(e), .B(b), .Y(ori_ori_n56_));
  NO2        o0028(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  INV        o0029(.A(d), .Y(ori_ori_n58_));
  NAi21      o0030(.An(i), .B(h), .Y(ori_ori_n59_));
  NAi41      o0031(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n60_));
  NA2        o0032(.A(o), .B(f), .Y(ori_ori_n61_));
  NAi21      o0033(.An(i), .B(j), .Y(ori_ori_n62_));
  NAi32      o0034(.An(n), .Bn(k), .C(m), .Y(ori_ori_n63_));
  NAi31      o0035(.An(l), .B(m), .C(k), .Y(ori_ori_n64_));
  NAi21      o0036(.An(e), .B(h), .Y(ori_ori_n65_));
  NAi41      o0037(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n66_));
  INV        o0038(.A(m), .Y(ori_ori_n67_));
  NOi21      o0039(.An(k), .B(l), .Y(ori_ori_n68_));
  NA2        o0040(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  AN4        o0041(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n70_));
  NOi21      o0042(.An(h), .B(f), .Y(ori_ori_n71_));
  NA2        o0043(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n72_));
  NAi32      o0044(.An(m), .Bn(k), .C(j), .Y(ori_ori_n73_));
  NOi32      o0045(.An(h), .Bn(o), .C(f), .Y(ori_ori_n74_));
  OR2        o0046(.A(ori_ori_n72_), .B(ori_ori_n69_), .Y(ori_ori_n75_));
  INV        o0047(.A(ori_ori_n75_), .Y(ori_ori_n76_));
  INV        o0048(.A(n), .Y(ori_ori_n77_));
  AN2        o0049(.A(e), .B(b), .Y(ori_ori_n78_));
  NA2        o0050(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  INV        o0051(.A(j), .Y(ori_ori_n80_));
  AN3        o0052(.A(m), .B(k), .C(i), .Y(ori_ori_n81_));
  NA3        o0053(.A(ori_ori_n81_), .B(ori_ori_n80_), .C(o), .Y(ori_ori_n82_));
  NO2        o0054(.A(ori_ori_n82_), .B(f), .Y(ori_ori_n83_));
  NAi32      o0055(.An(o), .Bn(f), .C(h), .Y(ori_ori_n84_));
  NAi31      o0056(.An(j), .B(m), .C(l), .Y(ori_ori_n85_));
  NO2        o0057(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  NA2        o0058(.A(m), .B(l), .Y(ori_ori_n87_));
  NAi31      o0059(.An(k), .B(j), .C(o), .Y(ori_ori_n88_));
  NO3        o0060(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(f), .Y(ori_ori_n89_));
  AN2        o0061(.A(j), .B(o), .Y(ori_ori_n90_));
  NOi32      o0062(.An(m), .Bn(l), .C(i), .Y(ori_ori_n91_));
  NOi21      o0063(.An(o), .B(i), .Y(ori_ori_n92_));
  NOi32      o0064(.An(m), .Bn(j), .C(k), .Y(ori_ori_n93_));
  AOI220     o0065(.A0(ori_ori_n93_), .A1(ori_ori_n92_), .B0(ori_ori_n91_), .B1(ori_ori_n90_), .Y(ori_ori_n94_));
  NO2        o0066(.A(ori_ori_n94_), .B(f), .Y(ori_ori_n95_));
  NAi41      o0067(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n96_));
  AN2        o0068(.A(e), .B(b), .Y(ori_ori_n97_));
  NOi21      o0069(.An(i), .B(h), .Y(ori_ori_n98_));
  INV        o0070(.A(a), .Y(ori_ori_n99_));
  NA2        o0071(.A(ori_ori_n97_), .B(ori_ori_n99_), .Y(ori_ori_n100_));
  INV        o0072(.A(l), .Y(ori_ori_n101_));
  NOi21      o0073(.An(m), .B(n), .Y(ori_ori_n102_));
  AN2        o0074(.A(k), .B(h), .Y(ori_ori_n103_));
  INV        o0075(.A(b), .Y(ori_ori_n104_));
  NA2        o0076(.A(l), .B(j), .Y(ori_ori_n105_));
  AN2        o0077(.A(k), .B(i), .Y(ori_ori_n106_));
  NA2        o0078(.A(ori_ori_n106_), .B(ori_ori_n105_), .Y(ori_ori_n107_));
  NA2        o0079(.A(o), .B(e), .Y(ori_ori_n108_));
  NOi32      o0080(.An(c), .Bn(a), .C(d), .Y(ori_ori_n109_));
  NA2        o0081(.A(ori_ori_n109_), .B(ori_ori_n102_), .Y(ori_ori_n110_));
  NO2        o0082(.A(ori_ori_n1155_), .B(ori_ori_n79_), .Y(ori_ori_n111_));
  NOi31      o0083(.An(k), .B(m), .C(j), .Y(ori_ori_n112_));
  NA3        o0084(.A(ori_ori_n112_), .B(ori_ori_n71_), .C(ori_ori_n70_), .Y(ori_ori_n113_));
  NOi31      o0085(.An(k), .B(m), .C(i), .Y(ori_ori_n114_));
  INV        o0086(.A(ori_ori_n113_), .Y(ori_ori_n115_));
  NOi32      o0087(.An(f), .Bn(b), .C(e), .Y(ori_ori_n116_));
  NAi21      o0088(.An(o), .B(h), .Y(ori_ori_n117_));
  NAi21      o0089(.An(m), .B(n), .Y(ori_ori_n118_));
  NAi41      o0090(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n119_));
  NAi31      o0091(.An(j), .B(k), .C(h), .Y(ori_ori_n120_));
  NO2        o0092(.A(k), .B(j), .Y(ori_ori_n121_));
  NO2        o0093(.A(ori_ori_n121_), .B(ori_ori_n118_), .Y(ori_ori_n122_));
  AN2        o0094(.A(k), .B(j), .Y(ori_ori_n123_));
  NAi21      o0095(.An(c), .B(b), .Y(ori_ori_n124_));
  NA2        o0096(.A(f), .B(d), .Y(ori_ori_n125_));
  NO4        o0097(.A(ori_ori_n125_), .B(ori_ori_n124_), .C(ori_ori_n123_), .D(ori_ori_n117_), .Y(ori_ori_n126_));
  NA2        o0098(.A(h), .B(c), .Y(ori_ori_n127_));
  NAi31      o0099(.An(f), .B(e), .C(b), .Y(ori_ori_n128_));
  NA2        o0100(.A(ori_ori_n126_), .B(ori_ori_n122_), .Y(ori_ori_n129_));
  NA2        o0101(.A(d), .B(b), .Y(ori_ori_n130_));
  NAi21      o0102(.An(e), .B(f), .Y(ori_ori_n131_));
  NO2        o0103(.A(ori_ori_n131_), .B(ori_ori_n130_), .Y(ori_ori_n132_));
  NA2        o0104(.A(b), .B(a), .Y(ori_ori_n133_));
  NAi21      o0105(.An(e), .B(o), .Y(ori_ori_n134_));
  NAi21      o0106(.An(c), .B(d), .Y(ori_ori_n135_));
  NAi31      o0107(.An(l), .B(k), .C(h), .Y(ori_ori_n136_));
  NO2        o0108(.A(ori_ori_n118_), .B(ori_ori_n136_), .Y(ori_ori_n137_));
  NA2        o0109(.A(ori_ori_n137_), .B(ori_ori_n132_), .Y(ori_ori_n138_));
  NAi31      o0110(.An(ori_ori_n115_), .B(ori_ori_n138_), .C(ori_ori_n129_), .Y(ori_ori_n139_));
  NAi31      o0111(.An(e), .B(f), .C(b), .Y(ori_ori_n140_));
  NOi21      o0112(.An(o), .B(d), .Y(ori_ori_n141_));
  NO2        o0113(.A(ori_ori_n141_), .B(ori_ori_n140_), .Y(ori_ori_n142_));
  NOi21      o0114(.An(h), .B(i), .Y(ori_ori_n143_));
  NOi21      o0115(.An(k), .B(m), .Y(ori_ori_n144_));
  NA3        o0116(.A(ori_ori_n144_), .B(ori_ori_n143_), .C(n), .Y(ori_ori_n145_));
  NOi21      o0117(.An(ori_ori_n142_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NOi21      o0118(.An(h), .B(o), .Y(ori_ori_n147_));
  NAi31      o0119(.An(l), .B(j), .C(h), .Y(ori_ori_n148_));
  NAi31      o0120(.An(d), .B(f), .C(c), .Y(ori_ori_n149_));
  NAi31      o0121(.An(e), .B(f), .C(c), .Y(ori_ori_n150_));
  NA2        o0122(.A(ori_ori_n150_), .B(ori_ori_n149_), .Y(ori_ori_n151_));
  NA2        o0123(.A(j), .B(h), .Y(ori_ori_n152_));
  OR3        o0124(.A(n), .B(m), .C(k), .Y(ori_ori_n153_));
  NO2        o0125(.A(ori_ori_n153_), .B(ori_ori_n152_), .Y(ori_ori_n154_));
  NAi32      o0126(.An(m), .Bn(k), .C(n), .Y(ori_ori_n155_));
  NO2        o0127(.A(ori_ori_n155_), .B(ori_ori_n152_), .Y(ori_ori_n156_));
  AOI220     o0128(.A0(ori_ori_n156_), .A1(ori_ori_n142_), .B0(ori_ori_n154_), .B1(ori_ori_n151_), .Y(ori_ori_n157_));
  NO2        o0129(.A(n), .B(m), .Y(ori_ori_n158_));
  NA2        o0130(.A(ori_ori_n158_), .B(ori_ori_n49_), .Y(ori_ori_n159_));
  NAi21      o0131(.An(f), .B(e), .Y(ori_ori_n160_));
  NA2        o0132(.A(d), .B(c), .Y(ori_ori_n161_));
  NO2        o0133(.A(ori_ori_n161_), .B(ori_ori_n160_), .Y(ori_ori_n162_));
  NOi21      o0134(.An(ori_ori_n162_), .B(ori_ori_n159_), .Y(ori_ori_n163_));
  NAi31      o0135(.An(m), .B(n), .C(b), .Y(ori_ori_n164_));
  NAi21      o0136(.An(h), .B(f), .Y(ori_ori_n165_));
  NO2        o0137(.A(ori_ori_n164_), .B(ori_ori_n135_), .Y(ori_ori_n166_));
  NOi32      o0138(.An(f), .Bn(c), .C(d), .Y(ori_ori_n167_));
  NOi32      o0139(.An(f), .Bn(c), .C(e), .Y(ori_ori_n168_));
  NO2        o0140(.A(ori_ori_n168_), .B(ori_ori_n167_), .Y(ori_ori_n169_));
  NO3        o0141(.A(n), .B(m), .C(j), .Y(ori_ori_n170_));
  NA2        o0142(.A(ori_ori_n170_), .B(ori_ori_n103_), .Y(ori_ori_n171_));
  AO210      o0143(.A0(ori_ori_n171_), .A1(ori_ori_n159_), .B0(ori_ori_n169_), .Y(ori_ori_n172_));
  NAi31      o0144(.An(ori_ori_n163_), .B(ori_ori_n172_), .C(ori_ori_n157_), .Y(ori_ori_n173_));
  OR3        o0145(.A(ori_ori_n173_), .B(ori_ori_n146_), .C(ori_ori_n139_), .Y(ori_ori_n174_));
  NO4        o0146(.A(ori_ori_n174_), .B(ori_ori_n111_), .C(ori_ori_n76_), .D(ori_ori_n54_), .Y(ori_ori_n175_));
  NA3        o0147(.A(m), .B(ori_ori_n101_), .C(j), .Y(ori_ori_n176_));
  NAi31      o0148(.An(n), .B(h), .C(o), .Y(ori_ori_n177_));
  NO2        o0149(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  NOi32      o0150(.An(m), .Bn(k), .C(l), .Y(ori_ori_n179_));
  NA3        o0151(.A(ori_ori_n179_), .B(ori_ori_n80_), .C(o), .Y(ori_ori_n180_));
  NO2        o0152(.A(ori_ori_n180_), .B(n), .Y(ori_ori_n181_));
  NOi21      o0153(.An(k), .B(j), .Y(ori_ori_n182_));
  NA4        o0154(.A(ori_ori_n182_), .B(ori_ori_n102_), .C(i), .D(o), .Y(ori_ori_n183_));
  AN2        o0155(.A(i), .B(o), .Y(ori_ori_n184_));
  NA3        o0156(.A(ori_ori_n68_), .B(ori_ori_n184_), .C(ori_ori_n102_), .Y(ori_ori_n185_));
  NA2        o0157(.A(ori_ori_n185_), .B(ori_ori_n183_), .Y(ori_ori_n186_));
  NO3        o0158(.A(ori_ori_n186_), .B(ori_ori_n181_), .C(ori_ori_n178_), .Y(ori_ori_n187_));
  NAi41      o0159(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n188_));
  INV        o0160(.A(ori_ori_n188_), .Y(ori_ori_n189_));
  INV        o0161(.A(f), .Y(ori_ori_n190_));
  INV        o0162(.A(o), .Y(ori_ori_n191_));
  NOi31      o0163(.An(i), .B(j), .C(h), .Y(ori_ori_n192_));
  NOi21      o0164(.An(l), .B(m), .Y(ori_ori_n193_));
  NA2        o0165(.A(ori_ori_n193_), .B(ori_ori_n192_), .Y(ori_ori_n194_));
  NO3        o0166(.A(ori_ori_n194_), .B(ori_ori_n191_), .C(ori_ori_n190_), .Y(ori_ori_n195_));
  NA2        o0167(.A(ori_ori_n195_), .B(ori_ori_n189_), .Y(ori_ori_n196_));
  OAI210     o0168(.A0(ori_ori_n187_), .A1(ori_ori_n31_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  NOi21      o0169(.An(n), .B(m), .Y(ori_ori_n198_));
  OR2        o0170(.A(ori_ori_n73_), .B(ori_ori_n72_), .Y(ori_ori_n199_));
  NAi21      o0171(.An(j), .B(h), .Y(ori_ori_n200_));
  XN2        o0172(.A(i), .B(h), .Y(ori_ori_n201_));
  NA2        o0173(.A(ori_ori_n201_), .B(ori_ori_n200_), .Y(ori_ori_n202_));
  NOi31      o0174(.An(k), .B(n), .C(m), .Y(ori_ori_n203_));
  NOi31      o0175(.An(ori_ori_n203_), .B(ori_ori_n161_), .C(ori_ori_n160_), .Y(ori_ori_n204_));
  NA2        o0176(.A(ori_ori_n204_), .B(ori_ori_n202_), .Y(ori_ori_n205_));
  NAi31      o0177(.An(f), .B(e), .C(c), .Y(ori_ori_n206_));
  NO4        o0178(.A(ori_ori_n206_), .B(ori_ori_n153_), .C(ori_ori_n152_), .D(ori_ori_n58_), .Y(ori_ori_n207_));
  NAi32      o0179(.An(m), .Bn(i), .C(k), .Y(ori_ori_n208_));
  INV        o0180(.A(k), .Y(ori_ori_n209_));
  INV        o0181(.A(ori_ori_n207_), .Y(ori_ori_n210_));
  NAi21      o0182(.An(n), .B(a), .Y(ori_ori_n211_));
  NO2        o0183(.A(ori_ori_n211_), .B(ori_ori_n130_), .Y(ori_ori_n212_));
  NAi41      o0184(.An(o), .B(m), .C(k), .D(h), .Y(ori_ori_n213_));
  NO2        o0185(.A(ori_ori_n213_), .B(e), .Y(ori_ori_n214_));
  NA2        o0186(.A(ori_ori_n214_), .B(ori_ori_n212_), .Y(ori_ori_n215_));
  AN4        o0187(.A(ori_ori_n215_), .B(ori_ori_n210_), .C(ori_ori_n205_), .D(ori_ori_n199_), .Y(ori_ori_n216_));
  NO2        o0188(.A(h), .B(ori_ori_n96_), .Y(ori_ori_n217_));
  NA2        o0189(.A(ori_ori_n217_), .B(ori_ori_n116_), .Y(ori_ori_n218_));
  NAi41      o0190(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n219_));
  NO2        o0191(.A(ori_ori_n219_), .B(ori_ori_n190_), .Y(ori_ori_n220_));
  NA2        o0192(.A(ori_ori_n144_), .B(ori_ori_n98_), .Y(ori_ori_n221_));
  NAi21      o0193(.An(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NO2        o0194(.A(n), .B(a), .Y(ori_ori_n223_));
  NAi31      o0195(.An(ori_ori_n213_), .B(ori_ori_n223_), .C(ori_ori_n97_), .Y(ori_ori_n224_));
  AN2        o0196(.A(ori_ori_n224_), .B(ori_ori_n222_), .Y(ori_ori_n225_));
  NAi21      o0197(.An(h), .B(i), .Y(ori_ori_n226_));
  NA2        o0198(.A(ori_ori_n158_), .B(k), .Y(ori_ori_n227_));
  NO2        o0199(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  NA2        o0200(.A(ori_ori_n228_), .B(ori_ori_n167_), .Y(ori_ori_n229_));
  NA3        o0201(.A(ori_ori_n229_), .B(ori_ori_n225_), .C(ori_ori_n218_), .Y(ori_ori_n230_));
  NOi21      o0202(.An(o), .B(e), .Y(ori_ori_n231_));
  NO2        o0203(.A(ori_ori_n66_), .B(ori_ori_n67_), .Y(ori_ori_n232_));
  NA2        o0204(.A(ori_ori_n232_), .B(ori_ori_n231_), .Y(ori_ori_n233_));
  NOi32      o0205(.An(l), .Bn(j), .C(i), .Y(ori_ori_n234_));
  AOI210     o0206(.A0(ori_ori_n68_), .A1(ori_ori_n80_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  NAi21      o0207(.An(f), .B(o), .Y(ori_ori_n236_));
  NO2        o0208(.A(ori_ori_n236_), .B(ori_ori_n60_), .Y(ori_ori_n237_));
  NO2        o0209(.A(ori_ori_n235_), .B(ori_ori_n233_), .Y(ori_ori_n238_));
  NOi41      o0210(.An(ori_ori_n216_), .B(ori_ori_n238_), .C(ori_ori_n230_), .D(ori_ori_n197_), .Y(ori_ori_n239_));
  NO4        o0211(.A(ori_ori_n178_), .B(ori_ori_n47_), .C(ori_ori_n42_), .D(ori_ori_n38_), .Y(ori_ori_n240_));
  NO2        o0212(.A(ori_ori_n240_), .B(ori_ori_n100_), .Y(ori_ori_n241_));
  NA3        o0213(.A(ori_ori_n58_), .B(c), .C(b), .Y(ori_ori_n242_));
  NO2        o0214(.A(ori_ori_n221_), .B(ori_ori_n236_), .Y(ori_ori_n243_));
  NAi31      o0215(.An(o), .B(k), .C(h), .Y(ori_ori_n244_));
  NA3        o0216(.A(ori_ori_n144_), .B(ori_ori_n143_), .C(ori_ori_n77_), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(ori_ori_n169_), .Y(ori_ori_n246_));
  INV        o0218(.A(ori_ori_n246_), .Y(ori_ori_n247_));
  NA3        o0219(.A(e), .B(c), .C(b), .Y(ori_ori_n248_));
  NAi32      o0220(.An(k), .Bn(i), .C(j), .Y(ori_ori_n249_));
  NAi31      o0221(.An(h), .B(l), .C(i), .Y(ori_ori_n250_));
  NA3        o0222(.A(ori_ori_n250_), .B(ori_ori_n249_), .C(ori_ori_n148_), .Y(ori_ori_n251_));
  NOi21      o0223(.An(ori_ori_n251_), .B(ori_ori_n48_), .Y(ori_ori_n252_));
  NA2        o0224(.A(ori_ori_n237_), .B(ori_ori_n252_), .Y(ori_ori_n253_));
  NAi21      o0225(.An(l), .B(k), .Y(ori_ori_n254_));
  NO2        o0226(.A(ori_ori_n254_), .B(ori_ori_n48_), .Y(ori_ori_n255_));
  NOi21      o0227(.An(l), .B(j), .Y(ori_ori_n256_));
  NA2        o0228(.A(ori_ori_n147_), .B(ori_ori_n256_), .Y(ori_ori_n257_));
  NAi32      o0229(.An(j), .Bn(h), .C(i), .Y(ori_ori_n258_));
  NAi21      o0230(.An(m), .B(l), .Y(ori_ori_n259_));
  NA2        o0231(.A(h), .B(o), .Y(ori_ori_n260_));
  NA2        o0232(.A(ori_ori_n253_), .B(ori_ori_n247_), .Y(ori_ori_n261_));
  NO2        o0233(.A(ori_ori_n128_), .B(d), .Y(ori_ori_n262_));
  NAi32      o0234(.An(n), .Bn(m), .C(l), .Y(ori_ori_n263_));
  NO2        o0235(.A(ori_ori_n263_), .B(ori_ori_n258_), .Y(ori_ori_n264_));
  NA2        o0236(.A(ori_ori_n264_), .B(ori_ori_n162_), .Y(ori_ori_n265_));
  NAi31      o0237(.An(k), .B(l), .C(j), .Y(ori_ori_n266_));
  OAI210     o0238(.A0(ori_ori_n254_), .A1(j), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  NOi21      o0239(.An(ori_ori_n267_), .B(ori_ori_n108_), .Y(ori_ori_n268_));
  NO3        o0240(.A(ori_ori_n1154_), .B(ori_ori_n261_), .C(ori_ori_n241_), .Y(ori_ori_n269_));
  NA2        o0241(.A(ori_ori_n228_), .B(ori_ori_n168_), .Y(ori_ori_n270_));
  NAi21      o0242(.An(m), .B(k), .Y(ori_ori_n271_));
  NO2        o0243(.A(ori_ori_n201_), .B(ori_ori_n271_), .Y(ori_ori_n272_));
  NAi41      o0244(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n273_));
  NO2        o0245(.A(ori_ori_n273_), .B(ori_ori_n134_), .Y(ori_ori_n274_));
  NA2        o0246(.A(ori_ori_n274_), .B(ori_ori_n272_), .Y(ori_ori_n275_));
  NA2        o0247(.A(e), .B(c), .Y(ori_ori_n276_));
  NO3        o0248(.A(ori_ori_n276_), .B(n), .C(d), .Y(ori_ori_n277_));
  NOi21      o0249(.An(f), .B(h), .Y(ori_ori_n278_));
  NA2        o0250(.A(ori_ori_n278_), .B(ori_ori_n106_), .Y(ori_ori_n279_));
  NO2        o0251(.A(ori_ori_n279_), .B(ori_ori_n191_), .Y(ori_ori_n280_));
  NAi31      o0252(.An(d), .B(e), .C(b), .Y(ori_ori_n281_));
  NA2        o0253(.A(ori_ori_n275_), .B(ori_ori_n270_), .Y(ori_ori_n282_));
  NO4        o0254(.A(ori_ori_n273_), .B(ori_ori_n73_), .C(ori_ori_n65_), .D(ori_ori_n191_), .Y(ori_ori_n283_));
  NA2        o0255(.A(ori_ori_n223_), .B(ori_ori_n97_), .Y(ori_ori_n284_));
  NOi31      o0256(.An(l), .B(n), .C(m), .Y(ori_ori_n285_));
  NA2        o0257(.A(ori_ori_n285_), .B(ori_ori_n192_), .Y(ori_ori_n286_));
  NO2        o0258(.A(ori_ori_n286_), .B(ori_ori_n169_), .Y(ori_ori_n287_));
  OR2        o0259(.A(ori_ori_n287_), .B(ori_ori_n283_), .Y(ori_ori_n288_));
  NAi32      o0260(.An(m), .Bn(j), .C(k), .Y(ori_ori_n289_));
  NAi41      o0261(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n290_));
  NOi31      o0262(.An(j), .B(m), .C(k), .Y(ori_ori_n291_));
  NO2        o0263(.A(ori_ori_n112_), .B(ori_ori_n291_), .Y(ori_ori_n292_));
  AN3        o0264(.A(h), .B(o), .C(f), .Y(ori_ori_n293_));
  NOi32      o0265(.An(m), .Bn(j), .C(l), .Y(ori_ori_n294_));
  NO2        o0266(.A(ori_ori_n259_), .B(ori_ori_n258_), .Y(ori_ori_n295_));
  NO2        o0267(.A(ori_ori_n194_), .B(o), .Y(ori_ori_n296_));
  NO2        o0268(.A(ori_ori_n140_), .B(ori_ori_n77_), .Y(ori_ori_n297_));
  AOI220     o0269(.A0(ori_ori_n297_), .A1(ori_ori_n296_), .B0(ori_ori_n220_), .B1(ori_ori_n295_), .Y(ori_ori_n298_));
  INV        o0270(.A(ori_ori_n298_), .Y(ori_ori_n299_));
  NA3        o0271(.A(h), .B(o), .C(f), .Y(ori_ori_n300_));
  NO2        o0272(.A(ori_ori_n300_), .B(ori_ori_n69_), .Y(ori_ori_n301_));
  NA2        o0273(.A(ori_ori_n290_), .B(ori_ori_n188_), .Y(ori_ori_n302_));
  NA2        o0274(.A(ori_ori_n147_), .B(e), .Y(ori_ori_n303_));
  NO2        o0275(.A(ori_ori_n303_), .B(ori_ori_n40_), .Y(ori_ori_n304_));
  NA2        o0276(.A(ori_ori_n302_), .B(ori_ori_n301_), .Y(ori_ori_n305_));
  NOi32      o0277(.An(j), .Bn(o), .C(i), .Y(ori_ori_n306_));
  NA3        o0278(.A(ori_ori_n306_), .B(ori_ori_n254_), .C(ori_ori_n102_), .Y(ori_ori_n307_));
  AO210      o0279(.A0(ori_ori_n100_), .A1(ori_ori_n31_), .B0(ori_ori_n307_), .Y(ori_ori_n308_));
  NOi32      o0280(.An(e), .Bn(b), .C(a), .Y(ori_ori_n309_));
  AN2        o0281(.A(l), .B(j), .Y(ori_ori_n310_));
  NA3        o0282(.A(ori_ori_n185_), .B(ori_ori_n183_), .C(ori_ori_n34_), .Y(ori_ori_n311_));
  NA2        o0283(.A(ori_ori_n311_), .B(ori_ori_n309_), .Y(ori_ori_n312_));
  NA2        o0284(.A(ori_ori_n184_), .B(k), .Y(ori_ori_n313_));
  NA3        o0285(.A(m), .B(ori_ori_n101_), .C(ori_ori_n190_), .Y(ori_ori_n314_));
  NA4        o0286(.A(ori_ori_n179_), .B(ori_ori_n80_), .C(o), .D(ori_ori_n190_), .Y(ori_ori_n315_));
  NA2        o0287(.A(ori_ori_n50_), .B(ori_ori_n102_), .Y(ori_ori_n316_));
  NA3        o0288(.A(ori_ori_n312_), .B(ori_ori_n308_), .C(ori_ori_n305_), .Y(ori_ori_n317_));
  NO4        o0289(.A(ori_ori_n317_), .B(ori_ori_n299_), .C(ori_ori_n288_), .D(ori_ori_n282_), .Y(ori_ori_n318_));
  NA4        o0290(.A(ori_ori_n318_), .B(ori_ori_n269_), .C(ori_ori_n239_), .D(ori_ori_n175_), .Y(ori10));
  NA3        o0291(.A(m), .B(k), .C(i), .Y(ori_ori_n320_));
  NOi21      o0292(.An(e), .B(f), .Y(ori_ori_n321_));
  NAi31      o0293(.An(b), .B(f), .C(c), .Y(ori_ori_n322_));
  INV        o0294(.A(ori_ori_n322_), .Y(ori_ori_n323_));
  NOi32      o0295(.An(k), .Bn(h), .C(j), .Y(ori_ori_n324_));
  NA2        o0296(.A(ori_ori_n324_), .B(ori_ori_n198_), .Y(ori_ori_n325_));
  NA2        o0297(.A(ori_ori_n145_), .B(ori_ori_n325_), .Y(ori_ori_n326_));
  NA2        o0298(.A(ori_ori_n326_), .B(ori_ori_n323_), .Y(ori_ori_n327_));
  AN2        o0299(.A(j), .B(h), .Y(ori_ori_n328_));
  NO3        o0300(.A(n), .B(m), .C(k), .Y(ori_ori_n329_));
  NA2        o0301(.A(ori_ori_n329_), .B(ori_ori_n328_), .Y(ori_ori_n330_));
  NO3        o0302(.A(ori_ori_n330_), .B(ori_ori_n135_), .C(ori_ori_n190_), .Y(ori_ori_n331_));
  OR2        o0303(.A(m), .B(k), .Y(ori_ori_n332_));
  NO2        o0304(.A(ori_ori_n152_), .B(ori_ori_n332_), .Y(ori_ori_n333_));
  NA4        o0305(.A(n), .B(f), .C(c), .D(ori_ori_n104_), .Y(ori_ori_n334_));
  NOi21      o0306(.An(ori_ori_n333_), .B(ori_ori_n334_), .Y(ori_ori_n335_));
  NOi32      o0307(.An(d), .Bn(a), .C(c), .Y(ori_ori_n336_));
  NA2        o0308(.A(ori_ori_n336_), .B(ori_ori_n160_), .Y(ori_ori_n337_));
  NAi21      o0309(.An(i), .B(o), .Y(ori_ori_n338_));
  NAi31      o0310(.An(k), .B(m), .C(j), .Y(ori_ori_n339_));
  NO3        o0311(.A(ori_ori_n339_), .B(ori_ori_n338_), .C(n), .Y(ori_ori_n340_));
  NOi21      o0312(.An(ori_ori_n340_), .B(ori_ori_n337_), .Y(ori_ori_n341_));
  NO3        o0313(.A(ori_ori_n341_), .B(ori_ori_n335_), .C(ori_ori_n331_), .Y(ori_ori_n342_));
  NO2        o0314(.A(ori_ori_n334_), .B(ori_ori_n259_), .Y(ori_ori_n343_));
  NOi32      o0315(.An(f), .Bn(d), .C(c), .Y(ori_ori_n344_));
  AOI220     o0316(.A0(ori_ori_n344_), .A1(ori_ori_n264_), .B0(ori_ori_n343_), .B1(ori_ori_n192_), .Y(ori_ori_n345_));
  NA3        o0317(.A(ori_ori_n345_), .B(ori_ori_n342_), .C(ori_ori_n327_), .Y(ori_ori_n346_));
  NO2        o0318(.A(ori_ori_n58_), .B(ori_ori_n104_), .Y(ori_ori_n347_));
  NA2        o0319(.A(ori_ori_n223_), .B(ori_ori_n347_), .Y(ori_ori_n348_));
  INV        o0320(.A(e), .Y(ori_ori_n349_));
  NO2        o0321(.A(ori_ori_n82_), .B(ori_ori_n349_), .Y(ori_ori_n350_));
  INV        o0322(.A(ori_ori_n350_), .Y(ori_ori_n351_));
  NOi21      o0323(.An(o), .B(h), .Y(ori_ori_n352_));
  AN3        o0324(.A(m), .B(l), .C(i), .Y(ori_ori_n353_));
  AN3        o0325(.A(h), .B(o), .C(e), .Y(ori_ori_n354_));
  NO2        o0326(.A(ori_ori_n351_), .B(ori_ori_n348_), .Y(ori_ori_n355_));
  NA3        o0327(.A(ori_ori_n36_), .B(ori_ori_n35_), .C(e), .Y(ori_ori_n356_));
  NO2        o0328(.A(ori_ori_n356_), .B(ori_ori_n348_), .Y(ori_ori_n357_));
  NA3        o0329(.A(ori_ori_n336_), .B(ori_ori_n160_), .C(ori_ori_n77_), .Y(ori_ori_n358_));
  NAi31      o0330(.An(b), .B(c), .C(a), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n359_), .B(n), .Y(ori_ori_n360_));
  NO3        o0332(.A(ori_ori_n357_), .B(ori_ori_n355_), .C(ori_ori_n346_), .Y(ori_ori_n361_));
  NA2        o0333(.A(i), .B(o), .Y(ori_ori_n362_));
  NOi21      o0334(.An(a), .B(n), .Y(ori_ori_n363_));
  NOi21      o0335(.An(d), .B(c), .Y(ori_ori_n364_));
  NA2        o0336(.A(ori_ori_n364_), .B(ori_ori_n363_), .Y(ori_ori_n365_));
  NA3        o0337(.A(i), .B(o), .C(f), .Y(ori_ori_n366_));
  OR2        o0338(.A(ori_ori_n366_), .B(ori_ori_n64_), .Y(ori_ori_n367_));
  NA3        o0339(.A(ori_ori_n353_), .B(ori_ori_n352_), .C(ori_ori_n160_), .Y(ori_ori_n368_));
  AOI210     o0340(.A0(ori_ori_n368_), .A1(ori_ori_n367_), .B0(ori_ori_n365_), .Y(ori_ori_n369_));
  INV        o0341(.A(ori_ori_n369_), .Y(ori_ori_n370_));
  OR2        o0342(.A(n), .B(m), .Y(ori_ori_n371_));
  NO2        o0343(.A(ori_ori_n371_), .B(ori_ori_n136_), .Y(ori_ori_n372_));
  NO2        o0344(.A(ori_ori_n161_), .B(ori_ori_n131_), .Y(ori_ori_n373_));
  OAI210     o0345(.A0(ori_ori_n372_), .A1(ori_ori_n154_), .B0(ori_ori_n373_), .Y(ori_ori_n374_));
  INV        o0346(.A(ori_ori_n316_), .Y(ori_ori_n375_));
  NA3        o0347(.A(ori_ori_n375_), .B(ori_ori_n309_), .C(d), .Y(ori_ori_n376_));
  NO2        o0348(.A(ori_ori_n359_), .B(ori_ori_n48_), .Y(ori_ori_n377_));
  NO3        o0349(.A(ori_ori_n61_), .B(ori_ori_n101_), .C(e), .Y(ori_ori_n378_));
  NAi21      o0350(.An(k), .B(j), .Y(ori_ori_n379_));
  NA2        o0351(.A(ori_ori_n226_), .B(ori_ori_n379_), .Y(ori_ori_n380_));
  NA3        o0352(.A(ori_ori_n380_), .B(ori_ori_n378_), .C(ori_ori_n377_), .Y(ori_ori_n381_));
  NAi21      o0353(.An(e), .B(d), .Y(ori_ori_n382_));
  INV        o0354(.A(ori_ori_n382_), .Y(ori_ori_n383_));
  NO2        o0355(.A(ori_ori_n227_), .B(ori_ori_n190_), .Y(ori_ori_n384_));
  NA3        o0356(.A(ori_ori_n384_), .B(ori_ori_n383_), .C(ori_ori_n202_), .Y(ori_ori_n385_));
  NA4        o0357(.A(ori_ori_n385_), .B(ori_ori_n381_), .C(ori_ori_n376_), .D(ori_ori_n374_), .Y(ori_ori_n386_));
  NO2        o0358(.A(ori_ori_n286_), .B(ori_ori_n190_), .Y(ori_ori_n387_));
  NA2        o0359(.A(ori_ori_n387_), .B(ori_ori_n383_), .Y(ori_ori_n388_));
  NOi31      o0360(.An(n), .B(m), .C(k), .Y(ori_ori_n389_));
  AOI220     o0361(.A0(ori_ori_n389_), .A1(ori_ori_n328_), .B0(ori_ori_n198_), .B1(ori_ori_n49_), .Y(ori_ori_n390_));
  NAi31      o0362(.An(o), .B(f), .C(c), .Y(ori_ori_n391_));
  OR3        o0363(.A(ori_ori_n391_), .B(ori_ori_n390_), .C(e), .Y(ori_ori_n392_));
  NA3        o0364(.A(ori_ori_n392_), .B(ori_ori_n388_), .C(ori_ori_n265_), .Y(ori_ori_n393_));
  NOi41      o0365(.An(ori_ori_n370_), .B(ori_ori_n393_), .C(ori_ori_n386_), .D(ori_ori_n238_), .Y(ori_ori_n394_));
  NOi32      o0366(.An(c), .Bn(a), .C(b), .Y(ori_ori_n395_));
  NA2        o0367(.A(ori_ori_n395_), .B(ori_ori_n102_), .Y(ori_ori_n396_));
  INV        o0368(.A(ori_ori_n244_), .Y(ori_ori_n397_));
  AN2        o0369(.A(e), .B(d), .Y(ori_ori_n398_));
  INV        o0370(.A(ori_ori_n131_), .Y(ori_ori_n399_));
  NO2        o0371(.A(ori_ori_n117_), .B(ori_ori_n40_), .Y(ori_ori_n400_));
  NO2        o0372(.A(ori_ori_n61_), .B(e), .Y(ori_ori_n401_));
  NOi31      o0373(.An(j), .B(k), .C(i), .Y(ori_ori_n402_));
  NOi21      o0374(.An(ori_ori_n148_), .B(ori_ori_n402_), .Y(ori_ori_n403_));
  NA3        o0375(.A(ori_ori_n403_), .B(ori_ori_n235_), .C(ori_ori_n107_), .Y(ori_ori_n404_));
  AOI220     o0376(.A0(ori_ori_n404_), .A1(ori_ori_n401_), .B0(ori_ori_n400_), .B1(ori_ori_n399_), .Y(ori_ori_n405_));
  NO2        o0377(.A(ori_ori_n405_), .B(ori_ori_n396_), .Y(ori_ori_n406_));
  NO2        o0378(.A(ori_ori_n186_), .B(ori_ori_n181_), .Y(ori_ori_n407_));
  NOi21      o0379(.An(a), .B(b), .Y(ori_ori_n408_));
  NA3        o0380(.A(e), .B(d), .C(c), .Y(ori_ori_n409_));
  NAi21      o0381(.An(ori_ori_n409_), .B(ori_ori_n408_), .Y(ori_ori_n410_));
  NO2        o0382(.A(ori_ori_n358_), .B(ori_ori_n180_), .Y(ori_ori_n411_));
  NOi21      o0383(.An(ori_ori_n410_), .B(ori_ori_n411_), .Y(ori_ori_n412_));
  AOI210     o0384(.A0(ori_ori_n240_), .A1(ori_ori_n407_), .B0(ori_ori_n412_), .Y(ori_ori_n413_));
  NO4        o0385(.A(ori_ori_n165_), .B(ori_ori_n96_), .C(ori_ori_n55_), .D(b), .Y(ori_ori_n414_));
  NA2        o0386(.A(ori_ori_n323_), .B(ori_ori_n137_), .Y(ori_ori_n415_));
  OR2        o0387(.A(k), .B(j), .Y(ori_ori_n416_));
  NA2        o0388(.A(l), .B(k), .Y(ori_ori_n417_));
  NA3        o0389(.A(ori_ori_n417_), .B(ori_ori_n416_), .C(ori_ori_n198_), .Y(ori_ori_n418_));
  AOI210     o0390(.A0(ori_ori_n208_), .A1(ori_ori_n289_), .B0(ori_ori_n77_), .Y(ori_ori_n419_));
  NOi21      o0391(.An(ori_ori_n418_), .B(ori_ori_n419_), .Y(ori_ori_n420_));
  OR3        o0392(.A(ori_ori_n420_), .B(ori_ori_n127_), .C(ori_ori_n119_), .Y(ori_ori_n421_));
  INV        o0393(.A(ori_ori_n113_), .Y(ori_ori_n422_));
  NO3        o0394(.A(ori_ori_n358_), .B(ori_ori_n85_), .C(ori_ori_n117_), .Y(ori_ori_n423_));
  NO2        o0395(.A(ori_ori_n423_), .B(ori_ori_n422_), .Y(ori_ori_n424_));
  NA3        o0396(.A(ori_ori_n424_), .B(ori_ori_n421_), .C(ori_ori_n415_), .Y(ori_ori_n425_));
  NO4        o0397(.A(ori_ori_n425_), .B(ori_ori_n414_), .C(ori_ori_n413_), .D(ori_ori_n406_), .Y(ori_ori_n426_));
  INV        o0398(.A(e), .Y(ori_ori_n427_));
  NO2        o0399(.A(ori_ori_n165_), .B(ori_ori_n55_), .Y(ori_ori_n428_));
  NAi31      o0400(.An(j), .B(l), .C(i), .Y(ori_ori_n429_));
  OAI210     o0401(.A0(ori_ori_n429_), .A1(ori_ori_n118_), .B0(ori_ori_n96_), .Y(ori_ori_n430_));
  NA3        o0402(.A(ori_ori_n430_), .B(ori_ori_n428_), .C(ori_ori_n427_), .Y(ori_ori_n431_));
  NO2        o0403(.A(ori_ori_n337_), .B(ori_ori_n316_), .Y(ori_ori_n432_));
  NO2        o0404(.A(ori_ori_n432_), .B(ori_ori_n163_), .Y(ori_ori_n433_));
  NA3        o0405(.A(ori_ori_n433_), .B(ori_ori_n431_), .C(ori_ori_n216_), .Y(ori_ori_n434_));
  OAI210     o0406(.A0(ori_ori_n114_), .A1(ori_ori_n112_), .B0(n), .Y(ori_ori_n435_));
  XO2        o0407(.A(i), .B(h), .Y(ori_ori_n436_));
  NA3        o0408(.A(ori_ori_n436_), .B(ori_ori_n144_), .C(n), .Y(ori_ori_n437_));
  NA3        o0409(.A(ori_ori_n437_), .B(ori_ori_n390_), .C(ori_ori_n325_), .Y(ori_ori_n438_));
  NAi31      o0410(.An(c), .B(f), .C(d), .Y(ori_ori_n439_));
  AOI210     o0411(.A0(ori_ori_n245_), .A1(ori_ori_n171_), .B0(ori_ori_n439_), .Y(ori_ori_n440_));
  NOi21      o0412(.An(ori_ori_n75_), .B(ori_ori_n440_), .Y(ori_ori_n441_));
  NA2        o0413(.A(ori_ori_n203_), .B(ori_ori_n98_), .Y(ori_ori_n442_));
  AOI210     o0414(.A0(ori_ori_n442_), .A1(ori_ori_n159_), .B0(ori_ori_n439_), .Y(ori_ori_n443_));
  AOI210     o0415(.A0(ori_ori_n307_), .A1(ori_ori_n34_), .B0(ori_ori_n410_), .Y(ori_ori_n444_));
  NO2        o0416(.A(ori_ori_n444_), .B(ori_ori_n443_), .Y(ori_ori_n445_));
  AN2        o0417(.A(ori_ori_n252_), .B(ori_ori_n237_), .Y(ori_ori_n446_));
  NA3        o0418(.A(ori_ori_n36_), .B(ori_ori_n35_), .C(f), .Y(ori_ori_n447_));
  NAi31      o0419(.An(ori_ori_n446_), .B(ori_ori_n445_), .C(ori_ori_n441_), .Y(ori_ori_n448_));
  NO2        o0420(.A(ori_ori_n448_), .B(ori_ori_n434_), .Y(ori_ori_n449_));
  NA4        o0421(.A(ori_ori_n449_), .B(ori_ori_n426_), .C(ori_ori_n394_), .D(ori_ori_n361_), .Y(ori11));
  NO2        o0422(.A(ori_ori_n66_), .B(f), .Y(ori_ori_n451_));
  NA2        o0423(.A(j), .B(o), .Y(ori_ori_n452_));
  NAi31      o0424(.An(i), .B(m), .C(l), .Y(ori_ori_n453_));
  NA3        o0425(.A(m), .B(k), .C(j), .Y(ori_ori_n454_));
  OAI220     o0426(.A0(ori_ori_n454_), .A1(ori_ori_n117_), .B0(ori_ori_n453_), .B1(ori_ori_n452_), .Y(ori_ori_n455_));
  NA2        o0427(.A(ori_ori_n455_), .B(ori_ori_n451_), .Y(ori_ori_n456_));
  NOi32      o0428(.An(e), .Bn(b), .C(f), .Y(ori_ori_n457_));
  NA2        o0429(.A(ori_ori_n45_), .B(j), .Y(ori_ori_n458_));
  NAi31      o0430(.An(d), .B(e), .C(a), .Y(ori_ori_n459_));
  NO2        o0431(.A(ori_ori_n459_), .B(n), .Y(ori_ori_n460_));
  NA2        o0432(.A(ori_ori_n460_), .B(ori_ori_n95_), .Y(ori_ori_n461_));
  NA2        o0433(.A(j), .B(i), .Y(ori_ori_n462_));
  NAi31      o0434(.An(n), .B(m), .C(k), .Y(ori_ori_n463_));
  NO3        o0435(.A(ori_ori_n463_), .B(ori_ori_n462_), .C(ori_ori_n101_), .Y(ori_ori_n464_));
  NO4        o0436(.A(n), .B(d), .C(ori_ori_n104_), .D(a), .Y(ori_ori_n465_));
  OR2        o0437(.A(n), .B(c), .Y(ori_ori_n466_));
  NO2        o0438(.A(ori_ori_n466_), .B(ori_ori_n133_), .Y(ori_ori_n467_));
  NO2        o0439(.A(ori_ori_n467_), .B(ori_ori_n465_), .Y(ori_ori_n468_));
  NOi32      o0440(.An(o), .Bn(f), .C(i), .Y(ori_ori_n469_));
  AOI220     o0441(.A0(ori_ori_n469_), .A1(ori_ori_n93_), .B0(ori_ori_n455_), .B1(f), .Y(ori_ori_n470_));
  NO2        o0442(.A(ori_ori_n470_), .B(ori_ori_n468_), .Y(ori_ori_n471_));
  INV        o0443(.A(ori_ori_n471_), .Y(ori_ori_n472_));
  NA2        o0444(.A(ori_ori_n123_), .B(ori_ori_n33_), .Y(ori_ori_n473_));
  OAI220     o0445(.A0(ori_ori_n473_), .A1(m), .B0(ori_ori_n458_), .B1(ori_ori_n208_), .Y(ori_ori_n474_));
  NOi41      o0446(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n475_));
  NAi32      o0447(.An(e), .Bn(b), .C(c), .Y(ori_ori_n476_));
  OR2        o0448(.A(ori_ori_n476_), .B(ori_ori_n77_), .Y(ori_ori_n477_));
  AN2        o0449(.A(ori_ori_n290_), .B(ori_ori_n273_), .Y(ori_ori_n478_));
  NA2        o0450(.A(ori_ori_n478_), .B(ori_ori_n477_), .Y(ori_ori_n479_));
  OA210      o0451(.A0(ori_ori_n479_), .A1(ori_ori_n475_), .B0(ori_ori_n474_), .Y(ori_ori_n480_));
  OAI220     o0452(.A0(ori_ori_n339_), .A1(ori_ori_n338_), .B0(ori_ori_n453_), .B1(ori_ori_n452_), .Y(ori_ori_n481_));
  NO2        o0453(.A(ori_ori_n206_), .B(ori_ori_n99_), .Y(ori_ori_n482_));
  NA2        o0454(.A(ori_ori_n340_), .B(ori_ori_n482_), .Y(ori_ori_n483_));
  INV        o0455(.A(ori_ori_n483_), .Y(ori_ori_n484_));
  INV        o0456(.A(ori_ori_n360_), .Y(ori_ori_n485_));
  NA2        o0457(.A(ori_ori_n481_), .B(f), .Y(ori_ori_n486_));
  NAi32      o0458(.An(d), .Bn(a), .C(b), .Y(ori_ori_n487_));
  NO2        o0459(.A(ori_ori_n487_), .B(ori_ori_n48_), .Y(ori_ori_n488_));
  NA2        o0460(.A(h), .B(f), .Y(ori_ori_n489_));
  NO2        o0461(.A(ori_ori_n489_), .B(ori_ori_n88_), .Y(ori_ori_n490_));
  NO3        o0462(.A(ori_ori_n155_), .B(ori_ori_n152_), .C(o), .Y(ori_ori_n491_));
  AOI220     o0463(.A0(ori_ori_n491_), .A1(ori_ori_n57_), .B0(ori_ori_n490_), .B1(ori_ori_n488_), .Y(ori_ori_n492_));
  OAI210     o0464(.A0(ori_ori_n486_), .A1(ori_ori_n485_), .B0(ori_ori_n492_), .Y(ori_ori_n493_));
  AN3        o0465(.A(j), .B(h), .C(o), .Y(ori_ori_n494_));
  NA3        o0466(.A(f), .B(d), .C(b), .Y(ori_ori_n495_));
  NO4        o0467(.A(ori_ori_n495_), .B(ori_ori_n155_), .C(ori_ori_n152_), .D(o), .Y(ori_ori_n496_));
  NO4        o0468(.A(ori_ori_n496_), .B(ori_ori_n493_), .C(ori_ori_n484_), .D(ori_ori_n480_), .Y(ori_ori_n497_));
  AN4        o0469(.A(ori_ori_n497_), .B(ori_ori_n472_), .C(ori_ori_n461_), .D(ori_ori_n456_), .Y(ori_ori_n498_));
  INV        o0470(.A(k), .Y(ori_ori_n499_));
  NA3        o0471(.A(l), .B(ori_ori_n499_), .C(i), .Y(ori_ori_n500_));
  INV        o0472(.A(ori_ori_n500_), .Y(ori_ori_n501_));
  NAi32      o0473(.An(h), .Bn(f), .C(o), .Y(ori_ori_n502_));
  NAi41      o0474(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n503_));
  OAI210     o0475(.A0(ori_ori_n459_), .A1(n), .B0(ori_ori_n503_), .Y(ori_ori_n504_));
  NA2        o0476(.A(ori_ori_n504_), .B(m), .Y(ori_ori_n505_));
  NAi31      o0477(.An(h), .B(o), .C(f), .Y(ori_ori_n506_));
  NO3        o0478(.A(ori_ori_n502_), .B(ori_ori_n66_), .C(ori_ori_n67_), .Y(ori_ori_n507_));
  NO4        o0479(.A(ori_ori_n506_), .B(ori_ori_n466_), .C(ori_ori_n133_), .D(ori_ori_n67_), .Y(ori_ori_n508_));
  OR2        o0480(.A(ori_ori_n508_), .B(ori_ori_n507_), .Y(ori_ori_n509_));
  NAi31      o0481(.An(f), .B(h), .C(o), .Y(ori_ori_n510_));
  NOi32      o0482(.An(d), .Bn(a), .C(e), .Y(ori_ori_n511_));
  NO2        o0483(.A(n), .B(c), .Y(ori_ori_n512_));
  NA3        o0484(.A(ori_ori_n512_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n513_));
  INV        o0485(.A(ori_ori_n513_), .Y(ori_ori_n514_));
  NOi32      o0486(.An(e), .Bn(a), .C(d), .Y(ori_ori_n515_));
  AOI210     o0487(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n515_), .Y(ori_ori_n516_));
  INV        o0488(.A(ori_ori_n473_), .Y(ori_ori_n517_));
  NA2        o0489(.A(ori_ori_n517_), .B(ori_ori_n514_), .Y(ori_ori_n518_));
  OAI210     o0490(.A0(ori_ori_n222_), .A1(ori_ori_n80_), .B0(ori_ori_n518_), .Y(ori_ori_n519_));
  AOI210     o0491(.A0(ori_ori_n509_), .A1(ori_ori_n501_), .B0(ori_ori_n519_), .Y(ori_ori_n520_));
  NO3        o0492(.A(ori_ori_n271_), .B(ori_ori_n59_), .C(n), .Y(ori_ori_n521_));
  NA3        o0493(.A(ori_ori_n439_), .B(ori_ori_n150_), .C(ori_ori_n149_), .Y(ori_ori_n522_));
  NA2        o0494(.A(ori_ori_n391_), .B(ori_ori_n206_), .Y(ori_ori_n523_));
  OR2        o0495(.A(ori_ori_n523_), .B(ori_ori_n522_), .Y(ori_ori_n524_));
  NA2        o0496(.A(ori_ori_n524_), .B(ori_ori_n521_), .Y(ori_ori_n525_));
  NO2        o0497(.A(ori_ori_n525_), .B(ori_ori_n80_), .Y(ori_ori_n526_));
  NA3        o0498(.A(ori_ori_n475_), .B(ori_ori_n291_), .C(ori_ori_n45_), .Y(ori_ori_n527_));
  NOi32      o0499(.An(e), .Bn(c), .C(f), .Y(ori_ori_n528_));
  NOi21      o0500(.An(f), .B(o), .Y(ori_ori_n529_));
  NO2        o0501(.A(ori_ori_n529_), .B(ori_ori_n188_), .Y(ori_ori_n530_));
  AOI220     o0502(.A0(ori_ori_n530_), .A1(ori_ori_n333_), .B0(ori_ori_n528_), .B1(ori_ori_n154_), .Y(ori_ori_n531_));
  NA3        o0503(.A(ori_ori_n531_), .B(ori_ori_n527_), .C(ori_ori_n157_), .Y(ori_ori_n532_));
  NOi21      o0504(.An(j), .B(l), .Y(ori_ori_n533_));
  NAi21      o0505(.An(k), .B(h), .Y(ori_ori_n534_));
  NO2        o0506(.A(ori_ori_n534_), .B(ori_ori_n236_), .Y(ori_ori_n535_));
  NA2        o0507(.A(ori_ori_n535_), .B(ori_ori_n533_), .Y(ori_ori_n536_));
  OR2        o0508(.A(ori_ori_n536_), .B(ori_ori_n505_), .Y(ori_ori_n537_));
  NO2        o0509(.A(ori_ori_n266_), .B(ori_ori_n510_), .Y(ori_ori_n538_));
  NO2        o0510(.A(ori_ori_n459_), .B(ori_ori_n48_), .Y(ori_ori_n539_));
  NA2        o0511(.A(ori_ori_n539_), .B(ori_ori_n538_), .Y(ori_ori_n540_));
  NA2        o0512(.A(ori_ori_n540_), .B(ori_ori_n537_), .Y(ori_ori_n541_));
  NA2        o0513(.A(ori_ori_n98_), .B(ori_ori_n35_), .Y(ori_ori_n542_));
  INV        o0514(.A(ori_ori_n309_), .Y(ori_ori_n543_));
  NO2        o0515(.A(ori_ori_n543_), .B(n), .Y(ori_ori_n544_));
  NO2        o0516(.A(ori_ori_n458_), .B(ori_ori_n155_), .Y(ori_ori_n545_));
  NA3        o0517(.A(ori_ori_n476_), .B(ori_ori_n242_), .C(ori_ori_n128_), .Y(ori_ori_n546_));
  NA2        o0518(.A(ori_ori_n436_), .B(ori_ori_n144_), .Y(ori_ori_n547_));
  NO3        o0519(.A(ori_ori_n334_), .B(ori_ori_n547_), .C(ori_ori_n80_), .Y(ori_ori_n548_));
  AOI210     o0520(.A0(ori_ori_n546_), .A1(ori_ori_n545_), .B0(ori_ori_n548_), .Y(ori_ori_n549_));
  AN3        o0521(.A(f), .B(d), .C(b), .Y(ori_ori_n550_));
  NAi31      o0522(.An(m), .B(n), .C(k), .Y(ori_ori_n551_));
  OR2        o0523(.A(ori_ori_n119_), .B(ori_ori_n59_), .Y(ori_ori_n552_));
  OAI210     o0524(.A0(ori_ori_n552_), .A1(ori_ori_n551_), .B0(ori_ori_n224_), .Y(ori_ori_n553_));
  NA2        o0525(.A(ori_ori_n553_), .B(j), .Y(ori_ori_n554_));
  NA2        o0526(.A(ori_ori_n554_), .B(ori_ori_n549_), .Y(ori_ori_n555_));
  NO4        o0527(.A(ori_ori_n555_), .B(ori_ori_n541_), .C(ori_ori_n532_), .D(ori_ori_n526_), .Y(ori_ori_n556_));
  NAi31      o0528(.An(o), .B(h), .C(f), .Y(ori_ori_n557_));
  OA210      o0529(.A0(ori_ori_n459_), .A1(n), .B0(ori_ori_n503_), .Y(ori_ori_n558_));
  NO3        o0530(.A(o), .B(ori_ori_n190_), .C(ori_ori_n55_), .Y(ori_ori_n559_));
  NA2        o0531(.A(ori_ori_n333_), .B(ori_ori_n559_), .Y(ori_ori_n560_));
  OR2        o0532(.A(ori_ori_n66_), .B(ori_ori_n67_), .Y(ori_ori_n561_));
  OR2        o0533(.A(ori_ori_n536_), .B(ori_ori_n561_), .Y(ori_ori_n562_));
  AN2        o0534(.A(h), .B(f), .Y(ori_ori_n563_));
  NA2        o0535(.A(ori_ori_n563_), .B(ori_ori_n36_), .Y(ori_ori_n564_));
  NO2        o0536(.A(ori_ori_n564_), .B(ori_ori_n396_), .Y(ori_ori_n565_));
  AOI210     o0537(.A0(ori_ori_n487_), .A1(ori_ori_n359_), .B0(ori_ori_n48_), .Y(ori_ori_n566_));
  OAI220     o0538(.A0(ori_ori_n506_), .A1(ori_ori_n500_), .B0(ori_ori_n279_), .B1(ori_ori_n452_), .Y(ori_ori_n567_));
  AOI210     o0539(.A0(ori_ori_n567_), .A1(ori_ori_n566_), .B0(ori_ori_n565_), .Y(ori_ori_n568_));
  NA3        o0540(.A(ori_ori_n568_), .B(ori_ori_n562_), .C(ori_ori_n560_), .Y(ori_ori_n569_));
  NA2        o0541(.A(ori_ori_n118_), .B(ori_ori_n48_), .Y(ori_ori_n570_));
  AOI220     o0542(.A0(ori_ori_n570_), .A1(ori_ori_n457_), .B0(ori_ori_n309_), .B1(ori_ori_n102_), .Y(ori_ori_n571_));
  OR2        o0543(.A(ori_ori_n571_), .B(ori_ori_n473_), .Y(ori_ori_n572_));
  INV        o0544(.A(ori_ori_n572_), .Y(ori_ori_n573_));
  NO3        o0545(.A(ori_ori_n344_), .B(ori_ori_n168_), .C(ori_ori_n167_), .Y(ori_ori_n574_));
  NA2        o0546(.A(ori_ori_n574_), .B(ori_ori_n206_), .Y(ori_ori_n575_));
  NA3        o0547(.A(ori_ori_n575_), .B(ori_ori_n228_), .C(j), .Y(ori_ori_n576_));
  NO3        o0548(.A(ori_ori_n391_), .B(ori_ori_n152_), .C(i), .Y(ori_ori_n577_));
  NA2        o0549(.A(ori_ori_n395_), .B(ori_ori_n77_), .Y(ori_ori_n578_));
  NO4        o0550(.A(ori_ori_n454_), .B(ori_ori_n578_), .C(ori_ori_n117_), .D(ori_ori_n190_), .Y(ori_ori_n579_));
  INV        o0551(.A(ori_ori_n579_), .Y(ori_ori_n580_));
  NA3        o0552(.A(ori_ori_n580_), .B(ori_ori_n576_), .C(ori_ori_n342_), .Y(ori_ori_n581_));
  NO3        o0553(.A(ori_ori_n581_), .B(ori_ori_n573_), .C(ori_ori_n569_), .Y(ori_ori_n582_));
  NA4        o0554(.A(ori_ori_n582_), .B(ori_ori_n556_), .C(ori_ori_n520_), .D(ori_ori_n498_), .Y(ori08));
  NO2        o0555(.A(k), .B(h), .Y(ori_ori_n584_));
  AO210      o0556(.A0(ori_ori_n226_), .A1(ori_ori_n379_), .B0(ori_ori_n584_), .Y(ori_ori_n585_));
  NO2        o0557(.A(ori_ori_n585_), .B(ori_ori_n259_), .Y(ori_ori_n586_));
  NA2        o0558(.A(ori_ori_n528_), .B(ori_ori_n77_), .Y(ori_ori_n587_));
  NA2        o0559(.A(ori_ori_n587_), .B(ori_ori_n391_), .Y(ori_ori_n588_));
  AOI210     o0560(.A0(ori_ori_n588_), .A1(ori_ori_n586_), .B0(ori_ori_n423_), .Y(ori_ori_n589_));
  NA2        o0561(.A(ori_ori_n77_), .B(ori_ori_n99_), .Y(ori_ori_n590_));
  NO2        o0562(.A(ori_ori_n590_), .B(ori_ori_n56_), .Y(ori_ori_n591_));
  NO4        o0563(.A(ori_ori_n320_), .B(ori_ori_n101_), .C(j), .D(ori_ori_n191_), .Y(ori_ori_n592_));
  NA2        o0564(.A(ori_ori_n592_), .B(ori_ori_n591_), .Y(ori_ori_n593_));
  AOI210     o0565(.A0(ori_ori_n495_), .A1(ori_ori_n140_), .B0(ori_ori_n77_), .Y(ori_ori_n594_));
  NA4        o0566(.A(ori_ori_n193_), .B(ori_ori_n123_), .C(ori_ori_n44_), .D(h), .Y(ori_ori_n595_));
  AN2        o0567(.A(l), .B(k), .Y(ori_ori_n596_));
  NA4        o0568(.A(ori_ori_n596_), .B(ori_ori_n98_), .C(ori_ori_n67_), .D(ori_ori_n191_), .Y(ori_ori_n597_));
  OAI210     o0569(.A0(ori_ori_n595_), .A1(o), .B0(ori_ori_n597_), .Y(ori_ori_n598_));
  NA2        o0570(.A(ori_ori_n598_), .B(ori_ori_n594_), .Y(ori_ori_n599_));
  NA4        o0571(.A(ori_ori_n599_), .B(ori_ori_n593_), .C(ori_ori_n589_), .D(ori_ori_n298_), .Y(ori_ori_n600_));
  AN2        o0572(.A(ori_ori_n460_), .B(ori_ori_n89_), .Y(ori_ori_n601_));
  NO4        o0573(.A(ori_ori_n152_), .B(ori_ori_n332_), .C(ori_ori_n101_), .D(o), .Y(ori_ori_n602_));
  NO2        o0574(.A(ori_ori_n37_), .B(ori_ori_n190_), .Y(ori_ori_n603_));
  NA2        o0575(.A(ori_ori_n530_), .B(ori_ori_n295_), .Y(ori_ori_n604_));
  NAi21      o0576(.An(ori_ori_n601_), .B(ori_ori_n604_), .Y(ori_ori_n605_));
  OAI210     o0577(.A0(ori_ori_n476_), .A1(ori_ori_n46_), .B0(ori_ori_n552_), .Y(ori_ori_n606_));
  NO2        o0578(.A(ori_ori_n417_), .B(ori_ori_n118_), .Y(ori_ori_n607_));
  NA2        o0579(.A(ori_ori_n607_), .B(ori_ori_n606_), .Y(ori_ori_n608_));
  NO3        o0580(.A(ori_ori_n271_), .B(ori_ori_n117_), .C(ori_ori_n40_), .Y(ori_ori_n609_));
  NAi21      o0581(.An(ori_ori_n609_), .B(ori_ori_n597_), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n585_), .B(ori_ori_n120_), .Y(ori_ori_n611_));
  AOI220     o0583(.A0(ori_ori_n611_), .A1(ori_ori_n343_), .B0(ori_ori_n610_), .B1(ori_ori_n70_), .Y(ori_ori_n612_));
  NA2        o0584(.A(ori_ori_n608_), .B(ori_ori_n612_), .Y(ori_ori_n613_));
  NA3        o0585(.A(ori_ori_n575_), .B(ori_ori_n285_), .C(ori_ori_n324_), .Y(ori_ori_n614_));
  NA3        o0586(.A(m), .B(l), .C(k), .Y(ori_ori_n615_));
  INV        o0587(.A(ori_ori_n614_), .Y(ori_ori_n616_));
  NO4        o0588(.A(ori_ori_n616_), .B(ori_ori_n613_), .C(ori_ori_n605_), .D(ori_ori_n600_), .Y(ori_ori_n617_));
  NO3        o0589(.A(ori_ori_n337_), .B(ori_ori_n452_), .C(h), .Y(ori_ori_n618_));
  NA2        o0590(.A(ori_ori_n618_), .B(ori_ori_n102_), .Y(ori_ori_n619_));
  NA2        o0591(.A(ori_ori_n619_), .B(ori_ori_n225_), .Y(ori_ori_n620_));
  NA2        o0592(.A(ori_ori_n596_), .B(ori_ori_n67_), .Y(ori_ori_n621_));
  NO4        o0593(.A(ori_ori_n574_), .B(ori_ori_n152_), .C(n), .D(i), .Y(ori_ori_n622_));
  NOi21      o0594(.An(h), .B(j), .Y(ori_ori_n623_));
  NA2        o0595(.A(ori_ori_n623_), .B(f), .Y(ori_ori_n624_));
  NO2        o0596(.A(ori_ori_n622_), .B(ori_ori_n577_), .Y(ori_ori_n625_));
  NO2        o0597(.A(ori_ori_n625_), .B(ori_ori_n621_), .Y(ori_ori_n626_));
  AOI210     o0598(.A0(ori_ori_n620_), .A1(l), .B0(ori_ori_n626_), .Y(ori_ori_n627_));
  NO2        o0599(.A(j), .B(i), .Y(ori_ori_n628_));
  NA3        o0600(.A(ori_ori_n628_), .B(ori_ori_n74_), .C(l), .Y(ori_ori_n629_));
  NA2        o0601(.A(ori_ori_n628_), .B(ori_ori_n32_), .Y(ori_ori_n630_));
  OR2        o0602(.A(ori_ori_n629_), .B(ori_ori_n505_), .Y(ori_ori_n631_));
  NO3        o0603(.A(ori_ori_n135_), .B(ori_ori_n48_), .C(ori_ori_n99_), .Y(ori_ori_n632_));
  NO3        o0604(.A(ori_ori_n466_), .B(ori_ori_n133_), .C(ori_ori_n67_), .Y(ori_ori_n633_));
  NO3        o0605(.A(ori_ori_n417_), .B(ori_ori_n366_), .C(j), .Y(ori_ori_n634_));
  OAI210     o0606(.A0(ori_ori_n633_), .A1(ori_ori_n632_), .B0(ori_ori_n634_), .Y(ori_ori_n635_));
  INV        o0607(.A(ori_ori_n635_), .Y(ori_ori_n636_));
  INV        o0608(.A(j), .Y(ori_ori_n637_));
  NO3        o0609(.A(ori_ori_n259_), .B(ori_ori_n637_), .C(ori_ori_n39_), .Y(ori_ori_n638_));
  AOI210     o0610(.A0(ori_ori_n457_), .A1(n), .B0(ori_ori_n475_), .Y(ori_ori_n639_));
  NA2        o0611(.A(ori_ori_n639_), .B(ori_ori_n478_), .Y(ori_ori_n640_));
  AN3        o0612(.A(ori_ori_n640_), .B(ori_ori_n638_), .C(ori_ori_n92_), .Y(ori_ori_n641_));
  NO3        o0613(.A(ori_ori_n152_), .B(ori_ori_n332_), .C(ori_ori_n101_), .Y(ori_ori_n642_));
  AOI220     o0614(.A0(ori_ori_n642_), .A1(ori_ori_n220_), .B0(ori_ori_n523_), .B1(ori_ori_n264_), .Y(ori_ori_n643_));
  NAi31      o0615(.An(ori_ori_n516_), .B(ori_ori_n86_), .C(ori_ori_n77_), .Y(ori_ori_n644_));
  NA2        o0616(.A(ori_ori_n644_), .B(ori_ori_n643_), .Y(ori_ori_n645_));
  NA2        o0617(.A(ori_ori_n609_), .B(ori_ori_n594_), .Y(ori_ori_n646_));
  NO2        o0618(.A(ori_ori_n615_), .B(ori_ori_n84_), .Y(ori_ori_n647_));
  NA2        o0619(.A(ori_ori_n647_), .B(ori_ori_n504_), .Y(ori_ori_n648_));
  NO2        o0620(.A(ori_ori_n506_), .B(ori_ori_n105_), .Y(ori_ori_n649_));
  OAI210     o0621(.A0(ori_ori_n649_), .A1(ori_ori_n634_), .B0(ori_ori_n566_), .Y(ori_ori_n650_));
  NA3        o0622(.A(ori_ori_n650_), .B(ori_ori_n648_), .C(ori_ori_n646_), .Y(ori_ori_n651_));
  OR4        o0623(.A(ori_ori_n651_), .B(ori_ori_n645_), .C(ori_ori_n641_), .D(ori_ori_n636_), .Y(ori_ori_n652_));
  NA3        o0624(.A(ori_ori_n639_), .B(ori_ori_n478_), .C(ori_ori_n477_), .Y(ori_ori_n653_));
  NA4        o0625(.A(ori_ori_n653_), .B(ori_ori_n193_), .C(ori_ori_n379_), .D(ori_ori_n33_), .Y(ori_ori_n654_));
  NO4        o0626(.A(ori_ori_n417_), .B(ori_ori_n362_), .C(j), .D(f), .Y(ori_ori_n655_));
  NA3        o0627(.A(ori_ori_n469_), .B(ori_ori_n256_), .C(h), .Y(ori_ori_n656_));
  NOi21      o0628(.An(ori_ori_n566_), .B(ori_ori_n656_), .Y(ori_ori_n657_));
  OAI220     o0629(.A0(ori_ori_n656_), .A1(ori_ori_n513_), .B0(ori_ori_n629_), .B1(ori_ori_n561_), .Y(ori_ori_n658_));
  INV        o0630(.A(ori_ori_n658_), .Y(ori_ori_n659_));
  NAi31      o0631(.An(ori_ori_n657_), .B(ori_ori_n659_), .C(ori_ori_n654_), .Y(ori_ori_n660_));
  BUFFER     o0632(.A(ori_ori_n647_), .Y(ori_ori_n661_));
  NA2        o0633(.A(ori_ori_n661_), .B(ori_ori_n212_), .Y(ori_ori_n662_));
  NO2        o0634(.A(ori_ori_n558_), .B(ori_ori_n67_), .Y(ori_ori_n663_));
  AOI210     o0635(.A0(ori_ori_n655_), .A1(ori_ori_n663_), .B0(ori_ori_n287_), .Y(ori_ori_n664_));
  OAI210     o0636(.A0(ori_ori_n615_), .A1(ori_ori_n557_), .B0(ori_ori_n447_), .Y(ori_ori_n665_));
  NA3        o0637(.A(ori_ori_n223_), .B(ori_ori_n58_), .C(b), .Y(ori_ori_n666_));
  AOI220     o0638(.A0(ori_ori_n512_), .A1(ori_ori_n29_), .B0(ori_ori_n395_), .B1(ori_ori_n77_), .Y(ori_ori_n667_));
  NA2        o0639(.A(ori_ori_n667_), .B(ori_ori_n666_), .Y(ori_ori_n668_));
  NA2        o0640(.A(ori_ori_n668_), .B(ori_ori_n665_), .Y(ori_ori_n669_));
  NA3        o0641(.A(ori_ori_n669_), .B(ori_ori_n664_), .C(ori_ori_n662_), .Y(ori_ori_n670_));
  NOi41      o0642(.An(ori_ori_n631_), .B(ori_ori_n670_), .C(ori_ori_n660_), .D(ori_ori_n652_), .Y(ori_ori_n671_));
  NO3        o0643(.A(ori_ori_n292_), .B(ori_ori_n260_), .C(ori_ori_n101_), .Y(ori_ori_n672_));
  NA2        o0644(.A(ori_ori_n672_), .B(ori_ori_n640_), .Y(ori_ori_n673_));
  NA2        o0645(.A(ori_ori_n673_), .B(ori_ori_n345_), .Y(ori_ori_n674_));
  OR2        o0646(.A(ori_ori_n557_), .B(ori_ori_n85_), .Y(ori_ori_n675_));
  NOi31      o0647(.An(b), .B(d), .C(a), .Y(ori_ori_n676_));
  NO2        o0648(.A(ori_ori_n676_), .B(ori_ori_n511_), .Y(ori_ori_n677_));
  NO2        o0649(.A(ori_ori_n677_), .B(n), .Y(ori_ori_n678_));
  NOi21      o0650(.An(ori_ori_n667_), .B(ori_ori_n678_), .Y(ori_ori_n679_));
  NO2        o0651(.A(ori_ori_n679_), .B(ori_ori_n675_), .Y(ori_ori_n680_));
  NO2        o0652(.A(ori_ori_n476_), .B(ori_ori_n77_), .Y(ori_ori_n681_));
  NA2        o0653(.A(ori_ori_n672_), .B(ori_ori_n681_), .Y(ori_ori_n682_));
  OAI210     o0654(.A0(ori_ori_n595_), .A1(ori_ori_n334_), .B0(ori_ori_n682_), .Y(ori_ori_n683_));
  NO2        o0655(.A(ori_ori_n574_), .B(n), .Y(ori_ori_n684_));
  NA2        o0656(.A(ori_ori_n684_), .B(ori_ori_n586_), .Y(ori_ori_n685_));
  NO2        o0657(.A(ori_ori_n276_), .B(ori_ori_n211_), .Y(ori_ori_n686_));
  OAI210     o0658(.A0(ori_ori_n89_), .A1(ori_ori_n86_), .B0(ori_ori_n686_), .Y(ori_ori_n687_));
  INV        o0659(.A(ori_ori_n687_), .Y(ori_ori_n688_));
  NA2        o0660(.A(ori_ori_n602_), .B(ori_ori_n297_), .Y(ori_ori_n689_));
  OAI210     o0661(.A0(ori_ori_n508_), .A1(ori_ori_n507_), .B0(ori_ori_n310_), .Y(ori_ori_n690_));
  AN2        o0662(.A(ori_ori_n690_), .B(ori_ori_n689_), .Y(ori_ori_n691_));
  NAi31      o0663(.An(ori_ori_n688_), .B(ori_ori_n691_), .C(ori_ori_n685_), .Y(ori_ori_n692_));
  NO4        o0664(.A(ori_ori_n692_), .B(ori_ori_n683_), .C(ori_ori_n680_), .D(ori_ori_n674_), .Y(ori_ori_n693_));
  NA4        o0665(.A(ori_ori_n693_), .B(ori_ori_n671_), .C(ori_ori_n627_), .D(ori_ori_n617_), .Y(ori09));
  INV        o0666(.A(ori_ori_n110_), .Y(ori_ori_n695_));
  NA2        o0667(.A(f), .B(e), .Y(ori_ori_n696_));
  NO2        o0668(.A(ori_ori_n201_), .B(ori_ori_n101_), .Y(ori_ori_n697_));
  NA4        o0669(.A(ori_ori_n266_), .B(ori_ori_n403_), .C(ori_ori_n235_), .D(ori_ori_n107_), .Y(ori_ori_n698_));
  AOI210     o0670(.A0(ori_ori_n698_), .A1(o), .B0(ori_ori_n400_), .Y(ori_ori_n699_));
  NO2        o0671(.A(ori_ori_n699_), .B(ori_ori_n696_), .Y(ori_ori_n700_));
  NA2        o0672(.A(ori_ori_n372_), .B(e), .Y(ori_ori_n701_));
  NO2        o0673(.A(ori_ori_n701_), .B(ori_ori_n439_), .Y(ori_ori_n702_));
  AOI210     o0674(.A0(ori_ori_n700_), .A1(ori_ori_n695_), .B0(ori_ori_n702_), .Y(ori_ori_n703_));
  NA3        o0675(.A(m), .B(l), .C(i), .Y(ori_ori_n704_));
  OAI220     o0676(.A0(ori_ori_n506_), .A1(ori_ori_n704_), .B0(ori_ori_n300_), .B1(ori_ori_n453_), .Y(ori_ori_n705_));
  NA4        o0677(.A(ori_ori_n81_), .B(ori_ori_n80_), .C(o), .D(f), .Y(ori_ori_n706_));
  NAi31      o0678(.An(ori_ori_n705_), .B(ori_ori_n706_), .C(ori_ori_n367_), .Y(ori_ori_n707_));
  NA3        o0679(.A(ori_ori_n675_), .B(ori_ori_n486_), .C(ori_ori_n447_), .Y(ori_ori_n708_));
  OA210      o0680(.A0(ori_ori_n708_), .A1(ori_ori_n707_), .B0(ori_ori_n678_), .Y(ori_ori_n709_));
  INV        o0681(.A(ori_ori_n290_), .Y(ori_ori_n710_));
  NO2        o0682(.A(ori_ori_n114_), .B(ori_ori_n112_), .Y(ori_ori_n711_));
  NOi31      o0683(.An(k), .B(m), .C(l), .Y(ori_ori_n712_));
  NO2        o0684(.A(ori_ori_n291_), .B(ori_ori_n712_), .Y(ori_ori_n713_));
  AOI210     o0685(.A0(ori_ori_n713_), .A1(ori_ori_n711_), .B0(ori_ori_n510_), .Y(ori_ori_n714_));
  NA2        o0686(.A(ori_ori_n666_), .B(ori_ori_n284_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n293_), .B(ori_ori_n294_), .Y(ori_ori_n716_));
  OAI210     o0688(.A0(ori_ori_n180_), .A1(ori_ori_n190_), .B0(ori_ori_n716_), .Y(ori_ori_n717_));
  AOI220     o0689(.A0(ori_ori_n717_), .A1(ori_ori_n715_), .B0(ori_ori_n714_), .B1(ori_ori_n710_), .Y(ori_ori_n718_));
  NA3        o0690(.A(ori_ori_n718_), .B(ori_ori_n531_), .C(ori_ori_n75_), .Y(ori_ori_n719_));
  NO2        o0691(.A(ori_ori_n502_), .B(ori_ori_n429_), .Y(ori_ori_n720_));
  NA2        o0692(.A(ori_ori_n720_), .B(ori_ori_n166_), .Y(ori_ori_n721_));
  NOi21      o0693(.An(f), .B(d), .Y(ori_ori_n722_));
  NA2        o0694(.A(ori_ori_n722_), .B(m), .Y(ori_ori_n723_));
  NO2        o0695(.A(ori_ori_n723_), .B(ori_ori_n51_), .Y(ori_ori_n724_));
  NOi32      o0696(.An(o), .Bn(f), .C(d), .Y(ori_ori_n725_));
  NA4        o0697(.A(ori_ori_n725_), .B(ori_ori_n512_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n726_));
  NOi21      o0698(.An(ori_ori_n267_), .B(ori_ori_n726_), .Y(ori_ori_n727_));
  AOI210     o0699(.A0(ori_ori_n724_), .A1(ori_ori_n467_), .B0(ori_ori_n727_), .Y(ori_ori_n728_));
  NA2        o0700(.A(ori_ori_n235_), .B(ori_ori_n107_), .Y(ori_ori_n729_));
  AN2        o0701(.A(f), .B(d), .Y(ori_ori_n730_));
  NA3        o0702(.A(ori_ori_n408_), .B(ori_ori_n730_), .C(ori_ori_n77_), .Y(ori_ori_n731_));
  NO3        o0703(.A(ori_ori_n731_), .B(ori_ori_n67_), .C(ori_ori_n191_), .Y(ori_ori_n732_));
  NA2        o0704(.A(ori_ori_n729_), .B(ori_ori_n732_), .Y(ori_ori_n733_));
  NAi41      o0705(.An(ori_ori_n422_), .B(ori_ori_n733_), .C(ori_ori_n728_), .D(ori_ori_n721_), .Y(ori_ori_n734_));
  NO4        o0706(.A(ori_ori_n529_), .B(ori_ori_n118_), .C(ori_ori_n281_), .D(ori_ori_n136_), .Y(ori_ori_n735_));
  INV        o0707(.A(ori_ori_n735_), .Y(ori_ori_n736_));
  NA2        o0708(.A(c), .B(ori_ori_n104_), .Y(ori_ori_n737_));
  NO2        o0709(.A(ori_ori_n737_), .B(ori_ori_n349_), .Y(ori_ori_n738_));
  NA3        o0710(.A(ori_ori_n738_), .B(ori_ori_n438_), .C(f), .Y(ori_ori_n739_));
  OR2        o0711(.A(ori_ori_n557_), .B(ori_ori_n463_), .Y(ori_ori_n740_));
  INV        o0712(.A(ori_ori_n740_), .Y(ori_ori_n741_));
  NA2        o0713(.A(ori_ori_n677_), .B(ori_ori_n100_), .Y(ori_ori_n742_));
  NA2        o0714(.A(ori_ori_n742_), .B(ori_ori_n741_), .Y(ori_ori_n743_));
  NA4        o0715(.A(ori_ori_n743_), .B(ori_ori_n739_), .C(ori_ori_n199_), .D(ori_ori_n736_), .Y(ori_ori_n744_));
  NO4        o0716(.A(ori_ori_n744_), .B(ori_ori_n734_), .C(ori_ori_n719_), .D(ori_ori_n709_), .Y(ori_ori_n745_));
  OR2        o0717(.A(ori_ori_n731_), .B(ori_ori_n67_), .Y(ori_ori_n746_));
  NA2        o0718(.A(ori_ori_n697_), .B(o), .Y(ori_ori_n747_));
  AOI210     o0719(.A0(ori_ori_n747_), .A1(ori_ori_n257_), .B0(ori_ori_n746_), .Y(ori_ori_n748_));
  NO2        o0720(.A(ori_ori_n284_), .B(ori_ori_n706_), .Y(ori_ori_n749_));
  NO2        o0721(.A(ori_ori_n120_), .B(ori_ori_n118_), .Y(ori_ori_n750_));
  NO2        o0722(.A(ori_ori_n206_), .B(ori_ori_n200_), .Y(ori_ori_n751_));
  AOI220     o0723(.A0(ori_ori_n751_), .A1(ori_ori_n203_), .B0(ori_ori_n262_), .B1(ori_ori_n750_), .Y(ori_ori_n752_));
  INV        o0724(.A(ori_ori_n752_), .Y(ori_ori_n753_));
  NA2        o0725(.A(e), .B(d), .Y(ori_ori_n754_));
  OAI220     o0726(.A0(ori_ori_n754_), .A1(c), .B0(ori_ori_n276_), .B1(d), .Y(ori_ori_n755_));
  NA3        o0727(.A(ori_ori_n755_), .B(ori_ori_n384_), .C(ori_ori_n436_), .Y(ori_ori_n756_));
  AOI210     o0728(.A0(ori_ori_n442_), .A1(ori_ori_n159_), .B0(ori_ori_n206_), .Y(ori_ori_n757_));
  AOI210     o0729(.A0(ori_ori_n530_), .A1(ori_ori_n295_), .B0(ori_ori_n757_), .Y(ori_ori_n758_));
  NA2        o0730(.A(ori_ori_n249_), .B(ori_ori_n148_), .Y(ori_ori_n759_));
  NA2        o0731(.A(ori_ori_n732_), .B(ori_ori_n759_), .Y(ori_ori_n760_));
  NA3        o0732(.A(ori_ori_n760_), .B(ori_ori_n758_), .C(ori_ori_n756_), .Y(ori_ori_n761_));
  NO4        o0733(.A(ori_ori_n761_), .B(ori_ori_n753_), .C(ori_ori_n749_), .D(ori_ori_n748_), .Y(ori_ori_n762_));
  OR2        o0734(.A(ori_ori_n587_), .B(ori_ori_n194_), .Y(ori_ori_n763_));
  NA2        o0735(.A(ori_ori_n521_), .B(ori_ori_n528_), .Y(ori_ori_n764_));
  NO2        o0736(.A(ori_ori_n701_), .B(ori_ori_n149_), .Y(ori_ori_n765_));
  OAI210     o0737(.A0(ori_ori_n697_), .A1(ori_ori_n759_), .B0(ori_ori_n725_), .Y(ori_ori_n766_));
  NO2        o0738(.A(ori_ori_n766_), .B(ori_ori_n513_), .Y(ori_ori_n767_));
  AOI210     o0739(.A0(ori_ori_n106_), .A1(ori_ori_n105_), .B0(ori_ori_n234_), .Y(ori_ori_n768_));
  NO2        o0740(.A(ori_ori_n768_), .B(ori_ori_n726_), .Y(ori_ori_n769_));
  BUFFER     o0741(.A(ori_ori_n769_), .Y(ori_ori_n770_));
  NOi31      o0742(.An(ori_ori_n467_), .B(ori_ori_n723_), .C(ori_ori_n257_), .Y(ori_ori_n771_));
  NO4        o0743(.A(ori_ori_n771_), .B(ori_ori_n770_), .C(ori_ori_n767_), .D(ori_ori_n765_), .Y(ori_ori_n772_));
  AO220      o0744(.A0(ori_ori_n384_), .A1(ori_ori_n623_), .B0(ori_ori_n154_), .B1(f), .Y(ori_ori_n773_));
  OAI210     o0745(.A0(ori_ori_n773_), .A1(ori_ori_n387_), .B0(ori_ori_n755_), .Y(ori_ori_n774_));
  NO2        o0746(.A(ori_ori_n366_), .B(ori_ori_n64_), .Y(ori_ori_n775_));
  NA2        o0747(.A(ori_ori_n775_), .B(ori_ori_n591_), .Y(ori_ori_n776_));
  AN4        o0748(.A(ori_ori_n776_), .B(ori_ori_n774_), .C(ori_ori_n772_), .D(ori_ori_n763_), .Y(ori_ori_n777_));
  NA4        o0749(.A(ori_ori_n777_), .B(ori_ori_n762_), .C(ori_ori_n745_), .D(ori_ori_n703_), .Y(ori12));
  NO2        o0750(.A(ori_ori_n382_), .B(c), .Y(ori_ori_n779_));
  NO4        o0751(.A(ori_ori_n371_), .B(ori_ori_n226_), .C(ori_ori_n499_), .D(ori_ori_n191_), .Y(ori_ori_n780_));
  NA2        o0752(.A(ori_ori_n780_), .B(ori_ori_n779_), .Y(ori_ori_n781_));
  NA2        o0753(.A(ori_ori_n467_), .B(ori_ori_n775_), .Y(ori_ori_n782_));
  NO2        o0754(.A(ori_ori_n382_), .B(ori_ori_n104_), .Y(ori_ori_n783_));
  NO2        o0755(.A(ori_ori_n711_), .B(ori_ori_n300_), .Y(ori_ori_n784_));
  NO2        o0756(.A(ori_ori_n557_), .B(ori_ori_n320_), .Y(ori_ori_n785_));
  AOI220     o0757(.A0(ori_ori_n785_), .A1(ori_ori_n465_), .B0(ori_ori_n784_), .B1(ori_ori_n783_), .Y(ori_ori_n786_));
  NA4        o0758(.A(ori_ori_n786_), .B(ori_ori_n782_), .C(ori_ori_n781_), .D(ori_ori_n370_), .Y(ori_ori_n787_));
  AOI210     o0759(.A0(ori_ori_n208_), .A1(ori_ori_n289_), .B0(ori_ori_n177_), .Y(ori_ori_n788_));
  OR2        o0760(.A(ori_ori_n788_), .B(ori_ori_n780_), .Y(ori_ori_n789_));
  AOI210     o0761(.A0(ori_ori_n286_), .A1(ori_ori_n330_), .B0(ori_ori_n191_), .Y(ori_ori_n790_));
  OAI210     o0762(.A0(ori_ori_n790_), .A1(ori_ori_n789_), .B0(ori_ori_n344_), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n542_), .B(ori_ori_n236_), .Y(ori_ori_n792_));
  NO2        o0764(.A(ori_ori_n506_), .B(ori_ori_n704_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n135_), .B(ori_ori_n211_), .Y(ori_ori_n794_));
  NA3        o0766(.A(ori_ori_n794_), .B(ori_ori_n214_), .C(i), .Y(ori_ori_n795_));
  NA2        o0767(.A(ori_ori_n795_), .B(ori_ori_n791_), .Y(ori_ori_n796_));
  OR2        o0768(.A(ori_ori_n277_), .B(ori_ori_n783_), .Y(ori_ori_n797_));
  NA2        o0769(.A(ori_ori_n797_), .B(ori_ori_n301_), .Y(ori_ori_n798_));
  NO3        o0770(.A(ori_ori_n118_), .B(ori_ori_n136_), .C(ori_ori_n191_), .Y(ori_ori_n799_));
  NA2        o0771(.A(ori_ori_n799_), .B(ori_ori_n457_), .Y(ori_ori_n800_));
  NA4        o0772(.A(ori_ori_n372_), .B(ori_ori_n364_), .C(ori_ori_n160_), .D(o), .Y(ori_ori_n801_));
  NA3        o0773(.A(ori_ori_n801_), .B(ori_ori_n800_), .C(ori_ori_n798_), .Y(ori_ori_n802_));
  NO3        o0774(.A(ori_ori_n802_), .B(ori_ori_n796_), .C(ori_ori_n787_), .Y(ori_ori_n803_));
  NO2        o0775(.A(ori_ori_n314_), .B(ori_ori_n313_), .Y(ori_ori_n804_));
  INV        o0776(.A(ori_ori_n66_), .Y(ori_ori_n805_));
  NA2        o0777(.A(ori_ori_n476_), .B(ori_ori_n128_), .Y(ori_ori_n806_));
  NOi21      o0778(.An(ori_ori_n33_), .B(ori_ori_n551_), .Y(ori_ori_n807_));
  AOI220     o0779(.A0(ori_ori_n807_), .A1(ori_ori_n806_), .B0(ori_ori_n805_), .B1(ori_ori_n804_), .Y(ori_ori_n808_));
  OAI210     o0780(.A0(ori_ori_n224_), .A1(ori_ori_n44_), .B0(ori_ori_n808_), .Y(ori_ori_n809_));
  INV        o0781(.A(ori_ori_n275_), .Y(ori_ori_n810_));
  NO2        o0782(.A(ori_ori_n48_), .B(ori_ori_n44_), .Y(ori_ori_n811_));
  NO2        o0783(.A(ori_ori_n435_), .B(ori_ori_n260_), .Y(ori_ori_n812_));
  INV        o0784(.A(ori_ori_n812_), .Y(ori_ori_n813_));
  NO2        o0785(.A(ori_ori_n813_), .B(ori_ori_n128_), .Y(ori_ori_n814_));
  INV        o0786(.A(ori_ori_n312_), .Y(ori_ori_n815_));
  NO4        o0787(.A(ori_ori_n815_), .B(ori_ori_n814_), .C(ori_ori_n810_), .D(ori_ori_n809_), .Y(ori_ori_n816_));
  NA2        o0788(.A(ori_ori_n295_), .B(o), .Y(ori_ori_n817_));
  NO2        o0789(.A(ori_ori_n128_), .B(ori_ori_n77_), .Y(ori_ori_n818_));
  OR2        o0790(.A(ori_ori_n818_), .B(ori_ori_n475_), .Y(ori_ori_n819_));
  NA2        o0791(.A(ori_ori_n476_), .B(ori_ori_n322_), .Y(ori_ori_n820_));
  AOI210     o0792(.A0(ori_ori_n820_), .A1(n), .B0(ori_ori_n819_), .Y(ori_ori_n821_));
  NO2        o0793(.A(ori_ori_n821_), .B(ori_ori_n817_), .Y(ori_ori_n822_));
  NO2        o0794(.A(ori_ori_n557_), .B(ori_ori_n429_), .Y(ori_ori_n823_));
  NA3        o0795(.A(ori_ori_n293_), .B(ori_ori_n533_), .C(i), .Y(ori_ori_n824_));
  OAI210     o0796(.A0(ori_ori_n366_), .A1(ori_ori_n266_), .B0(ori_ori_n824_), .Y(ori_ori_n825_));
  OAI220     o0797(.A0(ori_ori_n825_), .A1(ori_ori_n823_), .B0(ori_ori_n566_), .B1(ori_ori_n633_), .Y(ori_ori_n826_));
  NA2        o0798(.A(ori_ori_n515_), .B(ori_ori_n102_), .Y(ori_ori_n827_));
  OR3        o0799(.A(ori_ori_n266_), .B(ori_ori_n362_), .C(f), .Y(ori_ori_n828_));
  NA3        o0800(.A(ori_ori_n533_), .B(ori_ori_n74_), .C(i), .Y(ori_ori_n829_));
  OA220      o0801(.A0(ori_ori_n829_), .A1(ori_ori_n827_), .B0(ori_ori_n828_), .B1(ori_ori_n505_), .Y(ori_ori_n830_));
  NA3        o0802(.A(ori_ori_n278_), .B(ori_ori_n106_), .C(o), .Y(ori_ori_n831_));
  AOI210     o0803(.A0(ori_ori_n564_), .A1(ori_ori_n831_), .B0(m), .Y(ori_ori_n832_));
  OAI210     o0804(.A0(ori_ori_n832_), .A1(ori_ori_n784_), .B0(ori_ori_n277_), .Y(ori_ori_n833_));
  INV        o0805(.A(ori_ori_n578_), .Y(ori_ori_n834_));
  NA2        o0806(.A(ori_ori_n706_), .B(ori_ori_n367_), .Y(ori_ori_n835_));
  INV        o0807(.A(ori_ori_n829_), .Y(ori_ori_n836_));
  AOI220     o0808(.A0(ori_ori_n836_), .A1(ori_ori_n232_), .B0(ori_ori_n835_), .B1(ori_ori_n834_), .Y(ori_ori_n837_));
  NA4        o0809(.A(ori_ori_n837_), .B(ori_ori_n833_), .C(ori_ori_n830_), .D(ori_ori_n826_), .Y(ori_ori_n838_));
  NO2        o0810(.A(ori_ori_n320_), .B(ori_ori_n84_), .Y(ori_ori_n839_));
  OAI210     o0811(.A0(ori_ori_n839_), .A1(ori_ori_n792_), .B0(ori_ori_n212_), .Y(ori_ori_n840_));
  NO2        o0812(.A(ori_ori_n390_), .B(ori_ori_n191_), .Y(ori_ori_n841_));
  AOI220     o0813(.A0(ori_ori_n841_), .A1(ori_ori_n323_), .B0(ori_ori_n797_), .B1(ori_ori_n195_), .Y(ori_ori_n842_));
  AOI220     o0814(.A0(ori_ori_n785_), .A1(ori_ori_n794_), .B0(ori_ori_n504_), .B1(ori_ori_n83_), .Y(ori_ori_n843_));
  NA3        o0815(.A(ori_ori_n843_), .B(ori_ori_n842_), .C(ori_ori_n840_), .Y(ori_ori_n844_));
  OAI210     o0816(.A0(ori_ori_n835_), .A1(ori_ori_n793_), .B0(ori_ori_n465_), .Y(ori_ori_n845_));
  NA2        o0817(.A(ori_ori_n832_), .B(ori_ori_n783_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n545_), .B(ori_ori_n457_), .Y(ori_ori_n847_));
  NA3        o0819(.A(ori_ori_n847_), .B(ori_ori_n846_), .C(ori_ori_n845_), .Y(ori_ori_n848_));
  NO4        o0820(.A(ori_ori_n848_), .B(ori_ori_n844_), .C(ori_ori_n838_), .D(ori_ori_n822_), .Y(ori_ori_n849_));
  NAi31      o0821(.An(ori_ori_n124_), .B(ori_ori_n354_), .C(n), .Y(ori_ori_n850_));
  NO3        o0822(.A(ori_ori_n112_), .B(ori_ori_n291_), .C(ori_ori_n712_), .Y(ori_ori_n851_));
  NO2        o0823(.A(ori_ori_n851_), .B(ori_ori_n850_), .Y(ori_ori_n852_));
  INV        o0824(.A(ori_ori_n852_), .Y(ori_ori_n853_));
  NA2        o0825(.A(ori_ori_n423_), .B(i), .Y(ori_ori_n854_));
  NA2        o0826(.A(ori_ori_n854_), .B(ori_ori_n853_), .Y(ori_ori_n855_));
  NA2        o0827(.A(ori_ori_n206_), .B(ori_ori_n150_), .Y(ori_ori_n856_));
  NO3        o0828(.A(ori_ori_n264_), .B(ori_ori_n372_), .C(ori_ori_n154_), .Y(ori_ori_n857_));
  NOi31      o0829(.An(ori_ori_n856_), .B(ori_ori_n857_), .C(ori_ori_n191_), .Y(ori_ori_n858_));
  NAi21      o0830(.An(ori_ori_n476_), .B(ori_ori_n841_), .Y(ori_ori_n859_));
  NA2        o0831(.A(ori_ori_n414_), .B(o), .Y(ori_ori_n860_));
  NA2        o0832(.A(ori_ori_n860_), .B(ori_ori_n859_), .Y(ori_ori_n861_));
  NA2        o0833(.A(ori_ori_n788_), .B(ori_ori_n779_), .Y(ori_ori_n862_));
  OAI220     o0834(.A0(ori_ori_n785_), .A1(ori_ori_n793_), .B0(ori_ori_n467_), .B1(ori_ori_n360_), .Y(ori_ori_n863_));
  NA3        o0835(.A(ori_ori_n863_), .B(ori_ori_n862_), .C(ori_ori_n527_), .Y(ori_ori_n864_));
  OAI210     o0836(.A0(ori_ori_n788_), .A1(ori_ori_n780_), .B0(ori_ori_n856_), .Y(ori_ori_n865_));
  NA3        o0837(.A(ori_ori_n820_), .B(ori_ori_n419_), .C(ori_ori_n45_), .Y(ori_ori_n866_));
  INV        o0838(.A(ori_ori_n283_), .Y(ori_ori_n867_));
  NA3        o0839(.A(ori_ori_n867_), .B(ori_ori_n866_), .C(ori_ori_n865_), .Y(ori_ori_n868_));
  OR2        o0840(.A(ori_ori_n868_), .B(ori_ori_n864_), .Y(ori_ori_n869_));
  NO4        o0841(.A(ori_ori_n869_), .B(ori_ori_n861_), .C(ori_ori_n858_), .D(ori_ori_n855_), .Y(ori_ori_n870_));
  NA4        o0842(.A(ori_ori_n870_), .B(ori_ori_n849_), .C(ori_ori_n816_), .D(ori_ori_n803_), .Y(ori13));
  NAi32      o0843(.An(d), .Bn(c), .C(e), .Y(ori_ori_n872_));
  AN2        o0844(.A(d), .B(c), .Y(ori_ori_n873_));
  NA2        o0845(.A(ori_ori_n873_), .B(ori_ori_n104_), .Y(ori_ori_n874_));
  NAi32      o0846(.An(f), .Bn(e), .C(c), .Y(ori_ori_n875_));
  NO3        o0847(.A(m), .B(i), .C(h), .Y(ori_ori_n876_));
  NA3        o0848(.A(k), .B(j), .C(i), .Y(ori_ori_n877_));
  NO2        o0849(.A(f), .B(c), .Y(ori_ori_n878_));
  NOi21      o0850(.An(ori_ori_n878_), .B(ori_ori_n371_), .Y(ori_ori_n879_));
  AN3        o0851(.A(o), .B(f), .C(c), .Y(ori_ori_n880_));
  NA3        o0852(.A(l), .B(k), .C(j), .Y(ori_ori_n881_));
  NA2        o0853(.A(i), .B(h), .Y(ori_ori_n882_));
  NO3        o0854(.A(ori_ori_n882_), .B(ori_ori_n881_), .C(ori_ori_n118_), .Y(ori_ori_n883_));
  NO3        o0855(.A(ori_ori_n125_), .B(ori_ori_n248_), .C(ori_ori_n191_), .Y(ori_ori_n884_));
  NA3        o0856(.A(c), .B(b), .C(a), .Y(ori_ori_n885_));
  NO2        o0857(.A(ori_ori_n453_), .B(ori_ori_n510_), .Y(ori_ori_n886_));
  NA4        o0858(.A(ori_ori_n81_), .B(ori_ori_n80_), .C(o), .D(ori_ori_n190_), .Y(ori_ori_n887_));
  NA4        o0859(.A(ori_ori_n494_), .B(m), .C(ori_ori_n101_), .D(ori_ori_n190_), .Y(ori_ori_n888_));
  NA3        o0860(.A(ori_ori_n888_), .B(ori_ori_n315_), .C(ori_ori_n887_), .Y(ori_ori_n889_));
  NO2        o0861(.A(ori_ori_n889_), .B(ori_ori_n886_), .Y(ori_ori_n890_));
  NOi41      o0862(.An(ori_ori_n675_), .B(ori_ori_n717_), .C(ori_ori_n707_), .D(ori_ori_n603_), .Y(ori_ori_n891_));
  OAI220     o0863(.A0(ori_ori_n891_), .A1(ori_ori_n578_), .B0(ori_ori_n890_), .B1(ori_ori_n503_), .Y(ori_ori_n892_));
  NOi31      o0864(.An(m), .B(n), .C(f), .Y(ori_ori_n893_));
  NA2        o0865(.A(ori_ori_n893_), .B(ori_ori_n50_), .Y(ori_ori_n894_));
  AN2        o0866(.A(e), .B(c), .Y(ori_ori_n895_));
  NA2        o0867(.A(ori_ori_n895_), .B(a), .Y(ori_ori_n896_));
  OAI220     o0868(.A0(ori_ori_n896_), .A1(ori_ori_n894_), .B0(ori_ori_n740_), .B1(ori_ori_n359_), .Y(ori_ori_n897_));
  NA2        o0869(.A(ori_ori_n436_), .B(l), .Y(ori_ori_n898_));
  NO2        o0870(.A(ori_ori_n80_), .B(o), .Y(ori_ori_n899_));
  NO4        o0871(.A(ori_ori_n897_), .B(ori_ori_n892_), .C(ori_ori_n688_), .D(ori_ori_n484_), .Y(ori_ori_n900_));
  NA2        o0872(.A(c), .B(b), .Y(ori_ori_n901_));
  NO2        o0873(.A(ori_ori_n590_), .B(ori_ori_n901_), .Y(ori_ori_n902_));
  OAI210     o0874(.A0(ori_ori_n723_), .A1(ori_ori_n699_), .B0(ori_ori_n351_), .Y(ori_ori_n903_));
  OAI210     o0875(.A0(ori_ori_n903_), .A1(ori_ori_n724_), .B0(ori_ori_n902_), .Y(ori_ori_n904_));
  NA3        o0876(.A(ori_ori_n360_), .B(ori_ori_n481_), .C(f), .Y(ori_ori_n905_));
  NA2        o0877(.A(ori_ori_n235_), .B(ori_ori_n107_), .Y(ori_ori_n906_));
  OAI210     o0878(.A0(ori_ori_n906_), .A1(ori_ori_n251_), .B0(o), .Y(ori_ori_n907_));
  NAi21      o0879(.An(f), .B(d), .Y(ori_ori_n908_));
  NO2        o0880(.A(ori_ori_n908_), .B(ori_ori_n885_), .Y(ori_ori_n909_));
  INV        o0881(.A(ori_ori_n909_), .Y(ori_ori_n910_));
  NO2        o0882(.A(ori_ori_n907_), .B(ori_ori_n910_), .Y(ori_ori_n911_));
  AOI210     o0883(.A0(ori_ori_n911_), .A1(ori_ori_n102_), .B0(ori_ori_n1156_), .Y(ori_ori_n912_));
  NA3        o0884(.A(ori_ori_n768_), .B(ori_ori_n898_), .C(ori_ori_n403_), .Y(ori_ori_n913_));
  NA2        o0885(.A(ori_ori_n375_), .B(ori_ori_n909_), .Y(ori_ori_n914_));
  NA4        o0886(.A(ori_ori_n914_), .B(ori_ori_n912_), .C(ori_ori_n904_), .D(ori_ori_n900_), .Y(ori00));
  NA2        o0887(.A(ori_ori_n438_), .B(f), .Y(ori_ori_n916_));
  OAI210     o0888(.A0(ori_ori_n851_), .A1(ori_ori_n39_), .B0(ori_ori_n547_), .Y(ori_ori_n917_));
  NA3        o0889(.A(ori_ori_n917_), .B(ori_ori_n231_), .C(n), .Y(ori_ori_n918_));
  AOI210     o0890(.A0(ori_ori_n918_), .A1(ori_ori_n916_), .B0(ori_ori_n874_), .Y(ori_ori_n919_));
  NO2        o0891(.A(ori_ori_n919_), .B(ori_ori_n601_), .Y(ori_ori_n920_));
  INV        o0892(.A(ori_ori_n771_), .Y(ori_ori_n921_));
  NO4        o0893(.A(ori_ori_n420_), .B(ori_ori_n303_), .C(ori_ori_n901_), .D(ori_ori_n58_), .Y(ori_ori_n922_));
  NA3        o0894(.A(ori_ori_n324_), .B(ori_ori_n198_), .C(o), .Y(ori_ori_n923_));
  NO2        o0895(.A(h), .B(o), .Y(ori_ori_n924_));
  OAI220     o0896(.A0(ori_ori_n453_), .A1(ori_ori_n510_), .B0(ori_ori_n85_), .B1(ori_ori_n84_), .Y(ori_ori_n925_));
  NA2        o0897(.A(ori_ori_n925_), .B(ori_ori_n460_), .Y(ori_ori_n926_));
  AOI220     o0898(.A0(ori_ori_n272_), .A1(ori_ori_n220_), .B0(ori_ori_n156_), .B1(ori_ori_n132_), .Y(ori_ori_n927_));
  NA2        o0899(.A(ori_ori_n927_), .B(ori_ori_n926_), .Y(ori_ori_n928_));
  NO3        o0900(.A(ori_ori_n928_), .B(ori_ori_n922_), .C(ori_ori_n238_), .Y(ori_ori_n929_));
  NA2        o0901(.A(ori_ori_n220_), .B(ori_ori_n295_), .Y(ori_ori_n930_));
  NA2        o0902(.A(ori_ori_n930_), .B(ori_ori_n138_), .Y(ori_ori_n931_));
  NO2        o0903(.A(ori_ori_n931_), .B(ori_ori_n446_), .Y(ori_ori_n932_));
  AN3        o0904(.A(ori_ori_n932_), .B(ori_ori_n929_), .C(ori_ori_n921_), .Y(ori_ori_n933_));
  NA2        o0905(.A(ori_ori_n460_), .B(ori_ori_n95_), .Y(ori_ori_n934_));
  NA3        o0906(.A(ori_ori_n893_), .B(ori_ori_n515_), .C(ori_ori_n397_), .Y(ori_ori_n935_));
  NA3        o0907(.A(ori_ori_n935_), .B(ori_ori_n934_), .C(ori_ori_n215_), .Y(ori_ori_n936_));
  NA2        o0908(.A(ori_ori_n889_), .B(ori_ori_n460_), .Y(ori_ori_n937_));
  NA4        o0909(.A(ori_ori_n550_), .B(ori_ori_n182_), .C(ori_ori_n198_), .D(ori_ori_n147_), .Y(ori_ori_n938_));
  NA2        o0910(.A(ori_ori_n938_), .B(ori_ori_n937_), .Y(ori_ori_n939_));
  OAI210     o0911(.A0(ori_ori_n396_), .A1(ori_ori_n108_), .B0(ori_ori_n726_), .Y(ori_ori_n940_));
  NA2        o0912(.A(ori_ori_n940_), .B(ori_ori_n913_), .Y(ori_ori_n941_));
  NO2        o0913(.A(ori_ori_n194_), .B(ori_ori_n191_), .Y(ori_ori_n942_));
  NA2        o0914(.A(n), .B(e), .Y(ori_ori_n943_));
  NO2        o0915(.A(ori_ori_n943_), .B(ori_ori_n130_), .Y(ori_ori_n944_));
  AOI220     o0916(.A0(ori_ori_n944_), .A1(ori_ori_n243_), .B0(ori_ori_n710_), .B1(ori_ori_n942_), .Y(ori_ori_n945_));
  OAI210     o0917(.A0(ori_ori_n304_), .A1(ori_ori_n268_), .B0(ori_ori_n377_), .Y(ori_ori_n946_));
  NA3        o0918(.A(ori_ori_n946_), .B(ori_ori_n945_), .C(ori_ori_n941_), .Y(ori_ori_n947_));
  NA2        o0919(.A(ori_ori_n944_), .B(ori_ori_n714_), .Y(ori_ori_n948_));
  NO2        o0920(.A(ori_ori_n62_), .B(h), .Y(ori_ori_n949_));
  NA2        o0921(.A(ori_ori_n948_), .B(ori_ori_n728_), .Y(ori_ori_n950_));
  NO4        o0922(.A(ori_ori_n950_), .B(ori_ori_n947_), .C(ori_ori_n939_), .D(ori_ori_n936_), .Y(ori_ori_n951_));
  NA2        o0923(.A(ori_ori_n700_), .B(ori_ori_n632_), .Y(ori_ori_n952_));
  NA4        o0924(.A(ori_ori_n952_), .B(ori_ori_n951_), .C(ori_ori_n933_), .D(ori_ori_n920_), .Y(ori01));
  NO2        o0925(.A(ori_ori_n411_), .B(ori_ori_n246_), .Y(ori_ori_n954_));
  NA2        o0926(.A(ori_ori_n335_), .B(i), .Y(ori_ori_n955_));
  NA3        o0927(.A(ori_ori_n955_), .B(ori_ori_n954_), .C(ori_ori_n862_), .Y(ori_ori_n956_));
  NA2        o0928(.A(ori_ori_n504_), .B(ori_ori_n83_), .Y(ori_ori_n957_));
  NA2        o0929(.A(ori_ori_n476_), .B(ori_ori_n242_), .Y(ori_ori_n958_));
  NA2        o0930(.A(ori_ori_n812_), .B(ori_ori_n958_), .Y(ori_ori_n959_));
  NA3        o0931(.A(ori_ori_n959_), .B(ori_ori_n957_), .C(ori_ori_n764_), .Y(ori_ori_n960_));
  NA2        o0932(.A(ori_ori_n44_), .B(f), .Y(ori_ori_n961_));
  NA2        o0933(.A(ori_ori_n596_), .B(ori_ori_n90_), .Y(ori_ori_n962_));
  NO2        o0934(.A(ori_ori_n962_), .B(ori_ori_n961_), .Y(ori_ori_n963_));
  OR2        o0935(.A(ori_ori_n558_), .B(ori_ori_n315_), .Y(ori_ori_n964_));
  NAi41      o0936(.An(ori_ori_n146_), .B(ori_ori_n964_), .C(ori_ori_n938_), .D(ori_ori_n752_), .Y(ori_ori_n965_));
  NO3        o0937(.A(ori_ori_n657_), .B(ori_ori_n565_), .C(ori_ori_n440_), .Y(ori_ori_n966_));
  NA4        o0938(.A(ori_ori_n596_), .B(ori_ori_n90_), .C(ori_ori_n44_), .D(ori_ori_n190_), .Y(ori_ori_n967_));
  OA220      o0939(.A0(ori_ori_n967_), .A1(ori_ori_n561_), .B0(ori_ori_n171_), .B1(ori_ori_n169_), .Y(ori_ori_n968_));
  NA2        o0940(.A(ori_ori_n968_), .B(ori_ori_n966_), .Y(ori_ori_n969_));
  NO4        o0941(.A(ori_ori_n969_), .B(ori_ori_n965_), .C(ori_ori_n960_), .D(ori_ori_n956_), .Y(ori_ori_n970_));
  INV        o0942(.A(ori_ori_n923_), .Y(ori_ori_n971_));
  NA2        o0943(.A(ori_ori_n971_), .B(ori_ori_n457_), .Y(ori_ori_n972_));
  AOI210     o0944(.A0(ori_ori_n180_), .A1(ori_ori_n82_), .B0(ori_ori_n190_), .Y(ori_ori_n973_));
  OAI210     o0945(.A0(ori_ori_n678_), .A1(ori_ori_n360_), .B0(ori_ori_n973_), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n974_), .B(ori_ori_n972_), .Y(ori_ori_n975_));
  NA2        o0947(.A(ori_ori_n509_), .B(ori_ori_n106_), .Y(ori_ori_n976_));
  INV        o0948(.A(ori_ori_n976_), .Y(ori_ori_n977_));
  NA2        o0949(.A(ori_ori_n245_), .B(ori_ori_n171_), .Y(ori_ori_n978_));
  NA2        o0950(.A(ori_ori_n978_), .B(ori_ori_n559_), .Y(ori_ori_n979_));
  OAI210     o0951(.A0(ori_ori_n963_), .A1(ori_ori_n280_), .B0(ori_ori_n566_), .Y(ori_ori_n980_));
  NA3        o0952(.A(ori_ori_n980_), .B(ori_ori_n979_), .C(ori_ori_n659_), .Y(ori_ori_n981_));
  NO3        o0953(.A(ori_ori_n981_), .B(ori_ori_n977_), .C(ori_ori_n975_), .Y(ori_ori_n982_));
  NA3        o0954(.A(ori_ori_n512_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n983_));
  NO2        o0955(.A(ori_ori_n983_), .B(ori_ori_n180_), .Y(ori_ori_n984_));
  INV        o0956(.A(ori_ori_n984_), .Y(ori_ori_n985_));
  OR3        o0957(.A(ori_ori_n962_), .B(ori_ori_n513_), .C(ori_ori_n961_), .Y(ori_ori_n986_));
  NO2        o0958(.A(ori_ori_n967_), .B(ori_ori_n827_), .Y(ori_ori_n987_));
  NO2        o0959(.A(ori_ori_n183_), .B(ori_ori_n100_), .Y(ori_ori_n988_));
  NO2        o0960(.A(ori_ori_n988_), .B(ori_ori_n987_), .Y(ori_ori_n989_));
  NA4        o0961(.A(ori_ori_n989_), .B(ori_ori_n986_), .C(ori_ori_n985_), .D(ori_ori_n631_), .Y(ori_ori_n990_));
  NA2        o0962(.A(ori_ori_n490_), .B(ori_ori_n488_), .Y(ori_ori_n991_));
  NO3        o0963(.A(ori_ori_n73_), .B(ori_ori_n260_), .C(ori_ori_n44_), .Y(ori_ori_n992_));
  NA2        o0964(.A(ori_ori_n992_), .B(ori_ori_n475_), .Y(ori_ori_n993_));
  NA3        o0965(.A(ori_ori_n993_), .B(ori_ori_n991_), .C(ori_ori_n562_), .Y(ori_ori_n994_));
  NO2        o0966(.A(ori_ori_n315_), .B(ori_ori_n66_), .Y(ori_ori_n995_));
  INV        o0967(.A(ori_ori_n995_), .Y(ori_ori_n996_));
  NA2        o0968(.A(ori_ori_n992_), .B(ori_ori_n681_), .Y(ori_ori_n997_));
  NA3        o0969(.A(ori_ori_n997_), .B(ori_ori_n996_), .C(ori_ori_n327_), .Y(ori_ori_n998_));
  NO3        o0970(.A(ori_ori_n998_), .B(ori_ori_n994_), .C(ori_ori_n990_), .Y(ori_ori_n999_));
  INV        o0971(.A(ori_ori_n119_), .Y(ori_ori_n1000_));
  NO3        o0972(.A(ori_ori_n882_), .B(ori_ori_n155_), .C(ori_ori_n80_), .Y(ori_ori_n1001_));
  AOI220     o0973(.A0(ori_ori_n1001_), .A1(ori_ori_n1000_), .B0(ori_ori_n992_), .B1(ori_ori_n818_), .Y(ori_ori_n1002_));
  INV        o0974(.A(ori_ori_n1002_), .Y(ori_ori_n1003_));
  NO2        o0975(.A(ori_ori_n523_), .B(ori_ori_n522_), .Y(ori_ori_n1004_));
  NO4        o0976(.A(ori_ori_n882_), .B(ori_ori_n1004_), .C(ori_ori_n153_), .D(ori_ori_n80_), .Y(ori_ori_n1005_));
  NO3        o0977(.A(ori_ori_n1005_), .B(ori_ori_n1003_), .C(ori_ori_n541_), .Y(ori_ori_n1006_));
  NA4        o0978(.A(ori_ori_n1006_), .B(ori_ori_n999_), .C(ori_ori_n982_), .D(ori_ori_n970_), .Y(ori06));
  NO2        o0979(.A(ori_ori_n200_), .B(ori_ori_n96_), .Y(ori_ori_n1008_));
  OAI210     o0980(.A0(ori_ori_n1008_), .A1(ori_ori_n1001_), .B0(ori_ori_n323_), .Y(ori_ori_n1009_));
  INV        o0981(.A(ori_ori_n676_), .Y(ori_ori_n1010_));
  OR2        o0982(.A(ori_ori_n1010_), .B(ori_ori_n740_), .Y(ori_ori_n1011_));
  NA2        o0983(.A(ori_ori_n1011_), .B(ori_ori_n1009_), .Y(ori_ori_n1012_));
  NO3        o0984(.A(ori_ori_n1012_), .B(ori_ori_n994_), .C(ori_ori_n230_), .Y(ori_ori_n1013_));
  NO2        o0985(.A(ori_ori_n260_), .B(ori_ori_n44_), .Y(ori_ori_n1014_));
  NA2        o0986(.A(ori_ori_n1014_), .B(ori_ori_n819_), .Y(ori_ori_n1015_));
  NA2        o0987(.A(ori_ori_n1014_), .B(ori_ori_n479_), .Y(ori_ori_n1016_));
  AOI210     o0988(.A0(ori_ori_n1016_), .A1(ori_ori_n1015_), .B0(ori_ori_n289_), .Y(ori_ori_n1017_));
  NO2        o0989(.A(ori_ori_n82_), .B(ori_ori_n39_), .Y(ori_ori_n1018_));
  NA2        o0990(.A(ori_ori_n1018_), .B(ori_ori_n544_), .Y(ori_ori_n1019_));
  NO2        o0991(.A(ori_ori_n516_), .B(ori_ori_n894_), .Y(ori_ori_n1020_));
  NO2        o0992(.A(ori_ori_n391_), .B(ori_ori_n221_), .Y(ori_ori_n1021_));
  NO2        o0993(.A(ori_ori_n1021_), .B(ori_ori_n1020_), .Y(ori_ori_n1022_));
  NA2        o0994(.A(ori_ori_n1022_), .B(ori_ori_n1019_), .Y(ori_ori_n1023_));
  NO2        o0995(.A(ori_ori_n624_), .B(ori_ori_n313_), .Y(ori_ori_n1024_));
  INV        o0996(.A(ori_ori_n566_), .Y(ori_ori_n1025_));
  NOi21      o0997(.An(ori_ori_n1024_), .B(ori_ori_n1025_), .Y(ori_ori_n1026_));
  AN2        o0998(.A(ori_ori_n807_), .B(ori_ori_n546_), .Y(ori_ori_n1027_));
  NO4        o0999(.A(ori_ori_n1027_), .B(ori_ori_n1026_), .C(ori_ori_n1023_), .D(ori_ori_n1017_), .Y(ori_ori_n1028_));
  OAI220     o1000(.A0(ori_ori_n587_), .A1(ori_ori_n221_), .B0(ori_ori_n439_), .B1(ori_ori_n442_), .Y(ori_ori_n1029_));
  INV        o1001(.A(k), .Y(ori_ori_n1030_));
  NO3        o1002(.A(ori_ori_n1030_), .B(ori_ori_n510_), .C(j), .Y(ori_ori_n1031_));
  NOi21      o1003(.An(ori_ori_n1031_), .B(ori_ori_n561_), .Y(ori_ori_n1032_));
  NO3        o1004(.A(ori_ori_n1032_), .B(ori_ori_n1029_), .C(ori_ori_n897_), .Y(ori_ori_n1033_));
  NA3        o1005(.A(ori_ori_n667_), .B(ori_ori_n666_), .C(ori_ori_n365_), .Y(ori_ori_n1034_));
  NAi31      o1006(.An(ori_ori_n624_), .B(ori_ori_n1034_), .C(ori_ori_n179_), .Y(ori_ori_n1035_));
  NA2        o1007(.A(ori_ori_n1035_), .B(ori_ori_n1033_), .Y(ori_ori_n1036_));
  OR3        o1008(.A(ori_ori_n1010_), .B(ori_ori_n656_), .C(ori_ori_n463_), .Y(ori_ori_n1037_));
  NA2        o1009(.A(ori_ori_n490_), .B(ori_ori_n377_), .Y(ori_ori_n1038_));
  NA2        o1010(.A(ori_ori_n1031_), .B(ori_ori_n663_), .Y(ori_ori_n1039_));
  NA3        o1011(.A(ori_ori_n1039_), .B(ori_ori_n1038_), .C(ori_ori_n1037_), .Y(ori_ori_n1040_));
  AN2        o1012(.A(ori_ori_n780_), .B(ori_ori_n779_), .Y(ori_ori_n1041_));
  NO3        o1013(.A(ori_ori_n1041_), .B(ori_ori_n432_), .C(ori_ori_n414_), .Y(ori_ori_n1042_));
  NA2        o1014(.A(ori_ori_n1042_), .B(ori_ori_n997_), .Y(ori_ori_n1043_));
  NAi21      o1015(.An(j), .B(i), .Y(ori_ori_n1044_));
  NO4        o1016(.A(ori_ori_n1004_), .B(ori_ori_n1044_), .C(ori_ori_n371_), .D(ori_ori_n209_), .Y(ori_ori_n1045_));
  NO4        o1017(.A(ori_ori_n1045_), .B(ori_ori_n1043_), .C(ori_ori_n1040_), .D(ori_ori_n1036_), .Y(ori_ori_n1046_));
  NA4        o1018(.A(ori_ori_n1046_), .B(ori_ori_n1028_), .C(ori_ori_n1013_), .D(ori_ori_n1006_), .Y(ori07));
  NAi32      o1019(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1048_));
  NO3        o1020(.A(ori_ori_n1048_), .B(o), .C(f), .Y(ori_ori_n1049_));
  NOi31      o1021(.An(n), .B(m), .C(b), .Y(ori_ori_n1050_));
  NO3        o1022(.A(ori_ori_n118_), .B(ori_ori_n379_), .C(h), .Y(ori_ori_n1051_));
  NO3        o1023(.A(n), .B(m), .C(h), .Y(ori_ori_n1052_));
  NO2        o1024(.A(ori_ori_n875_), .B(ori_ori_n371_), .Y(ori_ori_n1053_));
  INV        o1025(.A(ori_ori_n1053_), .Y(ori_ori_n1054_));
  NO2        o1026(.A(ori_ori_n877_), .B(ori_ori_n263_), .Y(ori_ori_n1055_));
  NA2        o1027(.A(ori_ori_n464_), .B(ori_ori_n74_), .Y(ori_ori_n1056_));
  NA2        o1028(.A(ori_ori_n949_), .B(ori_ori_n255_), .Y(ori_ori_n1057_));
  NA3        o1029(.A(ori_ori_n1057_), .B(ori_ori_n1056_), .C(ori_ori_n1054_), .Y(ori_ori_n1058_));
  NO2        o1030(.A(ori_ori_n1058_), .B(ori_ori_n1049_), .Y(ori_ori_n1059_));
  NO3        o1031(.A(e), .B(d), .C(c), .Y(ori_ori_n1060_));
  NO2        o1032(.A(ori_ori_n118_), .B(ori_ori_n191_), .Y(ori_ori_n1061_));
  NA2        o1033(.A(ori_ori_n1061_), .B(ori_ori_n1060_), .Y(ori_ori_n1062_));
  INV        o1034(.A(ori_ori_n1062_), .Y(ori_ori_n1063_));
  NA3        o1035(.A(ori_ori_n584_), .B(ori_ori_n570_), .C(ori_ori_n101_), .Y(ori_ori_n1064_));
  NO2        o1036(.A(ori_ori_n1064_), .B(ori_ori_n44_), .Y(ori_ori_n1065_));
  NO2        o1037(.A(l), .B(k), .Y(ori_ori_n1066_));
  NO3        o1038(.A(ori_ori_n371_), .B(d), .C(c), .Y(ori_ori_n1067_));
  NO2        o1039(.A(ori_ori_n1065_), .B(ori_ori_n1063_), .Y(ori_ori_n1068_));
  NO2        o1040(.A(o), .B(c), .Y(ori_ori_n1069_));
  NO2        o1041(.A(ori_ori_n382_), .B(a), .Y(ori_ori_n1070_));
  NA2        o1042(.A(ori_ori_n1070_), .B(ori_ori_n102_), .Y(ori_ori_n1071_));
  NO2        o1043(.A(ori_ori_n630_), .B(ori_ori_n165_), .Y(ori_ori_n1072_));
  NOi31      o1044(.An(m), .B(n), .C(b), .Y(ori_ori_n1073_));
  NOi31      o1045(.An(f), .B(d), .C(c), .Y(ori_ori_n1074_));
  NA2        o1046(.A(ori_ori_n1074_), .B(ori_ori_n1073_), .Y(ori_ori_n1075_));
  INV        o1047(.A(ori_ori_n1075_), .Y(ori_ori_n1076_));
  NO2        o1048(.A(ori_ori_n1076_), .B(ori_ori_n1072_), .Y(ori_ori_n1077_));
  NA2        o1049(.A(ori_ori_n880_), .B(ori_ori_n398_), .Y(ori_ori_n1078_));
  NO2        o1050(.A(ori_ori_n1078_), .B(ori_ori_n371_), .Y(ori_ori_n1079_));
  NO3        o1051(.A(ori_ori_n40_), .B(i), .C(h), .Y(ori_ori_n1080_));
  NO2        o1052(.A(ori_ori_n876_), .B(ori_ori_n1079_), .Y(ori_ori_n1081_));
  AN3        o1053(.A(ori_ori_n1081_), .B(ori_ori_n1077_), .C(ori_ori_n1071_), .Y(ori_ori_n1082_));
  NA2        o1054(.A(ori_ori_n1050_), .B(ori_ori_n321_), .Y(ori_ori_n1083_));
  INV        o1055(.A(ori_ori_n1083_), .Y(ori_ori_n1084_));
  INV        o1056(.A(ori_ori_n883_), .Y(ori_ori_n1085_));
  NAi21      o1057(.An(ori_ori_n1084_), .B(ori_ori_n1085_), .Y(ori_ori_n1086_));
  NO4        o1058(.A(ori_ori_n118_), .B(o), .C(f), .D(e), .Y(ori_ori_n1087_));
  NA2        o1059(.A(ori_ori_n1052_), .B(ori_ori_n1066_), .Y(ori_ori_n1088_));
  INV        o1060(.A(ori_ori_n1088_), .Y(ori_ori_n1089_));
  OR3        o1061(.A(ori_ori_n463_), .B(ori_ori_n462_), .C(ori_ori_n101_), .Y(ori_ori_n1090_));
  NA2        o1062(.A(ori_ori_n893_), .B(ori_ori_n349_), .Y(ori_ori_n1091_));
  NO2        o1063(.A(ori_ori_n1091_), .B(ori_ori_n364_), .Y(ori_ori_n1092_));
  AO210      o1064(.A0(ori_ori_n1092_), .A1(ori_ori_n104_), .B0(ori_ori_n1089_), .Y(ori_ori_n1093_));
  NO2        o1065(.A(ori_ori_n1093_), .B(ori_ori_n1086_), .Y(ori_ori_n1094_));
  NA4        o1066(.A(ori_ori_n1094_), .B(ori_ori_n1082_), .C(ori_ori_n1068_), .D(ori_ori_n1059_), .Y(ori_ori_n1095_));
  NO2        o1067(.A(ori_ori_n901_), .B(ori_ori_n99_), .Y(ori_ori_n1096_));
  NO2        o1068(.A(ori_ori_n332_), .B(j), .Y(ori_ori_n1097_));
  NA2        o1069(.A(ori_ori_n1080_), .B(ori_ori_n893_), .Y(ori_ori_n1098_));
  NA2        o1070(.A(ori_ori_n879_), .B(ori_ori_n134_), .Y(ori_ori_n1099_));
  NA2        o1071(.A(ori_ori_n1099_), .B(ori_ori_n1098_), .Y(ori_ori_n1100_));
  NA2        o1072(.A(ori_ori_n1097_), .B(ori_ori_n143_), .Y(ori_ori_n1101_));
  INV        o1073(.A(ori_ori_n1101_), .Y(ori_ori_n1102_));
  NO2        o1074(.A(ori_ori_n1102_), .B(ori_ori_n1100_), .Y(ori_ori_n1103_));
  INV        o1075(.A(ori_ori_n48_), .Y(ori_ori_n1104_));
  NA2        o1076(.A(ori_ori_n1104_), .B(ori_ori_n924_), .Y(ori_ori_n1105_));
  INV        o1077(.A(ori_ori_n1105_), .Y(ori_ori_n1106_));
  NO2        o1078(.A(ori_ori_n200_), .B(ori_ori_n155_), .Y(ori_ori_n1107_));
  NO2        o1079(.A(ori_ori_n1090_), .B(ori_ori_n300_), .Y(ori_ori_n1108_));
  NO3        o1080(.A(ori_ori_n1108_), .B(ori_ori_n1107_), .C(ori_ori_n1106_), .Y(ori_ori_n1109_));
  NA2        o1081(.A(ori_ori_n1096_), .B(f), .Y(ori_ori_n1110_));
  NO2        o1082(.A(ori_ori_n1151_), .B(ori_ori_n1110_), .Y(ori_ori_n1111_));
  NO2        o1083(.A(ori_ori_n1044_), .B(ori_ori_n153_), .Y(ori_ori_n1112_));
  NOi21      o1084(.An(d), .B(f), .Y(ori_ori_n1113_));
  NA2        o1085(.A(h), .B(ori_ori_n1112_), .Y(ori_ori_n1114_));
  INV        o1086(.A(ori_ori_n1114_), .Y(ori_ori_n1115_));
  NO2        o1087(.A(ori_ori_n1115_), .B(ori_ori_n1111_), .Y(ori_ori_n1116_));
  NA3        o1088(.A(ori_ori_n1116_), .B(ori_ori_n1109_), .C(ori_ori_n1103_), .Y(ori_ori_n1117_));
  NA2        o1089(.A(h), .B(ori_ori_n1055_), .Y(ori_ori_n1118_));
  OAI210     o1090(.A0(ori_ori_n1087_), .A1(ori_ori_n1050_), .B0(ori_ori_n737_), .Y(ori_ori_n1119_));
  NO2        o1091(.A(ori_ori_n872_), .B(ori_ori_n118_), .Y(ori_ori_n1120_));
  NA2        o1092(.A(ori_ori_n1120_), .B(ori_ori_n529_), .Y(ori_ori_n1121_));
  NA3        o1093(.A(ori_ori_n1121_), .B(ori_ori_n1119_), .C(ori_ori_n1118_), .Y(ori_ori_n1122_));
  NA2        o1094(.A(ori_ori_n1069_), .B(ori_ori_n1113_), .Y(ori_ori_n1123_));
  NO2        o1095(.A(ori_ori_n1123_), .B(m), .Y(ori_ori_n1124_));
  NA2        o1096(.A(ori_ori_n884_), .B(ori_ori_n198_), .Y(ori_ori_n1125_));
  NO2        o1097(.A(ori_ori_n135_), .B(ori_ori_n160_), .Y(ori_ori_n1126_));
  OAI210     o1098(.A0(ori_ori_n1126_), .A1(ori_ori_n99_), .B0(ori_ori_n1073_), .Y(ori_ori_n1127_));
  NA2        o1099(.A(ori_ori_n1127_), .B(ori_ori_n1125_), .Y(ori_ori_n1128_));
  NO3        o1100(.A(ori_ori_n1128_), .B(ori_ori_n1124_), .C(ori_ori_n1122_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(f), .B(e), .Y(ori_ori_n1130_));
  NA2        o1102(.A(ori_ori_n1130_), .B(ori_ori_n347_), .Y(ori_ori_n1131_));
  NO2        o1103(.A(ori_ori_n118_), .B(ori_ori_n1131_), .Y(ori_ori_n1132_));
  INV        o1104(.A(ori_ori_n1132_), .Y(ori_ori_n1133_));
  INV        o1105(.A(ori_ori_n1067_), .Y(ori_ori_n1134_));
  INV        o1106(.A(ori_ori_n899_), .Y(ori_ori_n1135_));
  OAI210     o1107(.A0(ori_ori_n1135_), .A1(ori_ori_n63_), .B0(ori_ori_n1134_), .Y(ori_ori_n1136_));
  OR2        o1108(.A(h), .B(ori_ori_n462_), .Y(ori_ori_n1137_));
  NO2        o1109(.A(ori_ori_n1137_), .B(ori_ori_n153_), .Y(ori_ori_n1138_));
  NO2        o1110(.A(ori_ori_n48_), .B(l), .Y(ori_ori_n1139_));
  INV        o1111(.A(ori_ori_n416_), .Y(ori_ori_n1140_));
  NA2        o1112(.A(ori_ori_n1140_), .B(ori_ori_n1139_), .Y(ori_ori_n1141_));
  INV        o1113(.A(ori_ori_n1141_), .Y(ori_ori_n1142_));
  NO3        o1114(.A(ori_ori_n1142_), .B(ori_ori_n1138_), .C(ori_ori_n1136_), .Y(ori_ori_n1143_));
  NA3        o1115(.A(ori_ori_n1143_), .B(ori_ori_n1133_), .C(ori_ori_n1129_), .Y(ori_ori_n1144_));
  NA3        o1116(.A(ori_ori_n811_), .B(ori_ori_n121_), .C(ori_ori_n45_), .Y(ori_ori_n1145_));
  NO2        o1117(.A(ori_ori_n1091_), .B(d), .Y(ori_ori_n1146_));
  NA3        o1118(.A(ori_ori_n1152_), .B(ori_ori_n1153_), .C(ori_ori_n1145_), .Y(ori_ori_n1147_));
  OR4        o1119(.A(ori_ori_n1147_), .B(ori_ori_n1144_), .C(ori_ori_n1117_), .D(ori_ori_n1095_), .Y(ori04));
  INV        o1120(.A(ori_ori_n102_), .Y(ori_ori_n1151_));
  INV        o1121(.A(ori_ori_n1146_), .Y(ori_ori_n1152_));
  INV        o1122(.A(ori_ori_n1051_), .Y(ori_ori_n1153_));
  INV        o1123(.A(ori_ori_n265_), .Y(ori_ori_n1154_));
  INV        o1124(.A(ori_ori_n89_), .Y(ori_ori_n1155_));
  INV        o1125(.A(ori_ori_n905_), .Y(ori_ori_n1156_));
  ZERO       o1126(.Y(ori02));
  ZERO       o1127(.Y(ori03));
  ZERO       o1128(.Y(ori05));
  NO2        m0000(.A(d), .B(c), .Y(mai_mai_n29_));
  AN2        m0001(.A(f), .B(e), .Y(mai_mai_n30_));
  NA3        m0002(.A(mai_mai_n30_), .B(mai_mai_n29_), .C(b), .Y(mai_mai_n31_));
  NOi32      m0003(.An(m), .Bn(l), .C(n), .Y(mai_mai_n32_));
  NOi32      m0004(.An(i), .Bn(m), .C(h), .Y(mai_mai_n33_));
  NA2        m0005(.A(mai_mai_n33_), .B(mai_mai_n32_), .Y(mai_mai_n34_));
  AN2        m0006(.A(m), .B(l), .Y(mai_mai_n35_));
  NOi32      m0007(.An(j), .Bn(m), .C(k), .Y(mai_mai_n36_));
  NA2        m0008(.A(mai_mai_n36_), .B(mai_mai_n35_), .Y(mai_mai_n37_));
  NO2        m0009(.A(mai_mai_n37_), .B(n), .Y(mai_mai_n38_));
  INV        m0010(.A(h), .Y(mai_mai_n39_));
  NAi21      m0011(.An(j), .B(l), .Y(mai_mai_n40_));
  NAi32      m0012(.An(n), .Bn(m), .C(m), .Y(mai_mai_n41_));
  NO3        m0013(.A(mai_mai_n41_), .B(mai_mai_n40_), .C(mai_mai_n39_), .Y(mai_mai_n42_));
  INV        m0014(.A(i), .Y(mai_mai_n43_));
  AN2        m0015(.A(h), .B(m), .Y(mai_mai_n44_));
  NA2        m0016(.A(mai_mai_n44_), .B(mai_mai_n43_), .Y(mai_mai_n45_));
  NAi21      m0017(.An(n), .B(m), .Y(mai_mai_n46_));
  NOi32      m0018(.An(k), .Bn(h), .C(l), .Y(mai_mai_n47_));
  NOi32      m0019(.An(k), .Bn(h), .C(m), .Y(mai_mai_n48_));
  INV        m0020(.A(mai_mai_n38_), .Y(mai_mai_n49_));
  NO2        m0021(.A(mai_mai_n49_), .B(mai_mai_n31_), .Y(mai_mai_n50_));
  INV        m0022(.A(c), .Y(mai_mai_n51_));
  NA2        m0023(.A(e), .B(b), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  INV        m0025(.A(d), .Y(mai_mai_n54_));
  NAi21      m0026(.An(i), .B(h), .Y(mai_mai_n55_));
  NAi31      m0027(.An(i), .B(l), .C(j), .Y(mai_mai_n56_));
  NA2        m0028(.A(m), .B(f), .Y(mai_mai_n57_));
  NAi21      m0029(.An(i), .B(j), .Y(mai_mai_n58_));
  NAi32      m0030(.An(n), .Bn(k), .C(m), .Y(mai_mai_n59_));
  NAi31      m0031(.An(l), .B(m), .C(k), .Y(mai_mai_n60_));
  NAi21      m0032(.An(e), .B(h), .Y(mai_mai_n61_));
  NAi41      m0033(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n62_));
  INV        m0034(.A(m), .Y(mai_mai_n63_));
  NA2        m0035(.A(k), .B(mai_mai_n63_), .Y(mai_mai_n64_));
  AN4        m0036(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n65_));
  NOi31      m0037(.An(h), .B(m), .C(f), .Y(mai_mai_n66_));
  NA2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi32      m0039(.An(m), .Bn(k), .C(j), .Y(mai_mai_n68_));
  NOi32      m0040(.An(h), .Bn(m), .C(f), .Y(mai_mai_n69_));
  NA2        m0041(.A(mai_mai_n69_), .B(mai_mai_n65_), .Y(mai_mai_n70_));
  OA220      m0042(.A0(mai_mai_n70_), .A1(mai_mai_n68_), .B0(mai_mai_n67_), .B1(mai_mai_n64_), .Y(mai_mai_n71_));
  INV        m0043(.A(mai_mai_n71_), .Y(mai_mai_n72_));
  INV        m0044(.A(n), .Y(mai_mai_n73_));
  NOi32      m0045(.An(e), .Bn(b), .C(d), .Y(mai_mai_n74_));
  NA2        m0046(.A(mai_mai_n74_), .B(mai_mai_n73_), .Y(mai_mai_n75_));
  INV        m0047(.A(j), .Y(mai_mai_n76_));
  AN3        m0048(.A(m), .B(k), .C(i), .Y(mai_mai_n77_));
  NA3        m0049(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(m), .Y(mai_mai_n78_));
  NAi32      m0050(.An(m), .Bn(f), .C(h), .Y(mai_mai_n79_));
  NAi31      m0051(.An(j), .B(m), .C(l), .Y(mai_mai_n80_));
  NA2        m0052(.A(m), .B(l), .Y(mai_mai_n81_));
  NAi31      m0053(.An(k), .B(j), .C(m), .Y(mai_mai_n82_));
  NO3        m0054(.A(mai_mai_n82_), .B(mai_mai_n81_), .C(f), .Y(mai_mai_n83_));
  AN2        m0055(.A(j), .B(m), .Y(mai_mai_n84_));
  NOi32      m0056(.An(m), .Bn(l), .C(i), .Y(mai_mai_n85_));
  NOi21      m0057(.An(m), .B(i), .Y(mai_mai_n86_));
  NOi32      m0058(.An(m), .Bn(j), .C(k), .Y(mai_mai_n87_));
  AOI220     m0059(.A0(mai_mai_n87_), .A1(mai_mai_n86_), .B0(mai_mai_n85_), .B1(mai_mai_n84_), .Y(mai_mai_n88_));
  NAi41      m0060(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n89_));
  AN2        m0061(.A(e), .B(b), .Y(mai_mai_n90_));
  NOi31      m0062(.An(c), .B(h), .C(f), .Y(mai_mai_n91_));
  NA2        m0063(.A(mai_mai_n91_), .B(mai_mai_n90_), .Y(mai_mai_n92_));
  NO2        m0064(.A(mai_mai_n92_), .B(mai_mai_n89_), .Y(mai_mai_n93_));
  NOi21      m0065(.An(i), .B(h), .Y(mai_mai_n94_));
  NA3        m0066(.A(mai_mai_n94_), .B(m), .C(mai_mai_n35_), .Y(mai_mai_n95_));
  INV        m0067(.A(a), .Y(mai_mai_n96_));
  NA2        m0068(.A(mai_mai_n90_), .B(mai_mai_n96_), .Y(mai_mai_n97_));
  INV        m0069(.A(l), .Y(mai_mai_n98_));
  NOi21      m0070(.An(m), .B(n), .Y(mai_mai_n99_));
  AN2        m0071(.A(k), .B(h), .Y(mai_mai_n100_));
  NO2        m0072(.A(mai_mai_n95_), .B(mai_mai_n75_), .Y(mai_mai_n101_));
  INV        m0073(.A(b), .Y(mai_mai_n102_));
  NA2        m0074(.A(l), .B(j), .Y(mai_mai_n103_));
  AN2        m0075(.A(k), .B(i), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NA2        m0077(.A(m), .B(e), .Y(mai_mai_n106_));
  NOi32      m0078(.An(c), .Bn(a), .C(d), .Y(mai_mai_n107_));
  NA2        m0079(.A(mai_mai_n107_), .B(mai_mai_n99_), .Y(mai_mai_n108_));
  NO2        m0080(.A(mai_mai_n101_), .B(mai_mai_n93_), .Y(mai_mai_n109_));
  OAI210     m0081(.A0(mai_mai_n88_), .A1(mai_mai_n75_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  NOi31      m0082(.An(k), .B(m), .C(j), .Y(mai_mai_n111_));
  NOi31      m0083(.An(k), .B(m), .C(i), .Y(mai_mai_n112_));
  NA3        m0084(.A(mai_mai_n112_), .B(mai_mai_n69_), .C(mai_mai_n65_), .Y(mai_mai_n113_));
  INV        m0085(.A(mai_mai_n113_), .Y(mai_mai_n114_));
  NOi32      m0086(.An(f), .Bn(b), .C(e), .Y(mai_mai_n115_));
  NAi21      m0087(.An(m), .B(h), .Y(mai_mai_n116_));
  NAi21      m0088(.An(m), .B(n), .Y(mai_mai_n117_));
  NAi21      m0089(.An(j), .B(k), .Y(mai_mai_n118_));
  NO3        m0090(.A(mai_mai_n118_), .B(mai_mai_n117_), .C(mai_mai_n116_), .Y(mai_mai_n119_));
  NAi41      m0091(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n120_));
  NAi31      m0092(.An(j), .B(k), .C(h), .Y(mai_mai_n121_));
  NO3        m0093(.A(mai_mai_n121_), .B(mai_mai_n120_), .C(mai_mai_n117_), .Y(mai_mai_n122_));
  AOI210     m0094(.A0(mai_mai_n119_), .A1(mai_mai_n115_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NO2        m0095(.A(k), .B(j), .Y(mai_mai_n124_));
  AN2        m0096(.A(k), .B(j), .Y(mai_mai_n125_));
  NAi21      m0097(.An(c), .B(b), .Y(mai_mai_n126_));
  NA2        m0098(.A(f), .B(d), .Y(mai_mai_n127_));
  NAi31      m0099(.An(f), .B(e), .C(b), .Y(mai_mai_n128_));
  NA2        m0100(.A(d), .B(b), .Y(mai_mai_n129_));
  NAi21      m0101(.An(e), .B(f), .Y(mai_mai_n130_));
  NA2        m0102(.A(b), .B(a), .Y(mai_mai_n131_));
  NAi21      m0103(.An(e), .B(m), .Y(mai_mai_n132_));
  NAi21      m0104(.An(c), .B(d), .Y(mai_mai_n133_));
  NAi31      m0105(.An(l), .B(k), .C(h), .Y(mai_mai_n134_));
  NAi21      m0106(.An(mai_mai_n114_), .B(mai_mai_n123_), .Y(mai_mai_n135_));
  NAi31      m0107(.An(e), .B(f), .C(b), .Y(mai_mai_n136_));
  NOi21      m0108(.An(m), .B(d), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n138_));
  NOi21      m0110(.An(h), .B(i), .Y(mai_mai_n139_));
  NOi21      m0111(.An(k), .B(m), .Y(mai_mai_n140_));
  NA3        m0112(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(n), .Y(mai_mai_n141_));
  NOi21      m0113(.An(h), .B(m), .Y(mai_mai_n142_));
  NO2        m0114(.A(mai_mai_n127_), .B(mai_mai_n126_), .Y(mai_mai_n143_));
  NA2        m0115(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NOi32      m0116(.An(n), .Bn(k), .C(m), .Y(mai_mai_n145_));
  NA2        m0117(.A(l), .B(i), .Y(mai_mai_n146_));
  NA2        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n147_), .B(mai_mai_n144_), .Y(mai_mai_n148_));
  NAi31      m0120(.An(d), .B(f), .C(c), .Y(mai_mai_n149_));
  NAi31      m0121(.An(e), .B(f), .C(c), .Y(mai_mai_n150_));
  NA2        m0122(.A(mai_mai_n150_), .B(mai_mai_n149_), .Y(mai_mai_n151_));
  NA2        m0123(.A(j), .B(h), .Y(mai_mai_n152_));
  OR3        m0124(.A(n), .B(m), .C(k), .Y(mai_mai_n153_));
  NO2        m0125(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NAi32      m0126(.An(m), .Bn(k), .C(n), .Y(mai_mai_n155_));
  NO2        m0127(.A(mai_mai_n155_), .B(mai_mai_n152_), .Y(mai_mai_n156_));
  AOI220     m0128(.A0(mai_mai_n156_), .A1(mai_mai_n138_), .B0(mai_mai_n154_), .B1(mai_mai_n151_), .Y(mai_mai_n157_));
  NO2        m0129(.A(n), .B(m), .Y(mai_mai_n158_));
  NA2        m0130(.A(mai_mai_n158_), .B(mai_mai_n47_), .Y(mai_mai_n159_));
  NAi21      m0131(.An(f), .B(e), .Y(mai_mai_n160_));
  NA2        m0132(.A(d), .B(c), .Y(mai_mai_n161_));
  NO2        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .Y(mai_mai_n162_));
  NOi21      m0134(.An(mai_mai_n162_), .B(mai_mai_n159_), .Y(mai_mai_n163_));
  NAi21      m0135(.An(d), .B(c), .Y(mai_mai_n164_));
  NAi31      m0136(.An(m), .B(n), .C(b), .Y(mai_mai_n165_));
  NA2        m0137(.A(k), .B(i), .Y(mai_mai_n166_));
  NAi21      m0138(.An(h), .B(f), .Y(mai_mai_n167_));
  NO2        m0139(.A(mai_mai_n167_), .B(mai_mai_n166_), .Y(mai_mai_n168_));
  NO2        m0140(.A(mai_mai_n165_), .B(mai_mai_n133_), .Y(mai_mai_n169_));
  NA2        m0141(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NOi32      m0142(.An(f), .Bn(c), .C(d), .Y(mai_mai_n171_));
  NOi32      m0143(.An(f), .Bn(c), .C(e), .Y(mai_mai_n172_));
  NO2        m0144(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  NO3        m0145(.A(n), .B(m), .C(j), .Y(mai_mai_n174_));
  NA2        m0146(.A(mai_mai_n174_), .B(mai_mai_n100_), .Y(mai_mai_n175_));
  AO210      m0147(.A0(mai_mai_n175_), .A1(mai_mai_n159_), .B0(mai_mai_n173_), .Y(mai_mai_n176_));
  NAi41      m0148(.An(mai_mai_n163_), .B(mai_mai_n176_), .C(mai_mai_n170_), .D(mai_mai_n157_), .Y(mai_mai_n177_));
  OR3        m0149(.A(mai_mai_n177_), .B(mai_mai_n148_), .C(mai_mai_n135_), .Y(mai_mai_n178_));
  NO4        m0150(.A(mai_mai_n178_), .B(mai_mai_n110_), .C(mai_mai_n72_), .D(mai_mai_n50_), .Y(mai_mai_n179_));
  NA3        m0151(.A(m), .B(mai_mai_n98_), .C(j), .Y(mai_mai_n180_));
  NAi31      m0152(.An(n), .B(h), .C(m), .Y(mai_mai_n181_));
  NO2        m0153(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NOi32      m0154(.An(m), .Bn(k), .C(l), .Y(mai_mai_n183_));
  NA3        m0155(.A(mai_mai_n183_), .B(mai_mai_n76_), .C(m), .Y(mai_mai_n184_));
  AN2        m0156(.A(i), .B(m), .Y(mai_mai_n185_));
  NA3        m0157(.A(k), .B(mai_mai_n185_), .C(mai_mai_n99_), .Y(mai_mai_n186_));
  NAi41      m0158(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n187_));
  INV        m0159(.A(f), .Y(mai_mai_n188_));
  INV        m0160(.A(m), .Y(mai_mai_n189_));
  NOi31      m0161(.An(i), .B(j), .C(h), .Y(mai_mai_n190_));
  NOi21      m0162(.An(l), .B(m), .Y(mai_mai_n191_));
  NA2        m0163(.A(mai_mai_n191_), .B(mai_mai_n190_), .Y(mai_mai_n192_));
  NO3        m0164(.A(mai_mai_n192_), .B(mai_mai_n189_), .C(mai_mai_n188_), .Y(mai_mai_n193_));
  NOi21      m0165(.An(n), .B(m), .Y(mai_mai_n194_));
  NOi32      m0166(.An(l), .Bn(i), .C(j), .Y(mai_mai_n195_));
  NA2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  OA220      m0168(.A0(mai_mai_n196_), .A1(mai_mai_n92_), .B0(mai_mai_n68_), .B1(mai_mai_n67_), .Y(mai_mai_n197_));
  NAi21      m0169(.An(j), .B(h), .Y(mai_mai_n198_));
  XN2        m0170(.A(i), .B(h), .Y(mai_mai_n199_));
  NA2        m0171(.A(mai_mai_n199_), .B(mai_mai_n198_), .Y(mai_mai_n200_));
  NOi31      m0172(.An(k), .B(n), .C(m), .Y(mai_mai_n201_));
  NOi31      m0173(.An(mai_mai_n201_), .B(mai_mai_n161_), .C(mai_mai_n160_), .Y(mai_mai_n202_));
  NA2        m0174(.A(mai_mai_n202_), .B(mai_mai_n200_), .Y(mai_mai_n203_));
  NAi31      m0175(.An(f), .B(e), .C(c), .Y(mai_mai_n204_));
  NO4        m0176(.A(mai_mai_n204_), .B(mai_mai_n153_), .C(mai_mai_n152_), .D(mai_mai_n54_), .Y(mai_mai_n205_));
  NA4        m0177(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n206_));
  NAi32      m0178(.An(m), .Bn(i), .C(k), .Y(mai_mai_n207_));
  INV        m0179(.A(k), .Y(mai_mai_n208_));
  INV        m0180(.A(mai_mai_n205_), .Y(mai_mai_n209_));
  NAi21      m0181(.An(n), .B(a), .Y(mai_mai_n210_));
  NO2        m0182(.A(mai_mai_n210_), .B(mai_mai_n129_), .Y(mai_mai_n211_));
  NAi41      m0183(.An(m), .B(m), .C(k), .D(h), .Y(mai_mai_n212_));
  AN3        m0184(.A(mai_mai_n209_), .B(mai_mai_n203_), .C(mai_mai_n197_), .Y(mai_mai_n213_));
  OR2        m0185(.A(h), .B(m), .Y(mai_mai_n214_));
  NO2        m0186(.A(mai_mai_n214_), .B(mai_mai_n89_), .Y(mai_mai_n215_));
  NA2        m0187(.A(mai_mai_n215_), .B(mai_mai_n115_), .Y(mai_mai_n216_));
  NAi31      m0188(.An(e), .B(d), .C(b), .Y(mai_mai_n217_));
  NA2        m0189(.A(mai_mai_n140_), .B(mai_mai_n94_), .Y(mai_mai_n218_));
  NO2        m0190(.A(n), .B(a), .Y(mai_mai_n219_));
  NAi31      m0191(.An(mai_mai_n212_), .B(mai_mai_n219_), .C(mai_mai_n90_), .Y(mai_mai_n220_));
  NAi21      m0192(.An(h), .B(i), .Y(mai_mai_n221_));
  NA2        m0193(.A(mai_mai_n158_), .B(k), .Y(mai_mai_n222_));
  NO2        m0194(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n223_));
  NA2        m0195(.A(mai_mai_n223_), .B(mai_mai_n171_), .Y(mai_mai_n224_));
  NA3        m0196(.A(mai_mai_n224_), .B(mai_mai_n220_), .C(mai_mai_n216_), .Y(mai_mai_n225_));
  NOi21      m0197(.An(m), .B(e), .Y(mai_mai_n226_));
  NO2        m0198(.A(mai_mai_n62_), .B(mai_mai_n63_), .Y(mai_mai_n227_));
  AOI210     m0199(.A0(k), .A1(mai_mai_n76_), .B0(j), .Y(mai_mai_n228_));
  NAi21      m0200(.An(f), .B(m), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n59_), .B(mai_mai_n103_), .Y(mai_mai_n230_));
  NOi21      m0202(.An(mai_mai_n213_), .B(mai_mai_n225_), .Y(mai_mai_n231_));
  NO3        m0203(.A(mai_mai_n182_), .B(mai_mai_n42_), .C(mai_mai_n38_), .Y(mai_mai_n232_));
  NO2        m0204(.A(mai_mai_n232_), .B(mai_mai_n97_), .Y(mai_mai_n233_));
  NA3        m0205(.A(mai_mai_n54_), .B(c), .C(b), .Y(mai_mai_n234_));
  NAi21      m0206(.An(h), .B(m), .Y(mai_mai_n235_));
  OR4        m0207(.A(mai_mai_n235_), .B(mai_mai_n234_), .C(mai_mai_n196_), .D(e), .Y(mai_mai_n236_));
  NO2        m0208(.A(mai_mai_n218_), .B(mai_mai_n229_), .Y(mai_mai_n237_));
  NAi31      m0209(.An(m), .B(k), .C(h), .Y(mai_mai_n238_));
  NO3        m0210(.A(mai_mai_n117_), .B(mai_mai_n238_), .C(l), .Y(mai_mai_n239_));
  NAi31      m0211(.An(e), .B(d), .C(a), .Y(mai_mai_n240_));
  NA2        m0212(.A(mai_mai_n239_), .B(mai_mai_n115_), .Y(mai_mai_n241_));
  NA2        m0213(.A(mai_mai_n241_), .B(mai_mai_n236_), .Y(mai_mai_n242_));
  NA4        m0214(.A(mai_mai_n140_), .B(mai_mai_n69_), .C(mai_mai_n65_), .D(mai_mai_n103_), .Y(mai_mai_n243_));
  NA3        m0215(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n73_), .Y(mai_mai_n244_));
  NO2        m0216(.A(mai_mai_n244_), .B(mai_mai_n173_), .Y(mai_mai_n245_));
  NOi21      m0217(.An(mai_mai_n243_), .B(mai_mai_n245_), .Y(mai_mai_n246_));
  NA3        m0218(.A(e), .B(c), .C(b), .Y(mai_mai_n247_));
  NAi21      m0219(.An(l), .B(k), .Y(mai_mai_n248_));
  NO2        m0220(.A(mai_mai_n248_), .B(mai_mai_n46_), .Y(mai_mai_n249_));
  NOi21      m0221(.An(l), .B(j), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n142_), .B(mai_mai_n250_), .Y(mai_mai_n251_));
  OR3        m0223(.A(mai_mai_n62_), .B(mai_mai_n63_), .C(e), .Y(mai_mai_n252_));
  AOI210     m0224(.A0(mai_mai_n1410_), .A1(mai_mai_n251_), .B0(mai_mai_n252_), .Y(mai_mai_n253_));
  INV        m0225(.A(mai_mai_n253_), .Y(mai_mai_n254_));
  NAi32      m0226(.An(j), .Bn(h), .C(i), .Y(mai_mai_n255_));
  NAi21      m0227(.An(m), .B(l), .Y(mai_mai_n256_));
  NO3        m0228(.A(mai_mai_n256_), .B(mai_mai_n255_), .C(mai_mai_n73_), .Y(mai_mai_n257_));
  NA2        m0229(.A(h), .B(m), .Y(mai_mai_n258_));
  NA2        m0230(.A(mai_mai_n145_), .B(mai_mai_n43_), .Y(mai_mai_n259_));
  NO2        m0231(.A(mai_mai_n259_), .B(mai_mai_n258_), .Y(mai_mai_n260_));
  NA2        m0232(.A(mai_mai_n257_), .B(mai_mai_n143_), .Y(mai_mai_n261_));
  NA3        m0233(.A(mai_mai_n261_), .B(mai_mai_n254_), .C(mai_mai_n246_), .Y(mai_mai_n262_));
  NO2        m0234(.A(mai_mai_n92_), .B(mai_mai_n89_), .Y(mai_mai_n263_));
  NAi32      m0235(.An(n), .Bn(m), .C(l), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n264_), .B(mai_mai_n255_), .Y(mai_mai_n265_));
  NA2        m0237(.A(mai_mai_n265_), .B(mai_mai_n162_), .Y(mai_mai_n266_));
  NO2        m0238(.A(mai_mai_n108_), .B(mai_mai_n102_), .Y(mai_mai_n267_));
  NAi31      m0239(.An(k), .B(l), .C(j), .Y(mai_mai_n268_));
  NA2        m0240(.A(mai_mai_n248_), .B(mai_mai_n268_), .Y(mai_mai_n269_));
  NOi21      m0241(.An(mai_mai_n269_), .B(mai_mai_n106_), .Y(mai_mai_n270_));
  NA2        m0242(.A(mai_mai_n270_), .B(mai_mai_n267_), .Y(mai_mai_n271_));
  NA2        m0243(.A(mai_mai_n271_), .B(mai_mai_n266_), .Y(mai_mai_n272_));
  NO4        m0244(.A(mai_mai_n272_), .B(mai_mai_n262_), .C(mai_mai_n242_), .D(mai_mai_n233_), .Y(mai_mai_n273_));
  NA2        m0245(.A(mai_mai_n223_), .B(mai_mai_n172_), .Y(mai_mai_n274_));
  NAi21      m0246(.An(m), .B(k), .Y(mai_mai_n275_));
  NAi41      m0247(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n276_));
  NA2        m0248(.A(e), .B(c), .Y(mai_mai_n277_));
  NO3        m0249(.A(mai_mai_n277_), .B(n), .C(d), .Y(mai_mai_n278_));
  NA2        m0250(.A(f), .B(mai_mai_n104_), .Y(mai_mai_n279_));
  NO2        m0251(.A(mai_mai_n279_), .B(mai_mai_n189_), .Y(mai_mai_n280_));
  NAi31      m0252(.An(d), .B(e), .C(b), .Y(mai_mai_n281_));
  NO2        m0253(.A(mai_mai_n117_), .B(mai_mai_n281_), .Y(mai_mai_n282_));
  NA2        m0254(.A(mai_mai_n282_), .B(mai_mai_n280_), .Y(mai_mai_n283_));
  NA2        m0255(.A(mai_mai_n283_), .B(mai_mai_n274_), .Y(mai_mai_n284_));
  NO4        m0256(.A(mai_mai_n276_), .B(mai_mai_n68_), .C(mai_mai_n61_), .D(mai_mai_n189_), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n219_), .B(mai_mai_n90_), .Y(mai_mai_n286_));
  OR2        m0258(.A(mai_mai_n286_), .B(mai_mai_n184_), .Y(mai_mai_n287_));
  NOi31      m0259(.An(l), .B(n), .C(m), .Y(mai_mai_n288_));
  NA2        m0260(.A(mai_mai_n288_), .B(mai_mai_n190_), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n289_), .B(mai_mai_n173_), .Y(mai_mai_n290_));
  NAi32      m0262(.An(mai_mai_n290_), .Bn(mai_mai_n285_), .C(mai_mai_n287_), .Y(mai_mai_n291_));
  NAi32      m0263(.An(m), .Bn(j), .C(k), .Y(mai_mai_n292_));
  NAi41      m0264(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n293_));
  NA2        m0265(.A(mai_mai_n187_), .B(mai_mai_n293_), .Y(mai_mai_n294_));
  NOi31      m0266(.An(j), .B(m), .C(k), .Y(mai_mai_n295_));
  NO2        m0267(.A(mai_mai_n111_), .B(mai_mai_n295_), .Y(mai_mai_n296_));
  AN3        m0268(.A(h), .B(m), .C(f), .Y(mai_mai_n297_));
  NAi31      m0269(.An(mai_mai_n296_), .B(mai_mai_n297_), .C(mai_mai_n294_), .Y(mai_mai_n298_));
  NOi32      m0270(.An(m), .Bn(j), .C(l), .Y(mai_mai_n299_));
  NO2        m0271(.A(mai_mai_n299_), .B(mai_mai_n85_), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n256_), .B(mai_mai_n255_), .Y(mai_mai_n301_));
  NO2        m0273(.A(mai_mai_n192_), .B(m), .Y(mai_mai_n302_));
  INV        m0274(.A(mai_mai_n298_), .Y(mai_mai_n303_));
  NA3        m0275(.A(h), .B(m), .C(f), .Y(mai_mai_n304_));
  NO2        m0276(.A(mai_mai_n304_), .B(mai_mai_n64_), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n293_), .B(mai_mai_n187_), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n142_), .B(e), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n307_), .B(mai_mai_n40_), .Y(mai_mai_n308_));
  AOI220     m0280(.A0(mai_mai_n308_), .A1(mai_mai_n267_), .B0(mai_mai_n306_), .B1(mai_mai_n305_), .Y(mai_mai_n309_));
  NOi32      m0281(.An(j), .Bn(m), .C(i), .Y(mai_mai_n310_));
  NA3        m0282(.A(mai_mai_n310_), .B(mai_mai_n248_), .C(mai_mai_n99_), .Y(mai_mai_n311_));
  NOi32      m0283(.An(e), .Bn(b), .C(a), .Y(mai_mai_n312_));
  INV        m0284(.A(mai_mai_n275_), .Y(mai_mai_n313_));
  NO3        m0285(.A(mai_mai_n276_), .B(mai_mai_n61_), .C(mai_mai_n189_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n186_), .B(mai_mai_n34_), .Y(mai_mai_n315_));
  AOI220     m0287(.A0(mai_mai_n315_), .A1(mai_mai_n312_), .B0(mai_mai_n314_), .B1(mai_mai_n313_), .Y(mai_mai_n316_));
  NO2        m0288(.A(mai_mai_n281_), .B(n), .Y(mai_mai_n317_));
  NA2        m0289(.A(mai_mai_n185_), .B(k), .Y(mai_mai_n318_));
  NA3        m0290(.A(m), .B(mai_mai_n98_), .C(mai_mai_n188_), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n320_));
  NAi41      m0292(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n48_), .B(mai_mai_n99_), .Y(mai_mai_n322_));
  NO2        m0294(.A(mai_mai_n322_), .B(mai_mai_n321_), .Y(mai_mai_n323_));
  AOI220     m0295(.A0(mai_mai_n323_), .A1(b), .B0(mai_mai_n320_), .B1(mai_mai_n317_), .Y(mai_mai_n324_));
  NA3        m0296(.A(mai_mai_n324_), .B(mai_mai_n316_), .C(mai_mai_n309_), .Y(mai_mai_n325_));
  NO4        m0297(.A(mai_mai_n325_), .B(mai_mai_n303_), .C(mai_mai_n291_), .D(mai_mai_n284_), .Y(mai_mai_n326_));
  NA4        m0298(.A(mai_mai_n326_), .B(mai_mai_n273_), .C(mai_mai_n231_), .D(mai_mai_n179_), .Y(mai10));
  NA3        m0299(.A(m), .B(k), .C(i), .Y(mai_mai_n328_));
  NO3        m0300(.A(mai_mai_n328_), .B(j), .C(mai_mai_n189_), .Y(mai_mai_n329_));
  NOi21      m0301(.An(e), .B(f), .Y(mai_mai_n330_));
  NO4        m0302(.A(mai_mai_n133_), .B(mai_mai_n330_), .C(n), .D(mai_mai_n96_), .Y(mai_mai_n331_));
  NAi31      m0303(.An(b), .B(f), .C(c), .Y(mai_mai_n332_));
  INV        m0304(.A(mai_mai_n332_), .Y(mai_mai_n333_));
  NOi32      m0305(.An(k), .Bn(h), .C(j), .Y(mai_mai_n334_));
  NA2        m0306(.A(mai_mai_n334_), .B(mai_mai_n194_), .Y(mai_mai_n335_));
  NA2        m0307(.A(mai_mai_n141_), .B(mai_mai_n335_), .Y(mai_mai_n336_));
  AOI220     m0308(.A0(mai_mai_n336_), .A1(mai_mai_n333_), .B0(mai_mai_n331_), .B1(mai_mai_n329_), .Y(mai_mai_n337_));
  AN2        m0309(.A(j), .B(h), .Y(mai_mai_n338_));
  NO3        m0310(.A(n), .B(m), .C(k), .Y(mai_mai_n339_));
  NA2        m0311(.A(mai_mai_n339_), .B(mai_mai_n338_), .Y(mai_mai_n340_));
  NO3        m0312(.A(mai_mai_n340_), .B(mai_mai_n133_), .C(mai_mai_n188_), .Y(mai_mai_n341_));
  OR2        m0313(.A(m), .B(k), .Y(mai_mai_n342_));
  NO2        m0314(.A(mai_mai_n152_), .B(mai_mai_n342_), .Y(mai_mai_n343_));
  NA4        m0315(.A(n), .B(f), .C(c), .D(mai_mai_n102_), .Y(mai_mai_n344_));
  NOi21      m0316(.An(mai_mai_n343_), .B(mai_mai_n344_), .Y(mai_mai_n345_));
  NOi32      m0317(.An(d), .Bn(a), .C(c), .Y(mai_mai_n346_));
  NA2        m0318(.A(mai_mai_n346_), .B(mai_mai_n160_), .Y(mai_mai_n347_));
  NAi21      m0319(.An(i), .B(m), .Y(mai_mai_n348_));
  NAi31      m0320(.An(k), .B(m), .C(j), .Y(mai_mai_n349_));
  NO2        m0321(.A(mai_mai_n345_), .B(mai_mai_n341_), .Y(mai_mai_n350_));
  NO2        m0322(.A(mai_mai_n344_), .B(mai_mai_n256_), .Y(mai_mai_n351_));
  NOi32      m0323(.An(f), .Bn(d), .C(c), .Y(mai_mai_n352_));
  AOI220     m0324(.A0(mai_mai_n352_), .A1(mai_mai_n265_), .B0(mai_mai_n351_), .B1(mai_mai_n190_), .Y(mai_mai_n353_));
  NA3        m0325(.A(mai_mai_n353_), .B(mai_mai_n350_), .C(mai_mai_n337_), .Y(mai_mai_n354_));
  NO2        m0326(.A(mai_mai_n54_), .B(mai_mai_n102_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n219_), .B(mai_mai_n355_), .Y(mai_mai_n356_));
  INV        m0328(.A(e), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n44_), .B(e), .Y(mai_mai_n358_));
  OAI220     m0330(.A0(mai_mai_n358_), .A1(mai_mai_n180_), .B0(mai_mai_n184_), .B1(mai_mai_n357_), .Y(mai_mai_n359_));
  AN2        m0331(.A(m), .B(e), .Y(mai_mai_n360_));
  NA3        m0332(.A(mai_mai_n360_), .B(mai_mai_n183_), .C(i), .Y(mai_mai_n361_));
  INV        m0333(.A(mai_mai_n361_), .Y(mai_mai_n362_));
  NO2        m0334(.A(mai_mai_n88_), .B(mai_mai_n357_), .Y(mai_mai_n363_));
  NO3        m0335(.A(mai_mai_n363_), .B(mai_mai_n362_), .C(mai_mai_n359_), .Y(mai_mai_n364_));
  NOi32      m0336(.An(h), .Bn(e), .C(m), .Y(mai_mai_n365_));
  NA3        m0337(.A(mai_mai_n365_), .B(mai_mai_n250_), .C(m), .Y(mai_mai_n366_));
  NOi21      m0338(.An(m), .B(h), .Y(mai_mai_n367_));
  AN3        m0339(.A(m), .B(l), .C(i), .Y(mai_mai_n368_));
  NA3        m0340(.A(mai_mai_n368_), .B(mai_mai_n367_), .C(e), .Y(mai_mai_n369_));
  AN3        m0341(.A(h), .B(m), .C(e), .Y(mai_mai_n370_));
  NA2        m0342(.A(mai_mai_n370_), .B(mai_mai_n85_), .Y(mai_mai_n371_));
  AN3        m0343(.A(mai_mai_n371_), .B(mai_mai_n369_), .C(mai_mai_n366_), .Y(mai_mai_n372_));
  AOI210     m0344(.A0(mai_mai_n372_), .A1(mai_mai_n364_), .B0(mai_mai_n356_), .Y(mai_mai_n373_));
  NA3        m0345(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(e), .Y(mai_mai_n374_));
  NO2        m0346(.A(mai_mai_n374_), .B(mai_mai_n356_), .Y(mai_mai_n375_));
  NA3        m0347(.A(mai_mai_n346_), .B(mai_mai_n160_), .C(mai_mai_n73_), .Y(mai_mai_n376_));
  NAi31      m0348(.An(b), .B(c), .C(a), .Y(mai_mai_n377_));
  NO2        m0349(.A(mai_mai_n377_), .B(n), .Y(mai_mai_n378_));
  OAI210     m0350(.A0(mai_mai_n48_), .A1(mai_mai_n47_), .B0(m), .Y(mai_mai_n379_));
  NO2        m0351(.A(mai_mai_n379_), .B(mai_mai_n130_), .Y(mai_mai_n380_));
  NA2        m0352(.A(mai_mai_n380_), .B(mai_mai_n378_), .Y(mai_mai_n381_));
  INV        m0353(.A(mai_mai_n381_), .Y(mai_mai_n382_));
  NO4        m0354(.A(mai_mai_n382_), .B(mai_mai_n375_), .C(mai_mai_n373_), .D(mai_mai_n354_), .Y(mai_mai_n383_));
  NA2        m0355(.A(i), .B(m), .Y(mai_mai_n384_));
  NO3        m0356(.A(mai_mai_n240_), .B(mai_mai_n384_), .C(c), .Y(mai_mai_n385_));
  NOi21      m0357(.An(a), .B(n), .Y(mai_mai_n386_));
  NOi21      m0358(.An(d), .B(c), .Y(mai_mai_n387_));
  NA2        m0359(.A(mai_mai_n387_), .B(mai_mai_n386_), .Y(mai_mai_n388_));
  NA3        m0360(.A(i), .B(m), .C(f), .Y(mai_mai_n389_));
  OR2        m0361(.A(mai_mai_n389_), .B(mai_mai_n60_), .Y(mai_mai_n390_));
  NA3        m0362(.A(mai_mai_n368_), .B(mai_mai_n367_), .C(mai_mai_n160_), .Y(mai_mai_n391_));
  AOI210     m0363(.A0(mai_mai_n391_), .A1(mai_mai_n390_), .B0(mai_mai_n388_), .Y(mai_mai_n392_));
  AOI210     m0364(.A0(mai_mai_n385_), .A1(mai_mai_n249_), .B0(mai_mai_n392_), .Y(mai_mai_n393_));
  OR2        m0365(.A(n), .B(m), .Y(mai_mai_n394_));
  NO2        m0366(.A(mai_mai_n394_), .B(mai_mai_n134_), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n161_), .B(mai_mai_n130_), .Y(mai_mai_n396_));
  OAI210     m0368(.A0(mai_mai_n395_), .A1(mai_mai_n154_), .B0(mai_mai_n396_), .Y(mai_mai_n397_));
  INV        m0369(.A(mai_mai_n322_), .Y(mai_mai_n398_));
  NA3        m0370(.A(mai_mai_n398_), .B(mai_mai_n312_), .C(d), .Y(mai_mai_n399_));
  NO2        m0371(.A(mai_mai_n377_), .B(mai_mai_n46_), .Y(mai_mai_n400_));
  NAi21      m0372(.An(k), .B(j), .Y(mai_mai_n401_));
  NAi21      m0373(.An(e), .B(d), .Y(mai_mai_n402_));
  INV        m0374(.A(mai_mai_n402_), .Y(mai_mai_n403_));
  NO2        m0375(.A(mai_mai_n222_), .B(mai_mai_n188_), .Y(mai_mai_n404_));
  NA3        m0376(.A(mai_mai_n404_), .B(mai_mai_n403_), .C(mai_mai_n200_), .Y(mai_mai_n405_));
  NA3        m0377(.A(mai_mai_n405_), .B(mai_mai_n399_), .C(mai_mai_n397_), .Y(mai_mai_n406_));
  NO2        m0378(.A(mai_mai_n289_), .B(mai_mai_n188_), .Y(mai_mai_n407_));
  NA2        m0379(.A(mai_mai_n407_), .B(mai_mai_n403_), .Y(mai_mai_n408_));
  NOi31      m0380(.An(n), .B(m), .C(k), .Y(mai_mai_n409_));
  AOI220     m0381(.A0(mai_mai_n409_), .A1(mai_mai_n338_), .B0(mai_mai_n194_), .B1(mai_mai_n47_), .Y(mai_mai_n410_));
  NAi31      m0382(.An(m), .B(f), .C(c), .Y(mai_mai_n411_));
  OR3        m0383(.A(mai_mai_n411_), .B(mai_mai_n410_), .C(e), .Y(mai_mai_n412_));
  NA3        m0384(.A(mai_mai_n412_), .B(mai_mai_n408_), .C(mai_mai_n266_), .Y(mai_mai_n413_));
  NOi31      m0385(.An(mai_mai_n393_), .B(mai_mai_n413_), .C(mai_mai_n406_), .Y(mai_mai_n414_));
  NOi32      m0386(.An(c), .Bn(a), .C(b), .Y(mai_mai_n415_));
  NA2        m0387(.A(mai_mai_n415_), .B(mai_mai_n99_), .Y(mai_mai_n416_));
  INV        m0388(.A(mai_mai_n238_), .Y(mai_mai_n417_));
  AN2        m0389(.A(e), .B(d), .Y(mai_mai_n418_));
  NA2        m0390(.A(mai_mai_n418_), .B(mai_mai_n417_), .Y(mai_mai_n419_));
  INV        m0391(.A(mai_mai_n130_), .Y(mai_mai_n420_));
  NO2        m0392(.A(mai_mai_n116_), .B(mai_mai_n40_), .Y(mai_mai_n421_));
  NO2        m0393(.A(mai_mai_n57_), .B(e), .Y(mai_mai_n422_));
  NA2        m0394(.A(i), .B(mai_mai_n105_), .Y(mai_mai_n423_));
  AOI220     m0395(.A0(mai_mai_n423_), .A1(mai_mai_n422_), .B0(mai_mai_n421_), .B1(mai_mai_n420_), .Y(mai_mai_n424_));
  AOI210     m0396(.A0(mai_mai_n424_), .A1(mai_mai_n419_), .B0(mai_mai_n416_), .Y(mai_mai_n425_));
  NOi21      m0397(.An(a), .B(b), .Y(mai_mai_n426_));
  NA3        m0398(.A(e), .B(d), .C(c), .Y(mai_mai_n427_));
  NAi21      m0399(.An(mai_mai_n427_), .B(mai_mai_n426_), .Y(mai_mai_n428_));
  NO2        m0400(.A(mai_mai_n376_), .B(mai_mai_n184_), .Y(mai_mai_n429_));
  NO4        m0401(.A(mai_mai_n167_), .B(mai_mai_n89_), .C(mai_mai_n51_), .D(b), .Y(mai_mai_n430_));
  OR2        m0402(.A(k), .B(j), .Y(mai_mai_n431_));
  NA2        m0403(.A(l), .B(k), .Y(mai_mai_n432_));
  AOI210     m0404(.A0(mai_mai_n207_), .A1(mai_mai_n292_), .B0(mai_mai_n73_), .Y(mai_mai_n433_));
  NA2        m0405(.A(mai_mai_n243_), .B(mai_mai_n113_), .Y(mai_mai_n434_));
  NA2        m0406(.A(mai_mai_n346_), .B(mai_mai_n99_), .Y(mai_mai_n435_));
  NO4        m0407(.A(mai_mai_n435_), .B(mai_mai_n82_), .C(mai_mai_n98_), .D(e), .Y(mai_mai_n436_));
  NO2        m0408(.A(mai_mai_n436_), .B(mai_mai_n434_), .Y(mai_mai_n437_));
  INV        m0409(.A(mai_mai_n437_), .Y(mai_mai_n438_));
  NO4        m0410(.A(mai_mai_n438_), .B(mai_mai_n430_), .C(mai_mai_n429_), .D(mai_mai_n425_), .Y(mai_mai_n439_));
  NOi21      m0411(.An(d), .B(e), .Y(mai_mai_n440_));
  NAi31      m0412(.An(j), .B(l), .C(i), .Y(mai_mai_n441_));
  OAI210     m0413(.A0(mai_mai_n441_), .A1(mai_mai_n117_), .B0(mai_mai_n89_), .Y(mai_mai_n442_));
  NO3        m0414(.A(mai_mai_n347_), .B(mai_mai_n300_), .C(mai_mai_n181_), .Y(mai_mai_n443_));
  NO2        m0415(.A(mai_mai_n347_), .B(mai_mai_n322_), .Y(mai_mai_n444_));
  NO4        m0416(.A(mai_mai_n444_), .B(mai_mai_n443_), .C(mai_mai_n163_), .D(mai_mai_n263_), .Y(mai_mai_n445_));
  NA2        m0417(.A(mai_mai_n445_), .B(mai_mai_n213_), .Y(mai_mai_n446_));
  OAI210     m0418(.A0(mai_mai_n112_), .A1(mai_mai_n111_), .B0(n), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n447_), .B(mai_mai_n116_), .Y(mai_mai_n448_));
  OA210      m0420(.A0(mai_mai_n215_), .A1(mai_mai_n448_), .B0(mai_mai_n172_), .Y(mai_mai_n449_));
  XO2        m0421(.A(i), .B(h), .Y(mai_mai_n450_));
  NA3        m0422(.A(mai_mai_n450_), .B(mai_mai_n140_), .C(n), .Y(mai_mai_n451_));
  NAi41      m0423(.An(mai_mai_n257_), .B(mai_mai_n451_), .C(mai_mai_n410_), .D(mai_mai_n335_), .Y(mai_mai_n452_));
  NOi32      m0424(.An(mai_mai_n452_), .Bn(mai_mai_n422_), .C(mai_mai_n234_), .Y(mai_mai_n453_));
  NAi31      m0425(.An(c), .B(f), .C(d), .Y(mai_mai_n454_));
  AOI210     m0426(.A0(mai_mai_n244_), .A1(mai_mai_n175_), .B0(mai_mai_n454_), .Y(mai_mai_n455_));
  NOi21      m0427(.An(mai_mai_n71_), .B(mai_mai_n455_), .Y(mai_mai_n456_));
  NA3        m0428(.A(mai_mai_n331_), .B(mai_mai_n85_), .C(mai_mai_n84_), .Y(mai_mai_n457_));
  NA2        m0429(.A(mai_mai_n201_), .B(mai_mai_n94_), .Y(mai_mai_n458_));
  AOI210     m0430(.A0(mai_mai_n458_), .A1(mai_mai_n159_), .B0(mai_mai_n454_), .Y(mai_mai_n459_));
  AOI210     m0431(.A0(mai_mai_n311_), .A1(mai_mai_n34_), .B0(mai_mai_n428_), .Y(mai_mai_n460_));
  NOi31      m0432(.An(mai_mai_n457_), .B(mai_mai_n460_), .C(mai_mai_n459_), .Y(mai_mai_n461_));
  NA3        m0433(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(f), .Y(mai_mai_n462_));
  NO2        m0434(.A(mai_mai_n462_), .B(mai_mai_n388_), .Y(mai_mai_n463_));
  NO2        m0435(.A(mai_mai_n463_), .B(mai_mai_n253_), .Y(mai_mai_n464_));
  NA3        m0436(.A(mai_mai_n464_), .B(mai_mai_n461_), .C(mai_mai_n456_), .Y(mai_mai_n465_));
  NO4        m0437(.A(mai_mai_n465_), .B(mai_mai_n453_), .C(mai_mai_n449_), .D(mai_mai_n446_), .Y(mai_mai_n466_));
  NA4        m0438(.A(mai_mai_n466_), .B(mai_mai_n439_), .C(mai_mai_n414_), .D(mai_mai_n383_), .Y(mai11));
  NO2        m0439(.A(mai_mai_n62_), .B(f), .Y(mai_mai_n468_));
  NA2        m0440(.A(j), .B(m), .Y(mai_mai_n469_));
  NAi31      m0441(.An(i), .B(m), .C(l), .Y(mai_mai_n470_));
  NA3        m0442(.A(m), .B(k), .C(j), .Y(mai_mai_n471_));
  NOi32      m0443(.An(e), .Bn(b), .C(f), .Y(mai_mai_n472_));
  NA2        m0444(.A(j), .B(mai_mai_n99_), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n44_), .B(j), .Y(mai_mai_n474_));
  NO2        m0446(.A(mai_mai_n474_), .B(mai_mai_n259_), .Y(mai_mai_n475_));
  NAi31      m0447(.An(d), .B(e), .C(a), .Y(mai_mai_n476_));
  NO2        m0448(.A(mai_mai_n476_), .B(n), .Y(mai_mai_n477_));
  NA2        m0449(.A(mai_mai_n475_), .B(mai_mai_n472_), .Y(mai_mai_n478_));
  NAi41      m0450(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n479_));
  AN2        m0451(.A(mai_mai_n479_), .B(mai_mai_n321_), .Y(mai_mai_n480_));
  AOI210     m0452(.A0(mai_mai_n480_), .A1(mai_mai_n347_), .B0(mai_mai_n235_), .Y(mai_mai_n481_));
  NA2        m0453(.A(j), .B(i), .Y(mai_mai_n482_));
  NAi31      m0454(.An(n), .B(m), .C(k), .Y(mai_mai_n483_));
  NO3        m0455(.A(mai_mai_n483_), .B(mai_mai_n482_), .C(mai_mai_n98_), .Y(mai_mai_n484_));
  NO4        m0456(.A(n), .B(d), .C(mai_mai_n102_), .D(a), .Y(mai_mai_n485_));
  OR2        m0457(.A(n), .B(c), .Y(mai_mai_n486_));
  NOi32      m0458(.An(m), .Bn(f), .C(i), .Y(mai_mai_n487_));
  NO2        m0459(.A(mai_mai_n238_), .B(mai_mai_n46_), .Y(mai_mai_n488_));
  NA2        m0460(.A(mai_mai_n125_), .B(mai_mai_n33_), .Y(mai_mai_n489_));
  OAI220     m0461(.A0(mai_mai_n489_), .A1(m), .B0(mai_mai_n474_), .B1(mai_mai_n207_), .Y(mai_mai_n490_));
  NOi41      m0462(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n491_));
  NAi32      m0463(.An(e), .Bn(b), .C(c), .Y(mai_mai_n492_));
  OR2        m0464(.A(mai_mai_n492_), .B(mai_mai_n73_), .Y(mai_mai_n493_));
  AN2        m0465(.A(mai_mai_n293_), .B(mai_mai_n276_), .Y(mai_mai_n494_));
  NA2        m0466(.A(mai_mai_n494_), .B(mai_mai_n493_), .Y(mai_mai_n495_));
  OA210      m0467(.A0(mai_mai_n495_), .A1(mai_mai_n491_), .B0(mai_mai_n490_), .Y(mai_mai_n496_));
  OAI220     m0468(.A0(mai_mai_n349_), .A1(mai_mai_n348_), .B0(mai_mai_n470_), .B1(mai_mai_n469_), .Y(mai_mai_n497_));
  NAi31      m0469(.An(d), .B(c), .C(a), .Y(mai_mai_n498_));
  NO2        m0470(.A(mai_mai_n498_), .B(n), .Y(mai_mai_n499_));
  NA3        m0471(.A(mai_mai_n499_), .B(mai_mai_n497_), .C(e), .Y(mai_mai_n500_));
  NO3        m0472(.A(mai_mai_n56_), .B(mai_mai_n46_), .C(mai_mai_n189_), .Y(mai_mai_n501_));
  NO2        m0473(.A(mai_mai_n204_), .B(mai_mai_n96_), .Y(mai_mai_n502_));
  NA2        m0474(.A(mai_mai_n501_), .B(mai_mai_n502_), .Y(mai_mai_n503_));
  NA2        m0475(.A(mai_mai_n503_), .B(mai_mai_n500_), .Y(mai_mai_n504_));
  NO2        m0476(.A(mai_mai_n240_), .B(n), .Y(mai_mai_n505_));
  NO2        m0477(.A(mai_mai_n378_), .B(mai_mai_n505_), .Y(mai_mai_n506_));
  NA2        m0478(.A(mai_mai_n497_), .B(f), .Y(mai_mai_n507_));
  NAi32      m0479(.An(d), .Bn(a), .C(b), .Y(mai_mai_n508_));
  NO2        m0480(.A(mai_mai_n508_), .B(mai_mai_n46_), .Y(mai_mai_n509_));
  NA2        m0481(.A(h), .B(f), .Y(mai_mai_n510_));
  NO2        m0482(.A(mai_mai_n510_), .B(mai_mai_n82_), .Y(mai_mai_n511_));
  NO3        m0483(.A(mai_mai_n155_), .B(mai_mai_n152_), .C(m), .Y(mai_mai_n512_));
  AOI220     m0484(.A0(mai_mai_n512_), .A1(mai_mai_n53_), .B0(mai_mai_n511_), .B1(mai_mai_n509_), .Y(mai_mai_n513_));
  OAI210     m0485(.A0(mai_mai_n507_), .A1(mai_mai_n506_), .B0(mai_mai_n513_), .Y(mai_mai_n514_));
  AN3        m0486(.A(j), .B(h), .C(m), .Y(mai_mai_n515_));
  NO2        m0487(.A(mai_mai_n129_), .B(c), .Y(mai_mai_n516_));
  NA3        m0488(.A(mai_mai_n516_), .B(mai_mai_n515_), .C(mai_mai_n409_), .Y(mai_mai_n517_));
  NA3        m0489(.A(f), .B(d), .C(b), .Y(mai_mai_n518_));
  NO4        m0490(.A(mai_mai_n518_), .B(mai_mai_n155_), .C(mai_mai_n152_), .D(m), .Y(mai_mai_n519_));
  INV        m0491(.A(mai_mai_n517_), .Y(mai_mai_n520_));
  NO4        m0492(.A(mai_mai_n520_), .B(mai_mai_n514_), .C(mai_mai_n504_), .D(mai_mai_n496_), .Y(mai_mai_n521_));
  AN2        m0493(.A(mai_mai_n521_), .B(mai_mai_n478_), .Y(mai_mai_n522_));
  INV        m0494(.A(k), .Y(mai_mai_n523_));
  NA3        m0495(.A(l), .B(mai_mai_n523_), .C(i), .Y(mai_mai_n524_));
  INV        m0496(.A(mai_mai_n524_), .Y(mai_mai_n525_));
  NA4        m0497(.A(mai_mai_n346_), .B(mai_mai_n367_), .C(mai_mai_n160_), .D(mai_mai_n99_), .Y(mai_mai_n526_));
  NAi32      m0498(.An(h), .Bn(f), .C(m), .Y(mai_mai_n527_));
  NAi41      m0499(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n528_));
  OAI210     m0500(.A0(mai_mai_n476_), .A1(n), .B0(mai_mai_n528_), .Y(mai_mai_n529_));
  NA2        m0501(.A(mai_mai_n529_), .B(m), .Y(mai_mai_n530_));
  NAi31      m0502(.An(h), .B(m), .C(f), .Y(mai_mai_n531_));
  OR3        m0503(.A(mai_mai_n531_), .B(mai_mai_n240_), .C(mai_mai_n46_), .Y(mai_mai_n532_));
  NA4        m0504(.A(mai_mai_n367_), .B(mai_mai_n107_), .C(mai_mai_n99_), .D(e), .Y(mai_mai_n533_));
  AN2        m0505(.A(mai_mai_n533_), .B(mai_mai_n532_), .Y(mai_mai_n534_));
  OA210      m0506(.A0(mai_mai_n530_), .A1(mai_mai_n527_), .B0(mai_mai_n534_), .Y(mai_mai_n535_));
  NA2        m0507(.A(mai_mai_n535_), .B(mai_mai_n526_), .Y(mai_mai_n536_));
  NAi31      m0508(.An(f), .B(h), .C(m), .Y(mai_mai_n537_));
  NO4        m0509(.A(mai_mai_n268_), .B(mai_mai_n537_), .C(mai_mai_n62_), .D(mai_mai_n63_), .Y(mai_mai_n538_));
  NOi32      m0510(.An(b), .Bn(a), .C(c), .Y(mai_mai_n539_));
  NOi41      m0511(.An(mai_mai_n539_), .B(mai_mai_n304_), .C(mai_mai_n59_), .D(mai_mai_n103_), .Y(mai_mai_n540_));
  OR2        m0512(.A(mai_mai_n540_), .B(mai_mai_n538_), .Y(mai_mai_n541_));
  NOi32      m0513(.An(d), .Bn(a), .C(e), .Y(mai_mai_n542_));
  NA2        m0514(.A(mai_mai_n542_), .B(mai_mai_n99_), .Y(mai_mai_n543_));
  NOi32      m0515(.An(e), .Bn(a), .C(d), .Y(mai_mai_n544_));
  AOI210     m0516(.A0(b), .A1(d), .B0(mai_mai_n544_), .Y(mai_mai_n545_));
  NO2        m0517(.A(mai_mai_n545_), .B(mai_mai_n489_), .Y(mai_mai_n546_));
  AOI210     m0518(.A0(mai_mai_n546_), .A1(mai_mai_n99_), .B0(mai_mai_n541_), .Y(mai_mai_n547_));
  INV        m0519(.A(mai_mai_n547_), .Y(mai_mai_n548_));
  AOI210     m0520(.A0(mai_mai_n536_), .A1(mai_mai_n525_), .B0(mai_mai_n548_), .Y(mai_mai_n549_));
  NO3        m0521(.A(mai_mai_n275_), .B(mai_mai_n55_), .C(n), .Y(mai_mai_n550_));
  NA3        m0522(.A(mai_mai_n454_), .B(mai_mai_n150_), .C(mai_mai_n149_), .Y(mai_mai_n551_));
  NA2        m0523(.A(mai_mai_n411_), .B(mai_mai_n204_), .Y(mai_mai_n552_));
  OR2        m0524(.A(mai_mai_n552_), .B(mai_mai_n551_), .Y(mai_mai_n553_));
  NA2        m0525(.A(k), .B(mai_mai_n99_), .Y(mai_mai_n554_));
  AOI220     m0526(.A0(mai_mai_n99_), .A1(mai_mai_n481_), .B0(mai_mai_n553_), .B1(mai_mai_n550_), .Y(mai_mai_n555_));
  NO2        m0527(.A(mai_mai_n555_), .B(mai_mai_n76_), .Y(mai_mai_n556_));
  NA3        m0528(.A(mai_mai_n491_), .B(mai_mai_n295_), .C(mai_mai_n44_), .Y(mai_mai_n557_));
  NOi32      m0529(.An(e), .Bn(c), .C(f), .Y(mai_mai_n558_));
  NOi21      m0530(.An(f), .B(m), .Y(mai_mai_n559_));
  NO2        m0531(.A(mai_mai_n559_), .B(mai_mai_n187_), .Y(mai_mai_n560_));
  AOI220     m0532(.A0(mai_mai_n560_), .A1(mai_mai_n343_), .B0(mai_mai_n558_), .B1(mai_mai_n154_), .Y(mai_mai_n561_));
  NA3        m0533(.A(mai_mai_n561_), .B(mai_mai_n557_), .C(mai_mai_n157_), .Y(mai_mai_n562_));
  AOI210     m0534(.A0(mai_mai_n480_), .A1(mai_mai_n347_), .B0(mai_mai_n258_), .Y(mai_mai_n563_));
  NA2        m0535(.A(mai_mai_n563_), .B(mai_mai_n230_), .Y(mai_mai_n564_));
  NOi21      m0536(.An(j), .B(l), .Y(mai_mai_n565_));
  NAi21      m0537(.An(k), .B(h), .Y(mai_mai_n566_));
  NO2        m0538(.A(mai_mai_n566_), .B(mai_mai_n229_), .Y(mai_mai_n567_));
  NOi31      m0539(.An(m), .B(n), .C(k), .Y(mai_mai_n568_));
  NA2        m0540(.A(mai_mai_n565_), .B(mai_mai_n568_), .Y(mai_mai_n569_));
  AOI210     m0541(.A0(mai_mai_n347_), .A1(mai_mai_n321_), .B0(mai_mai_n258_), .Y(mai_mai_n570_));
  NAi21      m0542(.An(mai_mai_n569_), .B(mai_mai_n570_), .Y(mai_mai_n571_));
  NO2        m0543(.A(mai_mai_n240_), .B(mai_mai_n46_), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n476_), .B(mai_mai_n46_), .Y(mai_mai_n573_));
  NA2        m0545(.A(mai_mai_n572_), .B(mai_mai_n511_), .Y(mai_mai_n574_));
  NA3        m0546(.A(mai_mai_n574_), .B(mai_mai_n571_), .C(mai_mai_n564_), .Y(mai_mai_n575_));
  NA2        m0547(.A(mai_mai_n94_), .B(mai_mai_n35_), .Y(mai_mai_n576_));
  NO2        m0548(.A(k), .B(mai_mai_n189_), .Y(mai_mai_n577_));
  NO2        m0549(.A(mai_mai_n472_), .B(mai_mai_n312_), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n578_), .B(n), .Y(mai_mai_n579_));
  NAi31      m0551(.An(mai_mai_n576_), .B(mai_mai_n579_), .C(mai_mai_n577_), .Y(mai_mai_n580_));
  NO2        m0552(.A(mai_mai_n474_), .B(mai_mai_n155_), .Y(mai_mai_n581_));
  NA3        m0553(.A(mai_mai_n492_), .B(mai_mai_n234_), .C(mai_mai_n128_), .Y(mai_mai_n582_));
  NA2        m0554(.A(mai_mai_n450_), .B(mai_mai_n140_), .Y(mai_mai_n583_));
  NO3        m0555(.A(mai_mai_n344_), .B(mai_mai_n583_), .C(mai_mai_n76_), .Y(mai_mai_n584_));
  AOI210     m0556(.A0(mai_mai_n582_), .A1(mai_mai_n581_), .B0(mai_mai_n584_), .Y(mai_mai_n585_));
  AN3        m0557(.A(f), .B(d), .C(b), .Y(mai_mai_n586_));
  OAI210     m0558(.A0(mai_mai_n586_), .A1(mai_mai_n115_), .B0(n), .Y(mai_mai_n587_));
  NA3        m0559(.A(mai_mai_n450_), .B(mai_mai_n140_), .C(mai_mai_n189_), .Y(mai_mai_n588_));
  AOI210     m0560(.A0(mai_mai_n587_), .A1(mai_mai_n206_), .B0(mai_mai_n588_), .Y(mai_mai_n589_));
  NAi31      m0561(.An(m), .B(n), .C(k), .Y(mai_mai_n590_));
  INV        m0562(.A(mai_mai_n220_), .Y(mai_mai_n591_));
  OAI210     m0563(.A0(mai_mai_n591_), .A1(mai_mai_n589_), .B0(j), .Y(mai_mai_n592_));
  NA3        m0564(.A(mai_mai_n592_), .B(mai_mai_n585_), .C(mai_mai_n580_), .Y(mai_mai_n593_));
  NO4        m0565(.A(mai_mai_n593_), .B(mai_mai_n575_), .C(mai_mai_n562_), .D(mai_mai_n556_), .Y(mai_mai_n594_));
  NA2        m0566(.A(mai_mai_n331_), .B(mai_mai_n142_), .Y(mai_mai_n595_));
  NAi31      m0567(.An(m), .B(h), .C(f), .Y(mai_mai_n596_));
  OR3        m0568(.A(mai_mai_n596_), .B(mai_mai_n240_), .C(n), .Y(mai_mai_n597_));
  OA210      m0569(.A0(mai_mai_n476_), .A1(n), .B0(mai_mai_n528_), .Y(mai_mai_n598_));
  NA3        m0570(.A(mai_mai_n365_), .B(mai_mai_n107_), .C(mai_mai_n73_), .Y(mai_mai_n599_));
  OAI210     m0571(.A0(mai_mai_n598_), .A1(mai_mai_n79_), .B0(mai_mai_n599_), .Y(mai_mai_n600_));
  NOi21      m0572(.An(mai_mai_n597_), .B(mai_mai_n600_), .Y(mai_mai_n601_));
  AOI210     m0573(.A0(mai_mai_n601_), .A1(mai_mai_n595_), .B0(mai_mai_n471_), .Y(mai_mai_n602_));
  NO3        m0574(.A(m), .B(mai_mai_n188_), .C(mai_mai_n51_), .Y(mai_mai_n603_));
  NAi21      m0575(.An(h), .B(j), .Y(mai_mai_n604_));
  NO2        m0576(.A(mai_mai_n458_), .B(mai_mai_n76_), .Y(mai_mai_n605_));
  OAI210     m0577(.A0(mai_mai_n605_), .A1(mai_mai_n343_), .B0(mai_mai_n603_), .Y(mai_mai_n606_));
  NA2        m0578(.A(mai_mai_n539_), .B(mai_mai_n297_), .Y(mai_mai_n607_));
  OR2        m0579(.A(mai_mai_n569_), .B(mai_mai_n607_), .Y(mai_mai_n608_));
  NA3        m0580(.A(mai_mai_n468_), .B(mai_mai_n87_), .C(mai_mai_n86_), .Y(mai_mai_n609_));
  NA2        m0581(.A(mai_mai_n87_), .B(mai_mai_n44_), .Y(mai_mai_n610_));
  NO2        m0582(.A(mai_mai_n610_), .B(mai_mai_n286_), .Y(mai_mai_n611_));
  AOI210     m0583(.A0(mai_mai_n508_), .A1(mai_mai_n377_), .B0(mai_mai_n46_), .Y(mai_mai_n612_));
  OAI220     m0584(.A0(mai_mai_n531_), .A1(mai_mai_n524_), .B0(mai_mai_n279_), .B1(mai_mai_n469_), .Y(mai_mai_n613_));
  AOI210     m0585(.A0(mai_mai_n613_), .A1(mai_mai_n612_), .B0(mai_mai_n611_), .Y(mai_mai_n614_));
  NA4        m0586(.A(mai_mai_n614_), .B(mai_mai_n609_), .C(mai_mai_n608_), .D(mai_mai_n606_), .Y(mai_mai_n615_));
  NO2        m0587(.A(mai_mai_n221_), .B(f), .Y(mai_mai_n616_));
  NO2        m0588(.A(mai_mai_n559_), .B(mai_mai_n55_), .Y(mai_mai_n617_));
  NO3        m0589(.A(mai_mai_n617_), .B(mai_mai_n616_), .C(mai_mai_n33_), .Y(mai_mai_n618_));
  NA2        m0590(.A(mai_mai_n282_), .B(mai_mai_n125_), .Y(mai_mai_n619_));
  NA2        m0591(.A(mai_mai_n117_), .B(mai_mai_n46_), .Y(mai_mai_n620_));
  NA2        m0592(.A(mai_mai_n620_), .B(mai_mai_n472_), .Y(mai_mai_n621_));
  OA220      m0593(.A0(mai_mai_n621_), .A1(mai_mai_n489_), .B0(mai_mai_n311_), .B1(mai_mai_n97_), .Y(mai_mai_n622_));
  OAI210     m0594(.A0(mai_mai_n619_), .A1(mai_mai_n618_), .B0(mai_mai_n622_), .Y(mai_mai_n623_));
  NO3        m0595(.A(mai_mai_n352_), .B(mai_mai_n172_), .C(mai_mai_n171_), .Y(mai_mai_n624_));
  NA2        m0596(.A(mai_mai_n624_), .B(mai_mai_n204_), .Y(mai_mai_n625_));
  NA3        m0597(.A(mai_mai_n625_), .B(mai_mai_n223_), .C(j), .Y(mai_mai_n626_));
  NA2        m0598(.A(mai_mai_n415_), .B(mai_mai_n73_), .Y(mai_mai_n627_));
  NO4        m0599(.A(mai_mai_n471_), .B(mai_mai_n627_), .C(mai_mai_n116_), .D(mai_mai_n188_), .Y(mai_mai_n628_));
  INV        m0600(.A(mai_mai_n628_), .Y(mai_mai_n629_));
  NA4        m0601(.A(mai_mai_n629_), .B(mai_mai_n626_), .C(mai_mai_n457_), .D(mai_mai_n350_), .Y(mai_mai_n630_));
  NO4        m0602(.A(mai_mai_n630_), .B(mai_mai_n623_), .C(mai_mai_n615_), .D(mai_mai_n602_), .Y(mai_mai_n631_));
  NA4        m0603(.A(mai_mai_n631_), .B(mai_mai_n594_), .C(mai_mai_n549_), .D(mai_mai_n522_), .Y(mai08));
  NO2        m0604(.A(k), .B(h), .Y(mai_mai_n633_));
  AO210      m0605(.A0(mai_mai_n221_), .A1(mai_mai_n401_), .B0(mai_mai_n633_), .Y(mai_mai_n634_));
  NO2        m0606(.A(mai_mai_n634_), .B(mai_mai_n256_), .Y(mai_mai_n635_));
  NA2        m0607(.A(mai_mai_n558_), .B(mai_mai_n73_), .Y(mai_mai_n636_));
  NA2        m0608(.A(mai_mai_n636_), .B(mai_mai_n411_), .Y(mai_mai_n637_));
  NA2        m0609(.A(mai_mai_n637_), .B(mai_mai_n635_), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n73_), .B(mai_mai_n96_), .Y(mai_mai_n639_));
  NO2        m0611(.A(mai_mai_n639_), .B(mai_mai_n52_), .Y(mai_mai_n640_));
  NA2        m0612(.A(mai_mai_n518_), .B(mai_mai_n206_), .Y(mai_mai_n641_));
  NA2        m0613(.A(mai_mai_n641_), .B(mai_mai_n302_), .Y(mai_mai_n642_));
  AOI210     m0614(.A0(mai_mai_n518_), .A1(mai_mai_n136_), .B0(mai_mai_n73_), .Y(mai_mai_n643_));
  NA4        m0615(.A(mai_mai_n191_), .B(mai_mai_n125_), .C(mai_mai_n43_), .D(h), .Y(mai_mai_n644_));
  AN2        m0616(.A(l), .B(k), .Y(mai_mai_n645_));
  NA4        m0617(.A(mai_mai_n645_), .B(mai_mai_n94_), .C(mai_mai_n63_), .D(mai_mai_n189_), .Y(mai_mai_n646_));
  OAI210     m0618(.A0(mai_mai_n644_), .A1(m), .B0(mai_mai_n646_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n647_), .B(mai_mai_n643_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n648_), .B(mai_mai_n642_), .C(mai_mai_n638_), .Y(mai_mai_n649_));
  NO4        m0621(.A(mai_mai_n152_), .B(mai_mai_n342_), .C(mai_mai_n98_), .D(m), .Y(mai_mai_n650_));
  AOI210     m0622(.A0(mai_mai_n650_), .A1(mai_mai_n641_), .B0(mai_mai_n463_), .Y(mai_mai_n651_));
  NO2        m0623(.A(mai_mai_n37_), .B(mai_mai_n188_), .Y(mai_mai_n652_));
  NA2        m0624(.A(mai_mai_n652_), .B(mai_mai_n505_), .Y(mai_mai_n653_));
  NA2        m0625(.A(mai_mai_n653_), .B(mai_mai_n651_), .Y(mai_mai_n654_));
  NO2        m0626(.A(mai_mai_n480_), .B(mai_mai_n34_), .Y(mai_mai_n655_));
  INV        m0627(.A(mai_mai_n655_), .Y(mai_mai_n656_));
  NA2        m0628(.A(mai_mai_n634_), .B(mai_mai_n121_), .Y(mai_mai_n657_));
  NA2        m0629(.A(mai_mai_n657_), .B(mai_mai_n351_), .Y(mai_mai_n658_));
  OAI210     m0630(.A0(mai_mai_n656_), .A1(mai_mai_n76_), .B0(mai_mai_n658_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n312_), .B(mai_mai_n42_), .Y(mai_mai_n660_));
  NA3        m0632(.A(mai_mai_n625_), .B(mai_mai_n288_), .C(mai_mai_n334_), .Y(mai_mai_n661_));
  NA2        m0633(.A(mai_mai_n645_), .B(mai_mai_n194_), .Y(mai_mai_n662_));
  NO2        m0634(.A(mai_mai_n662_), .B(mai_mai_n281_), .Y(mai_mai_n663_));
  AOI210     m0635(.A0(mai_mai_n663_), .A1(mai_mai_n616_), .B0(mai_mai_n436_), .Y(mai_mai_n664_));
  NA3        m0636(.A(m), .B(l), .C(k), .Y(mai_mai_n665_));
  AOI210     m0637(.A0(mai_mai_n599_), .A1(mai_mai_n597_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  NO2        m0638(.A(mai_mai_n479_), .B(mai_mai_n235_), .Y(mai_mai_n667_));
  NOi21      m0639(.An(mai_mai_n667_), .B(mai_mai_n473_), .Y(mai_mai_n668_));
  NA4        m0640(.A(mai_mai_n99_), .B(l), .C(k), .D(mai_mai_n76_), .Y(mai_mai_n669_));
  NA3        m0641(.A(mai_mai_n107_), .B(mai_mai_n360_), .C(i), .Y(mai_mai_n670_));
  NO2        m0642(.A(mai_mai_n670_), .B(mai_mai_n669_), .Y(mai_mai_n671_));
  NO3        m0643(.A(mai_mai_n671_), .B(mai_mai_n668_), .C(mai_mai_n666_), .Y(mai_mai_n672_));
  NA4        m0644(.A(mai_mai_n672_), .B(mai_mai_n664_), .C(mai_mai_n661_), .D(mai_mai_n660_), .Y(mai_mai_n673_));
  NO4        m0645(.A(mai_mai_n673_), .B(mai_mai_n659_), .C(mai_mai_n654_), .D(mai_mai_n649_), .Y(mai_mai_n674_));
  NA2        m0646(.A(mai_mai_n560_), .B(mai_mai_n343_), .Y(mai_mai_n675_));
  NA2        m0647(.A(mai_mai_n573_), .B(m), .Y(mai_mai_n676_));
  AO210      m0648(.A0(mai_mai_n676_), .A1(mai_mai_n532_), .B0(mai_mai_n482_), .Y(mai_mai_n677_));
  NO3        m0649(.A(mai_mai_n347_), .B(mai_mai_n469_), .C(h), .Y(mai_mai_n678_));
  AOI210     m0650(.A0(mai_mai_n678_), .A1(mai_mai_n99_), .B0(mai_mai_n444_), .Y(mai_mai_n679_));
  NA4        m0651(.A(mai_mai_n679_), .B(mai_mai_n677_), .C(mai_mai_n675_), .D(mai_mai_n220_), .Y(mai_mai_n680_));
  NA2        m0652(.A(mai_mai_n645_), .B(mai_mai_n63_), .Y(mai_mai_n681_));
  NO4        m0653(.A(mai_mai_n624_), .B(mai_mai_n152_), .C(n), .D(i), .Y(mai_mai_n682_));
  NOi21      m0654(.An(h), .B(j), .Y(mai_mai_n683_));
  NA2        m0655(.A(mai_mai_n683_), .B(f), .Y(mai_mai_n684_));
  NO2        m0656(.A(mai_mai_n684_), .B(mai_mai_n217_), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n685_), .B(mai_mai_n682_), .Y(mai_mai_n686_));
  OAI220     m0658(.A0(mai_mai_n686_), .A1(mai_mai_n681_), .B0(mai_mai_n534_), .B1(mai_mai_n56_), .Y(mai_mai_n687_));
  AOI210     m0659(.A0(mai_mai_n680_), .A1(l), .B0(mai_mai_n687_), .Y(mai_mai_n688_));
  NO2        m0660(.A(j), .B(i), .Y(mai_mai_n689_));
  NA2        m0661(.A(mai_mai_n689_), .B(mai_mai_n32_), .Y(mai_mai_n690_));
  NA2        m0662(.A(mai_mai_n370_), .B(mai_mai_n107_), .Y(mai_mai_n691_));
  OR2        m0663(.A(mai_mai_n691_), .B(mai_mai_n690_), .Y(mai_mai_n692_));
  NO3        m0664(.A(mai_mai_n133_), .B(mai_mai_n46_), .C(mai_mai_n96_), .Y(mai_mai_n693_));
  NO3        m0665(.A(mai_mai_n486_), .B(mai_mai_n131_), .C(mai_mai_n63_), .Y(mai_mai_n694_));
  NO2        m0666(.A(mai_mai_n432_), .B(mai_mai_n389_), .Y(mai_mai_n695_));
  NO2        m0667(.A(mai_mai_n676_), .B(mai_mai_n56_), .Y(mai_mai_n696_));
  NA2        m0668(.A(k), .B(j), .Y(mai_mai_n697_));
  NO3        m0669(.A(mai_mai_n256_), .B(mai_mai_n697_), .C(mai_mai_n39_), .Y(mai_mai_n698_));
  AOI210     m0670(.A0(mai_mai_n472_), .A1(n), .B0(mai_mai_n491_), .Y(mai_mai_n699_));
  NA2        m0671(.A(mai_mai_n699_), .B(mai_mai_n494_), .Y(mai_mai_n700_));
  AN3        m0672(.A(mai_mai_n700_), .B(mai_mai_n698_), .C(mai_mai_n86_), .Y(mai_mai_n701_));
  NA2        m0673(.A(mai_mai_n552_), .B(mai_mai_n265_), .Y(mai_mai_n702_));
  INV        m0674(.A(mai_mai_n702_), .Y(mai_mai_n703_));
  NO2        m0675(.A(mai_mai_n256_), .B(mai_mai_n121_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n704_), .B(mai_mai_n560_), .Y(mai_mai_n705_));
  NO2        m0677(.A(mai_mai_n665_), .B(mai_mai_n79_), .Y(mai_mai_n706_));
  NO2        m0678(.A(mai_mai_n531_), .B(mai_mai_n103_), .Y(mai_mai_n707_));
  OAI210     m0679(.A0(mai_mai_n707_), .A1(mai_mai_n695_), .B0(mai_mai_n612_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n708_), .B(mai_mai_n705_), .Y(mai_mai_n709_));
  OR4        m0681(.A(mai_mai_n709_), .B(mai_mai_n703_), .C(mai_mai_n701_), .D(mai_mai_n696_), .Y(mai_mai_n710_));
  NA3        m0682(.A(mai_mai_n699_), .B(mai_mai_n494_), .C(mai_mai_n493_), .Y(mai_mai_n711_));
  NA4        m0683(.A(mai_mai_n711_), .B(mai_mai_n191_), .C(mai_mai_n401_), .D(mai_mai_n33_), .Y(mai_mai_n712_));
  NO3        m0684(.A(mai_mai_n432_), .B(mai_mai_n384_), .C(j), .Y(mai_mai_n713_));
  OAI220     m0685(.A0(mai_mai_n644_), .A1(mai_mai_n636_), .B0(mai_mai_n286_), .B1(mai_mai_n37_), .Y(mai_mai_n714_));
  AOI210     m0686(.A0(mai_mai_n713_), .A1(mai_mai_n227_), .B0(mai_mai_n714_), .Y(mai_mai_n715_));
  NA3        m0687(.A(mai_mai_n487_), .B(mai_mai_n250_), .C(h), .Y(mai_mai_n716_));
  NOi21      m0688(.An(mai_mai_n612_), .B(mai_mai_n716_), .Y(mai_mai_n717_));
  NO2        m0689(.A(mai_mai_n80_), .B(mai_mai_n45_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n579_), .Y(mai_mai_n719_));
  NAi41      m0691(.An(mai_mai_n717_), .B(mai_mai_n719_), .C(mai_mai_n715_), .D(mai_mai_n712_), .Y(mai_mai_n720_));
  OR2        m0692(.A(mai_mai_n706_), .B(mai_mai_n83_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n721_), .B(mai_mai_n211_), .Y(mai_mai_n722_));
  INV        m0694(.A(mai_mai_n290_), .Y(mai_mai_n723_));
  NO2        m0695(.A(mai_mai_n716_), .B(mai_mai_n435_), .Y(mai_mai_n724_));
  INV        m0696(.A(mai_mai_n724_), .Y(mai_mai_n725_));
  NA3        m0697(.A(mai_mai_n725_), .B(mai_mai_n723_), .C(mai_mai_n722_), .Y(mai_mai_n726_));
  NOi41      m0698(.An(mai_mai_n692_), .B(mai_mai_n726_), .C(mai_mai_n720_), .D(mai_mai_n710_), .Y(mai_mai_n727_));
  OR3        m0699(.A(mai_mai_n644_), .B(mai_mai_n206_), .C(m), .Y(mai_mai_n728_));
  NO3        m0700(.A(mai_mai_n296_), .B(mai_mai_n258_), .C(mai_mai_n98_), .Y(mai_mai_n729_));
  NA2        m0701(.A(mai_mai_n729_), .B(mai_mai_n700_), .Y(mai_mai_n730_));
  INV        m0702(.A(mai_mai_n44_), .Y(mai_mai_n731_));
  NO3        m0703(.A(mai_mai_n731_), .B(mai_mai_n690_), .C(mai_mai_n240_), .Y(mai_mai_n732_));
  NO3        m0704(.A(mai_mai_n469_), .B(mai_mai_n81_), .C(h), .Y(mai_mai_n733_));
  AOI210     m0705(.A0(mai_mai_n733_), .A1(mai_mai_n640_), .B0(mai_mai_n732_), .Y(mai_mai_n734_));
  NA4        m0706(.A(mai_mai_n734_), .B(mai_mai_n730_), .C(mai_mai_n728_), .D(mai_mai_n353_), .Y(mai_mai_n735_));
  OR2        m0707(.A(mai_mai_n596_), .B(mai_mai_n80_), .Y(mai_mai_n736_));
  NOi31      m0708(.An(b), .B(d), .C(a), .Y(mai_mai_n737_));
  NO2        m0709(.A(mai_mai_n737_), .B(mai_mai_n542_), .Y(mai_mai_n738_));
  NO2        m0710(.A(mai_mai_n738_), .B(n), .Y(mai_mai_n739_));
  INV        m0711(.A(mai_mai_n739_), .Y(mai_mai_n740_));
  NO2        m0712(.A(mai_mai_n740_), .B(mai_mai_n736_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n492_), .B(mai_mai_n73_), .Y(mai_mai_n742_));
  NO3        m0714(.A(mai_mai_n559_), .B(mai_mai_n281_), .C(mai_mai_n103_), .Y(mai_mai_n743_));
  NOi21      m0715(.An(mai_mai_n743_), .B(mai_mai_n141_), .Y(mai_mai_n744_));
  AOI210     m0716(.A0(mai_mai_n729_), .A1(mai_mai_n742_), .B0(mai_mai_n744_), .Y(mai_mai_n745_));
  OAI210     m0717(.A0(mai_mai_n644_), .A1(mai_mai_n344_), .B0(mai_mai_n745_), .Y(mai_mai_n746_));
  NO2        m0718(.A(mai_mai_n624_), .B(n), .Y(mai_mai_n747_));
  AOI220     m0719(.A0(mai_mai_n704_), .A1(mai_mai_n603_), .B0(mai_mai_n747_), .B1(mai_mai_n635_), .Y(mai_mai_n748_));
  NO2        m0720(.A(mai_mai_n277_), .B(mai_mai_n210_), .Y(mai_mai_n749_));
  NA2        m0721(.A(mai_mai_n107_), .B(mai_mai_n73_), .Y(mai_mai_n750_));
  AOI210     m0722(.A0(mai_mai_n374_), .A1(mai_mai_n366_), .B0(mai_mai_n750_), .Y(mai_mai_n751_));
  NA2        m0723(.A(mai_mai_n663_), .B(mai_mai_n33_), .Y(mai_mai_n752_));
  NAi21      m0724(.An(mai_mai_n669_), .B(mai_mai_n385_), .Y(mai_mai_n753_));
  NO2        m0725(.A(mai_mai_n235_), .B(i), .Y(mai_mai_n754_));
  NAi41      m0726(.An(mai_mai_n751_), .B(mai_mai_n753_), .C(mai_mai_n752_), .D(mai_mai_n748_), .Y(mai_mai_n755_));
  NO4        m0727(.A(mai_mai_n755_), .B(mai_mai_n746_), .C(mai_mai_n741_), .D(mai_mai_n735_), .Y(mai_mai_n756_));
  NA4        m0728(.A(mai_mai_n756_), .B(mai_mai_n727_), .C(mai_mai_n688_), .D(mai_mai_n674_), .Y(mai09));
  INV        m0729(.A(mai_mai_n108_), .Y(mai_mai_n758_));
  NA2        m0730(.A(f), .B(e), .Y(mai_mai_n759_));
  NO2        m0731(.A(mai_mai_n199_), .B(mai_mai_n98_), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n760_), .B(m), .Y(mai_mai_n761_));
  NA3        m0733(.A(mai_mai_n268_), .B(mai_mai_n228_), .C(mai_mai_n105_), .Y(mai_mai_n762_));
  AOI210     m0734(.A0(mai_mai_n762_), .A1(m), .B0(mai_mai_n421_), .Y(mai_mai_n763_));
  AOI210     m0735(.A0(mai_mai_n763_), .A1(mai_mai_n761_), .B0(mai_mai_n759_), .Y(mai_mai_n764_));
  NA2        m0736(.A(mai_mai_n764_), .B(mai_mai_n758_), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n184_), .B(mai_mai_n188_), .Y(mai_mai_n766_));
  NA3        m0738(.A(m), .B(l), .C(i), .Y(mai_mai_n767_));
  OAI220     m0739(.A0(mai_mai_n531_), .A1(mai_mai_n767_), .B0(mai_mai_n304_), .B1(mai_mai_n470_), .Y(mai_mai_n768_));
  NA4        m0740(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(m), .D(f), .Y(mai_mai_n769_));
  NAi31      m0741(.An(mai_mai_n768_), .B(mai_mai_n769_), .C(mai_mai_n390_), .Y(mai_mai_n770_));
  OR2        m0742(.A(mai_mai_n770_), .B(mai_mai_n766_), .Y(mai_mai_n771_));
  NA3        m0743(.A(mai_mai_n736_), .B(mai_mai_n507_), .C(mai_mai_n462_), .Y(mai_mai_n772_));
  OA210      m0744(.A0(mai_mai_n772_), .A1(mai_mai_n771_), .B0(mai_mai_n739_), .Y(mai_mai_n773_));
  INV        m0745(.A(mai_mai_n293_), .Y(mai_mai_n774_));
  NO2        m0746(.A(mai_mai_n112_), .B(mai_mai_n111_), .Y(mai_mai_n775_));
  NOi31      m0747(.An(k), .B(m), .C(l), .Y(mai_mai_n776_));
  NO2        m0748(.A(mai_mai_n295_), .B(mai_mai_n776_), .Y(mai_mai_n777_));
  AOI210     m0749(.A0(mai_mai_n777_), .A1(mai_mai_n775_), .B0(mai_mai_n537_), .Y(mai_mai_n778_));
  INV        m0750(.A(mai_mai_n286_), .Y(mai_mai_n779_));
  NA2        m0751(.A(mai_mai_n297_), .B(mai_mai_n299_), .Y(mai_mai_n780_));
  OAI210     m0752(.A0(mai_mai_n184_), .A1(mai_mai_n188_), .B0(mai_mai_n780_), .Y(mai_mai_n781_));
  AOI220     m0753(.A0(mai_mai_n781_), .A1(mai_mai_n779_), .B0(mai_mai_n778_), .B1(mai_mai_n774_), .Y(mai_mai_n782_));
  NA2        m0754(.A(mai_mai_n146_), .B(mai_mai_n100_), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n783_), .B(mai_mai_n634_), .C(mai_mai_n121_), .Y(mai_mai_n784_));
  NA3        m0756(.A(mai_mai_n784_), .B(mai_mai_n169_), .C(mai_mai_n30_), .Y(mai_mai_n785_));
  NA4        m0757(.A(mai_mai_n785_), .B(mai_mai_n782_), .C(mai_mai_n561_), .D(mai_mai_n71_), .Y(mai_mai_n786_));
  NO2        m0758(.A(mai_mai_n527_), .B(mai_mai_n441_), .Y(mai_mai_n787_));
  NA2        m0759(.A(mai_mai_n787_), .B(mai_mai_n169_), .Y(mai_mai_n788_));
  NOi21      m0760(.An(f), .B(d), .Y(mai_mai_n789_));
  NA2        m0761(.A(mai_mai_n789_), .B(m), .Y(mai_mai_n790_));
  NOi32      m0762(.An(m), .Bn(f), .C(d), .Y(mai_mai_n791_));
  INV        m0763(.A(mai_mai_n228_), .Y(mai_mai_n792_));
  AN2        m0764(.A(f), .B(d), .Y(mai_mai_n793_));
  NA3        m0765(.A(mai_mai_n426_), .B(mai_mai_n793_), .C(mai_mai_n73_), .Y(mai_mai_n794_));
  NO3        m0766(.A(mai_mai_n794_), .B(mai_mai_n63_), .C(mai_mai_n189_), .Y(mai_mai_n795_));
  NO2        m0767(.A(i), .B(mai_mai_n51_), .Y(mai_mai_n796_));
  NA2        m0768(.A(mai_mai_n792_), .B(mai_mai_n795_), .Y(mai_mai_n797_));
  NAi31      m0769(.An(mai_mai_n434_), .B(mai_mai_n797_), .C(mai_mai_n788_), .Y(mai_mai_n798_));
  NO4        m0770(.A(mai_mai_n559_), .B(mai_mai_n117_), .C(mai_mai_n281_), .D(mai_mai_n134_), .Y(mai_mai_n799_));
  NO2        m0771(.A(mai_mai_n590_), .B(mai_mai_n281_), .Y(mai_mai_n800_));
  AN2        m0772(.A(mai_mai_n800_), .B(mai_mai_n616_), .Y(mai_mai_n801_));
  NO2        m0773(.A(mai_mai_n801_), .B(mai_mai_n799_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n542_), .B(mai_mai_n73_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n780_), .B(mai_mai_n803_), .Y(mai_mai_n804_));
  NA3        m0776(.A(mai_mai_n140_), .B(mai_mai_n94_), .C(m), .Y(mai_mai_n805_));
  OAI220     m0777(.A0(mai_mai_n794_), .A1(mai_mai_n379_), .B0(mai_mai_n293_), .B1(mai_mai_n805_), .Y(mai_mai_n806_));
  NOi41      m0778(.An(mai_mai_n197_), .B(mai_mai_n806_), .C(mai_mai_n804_), .D(mai_mai_n263_), .Y(mai_mai_n807_));
  NA2        m0779(.A(c), .B(mai_mai_n102_), .Y(mai_mai_n808_));
  NO2        m0780(.A(mai_mai_n808_), .B(mai_mai_n357_), .Y(mai_mai_n809_));
  NA3        m0781(.A(mai_mai_n809_), .B(mai_mai_n452_), .C(f), .Y(mai_mai_n810_));
  OR2        m0782(.A(mai_mai_n596_), .B(mai_mai_n483_), .Y(mai_mai_n811_));
  INV        m0783(.A(mai_mai_n811_), .Y(mai_mai_n812_));
  NA2        m0784(.A(mai_mai_n738_), .B(mai_mai_n97_), .Y(mai_mai_n813_));
  NA2        m0785(.A(mai_mai_n813_), .B(mai_mai_n812_), .Y(mai_mai_n814_));
  NA4        m0786(.A(mai_mai_n814_), .B(mai_mai_n810_), .C(mai_mai_n807_), .D(mai_mai_n802_), .Y(mai_mai_n815_));
  NO4        m0787(.A(mai_mai_n815_), .B(mai_mai_n798_), .C(mai_mai_n786_), .D(mai_mai_n773_), .Y(mai_mai_n816_));
  OR2        m0788(.A(mai_mai_n794_), .B(mai_mai_n63_), .Y(mai_mai_n817_));
  NA2        m0789(.A(mai_mai_n98_), .B(j), .Y(mai_mai_n818_));
  NA2        m0790(.A(mai_mai_n760_), .B(m), .Y(mai_mai_n819_));
  AOI210     m0791(.A0(mai_mai_n819_), .A1(mai_mai_n251_), .B0(mai_mai_n817_), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n204_), .B(mai_mai_n198_), .Y(mai_mai_n821_));
  NA2        m0793(.A(mai_mai_n821_), .B(mai_mai_n201_), .Y(mai_mai_n822_));
  NO2        m0794(.A(mai_mai_n379_), .B(mai_mai_n759_), .Y(mai_mai_n823_));
  NA2        m0795(.A(mai_mai_n823_), .B(mai_mai_n499_), .Y(mai_mai_n824_));
  NA2        m0796(.A(mai_mai_n824_), .B(mai_mai_n822_), .Y(mai_mai_n825_));
  NA2        m0797(.A(e), .B(d), .Y(mai_mai_n826_));
  OAI220     m0798(.A0(mai_mai_n826_), .A1(c), .B0(mai_mai_n277_), .B1(d), .Y(mai_mai_n827_));
  NA3        m0799(.A(mai_mai_n827_), .B(mai_mai_n404_), .C(mai_mai_n450_), .Y(mai_mai_n828_));
  AOI210     m0800(.A0(mai_mai_n458_), .A1(mai_mai_n159_), .B0(mai_mai_n204_), .Y(mai_mai_n829_));
  INV        m0801(.A(mai_mai_n829_), .Y(mai_mai_n830_));
  NA3        m0802(.A(mai_mai_n145_), .B(mai_mai_n74_), .C(mai_mai_n33_), .Y(mai_mai_n831_));
  NA3        m0803(.A(mai_mai_n831_), .B(mai_mai_n830_), .C(mai_mai_n828_), .Y(mai_mai_n832_));
  NO3        m0804(.A(mai_mai_n832_), .B(mai_mai_n825_), .C(mai_mai_n820_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n774_), .B(mai_mai_n30_), .Y(mai_mai_n834_));
  AO210      m0806(.A0(mai_mai_n834_), .A1(mai_mai_n636_), .B0(mai_mai_n192_), .Y(mai_mai_n835_));
  OAI220     m0807(.A0(mai_mai_n559_), .A1(mai_mai_n55_), .B0(mai_mai_n258_), .B1(j), .Y(mai_mai_n836_));
  AOI220     m0808(.A0(mai_mai_n836_), .A1(mai_mai_n800_), .B0(mai_mai_n550_), .B1(mai_mai_n558_), .Y(mai_mai_n837_));
  INV        m0809(.A(mai_mai_n837_), .Y(mai_mai_n838_));
  AN2        m0810(.A(mai_mai_n779_), .B(mai_mai_n768_), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n839_), .B(mai_mai_n838_), .Y(mai_mai_n840_));
  AO220      m0812(.A0(mai_mai_n404_), .A1(mai_mai_n683_), .B0(mai_mai_n154_), .B1(f), .Y(mai_mai_n841_));
  OAI210     m0813(.A0(mai_mai_n841_), .A1(mai_mai_n407_), .B0(mai_mai_n827_), .Y(mai_mai_n842_));
  NA2        m0814(.A(mai_mai_n772_), .B(mai_mai_n640_), .Y(mai_mai_n843_));
  AN4        m0815(.A(mai_mai_n843_), .B(mai_mai_n842_), .C(mai_mai_n840_), .D(mai_mai_n835_), .Y(mai_mai_n844_));
  NA4        m0816(.A(mai_mai_n844_), .B(mai_mai_n833_), .C(mai_mai_n816_), .D(mai_mai_n765_), .Y(mai12));
  NO2        m0817(.A(mai_mai_n402_), .B(c), .Y(mai_mai_n846_));
  NO4        m0818(.A(mai_mai_n394_), .B(mai_mai_n221_), .C(mai_mai_n523_), .D(mai_mai_n189_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n847_), .B(mai_mai_n846_), .Y(mai_mai_n848_));
  NO2        m0820(.A(mai_mai_n402_), .B(mai_mai_n102_), .Y(mai_mai_n849_));
  NO2        m0821(.A(mai_mai_n596_), .B(mai_mai_n328_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n848_), .B(mai_mai_n393_), .Y(mai_mai_n851_));
  AOI210     m0823(.A0(mai_mai_n207_), .A1(mai_mai_n292_), .B0(mai_mai_n181_), .Y(mai_mai_n852_));
  OR2        m0824(.A(mai_mai_n852_), .B(mai_mai_n847_), .Y(mai_mai_n853_));
  AOI210     m0825(.A0(mai_mai_n289_), .A1(mai_mai_n340_), .B0(mai_mai_n189_), .Y(mai_mai_n854_));
  OAI210     m0826(.A0(mai_mai_n854_), .A1(mai_mai_n853_), .B0(mai_mai_n352_), .Y(mai_mai_n855_));
  NO2        m0827(.A(mai_mai_n576_), .B(mai_mai_n229_), .Y(mai_mai_n856_));
  NO2        m0828(.A(mai_mai_n531_), .B(mai_mai_n767_), .Y(mai_mai_n857_));
  AOI220     m0829(.A0(mai_mai_n857_), .A1(mai_mai_n505_), .B0(mai_mai_n749_), .B1(mai_mai_n856_), .Y(mai_mai_n858_));
  NO2        m0830(.A(mai_mai_n133_), .B(mai_mai_n210_), .Y(mai_mai_n859_));
  NA2        m0831(.A(mai_mai_n858_), .B(mai_mai_n855_), .Y(mai_mai_n860_));
  OR2        m0832(.A(mai_mai_n278_), .B(mai_mai_n849_), .Y(mai_mai_n861_));
  NA2        m0833(.A(mai_mai_n861_), .B(mai_mai_n305_), .Y(mai_mai_n862_));
  NO3        m0834(.A(mai_mai_n117_), .B(mai_mai_n134_), .C(mai_mai_n189_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n863_), .B(mai_mai_n472_), .Y(mai_mai_n864_));
  NA2        m0836(.A(mai_mai_n864_), .B(mai_mai_n862_), .Y(mai_mai_n865_));
  NO3        m0837(.A(mai_mai_n601_), .B(mai_mai_n80_), .C(mai_mai_n43_), .Y(mai_mai_n866_));
  NO4        m0838(.A(mai_mai_n866_), .B(mai_mai_n865_), .C(mai_mai_n860_), .D(mai_mai_n851_), .Y(mai_mai_n867_));
  NO2        m0839(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n868_));
  NA2        m0840(.A(mai_mai_n528_), .B(mai_mai_n62_), .Y(mai_mai_n869_));
  NA2        m0841(.A(mai_mai_n492_), .B(mai_mai_n128_), .Y(mai_mai_n870_));
  NOi21      m0842(.An(mai_mai_n33_), .B(mai_mai_n590_), .Y(mai_mai_n871_));
  AOI220     m0843(.A0(mai_mai_n871_), .A1(mai_mai_n870_), .B0(mai_mai_n869_), .B1(mai_mai_n868_), .Y(mai_mai_n872_));
  OAI210     m0844(.A0(mai_mai_n220_), .A1(mai_mai_n43_), .B0(mai_mai_n872_), .Y(mai_mai_n873_));
  NA2        m0845(.A(mai_mai_n385_), .B(mai_mai_n230_), .Y(mai_mai_n874_));
  NO3        m0846(.A(mai_mai_n750_), .B(mai_mai_n78_), .C(mai_mai_n357_), .Y(mai_mai_n875_));
  NAi21      m0847(.An(mai_mai_n875_), .B(mai_mai_n874_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n46_), .B(mai_mai_n43_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n447_), .B(mai_mai_n258_), .Y(mai_mai_n878_));
  INV        m0850(.A(mai_mai_n878_), .Y(mai_mai_n879_));
  NO2        m0851(.A(mai_mai_n879_), .B(mai_mai_n128_), .Y(mai_mai_n880_));
  NA2        m0852(.A(mai_mai_n568_), .B(j), .Y(mai_mai_n881_));
  INV        m0853(.A(mai_mai_n316_), .Y(mai_mai_n882_));
  NO4        m0854(.A(mai_mai_n882_), .B(mai_mai_n880_), .C(mai_mai_n876_), .D(mai_mai_n873_), .Y(mai_mai_n883_));
  NA2        m0855(.A(mai_mai_n301_), .B(m), .Y(mai_mai_n884_));
  NA2        m0856(.A(mai_mai_n142_), .B(i), .Y(mai_mai_n885_));
  NA2        m0857(.A(mai_mai_n44_), .B(i), .Y(mai_mai_n886_));
  OAI220     m0858(.A0(mai_mai_n886_), .A1(mai_mai_n180_), .B0(mai_mai_n885_), .B1(mai_mai_n80_), .Y(mai_mai_n887_));
  AOI210     m0859(.A0(mai_mai_n368_), .A1(mai_mai_n36_), .B0(mai_mai_n887_), .Y(mai_mai_n888_));
  NO2        m0860(.A(mai_mai_n128_), .B(mai_mai_n73_), .Y(mai_mai_n889_));
  OR2        m0861(.A(mai_mai_n889_), .B(mai_mai_n491_), .Y(mai_mai_n890_));
  NA2        m0862(.A(mai_mai_n492_), .B(mai_mai_n332_), .Y(mai_mai_n891_));
  AOI210     m0863(.A0(mai_mai_n891_), .A1(n), .B0(mai_mai_n890_), .Y(mai_mai_n892_));
  OAI220     m0864(.A0(mai_mai_n892_), .A1(mai_mai_n884_), .B0(mai_mai_n888_), .B1(mai_mai_n286_), .Y(mai_mai_n893_));
  NO2        m0865(.A(mai_mai_n596_), .B(mai_mai_n441_), .Y(mai_mai_n894_));
  NA3        m0866(.A(mai_mai_n297_), .B(mai_mai_n565_), .C(i), .Y(mai_mai_n895_));
  OAI210     m0867(.A0(mai_mai_n389_), .A1(mai_mai_n268_), .B0(mai_mai_n895_), .Y(mai_mai_n896_));
  OAI220     m0868(.A0(mai_mai_n896_), .A1(mai_mai_n894_), .B0(mai_mai_n612_), .B1(mai_mai_n694_), .Y(mai_mai_n897_));
  OR3        m0869(.A(mai_mai_n268_), .B(mai_mai_n384_), .C(f), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n627_), .B(mai_mai_n803_), .Y(mai_mai_n899_));
  NA2        m0871(.A(mai_mai_n769_), .B(mai_mai_n390_), .Y(mai_mai_n900_));
  NA2        m0872(.A(mai_mai_n195_), .B(mai_mai_n66_), .Y(mai_mai_n901_));
  NA2        m0873(.A(mai_mai_n901_), .B(mai_mai_n898_), .Y(mai_mai_n902_));
  AOI220     m0874(.A0(mai_mai_n902_), .A1(mai_mai_n227_), .B0(mai_mai_n900_), .B1(mai_mai_n899_), .Y(mai_mai_n903_));
  NA2        m0875(.A(mai_mai_n903_), .B(mai_mai_n897_), .Y(mai_mai_n904_));
  NO2        m0876(.A(mai_mai_n328_), .B(mai_mai_n79_), .Y(mai_mai_n905_));
  OAI210     m0877(.A0(mai_mai_n905_), .A1(mai_mai_n856_), .B0(mai_mai_n211_), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n600_), .B(mai_mai_n77_), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n410_), .B(mai_mai_n189_), .Y(mai_mai_n908_));
  AOI220     m0880(.A0(mai_mai_n908_), .A1(mai_mai_n333_), .B0(mai_mai_n861_), .B1(mai_mai_n193_), .Y(mai_mai_n909_));
  NA2        m0881(.A(mai_mai_n850_), .B(mai_mai_n859_), .Y(mai_mai_n910_));
  NA4        m0882(.A(mai_mai_n910_), .B(mai_mai_n909_), .C(mai_mai_n907_), .D(mai_mai_n906_), .Y(mai_mai_n911_));
  OAI210     m0883(.A0(mai_mai_n900_), .A1(mai_mai_n857_), .B0(mai_mai_n485_), .Y(mai_mai_n912_));
  AOI210     m0884(.A0(mai_mai_n369_), .A1(mai_mai_n361_), .B0(mai_mai_n750_), .Y(mai_mai_n913_));
  OAI210     m0885(.A0(mai_mai_n319_), .A1(mai_mai_n318_), .B0(mai_mai_n95_), .Y(mai_mai_n914_));
  AOI210     m0886(.A0(mai_mai_n914_), .A1(mai_mai_n477_), .B0(mai_mai_n913_), .Y(mai_mai_n915_));
  NO3        m0887(.A(mai_mai_n818_), .B(mai_mai_n46_), .C(mai_mai_n43_), .Y(mai_mai_n916_));
  AOI220     m0888(.A0(mai_mai_n916_), .A1(mai_mai_n563_), .B0(mai_mai_n581_), .B1(mai_mai_n472_), .Y(mai_mai_n917_));
  NA3        m0889(.A(mai_mai_n917_), .B(mai_mai_n915_), .C(mai_mai_n912_), .Y(mai_mai_n918_));
  NO4        m0890(.A(mai_mai_n918_), .B(mai_mai_n911_), .C(mai_mai_n904_), .D(mai_mai_n893_), .Y(mai_mai_n919_));
  NAi31      m0891(.An(mai_mai_n126_), .B(mai_mai_n370_), .C(n), .Y(mai_mai_n920_));
  NO3        m0892(.A(mai_mai_n111_), .B(mai_mai_n295_), .C(mai_mai_n776_), .Y(mai_mai_n921_));
  NO2        m0893(.A(mai_mai_n921_), .B(mai_mai_n920_), .Y(mai_mai_n922_));
  NO3        m0894(.A(mai_mai_n235_), .B(mai_mai_n126_), .C(mai_mai_n357_), .Y(mai_mai_n923_));
  AOI210     m0895(.A0(mai_mai_n923_), .A1(mai_mai_n442_), .B0(mai_mai_n922_), .Y(mai_mai_n924_));
  INV        m0896(.A(mai_mai_n924_), .Y(mai_mai_n925_));
  NA2        m0897(.A(mai_mai_n204_), .B(mai_mai_n150_), .Y(mai_mai_n926_));
  NO3        m0898(.A(mai_mai_n265_), .B(mai_mai_n395_), .C(mai_mai_n154_), .Y(mai_mai_n927_));
  NOi31      m0899(.An(mai_mai_n926_), .B(mai_mai_n927_), .C(mai_mai_n189_), .Y(mai_mai_n928_));
  NAi21      m0900(.An(mai_mai_n492_), .B(mai_mai_n908_), .Y(mai_mai_n929_));
  NO3        m0901(.A(mai_mai_n389_), .B(mai_mai_n268_), .C(mai_mai_n63_), .Y(mai_mai_n930_));
  AOI220     m0902(.A0(mai_mai_n930_), .A1(mai_mai_n386_), .B0(mai_mai_n430_), .B1(m), .Y(mai_mai_n931_));
  NA2        m0903(.A(mai_mai_n931_), .B(mai_mai_n929_), .Y(mai_mai_n932_));
  OAI220     m0904(.A0(mai_mai_n920_), .A1(mai_mai_n207_), .B0(mai_mai_n895_), .B1(mai_mai_n543_), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n597_), .B(mai_mai_n328_), .Y(mai_mai_n934_));
  NA2        m0906(.A(mai_mai_n852_), .B(mai_mai_n846_), .Y(mai_mai_n935_));
  NO3        m0907(.A(mai_mai_n486_), .B(mai_mai_n131_), .C(mai_mai_n188_), .Y(mai_mai_n936_));
  OAI210     m0908(.A0(mai_mai_n936_), .A1(mai_mai_n468_), .B0(mai_mai_n329_), .Y(mai_mai_n937_));
  NA3        m0909(.A(mai_mai_n937_), .B(mai_mai_n935_), .C(mai_mai_n557_), .Y(mai_mai_n938_));
  OAI210     m0910(.A0(mai_mai_n852_), .A1(mai_mai_n847_), .B0(mai_mai_n926_), .Y(mai_mai_n939_));
  NA3        m0911(.A(mai_mai_n891_), .B(mai_mai_n433_), .C(mai_mai_n44_), .Y(mai_mai_n940_));
  AOI210     m0912(.A0(mai_mai_n331_), .A1(mai_mai_n329_), .B0(mai_mai_n285_), .Y(mai_mai_n941_));
  NA4        m0913(.A(mai_mai_n941_), .B(mai_mai_n940_), .C(mai_mai_n939_), .D(mai_mai_n236_), .Y(mai_mai_n942_));
  OR4        m0914(.A(mai_mai_n942_), .B(mai_mai_n938_), .C(mai_mai_n934_), .D(mai_mai_n933_), .Y(mai_mai_n943_));
  NO4        m0915(.A(mai_mai_n943_), .B(mai_mai_n932_), .C(mai_mai_n928_), .D(mai_mai_n925_), .Y(mai_mai_n944_));
  NA4        m0916(.A(mai_mai_n944_), .B(mai_mai_n919_), .C(mai_mai_n883_), .D(mai_mai_n867_), .Y(mai13));
  AN2        m0917(.A(c), .B(b), .Y(mai_mai_n946_));
  NA3        m0918(.A(mai_mai_n219_), .B(mai_mai_n946_), .C(m), .Y(mai_mai_n947_));
  NA2        m0919(.A(mai_mai_n440_), .B(f), .Y(mai_mai_n948_));
  NO3        m0920(.A(mai_mai_n948_), .B(mai_mai_n947_), .C(mai_mai_n524_), .Y(mai_mai_n949_));
  NAi32      m0921(.An(d), .Bn(c), .C(e), .Y(mai_mai_n950_));
  NA2        m0922(.A(mai_mai_n125_), .B(mai_mai_n43_), .Y(mai_mai_n951_));
  NO4        m0923(.A(mai_mai_n951_), .B(mai_mai_n950_), .C(mai_mai_n531_), .D(mai_mai_n264_), .Y(mai_mai_n952_));
  NA2        m0924(.A(mai_mai_n604_), .B(mai_mai_n198_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n360_), .B(mai_mai_n188_), .Y(mai_mai_n954_));
  AN2        m0926(.A(d), .B(c), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n955_), .B(mai_mai_n102_), .Y(mai_mai_n956_));
  NO4        m0928(.A(mai_mai_n956_), .B(mai_mai_n954_), .C(mai_mai_n155_), .D(mai_mai_n146_), .Y(mai_mai_n957_));
  NA2        m0929(.A(mai_mai_n440_), .B(c), .Y(mai_mai_n958_));
  NO4        m0930(.A(mai_mai_n951_), .B(mai_mai_n527_), .C(mai_mai_n958_), .D(mai_mai_n264_), .Y(mai_mai_n959_));
  AO210      m0931(.A0(mai_mai_n957_), .A1(mai_mai_n953_), .B0(mai_mai_n959_), .Y(mai_mai_n960_));
  OR3        m0932(.A(mai_mai_n960_), .B(mai_mai_n952_), .C(mai_mai_n949_), .Y(mai_mai_n961_));
  NAi32      m0933(.An(f), .Bn(e), .C(c), .Y(mai_mai_n962_));
  NO2        m0934(.A(mai_mai_n962_), .B(mai_mai_n129_), .Y(mai_mai_n963_));
  NA2        m0935(.A(mai_mai_n963_), .B(m), .Y(mai_mai_n964_));
  OR3        m0936(.A(mai_mai_n198_), .B(mai_mai_n155_), .C(mai_mai_n146_), .Y(mai_mai_n965_));
  NO2        m0937(.A(mai_mai_n965_), .B(mai_mai_n964_), .Y(mai_mai_n966_));
  NO2        m0938(.A(mai_mai_n958_), .B(mai_mai_n264_), .Y(mai_mai_n967_));
  NO2        m0939(.A(j), .B(mai_mai_n43_), .Y(mai_mai_n968_));
  NA2        m0940(.A(mai_mai_n567_), .B(mai_mai_n968_), .Y(mai_mai_n969_));
  NOi21      m0941(.An(mai_mai_n967_), .B(mai_mai_n969_), .Y(mai_mai_n970_));
  NO2        m0942(.A(mai_mai_n697_), .B(mai_mai_n98_), .Y(mai_mai_n971_));
  NOi41      m0943(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n972_));
  NA2        m0944(.A(mai_mai_n972_), .B(mai_mai_n971_), .Y(mai_mai_n973_));
  NO2        m0945(.A(mai_mai_n973_), .B(mai_mai_n964_), .Y(mai_mai_n974_));
  OR3        m0946(.A(e), .B(d), .C(c), .Y(mai_mai_n975_));
  NA3        m0947(.A(k), .B(j), .C(i), .Y(mai_mai_n976_));
  NO3        m0948(.A(mai_mai_n976_), .B(mai_mai_n264_), .C(mai_mai_n79_), .Y(mai_mai_n977_));
  NOi21      m0949(.An(mai_mai_n977_), .B(mai_mai_n975_), .Y(mai_mai_n978_));
  OR4        m0950(.A(mai_mai_n978_), .B(mai_mai_n974_), .C(mai_mai_n970_), .D(mai_mai_n966_), .Y(mai_mai_n979_));
  NA3        m0951(.A(mai_mai_n418_), .B(mai_mai_n288_), .C(mai_mai_n51_), .Y(mai_mai_n980_));
  NO2        m0952(.A(mai_mai_n980_), .B(mai_mai_n969_), .Y(mai_mai_n981_));
  NO4        m0953(.A(mai_mai_n980_), .B(mai_mai_n527_), .C(mai_mai_n401_), .D(mai_mai_n43_), .Y(mai_mai_n982_));
  NO2        m0954(.A(f), .B(c), .Y(mai_mai_n983_));
  NOi21      m0955(.An(mai_mai_n983_), .B(mai_mai_n394_), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n984_), .B(mai_mai_n54_), .Y(mai_mai_n985_));
  OR2        m0957(.A(k), .B(i), .Y(mai_mai_n986_));
  NO3        m0958(.A(mai_mai_n986_), .B(mai_mai_n214_), .C(l), .Y(mai_mai_n987_));
  NOi31      m0959(.An(mai_mai_n987_), .B(mai_mai_n985_), .C(j), .Y(mai_mai_n988_));
  OR3        m0960(.A(mai_mai_n988_), .B(mai_mai_n982_), .C(mai_mai_n981_), .Y(mai_mai_n989_));
  OR3        m0961(.A(mai_mai_n989_), .B(mai_mai_n979_), .C(mai_mai_n961_), .Y(mai02));
  OR2        m0962(.A(l), .B(k), .Y(mai_mai_n991_));
  OR3        m0963(.A(h), .B(m), .C(f), .Y(mai_mai_n992_));
  OR3        m0964(.A(n), .B(m), .C(i), .Y(mai_mai_n993_));
  NO4        m0965(.A(mai_mai_n993_), .B(mai_mai_n992_), .C(mai_mai_n991_), .D(mai_mai_n975_), .Y(mai_mai_n994_));
  NOi31      m0966(.An(e), .B(d), .C(c), .Y(mai_mai_n995_));
  AOI210     m0967(.A0(mai_mai_n977_), .A1(mai_mai_n995_), .B0(mai_mai_n952_), .Y(mai_mai_n996_));
  AN3        m0968(.A(m), .B(f), .C(c), .Y(mai_mai_n997_));
  NA3        m0969(.A(mai_mai_n997_), .B(mai_mai_n418_), .C(h), .Y(mai_mai_n998_));
  OR2        m0970(.A(mai_mai_n976_), .B(mai_mai_n264_), .Y(mai_mai_n999_));
  OR2        m0971(.A(mai_mai_n999_), .B(mai_mai_n998_), .Y(mai_mai_n1000_));
  NO3        m0972(.A(mai_mai_n980_), .B(mai_mai_n951_), .C(mai_mai_n527_), .Y(mai_mai_n1001_));
  NO2        m0973(.A(mai_mai_n1001_), .B(mai_mai_n966_), .Y(mai_mai_n1002_));
  NA3        m0974(.A(l), .B(k), .C(j), .Y(mai_mai_n1003_));
  NA2        m0975(.A(i), .B(h), .Y(mai_mai_n1004_));
  NO3        m0976(.A(mai_mai_n1004_), .B(mai_mai_n1003_), .C(mai_mai_n117_), .Y(mai_mai_n1005_));
  NO3        m0977(.A(mai_mai_n127_), .B(mai_mai_n247_), .C(mai_mai_n189_), .Y(mai_mai_n1006_));
  AOI210     m0978(.A0(mai_mai_n1006_), .A1(mai_mai_n1005_), .B0(mai_mai_n970_), .Y(mai_mai_n1007_));
  NA3        m0979(.A(c), .B(b), .C(a), .Y(mai_mai_n1008_));
  NO3        m0980(.A(mai_mai_n1008_), .B(mai_mai_n826_), .C(mai_mai_n188_), .Y(mai_mai_n1009_));
  NO3        m0981(.A(mai_mai_n976_), .B(mai_mai_n46_), .C(mai_mai_n98_), .Y(mai_mai_n1010_));
  AOI210     m0982(.A0(mai_mai_n1010_), .A1(mai_mai_n1009_), .B0(mai_mai_n981_), .Y(mai_mai_n1011_));
  AN4        m0983(.A(mai_mai_n1011_), .B(mai_mai_n1007_), .C(mai_mai_n1002_), .D(mai_mai_n1000_), .Y(mai_mai_n1012_));
  NO2        m0984(.A(mai_mai_n956_), .B(mai_mai_n954_), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n973_), .B(mai_mai_n965_), .Y(mai_mai_n1014_));
  AOI210     m0986(.A0(mai_mai_n1014_), .A1(mai_mai_n1013_), .B0(mai_mai_n949_), .Y(mai_mai_n1015_));
  NAi41      m0987(.An(mai_mai_n994_), .B(mai_mai_n1015_), .C(mai_mai_n1012_), .D(mai_mai_n996_), .Y(mai03));
  INV        m0988(.A(mai_mai_n914_), .Y(mai_mai_n1017_));
  NOi41      m0989(.An(mai_mai_n736_), .B(mai_mai_n781_), .C(mai_mai_n770_), .D(mai_mai_n652_), .Y(mai_mai_n1018_));
  OAI220     m0990(.A0(mai_mai_n1018_), .A1(mai_mai_n627_), .B0(mai_mai_n1017_), .B1(mai_mai_n528_), .Y(mai_mai_n1019_));
  NA4        m0991(.A(i), .B(mai_mai_n995_), .C(mai_mai_n297_), .D(mai_mai_n288_), .Y(mai_mai_n1020_));
  OAI210     m0992(.A0(mai_mai_n750_), .A1(mai_mai_n371_), .B0(mai_mai_n1020_), .Y(mai_mai_n1021_));
  NOi31      m0993(.An(m), .B(n), .C(f), .Y(mai_mai_n1022_));
  NA2        m0994(.A(mai_mai_n450_), .B(l), .Y(mai_mai_n1023_));
  NOi31      m0995(.An(mai_mai_n791_), .B(mai_mai_n947_), .C(mai_mai_n1023_), .Y(mai_mai_n1024_));
  NO3        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1021_), .C(mai_mai_n913_), .Y(mai_mai_n1025_));
  NO2        m0997(.A(mai_mai_n247_), .B(a), .Y(mai_mai_n1026_));
  INV        m0998(.A(mai_mai_n952_), .Y(mai_mai_n1027_));
  NO2        m0999(.A(mai_mai_n1004_), .B(mai_mai_n432_), .Y(mai_mai_n1028_));
  NO2        m1000(.A(mai_mai_n76_), .B(m), .Y(mai_mai_n1029_));
  AOI210     m1001(.A0(mai_mai_n1029_), .A1(mai_mai_n1028_), .B0(mai_mai_n987_), .Y(mai_mai_n1030_));
  OR2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n985_), .Y(mai_mai_n1031_));
  NA3        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1027_), .C(mai_mai_n1025_), .Y(mai_mai_n1032_));
  NO4        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1019_), .C(mai_mai_n751_), .D(mai_mai_n504_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(c), .B(b), .Y(mai_mai_n1034_));
  NO2        m1006(.A(mai_mai_n639_), .B(mai_mai_n1034_), .Y(mai_mai_n1035_));
  OAI210     m1007(.A0(mai_mai_n790_), .A1(mai_mai_n763_), .B0(mai_mai_n364_), .Y(mai_mai_n1036_));
  NA2        m1008(.A(mai_mai_n1036_), .B(mai_mai_n1035_), .Y(mai_mai_n1037_));
  NAi21      m1009(.An(mai_mai_n372_), .B(mai_mai_n1035_), .Y(mai_mai_n1038_));
  OAI210     m1010(.A0(mai_mai_n488_), .A1(mai_mai_n38_), .B0(mai_mai_n1026_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n1039_), .B(mai_mai_n1038_), .Y(mai_mai_n1040_));
  NAi21      m1012(.An(f), .B(d), .Y(mai_mai_n1041_));
  NO2        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1008_), .Y(mai_mai_n1042_));
  INV        m1014(.A(mai_mai_n1042_), .Y(mai_mai_n1043_));
  NO2        m1015(.A(mai_mai_n251_), .B(mai_mai_n1043_), .Y(mai_mai_n1044_));
  AOI210     m1016(.A0(mai_mai_n1044_), .A1(mai_mai_n99_), .B0(mai_mai_n1040_), .Y(mai_mai_n1045_));
  NA2        m1017(.A(mai_mai_n421_), .B(mai_mai_n420_), .Y(mai_mai_n1046_));
  NO2        m1018(.A(mai_mai_n161_), .B(mai_mai_n210_), .Y(mai_mai_n1047_));
  NA2        m1019(.A(mai_mai_n1047_), .B(m), .Y(mai_mai_n1048_));
  INV        m1020(.A(mai_mai_n422_), .Y(mai_mai_n1049_));
  AOI210     m1021(.A0(mai_mai_n1049_), .A1(mai_mai_n1046_), .B0(mai_mai_n1048_), .Y(mai_mai_n1050_));
  NA2        m1022(.A(mai_mai_n499_), .B(mai_mai_n359_), .Y(mai_mai_n1051_));
  NA2        m1023(.A(mai_mai_n139_), .B(mai_mai_n32_), .Y(mai_mai_n1052_));
  AOI210     m1024(.A0(mai_mai_n881_), .A1(mai_mai_n1052_), .B0(mai_mai_n189_), .Y(mai_mai_n1053_));
  OAI210     m1025(.A0(mai_mai_n1053_), .A1(mai_mai_n398_), .B0(mai_mai_n1042_), .Y(mai_mai_n1054_));
  NO2        m1026(.A(mai_mai_n322_), .B(mai_mai_n321_), .Y(mai_mai_n1055_));
  AOI210     m1027(.A0(mai_mai_n1047_), .A1(mai_mai_n380_), .B0(mai_mai_n875_), .Y(mai_mai_n1056_));
  NAi41      m1028(.An(mai_mai_n1055_), .B(mai_mai_n1056_), .C(mai_mai_n1054_), .D(mai_mai_n1051_), .Y(mai_mai_n1057_));
  NO2        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1050_), .Y(mai_mai_n1058_));
  NA4        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1045_), .C(mai_mai_n1037_), .D(mai_mai_n1033_), .Y(mai00));
  AOI210     m1031(.A0(mai_mai_n257_), .A1(mai_mai_n189_), .B0(mai_mai_n239_), .Y(mai_mai_n1060_));
  NO2        m1032(.A(mai_mai_n1060_), .B(mai_mai_n518_), .Y(mai_mai_n1061_));
  AOI210     m1033(.A0(mai_mai_n823_), .A1(mai_mai_n859_), .B0(mai_mai_n1021_), .Y(mai_mai_n1062_));
  NO2        m1034(.A(mai_mai_n1001_), .B(mai_mai_n875_), .Y(mai_mai_n1063_));
  NA3        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1062_), .C(mai_mai_n915_), .Y(mai_mai_n1064_));
  NA2        m1036(.A(mai_mai_n452_), .B(f), .Y(mai_mai_n1065_));
  OAI210     m1037(.A0(mai_mai_n921_), .A1(mai_mai_n39_), .B0(mai_mai_n583_), .Y(mai_mai_n1066_));
  NA3        m1038(.A(mai_mai_n1066_), .B(mai_mai_n226_), .C(n), .Y(mai_mai_n1067_));
  AOI210     m1039(.A0(mai_mai_n1067_), .A1(mai_mai_n1065_), .B0(mai_mai_n956_), .Y(mai_mai_n1068_));
  NO4        m1040(.A(mai_mai_n1068_), .B(mai_mai_n1064_), .C(mai_mai_n1061_), .D(mai_mai_n979_), .Y(mai_mai_n1069_));
  NA3        m1041(.A(mai_mai_n145_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n1070_));
  NA3        m1042(.A(d), .B(mai_mai_n51_), .C(b), .Y(mai_mai_n1071_));
  NOi31      m1043(.An(n), .B(m), .C(i), .Y(mai_mai_n1072_));
  NA3        m1044(.A(mai_mai_n1072_), .B(mai_mai_n586_), .C(mai_mai_n48_), .Y(mai_mai_n1073_));
  OAI210     m1045(.A0(mai_mai_n1071_), .A1(mai_mai_n1070_), .B0(mai_mai_n1073_), .Y(mai_mai_n1074_));
  INV        m1046(.A(mai_mai_n517_), .Y(mai_mai_n1075_));
  NO3        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1074_), .C(mai_mai_n1055_), .Y(mai_mai_n1076_));
  NA3        m1048(.A(mai_mai_n334_), .B(mai_mai_n194_), .C(m), .Y(mai_mai_n1077_));
  OA220      m1049(.A0(mai_mai_n1077_), .A1(mai_mai_n1071_), .B0(mai_mai_n335_), .B1(mai_mai_n120_), .Y(mai_mai_n1078_));
  NO2        m1050(.A(h), .B(m), .Y(mai_mai_n1079_));
  NA4        m1051(.A(mai_mai_n442_), .B(mai_mai_n418_), .C(mai_mai_n1079_), .D(mai_mai_n946_), .Y(mai_mai_n1080_));
  NA2        m1052(.A(mai_mai_n863_), .B(mai_mai_n516_), .Y(mai_mai_n1081_));
  NA3        m1053(.A(mai_mai_n1081_), .B(mai_mai_n1080_), .C(mai_mai_n1078_), .Y(mai_mai_n1082_));
  INV        m1054(.A(mai_mai_n1082_), .Y(mai_mai_n1083_));
  NO2        m1055(.A(mai_mai_n212_), .B(mai_mai_n160_), .Y(mai_mai_n1084_));
  NA2        m1056(.A(mai_mai_n1084_), .B(mai_mai_n378_), .Y(mai_mai_n1085_));
  NA3        m1057(.A(mai_mai_n158_), .B(mai_mai_n98_), .C(m), .Y(mai_mai_n1086_));
  NA3        m1058(.A(mai_mai_n418_), .B(mai_mai_n39_), .C(f), .Y(mai_mai_n1087_));
  NOi31      m1059(.An(mai_mai_n796_), .B(mai_mai_n1087_), .C(mai_mai_n1086_), .Y(mai_mai_n1088_));
  NAi31      m1060(.An(mai_mai_n165_), .B(mai_mai_n787_), .C(mai_mai_n418_), .Y(mai_mai_n1089_));
  NAi31      m1061(.An(mai_mai_n1088_), .B(mai_mai_n1089_), .C(mai_mai_n1085_), .Y(mai_mai_n1090_));
  NO2        m1062(.A(mai_mai_n238_), .B(mai_mai_n63_), .Y(mai_mai_n1091_));
  NO3        m1063(.A(mai_mai_n377_), .B(mai_mai_n759_), .C(n), .Y(mai_mai_n1092_));
  AOI210     m1064(.A0(mai_mai_n1092_), .A1(mai_mai_n1091_), .B0(mai_mai_n994_), .Y(mai_mai_n1093_));
  NAi21      m1065(.An(mai_mai_n959_), .B(mai_mai_n1093_), .Y(mai_mai_n1094_));
  NO3        m1066(.A(mai_mai_n1094_), .B(mai_mai_n1090_), .C(mai_mai_n519_), .Y(mai_mai_n1095_));
  AN3        m1067(.A(mai_mai_n1095_), .B(mai_mai_n1083_), .C(mai_mai_n1076_), .Y(mai_mai_n1096_));
  INV        m1068(.A(mai_mai_n500_), .Y(mai_mai_n1097_));
  NA2        m1069(.A(mai_mai_n499_), .B(mai_mai_n359_), .Y(mai_mai_n1098_));
  OR4        m1070(.A(mai_mai_n956_), .B(mai_mai_n235_), .C(mai_mai_n196_), .D(e), .Y(mai_mai_n1099_));
  NO2        m1071(.A(mai_mai_n192_), .B(mai_mai_n189_), .Y(mai_mai_n1100_));
  NA2        m1072(.A(n), .B(e), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n1101_), .B(mai_mai_n129_), .Y(mai_mai_n1102_));
  AOI220     m1074(.A0(mai_mai_n1102_), .A1(mai_mai_n237_), .B0(mai_mai_n774_), .B1(mai_mai_n1100_), .Y(mai_mai_n1103_));
  OAI210     m1075(.A0(mai_mai_n308_), .A1(mai_mai_n270_), .B0(mai_mai_n400_), .Y(mai_mai_n1104_));
  NA4        m1076(.A(mai_mai_n1104_), .B(mai_mai_n1103_), .C(mai_mai_n1099_), .D(mai_mai_n1098_), .Y(mai_mai_n1105_));
  AOI210     m1077(.A0(mai_mai_n1102_), .A1(mai_mai_n778_), .B0(mai_mai_n751_), .Y(mai_mai_n1106_));
  AOI220     m1078(.A0(mai_mai_n871_), .A1(mai_mai_n516_), .B0(mai_mai_n586_), .B1(mai_mai_n215_), .Y(mai_mai_n1107_));
  NO2        m1079(.A(mai_mai_n58_), .B(h), .Y(mai_mai_n1108_));
  NO3        m1080(.A(mai_mai_n956_), .B(mai_mai_n954_), .C(mai_mai_n662_), .Y(mai_mai_n1109_));
  NO2        m1081(.A(mai_mai_n991_), .B(mai_mai_n117_), .Y(mai_mai_n1110_));
  AN2        m1082(.A(mai_mai_n1110_), .B(mai_mai_n1006_), .Y(mai_mai_n1111_));
  OAI210     m1083(.A0(mai_mai_n1111_), .A1(mai_mai_n1109_), .B0(mai_mai_n1108_), .Y(mai_mai_n1112_));
  NA3        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1107_), .C(mai_mai_n1106_), .Y(mai_mai_n1113_));
  NO4        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1105_), .C(mai_mai_n253_), .D(mai_mai_n1097_), .Y(mai_mai_n1114_));
  NA2        m1086(.A(mai_mai_n764_), .B(mai_mai_n693_), .Y(mai_mai_n1115_));
  NA4        m1087(.A(mai_mai_n1115_), .B(mai_mai_n1114_), .C(mai_mai_n1096_), .D(mai_mai_n1069_), .Y(mai01));
  AN2        m1088(.A(mai_mai_n937_), .B(mai_mai_n935_), .Y(mai_mai_n1117_));
  NO4        m1089(.A(mai_mai_n732_), .B(mai_mai_n724_), .C(mai_mai_n429_), .D(mai_mai_n245_), .Y(mai_mai_n1118_));
  NO2        m1090(.A(mai_mai_n533_), .B(mai_mai_n248_), .Y(mai_mai_n1119_));
  OAI210     m1091(.A0(mai_mai_n1119_), .A1(mai_mai_n345_), .B0(i), .Y(mai_mai_n1120_));
  NA3        m1092(.A(mai_mai_n1120_), .B(mai_mai_n1118_), .C(mai_mai_n1117_), .Y(mai_mai_n1121_));
  NA2        m1093(.A(mai_mai_n492_), .B(mai_mai_n234_), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n878_), .B(mai_mai_n1122_), .Y(mai_mai_n1123_));
  NA3        m1095(.A(mai_mai_n1123_), .B(mai_mai_n837_), .C(mai_mai_n287_), .Y(mai_mai_n1124_));
  NA2        m1096(.A(mai_mai_n645_), .B(mai_mai_n84_), .Y(mai_mai_n1125_));
  NO2        m1097(.A(mai_mai_n1125_), .B(mai_mai_n1409_), .Y(mai_mai_n1126_));
  NA2        m1098(.A(mai_mai_n1126_), .B(mai_mai_n572_), .Y(mai_mai_n1127_));
  INV        m1099(.A(mai_mai_n104_), .Y(mai_mai_n1128_));
  OR2        m1100(.A(mai_mai_n1128_), .B(mai_mai_n526_), .Y(mai_mai_n1129_));
  NA3        m1101(.A(mai_mai_n1129_), .B(mai_mai_n1127_), .C(mai_mai_n822_), .Y(mai_mai_n1130_));
  NO3        m1102(.A(mai_mai_n717_), .B(mai_mai_n611_), .C(mai_mai_n455_), .Y(mai_mai_n1131_));
  OR2        m1103(.A(mai_mai_n175_), .B(mai_mai_n173_), .Y(mai_mai_n1132_));
  NA3        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1131_), .C(mai_mai_n123_), .Y(mai_mai_n1133_));
  NO4        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1130_), .C(mai_mai_n1124_), .D(mai_mai_n1121_), .Y(mai_mai_n1134_));
  INV        m1106(.A(mai_mai_n1077_), .Y(mai_mai_n1135_));
  OAI210     m1107(.A0(mai_mai_n1135_), .A1(mai_mai_n260_), .B0(mai_mai_n472_), .Y(mai_mai_n1136_));
  NA2        m1108(.A(mai_mai_n480_), .B(mai_mai_n347_), .Y(mai_mai_n1137_));
  NOi21      m1109(.An(mai_mai_n501_), .B(mai_mai_n523_), .Y(mai_mai_n1138_));
  NA2        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1137_), .Y(mai_mai_n1139_));
  AOI210     m1111(.A0(mai_mai_n184_), .A1(mai_mai_n78_), .B0(mai_mai_n188_), .Y(mai_mai_n1140_));
  OAI210     m1112(.A0(mai_mai_n739_), .A1(mai_mai_n378_), .B0(mai_mai_n1140_), .Y(mai_mai_n1141_));
  AN3        m1113(.A(m), .B(l), .C(k), .Y(mai_mai_n1142_));
  OAI210     m1114(.A0(mai_mai_n310_), .A1(mai_mai_n33_), .B0(mai_mai_n1142_), .Y(mai_mai_n1143_));
  NA2        m1115(.A(mai_mai_n183_), .B(mai_mai_n33_), .Y(mai_mai_n1144_));
  AO210      m1116(.A0(mai_mai_n1144_), .A1(mai_mai_n1143_), .B0(mai_mai_n286_), .Y(mai_mai_n1145_));
  NA4        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1141_), .C(mai_mai_n1139_), .D(mai_mai_n1136_), .Y(mai_mai_n1146_));
  INV        m1118(.A(mai_mai_n541_), .Y(mai_mai_n1147_));
  OAI210     m1119(.A0(mai_mai_n1128_), .A1(mai_mai_n535_), .B0(mai_mai_n1147_), .Y(mai_mai_n1148_));
  NA2        m1120(.A(mai_mai_n244_), .B(mai_mai_n175_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n1149_), .B(mai_mai_n603_), .Y(mai_mai_n1150_));
  NO3        m1122(.A(mai_mai_n750_), .B(mai_mai_n184_), .C(mai_mai_n357_), .Y(mai_mai_n1151_));
  NO2        m1123(.A(mai_mai_n1151_), .B(mai_mai_n875_), .Y(mai_mai_n1152_));
  OAI210     m1124(.A0(mai_mai_n1126_), .A1(mai_mai_n280_), .B0(mai_mai_n612_), .Y(mai_mai_n1153_));
  NA4        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1152_), .C(mai_mai_n1150_), .D(mai_mai_n719_), .Y(mai_mai_n1154_));
  NO3        m1126(.A(mai_mai_n1154_), .B(mai_mai_n1148_), .C(mai_mai_n1146_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n448_), .B(mai_mai_n53_), .Y(mai_mai_n1156_));
  INV        m1128(.A(mai_mai_n1074_), .Y(mai_mai_n1157_));
  NA3        m1129(.A(mai_mai_n1157_), .B(mai_mai_n1156_), .C(mai_mai_n692_), .Y(mai_mai_n1158_));
  NO2        m1130(.A(mai_mai_n885_), .B(mai_mai_n206_), .Y(mai_mai_n1159_));
  NO2        m1131(.A(mai_mai_n886_), .B(mai_mai_n494_), .Y(mai_mai_n1160_));
  OAI210     m1132(.A0(mai_mai_n1160_), .A1(mai_mai_n1159_), .B0(mai_mai_n295_), .Y(mai_mai_n1161_));
  NA2        m1133(.A(mai_mai_n511_), .B(mai_mai_n509_), .Y(mai_mai_n1162_));
  NO3        m1134(.A(mai_mai_n68_), .B(mai_mai_n258_), .C(mai_mai_n43_), .Y(mai_mai_n1163_));
  NA2        m1135(.A(mai_mai_n1163_), .B(mai_mai_n491_), .Y(mai_mai_n1164_));
  NA3        m1136(.A(mai_mai_n1164_), .B(mai_mai_n1162_), .C(mai_mai_n608_), .Y(mai_mai_n1165_));
  OR2        m1137(.A(mai_mai_n1077_), .B(mai_mai_n1071_), .Y(mai_mai_n1166_));
  NA2        m1138(.A(mai_mai_n1163_), .B(mai_mai_n742_), .Y(mai_mai_n1167_));
  NA3        m1139(.A(mai_mai_n1167_), .B(mai_mai_n1166_), .C(mai_mai_n337_), .Y(mai_mai_n1168_));
  NOi41      m1140(.An(mai_mai_n1161_), .B(mai_mai_n1168_), .C(mai_mai_n1165_), .D(mai_mai_n1158_), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n116_), .B(mai_mai_n43_), .Y(mai_mai_n1170_));
  NO2        m1142(.A(mai_mai_n43_), .B(mai_mai_n39_), .Y(mai_mai_n1171_));
  AO220      m1143(.A0(mai_mai_n1171_), .A1(mai_mai_n560_), .B0(mai_mai_n1170_), .B1(mai_mai_n643_), .Y(mai_mai_n1172_));
  NA2        m1144(.A(mai_mai_n1172_), .B(mai_mai_n295_), .Y(mai_mai_n1173_));
  NO3        m1145(.A(mai_mai_n1004_), .B(mai_mai_n155_), .C(mai_mai_n76_), .Y(mai_mai_n1174_));
  NA2        m1146(.A(mai_mai_n1163_), .B(mai_mai_n889_), .Y(mai_mai_n1175_));
  NA2        m1147(.A(mai_mai_n1175_), .B(mai_mai_n1173_), .Y(mai_mai_n1176_));
  NO2        m1148(.A(mai_mai_n552_), .B(mai_mai_n551_), .Y(mai_mai_n1177_));
  NO4        m1149(.A(mai_mai_n1004_), .B(mai_mai_n1177_), .C(mai_mai_n153_), .D(mai_mai_n76_), .Y(mai_mai_n1178_));
  NO3        m1150(.A(mai_mai_n1178_), .B(mai_mai_n1176_), .C(mai_mai_n575_), .Y(mai_mai_n1179_));
  NA4        m1151(.A(mai_mai_n1179_), .B(mai_mai_n1169_), .C(mai_mai_n1155_), .D(mai_mai_n1134_), .Y(mai06));
  NO2        m1152(.A(mai_mai_n358_), .B(mai_mai_n498_), .Y(mai_mai_n1181_));
  INV        m1153(.A(mai_mai_n669_), .Y(mai_mai_n1182_));
  NA2        m1154(.A(mai_mai_n1182_), .B(mai_mai_n1181_), .Y(mai_mai_n1183_));
  NO2        m1155(.A(mai_mai_n198_), .B(mai_mai_n89_), .Y(mai_mai_n1184_));
  OAI210     m1156(.A0(mai_mai_n1184_), .A1(mai_mai_n1174_), .B0(mai_mai_n333_), .Y(mai_mai_n1185_));
  NO3        m1157(.A(mai_mai_n539_), .B(mai_mai_n737_), .C(mai_mai_n542_), .Y(mai_mai_n1186_));
  OR2        m1158(.A(mai_mai_n1186_), .B(mai_mai_n811_), .Y(mai_mai_n1187_));
  NA4        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1185_), .C(mai_mai_n1183_), .D(mai_mai_n1161_), .Y(mai_mai_n1188_));
  NO3        m1160(.A(mai_mai_n1188_), .B(mai_mai_n1165_), .C(mai_mai_n225_), .Y(mai_mai_n1189_));
  NO2        m1161(.A(mai_mai_n258_), .B(mai_mai_n43_), .Y(mai_mai_n1190_));
  AOI210     m1162(.A0(mai_mai_n1190_), .A1(mai_mai_n890_), .B0(mai_mai_n1159_), .Y(mai_mai_n1191_));
  AOI210     m1163(.A0(mai_mai_n1190_), .A1(mai_mai_n495_), .B0(mai_mai_n1172_), .Y(mai_mai_n1192_));
  AOI210     m1164(.A0(mai_mai_n1192_), .A1(mai_mai_n1191_), .B0(mai_mai_n292_), .Y(mai_mai_n1193_));
  INV        m1165(.A(mai_mai_n610_), .Y(mai_mai_n1194_));
  NA2        m1166(.A(mai_mai_n1194_), .B(mai_mai_n579_), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n458_), .B(mai_mai_n150_), .Y(mai_mai_n1196_));
  NOi21      m1168(.An(mai_mai_n122_), .B(mai_mai_n43_), .Y(mai_mai_n1197_));
  OAI210     m1169(.A0(mai_mai_n411_), .A1(mai_mai_n218_), .B0(mai_mai_n831_), .Y(mai_mai_n1198_));
  NO3        m1170(.A(mai_mai_n1198_), .B(mai_mai_n1197_), .C(mai_mai_n1196_), .Y(mai_mai_n1199_));
  OR2        m1171(.A(mai_mai_n540_), .B(mai_mai_n538_), .Y(mai_mai_n1200_));
  INV        m1172(.A(mai_mai_n1200_), .Y(mai_mai_n1201_));
  NA3        m1173(.A(mai_mai_n1201_), .B(mai_mai_n1199_), .C(mai_mai_n1195_), .Y(mai_mai_n1202_));
  NO2        m1174(.A(mai_mai_n684_), .B(mai_mai_n318_), .Y(mai_mai_n1203_));
  NO3        m1175(.A(mai_mai_n612_), .B(mai_mai_n694_), .C(mai_mai_n572_), .Y(mai_mai_n1204_));
  NOi21      m1176(.An(mai_mai_n1203_), .B(mai_mai_n1204_), .Y(mai_mai_n1205_));
  AN2        m1177(.A(mai_mai_n871_), .B(mai_mai_n582_), .Y(mai_mai_n1206_));
  NO4        m1178(.A(mai_mai_n1206_), .B(mai_mai_n1205_), .C(mai_mai_n1202_), .D(mai_mai_n1193_), .Y(mai_mai_n1207_));
  NO2        m1179(.A(mai_mai_n198_), .B(mai_mai_n554_), .Y(mai_mai_n1208_));
  OAI210     m1180(.A0(mai_mai_n240_), .A1(c), .B0(mai_mai_n578_), .Y(mai_mai_n1209_));
  NA2        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1208_), .Y(mai_mai_n1210_));
  NO3        m1182(.A(mai_mai_n214_), .B(mai_mai_n89_), .C(mai_mai_n247_), .Y(mai_mai_n1211_));
  OAI220     m1183(.A0(mai_mai_n636_), .A1(mai_mai_n218_), .B0(mai_mai_n454_), .B1(mai_mai_n458_), .Y(mai_mai_n1212_));
  NO2        m1184(.A(mai_mai_n1212_), .B(mai_mai_n1211_), .Y(mai_mai_n1213_));
  INV        m1185(.A(mai_mai_n803_), .Y(mai_mai_n1214_));
  NAi31      m1186(.An(mai_mai_n684_), .B(mai_mai_n1214_), .C(mai_mai_n183_), .Y(mai_mai_n1215_));
  NA4        m1187(.A(mai_mai_n1215_), .B(mai_mai_n1213_), .C(mai_mai_n1210_), .D(mai_mai_n1107_), .Y(mai_mai_n1216_));
  NOi31      m1188(.An(mai_mai_n1186_), .B(mai_mai_n415_), .C(mai_mai_n346_), .Y(mai_mai_n1217_));
  OR3        m1189(.A(mai_mai_n1217_), .B(mai_mai_n716_), .C(mai_mai_n483_), .Y(mai_mai_n1218_));
  OR3        m1190(.A(mai_mai_n321_), .B(mai_mai_n198_), .C(mai_mai_n554_), .Y(mai_mai_n1219_));
  INV        m1191(.A(mai_mai_n323_), .Y(mai_mai_n1220_));
  NA3        m1192(.A(mai_mai_n1220_), .B(mai_mai_n1219_), .C(mai_mai_n1218_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n1203_), .B(mai_mai_n693_), .Y(mai_mai_n1222_));
  AN2        m1194(.A(mai_mai_n847_), .B(mai_mai_n846_), .Y(mai_mai_n1223_));
  NO4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n801_), .C(mai_mai_n444_), .D(mai_mai_n430_), .Y(mai_mai_n1224_));
  NA3        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1222_), .C(mai_mai_n1167_), .Y(mai_mai_n1225_));
  NAi21      m1197(.An(j), .B(i), .Y(mai_mai_n1226_));
  NO4        m1198(.A(mai_mai_n1177_), .B(mai_mai_n1226_), .C(mai_mai_n394_), .D(mai_mai_n208_), .Y(mai_mai_n1227_));
  NO4        m1199(.A(mai_mai_n1227_), .B(mai_mai_n1225_), .C(mai_mai_n1221_), .D(mai_mai_n1216_), .Y(mai_mai_n1228_));
  NA4        m1200(.A(mai_mai_n1228_), .B(mai_mai_n1207_), .C(mai_mai_n1189_), .D(mai_mai_n1179_), .Y(mai07));
  NOi21      m1201(.An(j), .B(k), .Y(mai_mai_n1230_));
  NA4        m1202(.A(mai_mai_n158_), .B(mai_mai_n94_), .C(mai_mai_n1230_), .D(f), .Y(mai_mai_n1231_));
  NAi32      m1203(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1232_));
  NO3        m1204(.A(mai_mai_n1232_), .B(m), .C(f), .Y(mai_mai_n1233_));
  OAI210     m1205(.A0(i), .A1(mai_mai_n431_), .B0(mai_mai_n1233_), .Y(mai_mai_n1234_));
  NAi21      m1206(.An(f), .B(c), .Y(mai_mai_n1235_));
  OR2        m1207(.A(e), .B(d), .Y(mai_mai_n1236_));
  OAI220     m1208(.A0(mai_mai_n1236_), .A1(mai_mai_n1235_), .B0(mai_mai_n566_), .B1(mai_mai_n277_), .Y(mai_mai_n1237_));
  NA3        m1209(.A(mai_mai_n1237_), .B(mai_mai_n968_), .C(mai_mai_n158_), .Y(mai_mai_n1238_));
  NOi31      m1210(.An(n), .B(m), .C(b), .Y(mai_mai_n1239_));
  NO3        m1211(.A(mai_mai_n117_), .B(mai_mai_n401_), .C(h), .Y(mai_mai_n1240_));
  NA3        m1212(.A(mai_mai_n1238_), .B(mai_mai_n1234_), .C(mai_mai_n1231_), .Y(mai_mai_n1241_));
  NOi41      m1213(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1242_));
  NO2        m1214(.A(k), .B(i), .Y(mai_mai_n1243_));
  NA3        m1215(.A(mai_mai_n1243_), .B(mai_mai_n821_), .C(mai_mai_n158_), .Y(mai_mai_n1244_));
  NA2        m1216(.A(mai_mai_n76_), .B(mai_mai_n43_), .Y(mai_mai_n1245_));
  NO2        m1217(.A(mai_mai_n962_), .B(mai_mai_n394_), .Y(mai_mai_n1246_));
  NA3        m1218(.A(mai_mai_n1246_), .B(mai_mai_n1245_), .C(mai_mai_n189_), .Y(mai_mai_n1247_));
  NO2        m1219(.A(mai_mai_n976_), .B(mai_mai_n264_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(mai_mai_n484_), .B(mai_mai_n69_), .Y(mai_mai_n1249_));
  NA2        m1221(.A(mai_mai_n1108_), .B(mai_mai_n249_), .Y(mai_mai_n1250_));
  NA4        m1222(.A(mai_mai_n1250_), .B(mai_mai_n1249_), .C(mai_mai_n1247_), .D(mai_mai_n1244_), .Y(mai_mai_n1251_));
  NO2        m1223(.A(mai_mai_n1251_), .B(mai_mai_n1241_), .Y(mai_mai_n1252_));
  NO3        m1224(.A(e), .B(d), .C(c), .Y(mai_mai_n1253_));
  NA2        m1225(.A(mai_mai_n1407_), .B(mai_mai_n1253_), .Y(mai_mai_n1254_));
  NO2        m1226(.A(mai_mai_n1254_), .B(mai_mai_n189_), .Y(mai_mai_n1255_));
  NO3        m1227(.A(n), .B(m), .C(i), .Y(mai_mai_n1256_));
  NA3        m1228(.A(mai_mai_n633_), .B(mai_mai_n620_), .C(mai_mai_n98_), .Y(mai_mai_n1257_));
  NO2        m1229(.A(mai_mai_n1257_), .B(mai_mai_n43_), .Y(mai_mai_n1258_));
  NA2        m1230(.A(mai_mai_n1256_), .B(mai_mai_n577_), .Y(mai_mai_n1259_));
  NO2        m1231(.A(l), .B(k), .Y(mai_mai_n1260_));
  NO3        m1232(.A(mai_mai_n394_), .B(d), .C(c), .Y(mai_mai_n1261_));
  NO2        m1233(.A(mai_mai_n1258_), .B(mai_mai_n1255_), .Y(mai_mai_n1262_));
  NO2        m1234(.A(mai_mai_n986_), .B(l), .Y(mai_mai_n1263_));
  NO2        m1235(.A(m), .B(c), .Y(mai_mai_n1264_));
  NA3        m1236(.A(mai_mai_n1264_), .B(mai_mai_n127_), .C(mai_mai_n166_), .Y(mai_mai_n1265_));
  NO2        m1237(.A(mai_mai_n1265_), .B(mai_mai_n1263_), .Y(mai_mai_n1266_));
  NA2        m1238(.A(mai_mai_n1266_), .B(mai_mai_n158_), .Y(mai_mai_n1267_));
  NO2        m1239(.A(mai_mai_n402_), .B(a), .Y(mai_mai_n1268_));
  NA3        m1240(.A(mai_mai_n1268_), .B(mai_mai_n1408_), .C(mai_mai_n99_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(i), .B(h), .Y(mai_mai_n1270_));
  NA2        m1242(.A(mai_mai_n1041_), .B(h), .Y(mai_mai_n1271_));
  NA2        m1243(.A(mai_mai_n124_), .B(mai_mai_n194_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n1272_), .B(mai_mai_n1271_), .Y(mai_mai_n1273_));
  NO2        m1245(.A(mai_mai_n690_), .B(mai_mai_n167_), .Y(mai_mai_n1274_));
  NOi31      m1246(.An(m), .B(n), .C(b), .Y(mai_mai_n1275_));
  NOi31      m1247(.An(f), .B(d), .C(c), .Y(mai_mai_n1276_));
  NA2        m1248(.A(mai_mai_n1276_), .B(mai_mai_n1275_), .Y(mai_mai_n1277_));
  INV        m1249(.A(mai_mai_n1277_), .Y(mai_mai_n1278_));
  NO3        m1250(.A(mai_mai_n1278_), .B(mai_mai_n1274_), .C(mai_mai_n1273_), .Y(mai_mai_n1279_));
  NA2        m1251(.A(mai_mai_n997_), .B(mai_mai_n418_), .Y(mai_mai_n1280_));
  NO4        m1252(.A(mai_mai_n1280_), .B(mai_mai_n971_), .C(mai_mai_n394_), .D(mai_mai_n43_), .Y(mai_mai_n1281_));
  OAI210     m1253(.A0(mai_mai_n161_), .A1(mai_mai_n469_), .B0(mai_mai_n972_), .Y(mai_mai_n1282_));
  INV        m1254(.A(mai_mai_n1282_), .Y(mai_mai_n1283_));
  NO2        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1281_), .Y(mai_mai_n1284_));
  AN4        m1256(.A(mai_mai_n1284_), .B(mai_mai_n1279_), .C(mai_mai_n1269_), .D(mai_mai_n1267_), .Y(mai_mai_n1285_));
  NA2        m1257(.A(mai_mai_n1239_), .B(mai_mai_n330_), .Y(mai_mai_n1286_));
  NO2        m1258(.A(mai_mai_n1286_), .B(mai_mai_n953_), .Y(mai_mai_n1287_));
  NA2        m1259(.A(mai_mai_n1261_), .B(mai_mai_n190_), .Y(mai_mai_n1288_));
  NO2        m1260(.A(mai_mai_n167_), .B(b), .Y(mai_mai_n1289_));
  AOI220     m1261(.A0(mai_mai_n1072_), .A1(mai_mai_n1289_), .B0(mai_mai_n1005_), .B1(mai_mai_n1280_), .Y(mai_mai_n1290_));
  NAi31      m1262(.An(mai_mai_n1287_), .B(mai_mai_n1290_), .C(mai_mai_n1288_), .Y(mai_mai_n1291_));
  NO4        m1263(.A(mai_mai_n117_), .B(m), .C(f), .D(e), .Y(mai_mai_n1292_));
  NA3        m1264(.A(mai_mai_n1243_), .B(mai_mai_n250_), .C(h), .Y(mai_mai_n1293_));
  OR2        m1265(.A(e), .B(a), .Y(mai_mai_n1294_));
  NO2        m1266(.A(mai_mai_n1236_), .B(mai_mai_n1235_), .Y(mai_mai_n1295_));
  AOI210     m1267(.A0(mai_mai_n29_), .A1(h), .B0(mai_mai_n1295_), .Y(mai_mai_n1296_));
  NO2        m1268(.A(mai_mai_n1296_), .B(mai_mai_n993_), .Y(mai_mai_n1297_));
  NA2        m1269(.A(mai_mai_n1242_), .B(mai_mai_n1260_), .Y(mai_mai_n1298_));
  INV        m1270(.A(mai_mai_n1298_), .Y(mai_mai_n1299_));
  OR3        m1271(.A(mai_mai_n483_), .B(mai_mai_n482_), .C(mai_mai_n98_), .Y(mai_mai_n1300_));
  NA2        m1272(.A(mai_mai_n1022_), .B(mai_mai_n357_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n1301_), .B(mai_mai_n387_), .Y(mai_mai_n1302_));
  AO210      m1274(.A0(mai_mai_n1302_), .A1(mai_mai_n102_), .B0(mai_mai_n1299_), .Y(mai_mai_n1303_));
  NO3        m1275(.A(mai_mai_n1303_), .B(mai_mai_n1297_), .C(mai_mai_n1291_), .Y(mai_mai_n1304_));
  NA4        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1285_), .C(mai_mai_n1262_), .D(mai_mai_n1252_), .Y(mai_mai_n1305_));
  NO2        m1277(.A(mai_mai_n1034_), .B(mai_mai_n96_), .Y(mai_mai_n1306_));
  NA2        m1278(.A(mai_mai_n330_), .B(mai_mai_n51_), .Y(mai_mai_n1307_));
  AOI210     m1279(.A0(mai_mai_n1307_), .A1(mai_mai_n962_), .B0(mai_mai_n1259_), .Y(mai_mai_n1308_));
  NO2        m1280(.A(mai_mai_n998_), .B(mai_mai_n993_), .Y(mai_mai_n1309_));
  NO2        m1281(.A(mai_mai_n1309_), .B(mai_mai_n1308_), .Y(mai_mai_n1310_));
  NO2        m1282(.A(mai_mai_n342_), .B(j), .Y(mai_mai_n1311_));
  NAi41      m1283(.An(mai_mai_n1270_), .B(mai_mai_n984_), .C(mai_mai_n146_), .D(mai_mai_n132_), .Y(mai_mai_n1312_));
  INV        m1284(.A(mai_mai_n1312_), .Y(mai_mai_n1313_));
  NA3        m1285(.A(m), .B(mai_mai_n1311_), .C(mai_mai_n139_), .Y(mai_mai_n1314_));
  INV        m1286(.A(mai_mai_n1314_), .Y(mai_mai_n1315_));
  NO3        m1287(.A(mai_mai_n684_), .B(mai_mai_n153_), .C(mai_mai_n360_), .Y(mai_mai_n1316_));
  NO3        m1288(.A(mai_mai_n1316_), .B(mai_mai_n1315_), .C(mai_mai_n1313_), .Y(mai_mai_n1317_));
  OR2        m1289(.A(n), .B(i), .Y(mai_mai_n1318_));
  OAI210     m1290(.A0(mai_mai_n1318_), .A1(mai_mai_n983_), .B0(mai_mai_n46_), .Y(mai_mai_n1319_));
  AOI220     m1291(.A0(mai_mai_n1319_), .A1(mai_mai_n1079_), .B0(mai_mai_n754_), .B1(mai_mai_n174_), .Y(mai_mai_n1320_));
  INV        m1292(.A(mai_mai_n1320_), .Y(mai_mai_n1321_));
  OAI220     m1293(.A0(mai_mai_n604_), .A1(m), .B0(mai_mai_n198_), .B1(c), .Y(mai_mai_n1322_));
  INV        m1294(.A(mai_mai_n1322_), .Y(mai_mai_n1323_));
  NO2        m1295(.A(mai_mai_n117_), .B(l), .Y(mai_mai_n1324_));
  NO2        m1296(.A(mai_mai_n198_), .B(k), .Y(mai_mai_n1325_));
  OAI210     m1297(.A0(mai_mai_n1325_), .A1(mai_mai_n1270_), .B0(mai_mai_n1324_), .Y(mai_mai_n1326_));
  OAI220     m1298(.A0(mai_mai_n1326_), .A1(mai_mai_n30_), .B0(mai_mai_n1323_), .B1(mai_mai_n155_), .Y(mai_mai_n1327_));
  NO3        m1299(.A(mai_mai_n1300_), .B(mai_mai_n418_), .C(mai_mai_n304_), .Y(mai_mai_n1328_));
  NO3        m1300(.A(mai_mai_n1328_), .B(mai_mai_n1327_), .C(mai_mai_n1321_), .Y(mai_mai_n1329_));
  NO3        m1301(.A(mai_mai_n1008_), .B(mai_mai_n1236_), .C(mai_mai_n46_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n993_), .B(h), .Y(mai_mai_n1331_));
  NA3        m1303(.A(mai_mai_n1331_), .B(d), .C(mai_mai_n954_), .Y(mai_mai_n1332_));
  NO2        m1304(.A(mai_mai_n1332_), .B(c), .Y(mai_mai_n1333_));
  NA3        m1305(.A(mai_mai_n1306_), .B(mai_mai_n418_), .C(f), .Y(mai_mai_n1334_));
  NA2        m1306(.A(mai_mai_n158_), .B(mai_mai_n98_), .Y(mai_mai_n1335_));
  NO2        m1307(.A(mai_mai_n41_), .B(mai_mai_n1334_), .Y(mai_mai_n1336_));
  NOi21      m1308(.An(d), .B(f), .Y(mai_mai_n1337_));
  NO2        m1309(.A(mai_mai_n1336_), .B(mai_mai_n1333_), .Y(mai_mai_n1338_));
  NA4        m1310(.A(mai_mai_n1338_), .B(mai_mai_n1329_), .C(mai_mai_n1317_), .D(mai_mai_n1310_), .Y(mai_mai_n1339_));
  NO3        m1311(.A(mai_mai_n997_), .B(mai_mai_n983_), .C(mai_mai_n39_), .Y(mai_mai_n1340_));
  NA2        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1248_), .Y(mai_mai_n1341_));
  OAI210     m1313(.A0(mai_mai_n1292_), .A1(mai_mai_n1239_), .B0(mai_mai_n808_), .Y(mai_mai_n1342_));
  NO2        m1314(.A(mai_mai_n950_), .B(mai_mai_n117_), .Y(mai_mai_n1343_));
  NA2        m1315(.A(mai_mai_n1343_), .B(mai_mai_n559_), .Y(mai_mai_n1344_));
  NA3        m1316(.A(mai_mai_n1344_), .B(mai_mai_n1342_), .C(mai_mai_n1341_), .Y(mai_mai_n1345_));
  NA2        m1317(.A(mai_mai_n1264_), .B(mai_mai_n1337_), .Y(mai_mai_n1346_));
  NO2        m1318(.A(mai_mai_n1346_), .B(m), .Y(mai_mai_n1347_));
  NO2        m1319(.A(mai_mai_n133_), .B(mai_mai_n160_), .Y(mai_mai_n1348_));
  OAI210     m1320(.A0(mai_mai_n1348_), .A1(mai_mai_n96_), .B0(mai_mai_n1275_), .Y(mai_mai_n1349_));
  INV        m1321(.A(mai_mai_n1349_), .Y(mai_mai_n1350_));
  NO3        m1322(.A(mai_mai_n1350_), .B(mai_mai_n1347_), .C(mai_mai_n1345_), .Y(mai_mai_n1351_));
  NO2        m1323(.A(mai_mai_n1235_), .B(e), .Y(mai_mai_n1352_));
  NA2        m1324(.A(mai_mai_n1352_), .B(mai_mai_n355_), .Y(mai_mai_n1353_));
  NA2        m1325(.A(mai_mai_n1029_), .B(mai_mai_n568_), .Y(mai_mai_n1354_));
  OR3        m1326(.A(mai_mai_n1325_), .B(mai_mai_n1108_), .C(mai_mai_n117_), .Y(mai_mai_n1355_));
  OAI220     m1327(.A0(mai_mai_n1355_), .A1(mai_mai_n1353_), .B0(mai_mai_n1354_), .B1(mai_mai_n396_), .Y(mai_mai_n1356_));
  INV        m1328(.A(mai_mai_n1356_), .Y(mai_mai_n1357_));
  NO2        m1329(.A(mai_mai_n160_), .B(c), .Y(mai_mai_n1358_));
  OAI210     m1330(.A0(mai_mai_n1358_), .A1(mai_mai_n1352_), .B0(mai_mai_n158_), .Y(mai_mai_n1359_));
  AOI220     m1331(.A0(mai_mai_n1359_), .A1(mai_mai_n985_), .B0(mai_mai_n474_), .B1(mai_mai_n318_), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n482_), .B(m), .Y(mai_mai_n1361_));
  AOI210     m1333(.A0(mai_mai_n1361_), .A1(mai_mai_n1261_), .B0(mai_mai_n1330_), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1294_), .B(f), .Y(mai_mai_n1363_));
  AOI210     m1335(.A0(mai_mai_n1029_), .A1(a), .B0(mai_mai_n1363_), .Y(mai_mai_n1364_));
  OAI220     m1336(.A0(mai_mai_n1364_), .A1(mai_mai_n59_), .B0(mai_mai_n1362_), .B1(mai_mai_n188_), .Y(mai_mai_n1365_));
  AOI210     m1337(.A0(mai_mai_n826_), .A1(mai_mai_n367_), .B0(mai_mai_n91_), .Y(mai_mai_n1366_));
  OR2        m1338(.A(mai_mai_n1366_), .B(mai_mai_n482_), .Y(mai_mai_n1367_));
  NA2        m1339(.A(mai_mai_n1363_), .B(mai_mai_n1245_), .Y(mai_mai_n1368_));
  OAI220     m1340(.A0(mai_mai_n1368_), .A1(mai_mai_n46_), .B0(mai_mai_n1367_), .B1(mai_mai_n153_), .Y(mai_mai_n1369_));
  NA4        m1341(.A(mai_mai_n1006_), .B(mai_mai_n1003_), .C(mai_mai_n194_), .D(mai_mai_n58_), .Y(mai_mai_n1370_));
  NA2        m1342(.A(mai_mai_n1240_), .B(mai_mai_n161_), .Y(mai_mai_n1371_));
  NO2        m1343(.A(mai_mai_n46_), .B(l), .Y(mai_mai_n1372_));
  OAI210     m1344(.A0(mai_mai_n1294_), .A1(mai_mai_n789_), .B0(mai_mai_n431_), .Y(mai_mai_n1373_));
  OAI210     m1345(.A0(mai_mai_n1373_), .A1(mai_mai_n1009_), .B0(mai_mai_n1372_), .Y(mai_mai_n1374_));
  NA3        m1346(.A(mai_mai_n1374_), .B(mai_mai_n1371_), .C(mai_mai_n1370_), .Y(mai_mai_n1375_));
  NO4        m1347(.A(mai_mai_n1375_), .B(mai_mai_n1369_), .C(mai_mai_n1365_), .D(mai_mai_n1360_), .Y(mai_mai_n1376_));
  NA3        m1348(.A(mai_mai_n1376_), .B(mai_mai_n1357_), .C(mai_mai_n1351_), .Y(mai_mai_n1377_));
  NA3        m1349(.A(mai_mai_n877_), .B(mai_mai_n124_), .C(mai_mai_n44_), .Y(mai_mai_n1378_));
  AOI210     m1350(.A0(d), .A1(c), .B0(mai_mai_n1378_), .Y(mai_mai_n1379_));
  INV        m1351(.A(mai_mai_n164_), .Y(mai_mai_n1380_));
  NA2        m1352(.A(mai_mai_n1380_), .B(mai_mai_n1331_), .Y(mai_mai_n1381_));
  INV        m1353(.A(mai_mai_n1381_), .Y(mai_mai_n1382_));
  NO2        m1354(.A(mai_mai_n1382_), .B(mai_mai_n1379_), .Y(mai_mai_n1383_));
  AOI210     m1355(.A0(mai_mai_n137_), .A1(mai_mai_n51_), .B0(mai_mai_n1352_), .Y(mai_mai_n1384_));
  NO2        m1356(.A(mai_mai_n1384_), .B(mai_mai_n1335_), .Y(mai_mai_n1385_));
  INV        m1357(.A(mai_mai_n1385_), .Y(mai_mai_n1386_));
  AN2        m1358(.A(mai_mai_n1006_), .B(mai_mai_n991_), .Y(mai_mai_n1387_));
  NA2        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1072_), .Y(mai_mai_n1388_));
  NO2        m1360(.A(mai_mai_n1334_), .B(mai_mai_n59_), .Y(mai_mai_n1389_));
  NA2        m1361(.A(mai_mai_n54_), .B(a), .Y(mai_mai_n1390_));
  NO2        m1362(.A(mai_mai_n1243_), .B(mai_mai_n104_), .Y(mai_mai_n1391_));
  OAI220     m1363(.A0(mai_mai_n1391_), .A1(mai_mai_n1286_), .B0(mai_mai_n1301_), .B1(mai_mai_n1390_), .Y(mai_mai_n1392_));
  NO2        m1364(.A(mai_mai_n1392_), .B(mai_mai_n1389_), .Y(mai_mai_n1393_));
  NA4        m1365(.A(mai_mai_n1393_), .B(mai_mai_n1388_), .C(mai_mai_n1386_), .D(mai_mai_n1383_), .Y(mai_mai_n1394_));
  OR4        m1366(.A(mai_mai_n1394_), .B(mai_mai_n1377_), .C(mai_mai_n1339_), .D(mai_mai_n1305_), .Y(mai04));
  NOi31      m1367(.An(mai_mai_n1292_), .B(mai_mai_n1293_), .C(mai_mai_n956_), .Y(mai_mai_n1396_));
  INV        m1368(.A(mai_mai_n754_), .Y(mai_mai_n1397_));
  NO3        m1369(.A(mai_mai_n1397_), .B(mai_mai_n947_), .C(mai_mai_n432_), .Y(mai_mai_n1398_));
  OR3        m1370(.A(mai_mai_n1398_), .B(mai_mai_n1396_), .C(mai_mai_n974_), .Y(mai_mai_n1399_));
  NO2        m1371(.A(mai_mai_n1245_), .B(mai_mai_n79_), .Y(mai_mai_n1400_));
  AOI210     m1372(.A0(mai_mai_n1400_), .A1(mai_mai_n967_), .B0(mai_mai_n1088_), .Y(mai_mai_n1401_));
  NA2        m1373(.A(mai_mai_n1401_), .B(mai_mai_n1112_), .Y(mai_mai_n1402_));
  NO4        m1374(.A(mai_mai_n1402_), .B(mai_mai_n1399_), .C(mai_mai_n982_), .D(mai_mai_n961_), .Y(mai_mai_n1403_));
  NA4        m1375(.A(mai_mai_n1403_), .B(mai_mai_n1031_), .C(mai_mai_n1020_), .D(mai_mai_n1012_), .Y(mai05));
  INV        m1376(.A(m), .Y(mai_mai_n1407_));
  INV        m1377(.A(i), .Y(mai_mai_n1408_));
  INV        m1378(.A(f), .Y(mai_mai_n1409_));
  INV        m1379(.A(m), .Y(mai_mai_n1410_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(u), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(u), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(u), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(u), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(u), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(u), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  NO2        u0034(.A(men_men_n61_), .B(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(u), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  AN4        u0048(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n77_));
  NOi31      u0049(.An(h), .B(u), .C(f), .Y(men_men_n78_));
  NOi32      u0050(.An(h), .Bn(u), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n74_), .B(men_men_n64_), .Y(men_men_n80_));
  INV        u0052(.A(n), .Y(men_men_n81_));
  NOi32      u0053(.An(e), .Bn(b), .C(d), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n81_), .Y(men_men_n83_));
  INV        u0055(.A(j), .Y(men_men_n84_));
  AN3        u0056(.A(m), .B(k), .C(i), .Y(men_men_n85_));
  NA3        u0057(.A(men_men_n85_), .B(men_men_n84_), .C(u), .Y(men_men_n86_));
  NO2        u0058(.A(men_men_n86_), .B(f), .Y(men_men_n87_));
  NAi32      u0059(.An(u), .Bn(f), .C(h), .Y(men_men_n88_));
  NAi31      u0060(.An(j), .B(m), .C(l), .Y(men_men_n89_));
  NO2        u0061(.A(men_men_n89_), .B(men_men_n88_), .Y(men_men_n90_));
  NA2        u0062(.A(m), .B(l), .Y(men_men_n91_));
  NAi31      u0063(.An(k), .B(j), .C(u), .Y(men_men_n92_));
  NO3        u0064(.A(men_men_n92_), .B(men_men_n91_), .C(f), .Y(men_men_n93_));
  AN2        u0065(.A(j), .B(u), .Y(men_men_n94_));
  NOi32      u0066(.An(m), .Bn(l), .C(i), .Y(men_men_n95_));
  NOi21      u0067(.An(u), .B(i), .Y(men_men_n96_));
  NOi32      u0068(.An(m), .Bn(j), .C(k), .Y(men_men_n97_));
  AOI220     u0069(.A0(men_men_n97_), .A1(men_men_n96_), .B0(men_men_n95_), .B1(men_men_n94_), .Y(men_men_n98_));
  NO2        u0070(.A(men_men_n98_), .B(f), .Y(men_men_n99_));
  NO4        u0071(.A(men_men_n99_), .B(men_men_n93_), .C(men_men_n90_), .D(men_men_n87_), .Y(men_men_n100_));
  NAi41      u0072(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n101_));
  AN2        u0073(.A(e), .B(b), .Y(men_men_n102_));
  NOi31      u0074(.An(c), .B(h), .C(f), .Y(men_men_n103_));
  NA2        u0075(.A(men_men_n103_), .B(men_men_n102_), .Y(men_men_n104_));
  NO2        u0076(.A(men_men_n104_), .B(men_men_n101_), .Y(men_men_n105_));
  NOi21      u0077(.An(u), .B(f), .Y(men_men_n106_));
  NOi21      u0078(.An(i), .B(h), .Y(men_men_n107_));
  NA3        u0079(.A(men_men_n107_), .B(men_men_n106_), .C(men_men_n36_), .Y(men_men_n108_));
  INV        u0080(.A(a), .Y(men_men_n109_));
  NA2        u0081(.A(men_men_n102_), .B(men_men_n109_), .Y(men_men_n110_));
  INV        u0082(.A(l), .Y(men_men_n111_));
  NOi21      u0083(.An(m), .B(n), .Y(men_men_n112_));
  AN2        u0084(.A(k), .B(h), .Y(men_men_n113_));
  NO2        u0085(.A(men_men_n108_), .B(men_men_n83_), .Y(men_men_n114_));
  INV        u0086(.A(b), .Y(men_men_n115_));
  NA2        u0087(.A(l), .B(j), .Y(men_men_n116_));
  AN2        u0088(.A(k), .B(i), .Y(men_men_n117_));
  NA2        u0089(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u0090(.A(u), .B(e), .Y(men_men_n119_));
  NOi32      u0091(.An(c), .Bn(a), .C(d), .Y(men_men_n120_));
  NA2        u0092(.A(men_men_n120_), .B(men_men_n112_), .Y(men_men_n121_));
  NO4        u0093(.A(men_men_n121_), .B(men_men_n119_), .C(men_men_n118_), .D(men_men_n115_), .Y(men_men_n122_));
  NO3        u0094(.A(men_men_n122_), .B(men_men_n114_), .C(men_men_n105_), .Y(men_men_n123_));
  OAI210     u0095(.A0(men_men_n100_), .A1(men_men_n83_), .B0(men_men_n123_), .Y(men_men_n124_));
  NOi31      u0096(.An(k), .B(m), .C(j), .Y(men_men_n125_));
  NA3        u0097(.A(men_men_n125_), .B(men_men_n78_), .C(men_men_n77_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(i), .Y(men_men_n127_));
  NA3        u0099(.A(men_men_n127_), .B(men_men_n79_), .C(men_men_n77_), .Y(men_men_n128_));
  NA2        u0100(.A(men_men_n128_), .B(men_men_n126_), .Y(men_men_n129_));
  NOi32      u0101(.An(f), .Bn(b), .C(e), .Y(men_men_n130_));
  NAi21      u0102(.An(u), .B(h), .Y(men_men_n131_));
  NAi21      u0103(.An(m), .B(n), .Y(men_men_n132_));
  NAi21      u0104(.An(j), .B(k), .Y(men_men_n133_));
  NO3        u0105(.A(men_men_n133_), .B(men_men_n132_), .C(men_men_n131_), .Y(men_men_n134_));
  NAi41      u0106(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n135_));
  NAi31      u0107(.An(j), .B(k), .C(h), .Y(men_men_n136_));
  NO3        u0108(.A(men_men_n136_), .B(men_men_n135_), .C(men_men_n132_), .Y(men_men_n137_));
  AOI210     u0109(.A0(men_men_n134_), .A1(men_men_n130_), .B0(men_men_n137_), .Y(men_men_n138_));
  NO2        u0110(.A(k), .B(j), .Y(men_men_n139_));
  NO2        u0111(.A(men_men_n139_), .B(men_men_n132_), .Y(men_men_n140_));
  AN2        u0112(.A(k), .B(j), .Y(men_men_n141_));
  NAi21      u0113(.An(c), .B(b), .Y(men_men_n142_));
  NA2        u0114(.A(f), .B(d), .Y(men_men_n143_));
  NO3        u0115(.A(men_men_n143_), .B(men_men_n142_), .C(men_men_n131_), .Y(men_men_n144_));
  NAi31      u0116(.An(f), .B(e), .C(b), .Y(men_men_n145_));
  NA2        u0117(.A(men_men_n144_), .B(men_men_n140_), .Y(men_men_n146_));
  NA2        u0118(.A(d), .B(b), .Y(men_men_n147_));
  NAi21      u0119(.An(e), .B(f), .Y(men_men_n148_));
  NO2        u0120(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n149_));
  NA2        u0121(.A(b), .B(a), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(u), .Y(men_men_n151_));
  NAi21      u0123(.An(c), .B(d), .Y(men_men_n152_));
  NAi31      u0124(.An(l), .B(k), .C(h), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n132_), .B(men_men_n153_), .Y(men_men_n154_));
  NA2        u0126(.A(men_men_n154_), .B(men_men_n149_), .Y(men_men_n155_));
  NAi41      u0127(.An(men_men_n129_), .B(men_men_n155_), .C(men_men_n146_), .D(men_men_n138_), .Y(men_men_n156_));
  NAi31      u0128(.An(e), .B(f), .C(b), .Y(men_men_n157_));
  NOi21      u0129(.An(u), .B(d), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NOi21      u0131(.An(h), .B(i), .Y(men_men_n160_));
  NOi21      u0132(.An(k), .B(m), .Y(men_men_n161_));
  NA3        u0133(.A(men_men_n161_), .B(men_men_n160_), .C(n), .Y(men_men_n162_));
  NOi21      u0134(.An(men_men_n159_), .B(men_men_n162_), .Y(men_men_n163_));
  NOi21      u0135(.An(h), .B(u), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n143_), .B(men_men_n142_), .Y(men_men_n165_));
  NAi31      u0137(.An(l), .B(j), .C(h), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n166_), .B(men_men_n49_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n67_), .Y(men_men_n168_));
  NOi32      u0140(.An(n), .Bn(k), .C(m), .Y(men_men_n169_));
  NA2        u0141(.A(l), .B(i), .Y(men_men_n170_));
  INV        u0142(.A(men_men_n168_), .Y(men_men_n171_));
  NAi31      u0143(.An(d), .B(f), .C(c), .Y(men_men_n172_));
  NAi31      u0144(.An(e), .B(f), .C(c), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NA2        u0146(.A(j), .B(h), .Y(men_men_n175_));
  OR3        u0147(.A(n), .B(m), .C(k), .Y(men_men_n176_));
  NO2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  NAi32      u0149(.An(m), .Bn(k), .C(n), .Y(men_men_n178_));
  NO2        u0150(.A(men_men_n178_), .B(men_men_n175_), .Y(men_men_n179_));
  AOI220     u0151(.A0(men_men_n179_), .A1(men_men_n159_), .B0(men_men_n177_), .B1(men_men_n174_), .Y(men_men_n180_));
  NO2        u0152(.A(n), .B(m), .Y(men_men_n181_));
  NA2        u0153(.A(men_men_n181_), .B(men_men_n50_), .Y(men_men_n182_));
  NAi21      u0154(.An(f), .B(e), .Y(men_men_n183_));
  NA2        u0155(.A(d), .B(c), .Y(men_men_n184_));
  NAi31      u0156(.An(m), .B(n), .C(b), .Y(men_men_n185_));
  NA2        u0157(.A(k), .B(i), .Y(men_men_n186_));
  NAi21      u0158(.An(h), .B(f), .Y(men_men_n187_));
  NO2        u0159(.A(men_men_n187_), .B(men_men_n186_), .Y(men_men_n188_));
  NO2        u0160(.A(men_men_n185_), .B(men_men_n152_), .Y(men_men_n189_));
  NA2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NOi32      u0162(.An(f), .Bn(c), .C(d), .Y(men_men_n191_));
  NOi32      u0163(.An(f), .Bn(c), .C(e), .Y(men_men_n192_));
  NO2        u0164(.A(men_men_n192_), .B(men_men_n191_), .Y(men_men_n193_));
  NO3        u0165(.A(n), .B(m), .C(j), .Y(men_men_n194_));
  NA2        u0166(.A(men_men_n194_), .B(men_men_n113_), .Y(men_men_n195_));
  AO210      u0167(.A0(men_men_n195_), .A1(men_men_n182_), .B0(men_men_n193_), .Y(men_men_n196_));
  NA3        u0168(.A(men_men_n196_), .B(men_men_n190_), .C(men_men_n180_), .Y(men_men_n197_));
  OR4        u0169(.A(men_men_n197_), .B(men_men_n171_), .C(men_men_n163_), .D(men_men_n156_), .Y(men_men_n198_));
  NO4        u0170(.A(men_men_n198_), .B(men_men_n124_), .C(men_men_n80_), .D(men_men_n55_), .Y(men_men_n199_));
  NA3        u0171(.A(m), .B(men_men_n111_), .C(j), .Y(men_men_n200_));
  NAi31      u0172(.An(n), .B(h), .C(u), .Y(men_men_n201_));
  NO2        u0173(.A(men_men_n201_), .B(men_men_n200_), .Y(men_men_n202_));
  NOi32      u0174(.An(m), .Bn(k), .C(l), .Y(men_men_n203_));
  NA3        u0175(.A(men_men_n203_), .B(men_men_n84_), .C(u), .Y(men_men_n204_));
  NO2        u0176(.A(men_men_n204_), .B(n), .Y(men_men_n205_));
  NOi21      u0177(.An(k), .B(j), .Y(men_men_n206_));
  NA4        u0178(.A(men_men_n206_), .B(men_men_n112_), .C(i), .D(u), .Y(men_men_n207_));
  AN2        u0179(.A(i), .B(u), .Y(men_men_n208_));
  NA3        u0180(.A(men_men_n76_), .B(men_men_n208_), .C(men_men_n112_), .Y(men_men_n209_));
  NA2        u0181(.A(men_men_n209_), .B(men_men_n207_), .Y(men_men_n210_));
  NO3        u0182(.A(men_men_n210_), .B(men_men_n205_), .C(men_men_n202_), .Y(men_men_n211_));
  NAi41      u0183(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n212_));
  INV        u0184(.A(men_men_n212_), .Y(men_men_n213_));
  INV        u0185(.A(f), .Y(men_men_n214_));
  INV        u0186(.A(u), .Y(men_men_n215_));
  NOi31      u0187(.An(i), .B(j), .C(h), .Y(men_men_n216_));
  NOi21      u0188(.An(l), .B(m), .Y(men_men_n217_));
  NA2        u0189(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  NO3        u0190(.A(men_men_n218_), .B(men_men_n215_), .C(men_men_n214_), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n213_), .Y(men_men_n220_));
  OAI210     u0192(.A0(men_men_n211_), .A1(men_men_n32_), .B0(men_men_n220_), .Y(men_men_n221_));
  NOi21      u0193(.An(n), .B(m), .Y(men_men_n222_));
  NOi32      u0194(.An(l), .Bn(i), .C(j), .Y(men_men_n223_));
  NA2        u0195(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  OR2        u0196(.A(men_men_n224_), .B(men_men_n104_), .Y(men_men_n225_));
  NAi21      u0197(.An(j), .B(h), .Y(men_men_n226_));
  XN2        u0198(.A(i), .B(h), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  NOi31      u0200(.An(k), .B(n), .C(m), .Y(men_men_n229_));
  NOi31      u0201(.An(men_men_n229_), .B(men_men_n184_), .C(men_men_n183_), .Y(men_men_n230_));
  NA2        u0202(.A(men_men_n230_), .B(men_men_n228_), .Y(men_men_n231_));
  NAi31      u0203(.An(f), .B(e), .C(c), .Y(men_men_n232_));
  NO4        u0204(.A(men_men_n232_), .B(men_men_n176_), .C(men_men_n175_), .D(men_men_n59_), .Y(men_men_n233_));
  NA4        u0205(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n234_));
  NAi32      u0206(.An(m), .Bn(i), .C(k), .Y(men_men_n235_));
  NO3        u0207(.A(men_men_n235_), .B(men_men_n88_), .C(men_men_n234_), .Y(men_men_n236_));
  INV        u0208(.A(k), .Y(men_men_n237_));
  NO2        u0209(.A(men_men_n236_), .B(men_men_n233_), .Y(men_men_n238_));
  NAi21      u0210(.An(n), .B(a), .Y(men_men_n239_));
  NO2        u0211(.A(men_men_n239_), .B(men_men_n147_), .Y(men_men_n240_));
  NAi41      u0212(.An(u), .B(m), .C(k), .D(h), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(e), .Y(men_men_n242_));
  NO3        u0214(.A(men_men_n148_), .B(men_men_n92_), .C(men_men_n91_), .Y(men_men_n243_));
  OAI210     u0215(.A0(men_men_n243_), .A1(men_men_n242_), .B0(men_men_n240_), .Y(men_men_n244_));
  AN4        u0216(.A(men_men_n244_), .B(men_men_n238_), .C(men_men_n231_), .D(men_men_n225_), .Y(men_men_n245_));
  OR2        u0217(.A(h), .B(u), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(men_men_n101_), .Y(men_men_n247_));
  NAi41      u0219(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n248_), .B(men_men_n214_), .Y(men_men_n249_));
  NA2        u0221(.A(men_men_n161_), .B(men_men_n107_), .Y(men_men_n250_));
  NAi21      u0222(.An(men_men_n250_), .B(men_men_n249_), .Y(men_men_n251_));
  NO2        u0223(.A(n), .B(a), .Y(men_men_n252_));
  NAi31      u0224(.An(men_men_n241_), .B(men_men_n252_), .C(men_men_n102_), .Y(men_men_n253_));
  AN2        u0225(.A(men_men_n253_), .B(men_men_n251_), .Y(men_men_n254_));
  NAi21      u0226(.An(h), .B(i), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n181_), .B(k), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  NA2        u0229(.A(men_men_n257_), .B(men_men_n191_), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n258_), .B(men_men_n254_), .Y(men_men_n259_));
  NOi21      u0231(.An(u), .B(e), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n261_));
  NOi32      u0233(.An(l), .Bn(j), .C(i), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n255_), .B(men_men_n44_), .Y(men_men_n263_));
  NAi21      u0235(.An(f), .B(u), .Y(men_men_n264_));
  NO2        u0236(.A(men_men_n264_), .B(men_men_n65_), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n69_), .B(men_men_n116_), .Y(men_men_n266_));
  AOI220     u0238(.A0(men_men_n266_), .A1(men_men_n265_), .B0(men_men_n263_), .B1(men_men_n67_), .Y(men_men_n267_));
  INV        u0239(.A(men_men_n267_), .Y(men_men_n268_));
  NO3        u0240(.A(men_men_n133_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n269_));
  NOi41      u0241(.An(men_men_n245_), .B(men_men_n268_), .C(men_men_n259_), .D(men_men_n221_), .Y(men_men_n270_));
  NO4        u0242(.A(men_men_n202_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n271_));
  NO2        u0243(.A(men_men_n271_), .B(men_men_n110_), .Y(men_men_n272_));
  NAi21      u0244(.An(h), .B(u), .Y(men_men_n273_));
  OR4        u0245(.A(men_men_n273_), .B(men_men_n1498_), .C(men_men_n224_), .D(e), .Y(men_men_n274_));
  NAi31      u0246(.An(u), .B(k), .C(h), .Y(men_men_n275_));
  NO3        u0247(.A(men_men_n132_), .B(men_men_n275_), .C(l), .Y(men_men_n276_));
  NAi31      u0248(.An(e), .B(d), .C(a), .Y(men_men_n277_));
  NA2        u0249(.A(men_men_n276_), .B(men_men_n130_), .Y(men_men_n278_));
  NA2        u0250(.A(men_men_n278_), .B(men_men_n274_), .Y(men_men_n279_));
  NA3        u0251(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n81_), .Y(men_men_n280_));
  NO2        u0252(.A(men_men_n280_), .B(men_men_n193_), .Y(men_men_n281_));
  INV        u0253(.A(men_men_n281_), .Y(men_men_n282_));
  NA3        u0254(.A(e), .B(c), .C(b), .Y(men_men_n283_));
  NO2        u0255(.A(men_men_n60_), .B(men_men_n283_), .Y(men_men_n284_));
  NAi32      u0256(.An(k), .Bn(i), .C(j), .Y(men_men_n285_));
  NAi31      u0257(.An(h), .B(l), .C(i), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n286_), .B(men_men_n285_), .C(men_men_n166_), .Y(men_men_n287_));
  NOi21      u0259(.An(men_men_n287_), .B(men_men_n49_), .Y(men_men_n288_));
  OAI210     u0260(.A0(men_men_n265_), .A1(men_men_n284_), .B0(men_men_n288_), .Y(men_men_n289_));
  NAi21      u0261(.An(l), .B(k), .Y(men_men_n290_));
  NO2        u0262(.A(men_men_n290_), .B(men_men_n49_), .Y(men_men_n291_));
  NOi21      u0263(.An(l), .B(j), .Y(men_men_n292_));
  NA2        u0264(.A(men_men_n164_), .B(men_men_n292_), .Y(men_men_n293_));
  NA3        u0265(.A(men_men_n117_), .B(men_men_n116_), .C(u), .Y(men_men_n294_));
  OR3        u0266(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n295_));
  AOI210     u0267(.A0(men_men_n294_), .A1(men_men_n293_), .B0(men_men_n295_), .Y(men_men_n296_));
  INV        u0268(.A(men_men_n296_), .Y(men_men_n297_));
  NAi32      u0269(.An(j), .Bn(h), .C(i), .Y(men_men_n298_));
  NAi21      u0270(.An(m), .B(l), .Y(men_men_n299_));
  NO3        u0271(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n81_), .Y(men_men_n300_));
  NA2        u0272(.A(h), .B(u), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n169_), .B(men_men_n45_), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n302_), .B(men_men_n301_), .Y(men_men_n303_));
  OAI210     u0275(.A0(men_men_n303_), .A1(men_men_n300_), .B0(men_men_n165_), .Y(men_men_n304_));
  NA4        u0276(.A(men_men_n304_), .B(men_men_n297_), .C(men_men_n289_), .D(men_men_n282_), .Y(men_men_n305_));
  NO2        u0277(.A(men_men_n145_), .B(d), .Y(men_men_n306_));
  NA2        u0278(.A(men_men_n306_), .B(men_men_n53_), .Y(men_men_n307_));
  NO2        u0279(.A(men_men_n104_), .B(men_men_n101_), .Y(men_men_n308_));
  NAi32      u0280(.An(n), .Bn(m), .C(l), .Y(men_men_n309_));
  NO2        u0281(.A(men_men_n121_), .B(men_men_n115_), .Y(men_men_n310_));
  NAi31      u0282(.An(k), .B(l), .C(j), .Y(men_men_n311_));
  OAI210     u0283(.A0(men_men_n290_), .A1(j), .B0(men_men_n311_), .Y(men_men_n312_));
  NOi21      u0284(.An(men_men_n312_), .B(men_men_n119_), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n310_), .Y(men_men_n314_));
  NA2        u0286(.A(men_men_n314_), .B(men_men_n307_), .Y(men_men_n315_));
  NO4        u0287(.A(men_men_n315_), .B(men_men_n305_), .C(men_men_n279_), .D(men_men_n272_), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n257_), .B(men_men_n192_), .Y(men_men_n317_));
  NAi21      u0289(.An(m), .B(k), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n227_), .B(men_men_n318_), .Y(men_men_n319_));
  NAi41      u0291(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n151_), .Y(men_men_n321_));
  NA2        u0293(.A(men_men_n321_), .B(men_men_n319_), .Y(men_men_n322_));
  NAi31      u0294(.An(i), .B(l), .C(h), .Y(men_men_n323_));
  NO4        u0295(.A(men_men_n323_), .B(men_men_n151_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n324_));
  NA2        u0296(.A(e), .B(c), .Y(men_men_n325_));
  NO3        u0297(.A(men_men_n325_), .B(n), .C(d), .Y(men_men_n326_));
  NOi21      u0298(.An(f), .B(h), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n327_), .B(men_men_n117_), .Y(men_men_n328_));
  NO2        u0300(.A(men_men_n328_), .B(men_men_n215_), .Y(men_men_n329_));
  NAi31      u0301(.An(d), .B(e), .C(b), .Y(men_men_n330_));
  NO2        u0302(.A(men_men_n132_), .B(men_men_n330_), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n331_), .B(men_men_n329_), .Y(men_men_n332_));
  NAi41      u0304(.An(men_men_n324_), .B(men_men_n332_), .C(men_men_n322_), .D(men_men_n317_), .Y(men_men_n333_));
  NA2        u0305(.A(men_men_n252_), .B(men_men_n102_), .Y(men_men_n334_));
  OR2        u0306(.A(men_men_n334_), .B(men_men_n204_), .Y(men_men_n335_));
  NOi31      u0307(.An(l), .B(n), .C(m), .Y(men_men_n336_));
  INV        u0308(.A(men_men_n335_), .Y(men_men_n337_));
  NAi32      u0309(.An(m), .Bn(j), .C(k), .Y(men_men_n338_));
  NAi41      u0310(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n339_));
  NA2        u0311(.A(men_men_n212_), .B(men_men_n339_), .Y(men_men_n340_));
  NOi31      u0312(.An(j), .B(m), .C(k), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n125_), .B(men_men_n341_), .Y(men_men_n342_));
  AN3        u0314(.A(h), .B(u), .C(f), .Y(men_men_n343_));
  NAi31      u0315(.An(men_men_n342_), .B(men_men_n343_), .C(men_men_n340_), .Y(men_men_n344_));
  NOi32      u0316(.An(m), .Bn(j), .C(l), .Y(men_men_n345_));
  NO2        u0317(.A(men_men_n345_), .B(men_men_n95_), .Y(men_men_n346_));
  NAi32      u0318(.An(men_men_n346_), .Bn(men_men_n201_), .C(men_men_n306_), .Y(men_men_n347_));
  NO2        u0319(.A(men_men_n299_), .B(men_men_n298_), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n218_), .B(u), .Y(men_men_n349_));
  NO2        u0321(.A(men_men_n157_), .B(men_men_n81_), .Y(men_men_n350_));
  AOI220     u0322(.A0(men_men_n350_), .A1(men_men_n349_), .B0(men_men_n249_), .B1(men_men_n348_), .Y(men_men_n351_));
  INV        u0323(.A(men_men_n235_), .Y(men_men_n352_));
  NA3        u0324(.A(men_men_n352_), .B(men_men_n343_), .C(men_men_n213_), .Y(men_men_n353_));
  NA4        u0325(.A(men_men_n353_), .B(men_men_n351_), .C(men_men_n347_), .D(men_men_n344_), .Y(men_men_n354_));
  NA3        u0326(.A(h), .B(u), .C(f), .Y(men_men_n355_));
  NA2        u0327(.A(men_men_n164_), .B(e), .Y(men_men_n356_));
  NOi32      u0328(.An(j), .Bn(u), .C(i), .Y(men_men_n357_));
  NA3        u0329(.A(men_men_n357_), .B(men_men_n290_), .C(men_men_n112_), .Y(men_men_n358_));
  AO210      u0330(.A0(men_men_n110_), .A1(men_men_n32_), .B0(men_men_n358_), .Y(men_men_n359_));
  NOi32      u0331(.An(e), .Bn(b), .C(a), .Y(men_men_n360_));
  AN2        u0332(.A(l), .B(j), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n318_), .B(men_men_n361_), .Y(men_men_n362_));
  NO3        u0334(.A(men_men_n320_), .B(men_men_n72_), .C(men_men_n215_), .Y(men_men_n363_));
  NA3        u0335(.A(men_men_n209_), .B(men_men_n207_), .C(men_men_n35_), .Y(men_men_n364_));
  AOI220     u0336(.A0(men_men_n364_), .A1(men_men_n360_), .B0(men_men_n363_), .B1(men_men_n362_), .Y(men_men_n365_));
  NO2        u0337(.A(men_men_n330_), .B(n), .Y(men_men_n366_));
  NA2        u0338(.A(men_men_n208_), .B(k), .Y(men_men_n367_));
  NA3        u0339(.A(m), .B(men_men_n111_), .C(men_men_n214_), .Y(men_men_n368_));
  NA4        u0340(.A(men_men_n203_), .B(men_men_n84_), .C(u), .D(men_men_n214_), .Y(men_men_n369_));
  OAI210     u0341(.A0(men_men_n368_), .A1(men_men_n367_), .B0(men_men_n369_), .Y(men_men_n370_));
  NAi41      u0342(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n371_));
  NA2        u0343(.A(men_men_n51_), .B(men_men_n112_), .Y(men_men_n372_));
  NO2        u0344(.A(men_men_n372_), .B(men_men_n371_), .Y(men_men_n373_));
  AOI220     u0345(.A0(men_men_n373_), .A1(b), .B0(men_men_n370_), .B1(men_men_n366_), .Y(men_men_n374_));
  NA3        u0346(.A(men_men_n374_), .B(men_men_n365_), .C(men_men_n359_), .Y(men_men_n375_));
  NO4        u0347(.A(men_men_n375_), .B(men_men_n354_), .C(men_men_n337_), .D(men_men_n333_), .Y(men_men_n376_));
  NA4        u0348(.A(men_men_n376_), .B(men_men_n316_), .C(men_men_n270_), .D(men_men_n199_), .Y(men10));
  NA3        u0349(.A(m), .B(k), .C(i), .Y(men_men_n378_));
  NO3        u0350(.A(men_men_n378_), .B(j), .C(men_men_n215_), .Y(men_men_n379_));
  NOi21      u0351(.An(e), .B(f), .Y(men_men_n380_));
  NO4        u0352(.A(men_men_n152_), .B(men_men_n380_), .C(n), .D(men_men_n109_), .Y(men_men_n381_));
  NAi31      u0353(.An(b), .B(f), .C(c), .Y(men_men_n382_));
  INV        u0354(.A(men_men_n382_), .Y(men_men_n383_));
  NOi32      u0355(.An(k), .Bn(h), .C(j), .Y(men_men_n384_));
  NA2        u0356(.A(men_men_n384_), .B(men_men_n222_), .Y(men_men_n385_));
  NA2        u0357(.A(men_men_n162_), .B(men_men_n385_), .Y(men_men_n386_));
  AOI220     u0358(.A0(men_men_n386_), .A1(men_men_n383_), .B0(men_men_n381_), .B1(men_men_n379_), .Y(men_men_n387_));
  AN2        u0359(.A(j), .B(h), .Y(men_men_n388_));
  NO3        u0360(.A(n), .B(m), .C(k), .Y(men_men_n389_));
  NA2        u0361(.A(men_men_n389_), .B(men_men_n388_), .Y(men_men_n390_));
  NO3        u0362(.A(men_men_n390_), .B(men_men_n152_), .C(men_men_n214_), .Y(men_men_n391_));
  OR2        u0363(.A(m), .B(k), .Y(men_men_n392_));
  NO2        u0364(.A(men_men_n175_), .B(men_men_n392_), .Y(men_men_n393_));
  NA4        u0365(.A(n), .B(f), .C(c), .D(men_men_n115_), .Y(men_men_n394_));
  NOi21      u0366(.An(men_men_n393_), .B(men_men_n394_), .Y(men_men_n395_));
  NOi32      u0367(.An(d), .Bn(a), .C(c), .Y(men_men_n396_));
  NA2        u0368(.A(men_men_n396_), .B(men_men_n183_), .Y(men_men_n397_));
  NAi21      u0369(.An(i), .B(u), .Y(men_men_n398_));
  NAi31      u0370(.An(k), .B(m), .C(j), .Y(men_men_n399_));
  NO3        u0371(.A(men_men_n399_), .B(men_men_n398_), .C(n), .Y(men_men_n400_));
  NOi21      u0372(.An(men_men_n400_), .B(men_men_n397_), .Y(men_men_n401_));
  NO3        u0373(.A(men_men_n401_), .B(men_men_n395_), .C(men_men_n391_), .Y(men_men_n402_));
  NO2        u0374(.A(men_men_n394_), .B(men_men_n299_), .Y(men_men_n403_));
  NOi32      u0375(.An(f), .Bn(d), .C(c), .Y(men_men_n404_));
  NA2        u0376(.A(men_men_n402_), .B(men_men_n387_), .Y(men_men_n405_));
  NO2        u0377(.A(men_men_n59_), .B(men_men_n115_), .Y(men_men_n406_));
  NA2        u0378(.A(men_men_n252_), .B(men_men_n406_), .Y(men_men_n407_));
  INV        u0379(.A(e), .Y(men_men_n408_));
  NA2        u0380(.A(men_men_n46_), .B(e), .Y(men_men_n409_));
  OAI220     u0381(.A0(men_men_n409_), .A1(men_men_n200_), .B0(men_men_n204_), .B1(men_men_n408_), .Y(men_men_n410_));
  AN2        u0382(.A(u), .B(e), .Y(men_men_n411_));
  NA3        u0383(.A(men_men_n411_), .B(men_men_n203_), .C(i), .Y(men_men_n412_));
  OAI210     u0384(.A0(men_men_n86_), .A1(men_men_n408_), .B0(men_men_n412_), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n98_), .B(men_men_n408_), .Y(men_men_n414_));
  NO3        u0386(.A(men_men_n414_), .B(men_men_n413_), .C(men_men_n410_), .Y(men_men_n415_));
  NOi32      u0387(.An(h), .Bn(e), .C(u), .Y(men_men_n416_));
  NA3        u0388(.A(men_men_n416_), .B(men_men_n292_), .C(m), .Y(men_men_n417_));
  NOi21      u0389(.An(u), .B(h), .Y(men_men_n418_));
  AN3        u0390(.A(m), .B(l), .C(i), .Y(men_men_n419_));
  NA3        u0391(.A(men_men_n419_), .B(men_men_n418_), .C(e), .Y(men_men_n420_));
  AN3        u0392(.A(h), .B(u), .C(e), .Y(men_men_n421_));
  NA2        u0393(.A(men_men_n421_), .B(men_men_n95_), .Y(men_men_n422_));
  AN3        u0394(.A(men_men_n422_), .B(men_men_n420_), .C(men_men_n417_), .Y(men_men_n423_));
  AOI210     u0395(.A0(men_men_n423_), .A1(men_men_n415_), .B0(men_men_n407_), .Y(men_men_n424_));
  NA3        u0396(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n425_));
  NA3        u0397(.A(men_men_n396_), .B(men_men_n183_), .C(men_men_n81_), .Y(men_men_n426_));
  NAi31      u0398(.An(b), .B(c), .C(a), .Y(men_men_n427_));
  NO2        u0399(.A(men_men_n427_), .B(n), .Y(men_men_n428_));
  OAI210     u0400(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n429_), .B(men_men_n148_), .Y(men_men_n430_));
  NA2        u0402(.A(men_men_n430_), .B(men_men_n428_), .Y(men_men_n431_));
  INV        u0403(.A(men_men_n431_), .Y(men_men_n432_));
  NO3        u0404(.A(men_men_n432_), .B(men_men_n424_), .C(men_men_n405_), .Y(men_men_n433_));
  NA2        u0405(.A(i), .B(u), .Y(men_men_n434_));
  NO3        u0406(.A(men_men_n277_), .B(men_men_n434_), .C(c), .Y(men_men_n435_));
  NOi21      u0407(.An(a), .B(n), .Y(men_men_n436_));
  NOi21      u0408(.An(d), .B(c), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n437_), .B(men_men_n436_), .Y(men_men_n438_));
  NA3        u0410(.A(i), .B(u), .C(f), .Y(men_men_n439_));
  OR2        u0411(.A(men_men_n439_), .B(men_men_n71_), .Y(men_men_n440_));
  NA2        u0412(.A(men_men_n435_), .B(men_men_n291_), .Y(men_men_n441_));
  OR2        u0413(.A(n), .B(m), .Y(men_men_n442_));
  NO2        u0414(.A(men_men_n442_), .B(men_men_n153_), .Y(men_men_n443_));
  NO2        u0415(.A(men_men_n184_), .B(men_men_n148_), .Y(men_men_n444_));
  OAI210     u0416(.A0(men_men_n443_), .A1(men_men_n177_), .B0(men_men_n444_), .Y(men_men_n445_));
  INV        u0417(.A(men_men_n372_), .Y(men_men_n446_));
  NA3        u0418(.A(men_men_n446_), .B(men_men_n360_), .C(d), .Y(men_men_n447_));
  NO2        u0419(.A(men_men_n427_), .B(men_men_n49_), .Y(men_men_n448_));
  NO3        u0420(.A(men_men_n66_), .B(men_men_n111_), .C(e), .Y(men_men_n449_));
  NAi21      u0421(.An(k), .B(j), .Y(men_men_n450_));
  NA3        u0422(.A(i), .B(men_men_n449_), .C(men_men_n448_), .Y(men_men_n451_));
  NAi21      u0423(.An(e), .B(d), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n452_), .Y(men_men_n453_));
  NO2        u0425(.A(men_men_n256_), .B(men_men_n214_), .Y(men_men_n454_));
  NA3        u0426(.A(men_men_n454_), .B(men_men_n453_), .C(men_men_n228_), .Y(men_men_n455_));
  NA4        u0427(.A(men_men_n455_), .B(men_men_n451_), .C(men_men_n447_), .D(men_men_n445_), .Y(men_men_n456_));
  NOi31      u0428(.An(n), .B(m), .C(k), .Y(men_men_n457_));
  AOI220     u0429(.A0(men_men_n457_), .A1(men_men_n388_), .B0(men_men_n222_), .B1(men_men_n50_), .Y(men_men_n458_));
  NAi31      u0430(.An(u), .B(f), .C(c), .Y(men_men_n459_));
  NOi31      u0431(.An(men_men_n441_), .B(men_men_n456_), .C(men_men_n268_), .Y(men_men_n460_));
  NOi32      u0432(.An(c), .Bn(a), .C(b), .Y(men_men_n461_));
  NA2        u0433(.A(men_men_n461_), .B(men_men_n112_), .Y(men_men_n462_));
  INV        u0434(.A(men_men_n275_), .Y(men_men_n463_));
  AN2        u0435(.A(e), .B(d), .Y(men_men_n464_));
  NA2        u0436(.A(men_men_n464_), .B(men_men_n463_), .Y(men_men_n465_));
  NO2        u0437(.A(men_men_n131_), .B(men_men_n41_), .Y(men_men_n466_));
  NO2        u0438(.A(men_men_n66_), .B(e), .Y(men_men_n467_));
  NOi31      u0439(.An(j), .B(k), .C(i), .Y(men_men_n468_));
  NOi21      u0440(.An(men_men_n166_), .B(men_men_n468_), .Y(men_men_n469_));
  NA2        u0441(.A(men_men_n323_), .B(men_men_n469_), .Y(men_men_n470_));
  NA2        u0442(.A(men_men_n470_), .B(men_men_n467_), .Y(men_men_n471_));
  AOI210     u0443(.A0(men_men_n471_), .A1(men_men_n465_), .B0(men_men_n462_), .Y(men_men_n472_));
  NO2        u0444(.A(men_men_n210_), .B(men_men_n205_), .Y(men_men_n473_));
  NOi21      u0445(.An(a), .B(b), .Y(men_men_n474_));
  NA3        u0446(.A(e), .B(d), .C(c), .Y(men_men_n475_));
  NAi21      u0447(.An(men_men_n475_), .B(men_men_n474_), .Y(men_men_n476_));
  AOI210     u0448(.A0(men_men_n271_), .A1(men_men_n473_), .B0(men_men_n476_), .Y(men_men_n477_));
  NO4        u0449(.A(men_men_n187_), .B(men_men_n101_), .C(men_men_n56_), .D(b), .Y(men_men_n478_));
  NA2        u0450(.A(men_men_n383_), .B(men_men_n154_), .Y(men_men_n479_));
  OR2        u0451(.A(k), .B(j), .Y(men_men_n480_));
  NA2        u0452(.A(l), .B(k), .Y(men_men_n481_));
  NA3        u0453(.A(men_men_n481_), .B(men_men_n480_), .C(men_men_n222_), .Y(men_men_n482_));
  AOI210     u0454(.A0(men_men_n235_), .A1(men_men_n338_), .B0(men_men_n81_), .Y(men_men_n483_));
  NOi21      u0455(.An(men_men_n482_), .B(men_men_n483_), .Y(men_men_n484_));
  NA2        u0456(.A(men_men_n128_), .B(men_men_n126_), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n396_), .B(men_men_n112_), .Y(men_men_n486_));
  NO4        u0458(.A(men_men_n486_), .B(men_men_n92_), .C(men_men_n111_), .D(e), .Y(men_men_n487_));
  NO3        u0459(.A(men_men_n426_), .B(men_men_n89_), .C(men_men_n131_), .Y(men_men_n488_));
  NO4        u0460(.A(men_men_n488_), .B(men_men_n487_), .C(men_men_n485_), .D(men_men_n324_), .Y(men_men_n489_));
  NA2        u0461(.A(men_men_n489_), .B(men_men_n479_), .Y(men_men_n490_));
  NO4        u0462(.A(men_men_n490_), .B(men_men_n478_), .C(men_men_n477_), .D(men_men_n472_), .Y(men_men_n491_));
  NA2        u0463(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n492_));
  NAi31      u0464(.An(j), .B(l), .C(i), .Y(men_men_n493_));
  OAI210     u0465(.A0(men_men_n493_), .A1(men_men_n132_), .B0(men_men_n101_), .Y(men_men_n494_));
  NO3        u0466(.A(men_men_n397_), .B(men_men_n346_), .C(men_men_n201_), .Y(men_men_n495_));
  NO2        u0467(.A(men_men_n397_), .B(men_men_n372_), .Y(men_men_n496_));
  NO3        u0468(.A(men_men_n496_), .B(men_men_n495_), .C(men_men_n308_), .Y(men_men_n497_));
  NA3        u0469(.A(men_men_n497_), .B(men_men_n492_), .C(men_men_n245_), .Y(men_men_n498_));
  OAI210     u0470(.A0(men_men_n127_), .A1(men_men_n125_), .B0(n), .Y(men_men_n499_));
  NO2        u0471(.A(men_men_n499_), .B(men_men_n131_), .Y(men_men_n500_));
  BUFFER     u0472(.A(men_men_n300_), .Y(men_men_n501_));
  OA210      u0473(.A0(men_men_n501_), .A1(men_men_n500_), .B0(men_men_n192_), .Y(men_men_n502_));
  XO2        u0474(.A(i), .B(h), .Y(men_men_n503_));
  NA3        u0475(.A(men_men_n503_), .B(men_men_n161_), .C(n), .Y(men_men_n504_));
  NAi41      u0476(.An(men_men_n300_), .B(men_men_n504_), .C(men_men_n458_), .D(men_men_n385_), .Y(men_men_n505_));
  NOi32      u0477(.An(men_men_n505_), .Bn(men_men_n467_), .C(men_men_n1498_), .Y(men_men_n506_));
  NAi31      u0478(.An(c), .B(f), .C(d), .Y(men_men_n507_));
  AOI210     u0479(.A0(men_men_n280_), .A1(men_men_n195_), .B0(men_men_n507_), .Y(men_men_n508_));
  INV        u0480(.A(men_men_n508_), .Y(men_men_n509_));
  NA3        u0481(.A(men_men_n381_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n510_));
  NA2        u0482(.A(men_men_n229_), .B(men_men_n107_), .Y(men_men_n511_));
  AOI210     u0483(.A0(men_men_n511_), .A1(men_men_n182_), .B0(men_men_n507_), .Y(men_men_n512_));
  NOi21      u0484(.An(men_men_n510_), .B(men_men_n512_), .Y(men_men_n513_));
  AO220      u0485(.A0(men_men_n288_), .A1(men_men_n265_), .B0(men_men_n167_), .B1(men_men_n67_), .Y(men_men_n514_));
  NA3        u0486(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n515_));
  NO2        u0487(.A(men_men_n515_), .B(men_men_n438_), .Y(men_men_n516_));
  NO2        u0488(.A(men_men_n516_), .B(men_men_n296_), .Y(men_men_n517_));
  NAi41      u0489(.An(men_men_n514_), .B(men_men_n517_), .C(men_men_n513_), .D(men_men_n509_), .Y(men_men_n518_));
  NO4        u0490(.A(men_men_n518_), .B(men_men_n506_), .C(men_men_n502_), .D(men_men_n498_), .Y(men_men_n519_));
  NA4        u0491(.A(men_men_n519_), .B(men_men_n491_), .C(men_men_n460_), .D(men_men_n433_), .Y(men11));
  NO2        u0492(.A(men_men_n73_), .B(f), .Y(men_men_n521_));
  NA2        u0493(.A(j), .B(u), .Y(men_men_n522_));
  NAi31      u0494(.An(i), .B(m), .C(l), .Y(men_men_n523_));
  NA3        u0495(.A(m), .B(k), .C(j), .Y(men_men_n524_));
  OAI220     u0496(.A0(men_men_n524_), .A1(men_men_n131_), .B0(men_men_n523_), .B1(men_men_n522_), .Y(men_men_n525_));
  NA2        u0497(.A(men_men_n525_), .B(men_men_n521_), .Y(men_men_n526_));
  NOi32      u0498(.An(e), .Bn(b), .C(f), .Y(men_men_n527_));
  NA2        u0499(.A(men_men_n262_), .B(men_men_n112_), .Y(men_men_n528_));
  NA2        u0500(.A(men_men_n46_), .B(j), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n302_), .Y(men_men_n530_));
  NAi31      u0502(.An(d), .B(e), .C(a), .Y(men_men_n531_));
  NO2        u0503(.A(men_men_n531_), .B(n), .Y(men_men_n532_));
  AOI220     u0504(.A0(men_men_n532_), .A1(men_men_n99_), .B0(men_men_n530_), .B1(men_men_n527_), .Y(men_men_n533_));
  NAi41      u0505(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n534_));
  AN2        u0506(.A(men_men_n534_), .B(men_men_n371_), .Y(men_men_n535_));
  AOI210     u0507(.A0(men_men_n535_), .A1(men_men_n397_), .B0(men_men_n273_), .Y(men_men_n536_));
  NA2        u0508(.A(j), .B(i), .Y(men_men_n537_));
  NAi31      u0509(.An(n), .B(m), .C(k), .Y(men_men_n538_));
  NO3        u0510(.A(men_men_n538_), .B(men_men_n537_), .C(men_men_n111_), .Y(men_men_n539_));
  NO4        u0511(.A(n), .B(d), .C(men_men_n115_), .D(a), .Y(men_men_n540_));
  OR2        u0512(.A(n), .B(c), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n541_), .B(men_men_n150_), .Y(men_men_n542_));
  NO2        u0514(.A(men_men_n542_), .B(men_men_n540_), .Y(men_men_n543_));
  NOi32      u0515(.An(u), .Bn(f), .C(i), .Y(men_men_n544_));
  AOI220     u0516(.A0(men_men_n544_), .A1(men_men_n97_), .B0(men_men_n525_), .B1(f), .Y(men_men_n545_));
  NO2        u0517(.A(men_men_n275_), .B(men_men_n49_), .Y(men_men_n546_));
  NO2        u0518(.A(men_men_n545_), .B(men_men_n543_), .Y(men_men_n547_));
  AOI210     u0519(.A0(men_men_n539_), .A1(men_men_n536_), .B0(men_men_n547_), .Y(men_men_n548_));
  NA2        u0520(.A(men_men_n141_), .B(men_men_n34_), .Y(men_men_n549_));
  NAi32      u0521(.An(e), .Bn(b), .C(c), .Y(men_men_n550_));
  AN2        u0522(.A(men_men_n339_), .B(men_men_n320_), .Y(men_men_n551_));
  OAI220     u0523(.A0(men_men_n399_), .A1(men_men_n398_), .B0(men_men_n523_), .B1(men_men_n522_), .Y(men_men_n552_));
  NAi31      u0524(.An(d), .B(c), .C(a), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n553_), .B(n), .Y(men_men_n554_));
  NA3        u0526(.A(men_men_n554_), .B(men_men_n552_), .C(e), .Y(men_men_n555_));
  NO3        u0527(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n215_), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n232_), .B(men_men_n109_), .Y(men_men_n557_));
  OAI210     u0529(.A0(men_men_n556_), .A1(men_men_n400_), .B0(men_men_n557_), .Y(men_men_n558_));
  NA2        u0530(.A(men_men_n558_), .B(men_men_n555_), .Y(men_men_n559_));
  NO2        u0531(.A(men_men_n277_), .B(n), .Y(men_men_n560_));
  INV        u0532(.A(men_men_n560_), .Y(men_men_n561_));
  NA2        u0533(.A(men_men_n552_), .B(f), .Y(men_men_n562_));
  NA2        u0534(.A(h), .B(f), .Y(men_men_n563_));
  NO2        u0535(.A(men_men_n563_), .B(men_men_n92_), .Y(men_men_n564_));
  NO2        u0536(.A(men_men_n562_), .B(men_men_n561_), .Y(men_men_n565_));
  AN3        u0537(.A(j), .B(h), .C(u), .Y(men_men_n566_));
  NO2        u0538(.A(men_men_n147_), .B(c), .Y(men_men_n567_));
  NA3        u0539(.A(men_men_n567_), .B(men_men_n566_), .C(men_men_n457_), .Y(men_men_n568_));
  NA3        u0540(.A(f), .B(d), .C(b), .Y(men_men_n569_));
  NO4        u0541(.A(men_men_n569_), .B(men_men_n178_), .C(men_men_n175_), .D(u), .Y(men_men_n570_));
  NAi21      u0542(.An(men_men_n570_), .B(men_men_n568_), .Y(men_men_n571_));
  NO3        u0543(.A(men_men_n571_), .B(men_men_n565_), .C(men_men_n559_), .Y(men_men_n572_));
  AN4        u0544(.A(men_men_n572_), .B(men_men_n548_), .C(men_men_n533_), .D(men_men_n526_), .Y(men_men_n573_));
  INV        u0545(.A(k), .Y(men_men_n574_));
  NA3        u0546(.A(l), .B(men_men_n574_), .C(i), .Y(men_men_n575_));
  INV        u0547(.A(men_men_n575_), .Y(men_men_n576_));
  NA4        u0548(.A(men_men_n396_), .B(men_men_n418_), .C(men_men_n183_), .D(men_men_n112_), .Y(men_men_n577_));
  NAi32      u0549(.An(h), .Bn(f), .C(u), .Y(men_men_n578_));
  NAi41      u0550(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n579_));
  OAI210     u0551(.A0(men_men_n531_), .A1(n), .B0(men_men_n579_), .Y(men_men_n580_));
  NA2        u0552(.A(men_men_n580_), .B(m), .Y(men_men_n581_));
  NAi31      u0553(.An(h), .B(u), .C(f), .Y(men_men_n582_));
  OR3        u0554(.A(men_men_n582_), .B(men_men_n277_), .C(men_men_n49_), .Y(men_men_n583_));
  NA4        u0555(.A(men_men_n418_), .B(men_men_n120_), .C(men_men_n112_), .D(e), .Y(men_men_n584_));
  AN2        u0556(.A(men_men_n584_), .B(men_men_n583_), .Y(men_men_n585_));
  OA210      u0557(.A0(men_men_n581_), .A1(men_men_n578_), .B0(men_men_n585_), .Y(men_men_n586_));
  NO3        u0558(.A(men_men_n578_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n587_));
  NO4        u0559(.A(men_men_n582_), .B(men_men_n541_), .C(men_men_n150_), .D(men_men_n75_), .Y(men_men_n588_));
  OR2        u0560(.A(men_men_n588_), .B(men_men_n587_), .Y(men_men_n589_));
  NAi31      u0561(.An(men_men_n589_), .B(men_men_n586_), .C(men_men_n577_), .Y(men_men_n590_));
  NAi31      u0562(.An(f), .B(h), .C(u), .Y(men_men_n591_));
  NOi32      u0563(.An(b), .Bn(a), .C(c), .Y(men_men_n592_));
  NOi32      u0564(.An(d), .Bn(a), .C(e), .Y(men_men_n593_));
  NA2        u0565(.A(men_men_n593_), .B(men_men_n112_), .Y(men_men_n594_));
  NO2        u0566(.A(n), .B(c), .Y(men_men_n595_));
  NA3        u0567(.A(men_men_n595_), .B(men_men_n29_), .C(m), .Y(men_men_n596_));
  NAi32      u0568(.An(n), .Bn(f), .C(m), .Y(men_men_n597_));
  NA3        u0569(.A(men_men_n597_), .B(men_men_n596_), .C(men_men_n594_), .Y(men_men_n598_));
  NOi32      u0570(.An(e), .Bn(a), .C(d), .Y(men_men_n599_));
  AOI210     u0571(.A0(men_men_n29_), .A1(d), .B0(men_men_n599_), .Y(men_men_n600_));
  AOI210     u0572(.A0(men_men_n600_), .A1(men_men_n214_), .B0(men_men_n549_), .Y(men_men_n601_));
  NA2        u0573(.A(men_men_n601_), .B(men_men_n598_), .Y(men_men_n602_));
  OAI210     u0574(.A0(men_men_n251_), .A1(men_men_n84_), .B0(men_men_n602_), .Y(men_men_n603_));
  AOI210     u0575(.A0(men_men_n590_), .A1(men_men_n576_), .B0(men_men_n603_), .Y(men_men_n604_));
  NO3        u0576(.A(men_men_n318_), .B(men_men_n61_), .C(n), .Y(men_men_n605_));
  NA3        u0577(.A(men_men_n507_), .B(men_men_n173_), .C(men_men_n172_), .Y(men_men_n606_));
  NA2        u0578(.A(men_men_n459_), .B(men_men_n232_), .Y(men_men_n607_));
  OR2        u0579(.A(men_men_n607_), .B(men_men_n606_), .Y(men_men_n608_));
  NA2        u0580(.A(men_men_n76_), .B(men_men_n112_), .Y(men_men_n609_));
  NO2        u0581(.A(men_men_n609_), .B(men_men_n45_), .Y(men_men_n610_));
  AOI220     u0582(.A0(men_men_n610_), .A1(men_men_n536_), .B0(men_men_n608_), .B1(men_men_n605_), .Y(men_men_n611_));
  NO2        u0583(.A(men_men_n611_), .B(men_men_n84_), .Y(men_men_n612_));
  NOi32      u0584(.An(e), .Bn(c), .C(f), .Y(men_men_n613_));
  NOi21      u0585(.An(f), .B(u), .Y(men_men_n614_));
  NO2        u0586(.A(men_men_n614_), .B(men_men_n212_), .Y(men_men_n615_));
  AOI220     u0587(.A0(men_men_n615_), .A1(men_men_n393_), .B0(men_men_n613_), .B1(men_men_n177_), .Y(men_men_n616_));
  NA2        u0588(.A(men_men_n616_), .B(men_men_n180_), .Y(men_men_n617_));
  AOI210     u0589(.A0(men_men_n535_), .A1(men_men_n397_), .B0(men_men_n301_), .Y(men_men_n618_));
  NAi21      u0590(.An(k), .B(h), .Y(men_men_n619_));
  NO2        u0591(.A(men_men_n619_), .B(men_men_n264_), .Y(men_men_n620_));
  NA2        u0592(.A(men_men_n620_), .B(j), .Y(men_men_n621_));
  OR2        u0593(.A(men_men_n621_), .B(men_men_n581_), .Y(men_men_n622_));
  NOi31      u0594(.An(m), .B(n), .C(k), .Y(men_men_n623_));
  NA2        u0595(.A(j), .B(men_men_n623_), .Y(men_men_n624_));
  AOI210     u0596(.A0(men_men_n397_), .A1(men_men_n371_), .B0(men_men_n301_), .Y(men_men_n625_));
  NAi21      u0597(.An(men_men_n624_), .B(men_men_n625_), .Y(men_men_n626_));
  NO2        u0598(.A(men_men_n277_), .B(men_men_n49_), .Y(men_men_n627_));
  NO2        u0599(.A(men_men_n531_), .B(men_men_n49_), .Y(men_men_n628_));
  NA2        u0600(.A(men_men_n627_), .B(men_men_n564_), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n629_), .B(men_men_n626_), .C(men_men_n622_), .Y(men_men_n630_));
  NA2        u0602(.A(men_men_n107_), .B(men_men_n36_), .Y(men_men_n631_));
  NO2        u0603(.A(k), .B(men_men_n215_), .Y(men_men_n632_));
  INV        u0604(.A(men_men_n360_), .Y(men_men_n633_));
  NO2        u0605(.A(men_men_n633_), .B(n), .Y(men_men_n634_));
  NAi31      u0606(.An(men_men_n631_), .B(men_men_n634_), .C(men_men_n632_), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n503_), .B(men_men_n161_), .Y(men_men_n636_));
  NO3        u0608(.A(men_men_n394_), .B(men_men_n636_), .C(men_men_n84_), .Y(men_men_n637_));
  INV        u0609(.A(men_men_n637_), .Y(men_men_n638_));
  AN3        u0610(.A(f), .B(d), .C(b), .Y(men_men_n639_));
  OAI210     u0611(.A0(men_men_n639_), .A1(men_men_n130_), .B0(n), .Y(men_men_n640_));
  NA3        u0612(.A(men_men_n503_), .B(men_men_n161_), .C(men_men_n215_), .Y(men_men_n641_));
  AOI210     u0613(.A0(men_men_n640_), .A1(men_men_n234_), .B0(men_men_n641_), .Y(men_men_n642_));
  NAi31      u0614(.An(m), .B(n), .C(k), .Y(men_men_n643_));
  OR2        u0615(.A(men_men_n135_), .B(men_men_n61_), .Y(men_men_n644_));
  OAI210     u0616(.A0(men_men_n644_), .A1(men_men_n643_), .B0(men_men_n253_), .Y(men_men_n645_));
  OAI210     u0617(.A0(men_men_n645_), .A1(men_men_n642_), .B0(j), .Y(men_men_n646_));
  NA3        u0618(.A(men_men_n646_), .B(men_men_n638_), .C(men_men_n635_), .Y(men_men_n647_));
  NO4        u0619(.A(men_men_n647_), .B(men_men_n630_), .C(men_men_n617_), .D(men_men_n612_), .Y(men_men_n648_));
  NA2        u0620(.A(men_men_n381_), .B(men_men_n164_), .Y(men_men_n649_));
  NAi31      u0621(.An(u), .B(h), .C(f), .Y(men_men_n650_));
  OR3        u0622(.A(men_men_n650_), .B(men_men_n277_), .C(n), .Y(men_men_n651_));
  OA210      u0623(.A0(men_men_n531_), .A1(n), .B0(men_men_n579_), .Y(men_men_n652_));
  NA3        u0624(.A(men_men_n416_), .B(men_men_n120_), .C(men_men_n81_), .Y(men_men_n653_));
  OAI210     u0625(.A0(men_men_n652_), .A1(men_men_n88_), .B0(men_men_n653_), .Y(men_men_n654_));
  NOi21      u0626(.An(men_men_n651_), .B(men_men_n654_), .Y(men_men_n655_));
  AOI210     u0627(.A0(men_men_n655_), .A1(men_men_n649_), .B0(men_men_n524_), .Y(men_men_n656_));
  NO3        u0628(.A(u), .B(men_men_n214_), .C(men_men_n56_), .Y(men_men_n657_));
  NO2        u0629(.A(men_men_n511_), .B(men_men_n84_), .Y(men_men_n658_));
  OAI210     u0630(.A0(men_men_n658_), .A1(men_men_n393_), .B0(men_men_n657_), .Y(men_men_n659_));
  OR2        u0631(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n660_));
  NA2        u0632(.A(men_men_n592_), .B(men_men_n343_), .Y(men_men_n661_));
  OA220      u0633(.A0(men_men_n624_), .A1(men_men_n661_), .B0(men_men_n621_), .B1(men_men_n660_), .Y(men_men_n662_));
  NA3        u0634(.A(men_men_n521_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n663_));
  AN2        u0635(.A(h), .B(f), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n664_), .B(men_men_n37_), .Y(men_men_n665_));
  NA2        u0637(.A(men_men_n97_), .B(men_men_n46_), .Y(men_men_n666_));
  OAI220     u0638(.A0(men_men_n666_), .A1(men_men_n334_), .B0(men_men_n665_), .B1(men_men_n462_), .Y(men_men_n667_));
  INV        u0639(.A(men_men_n667_), .Y(men_men_n668_));
  NA4        u0640(.A(men_men_n668_), .B(men_men_n663_), .C(men_men_n662_), .D(men_men_n659_), .Y(men_men_n669_));
  NO2        u0641(.A(men_men_n255_), .B(f), .Y(men_men_n670_));
  INV        u0642(.A(men_men_n61_), .Y(men_men_n671_));
  NO3        u0643(.A(men_men_n671_), .B(men_men_n670_), .C(men_men_n34_), .Y(men_men_n672_));
  NA2        u0644(.A(men_men_n331_), .B(men_men_n141_), .Y(men_men_n673_));
  NA2        u0645(.A(men_men_n132_), .B(men_men_n49_), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n360_), .B(men_men_n112_), .Y(men_men_n675_));
  OA220      u0647(.A0(men_men_n675_), .A1(men_men_n549_), .B0(men_men_n358_), .B1(men_men_n110_), .Y(men_men_n676_));
  OAI210     u0648(.A0(men_men_n673_), .A1(men_men_n672_), .B0(men_men_n676_), .Y(men_men_n677_));
  NO3        u0649(.A(men_men_n404_), .B(men_men_n192_), .C(men_men_n191_), .Y(men_men_n678_));
  NA2        u0650(.A(men_men_n678_), .B(men_men_n232_), .Y(men_men_n679_));
  NA3        u0651(.A(men_men_n679_), .B(men_men_n257_), .C(j), .Y(men_men_n680_));
  NO3        u0652(.A(men_men_n459_), .B(men_men_n175_), .C(i), .Y(men_men_n681_));
  NA3        u0653(.A(men_men_n680_), .B(men_men_n510_), .C(men_men_n402_), .Y(men_men_n682_));
  NO4        u0654(.A(men_men_n682_), .B(men_men_n677_), .C(men_men_n669_), .D(men_men_n656_), .Y(men_men_n683_));
  NA4        u0655(.A(men_men_n683_), .B(men_men_n648_), .C(men_men_n604_), .D(men_men_n573_), .Y(men08));
  NO2        u0656(.A(k), .B(h), .Y(men_men_n685_));
  AO210      u0657(.A0(men_men_n255_), .A1(men_men_n450_), .B0(men_men_n685_), .Y(men_men_n686_));
  NO2        u0658(.A(men_men_n686_), .B(men_men_n299_), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n613_), .B(men_men_n81_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n688_), .B(men_men_n459_), .Y(men_men_n689_));
  AOI210     u0661(.A0(men_men_n689_), .A1(men_men_n687_), .B0(men_men_n488_), .Y(men_men_n690_));
  NA2        u0662(.A(men_men_n81_), .B(men_men_n109_), .Y(men_men_n691_));
  NO2        u0663(.A(men_men_n691_), .B(men_men_n57_), .Y(men_men_n692_));
  NO4        u0664(.A(men_men_n378_), .B(men_men_n111_), .C(j), .D(men_men_n215_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n569_), .B(men_men_n234_), .Y(men_men_n694_));
  AOI220     u0666(.A0(men_men_n694_), .A1(men_men_n349_), .B0(men_men_n693_), .B1(men_men_n692_), .Y(men_men_n695_));
  AOI210     u0667(.A0(men_men_n569_), .A1(men_men_n157_), .B0(men_men_n81_), .Y(men_men_n696_));
  NA4        u0668(.A(men_men_n217_), .B(men_men_n141_), .C(men_men_n45_), .D(h), .Y(men_men_n697_));
  AN2        u0669(.A(l), .B(k), .Y(men_men_n698_));
  NA4        u0670(.A(men_men_n698_), .B(men_men_n107_), .C(men_men_n75_), .D(men_men_n215_), .Y(men_men_n699_));
  NA3        u0671(.A(men_men_n695_), .B(men_men_n690_), .C(men_men_n351_), .Y(men_men_n700_));
  AN2        u0672(.A(men_men_n532_), .B(men_men_n93_), .Y(men_men_n701_));
  NO4        u0673(.A(men_men_n175_), .B(men_men_n392_), .C(men_men_n111_), .D(u), .Y(men_men_n702_));
  AOI210     u0674(.A0(men_men_n702_), .A1(men_men_n694_), .B0(men_men_n516_), .Y(men_men_n703_));
  NO2        u0675(.A(men_men_n38_), .B(men_men_n214_), .Y(men_men_n704_));
  AOI220     u0676(.A0(men_men_n615_), .A1(men_men_n348_), .B0(men_men_n704_), .B1(men_men_n560_), .Y(men_men_n705_));
  NAi31      u0677(.An(men_men_n701_), .B(men_men_n705_), .C(men_men_n703_), .Y(men_men_n706_));
  NO2        u0678(.A(men_men_n535_), .B(men_men_n35_), .Y(men_men_n707_));
  OAI210     u0679(.A0(men_men_n550_), .A1(men_men_n47_), .B0(men_men_n644_), .Y(men_men_n708_));
  NO2        u0680(.A(men_men_n481_), .B(men_men_n132_), .Y(men_men_n709_));
  AOI210     u0681(.A0(men_men_n709_), .A1(men_men_n708_), .B0(men_men_n707_), .Y(men_men_n710_));
  NO3        u0682(.A(men_men_n318_), .B(men_men_n131_), .C(men_men_n41_), .Y(men_men_n711_));
  NAi21      u0683(.An(men_men_n711_), .B(men_men_n699_), .Y(men_men_n712_));
  NA2        u0684(.A(men_men_n686_), .B(men_men_n136_), .Y(men_men_n713_));
  AOI220     u0685(.A0(men_men_n713_), .A1(men_men_n403_), .B0(men_men_n712_), .B1(men_men_n77_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n710_), .B(men_men_n714_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n360_), .B(men_men_n43_), .Y(men_men_n716_));
  NA3        u0688(.A(men_men_n679_), .B(men_men_n336_), .C(men_men_n384_), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n698_), .B(men_men_n222_), .Y(men_men_n718_));
  NO2        u0690(.A(men_men_n718_), .B(men_men_n330_), .Y(men_men_n719_));
  AOI210     u0691(.A0(men_men_n719_), .A1(men_men_n670_), .B0(men_men_n487_), .Y(men_men_n720_));
  NA3        u0692(.A(m), .B(l), .C(k), .Y(men_men_n721_));
  AOI210     u0693(.A0(men_men_n653_), .A1(men_men_n651_), .B0(men_men_n721_), .Y(men_men_n722_));
  NO2        u0694(.A(men_men_n534_), .B(men_men_n273_), .Y(men_men_n723_));
  NOi21      u0695(.An(men_men_n723_), .B(men_men_n528_), .Y(men_men_n724_));
  NA4        u0696(.A(men_men_n112_), .B(l), .C(k), .D(men_men_n84_), .Y(men_men_n725_));
  NA3        u0697(.A(men_men_n120_), .B(men_men_n411_), .C(i), .Y(men_men_n726_));
  NO2        u0698(.A(men_men_n726_), .B(men_men_n725_), .Y(men_men_n727_));
  NO3        u0699(.A(men_men_n727_), .B(men_men_n724_), .C(men_men_n722_), .Y(men_men_n728_));
  NA4        u0700(.A(men_men_n728_), .B(men_men_n720_), .C(men_men_n717_), .D(men_men_n716_), .Y(men_men_n729_));
  NO4        u0701(.A(men_men_n729_), .B(men_men_n715_), .C(men_men_n706_), .D(men_men_n700_), .Y(men_men_n730_));
  NA2        u0702(.A(men_men_n615_), .B(men_men_n393_), .Y(men_men_n731_));
  NOi31      u0703(.An(u), .B(h), .C(f), .Y(men_men_n732_));
  NA2        u0704(.A(men_men_n628_), .B(men_men_n732_), .Y(men_men_n733_));
  AO210      u0705(.A0(men_men_n733_), .A1(men_men_n583_), .B0(men_men_n537_), .Y(men_men_n734_));
  INV        u0706(.A(men_men_n496_), .Y(men_men_n735_));
  NA4        u0707(.A(men_men_n735_), .B(men_men_n734_), .C(men_men_n731_), .D(men_men_n254_), .Y(men_men_n736_));
  NA2        u0708(.A(men_men_n698_), .B(men_men_n75_), .Y(men_men_n737_));
  NO3        u0709(.A(men_men_n678_), .B(men_men_n175_), .C(i), .Y(men_men_n738_));
  NOi21      u0710(.An(h), .B(j), .Y(men_men_n739_));
  NA2        u0711(.A(men_men_n739_), .B(f), .Y(men_men_n740_));
  NO2        u0712(.A(men_men_n740_), .B(men_men_n248_), .Y(men_men_n741_));
  NO3        u0713(.A(men_men_n741_), .B(men_men_n738_), .C(men_men_n681_), .Y(men_men_n742_));
  OAI220     u0714(.A0(men_men_n742_), .A1(men_men_n737_), .B0(men_men_n585_), .B1(men_men_n62_), .Y(men_men_n743_));
  AOI210     u0715(.A0(men_men_n736_), .A1(l), .B0(men_men_n743_), .Y(men_men_n744_));
  NO2        u0716(.A(j), .B(i), .Y(men_men_n745_));
  NA3        u0717(.A(men_men_n745_), .B(men_men_n79_), .C(l), .Y(men_men_n746_));
  NA2        u0718(.A(men_men_n745_), .B(men_men_n33_), .Y(men_men_n747_));
  NA2        u0719(.A(men_men_n421_), .B(men_men_n120_), .Y(men_men_n748_));
  OA220      u0720(.A0(men_men_n748_), .A1(men_men_n747_), .B0(men_men_n746_), .B1(men_men_n581_), .Y(men_men_n749_));
  NO3        u0721(.A(men_men_n152_), .B(men_men_n49_), .C(men_men_n109_), .Y(men_men_n750_));
  NO3        u0722(.A(men_men_n541_), .B(men_men_n150_), .C(men_men_n75_), .Y(men_men_n751_));
  NO3        u0723(.A(men_men_n481_), .B(men_men_n439_), .C(j), .Y(men_men_n752_));
  OAI210     u0724(.A0(men_men_n751_), .A1(men_men_n750_), .B0(men_men_n752_), .Y(men_men_n753_));
  OAI210     u0725(.A0(men_men_n733_), .A1(men_men_n62_), .B0(men_men_n753_), .Y(men_men_n754_));
  NA2        u0726(.A(k), .B(j), .Y(men_men_n755_));
  NO3        u0727(.A(men_men_n175_), .B(men_men_n392_), .C(men_men_n111_), .Y(men_men_n756_));
  NA2        u0728(.A(men_men_n756_), .B(men_men_n249_), .Y(men_men_n757_));
  NAi31      u0729(.An(men_men_n600_), .B(men_men_n90_), .C(men_men_n81_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n758_), .B(men_men_n757_), .Y(men_men_n759_));
  NO2        u0731(.A(men_men_n299_), .B(men_men_n136_), .Y(men_men_n760_));
  AOI220     u0732(.A0(men_men_n760_), .A1(men_men_n615_), .B0(men_men_n711_), .B1(men_men_n696_), .Y(men_men_n761_));
  NO2        u0733(.A(men_men_n721_), .B(men_men_n88_), .Y(men_men_n762_));
  NA2        u0734(.A(men_men_n762_), .B(men_men_n580_), .Y(men_men_n763_));
  NA2        u0735(.A(men_men_n763_), .B(men_men_n761_), .Y(men_men_n764_));
  OR3        u0736(.A(men_men_n764_), .B(men_men_n759_), .C(men_men_n754_), .Y(men_men_n765_));
  NO4        u0737(.A(men_men_n481_), .B(men_men_n434_), .C(j), .D(f), .Y(men_men_n766_));
  OAI220     u0738(.A0(men_men_n697_), .A1(men_men_n688_), .B0(men_men_n334_), .B1(men_men_n38_), .Y(men_men_n767_));
  AOI210     u0739(.A0(men_men_n766_), .A1(men_men_n261_), .B0(men_men_n767_), .Y(men_men_n768_));
  NA3        u0740(.A(men_men_n544_), .B(men_men_n292_), .C(h), .Y(men_men_n769_));
  NO2        u0741(.A(men_men_n89_), .B(men_men_n47_), .Y(men_men_n770_));
  OAI220     u0742(.A0(men_men_n769_), .A1(men_men_n596_), .B0(men_men_n746_), .B1(men_men_n660_), .Y(men_men_n771_));
  AOI210     u0743(.A0(men_men_n770_), .A1(men_men_n634_), .B0(men_men_n771_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n772_), .B(men_men_n768_), .Y(men_men_n773_));
  BUFFER     u0745(.A(men_men_n93_), .Y(men_men_n774_));
  AOI220     u0746(.A0(men_men_n774_), .A1(men_men_n240_), .B0(men_men_n752_), .B1(men_men_n627_), .Y(men_men_n775_));
  NO2        u0747(.A(men_men_n652_), .B(men_men_n75_), .Y(men_men_n776_));
  NA2        u0748(.A(men_men_n766_), .B(men_men_n776_), .Y(men_men_n777_));
  OAI210     u0749(.A0(men_men_n721_), .A1(men_men_n650_), .B0(men_men_n515_), .Y(men_men_n778_));
  NA3        u0750(.A(men_men_n252_), .B(men_men_n59_), .C(b), .Y(men_men_n779_));
  AOI220     u0751(.A0(men_men_n595_), .A1(men_men_n29_), .B0(men_men_n461_), .B1(men_men_n81_), .Y(men_men_n780_));
  NA2        u0752(.A(men_men_n780_), .B(men_men_n779_), .Y(men_men_n781_));
  NO2        u0753(.A(men_men_n769_), .B(men_men_n486_), .Y(men_men_n782_));
  AOI210     u0754(.A0(men_men_n781_), .A1(men_men_n778_), .B0(men_men_n782_), .Y(men_men_n783_));
  NA3        u0755(.A(men_men_n783_), .B(men_men_n777_), .C(men_men_n775_), .Y(men_men_n784_));
  NOi41      u0756(.An(men_men_n749_), .B(men_men_n784_), .C(men_men_n773_), .D(men_men_n765_), .Y(men_men_n785_));
  OR2        u0757(.A(men_men_n697_), .B(men_men_n234_), .Y(men_men_n786_));
  NA2        u0758(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n787_));
  NO3        u0759(.A(men_men_n787_), .B(men_men_n747_), .C(men_men_n277_), .Y(men_men_n788_));
  NO3        u0760(.A(men_men_n522_), .B(men_men_n91_), .C(h), .Y(men_men_n789_));
  AOI210     u0761(.A0(men_men_n789_), .A1(men_men_n692_), .B0(men_men_n788_), .Y(men_men_n790_));
  NA2        u0762(.A(men_men_n790_), .B(men_men_n786_), .Y(men_men_n791_));
  OR2        u0763(.A(men_men_n650_), .B(men_men_n89_), .Y(men_men_n792_));
  NOi31      u0764(.An(b), .B(d), .C(a), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n793_), .B(men_men_n593_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n794_), .B(n), .Y(men_men_n795_));
  BUFFER     u0767(.A(men_men_n780_), .Y(men_men_n796_));
  OAI220     u0768(.A0(men_men_n796_), .A1(men_men_n792_), .B0(men_men_n769_), .B1(men_men_n594_), .Y(men_men_n797_));
  NO2        u0769(.A(men_men_n330_), .B(men_men_n116_), .Y(men_men_n798_));
  NOi21      u0770(.An(men_men_n798_), .B(men_men_n162_), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n678_), .B(n), .Y(men_men_n800_));
  AOI220     u0772(.A0(men_men_n760_), .A1(men_men_n657_), .B0(men_men_n800_), .B1(men_men_n687_), .Y(men_men_n801_));
  NO2        u0773(.A(men_men_n325_), .B(men_men_n239_), .Y(men_men_n802_));
  OAI210     u0774(.A0(men_men_n93_), .A1(men_men_n90_), .B0(men_men_n802_), .Y(men_men_n803_));
  NA2        u0775(.A(men_men_n120_), .B(men_men_n81_), .Y(men_men_n804_));
  AOI210     u0776(.A0(men_men_n425_), .A1(men_men_n417_), .B0(men_men_n804_), .Y(men_men_n805_));
  NAi21      u0777(.An(men_men_n805_), .B(men_men_n803_), .Y(men_men_n806_));
  NA2        u0778(.A(men_men_n719_), .B(men_men_n34_), .Y(men_men_n807_));
  NAi21      u0779(.An(men_men_n725_), .B(men_men_n435_), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n273_), .B(i), .Y(men_men_n809_));
  NA2        u0781(.A(men_men_n702_), .B(men_men_n350_), .Y(men_men_n810_));
  OAI210     u0782(.A0(men_men_n588_), .A1(men_men_n587_), .B0(men_men_n361_), .Y(men_men_n811_));
  AN3        u0783(.A(men_men_n811_), .B(men_men_n810_), .C(men_men_n808_), .Y(men_men_n812_));
  NAi41      u0784(.An(men_men_n806_), .B(men_men_n812_), .C(men_men_n807_), .D(men_men_n801_), .Y(men_men_n813_));
  NO4        u0785(.A(men_men_n813_), .B(men_men_n799_), .C(men_men_n797_), .D(men_men_n791_), .Y(men_men_n814_));
  NA4        u0786(.A(men_men_n814_), .B(men_men_n785_), .C(men_men_n744_), .D(men_men_n730_), .Y(men09));
  INV        u0787(.A(men_men_n121_), .Y(men_men_n816_));
  NA2        u0788(.A(f), .B(e), .Y(men_men_n817_));
  NO2        u0789(.A(men_men_n227_), .B(men_men_n111_), .Y(men_men_n818_));
  NA2        u0790(.A(men_men_n818_), .B(u), .Y(men_men_n819_));
  NA3        u0791(.A(men_men_n311_), .B(men_men_n469_), .C(men_men_n118_), .Y(men_men_n820_));
  AOI210     u0792(.A0(men_men_n820_), .A1(u), .B0(men_men_n466_), .Y(men_men_n821_));
  AOI210     u0793(.A0(men_men_n821_), .A1(men_men_n819_), .B0(men_men_n817_), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n443_), .B(e), .Y(men_men_n823_));
  NO2        u0795(.A(men_men_n823_), .B(men_men_n507_), .Y(men_men_n824_));
  AOI210     u0796(.A0(men_men_n822_), .A1(men_men_n816_), .B0(men_men_n824_), .Y(men_men_n825_));
  NO2        u0797(.A(men_men_n204_), .B(men_men_n214_), .Y(men_men_n826_));
  NA3        u0798(.A(m), .B(l), .C(i), .Y(men_men_n827_));
  OAI220     u0799(.A0(men_men_n582_), .A1(men_men_n827_), .B0(men_men_n355_), .B1(men_men_n523_), .Y(men_men_n828_));
  NA4        u0800(.A(men_men_n85_), .B(men_men_n84_), .C(u), .D(f), .Y(men_men_n829_));
  OR2        u0801(.A(men_men_n828_), .B(men_men_n826_), .Y(men_men_n830_));
  NA3        u0802(.A(men_men_n792_), .B(men_men_n562_), .C(men_men_n515_), .Y(men_men_n831_));
  OA210      u0803(.A0(men_men_n831_), .A1(men_men_n830_), .B0(men_men_n795_), .Y(men_men_n832_));
  INV        u0804(.A(men_men_n339_), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n834_));
  NA2        u0806(.A(men_men_n779_), .B(men_men_n334_), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n343_), .B(men_men_n345_), .Y(men_men_n836_));
  INV        u0808(.A(men_men_n836_), .Y(men_men_n837_));
  NA2        u0809(.A(men_men_n837_), .B(men_men_n835_), .Y(men_men_n838_));
  INV        u0810(.A(men_men_n113_), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n839_), .B(men_men_n686_), .Y(men_men_n840_));
  NA3        u0812(.A(men_men_n840_), .B(men_men_n189_), .C(men_men_n31_), .Y(men_men_n841_));
  NA3        u0813(.A(men_men_n841_), .B(men_men_n838_), .C(men_men_n616_), .Y(men_men_n842_));
  NO2        u0814(.A(men_men_n578_), .B(men_men_n493_), .Y(men_men_n843_));
  NOi21      u0815(.An(f), .B(d), .Y(men_men_n844_));
  NA2        u0816(.A(men_men_n844_), .B(m), .Y(men_men_n845_));
  NO2        u0817(.A(men_men_n845_), .B(men_men_n52_), .Y(men_men_n846_));
  NOi32      u0818(.An(u), .Bn(f), .C(d), .Y(men_men_n847_));
  NA4        u0819(.A(men_men_n847_), .B(men_men_n595_), .C(men_men_n29_), .D(m), .Y(men_men_n848_));
  NOi21      u0820(.An(men_men_n312_), .B(men_men_n848_), .Y(men_men_n849_));
  AOI210     u0821(.A0(men_men_n846_), .A1(men_men_n542_), .B0(men_men_n849_), .Y(men_men_n850_));
  NA2        u0822(.A(men_men_n311_), .B(men_men_n118_), .Y(men_men_n851_));
  AN2        u0823(.A(f), .B(d), .Y(men_men_n852_));
  NA3        u0824(.A(men_men_n474_), .B(men_men_n852_), .C(men_men_n81_), .Y(men_men_n853_));
  NO3        u0825(.A(men_men_n853_), .B(men_men_n75_), .C(men_men_n215_), .Y(men_men_n854_));
  NO2        u0826(.A(men_men_n285_), .B(men_men_n56_), .Y(men_men_n855_));
  NA2        u0827(.A(men_men_n851_), .B(men_men_n854_), .Y(men_men_n856_));
  NAi31      u0828(.An(men_men_n485_), .B(men_men_n856_), .C(men_men_n850_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n643_), .B(men_men_n330_), .Y(men_men_n858_));
  AN2        u0830(.A(men_men_n858_), .B(men_men_n670_), .Y(men_men_n859_));
  NO2        u0831(.A(men_men_n859_), .B(men_men_n236_), .Y(men_men_n860_));
  NA2        u0832(.A(men_men_n593_), .B(men_men_n81_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n836_), .B(men_men_n861_), .Y(men_men_n862_));
  NA3        u0834(.A(men_men_n161_), .B(men_men_n107_), .C(men_men_n106_), .Y(men_men_n863_));
  OAI220     u0835(.A0(men_men_n853_), .A1(men_men_n429_), .B0(men_men_n339_), .B1(men_men_n863_), .Y(men_men_n864_));
  NOi41      u0836(.An(men_men_n225_), .B(men_men_n864_), .C(men_men_n862_), .D(men_men_n308_), .Y(men_men_n865_));
  NA2        u0837(.A(c), .B(men_men_n115_), .Y(men_men_n866_));
  NO2        u0838(.A(men_men_n866_), .B(men_men_n408_), .Y(men_men_n867_));
  NA3        u0839(.A(men_men_n867_), .B(men_men_n505_), .C(f), .Y(men_men_n868_));
  OR2        u0840(.A(men_men_n650_), .B(men_men_n538_), .Y(men_men_n869_));
  INV        u0841(.A(men_men_n869_), .Y(men_men_n870_));
  NA2        u0842(.A(men_men_n794_), .B(men_men_n110_), .Y(men_men_n871_));
  NA2        u0843(.A(men_men_n871_), .B(men_men_n870_), .Y(men_men_n872_));
  NA4        u0844(.A(men_men_n872_), .B(men_men_n868_), .C(men_men_n865_), .D(men_men_n860_), .Y(men_men_n873_));
  NO4        u0845(.A(men_men_n873_), .B(men_men_n857_), .C(men_men_n842_), .D(men_men_n832_), .Y(men_men_n874_));
  NA2        u0846(.A(men_men_n111_), .B(j), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n334_), .B(men_men_n829_), .Y(men_men_n876_));
  NO2        u0848(.A(men_men_n136_), .B(men_men_n132_), .Y(men_men_n877_));
  NO2        u0849(.A(men_men_n232_), .B(men_men_n226_), .Y(men_men_n878_));
  AOI220     u0850(.A0(men_men_n878_), .A1(men_men_n229_), .B0(men_men_n306_), .B1(men_men_n877_), .Y(men_men_n879_));
  NO2        u0851(.A(men_men_n429_), .B(men_men_n817_), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n880_), .B(men_men_n554_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n881_), .B(men_men_n879_), .Y(men_men_n882_));
  NA2        u0854(.A(e), .B(d), .Y(men_men_n883_));
  OAI220     u0855(.A0(men_men_n883_), .A1(c), .B0(men_men_n325_), .B1(d), .Y(men_men_n884_));
  NA3        u0856(.A(men_men_n884_), .B(men_men_n454_), .C(men_men_n503_), .Y(men_men_n885_));
  AOI210     u0857(.A0(men_men_n511_), .A1(men_men_n182_), .B0(men_men_n232_), .Y(men_men_n886_));
  AOI210     u0858(.A0(men_men_n615_), .A1(men_men_n348_), .B0(men_men_n886_), .Y(men_men_n887_));
  NA2        u0859(.A(men_men_n285_), .B(men_men_n166_), .Y(men_men_n888_));
  NA2        u0860(.A(men_men_n854_), .B(men_men_n888_), .Y(men_men_n889_));
  NA3        u0861(.A(men_men_n169_), .B(men_men_n82_), .C(men_men_n34_), .Y(men_men_n890_));
  NA4        u0862(.A(men_men_n890_), .B(men_men_n889_), .C(men_men_n887_), .D(men_men_n885_), .Y(men_men_n891_));
  NO3        u0863(.A(men_men_n891_), .B(men_men_n882_), .C(men_men_n876_), .Y(men_men_n892_));
  NA2        u0864(.A(men_men_n833_), .B(men_men_n31_), .Y(men_men_n893_));
  OR2        u0865(.A(men_men_n893_), .B(men_men_n218_), .Y(men_men_n894_));
  OAI220     u0866(.A0(men_men_n614_), .A1(men_men_n61_), .B0(men_men_n301_), .B1(j), .Y(men_men_n895_));
  AOI220     u0867(.A0(men_men_n895_), .A1(men_men_n858_), .B0(men_men_n605_), .B1(men_men_n613_), .Y(men_men_n896_));
  OAI210     u0868(.A0(men_men_n823_), .A1(men_men_n172_), .B0(men_men_n896_), .Y(men_men_n897_));
  OAI210     u0869(.A0(men_men_n818_), .A1(men_men_n888_), .B0(men_men_n847_), .Y(men_men_n898_));
  NO2        u0870(.A(men_men_n898_), .B(men_men_n596_), .Y(men_men_n899_));
  AOI210     u0871(.A0(men_men_n117_), .A1(men_men_n116_), .B0(men_men_n262_), .Y(men_men_n900_));
  NO2        u0872(.A(men_men_n900_), .B(men_men_n848_), .Y(men_men_n901_));
  AO210      u0873(.A0(men_men_n835_), .A1(men_men_n828_), .B0(men_men_n901_), .Y(men_men_n902_));
  NOi31      u0874(.An(men_men_n542_), .B(men_men_n845_), .C(men_men_n293_), .Y(men_men_n903_));
  NO4        u0875(.A(men_men_n903_), .B(men_men_n902_), .C(men_men_n899_), .D(men_men_n897_), .Y(men_men_n904_));
  AO220      u0876(.A0(men_men_n454_), .A1(men_men_n739_), .B0(men_men_n177_), .B1(f), .Y(men_men_n905_));
  NA2        u0877(.A(men_men_n905_), .B(men_men_n884_), .Y(men_men_n906_));
  NO2        u0878(.A(men_men_n439_), .B(men_men_n71_), .Y(men_men_n907_));
  OAI210     u0879(.A0(men_men_n831_), .A1(men_men_n907_), .B0(men_men_n692_), .Y(men_men_n908_));
  AN4        u0880(.A(men_men_n908_), .B(men_men_n906_), .C(men_men_n904_), .D(men_men_n894_), .Y(men_men_n909_));
  NA4        u0881(.A(men_men_n909_), .B(men_men_n892_), .C(men_men_n874_), .D(men_men_n825_), .Y(men12));
  NO4        u0882(.A(men_men_n442_), .B(men_men_n255_), .C(men_men_n574_), .D(men_men_n215_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n542_), .B(men_men_n907_), .Y(men_men_n912_));
  NO2        u0884(.A(men_men_n452_), .B(men_men_n115_), .Y(men_men_n913_));
  NO2        u0885(.A(men_men_n834_), .B(men_men_n355_), .Y(men_men_n914_));
  NO2        u0886(.A(men_men_n650_), .B(men_men_n378_), .Y(men_men_n915_));
  AOI220     u0887(.A0(men_men_n915_), .A1(men_men_n540_), .B0(men_men_n914_), .B1(men_men_n913_), .Y(men_men_n916_));
  NA3        u0888(.A(men_men_n916_), .B(men_men_n912_), .C(men_men_n441_), .Y(men_men_n917_));
  AOI210     u0889(.A0(men_men_n235_), .A1(men_men_n338_), .B0(men_men_n201_), .Y(men_men_n918_));
  OR2        u0890(.A(men_men_n918_), .B(men_men_n911_), .Y(men_men_n919_));
  NO2        u0891(.A(men_men_n390_), .B(men_men_n215_), .Y(men_men_n920_));
  OAI210     u0892(.A0(men_men_n920_), .A1(men_men_n919_), .B0(men_men_n404_), .Y(men_men_n921_));
  NO2        u0893(.A(men_men_n631_), .B(men_men_n264_), .Y(men_men_n922_));
  NO2        u0894(.A(men_men_n582_), .B(men_men_n827_), .Y(men_men_n923_));
  AOI220     u0895(.A0(men_men_n923_), .A1(men_men_n560_), .B0(men_men_n802_), .B1(men_men_n922_), .Y(men_men_n924_));
  NO2        u0896(.A(men_men_n152_), .B(men_men_n239_), .Y(men_men_n925_));
  NA3        u0897(.A(men_men_n925_), .B(men_men_n242_), .C(i), .Y(men_men_n926_));
  NA3        u0898(.A(men_men_n926_), .B(men_men_n924_), .C(men_men_n921_), .Y(men_men_n927_));
  NA4        u0899(.A(men_men_n443_), .B(men_men_n437_), .C(men_men_n183_), .D(u), .Y(men_men_n928_));
  INV        u0900(.A(men_men_n928_), .Y(men_men_n929_));
  NO3        u0901(.A(men_men_n655_), .B(men_men_n89_), .C(men_men_n45_), .Y(men_men_n930_));
  NO4        u0902(.A(men_men_n930_), .B(men_men_n929_), .C(men_men_n927_), .D(men_men_n917_), .Y(men_men_n931_));
  NO2        u0903(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n932_));
  INV        u0904(.A(men_men_n579_), .Y(men_men_n933_));
  NOi21      u0905(.An(men_men_n34_), .B(men_men_n643_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n933_), .B(men_men_n932_), .Y(men_men_n935_));
  OAI210     u0907(.A0(men_men_n253_), .A1(men_men_n45_), .B0(men_men_n935_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n435_), .B(men_men_n266_), .Y(men_men_n937_));
  NO3        u0909(.A(men_men_n804_), .B(men_men_n86_), .C(men_men_n408_), .Y(men_men_n938_));
  NAi31      u0910(.An(men_men_n938_), .B(men_men_n937_), .C(men_men_n322_), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n623_), .B(men_men_n361_), .Y(men_men_n941_));
  OAI210     u0913(.A0(men_men_n726_), .A1(men_men_n941_), .B0(men_men_n365_), .Y(men_men_n942_));
  NO3        u0914(.A(men_men_n942_), .B(men_men_n939_), .C(men_men_n936_), .Y(men_men_n943_));
  NA2        u0915(.A(men_men_n164_), .B(i), .Y(men_men_n944_));
  NA2        u0916(.A(men_men_n46_), .B(i), .Y(men_men_n945_));
  OAI220     u0917(.A0(men_men_n945_), .A1(men_men_n200_), .B0(men_men_n944_), .B1(men_men_n89_), .Y(men_men_n946_));
  AOI210     u0918(.A0(men_men_n419_), .A1(men_men_n37_), .B0(men_men_n946_), .Y(men_men_n947_));
  NA2        u0919(.A(men_men_n550_), .B(men_men_n382_), .Y(men_men_n948_));
  NO2        u0920(.A(men_men_n947_), .B(men_men_n334_), .Y(men_men_n949_));
  NA3        u0921(.A(men_men_n343_), .B(j), .C(i), .Y(men_men_n950_));
  NA2        u0922(.A(men_men_n599_), .B(men_men_n112_), .Y(men_men_n951_));
  OR3        u0923(.A(men_men_n311_), .B(men_men_n434_), .C(f), .Y(men_men_n952_));
  NA3        u0924(.A(j), .B(men_men_n79_), .C(i), .Y(men_men_n953_));
  OA220      u0925(.A0(men_men_n953_), .A1(men_men_n951_), .B0(men_men_n952_), .B1(men_men_n581_), .Y(men_men_n954_));
  NA3        u0926(.A(men_men_n327_), .B(men_men_n117_), .C(u), .Y(men_men_n955_));
  AOI210     u0927(.A0(men_men_n665_), .A1(men_men_n955_), .B0(m), .Y(men_men_n956_));
  OAI210     u0928(.A0(men_men_n956_), .A1(men_men_n914_), .B0(men_men_n326_), .Y(men_men_n957_));
  INV        u0929(.A(men_men_n861_), .Y(men_men_n958_));
  NA2        u0930(.A(men_men_n829_), .B(men_men_n440_), .Y(men_men_n959_));
  NA2        u0931(.A(men_men_n223_), .B(men_men_n78_), .Y(men_men_n960_));
  NA3        u0932(.A(men_men_n960_), .B(men_men_n953_), .C(men_men_n952_), .Y(men_men_n961_));
  AOI220     u0933(.A0(men_men_n961_), .A1(men_men_n261_), .B0(men_men_n959_), .B1(men_men_n958_), .Y(men_men_n962_));
  NA3        u0934(.A(men_men_n962_), .B(men_men_n957_), .C(men_men_n954_), .Y(men_men_n963_));
  NA2        u0935(.A(men_men_n654_), .B(men_men_n85_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n458_), .B(men_men_n215_), .Y(men_men_n965_));
  NA2        u0937(.A(men_men_n965_), .B(men_men_n383_), .Y(men_men_n966_));
  NA2        u0938(.A(men_men_n580_), .B(men_men_n87_), .Y(men_men_n967_));
  NA3        u0939(.A(men_men_n967_), .B(men_men_n966_), .C(men_men_n964_), .Y(men_men_n968_));
  AOI210     u0940(.A0(men_men_n420_), .A1(men_men_n412_), .B0(men_men_n804_), .Y(men_men_n969_));
  OAI210     u0941(.A0(men_men_n368_), .A1(men_men_n367_), .B0(men_men_n108_), .Y(men_men_n970_));
  AOI210     u0942(.A0(men_men_n970_), .A1(men_men_n532_), .B0(men_men_n969_), .Y(men_men_n971_));
  NA2        u0943(.A(men_men_n956_), .B(men_men_n913_), .Y(men_men_n972_));
  NO3        u0944(.A(men_men_n875_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n973_));
  NA2        u0945(.A(men_men_n973_), .B(men_men_n618_), .Y(men_men_n974_));
  NA3        u0946(.A(men_men_n974_), .B(men_men_n972_), .C(men_men_n971_), .Y(men_men_n975_));
  NO4        u0947(.A(men_men_n975_), .B(men_men_n968_), .C(men_men_n963_), .D(men_men_n949_), .Y(men_men_n976_));
  NAi31      u0948(.An(men_men_n142_), .B(men_men_n421_), .C(n), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n125_), .B(men_men_n341_), .Y(men_men_n978_));
  NO2        u0950(.A(men_men_n978_), .B(men_men_n977_), .Y(men_men_n979_));
  NO3        u0951(.A(men_men_n273_), .B(men_men_n142_), .C(men_men_n408_), .Y(men_men_n980_));
  AOI210     u0952(.A0(men_men_n980_), .A1(men_men_n494_), .B0(men_men_n979_), .Y(men_men_n981_));
  NA2        u0953(.A(men_men_n488_), .B(i), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n982_), .B(men_men_n981_), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n232_), .B(men_men_n173_), .Y(men_men_n984_));
  NO2        u0956(.A(men_men_n443_), .B(men_men_n177_), .Y(men_men_n985_));
  NOi31      u0957(.An(men_men_n984_), .B(men_men_n985_), .C(men_men_n215_), .Y(men_men_n986_));
  NA2        u0958(.A(men_men_n438_), .B(men_men_n861_), .Y(men_men_n987_));
  NO3        u0959(.A(men_men_n439_), .B(men_men_n311_), .C(men_men_n75_), .Y(men_men_n988_));
  AOI220     u0960(.A0(men_men_n988_), .A1(men_men_n987_), .B0(men_men_n478_), .B1(u), .Y(men_men_n989_));
  INV        u0961(.A(men_men_n989_), .Y(men_men_n990_));
  OAI220     u0962(.A0(men_men_n977_), .A1(men_men_n235_), .B0(men_men_n950_), .B1(men_men_n594_), .Y(men_men_n991_));
  NO2        u0963(.A(men_men_n651_), .B(men_men_n378_), .Y(men_men_n992_));
  NO3        u0964(.A(men_men_n541_), .B(men_men_n150_), .C(men_men_n214_), .Y(men_men_n993_));
  OAI210     u0965(.A0(men_men_n993_), .A1(men_men_n521_), .B0(men_men_n379_), .Y(men_men_n994_));
  OAI220     u0966(.A0(men_men_n915_), .A1(men_men_n923_), .B0(men_men_n542_), .B1(men_men_n428_), .Y(men_men_n995_));
  NA2        u0967(.A(men_men_n995_), .B(men_men_n994_), .Y(men_men_n996_));
  OAI210     u0968(.A0(men_men_n918_), .A1(men_men_n911_), .B0(men_men_n984_), .Y(men_men_n997_));
  NA3        u0969(.A(men_men_n948_), .B(men_men_n483_), .C(men_men_n46_), .Y(men_men_n998_));
  NA2        u0970(.A(men_men_n381_), .B(men_men_n379_), .Y(men_men_n999_));
  NA4        u0971(.A(men_men_n999_), .B(men_men_n998_), .C(men_men_n997_), .D(men_men_n274_), .Y(men_men_n1000_));
  OR4        u0972(.A(men_men_n1000_), .B(men_men_n996_), .C(men_men_n992_), .D(men_men_n991_), .Y(men_men_n1001_));
  NO4        u0973(.A(men_men_n1001_), .B(men_men_n990_), .C(men_men_n986_), .D(men_men_n983_), .Y(men_men_n1002_));
  NA4        u0974(.A(men_men_n1002_), .B(men_men_n976_), .C(men_men_n943_), .D(men_men_n931_), .Y(men13));
  NA2        u0975(.A(men_men_n46_), .B(men_men_n84_), .Y(men_men_n1004_));
  AN2        u0976(.A(c), .B(b), .Y(men_men_n1005_));
  NA3        u0977(.A(men_men_n252_), .B(men_men_n1005_), .C(m), .Y(men_men_n1006_));
  NO4        u0978(.A(e), .B(men_men_n1006_), .C(men_men_n1004_), .D(men_men_n575_), .Y(men_men_n1007_));
  NA2        u0979(.A(men_men_n266_), .B(men_men_n1005_), .Y(men_men_n1008_));
  NO4        u0980(.A(men_men_n1008_), .B(e), .C(men_men_n944_), .D(a), .Y(men_men_n1009_));
  NAi32      u0981(.An(d), .Bn(c), .C(e), .Y(men_men_n1010_));
  NA2        u0982(.A(men_men_n141_), .B(men_men_n45_), .Y(men_men_n1011_));
  NO4        u0983(.A(men_men_n1011_), .B(men_men_n1010_), .C(men_men_n582_), .D(men_men_n309_), .Y(men_men_n1012_));
  NA2        u0984(.A(men_men_n411_), .B(men_men_n214_), .Y(men_men_n1013_));
  AN2        u0985(.A(d), .B(c), .Y(men_men_n1014_));
  NA2        u0986(.A(men_men_n1014_), .B(men_men_n115_), .Y(men_men_n1015_));
  NO4        u0987(.A(men_men_n1015_), .B(men_men_n1013_), .C(men_men_n178_), .D(men_men_n170_), .Y(men_men_n1016_));
  NA2        u0988(.A(d), .B(c), .Y(men_men_n1017_));
  NO4        u0989(.A(men_men_n1011_), .B(men_men_n578_), .C(men_men_n1017_), .D(men_men_n309_), .Y(men_men_n1018_));
  OR2        u0990(.A(men_men_n1016_), .B(men_men_n1018_), .Y(men_men_n1019_));
  OR4        u0991(.A(men_men_n1019_), .B(men_men_n1012_), .C(men_men_n1009_), .D(men_men_n1007_), .Y(men_men_n1020_));
  NAi32      u0992(.An(f), .Bn(e), .C(c), .Y(men_men_n1021_));
  NO2        u0993(.A(men_men_n1021_), .B(men_men_n147_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n1022_), .B(u), .Y(men_men_n1023_));
  OR3        u0995(.A(men_men_n226_), .B(men_men_n178_), .C(men_men_n170_), .Y(men_men_n1024_));
  NO2        u0996(.A(men_men_n1024_), .B(men_men_n1023_), .Y(men_men_n1025_));
  NO2        u0997(.A(men_men_n1017_), .B(men_men_n309_), .Y(men_men_n1026_));
  NO2        u0998(.A(j), .B(men_men_n45_), .Y(men_men_n1027_));
  NA2        u0999(.A(men_men_n620_), .B(men_men_n1027_), .Y(men_men_n1028_));
  NOi21      u1000(.An(men_men_n1026_), .B(men_men_n1028_), .Y(men_men_n1029_));
  NO2        u1001(.A(men_men_n755_), .B(men_men_n111_), .Y(men_men_n1030_));
  NOi41      u1002(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1031_));
  NA2        u1003(.A(men_men_n1031_), .B(men_men_n1030_), .Y(men_men_n1032_));
  NO2        u1004(.A(men_men_n1032_), .B(men_men_n1023_), .Y(men_men_n1033_));
  OR3        u1005(.A(e), .B(d), .C(c), .Y(men_men_n1034_));
  NA3        u1006(.A(k), .B(j), .C(i), .Y(men_men_n1035_));
  NO3        u1007(.A(men_men_n1035_), .B(men_men_n309_), .C(men_men_n88_), .Y(men_men_n1036_));
  NOi21      u1008(.An(men_men_n1036_), .B(men_men_n1034_), .Y(men_men_n1037_));
  OR4        u1009(.A(men_men_n1037_), .B(men_men_n1033_), .C(men_men_n1029_), .D(men_men_n1025_), .Y(men_men_n1038_));
  NA3        u1010(.A(men_men_n464_), .B(men_men_n336_), .C(men_men_n56_), .Y(men_men_n1039_));
  NO2        u1011(.A(men_men_n1039_), .B(men_men_n1028_), .Y(men_men_n1040_));
  NO3        u1012(.A(men_men_n1039_), .B(men_men_n578_), .C(men_men_n450_), .Y(men_men_n1041_));
  NO2        u1013(.A(f), .B(c), .Y(men_men_n1042_));
  NOi21      u1014(.An(men_men_n1042_), .B(men_men_n442_), .Y(men_men_n1043_));
  NA2        u1015(.A(men_men_n1043_), .B(men_men_n59_), .Y(men_men_n1044_));
  NO3        u1016(.A(i), .B(men_men_n246_), .C(l), .Y(men_men_n1045_));
  NOi31      u1017(.An(men_men_n1045_), .B(men_men_n1044_), .C(j), .Y(men_men_n1046_));
  OR3        u1018(.A(men_men_n1046_), .B(men_men_n1041_), .C(men_men_n1040_), .Y(men_men_n1047_));
  OR3        u1019(.A(men_men_n1047_), .B(men_men_n1038_), .C(men_men_n1020_), .Y(men02));
  OR3        u1020(.A(h), .B(u), .C(f), .Y(men_men_n1049_));
  OR3        u1021(.A(n), .B(m), .C(i), .Y(men_men_n1050_));
  NO4        u1022(.A(men_men_n1050_), .B(men_men_n1049_), .C(l), .D(men_men_n1034_), .Y(men_men_n1051_));
  NOi31      u1023(.An(e), .B(d), .C(c), .Y(men_men_n1052_));
  AOI210     u1024(.A0(men_men_n1036_), .A1(men_men_n1052_), .B0(men_men_n1012_), .Y(men_men_n1053_));
  AN3        u1025(.A(u), .B(f), .C(c), .Y(men_men_n1054_));
  NA3        u1026(.A(men_men_n1054_), .B(men_men_n464_), .C(h), .Y(men_men_n1055_));
  OR2        u1027(.A(men_men_n1035_), .B(men_men_n309_), .Y(men_men_n1056_));
  OR2        u1028(.A(men_men_n1056_), .B(men_men_n1055_), .Y(men_men_n1057_));
  NO3        u1029(.A(men_men_n1039_), .B(men_men_n1011_), .C(men_men_n578_), .Y(men_men_n1058_));
  NO2        u1030(.A(men_men_n1058_), .B(men_men_n1025_), .Y(men_men_n1059_));
  NA3        u1031(.A(l), .B(k), .C(j), .Y(men_men_n1060_));
  NA2        u1032(.A(i), .B(h), .Y(men_men_n1061_));
  NO3        u1033(.A(men_men_n1061_), .B(men_men_n1060_), .C(men_men_n132_), .Y(men_men_n1062_));
  NO3        u1034(.A(men_men_n143_), .B(men_men_n283_), .C(men_men_n215_), .Y(men_men_n1063_));
  AOI210     u1035(.A0(men_men_n1063_), .A1(men_men_n1062_), .B0(men_men_n1029_), .Y(men_men_n1064_));
  NA3        u1036(.A(c), .B(b), .C(a), .Y(men_men_n1065_));
  NO3        u1037(.A(men_men_n1065_), .B(men_men_n883_), .C(men_men_n214_), .Y(men_men_n1066_));
  NO3        u1038(.A(men_men_n1035_), .B(men_men_n301_), .C(men_men_n49_), .Y(men_men_n1067_));
  AOI210     u1039(.A0(men_men_n1067_), .A1(men_men_n1066_), .B0(men_men_n1040_), .Y(men_men_n1068_));
  AN4        u1040(.A(men_men_n1068_), .B(men_men_n1064_), .C(men_men_n1059_), .D(men_men_n1057_), .Y(men_men_n1069_));
  NO2        u1041(.A(men_men_n1015_), .B(men_men_n1013_), .Y(men_men_n1070_));
  NA2        u1042(.A(men_men_n1032_), .B(men_men_n1024_), .Y(men_men_n1071_));
  AOI210     u1043(.A0(men_men_n1071_), .A1(men_men_n1070_), .B0(men_men_n1007_), .Y(men_men_n1072_));
  NAi41      u1044(.An(men_men_n1051_), .B(men_men_n1072_), .C(men_men_n1069_), .D(men_men_n1053_), .Y(men03));
  NO2        u1045(.A(men_men_n523_), .B(men_men_n591_), .Y(men_men_n1074_));
  NA4        u1046(.A(men_men_n85_), .B(men_men_n84_), .C(u), .D(men_men_n214_), .Y(men_men_n1075_));
  NA4        u1047(.A(men_men_n566_), .B(m), .C(men_men_n111_), .D(men_men_n214_), .Y(men_men_n1076_));
  NA3        u1048(.A(men_men_n1076_), .B(men_men_n369_), .C(men_men_n1075_), .Y(men_men_n1077_));
  NO3        u1049(.A(men_men_n1077_), .B(men_men_n1074_), .C(men_men_n970_), .Y(men_men_n1078_));
  NO2        u1050(.A(men_men_n1078_), .B(men_men_n579_), .Y(men_men_n1079_));
  NOi31      u1051(.An(i), .B(k), .C(j), .Y(men_men_n1080_));
  NA4        u1052(.A(men_men_n1080_), .B(men_men_n1052_), .C(men_men_n343_), .D(men_men_n336_), .Y(men_men_n1081_));
  OAI210     u1053(.A0(men_men_n804_), .A1(men_men_n422_), .B0(men_men_n1081_), .Y(men_men_n1082_));
  NOi31      u1054(.An(m), .B(n), .C(f), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n1083_), .B(men_men_n51_), .Y(men_men_n1084_));
  AN2        u1056(.A(e), .B(c), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n1085_), .B(a), .Y(men_men_n1086_));
  OAI220     u1058(.A0(men_men_n1086_), .A1(men_men_n1084_), .B0(men_men_n869_), .B1(men_men_n427_), .Y(men_men_n1087_));
  NA2        u1059(.A(men_men_n503_), .B(l), .Y(men_men_n1088_));
  NOi31      u1060(.An(men_men_n847_), .B(men_men_n1006_), .C(men_men_n1088_), .Y(men_men_n1089_));
  NO4        u1061(.A(men_men_n1089_), .B(men_men_n1087_), .C(men_men_n1082_), .D(men_men_n969_), .Y(men_men_n1090_));
  NO2        u1062(.A(men_men_n283_), .B(a), .Y(men_men_n1091_));
  INV        u1063(.A(men_men_n1012_), .Y(men_men_n1092_));
  NO2        u1064(.A(men_men_n1061_), .B(men_men_n481_), .Y(men_men_n1093_));
  NO2        u1065(.A(men_men_n84_), .B(u), .Y(men_men_n1094_));
  AOI210     u1066(.A0(men_men_n1094_), .A1(men_men_n1093_), .B0(men_men_n1045_), .Y(men_men_n1095_));
  OR2        u1067(.A(men_men_n1095_), .B(men_men_n1044_), .Y(men_men_n1096_));
  NA3        u1068(.A(men_men_n1096_), .B(men_men_n1092_), .C(men_men_n1090_), .Y(men_men_n1097_));
  NO4        u1069(.A(men_men_n1097_), .B(men_men_n1079_), .C(men_men_n806_), .D(men_men_n559_), .Y(men_men_n1098_));
  NA2        u1070(.A(c), .B(b), .Y(men_men_n1099_));
  NO2        u1071(.A(men_men_n691_), .B(men_men_n1099_), .Y(men_men_n1100_));
  INV        u1072(.A(men_men_n415_), .Y(men_men_n1101_));
  OAI210     u1073(.A0(men_men_n1101_), .A1(men_men_n846_), .B0(men_men_n1100_), .Y(men_men_n1102_));
  NAi21      u1074(.An(men_men_n423_), .B(men_men_n1100_), .Y(men_men_n1103_));
  NA3        u1075(.A(men_men_n428_), .B(men_men_n552_), .C(f), .Y(men_men_n1104_));
  OAI210     u1076(.A0(men_men_n546_), .A1(men_men_n39_), .B0(men_men_n1091_), .Y(men_men_n1105_));
  NA3        u1077(.A(men_men_n1105_), .B(men_men_n1104_), .C(men_men_n1103_), .Y(men_men_n1106_));
  OAI210     u1078(.A0(k), .A1(men_men_n287_), .B0(u), .Y(men_men_n1107_));
  NAi21      u1079(.An(f), .B(d), .Y(men_men_n1108_));
  NO2        u1080(.A(men_men_n1108_), .B(men_men_n1065_), .Y(men_men_n1109_));
  INV        u1081(.A(men_men_n1109_), .Y(men_men_n1110_));
  NO2        u1082(.A(men_men_n1107_), .B(men_men_n1110_), .Y(men_men_n1111_));
  AOI210     u1083(.A0(men_men_n1111_), .A1(men_men_n112_), .B0(men_men_n1106_), .Y(men_men_n1112_));
  INV        u1084(.A(men_men_n466_), .Y(men_men_n1113_));
  NO2        u1085(.A(men_men_n184_), .B(men_men_n239_), .Y(men_men_n1114_));
  NA2        u1086(.A(men_men_n1114_), .B(m), .Y(men_men_n1115_));
  NA3        u1087(.A(men_men_n900_), .B(men_men_n1088_), .C(men_men_n469_), .Y(men_men_n1116_));
  OAI210     u1088(.A0(men_men_n1116_), .A1(men_men_n312_), .B0(men_men_n467_), .Y(men_men_n1117_));
  AOI210     u1089(.A0(men_men_n1117_), .A1(men_men_n1113_), .B0(men_men_n1115_), .Y(men_men_n1118_));
  NA2        u1090(.A(men_men_n554_), .B(men_men_n410_), .Y(men_men_n1119_));
  NA2        u1091(.A(men_men_n160_), .B(men_men_n33_), .Y(men_men_n1120_));
  AOI210     u1092(.A0(men_men_n941_), .A1(men_men_n1120_), .B0(men_men_n215_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n1121_), .B(men_men_n1109_), .Y(men_men_n1122_));
  NO2        u1094(.A(men_men_n372_), .B(men_men_n371_), .Y(men_men_n1123_));
  AOI210     u1095(.A0(men_men_n1114_), .A1(men_men_n430_), .B0(men_men_n938_), .Y(men_men_n1124_));
  NAi41      u1096(.An(men_men_n1123_), .B(men_men_n1124_), .C(men_men_n1122_), .D(men_men_n1119_), .Y(men_men_n1125_));
  NO2        u1097(.A(men_men_n1125_), .B(men_men_n1118_), .Y(men_men_n1126_));
  NA4        u1098(.A(men_men_n1126_), .B(men_men_n1112_), .C(men_men_n1102_), .D(men_men_n1098_), .Y(men00));
  NO2        u1099(.A(men_men_n300_), .B(men_men_n276_), .Y(men_men_n1128_));
  NO2        u1100(.A(men_men_n1128_), .B(men_men_n569_), .Y(men_men_n1129_));
  AOI210     u1101(.A0(men_men_n880_), .A1(men_men_n925_), .B0(men_men_n1082_), .Y(men_men_n1130_));
  NO3        u1102(.A(men_men_n1058_), .B(men_men_n938_), .C(men_men_n701_), .Y(men_men_n1131_));
  NA3        u1103(.A(men_men_n1131_), .B(men_men_n1130_), .C(men_men_n971_), .Y(men_men_n1132_));
  NA2        u1104(.A(men_men_n505_), .B(f), .Y(men_men_n1133_));
  NO2        u1105(.A(men_men_n1133_), .B(men_men_n1015_), .Y(men_men_n1134_));
  NO4        u1106(.A(men_men_n1134_), .B(men_men_n1132_), .C(men_men_n1129_), .D(men_men_n1038_), .Y(men_men_n1135_));
  NA2        u1107(.A(men_men_n169_), .B(men_men_n46_), .Y(men_men_n1136_));
  NA3        u1108(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1137_));
  NOi31      u1109(.An(n), .B(m), .C(i), .Y(men_men_n1138_));
  NA3        u1110(.A(men_men_n1138_), .B(men_men_n639_), .C(men_men_n51_), .Y(men_men_n1139_));
  OAI210     u1111(.A0(men_men_n1137_), .A1(men_men_n1136_), .B0(men_men_n1139_), .Y(men_men_n1140_));
  INV        u1112(.A(men_men_n568_), .Y(men_men_n1141_));
  NO4        u1113(.A(men_men_n1141_), .B(men_men_n1140_), .C(men_men_n1123_), .D(men_men_n903_), .Y(men_men_n1142_));
  NO4        u1114(.A(men_men_n484_), .B(men_men_n356_), .C(men_men_n1099_), .D(men_men_n59_), .Y(men_men_n1143_));
  OR2        u1115(.A(men_men_n385_), .B(men_men_n135_), .Y(men_men_n1144_));
  NO2        u1116(.A(h), .B(u), .Y(men_men_n1145_));
  NA4        u1117(.A(men_men_n494_), .B(men_men_n464_), .C(men_men_n1145_), .D(men_men_n1005_), .Y(men_men_n1146_));
  OAI220     u1118(.A0(men_men_n523_), .A1(men_men_n591_), .B0(men_men_n89_), .B1(men_men_n88_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n1147_), .B(men_men_n532_), .Y(men_men_n1148_));
  AOI220     u1120(.A0(men_men_n319_), .A1(men_men_n249_), .B0(men_men_n179_), .B1(men_men_n149_), .Y(men_men_n1149_));
  NA4        u1121(.A(men_men_n1149_), .B(men_men_n1148_), .C(men_men_n1146_), .D(men_men_n1144_), .Y(men_men_n1150_));
  NO3        u1122(.A(men_men_n1150_), .B(men_men_n1143_), .C(men_men_n268_), .Y(men_men_n1151_));
  INV        u1123(.A(men_men_n324_), .Y(men_men_n1152_));
  AOI210     u1124(.A0(men_men_n249_), .A1(men_men_n348_), .B0(men_men_n570_), .Y(men_men_n1153_));
  NA3        u1125(.A(men_men_n1153_), .B(men_men_n1152_), .C(men_men_n155_), .Y(men_men_n1154_));
  NO2        u1126(.A(men_men_n241_), .B(men_men_n183_), .Y(men_men_n1155_));
  NA2        u1127(.A(men_men_n1155_), .B(men_men_n428_), .Y(men_men_n1156_));
  NA3        u1128(.A(men_men_n181_), .B(men_men_n111_), .C(u), .Y(men_men_n1157_));
  NA3        u1129(.A(men_men_n464_), .B(men_men_n40_), .C(f), .Y(men_men_n1158_));
  NOi31      u1130(.An(men_men_n855_), .B(men_men_n1158_), .C(men_men_n1157_), .Y(men_men_n1159_));
  NAi31      u1131(.An(men_men_n185_), .B(men_men_n843_), .C(men_men_n464_), .Y(men_men_n1160_));
  NAi31      u1132(.An(men_men_n1159_), .B(men_men_n1160_), .C(men_men_n1156_), .Y(men_men_n1161_));
  NO2        u1133(.A(men_men_n275_), .B(men_men_n75_), .Y(men_men_n1162_));
  NO3        u1134(.A(men_men_n427_), .B(men_men_n817_), .C(n), .Y(men_men_n1163_));
  AOI210     u1135(.A0(men_men_n1163_), .A1(men_men_n1162_), .B0(men_men_n1051_), .Y(men_men_n1164_));
  NAi31      u1136(.An(men_men_n1018_), .B(men_men_n1164_), .C(men_men_n74_), .Y(men_men_n1165_));
  NO4        u1137(.A(men_men_n1165_), .B(men_men_n1161_), .C(men_men_n1154_), .D(men_men_n514_), .Y(men_men_n1166_));
  AN3        u1138(.A(men_men_n1166_), .B(men_men_n1151_), .C(men_men_n1142_), .Y(men_men_n1167_));
  NA2        u1139(.A(men_men_n532_), .B(men_men_n99_), .Y(men_men_n1168_));
  NA3        u1140(.A(men_men_n1083_), .B(men_men_n599_), .C(men_men_n463_), .Y(men_men_n1169_));
  NA4        u1141(.A(men_men_n1169_), .B(men_men_n555_), .C(men_men_n1168_), .D(men_men_n244_), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n1077_), .B(men_men_n532_), .Y(men_men_n1171_));
  NA4        u1143(.A(men_men_n639_), .B(men_men_n206_), .C(men_men_n222_), .D(men_men_n164_), .Y(men_men_n1172_));
  NA3        u1144(.A(men_men_n1172_), .B(men_men_n1171_), .C(men_men_n297_), .Y(men_men_n1173_));
  OAI210     u1145(.A0(men_men_n462_), .A1(men_men_n119_), .B0(men_men_n848_), .Y(men_men_n1174_));
  AOI220     u1146(.A0(men_men_n1174_), .A1(men_men_n1116_), .B0(men_men_n554_), .B1(men_men_n410_), .Y(men_men_n1175_));
  OR3        u1147(.A(men_men_n1015_), .B(men_men_n273_), .C(men_men_n224_), .Y(men_men_n1176_));
  NA2        u1148(.A(men_men_n1176_), .B(men_men_n1175_), .Y(men_men_n1177_));
  INV        u1149(.A(men_men_n805_), .Y(men_men_n1178_));
  AOI220     u1150(.A0(men_men_n934_), .A1(men_men_n567_), .B0(men_men_n639_), .B1(men_men_n247_), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n68_), .B(h), .Y(men_men_n1180_));
  NO3        u1152(.A(men_men_n1015_), .B(men_men_n1013_), .C(men_men_n718_), .Y(men_men_n1181_));
  INV        u1153(.A(men_men_n132_), .Y(men_men_n1182_));
  AN2        u1154(.A(men_men_n1182_), .B(men_men_n1063_), .Y(men_men_n1183_));
  OAI210     u1155(.A0(men_men_n1183_), .A1(men_men_n1181_), .B0(men_men_n1180_), .Y(men_men_n1184_));
  NA4        u1156(.A(men_men_n1184_), .B(men_men_n1179_), .C(men_men_n1178_), .D(men_men_n850_), .Y(men_men_n1185_));
  NO4        u1157(.A(men_men_n1185_), .B(men_men_n1177_), .C(men_men_n1173_), .D(men_men_n1170_), .Y(men_men_n1186_));
  NA2        u1158(.A(men_men_n822_), .B(men_men_n750_), .Y(men_men_n1187_));
  NA4        u1159(.A(men_men_n1187_), .B(men_men_n1186_), .C(men_men_n1167_), .D(men_men_n1135_), .Y(men01));
  NO3        u1160(.A(men_men_n788_), .B(men_men_n782_), .C(men_men_n281_), .Y(men_men_n1189_));
  NA2        u1161(.A(men_men_n395_), .B(i), .Y(men_men_n1190_));
  NA3        u1162(.A(men_men_n1190_), .B(men_men_n1189_), .C(men_men_n994_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n580_), .B(men_men_n87_), .Y(men_men_n1192_));
  NA3        u1164(.A(men_men_n1192_), .B(men_men_n896_), .C(men_men_n335_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n698_), .B(men_men_n94_), .Y(men_men_n1194_));
  NO2        u1166(.A(men_men_n1194_), .B(i), .Y(men_men_n1195_));
  OAI210     u1167(.A0(men_men_n769_), .A1(men_men_n594_), .B0(men_men_n1172_), .Y(men_men_n1196_));
  AOI210     u1168(.A0(men_men_n1195_), .A1(men_men_n627_), .B0(men_men_n1196_), .Y(men_men_n1197_));
  INV        u1169(.A(men_men_n117_), .Y(men_men_n1198_));
  OA220      u1170(.A0(men_men_n1198_), .A1(men_men_n577_), .B0(men_men_n652_), .B1(men_men_n369_), .Y(men_men_n1199_));
  NAi41      u1171(.An(men_men_n163_), .B(men_men_n1199_), .C(men_men_n1197_), .D(men_men_n879_), .Y(men_men_n1200_));
  NO2        u1172(.A(men_men_n667_), .B(men_men_n508_), .Y(men_men_n1201_));
  NA3        u1173(.A(men_men_n698_), .B(men_men_n94_), .C(men_men_n214_), .Y(men_men_n1202_));
  OR2        u1174(.A(men_men_n195_), .B(men_men_n193_), .Y(men_men_n1203_));
  NA3        u1175(.A(men_men_n1203_), .B(men_men_n1201_), .C(men_men_n138_), .Y(men_men_n1204_));
  NO4        u1176(.A(men_men_n1204_), .B(men_men_n1200_), .C(men_men_n1193_), .D(men_men_n1191_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n303_), .B(men_men_n527_), .Y(men_men_n1206_));
  NA2        u1178(.A(men_men_n535_), .B(men_men_n397_), .Y(men_men_n1207_));
  NOi21      u1179(.An(men_men_n556_), .B(men_men_n574_), .Y(men_men_n1208_));
  NA2        u1180(.A(men_men_n1208_), .B(men_men_n1207_), .Y(men_men_n1209_));
  AN3        u1181(.A(m), .B(l), .C(k), .Y(men_men_n1210_));
  OAI210     u1182(.A0(men_men_n357_), .A1(men_men_n34_), .B0(men_men_n1210_), .Y(men_men_n1211_));
  NA2        u1183(.A(men_men_n203_), .B(men_men_n34_), .Y(men_men_n1212_));
  AO210      u1184(.A0(men_men_n1212_), .A1(men_men_n1211_), .B0(men_men_n334_), .Y(men_men_n1213_));
  NA3        u1185(.A(men_men_n1213_), .B(men_men_n1209_), .C(men_men_n1206_), .Y(men_men_n1214_));
  NA2        u1186(.A(men_men_n589_), .B(men_men_n117_), .Y(men_men_n1215_));
  OAI210     u1187(.A0(men_men_n1198_), .A1(men_men_n586_), .B0(men_men_n1215_), .Y(men_men_n1216_));
  NA2        u1188(.A(men_men_n280_), .B(men_men_n195_), .Y(men_men_n1217_));
  NA2        u1189(.A(men_men_n1217_), .B(men_men_n657_), .Y(men_men_n1218_));
  NO3        u1190(.A(men_men_n804_), .B(men_men_n204_), .C(men_men_n408_), .Y(men_men_n1219_));
  NO2        u1191(.A(men_men_n1219_), .B(men_men_n938_), .Y(men_men_n1220_));
  NA3        u1192(.A(men_men_n1220_), .B(men_men_n1218_), .C(men_men_n772_), .Y(men_men_n1221_));
  NO3        u1193(.A(men_men_n1221_), .B(men_men_n1216_), .C(men_men_n1214_), .Y(men_men_n1222_));
  NA3        u1194(.A(men_men_n595_), .B(men_men_n29_), .C(f), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n1223_), .B(men_men_n204_), .Y(men_men_n1224_));
  AOI210     u1196(.A0(men_men_n500_), .A1(men_men_n58_), .B0(men_men_n1224_), .Y(men_men_n1225_));
  OR3        u1197(.A(men_men_n1194_), .B(men_men_n596_), .C(i), .Y(men_men_n1226_));
  NO2        u1198(.A(men_men_n1202_), .B(men_men_n951_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n207_), .B(men_men_n110_), .Y(men_men_n1228_));
  NO3        u1200(.A(men_men_n1228_), .B(men_men_n1227_), .C(men_men_n1140_), .Y(men_men_n1229_));
  NA4        u1201(.A(men_men_n1229_), .B(men_men_n1226_), .C(men_men_n1225_), .D(men_men_n749_), .Y(men_men_n1230_));
  NO2        u1202(.A(men_men_n944_), .B(men_men_n234_), .Y(men_men_n1231_));
  NO2        u1203(.A(men_men_n945_), .B(men_men_n551_), .Y(men_men_n1232_));
  OAI210     u1204(.A0(men_men_n1232_), .A1(men_men_n1231_), .B0(men_men_n341_), .Y(men_men_n1233_));
  INV        u1205(.A(men_men_n662_), .Y(men_men_n1234_));
  NO2        u1206(.A(men_men_n369_), .B(men_men_n73_), .Y(men_men_n1235_));
  INV        u1207(.A(men_men_n1235_), .Y(men_men_n1236_));
  NA2        u1208(.A(men_men_n1236_), .B(men_men_n387_), .Y(men_men_n1237_));
  NOi41      u1209(.An(men_men_n1233_), .B(men_men_n1237_), .C(men_men_n1234_), .D(men_men_n1230_), .Y(men_men_n1238_));
  NO2        u1210(.A(men_men_n131_), .B(men_men_n45_), .Y(men_men_n1239_));
  NO2        u1211(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1240_));
  AO220      u1212(.A0(men_men_n1240_), .A1(men_men_n615_), .B0(men_men_n1239_), .B1(men_men_n696_), .Y(men_men_n1241_));
  NA2        u1213(.A(men_men_n1241_), .B(men_men_n341_), .Y(men_men_n1242_));
  INV        u1214(.A(men_men_n135_), .Y(men_men_n1243_));
  NO3        u1215(.A(men_men_n1061_), .B(men_men_n178_), .C(men_men_n84_), .Y(men_men_n1244_));
  NA2        u1216(.A(men_men_n1244_), .B(men_men_n1243_), .Y(men_men_n1245_));
  NA2        u1217(.A(men_men_n1245_), .B(men_men_n1242_), .Y(men_men_n1246_));
  NO2        u1218(.A(men_men_n607_), .B(men_men_n606_), .Y(men_men_n1247_));
  NO4        u1219(.A(men_men_n1061_), .B(men_men_n1247_), .C(men_men_n176_), .D(men_men_n84_), .Y(men_men_n1248_));
  NO3        u1220(.A(men_men_n1248_), .B(men_men_n1246_), .C(men_men_n630_), .Y(men_men_n1249_));
  NA4        u1221(.A(men_men_n1249_), .B(men_men_n1238_), .C(men_men_n1222_), .D(men_men_n1205_), .Y(men06));
  NO2        u1222(.A(men_men_n409_), .B(men_men_n553_), .Y(men_men_n1251_));
  NA2        u1223(.A(men_men_n269_), .B(men_men_n1251_), .Y(men_men_n1252_));
  NO2        u1224(.A(men_men_n226_), .B(men_men_n101_), .Y(men_men_n1253_));
  OAI210     u1225(.A0(men_men_n1253_), .A1(men_men_n1244_), .B0(men_men_n383_), .Y(men_men_n1254_));
  NO3        u1226(.A(men_men_n592_), .B(men_men_n793_), .C(men_men_n593_), .Y(men_men_n1255_));
  OR2        u1227(.A(men_men_n1255_), .B(men_men_n869_), .Y(men_men_n1256_));
  NA4        u1228(.A(men_men_n1256_), .B(men_men_n1254_), .C(men_men_n1252_), .D(men_men_n1233_), .Y(men_men_n1257_));
  NO3        u1229(.A(men_men_n1257_), .B(men_men_n1234_), .C(men_men_n259_), .Y(men_men_n1258_));
  INV        u1230(.A(men_men_n1231_), .Y(men_men_n1259_));
  INV        u1231(.A(men_men_n1241_), .Y(men_men_n1260_));
  AOI210     u1232(.A0(men_men_n1260_), .A1(men_men_n1259_), .B0(men_men_n338_), .Y(men_men_n1261_));
  OAI210     u1233(.A0(men_men_n86_), .A1(men_men_n40_), .B0(men_men_n666_), .Y(men_men_n1262_));
  NA2        u1234(.A(men_men_n1262_), .B(men_men_n634_), .Y(men_men_n1263_));
  NO2        u1235(.A(men_men_n511_), .B(men_men_n173_), .Y(men_men_n1264_));
  NOi21      u1236(.An(men_men_n137_), .B(men_men_n45_), .Y(men_men_n1265_));
  NO2        u1237(.A(men_men_n600_), .B(men_men_n1084_), .Y(men_men_n1266_));
  OAI210     u1238(.A0(men_men_n459_), .A1(men_men_n250_), .B0(men_men_n890_), .Y(men_men_n1267_));
  NO4        u1239(.A(men_men_n1267_), .B(men_men_n1266_), .C(men_men_n1265_), .D(men_men_n1264_), .Y(men_men_n1268_));
  NO2        u1240(.A(men_men_n368_), .B(men_men_n136_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n580_), .Y(men_men_n1270_));
  NA3        u1242(.A(men_men_n1270_), .B(men_men_n1268_), .C(men_men_n1263_), .Y(men_men_n1271_));
  NO2        u1243(.A(men_men_n740_), .B(men_men_n367_), .Y(men_men_n1272_));
  NO2        u1244(.A(men_men_n751_), .B(men_men_n627_), .Y(men_men_n1273_));
  NOi21      u1245(.An(men_men_n1272_), .B(men_men_n1273_), .Y(men_men_n1274_));
  NO3        u1246(.A(men_men_n1274_), .B(men_men_n1271_), .C(men_men_n1261_), .Y(men_men_n1275_));
  NO2        u1247(.A(men_men_n787_), .B(men_men_n277_), .Y(men_men_n1276_));
  OAI220     u1248(.A0(men_men_n725_), .A1(men_men_n47_), .B0(men_men_n226_), .B1(men_men_n609_), .Y(men_men_n1277_));
  OAI210     u1249(.A0(men_men_n277_), .A1(c), .B0(men_men_n633_), .Y(men_men_n1278_));
  AOI220     u1250(.A0(men_men_n1278_), .A1(men_men_n1277_), .B0(men_men_n1276_), .B1(men_men_n269_), .Y(men_men_n1279_));
  NO3        u1251(.A(men_men_n246_), .B(men_men_n101_), .C(men_men_n283_), .Y(men_men_n1280_));
  OAI220     u1252(.A0(men_men_n688_), .A1(men_men_n250_), .B0(men_men_n507_), .B1(men_men_n511_), .Y(men_men_n1281_));
  OAI210     u1253(.A0(l), .A1(i), .B0(k), .Y(men_men_n1282_));
  NO3        u1254(.A(men_men_n1282_), .B(men_men_n591_), .C(j), .Y(men_men_n1283_));
  NOi21      u1255(.An(men_men_n1283_), .B(men_men_n660_), .Y(men_men_n1284_));
  NO4        u1256(.A(men_men_n1284_), .B(men_men_n1281_), .C(men_men_n1280_), .D(men_men_n1087_), .Y(men_men_n1285_));
  NA4        u1257(.A(men_men_n780_), .B(men_men_n779_), .C(men_men_n438_), .D(men_men_n861_), .Y(men_men_n1286_));
  NAi31      u1258(.An(men_men_n740_), .B(men_men_n1286_), .C(men_men_n203_), .Y(men_men_n1287_));
  NA4        u1259(.A(men_men_n1287_), .B(men_men_n1285_), .C(men_men_n1279_), .D(men_men_n1179_), .Y(men_men_n1288_));
  OR3        u1260(.A(men_men_n1497_), .B(men_men_n769_), .C(men_men_n538_), .Y(men_men_n1289_));
  OR3        u1261(.A(men_men_n371_), .B(men_men_n226_), .C(men_men_n609_), .Y(men_men_n1290_));
  AOI210     u1262(.A0(men_men_n564_), .A1(men_men_n448_), .B0(men_men_n373_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n1283_), .B(men_men_n776_), .Y(men_men_n1292_));
  NA4        u1264(.A(men_men_n1292_), .B(men_men_n1291_), .C(men_men_n1290_), .D(men_men_n1289_), .Y(men_men_n1293_));
  AOI220     u1265(.A0(men_men_n1272_), .A1(men_men_n750_), .B0(men_men_n1269_), .B1(men_men_n240_), .Y(men_men_n1294_));
  NO3        u1266(.A(men_men_n859_), .B(men_men_n496_), .C(men_men_n478_), .Y(men_men_n1295_));
  NA2        u1267(.A(men_men_n1295_), .B(men_men_n1294_), .Y(men_men_n1296_));
  NAi21      u1268(.An(j), .B(i), .Y(men_men_n1297_));
  NO4        u1269(.A(men_men_n1247_), .B(men_men_n1297_), .C(men_men_n442_), .D(men_men_n237_), .Y(men_men_n1298_));
  NO4        u1270(.A(men_men_n1298_), .B(men_men_n1296_), .C(men_men_n1293_), .D(men_men_n1288_), .Y(men_men_n1299_));
  NA4        u1271(.A(men_men_n1299_), .B(men_men_n1275_), .C(men_men_n1258_), .D(men_men_n1249_), .Y(men07));
  NAi32      u1272(.An(m), .Bn(b), .C(n), .Y(men_men_n1301_));
  NO3        u1273(.A(men_men_n1301_), .B(u), .C(f), .Y(men_men_n1302_));
  OAI210     u1274(.A0(men_men_n323_), .A1(men_men_n480_), .B0(men_men_n1302_), .Y(men_men_n1303_));
  OR2        u1275(.A(e), .B(d), .Y(men_men_n1304_));
  NOi31      u1276(.An(n), .B(m), .C(b), .Y(men_men_n1305_));
  NO3        u1277(.A(men_men_n132_), .B(men_men_n450_), .C(h), .Y(men_men_n1306_));
  INV        u1278(.A(men_men_n1303_), .Y(men_men_n1307_));
  NOi41      u1279(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1308_));
  NA3        u1280(.A(men_men_n1308_), .B(men_men_n852_), .C(men_men_n411_), .Y(men_men_n1309_));
  NO2        u1281(.A(men_men_n1309_), .B(men_men_n56_), .Y(men_men_n1310_));
  NA2        u1282(.A(men_men_n1063_), .B(men_men_n222_), .Y(men_men_n1311_));
  NO2        u1283(.A(men_men_n1311_), .B(men_men_n61_), .Y(men_men_n1312_));
  NO2        u1284(.A(k), .B(i), .Y(men_men_n1313_));
  NA3        u1285(.A(men_men_n1313_), .B(men_men_n878_), .C(men_men_n181_), .Y(men_men_n1314_));
  NA2        u1286(.A(men_men_n84_), .B(men_men_n45_), .Y(men_men_n1315_));
  NO2        u1287(.A(men_men_n1021_), .B(men_men_n442_), .Y(men_men_n1316_));
  NA3        u1288(.A(men_men_n1316_), .B(men_men_n1315_), .C(men_men_n215_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n1035_), .B(men_men_n309_), .Y(men_men_n1318_));
  NA2        u1290(.A(men_men_n1180_), .B(men_men_n291_), .Y(men_men_n1319_));
  NA3        u1291(.A(men_men_n1319_), .B(men_men_n1317_), .C(men_men_n1314_), .Y(men_men_n1320_));
  NO4        u1292(.A(men_men_n1320_), .B(men_men_n1312_), .C(men_men_n1310_), .D(men_men_n1307_), .Y(men_men_n1321_));
  NO3        u1293(.A(e), .B(d), .C(c), .Y(men_men_n1322_));
  OAI210     u1294(.A0(men_men_n132_), .A1(men_men_n215_), .B0(men_men_n597_), .Y(men_men_n1323_));
  NA2        u1295(.A(men_men_n1323_), .B(men_men_n1322_), .Y(men_men_n1324_));
  INV        u1296(.A(men_men_n1324_), .Y(men_men_n1325_));
  OR2        u1297(.A(h), .B(f), .Y(men_men_n1326_));
  NO3        u1298(.A(n), .B(m), .C(i), .Y(men_men_n1327_));
  OAI210     u1299(.A0(men_men_n1085_), .A1(men_men_n158_), .B0(men_men_n1327_), .Y(men_men_n1328_));
  NO2        u1300(.A(i), .B(u), .Y(men_men_n1329_));
  OR3        u1301(.A(men_men_n1329_), .B(men_men_n1301_), .C(men_men_n72_), .Y(men_men_n1330_));
  OAI220     u1302(.A0(men_men_n1330_), .A1(men_men_n480_), .B0(men_men_n1328_), .B1(men_men_n1326_), .Y(men_men_n1331_));
  NA3        u1303(.A(men_men_n685_), .B(men_men_n674_), .C(men_men_n111_), .Y(men_men_n1332_));
  NA3        u1304(.A(men_men_n1305_), .B(men_men_n1030_), .C(men_men_n664_), .Y(men_men_n1333_));
  AOI210     u1305(.A0(men_men_n1333_), .A1(men_men_n1332_), .B0(men_men_n45_), .Y(men_men_n1334_));
  NO2        u1306(.A(l), .B(k), .Y(men_men_n1335_));
  NOi41      u1307(.An(men_men_n544_), .B(men_men_n1335_), .C(men_men_n475_), .D(men_men_n442_), .Y(men_men_n1336_));
  NO3        u1308(.A(men_men_n442_), .B(d), .C(c), .Y(men_men_n1337_));
  NO4        u1309(.A(men_men_n1336_), .B(men_men_n1334_), .C(men_men_n1331_), .D(men_men_n1325_), .Y(men_men_n1338_));
  NO2        u1310(.A(men_men_n148_), .B(h), .Y(men_men_n1339_));
  NO2        u1311(.A(i), .B(l), .Y(men_men_n1340_));
  NO2        u1312(.A(u), .B(c), .Y(men_men_n1341_));
  NA3        u1313(.A(men_men_n1341_), .B(men_men_n143_), .C(men_men_n186_), .Y(men_men_n1342_));
  NO2        u1314(.A(men_men_n1342_), .B(men_men_n1340_), .Y(men_men_n1343_));
  NA2        u1315(.A(men_men_n1343_), .B(men_men_n181_), .Y(men_men_n1344_));
  NO2        u1316(.A(men_men_n452_), .B(a), .Y(men_men_n1345_));
  NA3        u1317(.A(men_men_n1345_), .B(k), .C(men_men_n112_), .Y(men_men_n1346_));
  NO2        u1318(.A(i), .B(h), .Y(men_men_n1347_));
  NA2        u1319(.A(men_men_n1347_), .B(men_men_n222_), .Y(men_men_n1348_));
  NA2        u1320(.A(men_men_n1108_), .B(h), .Y(men_men_n1349_));
  NA2        u1321(.A(men_men_n139_), .B(men_men_n222_), .Y(men_men_n1350_));
  AOI210     u1322(.A0(men_men_n260_), .A1(men_men_n115_), .B0(men_men_n527_), .Y(men_men_n1351_));
  OAI220     u1323(.A0(men_men_n1351_), .A1(men_men_n1348_), .B0(men_men_n1350_), .B1(men_men_n1349_), .Y(men_men_n1352_));
  NO2        u1324(.A(men_men_n747_), .B(men_men_n187_), .Y(men_men_n1353_));
  NOi31      u1325(.An(m), .B(n), .C(b), .Y(men_men_n1354_));
  NOi31      u1326(.An(f), .B(d), .C(c), .Y(men_men_n1355_));
  NA2        u1327(.A(men_men_n1355_), .B(men_men_n1354_), .Y(men_men_n1356_));
  INV        u1328(.A(men_men_n1356_), .Y(men_men_n1357_));
  NO3        u1329(.A(men_men_n1357_), .B(men_men_n1353_), .C(men_men_n1352_), .Y(men_men_n1358_));
  NA2        u1330(.A(men_men_n1054_), .B(men_men_n464_), .Y(men_men_n1359_));
  OAI210     u1331(.A0(men_men_n184_), .A1(men_men_n522_), .B0(men_men_n1031_), .Y(men_men_n1360_));
  NO3        u1332(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1361_));
  AN4        u1333(.A(men_men_n1360_), .B(men_men_n1358_), .C(men_men_n1346_), .D(men_men_n1344_), .Y(men_men_n1362_));
  NA2        u1334(.A(men_men_n1305_), .B(men_men_n380_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n187_), .B(b), .Y(men_men_n1364_));
  NA2        u1336(.A(men_men_n1062_), .B(men_men_n1359_), .Y(men_men_n1365_));
  NO2        u1337(.A(i), .B(men_men_n214_), .Y(men_men_n1366_));
  NA4        u1338(.A(men_men_n1114_), .B(men_men_n1366_), .C(men_men_n102_), .D(m), .Y(men_men_n1367_));
  NA2        u1339(.A(men_men_n1367_), .B(men_men_n1365_), .Y(men_men_n1368_));
  NO4        u1340(.A(men_men_n132_), .B(u), .C(f), .D(e), .Y(men_men_n1369_));
  NA3        u1341(.A(men_men_n1313_), .B(men_men_n292_), .C(h), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n194_), .B(men_men_n96_), .Y(men_men_n1371_));
  NA2        u1343(.A(men_men_n30_), .B(h), .Y(men_men_n1372_));
  NO2        u1344(.A(men_men_n1372_), .B(men_men_n1050_), .Y(men_men_n1373_));
  NOi41      u1345(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1374_));
  NA2        u1346(.A(men_men_n1374_), .B(men_men_n112_), .Y(men_men_n1375_));
  INV        u1347(.A(men_men_n1375_), .Y(men_men_n1376_));
  OR3        u1348(.A(men_men_n538_), .B(men_men_n537_), .C(men_men_n111_), .Y(men_men_n1377_));
  NA2        u1349(.A(men_men_n1083_), .B(men_men_n408_), .Y(men_men_n1378_));
  OAI220     u1350(.A0(men_men_n1378_), .A1(men_men_n437_), .B0(men_men_n1377_), .B1(men_men_n301_), .Y(men_men_n1379_));
  AO210      u1351(.A0(men_men_n1379_), .A1(men_men_n115_), .B0(men_men_n1376_), .Y(men_men_n1380_));
  NO3        u1352(.A(men_men_n1380_), .B(men_men_n1373_), .C(men_men_n1368_), .Y(men_men_n1381_));
  NA4        u1353(.A(men_men_n1381_), .B(men_men_n1362_), .C(men_men_n1338_), .D(men_men_n1321_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n1099_), .B(men_men_n109_), .Y(men_men_n1383_));
  NA2        u1355(.A(men_men_n380_), .B(men_men_n56_), .Y(men_men_n1384_));
  NA2        u1356(.A(men_men_n216_), .B(men_men_n181_), .Y(men_men_n1385_));
  AOI210     u1357(.A0(men_men_n1385_), .A1(men_men_n1157_), .B0(men_men_n1384_), .Y(men_men_n1386_));
  NO2        u1358(.A(men_men_n392_), .B(j), .Y(men_men_n1387_));
  NA3        u1359(.A(men_men_n1361_), .B(men_men_n1304_), .C(men_men_n1083_), .Y(men_men_n1388_));
  INV        u1360(.A(men_men_n1388_), .Y(men_men_n1389_));
  NA3        u1361(.A(u), .B(men_men_n1387_), .C(men_men_n160_), .Y(men_men_n1390_));
  INV        u1362(.A(men_men_n1390_), .Y(men_men_n1391_));
  NO3        u1363(.A(men_men_n740_), .B(men_men_n176_), .C(men_men_n411_), .Y(men_men_n1392_));
  NO3        u1364(.A(men_men_n1392_), .B(men_men_n1391_), .C(men_men_n1389_), .Y(men_men_n1393_));
  NO3        u1365(.A(men_men_n1050_), .B(men_men_n574_), .C(u), .Y(men_men_n1394_));
  NOi21      u1366(.An(men_men_n1385_), .B(men_men_n1394_), .Y(men_men_n1395_));
  AOI210     u1367(.A0(men_men_n1395_), .A1(men_men_n1371_), .B0(men_men_n1021_), .Y(men_men_n1396_));
  OR2        u1368(.A(n), .B(i), .Y(men_men_n1397_));
  OAI210     u1369(.A0(men_men_n1397_), .A1(men_men_n1042_), .B0(men_men_n49_), .Y(men_men_n1398_));
  AOI220     u1370(.A0(men_men_n1398_), .A1(men_men_n1145_), .B0(men_men_n809_), .B1(men_men_n194_), .Y(men_men_n1399_));
  INV        u1371(.A(men_men_n1399_), .Y(men_men_n1400_));
  NA2        u1372(.A(men_men_n1364_), .B(men_men_n41_), .Y(men_men_n1401_));
  NO2        u1373(.A(men_men_n1401_), .B(men_men_n178_), .Y(men_men_n1402_));
  NO3        u1374(.A(men_men_n1402_), .B(men_men_n1400_), .C(men_men_n1396_), .Y(men_men_n1403_));
  INV        u1375(.A(men_men_n49_), .Y(men_men_n1404_));
  NO3        u1376(.A(men_men_n1065_), .B(men_men_n1304_), .C(men_men_n49_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1066_), .B(men_men_n1404_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1050_), .B(h), .Y(men_men_n1407_));
  NA3        u1379(.A(men_men_n1407_), .B(d), .C(men_men_n1013_), .Y(men_men_n1408_));
  OAI220     u1380(.A0(men_men_n1408_), .A1(c), .B0(men_men_n1406_), .B1(j), .Y(men_men_n1409_));
  NA3        u1381(.A(men_men_n1383_), .B(men_men_n464_), .C(f), .Y(men_men_n1410_));
  NO2        u1382(.A(j), .B(men_men_n42_), .Y(men_men_n1411_));
  NA2        u1383(.A(men_men_n112_), .B(men_men_n40_), .Y(men_men_n1412_));
  NO2        u1384(.A(men_men_n1412_), .B(men_men_n1410_), .Y(men_men_n1413_));
  AOI210     u1385(.A0(men_men_n522_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1414_));
  NA2        u1386(.A(men_men_n1414_), .B(men_men_n1345_), .Y(men_men_n1415_));
  NO2        u1387(.A(men_men_n1297_), .B(men_men_n176_), .Y(men_men_n1416_));
  NOi21      u1388(.An(d), .B(f), .Y(men_men_n1417_));
  NO2        u1389(.A(men_men_n1355_), .B(men_men_n1417_), .Y(men_men_n1418_));
  NA2        u1390(.A(men_men_n1418_), .B(men_men_n1416_), .Y(men_men_n1419_));
  NO2        u1391(.A(men_men_n1304_), .B(f), .Y(men_men_n1420_));
  NA2        u1392(.A(men_men_n1345_), .B(men_men_n1411_), .Y(men_men_n1421_));
  NO2        u1393(.A(men_men_n301_), .B(c), .Y(men_men_n1422_));
  NA2        u1394(.A(men_men_n1422_), .B(men_men_n539_), .Y(men_men_n1423_));
  NA4        u1395(.A(men_men_n1423_), .B(men_men_n1421_), .C(men_men_n1419_), .D(men_men_n1415_), .Y(men_men_n1424_));
  NO3        u1396(.A(men_men_n1424_), .B(men_men_n1413_), .C(men_men_n1409_), .Y(men_men_n1425_));
  NA4        u1397(.A(men_men_n1425_), .B(men_men_n1403_), .C(men_men_n1393_), .D(men_men_n1496_), .Y(men_men_n1426_));
  NO3        u1398(.A(men_men_n1054_), .B(men_men_n1042_), .C(men_men_n40_), .Y(men_men_n1427_));
  NO2        u1399(.A(men_men_n464_), .B(men_men_n301_), .Y(men_men_n1428_));
  OAI210     u1400(.A0(men_men_n1428_), .A1(men_men_n1427_), .B0(men_men_n1318_), .Y(men_men_n1429_));
  OAI210     u1401(.A0(men_men_n1369_), .A1(men_men_n1305_), .B0(men_men_n866_), .Y(men_men_n1430_));
  OAI220     u1402(.A0(men_men_n1010_), .A1(men_men_n132_), .B0(h), .B1(men_men_n176_), .Y(men_men_n1431_));
  NA2        u1403(.A(men_men_n1431_), .B(men_men_n614_), .Y(men_men_n1432_));
  NA3        u1404(.A(men_men_n1432_), .B(men_men_n1430_), .C(men_men_n1429_), .Y(men_men_n1433_));
  NA2        u1405(.A(men_men_n1341_), .B(men_men_n1417_), .Y(men_men_n1434_));
  NO2        u1406(.A(men_men_n1434_), .B(m), .Y(men_men_n1435_));
  NA3        u1407(.A(men_men_n1063_), .B(men_men_n107_), .C(men_men_n222_), .Y(men_men_n1436_));
  NO2        u1408(.A(men_men_n152_), .B(men_men_n183_), .Y(men_men_n1437_));
  OAI210     u1409(.A0(men_men_n1437_), .A1(men_men_n109_), .B0(men_men_n1354_), .Y(men_men_n1438_));
  NA2        u1410(.A(men_men_n1438_), .B(men_men_n1436_), .Y(men_men_n1439_));
  NO3        u1411(.A(men_men_n1439_), .B(men_men_n1435_), .C(men_men_n1433_), .Y(men_men_n1440_));
  NO2        u1412(.A(f), .B(e), .Y(men_men_n1441_));
  OAI210     u1413(.A0(men_men_n1420_), .A1(men_men_n1094_), .B0(men_men_n623_), .Y(men_men_n1442_));
  NO2        u1414(.A(men_men_n1442_), .B(men_men_n444_), .Y(men_men_n1443_));
  NO3        u1415(.A(men_men_n1377_), .B(men_men_n355_), .C(a), .Y(men_men_n1444_));
  NO2        u1416(.A(men_men_n1444_), .B(men_men_n1443_), .Y(men_men_n1445_));
  NO2        u1417(.A(men_men_n183_), .B(c), .Y(men_men_n1446_));
  OAI210     u1418(.A0(men_men_n1446_), .A1(men_men_n1441_), .B0(men_men_n181_), .Y(men_men_n1447_));
  AOI220     u1419(.A0(men_men_n1447_), .A1(men_men_n1044_), .B0(men_men_n529_), .B1(men_men_n367_), .Y(men_men_n1448_));
  NA2        u1420(.A(men_men_n537_), .B(u), .Y(men_men_n1449_));
  AOI210     u1421(.A0(men_men_n1449_), .A1(men_men_n1337_), .B0(men_men_n1405_), .Y(men_men_n1450_));
  NO2        u1422(.A(men_men_n1450_), .B(men_men_n214_), .Y(men_men_n1451_));
  AOI210     u1423(.A0(men_men_n883_), .A1(men_men_n418_), .B0(men_men_n103_), .Y(men_men_n1452_));
  NO2        u1424(.A(men_men_n1452_), .B(men_men_n176_), .Y(men_men_n1453_));
  NA2        u1425(.A(men_men_n1306_), .B(men_men_n184_), .Y(men_men_n1454_));
  NO2        u1426(.A(men_men_n49_), .B(l), .Y(men_men_n1455_));
  INV        u1427(.A(men_men_n480_), .Y(men_men_n1456_));
  OAI210     u1428(.A0(men_men_n1456_), .A1(men_men_n1066_), .B0(men_men_n1455_), .Y(men_men_n1457_));
  NO2        u1429(.A(men_men_n255_), .B(u), .Y(men_men_n1458_));
  NO2        u1430(.A(m), .B(i), .Y(men_men_n1459_));
  BUFFER     u1431(.A(men_men_n1459_), .Y(men_men_n1460_));
  AOI220     u1432(.A0(men_men_n1460_), .A1(men_men_n1339_), .B0(men_men_n1043_), .B1(men_men_n1458_), .Y(men_men_n1461_));
  NA3        u1433(.A(men_men_n1461_), .B(men_men_n1457_), .C(men_men_n1454_), .Y(men_men_n1462_));
  NO4        u1434(.A(men_men_n1462_), .B(men_men_n1453_), .C(men_men_n1451_), .D(men_men_n1448_), .Y(men_men_n1463_));
  NA3        u1435(.A(men_men_n1463_), .B(men_men_n1445_), .C(men_men_n1440_), .Y(men_men_n1464_));
  NA3        u1436(.A(men_men_n940_), .B(men_men_n139_), .C(men_men_n46_), .Y(men_men_n1465_));
  NO2        u1437(.A(men_men_n149_), .B(men_men_n1465_), .Y(men_men_n1466_));
  AO210      u1438(.A0(men_men_n133_), .A1(l), .B0(men_men_n1363_), .Y(men_men_n1467_));
  NO2        u1439(.A(men_men_n72_), .B(c), .Y(men_men_n1468_));
  NO4        u1440(.A(men_men_n1326_), .B(men_men_n185_), .C(men_men_n450_), .D(men_men_n45_), .Y(men_men_n1469_));
  AOI210     u1441(.A0(men_men_n1416_), .A1(men_men_n1468_), .B0(men_men_n1469_), .Y(men_men_n1470_));
  NA2        u1442(.A(men_men_n1470_), .B(men_men_n1467_), .Y(men_men_n1471_));
  NO2        u1443(.A(men_men_n1471_), .B(men_men_n1466_), .Y(men_men_n1472_));
  NO4        u1444(.A(men_men_n226_), .B(men_men_n185_), .C(men_men_n260_), .D(k), .Y(men_men_n1473_));
  NO2        u1445(.A(men_men_n1465_), .B(men_men_n109_), .Y(men_men_n1474_));
  NOi21      u1446(.An(men_men_n1306_), .B(e), .Y(men_men_n1475_));
  NO3        u1447(.A(men_men_n1475_), .B(men_men_n1474_), .C(men_men_n1473_), .Y(men_men_n1476_));
  NA2        u1448(.A(men_men_n1027_), .B(men_men_n161_), .Y(men_men_n1477_));
  NOi31      u1449(.An(men_men_n30_), .B(men_men_n1477_), .C(n), .Y(men_men_n1478_));
  INV        u1450(.A(men_men_n1478_), .Y(men_men_n1479_));
  NA2        u1451(.A(men_men_n59_), .B(a), .Y(men_men_n1480_));
  NO2        u1452(.A(men_men_n1378_), .B(men_men_n1480_), .Y(men_men_n1481_));
  NA4        u1453(.A(men_men_n1495_), .B(men_men_n1479_), .C(men_men_n1476_), .D(men_men_n1472_), .Y(men_men_n1482_));
  OR4        u1454(.A(men_men_n1482_), .B(men_men_n1464_), .C(men_men_n1426_), .D(men_men_n1382_), .Y(men04));
  NOi31      u1455(.An(men_men_n1369_), .B(men_men_n1370_), .C(men_men_n1015_), .Y(men_men_n1484_));
  NA2        u1456(.A(men_men_n1420_), .B(men_men_n809_), .Y(men_men_n1485_));
  NO4        u1457(.A(men_men_n1485_), .B(men_men_n1006_), .C(men_men_n481_), .D(j), .Y(men_men_n1486_));
  OR3        u1458(.A(men_men_n1486_), .B(men_men_n1484_), .C(men_men_n1033_), .Y(men_men_n1487_));
  NO3        u1459(.A(men_men_n1315_), .B(men_men_n88_), .C(k), .Y(men_men_n1488_));
  AOI210     u1460(.A0(men_men_n1488_), .A1(men_men_n1026_), .B0(men_men_n1159_), .Y(men_men_n1489_));
  NA2        u1461(.A(men_men_n1489_), .B(men_men_n1184_), .Y(men_men_n1490_));
  NO4        u1462(.A(men_men_n1490_), .B(men_men_n1487_), .C(men_men_n1041_), .D(men_men_n1020_), .Y(men_men_n1491_));
  NA4        u1463(.A(men_men_n1491_), .B(men_men_n1096_), .C(men_men_n1081_), .D(men_men_n1069_), .Y(men05));
  INV        u1464(.A(men_men_n1481_), .Y(men_men_n1495_));
  INV        u1465(.A(men_men_n1386_), .Y(men_men_n1496_));
  INV        u1466(.A(a), .Y(men_men_n1497_));
  INV        u1467(.A(c), .Y(men_men_n1498_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule