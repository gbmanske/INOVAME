// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n117_, new_new_n118_, new_new_n120_,
    new_new_n121_, new_new_n122_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n314_, new_new_n315_, new_new_n316_, new_new_n317_,
    new_new_n318_, new_new_n319_, new_new_n320_, new_new_n321_,
    new_new_n322_, new_new_n323_, new_new_n324_, new_new_n325_,
    new_new_n326_, new_new_n327_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n336_, new_new_n337_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n350_, new_new_n351_, new_new_n352_, new_new_n353_,
    new_new_n354_, new_new_n355_, new_new_n356_, new_new_n357_,
    new_new_n358_, new_new_n359_, new_new_n360_, new_new_n361_,
    new_new_n362_, new_new_n363_, new_new_n364_, new_new_n365_,
    new_new_n366_, new_new_n367_, new_new_n368_, new_new_n369_,
    new_new_n370_, new_new_n371_, new_new_n372_, new_new_n373_,
    new_new_n374_, new_new_n375_, new_new_n376_, new_new_n377_,
    new_new_n378_, new_new_n379_, new_new_n380_, new_new_n381_,
    new_new_n382_, new_new_n383_, new_new_n384_, new_new_n385_,
    new_new_n386_, new_new_n387_, new_new_n388_, new_new_n389_,
    new_new_n390_, new_new_n391_, new_new_n392_, new_new_n393_,
    new_new_n394_, new_new_n395_, new_new_n396_, new_new_n397_,
    new_new_n398_, new_new_n399_, new_new_n400_, new_new_n401_,
    new_new_n402_, new_new_n403_, new_new_n404_, new_new_n405_,
    new_new_n407_, new_new_n408_, new_new_n409_, new_new_n410_,
    new_new_n411_, new_new_n412_, new_new_n413_, new_new_n414_,
    new_new_n415_, new_new_n416_, new_new_n417_, new_new_n418_,
    new_new_n419_, new_new_n420_, new_new_n421_, new_new_n422_,
    new_new_n423_, new_new_n424_, new_new_n425_, new_new_n426_,
    new_new_n427_, new_new_n428_, new_new_n429_, new_new_n430_,
    new_new_n431_, new_new_n432_, new_new_n433_, new_new_n434_,
    new_new_n435_, new_new_n436_, new_new_n437_, new_new_n438_,
    new_new_n439_, new_new_n440_, new_new_n441_, new_new_n442_,
    new_new_n443_, new_new_n444_, new_new_n445_, new_new_n446_,
    new_new_n448_, new_new_n449_, new_new_n450_, new_new_n451_,
    new_new_n452_, new_new_n453_, new_new_n454_, new_new_n455_,
    new_new_n456_, new_new_n457_, new_new_n458_, new_new_n459_,
    new_new_n460_, new_new_n461_, new_new_n462_, new_new_n463_,
    new_new_n464_, new_new_n465_, new_new_n466_, new_new_n467_,
    new_new_n468_, new_new_n469_, new_new_n470_, new_new_n471_,
    new_new_n472_, new_new_n473_, new_new_n474_, new_new_n475_,
    new_new_n476_, new_new_n477_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n576_, new_new_n577_, new_new_n578_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(ori1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_5_), .A1(new_new_n46_), .B0(new_new_n45_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n50_), .B(new_new_n44_), .Y(new_new_n54_));
  NA3        g032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  OAI210     g035(.A0(new_new_n57_), .A1(new_new_n56_), .B0(new_new_n55_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi31      g043(.An(new_new_n65_), .B(new_new_n63_), .C(new_new_n59_), .Y(new_new_n66_));
  NA2        g044(.A(new_new_n49_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  INV        g053(.A(new_new_n75_), .Y(new_new_n76_));
  OAI210     g054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  INV        g057(.A(i_6_), .Y(new_new_n80_));
  NO2        g058(.A(i_2_), .B(i_7_), .Y(new_new_n81_));
  INV        g059(.A(new_new_n81_), .Y(new_new_n82_));
  OAI210     g060(.A0(i_1_), .A1(i_6_), .B0(new_new_n82_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_10_), .Y(new_new_n84_));
  NA2        g062(.A(i_6_), .B(i_9_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n84_), .B0(new_new_n61_), .Y(new_new_n86_));
  NA2        g064(.A(i_2_), .B(i_6_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n86_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n88_), .A1(new_new_n83_), .B0(new_new_n78_), .Y(new_new_n89_));
  AN3        g067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  INV        g069(.A(i_7_), .Y(new_new_n92_));
  NO2        g070(.A(i_0_), .B(i_5_), .Y(new_new_n93_));
  NO2        g071(.A(new_new_n93_), .B(new_new_n80_), .Y(new_new_n94_));
  NA2        g072(.A(i_12_), .B(i_3_), .Y(new_new_n95_));
  NAi21      g073(.An(i_7_), .B(i_11_), .Y(new_new_n96_));
  NO3        g074(.A(new_new_n96_), .B(new_new_n84_), .C(new_new_n51_), .Y(new_new_n97_));
  AN2        g075(.A(i_2_), .B(i_10_), .Y(new_new_n98_));
  NA2        g076(.A(i_12_), .B(i_7_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n100_));
  NA2        g078(.A(i_11_), .B(i_12_), .Y(new_new_n101_));
  NAi21      g079(.An(new_new_n97_), .B(new_new_n101_), .Y(new_new_n102_));
  NOi21      g080(.An(i_1_), .B(i_5_), .Y(new_new_n103_));
  NA2        g081(.A(new_new_n103_), .B(i_11_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n92_), .B(new_new_n37_), .Y(new_new_n105_));
  NA2        g083(.A(i_7_), .B(new_new_n25_), .Y(new_new_n106_));
  NA2        g084(.A(new_new_n106_), .B(new_new_n105_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n107_), .B(new_new_n45_), .Y(new_new_n108_));
  NA2        g086(.A(new_new_n85_), .B(new_new_n84_), .Y(new_new_n109_));
  NO2        g087(.A(i_1_), .B(new_new_n80_), .Y(new_new_n110_));
  NO2        g088(.A(i_6_), .B(i_5_), .Y(new_new_n111_));
  NA2        g089(.A(new_new_n111_), .B(i_3_), .Y(new_new_n112_));
  AO210      g090(.A0(new_new_n112_), .A1(new_new_n46_), .B0(new_new_n110_), .Y(new_new_n113_));
  OAI210     g091(.A0(new_new_n113_), .A1(new_new_n96_), .B0(new_new_n104_), .Y(new_new_n114_));
  NO3        g092(.A(new_new_n114_), .B(new_new_n102_), .C(new_new_n89_), .Y(new_new_n115_));
  NA3        g093(.A(new_new_n115_), .B(new_new_n77_), .C(new_new_n54_), .Y(ori2));
  NO2        g094(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n576_), .B(new_new_n117_), .Y(new_new_n118_));
  NA4        g096(.A(new_new_n118_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(ori0));
  NAi21      g097(.An(i_5_), .B(i_11_), .Y(new_new_n120_));
  NO2        g098(.A(i_0_), .B(i_1_), .Y(new_new_n121_));
  NA2        g099(.A(i_1_), .B(i_5_), .Y(new_new_n122_));
  NOi21      g100(.An(i_4_), .B(i_10_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(new_new_n40_), .Y(new_new_n124_));
  NOi21      g102(.An(i_4_), .B(i_9_), .Y(new_new_n125_));
  NOi21      g103(.An(i_11_), .B(i_13_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n126_), .B(new_new_n125_), .Y(new_new_n127_));
  NAi21      g105(.An(i_12_), .B(i_11_), .Y(new_new_n128_));
  NO2        g106(.A(new_new_n71_), .B(i_5_), .Y(new_new_n129_));
  NO2        g107(.A(i_2_), .B(i_1_), .Y(new_new_n130_));
  NAi21      g108(.An(i_4_), .B(i_12_), .Y(new_new_n131_));
  INV        g109(.A(i_8_), .Y(new_new_n132_));
  NO3        g110(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n133_));
  NO2        g111(.A(i_3_), .B(i_8_), .Y(new_new_n134_));
  NO3        g112(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n135_));
  NO2        g113(.A(new_new_n93_), .B(new_new_n56_), .Y(new_new_n136_));
  NO2        g114(.A(i_13_), .B(i_9_), .Y(new_new_n137_));
  NAi21      g115(.An(i_12_), .B(i_3_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n43_), .B(i_5_), .Y(new_new_n139_));
  NA3        g117(.A(i_13_), .B(new_new_n132_), .C(i_10_), .Y(new_new_n140_));
  NA2        g118(.A(i_0_), .B(i_5_), .Y(new_new_n141_));
  NAi31      g119(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n143_));
  NO2        g121(.A(new_new_n45_), .B(new_new_n61_), .Y(new_new_n144_));
  INV        g122(.A(i_13_), .Y(new_new_n145_));
  NO2        g123(.A(i_12_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g124(.A(i_12_), .B(new_new_n37_), .Y(new_new_n147_));
  INV        g125(.A(i_12_), .Y(new_new_n148_));
  NO3        g126(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n149_));
  NA2        g127(.A(i_2_), .B(i_1_), .Y(new_new_n150_));
  NO3        g128(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n151_));
  NAi21      g129(.An(i_4_), .B(i_3_), .Y(new_new_n152_));
  NO2        g130(.A(i_0_), .B(i_6_), .Y(new_new_n153_));
  NOi41      g131(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n154_));
  NO2        g132(.A(i_11_), .B(new_new_n145_), .Y(new_new_n155_));
  NOi21      g133(.An(i_1_), .B(i_6_), .Y(new_new_n156_));
  NAi21      g134(.An(i_3_), .B(i_7_), .Y(new_new_n157_));
  NA2        g135(.A(new_new_n148_), .B(i_9_), .Y(new_new_n158_));
  OR4        g136(.A(new_new_n158_), .B(new_new_n157_), .C(new_new_n156_), .D(new_new_n129_), .Y(new_new_n159_));
  NA2        g137(.A(new_new_n71_), .B(i_5_), .Y(new_new_n160_));
  NA2        g138(.A(i_3_), .B(i_9_), .Y(new_new_n161_));
  NAi21      g139(.An(i_7_), .B(i_10_), .Y(new_new_n162_));
  NO2        g140(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  NA3        g141(.A(new_new_n163_), .B(new_new_n160_), .C(new_new_n62_), .Y(new_new_n164_));
  NA2        g142(.A(new_new_n164_), .B(new_new_n159_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n155_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n152_), .B(i_2_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n155_), .B(i_9_), .Y(new_new_n168_));
  NO3        g146(.A(i_11_), .B(new_new_n145_), .C(new_new_n25_), .Y(new_new_n169_));
  NO3        g147(.A(i_12_), .B(new_new_n145_), .C(new_new_n37_), .Y(new_new_n170_));
  AN2        g148(.A(i_3_), .B(i_10_), .Y(new_new_n171_));
  NO2        g149(.A(i_5_), .B(new_new_n37_), .Y(new_new_n172_));
  NO3        g150(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n173_));
  NO2        g151(.A(i_2_), .B(i_3_), .Y(new_new_n174_));
  OR2        g152(.A(i_0_), .B(i_5_), .Y(new_new_n175_));
  NO2        g153(.A(i_12_), .B(i_10_), .Y(new_new_n176_));
  NOi21      g154(.An(i_5_), .B(i_0_), .Y(new_new_n177_));
  NO2        g155(.A(i_1_), .B(i_7_), .Y(new_new_n178_));
  NOi21      g156(.An(new_new_n122_), .B(new_new_n94_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n179_), .B(new_new_n106_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(i_3_), .Y(new_new_n181_));
  NO2        g159(.A(new_new_n132_), .B(i_9_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(new_new_n136_), .Y(new_new_n183_));
  NO2        g161(.A(new_new_n183_), .B(new_new_n45_), .Y(new_new_n184_));
  INV        g162(.A(new_new_n184_), .Y(new_new_n185_));
  AOI210     g163(.A0(new_new_n185_), .A1(new_new_n181_), .B0(new_new_n124_), .Y(new_new_n186_));
  INV        g164(.A(new_new_n186_), .Y(new_new_n187_));
  NOi32      g165(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n188_));
  INV        g166(.A(new_new_n188_), .Y(new_new_n189_));
  NOi32      g167(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n190_));
  NAi21      g168(.An(i_6_), .B(i_1_), .Y(new_new_n191_));
  NA3        g169(.A(new_new_n191_), .B(new_new_n190_), .C(new_new_n45_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n192_), .B(i_0_), .Y(new_new_n193_));
  NO2        g171(.A(i_1_), .B(new_new_n92_), .Y(new_new_n194_));
  NAi21      g172(.An(i_3_), .B(i_4_), .Y(new_new_n195_));
  NO2        g173(.A(new_new_n195_), .B(i_9_), .Y(new_new_n196_));
  AN2        g174(.A(i_6_), .B(i_7_), .Y(new_new_n197_));
  OAI210     g175(.A0(new_new_n197_), .A1(new_new_n194_), .B0(new_new_n196_), .Y(new_new_n198_));
  NA2        g176(.A(i_2_), .B(i_7_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n195_), .B(i_10_), .Y(new_new_n200_));
  NA3        g178(.A(new_new_n200_), .B(new_new_n199_), .C(new_new_n153_), .Y(new_new_n201_));
  AOI210     g179(.A0(new_new_n201_), .A1(new_new_n198_), .B0(new_new_n129_), .Y(new_new_n202_));
  AOI210     g180(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n203_));
  OAI210     g181(.A0(new_new_n203_), .A1(new_new_n130_), .B0(new_new_n200_), .Y(new_new_n204_));
  AOI220     g182(.A0(new_new_n200_), .A1(new_new_n178_), .B0(new_new_n149_), .B1(new_new_n130_), .Y(new_new_n205_));
  AOI210     g183(.A0(new_new_n205_), .A1(new_new_n204_), .B0(i_5_), .Y(new_new_n206_));
  NO3        g184(.A(new_new_n206_), .B(new_new_n202_), .C(new_new_n193_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n207_), .B(new_new_n189_), .Y(new_new_n208_));
  AN2        g186(.A(i_12_), .B(i_5_), .Y(new_new_n209_));
  INV        g187(.A(new_new_n209_), .Y(new_new_n210_));
  NO2        g188(.A(i_11_), .B(i_6_), .Y(new_new_n211_));
  NO2        g189(.A(i_5_), .B(i_10_), .Y(new_new_n212_));
  NO2        g190(.A(i_11_), .B(i_12_), .Y(new_new_n213_));
  NAi21      g191(.An(i_13_), .B(i_0_), .Y(new_new_n214_));
  NO3        g192(.A(i_1_), .B(i_12_), .C(new_new_n80_), .Y(new_new_n215_));
  NO2        g193(.A(i_0_), .B(i_11_), .Y(new_new_n216_));
  AN2        g194(.A(i_1_), .B(i_6_), .Y(new_new_n217_));
  NOi21      g195(.An(i_2_), .B(i_12_), .Y(new_new_n218_));
  NAi21      g196(.An(i_9_), .B(i_4_), .Y(new_new_n219_));
  OR2        g197(.A(i_13_), .B(i_10_), .Y(new_new_n220_));
  NO3        g198(.A(new_new_n220_), .B(new_new_n101_), .C(new_new_n219_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n127_), .B(new_new_n105_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n92_), .B(new_new_n25_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n170_), .B(new_new_n223_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n224_), .B(new_new_n179_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n132_), .B(i_10_), .Y(new_new_n226_));
  NA3        g204(.A(new_new_n160_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n226_), .Y(new_new_n228_));
  INV        g206(.A(new_new_n228_), .Y(new_new_n229_));
  NO2        g207(.A(new_new_n229_), .B(new_new_n168_), .Y(new_new_n230_));
  NO3        g208(.A(new_new_n230_), .B(new_new_n225_), .C(new_new_n208_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n71_), .B(i_13_), .Y(new_new_n232_));
  NO2        g210(.A(i_10_), .B(i_9_), .Y(new_new_n233_));
  INV        g211(.A(new_new_n91_), .Y(new_new_n234_));
  NA2        g212(.A(i_8_), .B(i_9_), .Y(new_new_n235_));
  NA2        g213(.A(new_new_n170_), .B(new_new_n136_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n155_), .B(new_new_n172_), .Y(new_new_n238_));
  NO3        g216(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n239_), .Y(new_new_n240_));
  NA3        g218(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n241_));
  NA4        g219(.A(new_new_n120_), .B(new_new_n100_), .C(new_new_n78_), .D(new_new_n23_), .Y(new_new_n242_));
  OAI220     g220(.A0(new_new_n242_), .A1(new_new_n241_), .B0(new_new_n240_), .B1(new_new_n238_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n243_), .B(new_new_n237_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n90_), .B(i_13_), .Y(new_new_n245_));
  NO3        g223(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n246_));
  NO2        g224(.A(i_6_), .B(i_7_), .Y(new_new_n247_));
  NO2        g225(.A(i_11_), .B(i_1_), .Y(new_new_n248_));
  NOi21      g226(.An(i_2_), .B(i_7_), .Y(new_new_n249_));
  NO2        g227(.A(i_6_), .B(i_10_), .Y(new_new_n250_));
  NA3        g228(.A(new_new_n154_), .B(new_new_n126_), .C(new_new_n111_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n45_), .B(new_new_n43_), .Y(new_new_n252_));
  NA2        g230(.A(new_new_n239_), .B(new_new_n212_), .Y(new_new_n253_));
  NAi21      g231(.An(new_new_n140_), .B(new_new_n213_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n178_), .B(new_new_n141_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n255_), .B(new_new_n254_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n27_), .B(i_10_), .Y(new_new_n257_));
  NA2        g235(.A(new_new_n173_), .B(new_new_n149_), .Y(new_new_n258_));
  OAI220     g236(.A0(new_new_n258_), .A1(new_new_n227_), .B0(new_new_n257_), .B1(new_new_n245_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n259_), .B(new_new_n256_), .Y(new_new_n260_));
  NA3        g238(.A(new_new_n260_), .B(new_new_n251_), .C(new_new_n244_), .Y(new_new_n261_));
  NA2        g239(.A(new_new_n209_), .B(new_new_n145_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n197_), .B(new_new_n190_), .Y(new_new_n263_));
  OR2        g241(.A(new_new_n262_), .B(new_new_n263_), .Y(new_new_n264_));
  AOI210     g242(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n221_), .Y(new_new_n265_));
  NA2        g243(.A(new_new_n265_), .B(new_new_n264_), .Y(new_new_n266_));
  INV        g244(.A(new_new_n266_), .Y(new_new_n267_));
  NA2        g245(.A(new_new_n160_), .B(new_new_n62_), .Y(new_new_n268_));
  OAI210     g246(.A0(i_8_), .A1(new_new_n268_), .B0(new_new_n113_), .Y(new_new_n269_));
  NA2        g247(.A(new_new_n269_), .B(new_new_n222_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n270_), .B(new_new_n267_), .Y(new_new_n271_));
  NO2        g249(.A(i_12_), .B(new_new_n132_), .Y(new_new_n272_));
  NA2        g250(.A(new_new_n43_), .B(i_10_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(i_6_), .Y(new_new_n274_));
  NO2        g252(.A(i_0_), .B(i_5_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n170_), .B(new_new_n79_), .Y(new_new_n276_));
  NO2        g254(.A(i_11_), .B(new_new_n276_), .Y(new_new_n277_));
  NA2        g255(.A(new_new_n144_), .B(new_new_n143_), .Y(new_new_n278_));
  NA2        g256(.A(new_new_n233_), .B(i_4_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n278_), .B(new_new_n279_), .Y(new_new_n280_));
  AOI210     g258(.A0(new_new_n191_), .A1(new_new_n45_), .B0(new_new_n194_), .Y(new_new_n281_));
  NA2        g259(.A(i_0_), .B(new_new_n47_), .Y(new_new_n282_));
  NA3        g260(.A(new_new_n272_), .B(new_new_n169_), .C(new_new_n282_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n281_), .B(new_new_n283_), .Y(new_new_n284_));
  NO3        g262(.A(new_new_n284_), .B(new_new_n280_), .C(new_new_n277_), .Y(new_new_n285_));
  NOi21      g263(.An(i_10_), .B(i_6_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n80_), .B(new_new_n25_), .Y(new_new_n287_));
  INV        g265(.A(new_new_n174_), .Y(new_new_n288_));
  NO2        g266(.A(i_12_), .B(new_new_n80_), .Y(new_new_n289_));
  NA3        g267(.A(new_new_n289_), .B(new_new_n169_), .C(new_new_n282_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n211_), .B(new_new_n170_), .C(new_new_n141_), .Y(new_new_n291_));
  AOI210     g269(.A0(new_new_n291_), .A1(new_new_n290_), .B0(new_new_n288_), .Y(new_new_n292_));
  OR2        g270(.A(i_2_), .B(i_5_), .Y(new_new_n293_));
  OR2        g271(.A(new_new_n293_), .B(new_new_n217_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n199_), .B(new_new_n153_), .Y(new_new_n295_));
  AOI210     g273(.A0(new_new_n295_), .A1(new_new_n294_), .B0(new_new_n254_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n296_), .B(new_new_n292_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n297_), .B(new_new_n285_), .Y(new_new_n298_));
  NO3        g276(.A(new_new_n298_), .B(new_new_n271_), .C(new_new_n261_), .Y(new_new_n299_));
  NA4        g277(.A(new_new_n299_), .B(new_new_n231_), .C(new_new_n187_), .D(new_new_n166_), .Y(ori7));
  NO2        g278(.A(new_new_n87_), .B(new_new_n52_), .Y(new_new_n301_));
  NA2        g279(.A(new_new_n250_), .B(new_new_n79_), .Y(new_new_n302_));
  NA2        g280(.A(i_11_), .B(new_new_n132_), .Y(new_new_n303_));
  NO2        g281(.A(i_13_), .B(new_new_n302_), .Y(new_new_n304_));
  NA3        g282(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n148_), .B(i_4_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n306_), .B(i_8_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n95_), .B(new_new_n305_), .Y(new_new_n308_));
  NA2        g286(.A(i_2_), .B(new_new_n80_), .Y(new_new_n309_));
  OAI210     g287(.A0(new_new_n81_), .A1(new_new_n134_), .B0(new_new_n135_), .Y(new_new_n310_));
  NO2        g288(.A(i_7_), .B(new_new_n37_), .Y(new_new_n311_));
  NA2        g289(.A(i_4_), .B(i_8_), .Y(new_new_n312_));
  AOI210     g290(.A0(new_new_n312_), .A1(new_new_n171_), .B0(new_new_n311_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n313_), .B(new_new_n309_), .Y(new_new_n314_));
  NO4        g292(.A(new_new_n314_), .B(new_new_n308_), .C(new_new_n304_), .D(new_new_n301_), .Y(new_new_n315_));
  OR2        g293(.A(i_6_), .B(i_10_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n316_), .B(new_new_n23_), .Y(new_new_n317_));
  OR3        g295(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n318_));
  INV        g296(.A(new_new_n133_), .Y(new_new_n319_));
  INV        g297(.A(new_new_n317_), .Y(new_new_n320_));
  OR2        g298(.A(new_new_n320_), .B(new_new_n288_), .Y(new_new_n321_));
  AOI210     g299(.A0(new_new_n321_), .A1(new_new_n315_), .B0(new_new_n61_), .Y(new_new_n322_));
  NOi21      g300(.An(i_11_), .B(i_7_), .Y(new_new_n323_));
  AO210      g301(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n324_), .B(new_new_n323_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n325_), .B(new_new_n137_), .Y(new_new_n326_));
  NA3        g304(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n326_), .B(new_new_n61_), .Y(new_new_n328_));
  NO3        g306(.A(new_new_n162_), .B(new_new_n138_), .C(new_new_n303_), .Y(new_new_n329_));
  OAI210     g307(.A0(new_new_n329_), .A1(new_new_n146_), .B0(new_new_n61_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n218_), .B(new_new_n31_), .Y(new_new_n331_));
  OR2        g309(.A(new_new_n138_), .B(new_new_n96_), .Y(new_new_n332_));
  NA2        g310(.A(new_new_n332_), .B(new_new_n331_), .Y(new_new_n333_));
  NO2        g311(.A(i_1_), .B(i_4_), .Y(new_new_n334_));
  NA2        g312(.A(new_new_n334_), .B(new_new_n333_), .Y(new_new_n335_));
  NO2        g313(.A(i_1_), .B(i_12_), .Y(new_new_n336_));
  NA3        g314(.A(new_new_n336_), .B(new_new_n98_), .C(new_new_n24_), .Y(new_new_n337_));
  BUFFER     g315(.A(new_new_n337_), .Y(new_new_n338_));
  NA3        g316(.A(new_new_n338_), .B(new_new_n335_), .C(new_new_n330_), .Y(new_new_n339_));
  OAI210     g317(.A0(new_new_n339_), .A1(new_new_n328_), .B0(i_6_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n327_), .B(new_new_n96_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n289_), .Y(new_new_n342_));
  NO2        g320(.A(i_6_), .B(i_11_), .Y(new_new_n343_));
  INV        g321(.A(new_new_n342_), .Y(new_new_n344_));
  NO3        g322(.A(new_new_n316_), .B(i_8_), .C(new_new_n23_), .Y(new_new_n345_));
  AOI210     g323(.A0(i_1_), .A1(new_new_n163_), .B0(new_new_n345_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n346_), .B(new_new_n43_), .Y(new_new_n347_));
  NA3        g325(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n348_));
  NA2        g326(.A(i_2_), .B(new_new_n43_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(new_new_n348_), .Y(new_new_n350_));
  AOI210     g328(.A0(new_new_n248_), .A1(new_new_n223_), .B0(new_new_n151_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n351_), .B(new_new_n309_), .Y(new_new_n352_));
  OR2        g330(.A(new_new_n352_), .B(new_new_n350_), .Y(new_new_n353_));
  NO3        g331(.A(new_new_n353_), .B(new_new_n347_), .C(new_new_n344_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n148_), .B(new_new_n92_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(new_new_n323_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n356_), .B(i_1_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(new_new_n318_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n219_), .B(new_new_n80_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n358_), .B(new_new_n45_), .Y(new_new_n360_));
  NA2        g338(.A(i_3_), .B(new_new_n132_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(new_new_n99_), .Y(new_new_n362_));
  AN2        g340(.A(new_new_n362_), .B(new_new_n274_), .Y(new_new_n363_));
  NO2        g341(.A(i_8_), .B(new_new_n43_), .Y(new_new_n364_));
  NA2        g342(.A(i_1_), .B(i_3_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n235_), .B(new_new_n87_), .Y(new_new_n366_));
  AOI210     g344(.A0(new_new_n364_), .A1(new_new_n286_), .B0(new_new_n366_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n365_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n368_), .B(new_new_n363_), .Y(new_new_n369_));
  NA4        g347(.A(new_new_n369_), .B(new_new_n360_), .C(new_new_n354_), .D(new_new_n340_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n197_), .B(new_new_n196_), .Y(new_new_n371_));
  NO3        g349(.A(new_new_n249_), .B(new_new_n312_), .C(new_new_n80_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n372_), .B(new_new_n25_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n373_), .B(new_new_n371_), .Y(new_new_n374_));
  NA2        g352(.A(new_new_n374_), .B(i_1_), .Y(new_new_n375_));
  INV        g353(.A(i_1_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n375_), .B(i_13_), .Y(new_new_n377_));
  OR2        g355(.A(i_11_), .B(i_7_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n52_), .B(i_12_), .Y(new_new_n379_));
  INV        g357(.A(new_new_n379_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n249_), .B(new_new_n24_), .Y(new_new_n381_));
  AOI220     g359(.A0(new_new_n381_), .A1(new_new_n359_), .B0(new_new_n154_), .B1(new_new_n110_), .Y(new_new_n382_));
  OAI220     g360(.A0(new_new_n382_), .A1(new_new_n41_), .B0(new_new_n380_), .B1(new_new_n87_), .Y(new_new_n383_));
  INV        g361(.A(new_new_n383_), .Y(new_new_n384_));
  NOi31      g362(.An(new_new_n577_), .B(new_new_n302_), .C(new_new_n43_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n109_), .B(i_13_), .Y(new_new_n386_));
  NO2        g364(.A(new_new_n348_), .B(new_new_n99_), .Y(new_new_n387_));
  INV        g365(.A(new_new_n387_), .Y(new_new_n388_));
  OAI220     g366(.A0(new_new_n388_), .A1(new_new_n69_), .B0(new_new_n386_), .B1(new_new_n376_), .Y(new_new_n389_));
  NO3        g367(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n92_), .Y(new_new_n390_));
  INV        g368(.A(new_new_n390_), .Y(new_new_n391_));
  AOI210     g369(.A0(new_new_n211_), .A1(i_2_), .B0(new_new_n86_), .Y(new_new_n392_));
  OAI220     g370(.A0(new_new_n392_), .A1(new_new_n307_), .B0(new_new_n391_), .B1(new_new_n319_), .Y(new_new_n393_));
  NO3        g371(.A(new_new_n393_), .B(new_new_n389_), .C(new_new_n385_), .Y(new_new_n394_));
  OR2        g372(.A(i_11_), .B(i_6_), .Y(new_new_n395_));
  NA3        g373(.A(new_new_n218_), .B(new_new_n311_), .C(new_new_n91_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n343_), .B(i_13_), .Y(new_new_n397_));
  NAi21      g375(.An(i_11_), .B(i_12_), .Y(new_new_n398_));
  NO3        g376(.A(new_new_n398_), .B(i_13_), .C(new_new_n80_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n289_), .B(new_new_n312_), .Y(new_new_n400_));
  AOI210     g378(.A0(new_new_n400_), .A1(new_new_n173_), .B0(new_new_n399_), .Y(new_new_n401_));
  NA3        g379(.A(new_new_n401_), .B(new_new_n397_), .C(new_new_n396_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n402_), .B(new_new_n61_), .Y(new_new_n403_));
  NO2        g381(.A(i_2_), .B(i_12_), .Y(new_new_n404_));
  NA3        g382(.A(new_new_n403_), .B(new_new_n394_), .C(new_new_n384_), .Y(new_new_n405_));
  OR4        g383(.A(new_new_n405_), .B(new_new_n377_), .C(new_new_n370_), .D(new_new_n322_), .Y(ori5));
  NA2        g384(.A(new_new_n356_), .B(new_new_n167_), .Y(new_new_n407_));
  NA3        g385(.A(new_new_n24_), .B(new_new_n404_), .C(new_new_n96_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n307_), .B(i_11_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n81_), .B(new_new_n409_), .Y(new_new_n410_));
  NA3        g388(.A(new_new_n410_), .B(new_new_n408_), .C(new_new_n407_), .Y(new_new_n411_));
  NO3        g389(.A(i_11_), .B(new_new_n148_), .C(i_13_), .Y(new_new_n412_));
  NO2        g390(.A(new_new_n106_), .B(new_new_n23_), .Y(new_new_n413_));
  NA2        g391(.A(i_12_), .B(i_8_), .Y(new_new_n414_));
  OAI210     g392(.A0(new_new_n45_), .A1(i_3_), .B0(new_new_n414_), .Y(new_new_n415_));
  INV        g393(.A(new_new_n233_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n415_), .B(new_new_n413_), .Y(new_new_n417_));
  INV        g395(.A(new_new_n417_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n418_), .B(new_new_n411_), .Y(new_new_n419_));
  INV        g397(.A(new_new_n126_), .Y(new_new_n420_));
  INV        g398(.A(new_new_n154_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n421_), .B(new_new_n420_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n235_), .B(new_new_n26_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n423_), .B(new_new_n223_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n424_), .B(i_2_), .Y(new_new_n425_));
  INV        g403(.A(new_new_n425_), .Y(new_new_n426_));
  AOI210     g404(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n220_), .Y(new_new_n427_));
  AOI210     g405(.A0(new_new_n427_), .A1(new_new_n426_), .B0(new_new_n422_), .Y(new_new_n428_));
  NO2        g406(.A(new_new_n131_), .B(new_new_n107_), .Y(new_new_n429_));
  OAI210     g407(.A0(new_new_n429_), .A1(new_new_n413_), .B0(i_2_), .Y(new_new_n430_));
  INV        g408(.A(new_new_n127_), .Y(new_new_n431_));
  NO3        g409(.A(new_new_n324_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n432_));
  AOI210     g410(.A0(new_new_n431_), .A1(new_new_n81_), .B0(new_new_n432_), .Y(new_new_n433_));
  AOI210     g411(.A0(new_new_n433_), .A1(new_new_n430_), .B0(new_new_n132_), .Y(new_new_n434_));
  OA210      g412(.A0(new_new_n325_), .A1(new_new_n108_), .B0(i_13_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n133_), .B(new_new_n134_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n199_), .Y(new_new_n437_));
  INV        g415(.A(new_new_n138_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n438_), .B(new_new_n223_), .Y(new_new_n439_));
  NA3        g417(.A(i_2_), .B(new_new_n171_), .C(new_new_n106_), .Y(new_new_n440_));
  NA2        g418(.A(new_new_n440_), .B(new_new_n439_), .Y(new_new_n441_));
  NO4        g419(.A(new_new_n441_), .B(new_new_n437_), .C(new_new_n435_), .D(new_new_n434_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n60_), .B(i_12_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n443_), .B(new_new_n108_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n444_), .B(new_new_n303_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n445_), .B(new_new_n36_), .Y(new_new_n446_));
  NA4        g424(.A(new_new_n446_), .B(new_new_n442_), .C(new_new_n428_), .D(new_new_n419_), .Y(ori6));
  NO2        g425(.A(new_new_n142_), .B(new_new_n252_), .Y(new_new_n448_));
  INV        g426(.A(new_new_n177_), .Y(new_new_n449_));
  OR2        g427(.A(new_new_n449_), .B(i_12_), .Y(new_new_n450_));
  INV        g428(.A(new_new_n176_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n73_), .B(new_new_n110_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n452_), .B(new_new_n451_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n156_), .B(i_9_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n454_), .B(new_new_n443_), .Y(new_new_n455_));
  AOI210     g433(.A0(new_new_n455_), .A1(new_new_n263_), .B0(new_new_n129_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n32_), .B(i_11_), .Y(new_new_n457_));
  NAi32      g435(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n458_));
  NO2        g436(.A(new_new_n395_), .B(new_new_n458_), .Y(new_new_n459_));
  OR3        g437(.A(new_new_n459_), .B(new_new_n456_), .C(new_new_n453_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n378_), .B(i_2_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n47_), .B(new_new_n37_), .Y(new_new_n462_));
  INV        g440(.A(new_new_n462_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n463_), .B(new_new_n461_), .Y(new_new_n464_));
  BUFFER     g442(.A(new_new_n325_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n465_), .B(new_new_n121_), .Y(new_new_n466_));
  AO210      g444(.A0(new_new_n253_), .A1(new_new_n416_), .B0(new_new_n36_), .Y(new_new_n467_));
  NA3        g445(.A(new_new_n467_), .B(new_new_n466_), .C(new_new_n464_), .Y(new_new_n468_));
  INV        g446(.A(new_new_n448_), .Y(new_new_n469_));
  NA3        g447(.A(new_new_n199_), .B(new_new_n149_), .C(new_new_n121_), .Y(new_new_n470_));
  NA3        g448(.A(new_new_n470_), .B(new_new_n469_), .C(new_new_n310_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n316_), .B(i_2_), .Y(new_new_n472_));
  OAI210     g450(.A0(new_new_n472_), .A1(new_new_n78_), .B0(new_new_n216_), .Y(new_new_n473_));
  INV        g451(.A(new_new_n294_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n474_), .B(new_new_n176_), .Y(new_new_n475_));
  NA2        g453(.A(new_new_n475_), .B(new_new_n473_), .Y(new_new_n476_));
  NO4        g454(.A(new_new_n476_), .B(new_new_n471_), .C(new_new_n468_), .D(new_new_n460_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n477_), .B(new_new_n450_), .C(new_new_n207_), .Y(ori3));
  NA2        g456(.A(i_12_), .B(i_10_), .Y(new_new_n479_));
  NO2        g457(.A(i_11_), .B(new_new_n148_), .Y(new_new_n480_));
  NA3        g458(.A(new_new_n470_), .B(new_new_n310_), .C(new_new_n198_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n481_), .B(new_new_n40_), .Y(new_new_n482_));
  NOi21      g460(.An(new_new_n90_), .B(new_new_n424_), .Y(new_new_n483_));
  NO3        g461(.A(new_new_n332_), .B(new_new_n235_), .C(new_new_n110_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n218_), .B(new_new_n44_), .Y(new_new_n485_));
  AN2        g463(.A(new_new_n234_), .B(new_new_n53_), .Y(new_new_n486_));
  NO3        g464(.A(new_new_n486_), .B(new_new_n484_), .C(new_new_n483_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n487_), .A1(new_new_n482_), .B0(new_new_n47_), .Y(new_new_n488_));
  NO4        g466(.A(new_new_n203_), .B(new_new_n209_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n129_), .B(new_new_n286_), .Y(new_new_n490_));
  NOi21      g468(.An(new_new_n490_), .B(new_new_n489_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n491_), .B(new_new_n61_), .Y(new_new_n492_));
  NOi21      g470(.An(i_5_), .B(i_9_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n232_), .Y(new_new_n494_));
  AOI210     g472(.A0(new_new_n578_), .A1(new_new_n248_), .B0(new_new_n372_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n495_), .B(new_new_n494_), .Y(new_new_n496_));
  NO3        g474(.A(new_new_n496_), .B(new_new_n492_), .C(new_new_n488_), .Y(new_new_n497_));
  BUFFER     g475(.A(i_0_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n287_), .B(i_0_), .Y(new_new_n499_));
  NO3        g477(.A(new_new_n499_), .B(new_new_n210_), .C(new_new_n81_), .Y(new_new_n500_));
  NO4        g478(.A(new_new_n293_), .B(i_12_), .C(new_new_n220_), .D(new_new_n217_), .Y(new_new_n501_));
  AOI210     g479(.A0(new_new_n501_), .A1(i_11_), .B0(new_new_n500_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n412_), .B(new_new_n177_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n81_), .B(new_new_n56_), .Y(new_new_n504_));
  NO2        g482(.A(new_new_n504_), .B(new_new_n503_), .Y(new_new_n505_));
  NO2        g483(.A(new_new_n158_), .B(new_new_n122_), .Y(new_new_n506_));
  NO4        g484(.A(new_new_n99_), .B(new_new_n56_), .C(new_new_n361_), .D(i_5_), .Y(new_new_n507_));
  AO220      g485(.A0(new_new_n507_), .A1(i_10_), .B0(new_new_n506_), .B1(i_6_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n508_), .B(new_new_n505_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n509_), .B(new_new_n502_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n511_));
  NA2        g489(.A(i_11_), .B(i_9_), .Y(new_new_n512_));
  NO3        g490(.A(i_12_), .B(new_new_n512_), .C(new_new_n309_), .Y(new_new_n513_));
  AN2        g491(.A(new_new_n513_), .B(new_new_n511_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n512_), .B(new_new_n71_), .Y(new_new_n515_));
  INV        g493(.A(new_new_n215_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n516_), .B(new_new_n494_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n517_), .B(new_new_n514_), .Y(new_new_n518_));
  INV        g496(.A(new_new_n175_), .Y(new_new_n519_));
  INV        g497(.A(new_new_n518_), .Y(new_new_n520_));
  INV        g498(.A(new_new_n479_), .Y(new_new_n521_));
  OA210      g499(.A0(new_new_n247_), .A1(new_new_n144_), .B0(new_new_n246_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n521_), .B(new_new_n515_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n381_), .B(new_new_n275_), .Y(new_new_n524_));
  NAi21      g502(.An(i_9_), .B(i_5_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n525_), .B(new_new_n214_), .Y(new_new_n526_));
  NA2        g504(.A(new_new_n526_), .B(new_new_n325_), .Y(new_new_n527_));
  OAI220     g505(.A0(new_new_n527_), .A1(new_new_n80_), .B0(new_new_n524_), .B1(new_new_n127_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n528_), .B(new_new_n266_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n529_), .B(new_new_n523_), .Y(new_new_n530_));
  NO3        g508(.A(new_new_n530_), .B(new_new_n520_), .C(new_new_n510_), .Y(new_new_n531_));
  NO2        g509(.A(new_new_n498_), .B(new_new_n398_), .Y(new_new_n532_));
  NA2        g510(.A(new_new_n153_), .B(new_new_n147_), .Y(new_new_n533_));
  AOI210     g511(.A0(new_new_n533_), .A1(new_new_n499_), .B0(new_new_n122_), .Y(new_new_n534_));
  NO3        g512(.A(new_new_n139_), .B(new_new_n209_), .C(i_0_), .Y(new_new_n535_));
  OAI210     g513(.A0(new_new_n535_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n536_));
  INV        g514(.A(new_new_n536_), .Y(new_new_n537_));
  NO2        g515(.A(new_new_n152_), .B(new_new_n87_), .Y(new_new_n538_));
  AOI210     g516(.A0(new_new_n538_), .A1(new_new_n532_), .B0(new_new_n97_), .Y(new_new_n539_));
  OR2        g517(.A(new_new_n539_), .B(i_5_), .Y(new_new_n540_));
  AOI210     g518(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n128_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n541_), .B(new_new_n522_), .Y(new_new_n542_));
  NO3        g520(.A(new_new_n485_), .B(new_new_n52_), .C(new_new_n47_), .Y(new_new_n543_));
  INV        g521(.A(new_new_n251_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n544_), .B(new_new_n543_), .Y(new_new_n545_));
  NA3        g523(.A(new_new_n212_), .B(new_new_n126_), .C(new_new_n125_), .Y(new_new_n546_));
  INV        g524(.A(new_new_n546_), .Y(new_new_n547_));
  NO3        g525(.A(new_new_n512_), .B(new_new_n141_), .C(new_new_n131_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n548_), .B(new_new_n547_), .Y(new_new_n549_));
  NA4        g527(.A(new_new_n549_), .B(new_new_n545_), .C(new_new_n542_), .D(new_new_n540_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n80_), .B(i_5_), .Y(new_new_n551_));
  NA3        g529(.A(new_new_n480_), .B(new_new_n98_), .C(new_new_n106_), .Y(new_new_n552_));
  INV        g530(.A(new_new_n552_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n553_), .B(new_new_n551_), .Y(new_new_n554_));
  NAi21      g532(.An(new_new_n151_), .B(new_new_n152_), .Y(new_new_n555_));
  NO4        g533(.A(new_new_n150_), .B(new_new_n139_), .C(i_0_), .D(i_12_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n556_), .B(new_new_n555_), .Y(new_new_n557_));
  NA2        g535(.A(new_new_n557_), .B(new_new_n554_), .Y(new_new_n558_));
  NO4        g536(.A(new_new_n558_), .B(new_new_n550_), .C(new_new_n537_), .D(new_new_n534_), .Y(new_new_n559_));
  OAI210     g537(.A0(new_new_n461_), .A1(new_new_n457_), .B0(new_new_n37_), .Y(new_new_n560_));
  INV        g538(.A(new_new_n560_), .Y(new_new_n561_));
  NA2        g539(.A(new_new_n561_), .B(new_new_n137_), .Y(new_new_n562_));
  NAi31      g540(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n68_), .B(new_new_n563_), .Y(new_new_n564_));
  AOI210     g542(.A0(new_new_n564_), .A1(new_new_n47_), .B0(new_new_n501_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n565_), .A1(new_new_n562_), .B0(new_new_n71_), .Y(new_new_n566_));
  INV        g544(.A(new_new_n206_), .Y(new_new_n567_));
  NO2        g545(.A(new_new_n567_), .B(new_new_n420_), .Y(new_new_n568_));
  NO3        g546(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n569_));
  OAI210     g547(.A0(new_new_n519_), .A1(new_new_n172_), .B0(new_new_n569_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n570_), .B(new_new_n398_), .Y(new_new_n571_));
  NO3        g549(.A(new_new_n571_), .B(new_new_n568_), .C(new_new_n566_), .Y(new_new_n572_));
  NA4        g550(.A(new_new_n572_), .B(new_new_n559_), .C(new_new_n531_), .D(new_new_n497_), .Y(ori4));
  INV        g551(.A(i_6_), .Y(new_new_n576_));
  INV        g552(.A(i_13_), .Y(new_new_n577_));
  INV        g553(.A(i_6_), .Y(new_new_n578_));
endmodule


