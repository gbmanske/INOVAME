library verilog;
use verilog.vl_types.all;
entity shiftreg4bits_vlg_vec_tst is
end shiftreg4bits_vlg_vec_tst;
