library verilog;
use verilog.vl_types.all;
entity tb_sum_4inputs is
end tb_sum_4inputs;
