//Benchmark atmr_max1024_476_0.5

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n234_, ori_ori_n235_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  INV        o003(.A(ori_ori_n19_), .Y(ori_ori_n20_));
  NA2        o004(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n21_));
  INV        o005(.A(x5), .Y(ori_ori_n22_));
  NA2        o006(.A(x7), .B(x6), .Y(ori_ori_n23_));
  NA2        o007(.A(x4), .B(x2), .Y(ori_ori_n24_));
  INV        o008(.A(ori_ori_n21_), .Y(ori_ori_n25_));
  NO2        o009(.A(x4), .B(x3), .Y(ori_ori_n26_));
  INV        o010(.A(ori_ori_n26_), .Y(ori_ori_n27_));
  NOi21      o011(.An(ori_ori_n20_), .B(ori_ori_n25_), .Y(ori00));
  NO2        o012(.A(x1), .B(x0), .Y(ori_ori_n29_));
  INV        o013(.A(x6), .Y(ori_ori_n30_));
  NA2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  NO2        o015(.A(ori_ori_n20_), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NO2        o016(.A(x2), .B(x0), .Y(ori_ori_n33_));
  INV        o017(.A(x3), .Y(ori_ori_n34_));
  NO2        o018(.A(ori_ori_n34_), .B(ori_ori_n18_), .Y(ori_ori_n35_));
  INV        o019(.A(ori_ori_n35_), .Y(ori_ori_n36_));
  NA2        o020(.A(ori_ori_n36_), .B(ori_ori_n33_), .Y(ori_ori_n37_));
  INV        o021(.A(x4), .Y(ori_ori_n38_));
  NA2        o022(.A(x0), .B(x2), .Y(ori_ori_n39_));
  INV        o023(.A(ori_ori_n37_), .Y(ori_ori_n40_));
  INV        o024(.A(ori_ori_n29_), .Y(ori_ori_n41_));
  INV        o025(.A(x2), .Y(ori_ori_n42_));
  NO2        o026(.A(ori_ori_n42_), .B(ori_ori_n17_), .Y(ori_ori_n43_));
  NA2        o027(.A(ori_ori_n34_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  NA2        o028(.A(ori_ori_n44_), .B(ori_ori_n43_), .Y(ori_ori_n45_));
  OAI210     o029(.A0(ori_ori_n41_), .A1(ori_ori_n27_), .B0(ori_ori_n45_), .Y(ori_ori_n46_));
  NO3        o030(.A(ori_ori_n46_), .B(ori_ori_n40_), .C(ori_ori_n32_), .Y(ori01));
  NA2        o031(.A(ori_ori_n34_), .B(x1), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(x5), .Y(ori_ori_n49_));
  OAI210     o033(.A0(ori_ori_n35_), .A1(ori_ori_n22_), .B0(ori_ori_n42_), .Y(ori_ori_n50_));
  NA2        o034(.A(ori_ori_n50_), .B(x4), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(x2), .Y(ori_ori_n52_));
  OAI210     o036(.A0(ori_ori_n52_), .A1(ori_ori_n44_), .B0(x0), .Y(ori_ori_n53_));
  NA2        o037(.A(x5), .B(x3), .Y(ori_ori_n54_));
  NAi21      o038(.An(x4), .B(x3), .Y(ori_ori_n55_));
  NO2        o039(.A(x4), .B(x2), .Y(ori_ori_n56_));
  NO2        o040(.A(ori_ori_n55_), .B(ori_ori_n18_), .Y(ori_ori_n57_));
  NO2        o041(.A(ori_ori_n57_), .B(ori_ori_n53_), .Y(ori_ori_n58_));
  NA2        o042(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n59_));
  NO2        o043(.A(ori_ori_n59_), .B(ori_ori_n22_), .Y(ori_ori_n60_));
  INV        o044(.A(x8), .Y(ori_ori_n61_));
  AOI210     o045(.A0(ori_ori_n44_), .A1(ori_ori_n22_), .B0(ori_ori_n42_), .Y(ori_ori_n62_));
  NO3        o046(.A(x4), .B(ori_ori_n62_), .C(ori_ori_n60_), .Y(ori_ori_n63_));
  NA2        o047(.A(x4), .B(ori_ori_n34_), .Y(ori_ori_n64_));
  NO2        o048(.A(ori_ori_n64_), .B(x1), .Y(ori_ori_n65_));
  NO2        o049(.A(x3), .B(x2), .Y(ori_ori_n66_));
  NA3        o050(.A(ori_ori_n66_), .B(ori_ori_n23_), .C(ori_ori_n22_), .Y(ori_ori_n67_));
  INV        o051(.A(ori_ori_n67_), .Y(ori_ori_n68_));
  NA2        o052(.A(ori_ori_n42_), .B(x1), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n69_), .A1(ori_ori_n31_), .B0(ori_ori_n17_), .Y(ori_ori_n70_));
  NO4        o054(.A(ori_ori_n70_), .B(ori_ori_n68_), .C(ori_ori_n65_), .D(ori_ori_n63_), .Y(ori_ori_n71_));
  AO210      o055(.A0(ori_ori_n58_), .A1(ori_ori_n51_), .B0(ori_ori_n71_), .Y(ori02));
  NO2        o056(.A(x4), .B(x1), .Y(ori_ori_n73_));
  NA2        o057(.A(ori_ori_n73_), .B(x2), .Y(ori_ori_n74_));
  NO2        o058(.A(ori_ori_n74_), .B(ori_ori_n54_), .Y(ori_ori_n75_));
  NO2        o059(.A(x5), .B(ori_ori_n38_), .Y(ori_ori_n76_));
  NA2        o060(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n77_));
  NO2        o061(.A(ori_ori_n77_), .B(x3), .Y(ori_ori_n78_));
  OAI210     o062(.A0(ori_ori_n78_), .A1(ori_ori_n29_), .B0(ori_ori_n76_), .Y(ori_ori_n79_));
  NO2        o063(.A(ori_ori_n38_), .B(x2), .Y(ori_ori_n80_));
  NA2        o064(.A(ori_ori_n79_), .B(ori_ori_n30_), .Y(ori_ori_n81_));
  NO2        o065(.A(ori_ori_n81_), .B(ori_ori_n75_), .Y(ori_ori_n82_));
  NO3        o066(.A(ori_ori_n54_), .B(ori_ori_n52_), .C(ori_ori_n21_), .Y(ori_ori_n83_));
  NO2        o067(.A(ori_ori_n24_), .B(ori_ori_n22_), .Y(ori_ori_n84_));
  NA2        o068(.A(x7), .B(x3), .Y(ori_ori_n85_));
  NO2        o069(.A(ori_ori_n64_), .B(x5), .Y(ori_ori_n86_));
  INV        o070(.A(x7), .Y(ori_ori_n87_));
  NO2        o071(.A(x4), .B(x2), .Y(ori_ori_n88_));
  INV        o072(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  OAI210     o073(.A0(ori_ori_n85_), .A1(ori_ori_n39_), .B0(ori_ori_n89_), .Y(ori_ori_n90_));
  NAi21      o074(.An(x2), .B(x7), .Y(ori_ori_n91_));
  INV        o075(.A(ori_ori_n91_), .Y(ori_ori_n92_));
  NA2        o076(.A(ori_ori_n92_), .B(ori_ori_n49_), .Y(ori_ori_n93_));
  NA2        o077(.A(ori_ori_n93_), .B(x6), .Y(ori_ori_n94_));
  NO3        o078(.A(ori_ori_n94_), .B(ori_ori_n90_), .C(ori_ori_n83_), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n95_), .B(ori_ori_n82_), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n22_), .B(ori_ori_n18_), .Y(ori_ori_n97_));
  NA2        o081(.A(ori_ori_n22_), .B(ori_ori_n17_), .Y(ori_ori_n98_));
  NA3        o082(.A(ori_ori_n98_), .B(ori_ori_n97_), .C(ori_ori_n21_), .Y(ori_ori_n99_));
  AN2        o083(.A(ori_ori_n99_), .B(ori_ori_n80_), .Y(ori_ori_n100_));
  NO2        o084(.A(ori_ori_n87_), .B(ori_ori_n22_), .Y(ori_ori_n101_));
  NA2        o085(.A(x2), .B(x0), .Y(ori_ori_n102_));
  NA2        o086(.A(x4), .B(x1), .Y(ori_ori_n103_));
  NAi21      o087(.An(ori_ori_n73_), .B(ori_ori_n103_), .Y(ori_ori_n104_));
  NOi21      o088(.An(ori_ori_n104_), .B(ori_ori_n102_), .Y(ori_ori_n105_));
  NO2        o089(.A(ori_ori_n105_), .B(ori_ori_n100_), .Y(ori_ori_n106_));
  NO2        o090(.A(ori_ori_n106_), .B(ori_ori_n34_), .Y(ori_ori_n107_));
  NO2        o091(.A(ori_ori_n99_), .B(ori_ori_n52_), .Y(ori_ori_n108_));
  INV        o092(.A(ori_ori_n76_), .Y(ori_ori_n109_));
  NO2        o093(.A(ori_ori_n69_), .B(ori_ori_n17_), .Y(ori_ori_n110_));
  INV        o094(.A(ori_ori_n110_), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n111_), .B(ori_ori_n109_), .Y(ori_ori_n112_));
  NA3        o096(.A(ori_ori_n104_), .B(ori_ori_n109_), .C(ori_ori_n33_), .Y(ori_ori_n113_));
  INV        o097(.A(ori_ori_n113_), .Y(ori_ori_n114_));
  NO3        o098(.A(ori_ori_n114_), .B(ori_ori_n112_), .C(ori_ori_n108_), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n115_), .B(x3), .Y(ori_ori_n116_));
  NO3        o100(.A(ori_ori_n116_), .B(ori_ori_n107_), .C(ori_ori_n96_), .Y(ori03));
  NO2        o101(.A(ori_ori_n38_), .B(x3), .Y(ori_ori_n118_));
  NO2        o102(.A(ori_ori_n235_), .B(x4), .Y(ori_ori_n119_));
  NO2        o103(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n120_));
  NA2        o104(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n121_));
  NO2        o105(.A(ori_ori_n121_), .B(ori_ori_n97_), .Y(ori_ori_n122_));
  NO3        o106(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n123_));
  NA2        o107(.A(ori_ori_n123_), .B(ori_ori_n38_), .Y(ori_ori_n124_));
  INV        o108(.A(ori_ori_n124_), .Y(ori_ori_n125_));
  NA2        o109(.A(x3), .B(ori_ori_n19_), .Y(ori_ori_n126_));
  NA2        o110(.A(ori_ori_n34_), .B(ori_ori_n42_), .Y(ori_ori_n127_));
  OAI210     o111(.A0(ori_ori_n127_), .A1(ori_ori_n22_), .B0(ori_ori_n98_), .Y(ori_ori_n128_));
  NO2        o112(.A(ori_ori_n103_), .B(x6), .Y(ori_ori_n129_));
  AOI220     o113(.A0(ori_ori_n129_), .A1(ori_ori_n128_), .B0(ori_ori_n80_), .B1(ori_ori_n60_), .Y(ori_ori_n130_));
  NA2        o114(.A(x6), .B(ori_ori_n38_), .Y(ori_ori_n131_));
  INV        o115(.A(x4), .Y(ori_ori_n132_));
  AOI210     o116(.A0(ori_ori_n132_), .A1(ori_ori_n131_), .B0(ori_ori_n54_), .Y(ori_ori_n133_));
  NA3        o117(.A(ori_ori_n121_), .B(ori_ori_n76_), .C(x6), .Y(ori_ori_n134_));
  INV        o118(.A(ori_ori_n49_), .Y(ori_ori_n135_));
  NA2        o119(.A(ori_ori_n135_), .B(ori_ori_n134_), .Y(ori_ori_n136_));
  OAI210     o120(.A0(ori_ori_n136_), .A1(ori_ori_n133_), .B0(x2), .Y(ori_ori_n137_));
  NA3        o121(.A(ori_ori_n137_), .B(ori_ori_n130_), .C(x7), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n125_), .B(ori_ori_n138_), .Y(ori_ori_n139_));
  INV        o123(.A(x3), .Y(ori_ori_n140_));
  NA2        o124(.A(ori_ori_n140_), .B(ori_ori_n119_), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n59_), .B(ori_ori_n22_), .Y(ori_ori_n142_));
  INV        o126(.A(ori_ori_n142_), .Y(ori_ori_n143_));
  AOI210     o127(.A0(ori_ori_n143_), .A1(ori_ori_n141_), .B0(x2), .Y(ori_ori_n144_));
  AOI210     o128(.A0(ori_ori_n119_), .A1(ori_ori_n110_), .B0(ori_ori_n49_), .Y(ori_ori_n145_));
  NA2        o129(.A(ori_ori_n34_), .B(ori_ori_n17_), .Y(ori_ori_n146_));
  NO2        o130(.A(ori_ori_n146_), .B(ori_ori_n22_), .Y(ori_ori_n147_));
  NA2        o131(.A(ori_ori_n147_), .B(ori_ori_n73_), .Y(ori_ori_n148_));
  NA2        o132(.A(ori_ori_n121_), .B(x6), .Y(ori_ori_n149_));
  NA2        o133(.A(ori_ori_n149_), .B(ori_ori_n84_), .Y(ori_ori_n150_));
  NA4        o134(.A(ori_ori_n150_), .B(ori_ori_n148_), .C(ori_ori_n145_), .D(ori_ori_n87_), .Y(ori_ori_n151_));
  AOI210     o135(.A0(x3), .A1(x2), .B0(ori_ori_n38_), .Y(ori_ori_n152_));
  NA2        o136(.A(x6), .B(x2), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n151_), .B(ori_ori_n144_), .Y(ori_ori_n154_));
  OAI210     o138(.A0(x0), .A1(x6), .B0(ori_ori_n35_), .Y(ori_ori_n155_));
  NO2        o139(.A(ori_ori_n155_), .B(ori_ori_n109_), .Y(ori_ori_n156_));
  NOi21      o140(.An(ori_ori_n153_), .B(ori_ori_n17_), .Y(ori_ori_n157_));
  AOI210     o141(.A0(ori_ori_n30_), .A1(ori_ori_n42_), .B0(x0), .Y(ori_ori_n158_));
  NA2        o142(.A(x3), .B(x2), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n158_), .B(ori_ori_n157_), .Y(ori_ori_n160_));
  INV        o144(.A(ori_ori_n122_), .Y(ori_ori_n161_));
  NO2        o145(.A(ori_ori_n131_), .B(ori_ori_n161_), .Y(ori_ori_n162_));
  AO210      o146(.A0(ori_ori_n160_), .A1(ori_ori_n86_), .B0(ori_ori_n162_), .Y(ori_ori_n163_));
  NO2        o147(.A(ori_ori_n163_), .B(ori_ori_n156_), .Y(ori_ori_n164_));
  OAI210     o148(.A0(ori_ori_n154_), .A1(ori_ori_n139_), .B0(ori_ori_n164_), .Y(ori04));
  NO2        o149(.A(x2), .B(x1), .Y(ori_ori_n166_));
  OAI210     o150(.A0(ori_ori_n146_), .A1(ori_ori_n166_), .B0(ori_ori_n30_), .Y(ori_ori_n167_));
  INV        o151(.A(x4), .Y(ori_ori_n168_));
  OAI210     o152(.A0(ori_ori_n42_), .A1(ori_ori_n168_), .B0(ori_ori_n140_), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n159_), .B(ori_ori_n120_), .Y(ori_ori_n170_));
  INV        o154(.A(ori_ori_n170_), .Y(ori_ori_n171_));
  NA3        o155(.A(ori_ori_n171_), .B(x6), .C(ori_ori_n169_), .Y(ori_ori_n172_));
  NA2        o156(.A(ori_ori_n172_), .B(ori_ori_n167_), .Y(ori_ori_n173_));
  NA2        o157(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n174_));
  BUFFER     o158(.A(x4), .Y(ori_ori_n175_));
  XO2        o159(.A(x4), .B(x0), .Y(ori_ori_n176_));
  INV        o160(.A(ori_ori_n175_), .Y(ori_ori_n177_));
  NO2        o161(.A(ori_ori_n177_), .B(x3), .Y(ori_ori_n178_));
  NO2        o162(.A(ori_ori_n61_), .B(x4), .Y(ori_ori_n179_));
  NA2        o163(.A(ori_ori_n179_), .B(ori_ori_n35_), .Y(ori_ori_n180_));
  NO2        o164(.A(ori_ori_n176_), .B(x2), .Y(ori_ori_n181_));
  INV        o165(.A(ori_ori_n181_), .Y(ori_ori_n182_));
  NA4        o166(.A(ori_ori_n182_), .B(ori_ori_n180_), .C(ori_ori_n126_), .D(x6), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n102_), .B(ori_ori_n61_), .Y(ori_ori_n184_));
  NA2        o168(.A(ori_ori_n184_), .B(ori_ori_n48_), .Y(ori_ori_n185_));
  INV        o169(.A(ori_ori_n55_), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n29_), .B(x2), .Y(ori_ori_n187_));
  NA2        o171(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NA2        o172(.A(ori_ori_n185_), .B(ori_ori_n188_), .Y(ori_ori_n189_));
  OAI220     o173(.A0(ori_ori_n189_), .A1(x6), .B0(ori_ori_n183_), .B1(ori_ori_n178_), .Y(ori_ori_n190_));
  AO220      o174(.A0(x7), .A1(ori_ori_n190_), .B0(ori_ori_n234_), .B1(ori_ori_n173_), .Y(ori_ori_n191_));
  NA2        o175(.A(ori_ori_n187_), .B(x6), .Y(ori_ori_n192_));
  NA2        o176(.A(ori_ori_n179_), .B(x0), .Y(ori_ori_n193_));
  NA2        o177(.A(ori_ori_n56_), .B(x6), .Y(ori_ori_n194_));
  OAI210     o178(.A0(ori_ori_n193_), .A1(ori_ori_n34_), .B0(ori_ori_n194_), .Y(ori_ori_n195_));
  NA2        o179(.A(ori_ori_n195_), .B(ori_ori_n192_), .Y(ori_ori_n196_));
  NA2        o180(.A(ori_ori_n196_), .B(ori_ori_n191_), .Y(ori_ori_n197_));
  INV        o181(.A(ori_ori_n174_), .Y(ori_ori_n198_));
  NA2        o182(.A(ori_ori_n198_), .B(ori_ori_n118_), .Y(ori_ori_n199_));
  NA3        o183(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n200_));
  NA2        o184(.A(x3), .B(x0), .Y(ori_ori_n201_));
  OAI220     o185(.A0(ori_ori_n201_), .A1(x2), .B0(ori_ori_n200_), .B1(x1), .Y(ori_ori_n202_));
  INV        o186(.A(ori_ori_n202_), .Y(ori_ori_n203_));
  AOI210     o187(.A0(ori_ori_n203_), .A1(ori_ori_n199_), .B0(ori_ori_n22_), .Y(ori_ori_n204_));
  NA2        o188(.A(ori_ori_n204_), .B(x6), .Y(ori_ori_n205_));
  NAi31      o189(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n206_));
  OAI210     o190(.A0(ori_ori_n206_), .A1(x4), .B0(ori_ori_n91_), .Y(ori_ori_n207_));
  NA2        o191(.A(ori_ori_n207_), .B(ori_ori_n85_), .Y(ori_ori_n208_));
  NA2        o192(.A(ori_ori_n186_), .B(ori_ori_n87_), .Y(ori_ori_n209_));
  NA4        o193(.A(ori_ori_n209_), .B(x1), .C(ori_ori_n208_), .D(ori_ori_n39_), .Y(ori_ori_n210_));
  NA2        o194(.A(x1), .B(ori_ori_n210_), .Y(ori_ori_n211_));
  NO2        o195(.A(x1), .B(x0), .Y(ori_ori_n212_));
  OAI210     o196(.A0(x4), .A1(ori_ori_n34_), .B0(ori_ori_n176_), .Y(ori_ori_n213_));
  INV        o197(.A(ori_ori_n200_), .Y(ori_ori_n214_));
  AOI220     o198(.A0(ori_ori_n214_), .A1(ori_ori_n61_), .B0(ori_ori_n213_), .B1(ori_ori_n87_), .Y(ori_ori_n215_));
  NO2        o199(.A(ori_ori_n215_), .B(ori_ori_n42_), .Y(ori_ori_n216_));
  NO2        o200(.A(ori_ori_n216_), .B(ori_ori_n212_), .Y(ori_ori_n217_));
  AOI210     o201(.A0(ori_ori_n217_), .A1(ori_ori_n211_), .B0(ori_ori_n22_), .Y(ori_ori_n218_));
  NA3        o202(.A(ori_ori_n26_), .B(x2), .C(ori_ori_n17_), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n220_));
  NA2        o204(.A(ori_ori_n220_), .B(ori_ori_n152_), .Y(ori_ori_n221_));
  NO2        o205(.A(ori_ori_n221_), .B(ori_ori_n66_), .Y(ori_ori_n222_));
  NA2        o206(.A(ori_ori_n222_), .B(x7), .Y(ori_ori_n223_));
  NA2        o207(.A(ori_ori_n223_), .B(ori_ori_n219_), .Y(ori_ori_n224_));
  OAI210     o208(.A0(ori_ori_n224_), .A1(ori_ori_n218_), .B0(ori_ori_n30_), .Y(ori_ori_n225_));
  NA2        o209(.A(ori_ori_n206_), .B(ori_ori_n59_), .Y(ori_ori_n226_));
  NA2        o210(.A(ori_ori_n226_), .B(ori_ori_n101_), .Y(ori_ori_n227_));
  NO2        o211(.A(ori_ori_n227_), .B(ori_ori_n131_), .Y(ori_ori_n228_));
  INV        o212(.A(ori_ori_n228_), .Y(ori_ori_n229_));
  NA3        o213(.A(ori_ori_n229_), .B(ori_ori_n225_), .C(ori_ori_n205_), .Y(ori_ori_n230_));
  AOI210     o214(.A0(ori_ori_n197_), .A1(ori_ori_n22_), .B0(ori_ori_n230_), .Y(ori05));
  INV        o215(.A(x7), .Y(ori_ori_n234_));
  INV        o216(.A(x6), .Y(ori_ori_n235_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  INV        m005(.A(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO3        m012(.A(mai_mai_n28_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  NA2        m021(.A(x7), .B(mai_mai_n37_), .Y(mai_mai_n38_));
  NA2        m022(.A(x4), .B(x3), .Y(mai_mai_n39_));
  AOI210     m023(.A0(mai_mai_n38_), .A1(mai_mai_n23_), .B0(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(x2), .B(x0), .Y(mai_mai_n41_));
  INV        m025(.A(x3), .Y(mai_mai_n42_));
  NO2        m026(.A(mai_mai_n42_), .B(mai_mai_n18_), .Y(mai_mai_n43_));
  INV        m027(.A(mai_mai_n43_), .Y(mai_mai_n44_));
  NO2        m028(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n45_));
  OAI210     m029(.A0(mai_mai_n45_), .A1(mai_mai_n44_), .B0(mai_mai_n41_), .Y(mai_mai_n46_));
  INV        m030(.A(x4), .Y(mai_mai_n47_));
  NO2        m031(.A(mai_mai_n47_), .B(mai_mai_n17_), .Y(mai_mai_n48_));
  NA2        m032(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n49_));
  OAI210     m033(.A0(mai_mai_n49_), .A1(mai_mai_n20_), .B0(mai_mai_n46_), .Y(mai_mai_n50_));
  INV        m034(.A(x2), .Y(mai_mai_n51_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n17_), .Y(mai_mai_n52_));
  NA2        m036(.A(mai_mai_n42_), .B(mai_mai_n18_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  OAI210     m038(.A0(mai_mai_n21_), .A1(mai_mai_n32_), .B0(mai_mai_n54_), .Y(mai_mai_n55_));
  NO3        m039(.A(mai_mai_n55_), .B(mai_mai_n50_), .C(mai_mai_n40_), .Y(mai01));
  NA2        m040(.A(x8), .B(x7), .Y(mai_mai_n57_));
  NA2        m041(.A(mai_mai_n42_), .B(x1), .Y(mai_mai_n58_));
  INV        m042(.A(x9), .Y(mai_mai_n59_));
  NO2        m043(.A(mai_mai_n59_), .B(mai_mai_n36_), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n36_), .B(mai_mai_n58_), .Y(mai_mai_n61_));
  NO2        m045(.A(mai_mai_n58_), .B(x5), .Y(mai_mai_n62_));
  OAI210     m046(.A0(mai_mai_n53_), .A1(mai_mai_n20_), .B0(x2), .Y(mai_mai_n63_));
  NAi31      m047(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n64_));
  NO2        m048(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n65_), .A1(mai_mai_n61_), .B0(x4), .Y(mai_mai_n66_));
  INV        m050(.A(x0), .Y(mai_mai_n67_));
  NA2        m051(.A(x5), .B(x3), .Y(mai_mai_n68_));
  NO2        m052(.A(x8), .B(x6), .Y(mai_mai_n69_));
  NO2        m053(.A(mai_mai_n68_), .B(mai_mai_n51_), .Y(mai_mai_n70_));
  NAi21      m054(.An(x4), .B(x3), .Y(mai_mai_n71_));
  INV        m055(.A(mai_mai_n71_), .Y(mai_mai_n72_));
  NO2        m056(.A(mai_mai_n72_), .B(mai_mai_n22_), .Y(mai_mai_n73_));
  NO2        m057(.A(x4), .B(x2), .Y(mai_mai_n74_));
  NO2        m058(.A(mai_mai_n74_), .B(x3), .Y(mai_mai_n75_));
  NO3        m059(.A(mai_mai_n75_), .B(mai_mai_n73_), .C(mai_mai_n18_), .Y(mai_mai_n76_));
  NO3        m060(.A(mai_mai_n76_), .B(mai_mai_n70_), .C(mai_mai_n67_), .Y(mai_mai_n77_));
  NO4        m061(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n42_), .D(x1), .Y(mai_mai_n78_));
  NA2        m062(.A(mai_mai_n78_), .B(mai_mai_n47_), .Y(mai_mai_n79_));
  NA2        m063(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n80_), .B(mai_mai_n25_), .Y(mai_mai_n81_));
  INV        m065(.A(x8), .Y(mai_mai_n82_));
  NA2        m066(.A(x2), .B(x1), .Y(mai_mai_n83_));
  NO2        m067(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(mai_mai_n81_), .Y(mai_mai_n85_));
  NO2        m069(.A(mai_mai_n85_), .B(mai_mai_n26_), .Y(mai_mai_n86_));
  AOI210     m070(.A0(mai_mai_n53_), .A1(mai_mai_n25_), .B0(mai_mai_n51_), .Y(mai_mai_n87_));
  OAI210     m071(.A0(mai_mai_n44_), .A1(mai_mai_n37_), .B0(mai_mai_n47_), .Y(mai_mai_n88_));
  NO3        m072(.A(mai_mai_n88_), .B(mai_mai_n87_), .C(mai_mai_n86_), .Y(mai_mai_n89_));
  NA2        m073(.A(x4), .B(mai_mai_n42_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n47_), .B(mai_mai_n51_), .Y(mai_mai_n91_));
  OAI210     m075(.A0(mai_mai_n91_), .A1(mai_mai_n42_), .B0(mai_mai_n18_), .Y(mai_mai_n92_));
  AOI210     m076(.A0(mai_mai_n90_), .A1(mai_mai_n36_), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  NO2        m077(.A(x3), .B(x2), .Y(mai_mai_n94_));
  NA2        m078(.A(mai_mai_n94_), .B(mai_mai_n25_), .Y(mai_mai_n95_));
  AOI210     m079(.A0(x8), .A1(x6), .B0(mai_mai_n95_), .Y(mai_mai_n96_));
  NA2        m080(.A(mai_mai_n51_), .B(x1), .Y(mai_mai_n97_));
  NO4        m081(.A(x0), .B(mai_mai_n96_), .C(mai_mai_n93_), .D(mai_mai_n89_), .Y(mai_mai_n98_));
  AO220      m082(.A0(mai_mai_n98_), .A1(mai_mai_n79_), .B0(mai_mai_n77_), .B1(mai_mai_n66_), .Y(mai02));
  NO2        m083(.A(x3), .B(mai_mai_n51_), .Y(mai_mai_n100_));
  NO2        m084(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n101_));
  NO3        m085(.A(x8), .B(x7), .C(x5), .Y(mai_mai_n102_));
  NA2        m086(.A(x9), .B(x2), .Y(mai_mai_n103_));
  OR2        m087(.A(x8), .B(x0), .Y(mai_mai_n104_));
  INV        m088(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NAi21      m089(.An(x2), .B(x8), .Y(mai_mai_n106_));
  NO2        m090(.A(x4), .B(x1), .Y(mai_mai_n107_));
  NOi21      m091(.An(x0), .B(x1), .Y(mai_mai_n108_));
  NO3        m092(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n109_));
  NOi21      m093(.An(x0), .B(x4), .Y(mai_mai_n110_));
  AOI220     m094(.A0(mai_mai_n354_), .A1(mai_mai_n110_), .B0(mai_mai_n109_), .B1(mai_mai_n108_), .Y(mai_mai_n111_));
  NO2        m095(.A(mai_mai_n111_), .B(mai_mai_n68_), .Y(mai_mai_n112_));
  NO2        m096(.A(x5), .B(mai_mai_n47_), .Y(mai_mai_n113_));
  OAI210     m097(.A0(mai_mai_n42_), .A1(mai_mai_n35_), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  NAi21      m098(.An(x0), .B(x4), .Y(mai_mai_n115_));
  NO2        m099(.A(mai_mai_n115_), .B(x1), .Y(mai_mai_n116_));
  NO2        m100(.A(x7), .B(x0), .Y(mai_mai_n117_));
  NO2        m101(.A(mai_mai_n74_), .B(mai_mai_n91_), .Y(mai_mai_n118_));
  OAI210     m102(.A0(mai_mai_n117_), .A1(mai_mai_n116_), .B0(mai_mai_n358_), .Y(mai_mai_n119_));
  NO2        m103(.A(mai_mai_n21_), .B(mai_mai_n42_), .Y(mai_mai_n120_));
  NA2        m104(.A(x5), .B(x0), .Y(mai_mai_n121_));
  NO2        m105(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n122_));
  NA2        m106(.A(mai_mai_n122_), .B(mai_mai_n120_), .Y(mai_mai_n123_));
  NA4        m107(.A(mai_mai_n123_), .B(mai_mai_n119_), .C(mai_mai_n114_), .D(mai_mai_n36_), .Y(mai_mai_n124_));
  NO3        m108(.A(mai_mai_n124_), .B(mai_mai_n112_), .C(mai_mai_n102_), .Y(mai_mai_n125_));
  AOI220     m109(.A0(mai_mai_n108_), .A1(x4), .B0(mai_mai_n62_), .B1(mai_mai_n17_), .Y(mai_mai_n126_));
  NO2        m110(.A(mai_mai_n126_), .B(mai_mai_n57_), .Y(mai_mai_n127_));
  NO2        m111(.A(mai_mai_n90_), .B(x5), .Y(mai_mai_n128_));
  NO2        m112(.A(x9), .B(x7), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n42_), .B(x2), .Y(mai_mai_n130_));
  INV        m114(.A(x7), .Y(mai_mai_n131_));
  AOI220     m115(.A0(x7), .A1(mai_mai_n130_), .B0(mai_mai_n100_), .B1(x7), .Y(mai_mai_n132_));
  NO2        m116(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n133_), .B(mai_mai_n110_), .Y(mai_mai_n134_));
  NO2        m118(.A(mai_mai_n134_), .B(mai_mai_n132_), .Y(mai_mai_n135_));
  NA2        m119(.A(x5), .B(x1), .Y(mai_mai_n136_));
  INV        m120(.A(mai_mai_n136_), .Y(mai_mai_n137_));
  AOI210     m121(.A0(mai_mai_n137_), .A1(mai_mai_n110_), .B0(mai_mai_n36_), .Y(mai_mai_n138_));
  NAi31      m122(.An(mai_mai_n68_), .B(x7), .C(mai_mai_n35_), .Y(mai_mai_n139_));
  NA2        m123(.A(mai_mai_n139_), .B(mai_mai_n138_), .Y(mai_mai_n140_));
  NO3        m124(.A(mai_mai_n140_), .B(mai_mai_n135_), .C(mai_mai_n127_), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n141_), .B(mai_mai_n125_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n121_), .B(mai_mai_n118_), .Y(mai_mai_n143_));
  NA2        m127(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n144_));
  NA2        m128(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n145_));
  NA2        m129(.A(x8), .B(x0), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n131_), .B(mai_mai_n25_), .Y(mai_mai_n147_));
  NO2        m131(.A(mai_mai_n108_), .B(x4), .Y(mai_mai_n148_));
  NA2        m132(.A(mai_mai_n148_), .B(mai_mai_n147_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n146_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  NA2        m134(.A(x2), .B(x0), .Y(mai_mai_n151_));
  NA2        m135(.A(x4), .B(x1), .Y(mai_mai_n152_));
  NAi21      m136(.An(mai_mai_n107_), .B(mai_mai_n152_), .Y(mai_mai_n153_));
  NOi31      m137(.An(mai_mai_n153_), .B(mai_mai_n133_), .C(mai_mai_n151_), .Y(mai_mai_n154_));
  NO3        m138(.A(mai_mai_n154_), .B(mai_mai_n150_), .C(mai_mai_n143_), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n155_), .B(mai_mai_n42_), .Y(mai_mai_n156_));
  INV        m140(.A(mai_mai_n113_), .Y(mai_mai_n157_));
  NA2        m141(.A(mai_mai_n153_), .B(mai_mai_n41_), .Y(mai_mai_n158_));
  NA2        m142(.A(mai_mai_n145_), .B(mai_mai_n158_), .Y(mai_mai_n159_));
  INV        m143(.A(mai_mai_n159_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(x3), .Y(mai_mai_n161_));
  NO3        m145(.A(mai_mai_n161_), .B(mai_mai_n156_), .C(mai_mai_n142_), .Y(mai03));
  NO2        m146(.A(mai_mai_n47_), .B(x3), .Y(mai_mai_n163_));
  NO2        m147(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n51_), .B(x1), .Y(mai_mai_n165_));
  OAI210     m149(.A0(mai_mai_n165_), .A1(mai_mai_n25_), .B0(mai_mai_n60_), .Y(mai_mai_n166_));
  NO2        m150(.A(mai_mai_n166_), .B(mai_mai_n17_), .Y(mai_mai_n167_));
  NA2        m151(.A(mai_mai_n167_), .B(mai_mai_n163_), .Y(mai_mai_n168_));
  NO2        m152(.A(mai_mai_n68_), .B(x6), .Y(mai_mai_n169_));
  NA2        m153(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n170_));
  NO2        m154(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n171_));
  NO2        m155(.A(mai_mai_n357_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  INV        m156(.A(mai_mai_n172_), .Y(mai_mai_n173_));
  NO3        m157(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n174_));
  NO2        m158(.A(x5), .B(x1), .Y(mai_mai_n175_));
  AOI220     m159(.A0(mai_mai_n175_), .A1(mai_mai_n17_), .B0(mai_mai_n94_), .B1(x5), .Y(mai_mai_n176_));
  NO3        m160(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n177_));
  NA2        m161(.A(mai_mai_n353_), .B(mai_mai_n47_), .Y(mai_mai_n178_));
  NA3        m162(.A(mai_mai_n178_), .B(mai_mai_n173_), .C(mai_mai_n168_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n47_), .B(mai_mai_n42_), .Y(mai_mai_n180_));
  NA2        m164(.A(mai_mai_n180_), .B(mai_mai_n19_), .Y(mai_mai_n181_));
  NO2        m165(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n182_));
  NO2        m166(.A(mai_mai_n182_), .B(x6), .Y(mai_mai_n183_));
  NOi21      m167(.An(mai_mai_n74_), .B(mai_mai_n183_), .Y(mai_mai_n184_));
  NO2        m168(.A(mai_mai_n184_), .B(mai_mai_n131_), .Y(mai_mai_n185_));
  AO210      m169(.A0(mai_mai_n185_), .A1(mai_mai_n181_), .B0(mai_mai_n147_), .Y(mai_mai_n186_));
  NA2        m170(.A(mai_mai_n42_), .B(mai_mai_n51_), .Y(mai_mai_n187_));
  NA2        m171(.A(mai_mai_n122_), .B(mai_mai_n81_), .Y(mai_mai_n188_));
  NA2        m172(.A(x6), .B(mai_mai_n47_), .Y(mai_mai_n189_));
  AOI210     m173(.A0(mai_mai_n104_), .A1(mai_mai_n189_), .B0(mai_mai_n68_), .Y(mai_mai_n190_));
  NA2        m174(.A(mai_mai_n164_), .B(mai_mai_n116_), .Y(mai_mai_n191_));
  NA2        m175(.A(mai_mai_n191_), .B(mai_mai_n144_), .Y(mai_mai_n192_));
  OAI210     m176(.A0(mai_mai_n192_), .A1(mai_mai_n190_), .B0(x2), .Y(mai_mai_n193_));
  NA3        m177(.A(mai_mai_n193_), .B(mai_mai_n188_), .C(mai_mai_n186_), .Y(mai_mai_n194_));
  AOI210     m178(.A0(mai_mai_n179_), .A1(x8), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  NA2        m179(.A(mai_mai_n183_), .B(mai_mai_n133_), .Y(mai_mai_n196_));
  NO2        m180(.A(mai_mai_n196_), .B(x2), .Y(mai_mai_n197_));
  NO2        m181(.A(x4), .B(mai_mai_n51_), .Y(mai_mai_n198_));
  NA2        m182(.A(mai_mai_n198_), .B(mai_mai_n62_), .Y(mai_mai_n199_));
  NA2        m183(.A(mai_mai_n42_), .B(mai_mai_n17_), .Y(mai_mai_n200_));
  OAI210     m184(.A0(x5), .A1(x3), .B0(mai_mai_n107_), .Y(mai_mai_n201_));
  NA3        m185(.A(mai_mai_n201_), .B(mai_mai_n199_), .C(mai_mai_n131_), .Y(mai_mai_n202_));
  NA2        m186(.A(mai_mai_n164_), .B(mai_mai_n182_), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n121_), .B(mai_mai_n18_), .Y(mai_mai_n204_));
  BUFFER     m188(.A(mai_mai_n204_), .Y(mai_mai_n205_));
  NO2        m189(.A(mai_mai_n47_), .B(mai_mai_n205_), .Y(mai_mai_n206_));
  NA2        m190(.A(mai_mai_n206_), .B(mai_mai_n203_), .Y(mai_mai_n207_));
  NA2        m191(.A(mai_mai_n59_), .B(x2), .Y(mai_mai_n208_));
  NO2        m192(.A(x9), .B(x6), .Y(mai_mai_n209_));
  NA2        m193(.A(x6), .B(x2), .Y(mai_mai_n210_));
  OAI220     m194(.A0(x6), .A1(mai_mai_n42_), .B0(mai_mai_n148_), .B1(mai_mai_n45_), .Y(mai_mai_n211_));
  OAI210     m195(.A0(mai_mai_n211_), .A1(mai_mai_n164_), .B0(mai_mai_n207_), .Y(mai_mai_n212_));
  NA2        m196(.A(x9), .B(mai_mai_n42_), .Y(mai_mai_n213_));
  OR2        m197(.A(mai_mai_n169_), .B(mai_mai_n128_), .Y(mai_mai_n214_));
  NA2        m198(.A(x4), .B(x0), .Y(mai_mai_n215_));
  NA2        m199(.A(mai_mai_n214_), .B(mai_mai_n41_), .Y(mai_mai_n216_));
  AOI210     m200(.A0(mai_mai_n216_), .A1(mai_mai_n212_), .B0(x8), .Y(mai_mai_n217_));
  OAI210     m201(.A0(mai_mai_n204_), .A1(mai_mai_n175_), .B0(x6), .Y(mai_mai_n218_));
  INV        m202(.A(mai_mai_n146_), .Y(mai_mai_n219_));
  OAI210     m203(.A0(mai_mai_n219_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n220_));
  AOI210     m204(.A0(mai_mai_n220_), .A1(mai_mai_n218_), .B0(mai_mai_n187_), .Y(mai_mai_n221_));
  NO4        m205(.A(mai_mai_n221_), .B(mai_mai_n217_), .C(mai_mai_n202_), .D(mai_mai_n197_), .Y(mai_mai_n222_));
  OAI210     m206(.A0(x6), .A1(x3), .B0(x2), .Y(mai_mai_n223_));
  OAI210     m207(.A0(mai_mai_n219_), .A1(x6), .B0(mai_mai_n43_), .Y(mai_mai_n224_));
  AOI210     m208(.A0(mai_mai_n224_), .A1(mai_mai_n223_), .B0(mai_mai_n157_), .Y(mai_mai_n225_));
  NOi21      m209(.An(mai_mai_n210_), .B(mai_mai_n17_), .Y(mai_mai_n226_));
  NA2        m210(.A(mai_mai_n226_), .B(mai_mai_n175_), .Y(mai_mai_n227_));
  AOI210     m211(.A0(mai_mai_n36_), .A1(mai_mai_n51_), .B0(x0), .Y(mai_mai_n228_));
  NA3        m212(.A(mai_mai_n228_), .B(mai_mai_n137_), .C(mai_mai_n32_), .Y(mai_mai_n229_));
  NA2        m213(.A(x3), .B(x2), .Y(mai_mai_n230_));
  AOI220     m214(.A0(mai_mai_n230_), .A1(mai_mai_n187_), .B0(mai_mai_n229_), .B1(mai_mai_n227_), .Y(mai_mai_n231_));
  NAi21      m215(.An(x4), .B(x0), .Y(mai_mai_n232_));
  NO3        m216(.A(mai_mai_n232_), .B(mai_mai_n43_), .C(x2), .Y(mai_mai_n233_));
  OAI210     m217(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n233_), .Y(mai_mai_n234_));
  OAI210     m218(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(x6), .Y(mai_mai_n235_));
  AOI220     m219(.A0(mai_mai_n235_), .A1(mai_mai_n72_), .B0(mai_mai_n18_), .B1(mai_mai_n31_), .Y(mai_mai_n236_));
  AOI210     m220(.A0(mai_mai_n236_), .A1(mai_mai_n234_), .B0(mai_mai_n25_), .Y(mai_mai_n237_));
  NA3        m221(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n238_));
  OAI210     m222(.A0(mai_mai_n228_), .A1(mai_mai_n226_), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NA2        m223(.A(mai_mai_n36_), .B(mai_mai_n42_), .Y(mai_mai_n240_));
  OR2        m224(.A(mai_mai_n240_), .B(mai_mai_n215_), .Y(mai_mai_n241_));
  NO2        m225(.A(mai_mai_n241_), .B(mai_mai_n136_), .Y(mai_mai_n242_));
  AO210      m226(.A0(mai_mai_n239_), .A1(mai_mai_n128_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  NO4        m227(.A(mai_mai_n243_), .B(mai_mai_n237_), .C(mai_mai_n231_), .D(mai_mai_n225_), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n222_), .A1(mai_mai_n195_), .B0(mai_mai_n244_), .Y(mai04));
  NA3        m229(.A(x1), .B(mai_mai_n209_), .C(mai_mai_n75_), .Y(mai_mai_n246_));
  NO2        m230(.A(x2), .B(x1), .Y(mai_mai_n247_));
  OAI210     m231(.A0(mai_mai_n200_), .A1(mai_mai_n247_), .B0(mai_mai_n36_), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n208_), .B(mai_mai_n80_), .Y(mai_mai_n249_));
  NO2        m233(.A(mai_mai_n249_), .B(mai_mai_n36_), .Y(mai_mai_n250_));
  INV        m234(.A(mai_mai_n250_), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n251_), .B(mai_mai_n248_), .Y(mai_mai_n252_));
  NA2        m236(.A(x6), .B(x3), .Y(mai_mai_n253_));
  BUFFER     m237(.A(x8), .Y(mai_mai_n254_));
  AOI210     m238(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n255_));
  OAI220     m239(.A0(mai_mai_n255_), .A1(mai_mai_n240_), .B0(mai_mai_n208_), .B1(mai_mai_n238_), .Y(mai_mai_n256_));
  AOI210     m240(.A0(mai_mai_n254_), .A1(mai_mai_n60_), .B0(mai_mai_n256_), .Y(mai_mai_n257_));
  NA2        m241(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n258_));
  OAI210     m242(.A0(mai_mai_n97_), .A1(mai_mai_n17_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  AOI220     m243(.A0(mai_mai_n259_), .A1(mai_mai_n69_), .B0(mai_mai_n249_), .B1(mai_mai_n82_), .Y(mai_mai_n260_));
  NA3        m244(.A(mai_mai_n260_), .B(mai_mai_n257_), .C(mai_mai_n253_), .Y(mai_mai_n261_));
  OAI210     m245(.A0(mai_mai_n101_), .A1(x3), .B0(mai_mai_n233_), .Y(mai_mai_n262_));
  NA2        m246(.A(mai_mai_n174_), .B(mai_mai_n74_), .Y(mai_mai_n263_));
  NA3        m247(.A(mai_mai_n263_), .B(mai_mai_n262_), .C(mai_mai_n131_), .Y(mai_mai_n264_));
  AOI210     m248(.A0(mai_mai_n261_), .A1(x4), .B0(mai_mai_n264_), .Y(mai_mai_n265_));
  NA2        m249(.A(mai_mai_n356_), .B(mai_mai_n82_), .Y(mai_mai_n266_));
  XO2        m250(.A(x4), .B(x0), .Y(mai_mai_n267_));
  NO2        m251(.A(mai_mai_n267_), .B(mai_mai_n103_), .Y(mai_mai_n268_));
  NA2        m252(.A(mai_mai_n268_), .B(x8), .Y(mai_mai_n269_));
  AOI210     m253(.A0(mai_mai_n269_), .A1(mai_mai_n266_), .B0(x3), .Y(mai_mai_n270_));
  NA2        m254(.A(x8), .B(mai_mai_n43_), .Y(mai_mai_n271_));
  NO2        m255(.A(mai_mai_n28_), .B(mai_mai_n24_), .Y(mai_mai_n272_));
  INV        m256(.A(mai_mai_n272_), .Y(mai_mai_n273_));
  NA4        m257(.A(mai_mai_n273_), .B(mai_mai_n271_), .C(mai_mai_n181_), .D(x6), .Y(mai_mai_n274_));
  NO2        m258(.A(mai_mai_n42_), .B(x0), .Y(mai_mai_n275_));
  NOi21      m259(.An(mai_mai_n107_), .B(mai_mai_n27_), .Y(mai_mai_n276_));
  INV        m260(.A(mai_mai_n276_), .Y(mai_mai_n277_));
  OAI210     m261(.A0(mai_mai_n232_), .A1(mai_mai_n59_), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  OAI220     m262(.A0(mai_mai_n278_), .A1(x6), .B0(mai_mai_n274_), .B1(mai_mai_n270_), .Y(mai_mai_n279_));
  OAI210     m263(.A0(mai_mai_n60_), .A1(mai_mai_n47_), .B0(mai_mai_n41_), .Y(mai_mai_n280_));
  OAI210     m264(.A0(mai_mai_n280_), .A1(mai_mai_n82_), .B0(mai_mai_n241_), .Y(mai_mai_n281_));
  AOI210     m265(.A0(mai_mai_n281_), .A1(mai_mai_n18_), .B0(mai_mai_n131_), .Y(mai_mai_n282_));
  AO220      m266(.A0(mai_mai_n282_), .A1(mai_mai_n279_), .B0(mai_mai_n265_), .B1(mai_mai_n252_), .Y(mai_mai_n283_));
  NA2        m267(.A(mai_mai_n74_), .B(x6), .Y(mai_mai_n284_));
  AOI220     m268(.A0(mai_mai_n351_), .A1(mai_mai_n35_), .B0(mai_mai_n177_), .B1(mai_mai_n48_), .Y(mai_mai_n285_));
  NA3        m269(.A(mai_mai_n285_), .B(mai_mai_n283_), .C(mai_mai_n246_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n165_), .A1(x8), .B0(mai_mai_n101_), .Y(mai_mai_n287_));
  INV        m271(.A(mai_mai_n287_), .Y(mai_mai_n288_));
  NA3        m272(.A(mai_mai_n288_), .B(mai_mai_n163_), .C(mai_mai_n131_), .Y(mai_mai_n289_));
  NA3        m273(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n290_), .B(x2), .Y(mai_mai_n291_));
  AOI210     m275(.A0(mai_mai_n129_), .A1(mai_mai_n105_), .B0(mai_mai_n291_), .Y(mai_mai_n292_));
  AOI210     m276(.A0(mai_mai_n292_), .A1(mai_mai_n289_), .B0(mai_mai_n25_), .Y(mai_mai_n293_));
  NA2        m277(.A(mai_mai_n163_), .B(mai_mai_n171_), .Y(mai_mai_n294_));
  NA3        m278(.A(mai_mai_n165_), .B(mai_mai_n182_), .C(x8), .Y(mai_mai_n295_));
  AOI210     m279(.A0(mai_mai_n295_), .A1(mai_mai_n294_), .B0(mai_mai_n25_), .Y(mai_mai_n296_));
  AOI210     m280(.A0(mai_mai_n106_), .A1(mai_mai_n104_), .B0(mai_mai_n41_), .Y(mai_mai_n297_));
  NOi21      m281(.An(mai_mai_n297_), .B(mai_mai_n152_), .Y(mai_mai_n298_));
  OAI210     m282(.A0(mai_mai_n298_), .A1(mai_mai_n296_), .B0(mai_mai_n129_), .Y(mai_mai_n299_));
  NAi21      m283(.An(mai_mai_n49_), .B(mai_mai_n147_), .Y(mai_mai_n300_));
  NA2        m284(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n301_));
  OAI210     m285(.A0(mai_mai_n301_), .A1(mai_mai_n293_), .B0(x6), .Y(mai_mai_n302_));
  NA3        m286(.A(mai_mai_n52_), .B(x7), .C(mai_mai_n31_), .Y(mai_mai_n303_));
  NO2        m287(.A(mai_mai_n303_), .B(mai_mai_n32_), .Y(mai_mai_n304_));
  NA2        m288(.A(mai_mai_n163_), .B(mai_mai_n131_), .Y(mai_mai_n305_));
  INV        m289(.A(x1), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n305_), .A1(x8), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  NO4        m291(.A(x8), .B(mai_mai_n232_), .C(x9), .D(x2), .Y(mai_mai_n308_));
  NO3        m292(.A(mai_mai_n109_), .B(mai_mai_n308_), .C(mai_mai_n18_), .Y(mai_mai_n309_));
  NO3        m293(.A(x9), .B(mai_mai_n131_), .C(x0), .Y(mai_mai_n310_));
  NA2        m294(.A(mai_mai_n309_), .B(mai_mai_n49_), .Y(mai_mai_n311_));
  OAI210     m295(.A0(mai_mai_n307_), .A1(mai_mai_n304_), .B0(mai_mai_n311_), .Y(mai_mai_n312_));
  AOI210     m296(.A0(x7), .A1(x9), .B0(mai_mai_n115_), .Y(mai_mai_n313_));
  NO3        m297(.A(mai_mai_n313_), .B(mai_mai_n109_), .C(mai_mai_n42_), .Y(mai_mai_n314_));
  NOi31      m298(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n315_));
  NO3        m299(.A(mai_mai_n355_), .B(mai_mai_n314_), .C(x2), .Y(mai_mai_n316_));
  INV        m300(.A(mai_mai_n316_), .Y(mai_mai_n317_));
  AOI210     m301(.A0(mai_mai_n317_), .A1(mai_mai_n312_), .B0(mai_mai_n25_), .Y(mai_mai_n318_));
  NA2        m302(.A(mai_mai_n352_), .B(mai_mai_n297_), .Y(mai_mai_n319_));
  NO2        m303(.A(mai_mai_n319_), .B(mai_mai_n94_), .Y(mai_mai_n320_));
  NO3        m304(.A(mai_mai_n208_), .B(mai_mai_n146_), .C(mai_mai_n39_), .Y(mai_mai_n321_));
  OAI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n320_), .B0(x7), .Y(mai_mai_n322_));
  NA2        m306(.A(x8), .B(x7), .Y(mai_mai_n323_));
  NA3        m307(.A(mai_mai_n323_), .B(mai_mai_n130_), .C(mai_mai_n116_), .Y(mai_mai_n324_));
  NA2        m308(.A(mai_mai_n324_), .B(mai_mai_n322_), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n325_), .A1(mai_mai_n318_), .B0(mai_mai_n36_), .Y(mai_mai_n326_));
  NO2        m310(.A(mai_mai_n310_), .B(mai_mai_n171_), .Y(mai_mai_n327_));
  NO4        m311(.A(mai_mai_n327_), .B(mai_mai_n68_), .C(x4), .D(mai_mai_n51_), .Y(mai_mai_n328_));
  NA2        m312(.A(mai_mai_n200_), .B(mai_mai_n21_), .Y(mai_mai_n329_));
  NO2        m313(.A(mai_mai_n136_), .B(mai_mai_n117_), .Y(mai_mai_n330_));
  NA2        m314(.A(mai_mai_n330_), .B(mai_mai_n329_), .Y(mai_mai_n331_));
  AOI210     m315(.A0(mai_mai_n331_), .A1(mai_mai_n139_), .B0(mai_mai_n28_), .Y(mai_mai_n332_));
  AOI220     m316(.A0(mai_mai_n275_), .A1(mai_mai_n82_), .B0(x8), .B1(mai_mai_n165_), .Y(mai_mai_n333_));
  NA2        m317(.A(mai_mai_n333_), .B(mai_mai_n80_), .Y(mai_mai_n334_));
  NA2        m318(.A(mai_mai_n334_), .B(mai_mai_n147_), .Y(mai_mai_n335_));
  OAI220     m319(.A0(mai_mai_n213_), .A1(x2), .B0(mai_mai_n136_), .B1(mai_mai_n42_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(x2), .A1(mai_mai_n27_), .B0(mai_mai_n64_), .Y(mai_mai_n337_));
  OAI210     m321(.A0(mai_mai_n129_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n338_));
  NO3        m322(.A(mai_mai_n315_), .B(x3), .C(mai_mai_n51_), .Y(mai_mai_n339_));
  AOI210     m323(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n337_), .Y(mai_mai_n340_));
  INV        m324(.A(mai_mai_n340_), .Y(mai_mai_n341_));
  AOI220     m325(.A0(mai_mai_n341_), .A1(x0), .B0(mai_mai_n336_), .B1(mai_mai_n117_), .Y(mai_mai_n342_));
  AOI210     m326(.A0(mai_mai_n342_), .A1(mai_mai_n335_), .B0(mai_mai_n189_), .Y(mai_mai_n343_));
  INV        m327(.A(x5), .Y(mai_mai_n344_));
  NO4        m328(.A(mai_mai_n97_), .B(mai_mai_n344_), .C(mai_mai_n57_), .D(mai_mai_n32_), .Y(mai_mai_n345_));
  NO4        m329(.A(mai_mai_n345_), .B(mai_mai_n343_), .C(mai_mai_n332_), .D(mai_mai_n328_), .Y(mai_mai_n346_));
  NA3        m330(.A(mai_mai_n346_), .B(mai_mai_n326_), .C(mai_mai_n302_), .Y(mai_mai_n347_));
  AOI210     m331(.A0(mai_mai_n286_), .A1(mai_mai_n25_), .B0(mai_mai_n347_), .Y(mai05));
  INV        m332(.A(mai_mai_n284_), .Y(mai_mai_n351_));
  INV        m333(.A(x4), .Y(mai_mai_n352_));
  INV        m334(.A(mai_mai_n176_), .Y(mai_mai_n353_));
  INV        m335(.A(x8), .Y(mai_mai_n354_));
  INV        m336(.A(x3), .Y(mai_mai_n355_));
  INV        m337(.A(x4), .Y(mai_mai_n356_));
  INV        m338(.A(x3), .Y(mai_mai_n357_));
  INV        m339(.A(x3), .Y(mai_mai_n358_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  NAi21      u004(.An(men_men_n20_), .B(men_men_n19_), .Y(men_men_n21_));
  NA2        u005(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n22_));
  INV        u006(.A(x5), .Y(men_men_n23_));
  NA2        u007(.A(x8), .B(x3), .Y(men_men_n24_));
  NA2        u008(.A(x4), .B(x2), .Y(men_men_n25_));
  NO2        u009(.A(men_men_n24_), .B(men_men_n23_), .Y(men_men_n26_));
  NO2        u010(.A(men_men_n26_), .B(men_men_n22_), .Y(men_men_n27_));
  NO2        u011(.A(x4), .B(x3), .Y(men_men_n28_));
  INV        u012(.A(men_men_n28_), .Y(men_men_n29_));
  NOi21      u013(.An(men_men_n21_), .B(men_men_n27_), .Y(men00));
  NO2        u014(.A(x1), .B(x0), .Y(men_men_n31_));
  INV        u015(.A(x6), .Y(men_men_n32_));
  NO2        u016(.A(men_men_n32_), .B(men_men_n23_), .Y(men_men_n33_));
  AN2        u017(.A(x8), .B(x7), .Y(men_men_n34_));
  NA2        u018(.A(men_men_n34_), .B(men_men_n31_), .Y(men_men_n35_));
  NA2        u019(.A(x4), .B(x3), .Y(men_men_n36_));
  AOI210     u020(.A0(men_men_n35_), .A1(men_men_n21_), .B0(men_men_n36_), .Y(men_men_n37_));
  NO2        u021(.A(x2), .B(x0), .Y(men_men_n38_));
  INV        u022(.A(x3), .Y(men_men_n39_));
  NO2        u023(.A(men_men_n39_), .B(men_men_n18_), .Y(men_men_n40_));
  NO2        u024(.A(men_men_n33_), .B(x4), .Y(men_men_n41_));
  NA2        u025(.A(men_men_n41_), .B(men_men_n38_), .Y(men_men_n42_));
  INV        u026(.A(x4), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n44_));
  NA2        u028(.A(men_men_n44_), .B(x2), .Y(men_men_n45_));
  NA2        u029(.A(men_men_n45_), .B(men_men_n42_), .Y(men_men_n46_));
  NA2        u030(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n47_));
  AOI220     u031(.A0(men_men_n47_), .A1(men_men_n31_), .B0(men_men_n20_), .B1(men_men_n19_), .Y(men_men_n48_));
  INV        u032(.A(x2), .Y(men_men_n49_));
  NO2        u033(.A(men_men_n49_), .B(men_men_n17_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n39_), .B(men_men_n18_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  OAI210     u036(.A0(men_men_n48_), .A1(men_men_n29_), .B0(men_men_n52_), .Y(men_men_n53_));
  NO3        u037(.A(men_men_n53_), .B(men_men_n46_), .C(men_men_n37_), .Y(men01));
  NA2        u038(.A(x8), .B(x7), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n39_), .B(x1), .Y(men_men_n56_));
  INV        u040(.A(x9), .Y(men_men_n57_));
  NO2        u041(.A(men_men_n57_), .B(men_men_n32_), .Y(men_men_n58_));
  INV        u042(.A(men_men_n58_), .Y(men_men_n59_));
  NO3        u043(.A(men_men_n59_), .B(men_men_n56_), .C(men_men_n55_), .Y(men_men_n60_));
  NO2        u044(.A(x7), .B(x6), .Y(men_men_n61_));
  NO2        u045(.A(men_men_n56_), .B(x5), .Y(men_men_n62_));
  NO2        u046(.A(x8), .B(x2), .Y(men_men_n63_));
  INV        u047(.A(men_men_n63_), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n64_), .B(x1), .Y(men_men_n65_));
  OA210      u049(.A0(men_men_n65_), .A1(men_men_n62_), .B0(men_men_n61_), .Y(men_men_n66_));
  OAI210     u050(.A0(men_men_n40_), .A1(men_men_n23_), .B0(men_men_n49_), .Y(men_men_n67_));
  NA2        u051(.A(men_men_n51_), .B(men_men_n67_), .Y(men_men_n68_));
  NAi31      u052(.An(x1), .B(x9), .C(x5), .Y(men_men_n69_));
  OAI220     u053(.A0(men_men_n69_), .A1(men_men_n39_), .B0(men_men_n68_), .B1(men_men_n66_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n70_), .A1(men_men_n60_), .B0(x4), .Y(men_men_n71_));
  NA2        u055(.A(men_men_n43_), .B(x2), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n72_), .A1(men_men_n51_), .B0(x0), .Y(men_men_n73_));
  NA2        u057(.A(x5), .B(x3), .Y(men_men_n74_));
  NO2        u058(.A(x8), .B(x6), .Y(men_men_n75_));
  NO4        u059(.A(men_men_n75_), .B(men_men_n74_), .C(men_men_n61_), .D(men_men_n49_), .Y(men_men_n76_));
  NAi21      u060(.An(x4), .B(x3), .Y(men_men_n77_));
  INV        u061(.A(men_men_n77_), .Y(men_men_n78_));
  NO2        u062(.A(men_men_n78_), .B(men_men_n20_), .Y(men_men_n79_));
  NO2        u063(.A(x4), .B(x2), .Y(men_men_n80_));
  NO2        u064(.A(men_men_n80_), .B(x3), .Y(men_men_n81_));
  NO3        u065(.A(men_men_n81_), .B(men_men_n79_), .C(men_men_n18_), .Y(men_men_n82_));
  NO3        u066(.A(men_men_n82_), .B(men_men_n76_), .C(men_men_n73_), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n39_), .B(x1), .Y(men_men_n84_));
  NA2        u068(.A(men_men_n57_), .B(men_men_n43_), .Y(men_men_n85_));
  INV        u069(.A(men_men_n85_), .Y(men_men_n86_));
  OAI210     u070(.A0(men_men_n84_), .A1(men_men_n62_), .B0(men_men_n86_), .Y(men_men_n87_));
  NA2        u071(.A(x3), .B(men_men_n18_), .Y(men_men_n88_));
  INV        u072(.A(x8), .Y(men_men_n89_));
  NA2        u073(.A(x2), .B(x1), .Y(men_men_n90_));
  OAI210     u074(.A0(men_men_n18_), .A1(men_men_n33_), .B0(men_men_n43_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(x2), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n43_), .B(men_men_n49_), .Y(men_men_n93_));
  INV        u077(.A(men_men_n47_), .Y(men_men_n94_));
  NO2        u078(.A(x3), .B(x2), .Y(men_men_n95_));
  NA2        u079(.A(men_men_n49_), .B(x1), .Y(men_men_n96_));
  OAI210     u080(.A0(men_men_n96_), .A1(men_men_n36_), .B0(men_men_n17_), .Y(men_men_n97_));
  NO3        u081(.A(men_men_n97_), .B(men_men_n94_), .C(men_men_n92_), .Y(men_men_n98_));
  AO220      u082(.A0(men_men_n98_), .A1(men_men_n87_), .B0(men_men_n83_), .B1(men_men_n71_), .Y(men02));
  NO2        u083(.A(x3), .B(men_men_n49_), .Y(men_men_n100_));
  NA2        u084(.A(men_men_n49_), .B(men_men_n17_), .Y(men_men_n101_));
  NA2        u085(.A(men_men_n39_), .B(x0), .Y(men_men_n102_));
  OAI210     u086(.A0(men_men_n85_), .A1(men_men_n101_), .B0(men_men_n102_), .Y(men_men_n103_));
  NA2        u087(.A(men_men_n103_), .B(x1), .Y(men_men_n104_));
  NO2        u088(.A(men_men_n104_), .B(x7), .Y(men_men_n105_));
  NA2        u089(.A(x9), .B(x2), .Y(men_men_n106_));
  OR2        u090(.A(x8), .B(x0), .Y(men_men_n107_));
  INV        u091(.A(men_men_n107_), .Y(men_men_n108_));
  NAi21      u092(.An(x2), .B(x8), .Y(men_men_n109_));
  INV        u093(.A(men_men_n109_), .Y(men_men_n110_));
  OAI220     u094(.A0(men_men_n110_), .A1(men_men_n108_), .B0(men_men_n106_), .B1(x7), .Y(men_men_n111_));
  NO2        u095(.A(x4), .B(x1), .Y(men_men_n112_));
  NA3        u096(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n55_), .Y(men_men_n113_));
  NOi21      u097(.An(x0), .B(x1), .Y(men_men_n114_));
  NO3        u098(.A(x9), .B(x8), .C(x7), .Y(men_men_n115_));
  NOi21      u099(.An(x0), .B(x4), .Y(men_men_n116_));
  NAi21      u100(.An(x8), .B(x7), .Y(men_men_n117_));
  NO2        u101(.A(men_men_n117_), .B(men_men_n57_), .Y(men_men_n118_));
  AOI220     u102(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n115_), .B1(men_men_n114_), .Y(men_men_n119_));
  AOI210     u103(.A0(men_men_n119_), .A1(men_men_n113_), .B0(men_men_n74_), .Y(men_men_n120_));
  NO2        u104(.A(x5), .B(men_men_n43_), .Y(men_men_n121_));
  NA2        u105(.A(x2), .B(men_men_n18_), .Y(men_men_n122_));
  NAi21      u106(.An(x0), .B(x4), .Y(men_men_n123_));
  NO2        u107(.A(men_men_n123_), .B(x1), .Y(men_men_n124_));
  NO2        u108(.A(x7), .B(x0), .Y(men_men_n125_));
  NO2        u109(.A(men_men_n80_), .B(men_men_n93_), .Y(men_men_n126_));
  NO2        u110(.A(men_men_n126_), .B(x3), .Y(men_men_n127_));
  OAI210     u111(.A0(men_men_n125_), .A1(men_men_n124_), .B0(men_men_n127_), .Y(men_men_n128_));
  NA2        u112(.A(x5), .B(x0), .Y(men_men_n129_));
  NO2        u113(.A(men_men_n43_), .B(x2), .Y(men_men_n130_));
  NA3        u114(.A(men_men_n130_), .B(men_men_n129_), .C(x3), .Y(men_men_n131_));
  NA3        u115(.A(men_men_n131_), .B(men_men_n128_), .C(men_men_n32_), .Y(men_men_n132_));
  NO3        u116(.A(men_men_n132_), .B(men_men_n120_), .C(men_men_n105_), .Y(men_men_n133_));
  NO3        u117(.A(men_men_n74_), .B(men_men_n72_), .C(men_men_n22_), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n25_), .B(men_men_n23_), .Y(men_men_n135_));
  AOI220     u119(.A0(men_men_n114_), .A1(men_men_n135_), .B0(men_men_n62_), .B1(men_men_n17_), .Y(men_men_n136_));
  NO3        u120(.A(men_men_n136_), .B(men_men_n55_), .C(men_men_n57_), .Y(men_men_n137_));
  NA2        u121(.A(x7), .B(x3), .Y(men_men_n138_));
  NO2        u122(.A(x9), .B(x7), .Y(men_men_n139_));
  NOi21      u123(.An(x8), .B(x0), .Y(men_men_n140_));
  OA210      u124(.A0(men_men_n139_), .A1(x1), .B0(men_men_n140_), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n39_), .B(x2), .Y(men_men_n142_));
  INV        u126(.A(x7), .Y(men_men_n143_));
  AOI220     u127(.A0(x1), .A1(men_men_n142_), .B0(men_men_n100_), .B1(men_men_n34_), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n23_), .B(x4), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n145_), .B(men_men_n116_), .Y(men_men_n146_));
  NO2        u130(.A(men_men_n146_), .B(men_men_n144_), .Y(men_men_n147_));
  AOI210     u131(.A0(men_men_n141_), .A1(x4), .B0(men_men_n147_), .Y(men_men_n148_));
  OAI210     u132(.A0(men_men_n138_), .A1(men_men_n45_), .B0(men_men_n148_), .Y(men_men_n149_));
  NA2        u133(.A(x5), .B(x1), .Y(men_men_n150_));
  INV        u134(.A(men_men_n150_), .Y(men_men_n151_));
  AOI210     u135(.A0(men_men_n151_), .A1(men_men_n116_), .B0(men_men_n32_), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n57_), .B(men_men_n89_), .Y(men_men_n153_));
  NAi21      u137(.An(x2), .B(x7), .Y(men_men_n154_));
  NO3        u138(.A(men_men_n154_), .B(men_men_n153_), .C(men_men_n43_), .Y(men_men_n155_));
  NA2        u139(.A(men_men_n155_), .B(men_men_n62_), .Y(men_men_n156_));
  NAi31      u140(.An(men_men_n74_), .B(men_men_n34_), .C(men_men_n31_), .Y(men_men_n157_));
  NA3        u141(.A(men_men_n157_), .B(men_men_n156_), .C(men_men_n152_), .Y(men_men_n158_));
  NO4        u142(.A(men_men_n158_), .B(men_men_n149_), .C(men_men_n137_), .D(men_men_n134_), .Y(men_men_n159_));
  NO2        u143(.A(men_men_n159_), .B(men_men_n133_), .Y(men_men_n160_));
  NO2        u144(.A(men_men_n129_), .B(men_men_n126_), .Y(men_men_n161_));
  NA2        u145(.A(men_men_n23_), .B(men_men_n18_), .Y(men_men_n162_));
  NA2        u146(.A(men_men_n23_), .B(men_men_n17_), .Y(men_men_n163_));
  NA3        u147(.A(men_men_n163_), .B(men_men_n162_), .C(men_men_n22_), .Y(men_men_n164_));
  AN2        u148(.A(men_men_n164_), .B(men_men_n130_), .Y(men_men_n165_));
  NA2        u149(.A(x8), .B(x0), .Y(men_men_n166_));
  NO2        u150(.A(men_men_n143_), .B(men_men_n23_), .Y(men_men_n167_));
  NO2        u151(.A(men_men_n114_), .B(x4), .Y(men_men_n168_));
  NA2        u152(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  AOI210     u153(.A0(men_men_n166_), .A1(men_men_n122_), .B0(men_men_n169_), .Y(men_men_n170_));
  NA2        u154(.A(x2), .B(x0), .Y(men_men_n171_));
  NA2        u155(.A(x4), .B(x1), .Y(men_men_n172_));
  NO3        u156(.A(men_men_n170_), .B(men_men_n165_), .C(men_men_n161_), .Y(men_men_n173_));
  NO2        u157(.A(men_men_n173_), .B(men_men_n39_), .Y(men_men_n174_));
  NO2        u158(.A(men_men_n164_), .B(men_men_n72_), .Y(men_men_n175_));
  INV        u159(.A(men_men_n121_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n96_), .B(men_men_n17_), .Y(men_men_n177_));
  AOI210     u161(.A0(men_men_n31_), .A1(men_men_n89_), .B0(men_men_n177_), .Y(men_men_n178_));
  NO3        u162(.A(men_men_n178_), .B(men_men_n176_), .C(x7), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n163_), .B(men_men_n126_), .Y(men_men_n180_));
  NO3        u164(.A(men_men_n180_), .B(men_men_n179_), .C(men_men_n175_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n181_), .B(x3), .Y(men_men_n182_));
  NO3        u166(.A(men_men_n182_), .B(men_men_n174_), .C(men_men_n160_), .Y(men03));
  NO2        u167(.A(men_men_n43_), .B(x3), .Y(men_men_n184_));
  NO2        u168(.A(x6), .B(men_men_n23_), .Y(men_men_n185_));
  NA2        u169(.A(men_men_n430_), .B(men_men_n184_), .Y(men_men_n186_));
  NO2        u170(.A(men_men_n74_), .B(x6), .Y(men_men_n187_));
  NA2        u171(.A(x6), .B(men_men_n23_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n188_), .B(x4), .Y(men_men_n189_));
  NO2        u173(.A(men_men_n18_), .B(x0), .Y(men_men_n190_));
  AO220      u174(.A0(men_men_n190_), .A1(men_men_n189_), .B0(men_men_n187_), .B1(men_men_n50_), .Y(men_men_n191_));
  NA2        u175(.A(men_men_n191_), .B(men_men_n57_), .Y(men_men_n192_));
  NA2        u176(.A(x3), .B(men_men_n17_), .Y(men_men_n193_));
  NO2        u177(.A(men_men_n193_), .B(men_men_n188_), .Y(men_men_n194_));
  NA2        u178(.A(x9), .B(men_men_n49_), .Y(men_men_n195_));
  NA2        u179(.A(men_men_n195_), .B(x4), .Y(men_men_n196_));
  NA2        u180(.A(men_men_n188_), .B(men_men_n77_), .Y(men_men_n197_));
  AOI210     u181(.A0(men_men_n23_), .A1(x3), .B0(men_men_n171_), .Y(men_men_n198_));
  AOI220     u182(.A0(men_men_n198_), .A1(men_men_n197_), .B0(men_men_n196_), .B1(men_men_n194_), .Y(men_men_n199_));
  NO2        u183(.A(x5), .B(x1), .Y(men_men_n200_));
  AOI220     u184(.A0(men_men_n200_), .A1(men_men_n17_), .B0(men_men_n95_), .B1(x5), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n193_), .B(men_men_n162_), .Y(men_men_n202_));
  INV        u186(.A(men_men_n202_), .Y(men_men_n203_));
  OAI210     u187(.A0(men_men_n201_), .A1(men_men_n59_), .B0(men_men_n203_), .Y(men_men_n204_));
  AOI220     u188(.A0(men_men_n204_), .A1(men_men_n43_), .B0(x1), .B1(men_men_n121_), .Y(men_men_n205_));
  NA4        u189(.A(men_men_n205_), .B(men_men_n199_), .C(men_men_n192_), .D(men_men_n186_), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n43_), .B(men_men_n39_), .Y(men_men_n207_));
  NO2        u191(.A(x3), .B(men_men_n17_), .Y(men_men_n208_));
  NO2        u192(.A(men_men_n208_), .B(x6), .Y(men_men_n209_));
  NOi21      u193(.An(men_men_n80_), .B(men_men_n209_), .Y(men_men_n210_));
  NA2        u194(.A(men_men_n57_), .B(men_men_n89_), .Y(men_men_n211_));
  NA3        u195(.A(men_men_n211_), .B(men_men_n208_), .C(x6), .Y(men_men_n212_));
  AOI210     u196(.A0(men_men_n212_), .A1(men_men_n210_), .B0(men_men_n143_), .Y(men_men_n213_));
  OR2        u197(.A(men_men_n213_), .B(men_men_n167_), .Y(men_men_n214_));
  NA2        u198(.A(men_men_n39_), .B(men_men_n49_), .Y(men_men_n215_));
  NO3        u199(.A(men_men_n172_), .B(men_men_n57_), .C(x6), .Y(men_men_n216_));
  NA2        u200(.A(x6), .B(men_men_n43_), .Y(men_men_n217_));
  OAI210     u201(.A0(men_men_n108_), .A1(men_men_n75_), .B0(x4), .Y(men_men_n218_));
  NO2        u202(.A(men_men_n218_), .B(men_men_n74_), .Y(men_men_n219_));
  NO2        u203(.A(men_men_n57_), .B(x6), .Y(men_men_n220_));
  OAI210     u204(.A0(x1), .A1(men_men_n202_), .B0(men_men_n220_), .Y(men_men_n221_));
  NA2        u205(.A(men_men_n185_), .B(men_men_n124_), .Y(men_men_n222_));
  NA3        u206(.A(men_men_n193_), .B(men_men_n121_), .C(x6), .Y(men_men_n223_));
  OAI210     u207(.A0(men_men_n89_), .A1(men_men_n32_), .B0(men_men_n62_), .Y(men_men_n224_));
  NA4        u208(.A(men_men_n224_), .B(men_men_n223_), .C(men_men_n222_), .D(men_men_n221_), .Y(men_men_n225_));
  OAI210     u209(.A0(men_men_n225_), .A1(men_men_n219_), .B0(x2), .Y(men_men_n226_));
  NA3        u210(.A(men_men_n226_), .B(men_men_n429_), .C(men_men_n214_), .Y(men_men_n227_));
  AOI210     u211(.A0(men_men_n206_), .A1(x8), .B0(men_men_n227_), .Y(men_men_n228_));
  NO2        u212(.A(men_men_n89_), .B(x3), .Y(men_men_n229_));
  NA2        u213(.A(men_men_n229_), .B(men_men_n189_), .Y(men_men_n230_));
  NO3        u214(.A(men_men_n88_), .B(men_men_n75_), .C(men_men_n23_), .Y(men_men_n231_));
  AOI210     u215(.A0(men_men_n209_), .A1(men_men_n145_), .B0(men_men_n231_), .Y(men_men_n232_));
  AOI210     u216(.A0(men_men_n232_), .A1(men_men_n230_), .B0(x2), .Y(men_men_n233_));
  NO2        u217(.A(x4), .B(men_men_n49_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n189_), .B(men_men_n177_), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n57_), .B(x6), .Y(men_men_n236_));
  NA3        u220(.A(men_men_n23_), .B(x3), .C(x2), .Y(men_men_n237_));
  AOI210     u221(.A0(men_men_n237_), .A1(men_men_n129_), .B0(men_men_n236_), .Y(men_men_n238_));
  NA2        u222(.A(men_men_n238_), .B(men_men_n112_), .Y(men_men_n239_));
  NO2        u223(.A(men_men_n193_), .B(x6), .Y(men_men_n240_));
  NAi21      u224(.An(men_men_n153_), .B(men_men_n240_), .Y(men_men_n241_));
  NA2        u225(.A(men_men_n241_), .B(men_men_n135_), .Y(men_men_n242_));
  NA4        u226(.A(men_men_n242_), .B(men_men_n239_), .C(men_men_n235_), .D(men_men_n143_), .Y(men_men_n243_));
  NA2        u227(.A(men_men_n185_), .B(men_men_n208_), .Y(men_men_n244_));
  NO2        u228(.A(x9), .B(x6), .Y(men_men_n245_));
  NO2        u229(.A(men_men_n129_), .B(men_men_n18_), .Y(men_men_n246_));
  NAi21      u230(.An(men_men_n246_), .B(men_men_n237_), .Y(men_men_n247_));
  NAi21      u231(.An(x1), .B(x4), .Y(men_men_n248_));
  OAI210     u232(.A0(men_men_n129_), .A1(x3), .B0(x4), .Y(men_men_n249_));
  AOI220     u233(.A0(men_men_n249_), .A1(men_men_n248_), .B0(men_men_n247_), .B1(men_men_n245_), .Y(men_men_n250_));
  NA2        u234(.A(men_men_n250_), .B(men_men_n244_), .Y(men_men_n251_));
  NA2        u235(.A(men_men_n57_), .B(x2), .Y(men_men_n252_));
  NO2        u236(.A(men_men_n252_), .B(men_men_n244_), .Y(men_men_n253_));
  NO3        u237(.A(x9), .B(x6), .C(x0), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n96_), .B(men_men_n23_), .Y(men_men_n255_));
  NA2        u239(.A(x6), .B(x2), .Y(men_men_n256_));
  NO2        u240(.A(men_men_n256_), .B(men_men_n162_), .Y(men_men_n257_));
  AOI210     u241(.A0(men_men_n255_), .A1(men_men_n254_), .B0(men_men_n257_), .Y(men_men_n258_));
  OAI220     u242(.A0(men_men_n258_), .A1(men_men_n39_), .B0(men_men_n168_), .B1(men_men_n41_), .Y(men_men_n259_));
  OAI210     u243(.A0(men_men_n259_), .A1(men_men_n253_), .B0(men_men_n251_), .Y(men_men_n260_));
  NO2        u244(.A(men_men_n427_), .B(men_men_n188_), .Y(men_men_n261_));
  OR2        u245(.A(men_men_n261_), .B(x4), .Y(men_men_n262_));
  NA2        u246(.A(x4), .B(x0), .Y(men_men_n263_));
  NO3        u247(.A(men_men_n69_), .B(men_men_n263_), .C(x6), .Y(men_men_n264_));
  AOI210     u248(.A0(men_men_n262_), .A1(men_men_n38_), .B0(men_men_n264_), .Y(men_men_n265_));
  AOI210     u249(.A0(men_men_n265_), .A1(men_men_n260_), .B0(x8), .Y(men_men_n266_));
  INV        u250(.A(men_men_n236_), .Y(men_men_n267_));
  OAI210     u251(.A0(men_men_n246_), .A1(men_men_n200_), .B0(men_men_n267_), .Y(men_men_n268_));
  NO2        u252(.A(men_men_n268_), .B(men_men_n215_), .Y(men_men_n269_));
  NO4        u253(.A(men_men_n269_), .B(men_men_n266_), .C(men_men_n243_), .D(men_men_n233_), .Y(men_men_n270_));
  NO2        u254(.A(men_men_n153_), .B(x1), .Y(men_men_n271_));
  NO3        u255(.A(men_men_n271_), .B(x3), .C(men_men_n32_), .Y(men_men_n272_));
  OAI210     u256(.A0(men_men_n272_), .A1(men_men_n240_), .B0(x2), .Y(men_men_n273_));
  NO2        u257(.A(men_men_n273_), .B(men_men_n176_), .Y(men_men_n274_));
  NOi21      u258(.An(men_men_n256_), .B(men_men_n17_), .Y(men_men_n275_));
  NA3        u259(.A(men_men_n275_), .B(men_men_n200_), .C(men_men_n36_), .Y(men_men_n276_));
  AOI210     u260(.A0(men_men_n32_), .A1(men_men_n49_), .B0(x0), .Y(men_men_n277_));
  NA3        u261(.A(men_men_n277_), .B(men_men_n151_), .C(men_men_n29_), .Y(men_men_n278_));
  NA2        u262(.A(x3), .B(x2), .Y(men_men_n279_));
  AOI220     u263(.A0(men_men_n279_), .A1(men_men_n215_), .B0(men_men_n278_), .B1(men_men_n276_), .Y(men_men_n280_));
  NAi21      u264(.An(x4), .B(x0), .Y(men_men_n281_));
  NO3        u265(.A(men_men_n281_), .B(men_men_n40_), .C(x2), .Y(men_men_n282_));
  OAI210     u266(.A0(x6), .A1(men_men_n18_), .B0(men_men_n282_), .Y(men_men_n283_));
  OAI220     u267(.A0(men_men_n22_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n284_));
  NO2        u268(.A(x9), .B(x8), .Y(men_men_n285_));
  NA3        u269(.A(men_men_n285_), .B(men_men_n32_), .C(men_men_n49_), .Y(men_men_n286_));
  OAI210     u270(.A0(men_men_n277_), .A1(men_men_n275_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI220     u271(.A0(men_men_n287_), .A1(men_men_n78_), .B0(men_men_n284_), .B1(men_men_n28_), .Y(men_men_n288_));
  AOI210     u272(.A0(men_men_n288_), .A1(men_men_n283_), .B0(men_men_n23_), .Y(men_men_n289_));
  NA2        u273(.A(men_men_n32_), .B(men_men_n39_), .Y(men_men_n290_));
  OR2        u274(.A(men_men_n290_), .B(men_men_n263_), .Y(men_men_n291_));
  NO2        u275(.A(men_men_n291_), .B(men_men_n150_), .Y(men_men_n292_));
  NO4        u276(.A(men_men_n292_), .B(men_men_n289_), .C(men_men_n280_), .D(men_men_n274_), .Y(men_men_n293_));
  OAI210     u277(.A0(men_men_n270_), .A1(men_men_n228_), .B0(men_men_n293_), .Y(men04));
  OAI210     u278(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n295_));
  NA3        u279(.A(men_men_n295_), .B(men_men_n254_), .C(men_men_n81_), .Y(men_men_n296_));
  NO2        u280(.A(x2), .B(x1), .Y(men_men_n297_));
  NO2        u281(.A(men_men_n297_), .B(men_men_n281_), .Y(men_men_n298_));
  NO2        u282(.A(men_men_n279_), .B(men_men_n190_), .Y(men_men_n299_));
  NA2        u283(.A(x9), .B(x0), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n88_), .A1(men_men_n72_), .B0(men_men_n300_), .Y(men_men_n301_));
  OAI210     u285(.A0(men_men_n301_), .A1(men_men_n299_), .B0(men_men_n89_), .Y(men_men_n302_));
  NO2        u286(.A(men_men_n195_), .B(men_men_n102_), .Y(men_men_n303_));
  NO3        u287(.A(men_men_n236_), .B(men_men_n109_), .C(men_men_n18_), .Y(men_men_n304_));
  NO2        u288(.A(men_men_n304_), .B(men_men_n303_), .Y(men_men_n305_));
  OAI210     u289(.A0(men_men_n107_), .A1(men_men_n96_), .B0(men_men_n166_), .Y(men_men_n306_));
  NA3        u290(.A(men_men_n306_), .B(x6), .C(x3), .Y(men_men_n307_));
  NOi21      u291(.An(men_men_n140_), .B(men_men_n122_), .Y(men_men_n308_));
  AOI210     u292(.A0(men_men_n308_), .A1(men_men_n58_), .B0(men_men_n32_), .Y(men_men_n309_));
  NA3        u293(.A(men_men_n309_), .B(men_men_n307_), .C(men_men_n305_), .Y(men_men_n310_));
  OAI210     u294(.A0(x1), .A1(x3), .B0(men_men_n282_), .Y(men_men_n311_));
  NA3        u295(.A(men_men_n211_), .B(x1), .C(men_men_n80_), .Y(men_men_n312_));
  NA3        u296(.A(men_men_n312_), .B(men_men_n311_), .C(men_men_n143_), .Y(men_men_n313_));
  AOI210     u297(.A0(men_men_n310_), .A1(x4), .B0(men_men_n313_), .Y(men_men_n314_));
  NA3        u298(.A(men_men_n298_), .B(men_men_n195_), .C(men_men_n89_), .Y(men_men_n315_));
  NOi21      u299(.An(x4), .B(x0), .Y(men_men_n316_));
  XO2        u300(.A(x4), .B(x0), .Y(men_men_n317_));
  OAI210     u301(.A0(men_men_n317_), .A1(men_men_n106_), .B0(men_men_n248_), .Y(men_men_n318_));
  AOI220     u302(.A0(men_men_n318_), .A1(x8), .B0(men_men_n316_), .B1(men_men_n90_), .Y(men_men_n319_));
  AOI210     u303(.A0(men_men_n319_), .A1(men_men_n315_), .B0(x3), .Y(men_men_n320_));
  INV        u304(.A(men_men_n90_), .Y(men_men_n321_));
  NO2        u305(.A(men_men_n89_), .B(x4), .Y(men_men_n322_));
  NA2        u306(.A(men_men_n116_), .B(men_men_n321_), .Y(men_men_n323_));
  NO3        u307(.A(men_men_n317_), .B(men_men_n153_), .C(x2), .Y(men_men_n324_));
  NO3        u308(.A(men_men_n211_), .B(men_men_n25_), .C(men_men_n22_), .Y(men_men_n325_));
  NO2        u309(.A(men_men_n325_), .B(men_men_n324_), .Y(men_men_n326_));
  NA3        u310(.A(men_men_n326_), .B(men_men_n323_), .C(x6), .Y(men_men_n327_));
  OAI220     u311(.A0(men_men_n281_), .A1(men_men_n88_), .B0(men_men_n171_), .B1(men_men_n89_), .Y(men_men_n328_));
  OR2        u312(.A(men_men_n322_), .B(x3), .Y(men_men_n329_));
  NO2        u313(.A(men_men_n140_), .B(men_men_n96_), .Y(men_men_n330_));
  AOI220     u314(.A0(men_men_n330_), .A1(men_men_n329_), .B0(men_men_n328_), .B1(men_men_n56_), .Y(men_men_n331_));
  NO2        u315(.A(men_men_n140_), .B(men_men_n77_), .Y(men_men_n332_));
  NOi21      u316(.An(men_men_n112_), .B(men_men_n24_), .Y(men_men_n333_));
  AOI210     u317(.A0(men_men_n428_), .A1(men_men_n332_), .B0(men_men_n333_), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n331_), .A1(men_men_n57_), .B0(men_men_n334_), .Y(men_men_n335_));
  OAI220     u319(.A0(men_men_n335_), .A1(x6), .B0(men_men_n327_), .B1(men_men_n320_), .Y(men_men_n336_));
  OAI210     u320(.A0(men_men_n426_), .A1(men_men_n89_), .B0(men_men_n291_), .Y(men_men_n337_));
  AOI210     u321(.A0(men_men_n337_), .A1(men_men_n18_), .B0(men_men_n143_), .Y(men_men_n338_));
  AO220      u322(.A0(men_men_n338_), .A1(men_men_n336_), .B0(men_men_n314_), .B1(men_men_n302_), .Y(men_men_n339_));
  NA2        u323(.A(x6), .B(x1), .Y(men_men_n340_));
  NA2        u324(.A(men_men_n322_), .B(x0), .Y(men_men_n341_));
  NO2        u325(.A(men_men_n341_), .B(men_men_n340_), .Y(men_men_n342_));
  INV        u326(.A(men_men_n342_), .Y(men_men_n343_));
  NA3        u327(.A(men_men_n343_), .B(men_men_n339_), .C(men_men_n296_), .Y(men_men_n344_));
  NA2        u328(.A(men_men_n184_), .B(men_men_n143_), .Y(men_men_n345_));
  OAI210     u329(.A0(men_men_n25_), .A1(x1), .B0(men_men_n215_), .Y(men_men_n346_));
  AO220      u330(.A0(men_men_n346_), .A1(men_men_n139_), .B0(men_men_n100_), .B1(x4), .Y(men_men_n347_));
  NA3        u331(.A(x7), .B(x3), .C(x0), .Y(men_men_n348_));
  NO2        u332(.A(men_men_n43_), .B(men_men_n195_), .Y(men_men_n349_));
  AOI210     u333(.A0(men_men_n347_), .A1(men_men_n108_), .B0(men_men_n349_), .Y(men_men_n350_));
  AOI210     u334(.A0(men_men_n350_), .A1(men_men_n345_), .B0(men_men_n23_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n110_), .B(men_men_n207_), .C(x0), .Y(men_men_n352_));
  OAI210     u336(.A0(men_men_n184_), .A1(men_men_n63_), .B0(men_men_n190_), .Y(men_men_n353_));
  NO2        u337(.A(men_men_n353_), .B(men_men_n23_), .Y(men_men_n354_));
  AOI210     u338(.A0(men_men_n109_), .A1(men_men_n107_), .B0(men_men_n38_), .Y(men_men_n355_));
  NOi31      u339(.An(men_men_n355_), .B(x3), .C(men_men_n172_), .Y(men_men_n356_));
  OAI210     u340(.A0(men_men_n356_), .A1(men_men_n354_), .B0(men_men_n139_), .Y(men_men_n357_));
  NAi31      u341(.An(men_men_n45_), .B(men_men_n271_), .C(men_men_n167_), .Y(men_men_n358_));
  NA3        u342(.A(men_men_n358_), .B(men_men_n357_), .C(men_men_n352_), .Y(men_men_n359_));
  OAI210     u343(.A0(men_men_n359_), .A1(men_men_n351_), .B0(x6), .Y(men_men_n360_));
  OAI210     u344(.A0(men_men_n153_), .A1(men_men_n43_), .B0(men_men_n125_), .Y(men_men_n361_));
  NA3        u345(.A(men_men_n50_), .B(men_men_n34_), .C(men_men_n28_), .Y(men_men_n362_));
  AOI220     u346(.A0(men_men_n362_), .A1(men_men_n361_), .B0(men_men_n36_), .B1(men_men_n29_), .Y(men_men_n363_));
  NO2        u347(.A(men_men_n143_), .B(x0), .Y(men_men_n364_));
  AOI220     u348(.A0(men_men_n364_), .A1(men_men_n207_), .B0(men_men_n184_), .B1(men_men_n143_), .Y(men_men_n365_));
  AOI210     u349(.A0(men_men_n118_), .A1(men_men_n234_), .B0(x1), .Y(men_men_n366_));
  OAI210     u350(.A0(men_men_n365_), .A1(x8), .B0(men_men_n366_), .Y(men_men_n367_));
  NAi31      u351(.An(x2), .B(x8), .C(x0), .Y(men_men_n368_));
  OAI210     u352(.A0(men_men_n368_), .A1(x4), .B0(men_men_n154_), .Y(men_men_n369_));
  NA3        u353(.A(men_men_n369_), .B(men_men_n138_), .C(x9), .Y(men_men_n370_));
  NO4        u354(.A(men_men_n117_), .B(men_men_n281_), .C(x9), .D(x2), .Y(men_men_n371_));
  NOi21      u355(.An(men_men_n115_), .B(men_men_n171_), .Y(men_men_n372_));
  NO3        u356(.A(men_men_n372_), .B(men_men_n371_), .C(men_men_n18_), .Y(men_men_n373_));
  NO3        u357(.A(x9), .B(men_men_n143_), .C(x0), .Y(men_men_n374_));
  AOI220     u358(.A0(men_men_n374_), .A1(men_men_n229_), .B0(men_men_n332_), .B1(men_men_n143_), .Y(men_men_n375_));
  NA4        u359(.A(men_men_n375_), .B(men_men_n373_), .C(men_men_n370_), .D(men_men_n45_), .Y(men_men_n376_));
  OAI210     u360(.A0(men_men_n367_), .A1(men_men_n363_), .B0(men_men_n376_), .Y(men_men_n377_));
  NOi31      u361(.An(men_men_n364_), .B(men_men_n29_), .C(x8), .Y(men_men_n378_));
  AOI210     u362(.A0(men_men_n34_), .A1(x9), .B0(men_men_n123_), .Y(men_men_n379_));
  NO3        u363(.A(men_men_n379_), .B(men_men_n115_), .C(men_men_n39_), .Y(men_men_n380_));
  NOi31      u364(.An(x1), .B(x8), .C(x7), .Y(men_men_n381_));
  AOI220     u365(.A0(men_men_n381_), .A1(men_men_n316_), .B0(men_men_n116_), .B1(x3), .Y(men_men_n382_));
  AOI210     u366(.A0(men_men_n248_), .A1(men_men_n55_), .B0(men_men_n114_), .Y(men_men_n383_));
  OAI210     u367(.A0(men_men_n383_), .A1(x3), .B0(men_men_n382_), .Y(men_men_n384_));
  NO3        u368(.A(men_men_n384_), .B(men_men_n380_), .C(x2), .Y(men_men_n385_));
  OAI220     u369(.A0(men_men_n317_), .A1(men_men_n285_), .B0(men_men_n281_), .B1(men_men_n39_), .Y(men_men_n386_));
  AOI210     u370(.A0(x9), .A1(men_men_n43_), .B0(men_men_n348_), .Y(men_men_n387_));
  AOI220     u371(.A0(men_men_n387_), .A1(men_men_n89_), .B0(men_men_n386_), .B1(men_men_n143_), .Y(men_men_n388_));
  NO2        u372(.A(men_men_n388_), .B(men_men_n49_), .Y(men_men_n389_));
  NO3        u373(.A(men_men_n389_), .B(men_men_n385_), .C(men_men_n378_), .Y(men_men_n390_));
  AOI210     u374(.A0(men_men_n390_), .A1(men_men_n377_), .B0(men_men_n23_), .Y(men_men_n391_));
  NO3        u375(.A(men_men_n57_), .B(x4), .C(x1), .Y(men_men_n392_));
  NO3        u376(.A(men_men_n63_), .B(men_men_n18_), .C(x0), .Y(men_men_n393_));
  AOI220     u377(.A0(men_men_n393_), .A1(x4), .B0(men_men_n392_), .B1(men_men_n355_), .Y(men_men_n394_));
  NO2        u378(.A(men_men_n394_), .B(men_men_n95_), .Y(men_men_n395_));
  NO3        u379(.A(men_men_n252_), .B(men_men_n166_), .C(men_men_n36_), .Y(men_men_n396_));
  OAI210     u380(.A0(men_men_n396_), .A1(men_men_n395_), .B0(x7), .Y(men_men_n397_));
  NA3        u381(.A(men_men_n57_), .B(men_men_n142_), .C(men_men_n124_), .Y(men_men_n398_));
  NA2        u382(.A(men_men_n398_), .B(men_men_n397_), .Y(men_men_n399_));
  OAI210     u383(.A0(men_men_n399_), .A1(men_men_n391_), .B0(men_men_n32_), .Y(men_men_n400_));
  NO2        u384(.A(men_men_n374_), .B(men_men_n190_), .Y(men_men_n401_));
  NO4        u385(.A(men_men_n401_), .B(men_men_n74_), .C(x4), .D(men_men_n49_), .Y(men_men_n402_));
  INV        u386(.A(x7), .Y(men_men_n403_));
  NO2        u387(.A(men_men_n150_), .B(men_men_n125_), .Y(men_men_n404_));
  NA2        u388(.A(men_men_n404_), .B(men_men_n403_), .Y(men_men_n405_));
  AOI210     u389(.A0(men_men_n405_), .A1(men_men_n157_), .B0(men_men_n25_), .Y(men_men_n406_));
  AOI220     u390(.A0(x3), .A1(men_men_n89_), .B0(men_men_n140_), .B1(x2), .Y(men_men_n407_));
  NA2        u391(.A(men_men_n407_), .B(men_men_n368_), .Y(men_men_n408_));
  NA2        u392(.A(men_men_n408_), .B(men_men_n167_), .Y(men_men_n409_));
  OAI220     u393(.A0(men_men_n427_), .A1(men_men_n64_), .B0(men_men_n150_), .B1(men_men_n39_), .Y(men_men_n410_));
  NA2        u394(.A(x3), .B(men_men_n49_), .Y(men_men_n411_));
  AOI210     u395(.A0(men_men_n154_), .A1(men_men_n24_), .B0(men_men_n69_), .Y(men_men_n412_));
  OAI210     u396(.A0(men_men_n139_), .A1(men_men_n18_), .B0(x7), .Y(men_men_n413_));
  NO3        u397(.A(men_men_n381_), .B(x3), .C(men_men_n49_), .Y(men_men_n414_));
  AOI210     u398(.A0(men_men_n414_), .A1(men_men_n413_), .B0(men_men_n412_), .Y(men_men_n415_));
  OAI210     u399(.A0(x1), .A1(men_men_n411_), .B0(men_men_n415_), .Y(men_men_n416_));
  AOI220     u400(.A0(men_men_n416_), .A1(x0), .B0(men_men_n410_), .B1(men_men_n125_), .Y(men_men_n417_));
  AOI210     u401(.A0(men_men_n417_), .A1(men_men_n409_), .B0(men_men_n217_), .Y(men_men_n418_));
  NA2        u402(.A(x9), .B(x5), .Y(men_men_n419_));
  NO4        u403(.A(men_men_n96_), .B(men_men_n419_), .C(men_men_n55_), .D(men_men_n29_), .Y(men_men_n420_));
  NO4        u404(.A(men_men_n420_), .B(men_men_n418_), .C(men_men_n406_), .D(men_men_n402_), .Y(men_men_n421_));
  NA3        u405(.A(men_men_n421_), .B(men_men_n400_), .C(men_men_n360_), .Y(men_men_n422_));
  AOI210     u406(.A0(men_men_n344_), .A1(men_men_n23_), .B0(men_men_n422_), .Y(men05));
  INV        u407(.A(men_men_n38_), .Y(men_men_n426_));
  INV        u408(.A(x9), .Y(men_men_n427_));
  INV        u409(.A(x2), .Y(men_men_n428_));
  INV        u410(.A(men_men_n216_), .Y(men_men_n429_));
  INV        u411(.A(men_men_n23_), .Y(men_men_n430_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule