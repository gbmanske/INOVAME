library verilog;
use verilog.vl_types.all;
entity contador8_vlg_vec_tst is
end contador8_vlg_vec_tst;
