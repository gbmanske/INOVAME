// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n130_, new_new_n131_,
    new_new_n132_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n667_, new_new_n668_, new_new_n669_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n712_, new_new_n713_, new_new_n714_, new_new_n715_,
    new_new_n716_, new_new_n717_, new_new_n718_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n933_, new_new_n934_, new_new_n935_,
    new_new_n936_, new_new_n937_, new_new_n938_, new_new_n939_,
    new_new_n940_, new_new_n941_, new_new_n942_, new_new_n943_,
    new_new_n944_, new_new_n945_, new_new_n946_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA3        g029(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n52_));
  NO2        g030(.A(i_1_), .B(i_6_), .Y(new_new_n53_));
  NA2        g031(.A(i_8_), .B(i_7_), .Y(new_new_n54_));
  OAI210     g032(.A0(new_new_n54_), .A1(new_new_n53_), .B0(new_new_n52_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n55_), .B(i_12_), .Y(new_new_n56_));
  INV        g034(.A(i_1_), .Y(new_new_n57_));
  NA2        g035(.A(i_1_), .B(i_10_), .Y(new_new_n58_));
  NO2        g036(.A(new_new_n58_), .B(i_6_), .Y(new_new_n59_));
  NAi31      g037(.An(new_new_n59_), .B(new_new_n946_), .C(new_new_n56_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n50_), .B(i_2_), .Y(new_new_n61_));
  AOI210     g039(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n62_));
  NA2        g040(.A(i_1_), .B(i_6_), .Y(new_new_n63_));
  NO2        g041(.A(new_new_n63_), .B(new_new_n25_), .Y(new_new_n64_));
  INV        g042(.A(i_0_), .Y(new_new_n65_));
  NAi21      g043(.An(i_5_), .B(i_10_), .Y(new_new_n66_));
  NA2        g044(.A(i_5_), .B(i_9_), .Y(new_new_n67_));
  AOI210     g045(.A0(new_new_n67_), .A1(new_new_n66_), .B0(new_new_n65_), .Y(new_new_n68_));
  NO2        g046(.A(new_new_n68_), .B(new_new_n64_), .Y(new_new_n69_));
  INV        g047(.A(new_new_n69_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n70_), .A1(new_new_n60_), .B0(i_0_), .Y(new_new_n71_));
  NA2        g049(.A(i_12_), .B(i_5_), .Y(new_new_n72_));
  NA2        g050(.A(i_2_), .B(i_8_), .Y(new_new_n73_));
  NO2        g051(.A(new_new_n73_), .B(new_new_n53_), .Y(new_new_n74_));
  NO2        g052(.A(i_3_), .B(i_9_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_7_), .Y(new_new_n76_));
  INV        g054(.A(i_6_), .Y(new_new_n77_));
  OR4        g055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n78_));
  INV        g056(.A(new_new_n78_), .Y(new_new_n79_));
  NO2        g057(.A(i_2_), .B(i_7_), .Y(new_new_n80_));
  NAi21      g058(.An(i_6_), .B(i_10_), .Y(new_new_n81_));
  NA2        g059(.A(i_6_), .B(i_9_), .Y(new_new_n82_));
  AOI210     g060(.A0(new_new_n82_), .A1(new_new_n81_), .B0(new_new_n57_), .Y(new_new_n83_));
  NA2        g061(.A(i_2_), .B(i_6_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n83_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n936_), .B0(new_new_n72_), .Y(new_new_n86_));
  AN3        g064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_11_), .Y(new_new_n88_));
  NO2        g066(.A(i_5_), .B(i_8_), .Y(new_new_n89_));
  NOi21      g067(.An(new_new_n89_), .B(new_new_n88_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n87_), .A1(new_new_n32_), .B0(new_new_n90_), .Y(new_new_n91_));
  INV        g069(.A(i_7_), .Y(new_new_n92_));
  NA2        g070(.A(new_new_n46_), .B(new_new_n92_), .Y(new_new_n93_));
  NO2        g071(.A(i_0_), .B(i_5_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n94_), .B(new_new_n77_), .Y(new_new_n95_));
  NA2        g073(.A(i_12_), .B(i_3_), .Y(new_new_n96_));
  INV        g074(.A(new_new_n96_), .Y(new_new_n97_));
  NA3        g075(.A(new_new_n97_), .B(new_new_n95_), .C(new_new_n93_), .Y(new_new_n98_));
  NAi21      g076(.An(i_7_), .B(i_11_), .Y(new_new_n99_));
  NO3        g077(.A(new_new_n99_), .B(new_new_n81_), .C(new_new_n51_), .Y(new_new_n100_));
  AN2        g078(.A(i_2_), .B(i_10_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(i_7_), .Y(new_new_n102_));
  OR2        g080(.A(new_new_n72_), .B(new_new_n53_), .Y(new_new_n103_));
  NO2        g081(.A(i_8_), .B(new_new_n92_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n103_), .C(new_new_n102_), .Y(new_new_n105_));
  NA2        g083(.A(i_12_), .B(i_7_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n57_), .B(new_new_n26_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n107_), .B(i_0_), .Y(new_new_n108_));
  NA2        g086(.A(i_11_), .B(i_12_), .Y(new_new_n109_));
  OAI210     g087(.A0(new_new_n108_), .A1(new_new_n106_), .B0(new_new_n109_), .Y(new_new_n110_));
  NO2        g088(.A(new_new_n110_), .B(new_new_n105_), .Y(new_new_n111_));
  NAi41      g089(.An(new_new_n100_), .B(new_new_n111_), .C(new_new_n98_), .D(new_new_n91_), .Y(new_new_n112_));
  NOi21      g090(.An(i_1_), .B(i_5_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n113_), .B(i_11_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n92_), .B(new_new_n37_), .Y(new_new_n115_));
  NA2        g093(.A(i_7_), .B(new_new_n25_), .Y(new_new_n116_));
  NA2        g094(.A(new_new_n116_), .B(new_new_n115_), .Y(new_new_n117_));
  NO2        g095(.A(new_new_n117_), .B(new_new_n46_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n82_), .B(new_new_n81_), .Y(new_new_n119_));
  NAi21      g097(.An(i_3_), .B(i_8_), .Y(new_new_n120_));
  INV        g098(.A(new_new_n120_), .Y(new_new_n121_));
  NOi21      g099(.An(new_new_n121_), .B(new_new_n119_), .Y(new_new_n122_));
  NO2        g100(.A(i_1_), .B(new_new_n77_), .Y(new_new_n123_));
  NO2        g101(.A(i_6_), .B(i_5_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(i_3_), .Y(new_new_n125_));
  AO210      g103(.A0(new_new_n125_), .A1(new_new_n47_), .B0(new_new_n123_), .Y(new_new_n126_));
  OAI220     g104(.A0(new_new_n126_), .A1(new_new_n99_), .B0(new_new_n122_), .B1(new_new_n114_), .Y(new_new_n127_));
  NO3        g105(.A(new_new_n127_), .B(new_new_n112_), .C(new_new_n86_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n71_), .Y(mai2));
  NO2        g107(.A(new_new_n57_), .B(new_new_n37_), .Y(new_new_n130_));
  NA2        g108(.A(i_6_), .B(new_new_n25_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(new_new_n130_), .Y(new_new_n132_));
  NA4        g110(.A(new_new_n132_), .B(new_new_n69_), .C(new_new_n61_), .D(new_new_n30_), .Y(mai0));
  AN2        g111(.A(i_8_), .B(i_7_), .Y(new_new_n134_));
  NA2        g112(.A(new_new_n134_), .B(i_6_), .Y(new_new_n135_));
  NO2        g113(.A(i_12_), .B(i_13_), .Y(new_new_n136_));
  NAi21      g114(.An(i_5_), .B(i_11_), .Y(new_new_n137_));
  NOi21      g115(.An(new_new_n136_), .B(new_new_n137_), .Y(new_new_n138_));
  NO2        g116(.A(i_0_), .B(i_1_), .Y(new_new_n139_));
  NA2        g117(.A(i_2_), .B(i_3_), .Y(new_new_n140_));
  NO2        g118(.A(new_new_n140_), .B(i_4_), .Y(new_new_n141_));
  NA2        g119(.A(new_new_n141_), .B(new_new_n138_), .Y(new_new_n142_));
  AN2        g120(.A(new_new_n136_), .B(new_new_n75_), .Y(new_new_n143_));
  NA2        g121(.A(i_1_), .B(i_5_), .Y(new_new_n144_));
  NA2        g122(.A(i_0_), .B(new_new_n36_), .Y(new_new_n145_));
  NO3        g123(.A(new_new_n145_), .B(new_new_n144_), .C(i_13_), .Y(new_new_n146_));
  OR2        g124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NO3        g125(.A(new_new_n147_), .B(new_new_n72_), .C(i_13_), .Y(new_new_n148_));
  NAi32      g126(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n149_));
  NAi21      g127(.An(new_new_n149_), .B(new_new_n148_), .Y(new_new_n150_));
  NOi21      g128(.An(i_4_), .B(i_10_), .Y(new_new_n151_));
  NA2        g129(.A(new_new_n151_), .B(new_new_n40_), .Y(new_new_n152_));
  NO2        g130(.A(i_3_), .B(i_5_), .Y(new_new_n153_));
  NO3        g131(.A(new_new_n65_), .B(i_2_), .C(i_1_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n154_), .B(new_new_n153_), .Y(new_new_n155_));
  OAI210     g133(.A0(new_new_n155_), .A1(new_new_n152_), .B0(new_new_n150_), .Y(new_new_n156_));
  NO2        g134(.A(new_new_n156_), .B(new_new_n146_), .Y(new_new_n157_));
  AOI210     g135(.A0(new_new_n157_), .A1(new_new_n142_), .B0(new_new_n135_), .Y(new_new_n158_));
  NA3        g136(.A(new_new_n65_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n159_));
  NA2        g137(.A(i_3_), .B(new_new_n48_), .Y(new_new_n160_));
  NOi21      g138(.An(i_4_), .B(i_9_), .Y(new_new_n161_));
  NOi21      g139(.An(i_11_), .B(i_13_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  OR2        g141(.A(new_new_n163_), .B(new_new_n160_), .Y(new_new_n164_));
  NO2        g142(.A(i_4_), .B(i_5_), .Y(new_new_n165_));
  NAi21      g143(.An(i_12_), .B(i_11_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n166_), .B(i_13_), .Y(new_new_n167_));
  NA3        g145(.A(new_new_n167_), .B(new_new_n165_), .C(new_new_n75_), .Y(new_new_n168_));
  AOI210     g146(.A0(new_new_n168_), .A1(new_new_n164_), .B0(new_new_n159_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n65_), .B(new_new_n57_), .Y(new_new_n170_));
  NA2        g148(.A(new_new_n170_), .B(new_new_n46_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n36_), .B(i_5_), .Y(new_new_n172_));
  NAi31      g150(.An(new_new_n172_), .B(new_new_n143_), .C(i_11_), .Y(new_new_n173_));
  NA2        g151(.A(i_3_), .B(i_5_), .Y(new_new_n174_));
  OR2        g152(.A(new_new_n174_), .B(new_new_n163_), .Y(new_new_n175_));
  AOI210     g153(.A0(new_new_n175_), .A1(new_new_n173_), .B0(new_new_n171_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n65_), .B(i_5_), .Y(new_new_n177_));
  NO2        g155(.A(i_13_), .B(i_10_), .Y(new_new_n178_));
  NA3        g156(.A(new_new_n178_), .B(new_new_n177_), .C(new_new_n44_), .Y(new_new_n179_));
  NO2        g157(.A(i_2_), .B(i_1_), .Y(new_new_n180_));
  NAi21      g158(.An(i_4_), .B(i_12_), .Y(new_new_n181_));
  NO3        g159(.A(new_new_n181_), .B(new_new_n944_), .C(new_new_n179_), .Y(new_new_n182_));
  NO3        g160(.A(new_new_n182_), .B(new_new_n176_), .C(new_new_n169_), .Y(new_new_n183_));
  INV        g161(.A(i_8_), .Y(new_new_n184_));
  INV        g162(.A(i_6_), .Y(new_new_n185_));
  NO3        g163(.A(i_3_), .B(new_new_n77_), .C(new_new_n48_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n186_), .B(new_new_n104_), .Y(new_new_n187_));
  NO3        g165(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n188_));
  NA3        g166(.A(new_new_n188_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n189_));
  NO3        g167(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n190_));
  NO2        g168(.A(i_13_), .B(new_new_n187_), .Y(new_new_n191_));
  NO2        g169(.A(i_3_), .B(i_8_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n40_), .Y(new_new_n194_));
  NO2        g172(.A(i_13_), .B(i_9_), .Y(new_new_n195_));
  NAi21      g173(.An(i_12_), .B(i_3_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n44_), .B(i_5_), .Y(new_new_n197_));
  NO3        g175(.A(i_0_), .B(i_2_), .C(new_new_n57_), .Y(new_new_n198_));
  NA3        g176(.A(new_new_n198_), .B(new_new_n197_), .C(i_10_), .Y(new_new_n199_));
  OAI220     g177(.A0(new_new_n199_), .A1(i_13_), .B0(new_new_n53_), .B1(new_new_n194_), .Y(new_new_n200_));
  AOI210     g178(.A0(new_new_n200_), .A1(i_7_), .B0(new_new_n191_), .Y(new_new_n201_));
  OAI220     g179(.A0(new_new_n201_), .A1(i_4_), .B0(new_new_n185_), .B1(new_new_n183_), .Y(new_new_n202_));
  NA3        g180(.A(i_13_), .B(new_new_n184_), .C(i_10_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n203_), .B(i_12_), .Y(new_new_n204_));
  NA2        g182(.A(i_0_), .B(i_5_), .Y(new_new_n205_));
  NAi31      g183(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n36_), .B(i_13_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n46_), .B(new_new_n57_), .Y(new_new_n208_));
  NA3        g186(.A(new_new_n208_), .B(i_3_), .C(new_new_n207_), .Y(new_new_n209_));
  INV        g187(.A(i_13_), .Y(new_new_n210_));
  NO2        g188(.A(i_12_), .B(new_new_n210_), .Y(new_new_n211_));
  NA3        g189(.A(new_new_n211_), .B(new_new_n188_), .C(new_new_n186_), .Y(new_new_n212_));
  OAI210     g190(.A0(new_new_n209_), .A1(new_new_n206_), .B0(new_new_n212_), .Y(new_new_n213_));
  AOI220     g191(.A0(new_new_n213_), .A1(new_new_n134_), .B0(i_3_), .B1(new_new_n204_), .Y(new_new_n214_));
  NO2        g192(.A(i_12_), .B(new_new_n37_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n174_), .B(i_4_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  OR2        g195(.A(i_8_), .B(i_7_), .Y(new_new_n218_));
  NO2        g196(.A(new_new_n218_), .B(new_new_n77_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n51_), .B(i_1_), .Y(new_new_n220_));
  INV        g198(.A(i_12_), .Y(new_new_n221_));
  NO3        g199(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n222_));
  NA2        g200(.A(i_2_), .B(i_1_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n51_), .B(new_new_n217_), .Y(new_new_n224_));
  NO3        g202(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n225_));
  NAi21      g203(.An(i_4_), .B(i_3_), .Y(new_new_n226_));
  NO2        g204(.A(i_0_), .B(i_6_), .Y(new_new_n227_));
  NOi41      g205(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n228_));
  NA2        g206(.A(new_new_n228_), .B(new_new_n227_), .Y(new_new_n229_));
  AOI210     g207(.A0(new_new_n940_), .A1(new_new_n40_), .B0(new_new_n224_), .Y(new_new_n230_));
  NO2        g208(.A(i_11_), .B(new_new_n210_), .Y(new_new_n231_));
  NOi21      g209(.An(i_1_), .B(i_6_), .Y(new_new_n232_));
  NAi21      g210(.An(i_3_), .B(i_7_), .Y(new_new_n233_));
  NO2        g211(.A(i_12_), .B(i_3_), .Y(new_new_n234_));
  NA3        g212(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n135_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n221_), .B(i_13_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n67_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n236_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n218_), .B(new_new_n37_), .Y(new_new_n240_));
  NA2        g218(.A(i_12_), .B(i_6_), .Y(new_new_n241_));
  OR2        g219(.A(i_13_), .B(i_9_), .Y(new_new_n242_));
  NO3        g220(.A(new_new_n242_), .B(new_new_n241_), .C(new_new_n48_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n226_), .B(i_2_), .Y(new_new_n244_));
  NA3        g222(.A(new_new_n244_), .B(new_new_n243_), .C(new_new_n44_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n231_), .B(i_9_), .Y(new_new_n246_));
  OAI210     g224(.A0(new_new_n57_), .A1(new_new_n246_), .B0(new_new_n245_), .Y(new_new_n247_));
  NO3        g225(.A(i_11_), .B(new_new_n210_), .C(new_new_n25_), .Y(new_new_n248_));
  NO2        g226(.A(new_new_n233_), .B(i_8_), .Y(new_new_n249_));
  NO2        g227(.A(i_6_), .B(new_new_n48_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n247_), .B(new_new_n240_), .Y(new_new_n251_));
  NA4        g229(.A(new_new_n251_), .B(new_new_n239_), .C(new_new_n230_), .D(new_new_n214_), .Y(new_new_n252_));
  NO3        g230(.A(i_12_), .B(new_new_n210_), .C(new_new_n37_), .Y(new_new_n253_));
  INV        g231(.A(new_new_n253_), .Y(new_new_n254_));
  NA2        g232(.A(i_8_), .B(new_new_n92_), .Y(new_new_n255_));
  NO3        g233(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n256_));
  NO2        g234(.A(new_new_n223_), .B(i_0_), .Y(new_new_n257_));
  NA2        g235(.A(new_new_n250_), .B(new_new_n26_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n258_), .B(new_new_n941_), .Y(new_new_n259_));
  NA2        g237(.A(i_0_), .B(i_1_), .Y(new_new_n260_));
  NO2        g238(.A(new_new_n260_), .B(i_2_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n54_), .B(i_6_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n262_), .B(new_new_n261_), .Y(new_new_n263_));
  OAI210     g241(.A0(new_new_n155_), .A1(new_new_n135_), .B0(new_new_n263_), .Y(new_new_n264_));
  NO2        g242(.A(new_new_n264_), .B(new_new_n259_), .Y(new_new_n265_));
  NO2        g243(.A(i_3_), .B(i_10_), .Y(new_new_n266_));
  NA3        g244(.A(new_new_n266_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n267_));
  NO2        g245(.A(i_2_), .B(new_new_n92_), .Y(new_new_n268_));
  NA2        g246(.A(i_1_), .B(new_new_n36_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n269_), .B(i_8_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n270_), .B(new_new_n268_), .Y(new_new_n271_));
  AN2        g249(.A(i_3_), .B(i_10_), .Y(new_new_n272_));
  NA3        g250(.A(new_new_n272_), .B(new_new_n167_), .C(new_new_n165_), .Y(new_new_n273_));
  NO2        g251(.A(i_5_), .B(new_new_n37_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n275_));
  OR2        g253(.A(new_new_n271_), .B(new_new_n267_), .Y(new_new_n276_));
  OAI220     g254(.A0(new_new_n276_), .A1(i_6_), .B0(new_new_n265_), .B1(new_new_n254_), .Y(new_new_n277_));
  NO4        g255(.A(new_new_n277_), .B(new_new_n252_), .C(new_new_n202_), .D(new_new_n158_), .Y(new_new_n278_));
  NO3        g256(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n279_));
  NO3        g257(.A(i_6_), .B(new_new_n184_), .C(i_7_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n280_), .B(new_new_n188_), .Y(new_new_n281_));
  AOI210     g259(.A0(new_new_n281_), .A1(new_new_n223_), .B0(new_new_n160_), .Y(new_new_n282_));
  NO2        g260(.A(i_2_), .B(i_3_), .Y(new_new_n283_));
  OR2        g261(.A(i_0_), .B(i_5_), .Y(new_new_n284_));
  NA3        g262(.A(new_new_n219_), .B(new_new_n283_), .C(i_1_), .Y(new_new_n285_));
  NA2        g263(.A(new_new_n257_), .B(new_new_n104_), .Y(new_new_n286_));
  NAi21      g264(.An(i_8_), .B(i_7_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(i_6_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n147_), .B(new_new_n46_), .Y(new_new_n289_));
  NA2        g267(.A(new_new_n289_), .B(new_new_n288_), .Y(new_new_n290_));
  NA3        g268(.A(new_new_n290_), .B(new_new_n286_), .C(new_new_n285_), .Y(new_new_n291_));
  OAI210     g269(.A0(new_new_n291_), .A1(new_new_n282_), .B0(i_4_), .Y(new_new_n292_));
  NO2        g270(.A(i_12_), .B(i_10_), .Y(new_new_n293_));
  NOi21      g271(.An(i_5_), .B(i_0_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n269_), .B(new_new_n120_), .Y(new_new_n295_));
  NA4        g273(.A(new_new_n76_), .B(new_new_n36_), .C(new_new_n77_), .D(i_8_), .Y(new_new_n296_));
  NA2        g274(.A(new_new_n295_), .B(new_new_n293_), .Y(new_new_n297_));
  NO2        g275(.A(i_6_), .B(i_8_), .Y(new_new_n298_));
  NOi21      g276(.An(i_0_), .B(i_2_), .Y(new_new_n299_));
  AN2        g277(.A(new_new_n299_), .B(new_new_n298_), .Y(new_new_n300_));
  NO2        g278(.A(i_1_), .B(i_7_), .Y(new_new_n301_));
  AO220      g279(.A0(new_new_n301_), .A1(new_new_n300_), .B0(new_new_n288_), .B1(new_new_n220_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n302_), .B(i_4_), .Y(new_new_n303_));
  NA3        g281(.A(new_new_n303_), .B(new_new_n297_), .C(new_new_n292_), .Y(new_new_n304_));
  NO3        g282(.A(new_new_n218_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n305_));
  NO3        g283(.A(new_new_n287_), .B(i_2_), .C(i_1_), .Y(new_new_n306_));
  OAI210     g284(.A0(new_new_n306_), .A1(new_new_n305_), .B0(i_6_), .Y(new_new_n307_));
  NA2        g285(.A(new_new_n268_), .B(new_new_n184_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n308_), .B(new_new_n307_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n309_), .B(i_3_), .Y(new_new_n310_));
  INV        g288(.A(new_new_n76_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n84_), .B(new_new_n184_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n73_), .B(new_new_n311_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n184_), .B(i_9_), .Y(new_new_n314_));
  NA2        g292(.A(new_new_n314_), .B(i_0_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n313_), .B(new_new_n259_), .Y(new_new_n316_));
  AOI210     g294(.A0(new_new_n316_), .A1(new_new_n310_), .B0(new_new_n152_), .Y(new_new_n317_));
  AOI210     g295(.A0(new_new_n304_), .A1(new_new_n279_), .B0(new_new_n317_), .Y(new_new_n318_));
  NOi32      g296(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n319_));
  INV        g297(.A(new_new_n319_), .Y(new_new_n320_));
  NAi21      g298(.An(i_0_), .B(i_6_), .Y(new_new_n321_));
  NAi21      g299(.An(i_1_), .B(i_5_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n322_), .B(new_new_n321_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n323_), .B(new_new_n25_), .Y(new_new_n324_));
  OAI210     g302(.A0(new_new_n324_), .A1(new_new_n149_), .B0(new_new_n229_), .Y(new_new_n325_));
  NAi41      g303(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n326_));
  OAI220     g304(.A0(new_new_n326_), .A1(new_new_n322_), .B0(new_new_n206_), .B1(new_new_n149_), .Y(new_new_n327_));
  AOI210     g305(.A0(new_new_n326_), .A1(new_new_n149_), .B0(new_new_n147_), .Y(new_new_n328_));
  NOi32      g306(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n329_));
  NAi21      g307(.An(i_6_), .B(i_1_), .Y(new_new_n330_));
  NA3        g308(.A(new_new_n330_), .B(new_new_n329_), .C(new_new_n46_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n331_), .B(i_0_), .Y(new_new_n332_));
  OR3        g310(.A(new_new_n332_), .B(new_new_n328_), .C(new_new_n327_), .Y(new_new_n333_));
  NO2        g311(.A(i_1_), .B(new_new_n92_), .Y(new_new_n334_));
  NAi21      g312(.An(i_3_), .B(i_4_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n335_), .B(i_9_), .Y(new_new_n336_));
  AN2        g314(.A(i_6_), .B(i_7_), .Y(new_new_n337_));
  NA2        g315(.A(i_2_), .B(i_7_), .Y(new_new_n338_));
  NO2        g316(.A(new_new_n335_), .B(i_10_), .Y(new_new_n339_));
  NA3        g317(.A(new_new_n339_), .B(new_new_n338_), .C(new_new_n227_), .Y(new_new_n340_));
  INV        g318(.A(new_new_n340_), .Y(new_new_n341_));
  AOI210     g319(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n342_));
  OAI210     g320(.A0(new_new_n342_), .A1(new_new_n180_), .B0(new_new_n339_), .Y(new_new_n343_));
  AOI220     g321(.A0(new_new_n339_), .A1(new_new_n301_), .B0(new_new_n222_), .B1(new_new_n180_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(i_5_), .Y(new_new_n345_));
  NO4        g323(.A(new_new_n345_), .B(new_new_n341_), .C(new_new_n333_), .D(new_new_n325_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n346_), .B(new_new_n320_), .Y(new_new_n347_));
  NO2        g325(.A(new_new_n54_), .B(new_new_n25_), .Y(new_new_n348_));
  AN2        g326(.A(i_12_), .B(i_5_), .Y(new_new_n349_));
  NO2        g327(.A(i_4_), .B(new_new_n26_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n350_), .B(new_new_n349_), .Y(new_new_n351_));
  NO2        g329(.A(i_11_), .B(i_6_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n352_), .B(new_new_n289_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n353_), .B(new_new_n351_), .Y(new_new_n354_));
  NO2        g332(.A(new_new_n226_), .B(i_5_), .Y(new_new_n355_));
  NO2        g333(.A(i_5_), .B(i_10_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n136_), .B(new_new_n45_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(new_new_n226_), .Y(new_new_n358_));
  OAI210     g336(.A0(new_new_n358_), .A1(new_new_n354_), .B0(new_new_n348_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n360_));
  NA2        g338(.A(new_new_n354_), .B(new_new_n360_), .Y(new_new_n361_));
  NO3        g339(.A(new_new_n77_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n362_));
  NO2        g340(.A(i_11_), .B(i_12_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n356_), .B(new_new_n221_), .Y(new_new_n364_));
  NA2        g342(.A(new_new_n104_), .B(i_4_), .Y(new_new_n365_));
  OAI220     g343(.A0(new_new_n365_), .A1(new_new_n206_), .B0(new_new_n364_), .B1(new_new_n296_), .Y(new_new_n366_));
  NAi21      g344(.An(i_13_), .B(i_0_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n367_), .B(new_new_n223_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n366_), .B(new_new_n368_), .Y(new_new_n369_));
  NA3        g347(.A(new_new_n369_), .B(new_new_n361_), .C(new_new_n359_), .Y(new_new_n370_));
  NO2        g348(.A(i_0_), .B(i_11_), .Y(new_new_n371_));
  AN2        g349(.A(i_1_), .B(i_6_), .Y(new_new_n372_));
  NOi21      g350(.An(i_2_), .B(i_12_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n373_), .B(new_new_n372_), .Y(new_new_n374_));
  INV        g352(.A(new_new_n374_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n134_), .B(i_9_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(i_4_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n375_), .B(new_new_n377_), .Y(new_new_n378_));
  OR2        g356(.A(i_13_), .B(i_10_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n163_), .B(new_new_n115_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n92_), .B(new_new_n25_), .Y(new_new_n381_));
  INV        g359(.A(new_new_n285_), .Y(new_new_n382_));
  AOI220     g360(.A0(new_new_n262_), .A1(new_new_n256_), .B0(new_new_n257_), .B1(i_8_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n160_), .Y(new_new_n384_));
  NO2        g362(.A(i_2_), .B(new_new_n255_), .Y(new_new_n385_));
  NO3        g363(.A(new_new_n385_), .B(new_new_n384_), .C(new_new_n382_), .Y(new_new_n386_));
  NO2        g364(.A(i_3_), .B(new_new_n287_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n262_), .B(new_new_n220_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n388_), .B(new_new_n174_), .Y(new_new_n389_));
  NA3        g367(.A(new_new_n301_), .B(new_new_n300_), .C(i_5_), .Y(new_new_n390_));
  INV        g368(.A(new_new_n390_), .Y(new_new_n391_));
  NO3        g369(.A(new_new_n391_), .B(new_new_n389_), .C(new_new_n387_), .Y(new_new_n392_));
  AOI210     g370(.A0(new_new_n392_), .A1(new_new_n386_), .B0(new_new_n246_), .Y(new_new_n393_));
  NO4        g371(.A(new_new_n393_), .B(new_new_n943_), .C(new_new_n370_), .D(new_new_n347_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n57_), .B(i_4_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n65_), .B(i_13_), .Y(new_new_n396_));
  NA3        g374(.A(new_new_n396_), .B(new_new_n395_), .C(i_2_), .Y(new_new_n397_));
  NO2        g375(.A(i_10_), .B(i_9_), .Y(new_new_n398_));
  NAi21      g376(.An(i_12_), .B(i_8_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n399_), .B(i_3_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n400_), .B(new_new_n398_), .Y(new_new_n401_));
  NA2        g379(.A(i_2_), .B(new_new_n95_), .Y(new_new_n402_));
  OAI220     g380(.A0(new_new_n402_), .A1(new_new_n194_), .B0(new_new_n401_), .B1(new_new_n397_), .Y(new_new_n403_));
  NA2        g381(.A(new_new_n275_), .B(i_0_), .Y(new_new_n404_));
  NO3        g382(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n241_), .B(new_new_n88_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n406_), .B(new_new_n405_), .Y(new_new_n407_));
  NA2        g385(.A(i_8_), .B(i_9_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n407_), .B(new_new_n404_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n231_), .B(new_new_n274_), .Y(new_new_n410_));
  NO3        g388(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n411_));
  INV        g389(.A(new_new_n411_), .Y(new_new_n412_));
  NA3        g390(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n413_));
  NA4        g391(.A(new_new_n137_), .B(new_new_n107_), .C(new_new_n72_), .D(new_new_n23_), .Y(new_new_n414_));
  OAI220     g392(.A0(new_new_n414_), .A1(new_new_n413_), .B0(new_new_n412_), .B1(new_new_n410_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n409_), .C(new_new_n403_), .Y(new_new_n416_));
  OR2        g394(.A(new_new_n260_), .B(i_13_), .Y(new_new_n417_));
  OA210      g395(.A0(new_new_n315_), .A1(new_new_n92_), .B0(new_new_n263_), .Y(new_new_n418_));
  OA220      g396(.A0(new_new_n418_), .A1(new_new_n152_), .B0(new_new_n417_), .B1(new_new_n217_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n87_), .B(i_13_), .Y(new_new_n420_));
  NA2        g398(.A(i_3_), .B(new_new_n348_), .Y(new_new_n421_));
  NO2        g399(.A(i_2_), .B(i_13_), .Y(new_new_n422_));
  NA3        g400(.A(new_new_n422_), .B(new_new_n151_), .C(new_new_n90_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n421_), .B(new_new_n420_), .Y(new_new_n424_));
  NO3        g402(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n425_));
  NO2        g403(.A(i_6_), .B(i_7_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n426_), .B(new_new_n425_), .Y(new_new_n427_));
  NO2        g405(.A(i_11_), .B(i_1_), .Y(new_new_n428_));
  OR2        g406(.A(i_11_), .B(i_8_), .Y(new_new_n429_));
  NOi21      g407(.An(i_2_), .B(i_7_), .Y(new_new_n430_));
  NAi31      g408(.An(new_new_n429_), .B(new_new_n430_), .C(i_0_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n945_), .B(new_new_n395_), .Y(new_new_n432_));
  NO2        g410(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n433_));
  NO2        g411(.A(i_3_), .B(new_new_n184_), .Y(new_new_n434_));
  NO2        g412(.A(i_6_), .B(i_10_), .Y(new_new_n435_));
  NA3        g413(.A(new_new_n435_), .B(new_new_n279_), .C(new_new_n434_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n436_), .B(new_new_n145_), .Y(new_new_n437_));
  NO2        g415(.A(new_new_n147_), .B(i_3_), .Y(new_new_n438_));
  NA3        g416(.A(new_new_n360_), .B(new_new_n170_), .C(new_new_n141_), .Y(new_new_n439_));
  INV        g417(.A(new_new_n439_), .Y(new_new_n440_));
  NO4        g418(.A(new_new_n440_), .B(new_new_n437_), .C(new_new_n433_), .D(new_new_n424_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n411_), .B(new_new_n356_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n442_), .B(new_new_n209_), .Y(new_new_n443_));
  NAi21      g421(.An(new_new_n203_), .B(new_new_n363_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n26_), .B(i_5_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n942_), .B(new_new_n445_), .C(new_new_n134_), .Y(new_new_n446_));
  OR3        g424(.A(new_new_n269_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n447_), .B(new_new_n446_), .Y(new_new_n448_));
  NA3        g426(.A(new_new_n272_), .B(new_new_n208_), .C(new_new_n65_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n449_), .B(new_new_n427_), .Y(new_new_n450_));
  NO3        g428(.A(new_new_n450_), .B(new_new_n448_), .C(new_new_n443_), .Y(new_new_n451_));
  NA4        g429(.A(new_new_n451_), .B(new_new_n441_), .C(new_new_n419_), .D(new_new_n416_), .Y(new_new_n452_));
  NA3        g430(.A(new_new_n272_), .B(new_new_n167_), .C(new_new_n165_), .Y(new_new_n453_));
  INV        g431(.A(new_new_n453_), .Y(new_new_n454_));
  BUFFER     g432(.A(new_new_n256_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  AN2        g434(.A(i_12_), .B(new_new_n405_), .Y(new_new_n457_));
  OAI210     g435(.A0(new_new_n65_), .A1(new_new_n217_), .B0(new_new_n273_), .Y(new_new_n458_));
  AOI220     g436(.A0(new_new_n458_), .A1(new_new_n288_), .B0(new_new_n457_), .B1(new_new_n275_), .Y(new_new_n459_));
  NA4        g437(.A(new_new_n396_), .B(new_new_n395_), .C(new_new_n192_), .D(i_2_), .Y(new_new_n460_));
  INV        g438(.A(new_new_n460_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n319_), .B(new_new_n65_), .Y(new_new_n462_));
  INV        g440(.A(new_new_n329_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n36_), .B(i_8_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n39_), .B(i_13_), .Y(new_new_n465_));
  INV        g443(.A(new_new_n465_), .Y(new_new_n466_));
  AOI210     g444(.A0(new_new_n461_), .A1(new_new_n193_), .B0(new_new_n466_), .Y(new_new_n467_));
  OAI210     g445(.A0(i_8_), .A1(new_new_n57_), .B0(new_new_n126_), .Y(new_new_n468_));
  NO2        g446(.A(i_7_), .B(new_new_n189_), .Y(new_new_n469_));
  OR2        g447(.A(new_new_n174_), .B(i_4_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n77_), .Y(new_new_n471_));
  AOI220     g449(.A0(new_new_n471_), .A1(new_new_n469_), .B0(new_new_n468_), .B1(new_new_n380_), .Y(new_new_n472_));
  NA4        g450(.A(new_new_n472_), .B(new_new_n467_), .C(new_new_n459_), .D(new_new_n456_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n355_), .B(new_new_n261_), .Y(new_new_n474_));
  OAI210     g452(.A0(new_new_n351_), .A1(new_new_n159_), .B0(new_new_n474_), .Y(new_new_n475_));
  NO2        g453(.A(i_12_), .B(new_new_n184_), .Y(new_new_n476_));
  NA2        g454(.A(new_new_n476_), .B(new_new_n210_), .Y(new_new_n477_));
  NO2        g455(.A(i_6_), .B(new_new_n477_), .Y(new_new_n478_));
  NOi21      g456(.An(new_new_n280_), .B(new_new_n38_), .Y(new_new_n479_));
  OAI210     g457(.A0(new_new_n479_), .A1(new_new_n478_), .B0(new_new_n475_), .Y(new_new_n480_));
  NO2        g458(.A(i_8_), .B(i_7_), .Y(new_new_n481_));
  INV        g459(.A(new_new_n208_), .Y(new_new_n482_));
  OAI220     g460(.A0(new_new_n46_), .A1(new_new_n470_), .B0(new_new_n482_), .B1(new_new_n226_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n44_), .B(i_10_), .Y(new_new_n484_));
  NO2        g462(.A(new_new_n484_), .B(i_6_), .Y(new_new_n485_));
  NA3        g463(.A(new_new_n485_), .B(new_new_n483_), .C(new_new_n481_), .Y(new_new_n486_));
  NO2        g464(.A(new_new_n420_), .B(new_new_n125_), .Y(new_new_n487_));
  NA2        g465(.A(new_new_n487_), .B(new_new_n240_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n267_), .B(new_new_n172_), .Y(new_new_n489_));
  NA3        g467(.A(new_new_n272_), .B(new_new_n165_), .C(new_new_n87_), .Y(new_new_n490_));
  NO2        g468(.A(new_new_n207_), .B(new_new_n44_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n147_), .B(i_5_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n492_), .B(new_new_n283_), .Y(new_new_n493_));
  OAI210     g471(.A0(new_new_n493_), .A1(new_new_n491_), .B0(new_new_n490_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n494_), .A1(new_new_n489_), .B0(new_new_n411_), .Y(new_new_n495_));
  NA4        g473(.A(new_new_n495_), .B(new_new_n488_), .C(new_new_n486_), .D(new_new_n480_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n253_), .B(new_new_n76_), .Y(new_new_n497_));
  NO2        g475(.A(new_new_n73_), .B(new_new_n497_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n256_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n499_), .B(new_new_n164_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n208_), .B(i_3_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n398_), .B(new_new_n207_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n501_), .B(new_new_n502_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n476_), .B(new_new_n248_), .Y(new_new_n504_));
  NO2        g482(.A(new_new_n92_), .B(new_new_n504_), .Y(new_new_n505_));
  NO4        g483(.A(new_new_n505_), .B(new_new_n503_), .C(new_new_n500_), .D(new_new_n498_), .Y(new_new_n506_));
  NO4        g484(.A(new_new_n232_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n507_));
  NO3        g485(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n218_), .B(new_new_n36_), .Y(new_new_n509_));
  AN2        g487(.A(new_new_n509_), .B(new_new_n508_), .Y(new_new_n510_));
  OA210      g488(.A0(new_new_n510_), .A1(new_new_n507_), .B0(new_new_n319_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n379_), .B(i_1_), .Y(new_new_n512_));
  NOi31      g490(.An(new_new_n512_), .B(new_new_n406_), .C(new_new_n65_), .Y(new_new_n513_));
  AN3        g491(.A(new_new_n513_), .B(new_new_n377_), .C(new_new_n445_), .Y(new_new_n514_));
  NO2        g492(.A(new_new_n383_), .B(new_new_n168_), .Y(new_new_n515_));
  NO3        g493(.A(new_new_n515_), .B(new_new_n514_), .C(new_new_n511_), .Y(new_new_n516_));
  NOi21      g494(.An(i_10_), .B(i_6_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n77_), .B(new_new_n25_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n248_), .B(new_new_n517_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n519_), .B(new_new_n404_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n106_), .B(new_new_n23_), .Y(new_new_n521_));
  INV        g499(.A(new_new_n280_), .Y(new_new_n522_));
  AOI220     g500(.A0(new_new_n522_), .A1(new_new_n388_), .B0(new_new_n175_), .B1(new_new_n173_), .Y(new_new_n523_));
  NOi21      g501(.An(new_new_n138_), .B(new_new_n296_), .Y(new_new_n524_));
  NO3        g502(.A(new_new_n524_), .B(new_new_n523_), .C(new_new_n520_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n462_), .B(new_new_n344_), .Y(new_new_n526_));
  INV        g504(.A(new_new_n283_), .Y(new_new_n527_));
  NO2        g505(.A(i_12_), .B(new_new_n77_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n528_), .B(new_new_n248_), .Y(new_new_n529_));
  NA2        g507(.A(new_new_n352_), .B(new_new_n253_), .Y(new_new_n530_));
  AOI210     g508(.A0(new_new_n530_), .A1(new_new_n529_), .B0(new_new_n527_), .Y(new_new_n531_));
  NO3        g509(.A(i_4_), .B(new_new_n307_), .C(new_new_n267_), .Y(new_new_n532_));
  NO2        g510(.A(i_2_), .B(new_new_n444_), .Y(new_new_n533_));
  NO4        g511(.A(new_new_n533_), .B(new_new_n532_), .C(new_new_n531_), .D(new_new_n526_), .Y(new_new_n534_));
  NA4        g512(.A(new_new_n534_), .B(new_new_n525_), .C(new_new_n516_), .D(new_new_n506_), .Y(new_new_n535_));
  NO4        g513(.A(new_new_n535_), .B(new_new_n496_), .C(new_new_n473_), .D(new_new_n452_), .Y(new_new_n536_));
  NA4        g514(.A(new_new_n536_), .B(new_new_n394_), .C(new_new_n318_), .D(new_new_n278_), .Y(mai7));
  NA2        g515(.A(new_new_n435_), .B(new_new_n76_), .Y(new_new_n538_));
  NA2        g516(.A(new_new_n136_), .B(i_8_), .Y(new_new_n539_));
  NO2        g517(.A(new_new_n539_), .B(new_new_n538_), .Y(new_new_n540_));
  NA3        g518(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n221_), .B(i_4_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n542_), .B(i_8_), .Y(new_new_n543_));
  NA2        g521(.A(i_2_), .B(new_new_n77_), .Y(new_new_n544_));
  OAI210     g522(.A0(new_new_n80_), .A1(new_new_n192_), .B0(new_new_n193_), .Y(new_new_n545_));
  NA2        g523(.A(i_4_), .B(i_8_), .Y(new_new_n546_));
  OAI220     g524(.A0(new_new_n37_), .A1(new_new_n544_), .B0(new_new_n545_), .B1(i_13_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n547_), .B(new_new_n540_), .Y(new_new_n548_));
  OR2        g526(.A(i_6_), .B(i_10_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n549_), .B(new_new_n23_), .Y(new_new_n550_));
  OR3        g528(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n551_));
  NO3        g529(.A(new_new_n551_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n552_));
  INV        g530(.A(new_new_n190_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n552_), .B(new_new_n550_), .Y(new_new_n554_));
  OR2        g532(.A(new_new_n554_), .B(new_new_n527_), .Y(new_new_n555_));
  AOI210     g533(.A0(new_new_n555_), .A1(new_new_n548_), .B0(new_new_n57_), .Y(new_new_n556_));
  NOi21      g534(.An(i_11_), .B(i_7_), .Y(new_new_n557_));
  AO210      g535(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n558_), .B(new_new_n557_), .Y(new_new_n559_));
  NA3        g537(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n560_));
  NAi31      g538(.An(new_new_n560_), .B(i_12_), .C(i_11_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n561_), .B(new_new_n57_), .Y(new_new_n562_));
  NA2        g540(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n563_));
  AO210      g541(.A0(new_new_n563_), .A1(new_new_n344_), .B0(new_new_n41_), .Y(new_new_n564_));
  NA2        g542(.A(new_new_n211_), .B(new_new_n57_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n373_), .B(new_new_n31_), .Y(new_new_n566_));
  OR2        g544(.A(new_new_n196_), .B(new_new_n99_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n567_), .B(new_new_n566_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n57_), .B(i_9_), .Y(new_new_n569_));
  NA2        g547(.A(new_new_n57_), .B(new_new_n568_), .Y(new_new_n570_));
  NO2        g548(.A(i_1_), .B(i_12_), .Y(new_new_n571_));
  NA3        g549(.A(new_new_n570_), .B(new_new_n565_), .C(new_new_n564_), .Y(new_new_n572_));
  OAI210     g550(.A0(new_new_n572_), .A1(new_new_n562_), .B0(i_6_), .Y(new_new_n573_));
  NO2        g551(.A(i_6_), .B(i_11_), .Y(new_new_n574_));
  INV        g552(.A(new_new_n407_), .Y(new_new_n575_));
  NO4        g553(.A(i_12_), .B(new_new_n120_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n576_));
  NA2        g554(.A(new_new_n576_), .B(new_new_n569_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n221_), .B(i_6_), .Y(new_new_n578_));
  INV        g556(.A(new_new_n577_), .Y(new_new_n579_));
  NA3        g557(.A(new_new_n481_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n580_));
  NA2        g558(.A(new_new_n130_), .B(i_9_), .Y(new_new_n581_));
  NA3        g559(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n46_), .B(i_1_), .Y(new_new_n583_));
  NA3        g561(.A(new_new_n583_), .B(new_new_n241_), .C(new_new_n44_), .Y(new_new_n584_));
  OAI220     g562(.A0(new_new_n584_), .A1(new_new_n582_), .B0(new_new_n581_), .B1(new_new_n933_), .Y(new_new_n585_));
  NA3        g563(.A(new_new_n569_), .B(new_new_n283_), .C(i_6_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n586_), .B(new_new_n23_), .Y(new_new_n587_));
  AOI210     g565(.A0(new_new_n428_), .A1(new_new_n381_), .B0(new_new_n225_), .Y(new_new_n588_));
  NO2        g566(.A(new_new_n588_), .B(new_new_n544_), .Y(new_new_n589_));
  NAi21      g567(.An(new_new_n580_), .B(new_new_n83_), .Y(new_new_n590_));
  NO2        g568(.A(i_11_), .B(new_new_n37_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n24_), .Y(new_new_n592_));
  INV        g570(.A(new_new_n590_), .Y(new_new_n593_));
  OR4        g571(.A(new_new_n593_), .B(new_new_n589_), .C(new_new_n587_), .D(new_new_n585_), .Y(new_new_n594_));
  NO3        g572(.A(new_new_n594_), .B(new_new_n579_), .C(new_new_n575_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n221_), .B(new_new_n92_), .Y(new_new_n596_));
  NO2        g574(.A(new_new_n596_), .B(new_new_n557_), .Y(new_new_n597_));
  NA2        g575(.A(new_new_n597_), .B(i_1_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n598_), .B(new_new_n551_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n599_), .B(new_new_n46_), .Y(new_new_n600_));
  NA2        g578(.A(i_3_), .B(new_new_n184_), .Y(new_new_n601_));
  NO2        g579(.A(new_new_n601_), .B(new_new_n106_), .Y(new_new_n602_));
  AN2        g580(.A(new_new_n602_), .B(new_new_n485_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n77_), .B(i_9_), .Y(new_new_n604_));
  NA2        g582(.A(i_1_), .B(i_3_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n408_), .B(new_new_n84_), .Y(new_new_n606_));
  AOI210     g584(.A0(i_11_), .A1(new_new_n517_), .B0(new_new_n606_), .Y(new_new_n607_));
  NO2        g585(.A(new_new_n607_), .B(new_new_n605_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n608_), .B(new_new_n603_), .Y(new_new_n609_));
  NA4        g587(.A(new_new_n609_), .B(new_new_n600_), .C(new_new_n595_), .D(new_new_n573_), .Y(new_new_n610_));
  NO3        g588(.A(new_new_n429_), .B(i_3_), .C(i_7_), .Y(new_new_n611_));
  NOi21      g589(.An(new_new_n611_), .B(i_10_), .Y(new_new_n612_));
  OA210      g590(.A0(new_new_n612_), .A1(new_new_n228_), .B0(new_new_n77_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n337_), .B(new_new_n336_), .Y(new_new_n614_));
  NA3        g592(.A(new_new_n435_), .B(new_new_n464_), .C(new_new_n46_), .Y(new_new_n615_));
  NO3        g593(.A(new_new_n430_), .B(new_new_n546_), .C(new_new_n77_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(new_new_n25_), .Y(new_new_n617_));
  NA3        g595(.A(new_new_n151_), .B(new_new_n76_), .C(new_new_n77_), .Y(new_new_n618_));
  NA4        g596(.A(new_new_n618_), .B(new_new_n617_), .C(new_new_n615_), .D(new_new_n614_), .Y(new_new_n619_));
  OAI210     g597(.A0(new_new_n619_), .A1(new_new_n613_), .B0(i_1_), .Y(new_new_n620_));
  AOI210     g598(.A0(new_new_n241_), .A1(new_new_n88_), .B0(i_1_), .Y(new_new_n621_));
  NO2        g599(.A(new_new_n335_), .B(i_2_), .Y(new_new_n622_));
  NA2        g600(.A(new_new_n622_), .B(new_new_n621_), .Y(new_new_n623_));
  AOI210     g601(.A0(new_new_n623_), .A1(new_new_n620_), .B0(i_13_), .Y(new_new_n624_));
  OR2        g602(.A(i_11_), .B(i_7_), .Y(new_new_n625_));
  AOI220     g603(.A0(new_new_n422_), .A1(new_new_n151_), .B0(i_2_), .B1(new_new_n130_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n626_), .B(new_new_n44_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n228_), .B(new_new_n123_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n41_), .Y(new_new_n629_));
  AOI210     g607(.A0(new_new_n627_), .A1(new_new_n298_), .B0(new_new_n629_), .Y(new_new_n630_));
  INV        g608(.A(new_new_n106_), .Y(new_new_n631_));
  AOI220     g609(.A0(new_new_n631_), .A1(new_new_n64_), .B0(new_new_n352_), .B1(new_new_n583_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n226_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n399_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n634_));
  NOi31      g612(.An(new_new_n634_), .B(new_new_n538_), .C(new_new_n44_), .Y(new_new_n635_));
  NA2        g613(.A(new_new_n119_), .B(i_13_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n582_), .B(new_new_n106_), .Y(new_new_n637_));
  INV        g615(.A(new_new_n637_), .Y(new_new_n638_));
  OAI220     g616(.A0(new_new_n638_), .A1(new_new_n63_), .B0(new_new_n636_), .B1(new_new_n621_), .Y(new_new_n639_));
  NO3        g617(.A(new_new_n63_), .B(new_new_n32_), .C(new_new_n92_), .Y(new_new_n640_));
  NA2        g618(.A(new_new_n26_), .B(new_new_n184_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(i_7_), .Y(new_new_n642_));
  NO3        g620(.A(new_new_n430_), .B(new_new_n221_), .C(new_new_n77_), .Y(new_new_n643_));
  AOI210     g621(.A0(new_new_n643_), .A1(new_new_n642_), .B0(new_new_n640_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n553_), .Y(new_new_n645_));
  NO4        g623(.A(new_new_n645_), .B(new_new_n639_), .C(new_new_n635_), .D(new_new_n633_), .Y(new_new_n646_));
  OR2        g624(.A(i_11_), .B(i_6_), .Y(new_new_n647_));
  NA3        g625(.A(new_new_n542_), .B(new_new_n641_), .C(i_7_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n648_), .A1(new_new_n638_), .B0(new_new_n647_), .Y(new_new_n649_));
  NA3        g627(.A(new_new_n373_), .B(i_10_), .C(new_new_n88_), .Y(new_new_n650_));
  NA2        g628(.A(new_new_n574_), .B(i_13_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n93_), .B(new_new_n641_), .Y(new_new_n652_));
  NAi21      g630(.An(i_11_), .B(i_12_), .Y(new_new_n653_));
  NOi41      g631(.An(new_new_n102_), .B(new_new_n653_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n654_));
  NO3        g632(.A(new_new_n430_), .B(new_new_n528_), .C(new_new_n546_), .Y(new_new_n655_));
  AOI220     g633(.A0(new_new_n655_), .A1(new_new_n279_), .B0(new_new_n654_), .B1(new_new_n652_), .Y(new_new_n656_));
  NA3        g634(.A(new_new_n656_), .B(new_new_n651_), .C(new_new_n650_), .Y(new_new_n657_));
  OAI210     g635(.A0(new_new_n657_), .A1(new_new_n649_), .B0(new_new_n57_), .Y(new_new_n658_));
  NO2        g636(.A(i_2_), .B(i_12_), .Y(new_new_n659_));
  NA2        g637(.A(new_new_n221_), .B(new_new_n334_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n120_), .B(i_2_), .Y(new_new_n661_));
  NA2        g639(.A(new_new_n661_), .B(new_new_n571_), .Y(new_new_n662_));
  NA2        g640(.A(new_new_n662_), .B(new_new_n660_), .Y(new_new_n663_));
  NA3        g641(.A(new_new_n663_), .B(new_new_n45_), .C(new_new_n210_), .Y(new_new_n664_));
  NA4        g642(.A(new_new_n664_), .B(new_new_n658_), .C(new_new_n646_), .D(new_new_n630_), .Y(new_new_n665_));
  OR4        g643(.A(new_new_n665_), .B(new_new_n624_), .C(new_new_n610_), .D(new_new_n556_), .Y(mai5));
  AOI210     g644(.A0(new_new_n597_), .A1(new_new_n244_), .B0(new_new_n380_), .Y(new_new_n667_));
  AN2        g645(.A(new_new_n24_), .B(i_10_), .Y(new_new_n668_));
  NA3        g646(.A(new_new_n668_), .B(new_new_n659_), .C(new_new_n99_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n543_), .B(i_11_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n80_), .B(new_new_n670_), .Y(new_new_n671_));
  NA3        g649(.A(new_new_n671_), .B(new_new_n669_), .C(new_new_n667_), .Y(new_new_n672_));
  NO3        g650(.A(i_11_), .B(new_new_n221_), .C(i_13_), .Y(new_new_n673_));
  NA2        g651(.A(i_12_), .B(i_8_), .Y(new_new_n674_));
  INV        g652(.A(new_new_n398_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n283_), .B(new_new_n521_), .Y(new_new_n676_));
  INV        g654(.A(new_new_n676_), .Y(new_new_n677_));
  NO2        g655(.A(new_new_n677_), .B(new_new_n672_), .Y(new_new_n678_));
  INV        g656(.A(new_new_n162_), .Y(new_new_n679_));
  OAI210     g657(.A0(new_new_n622_), .A1(new_new_n400_), .B0(new_new_n102_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n680_), .B(new_new_n679_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n408_), .B(new_new_n26_), .Y(new_new_n682_));
  AOI210     g660(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n379_), .Y(new_new_n683_));
  AOI210     g661(.A0(new_new_n683_), .A1(i_2_), .B0(new_new_n681_), .Y(new_new_n684_));
  INV        g662(.A(new_new_n163_), .Y(new_new_n685_));
  NO3        g663(.A(new_new_n558_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n686_));
  AOI210     g664(.A0(new_new_n685_), .A1(new_new_n80_), .B0(new_new_n686_), .Y(new_new_n687_));
  NO2        g665(.A(new_new_n687_), .B(new_new_n184_), .Y(new_new_n688_));
  OA210      g666(.A0(new_new_n559_), .A1(new_new_n118_), .B0(i_13_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n190_), .B(new_new_n192_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n143_), .B(i_8_), .Y(new_new_n691_));
  AOI210     g669(.A0(new_new_n691_), .A1(new_new_n690_), .B0(new_new_n338_), .Y(new_new_n692_));
  AOI210     g670(.A0(new_new_n196_), .A1(new_new_n140_), .B0(new_new_n464_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n693_), .B(new_new_n381_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n93_), .B(new_new_n44_), .Y(new_new_n695_));
  INV        g673(.A(new_new_n268_), .Y(new_new_n696_));
  NA4        g674(.A(new_new_n696_), .B(new_new_n272_), .C(new_new_n116_), .D(new_new_n42_), .Y(new_new_n697_));
  OAI210     g675(.A0(new_new_n697_), .A1(new_new_n695_), .B0(new_new_n694_), .Y(new_new_n698_));
  NO4        g676(.A(new_new_n698_), .B(new_new_n692_), .C(new_new_n689_), .D(new_new_n688_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n521_), .B(new_new_n28_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n673_), .B(new_new_n249_), .Y(new_new_n701_));
  NA2        g679(.A(new_new_n701_), .B(new_new_n700_), .Y(new_new_n702_));
  NA2        g680(.A(new_new_n702_), .B(new_new_n46_), .Y(new_new_n703_));
  NA4        g681(.A(new_new_n703_), .B(new_new_n699_), .C(new_new_n684_), .D(new_new_n678_), .Y(mai6));
  NO3        g682(.A(i_9_), .B(new_new_n274_), .C(i_1_), .Y(new_new_n705_));
  NO2        g683(.A(new_new_n177_), .B(new_new_n131_), .Y(new_new_n706_));
  OAI210     g684(.A0(new_new_n706_), .A1(new_new_n705_), .B0(new_new_n661_), .Y(new_new_n707_));
  NA4        g685(.A(new_new_n356_), .B(new_new_n434_), .C(new_new_n63_), .D(new_new_n92_), .Y(new_new_n708_));
  INV        g686(.A(new_new_n708_), .Y(new_new_n709_));
  NO2        g687(.A(i_11_), .B(i_9_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n709_), .B(new_new_n294_), .Y(new_new_n711_));
  AO210      g689(.A0(new_new_n711_), .A1(new_new_n707_), .B0(i_12_), .Y(new_new_n712_));
  NA2        g690(.A(new_new_n339_), .B(new_new_n301_), .Y(new_new_n713_));
  NA2        g691(.A(new_new_n528_), .B(new_new_n57_), .Y(new_new_n714_));
  NA2        g692(.A(new_new_n612_), .B(new_new_n63_), .Y(new_new_n715_));
  NA4        g693(.A(new_new_n563_), .B(new_new_n715_), .C(new_new_n714_), .D(new_new_n713_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n187_), .Y(new_new_n717_));
  AOI220     g695(.A0(new_new_n717_), .A1(new_new_n710_), .B0(new_new_n716_), .B1(new_new_n65_), .Y(new_new_n718_));
  INV        g696(.A(new_new_n293_), .Y(new_new_n719_));
  NA2        g697(.A(new_new_n67_), .B(new_new_n123_), .Y(new_new_n720_));
  INV        g698(.A(new_new_n116_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n721_), .B(new_new_n46_), .Y(new_new_n722_));
  AOI210     g700(.A0(new_new_n722_), .A1(new_new_n720_), .B0(new_new_n719_), .Y(new_new_n723_));
  NO2        g701(.A(new_new_n32_), .B(i_11_), .Y(new_new_n724_));
  NA3        g702(.A(new_new_n724_), .B(new_new_n426_), .C(new_new_n356_), .Y(new_new_n725_));
  OAI210     g703(.A0(new_new_n611_), .A1(new_new_n509_), .B0(new_new_n508_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n726_), .B(new_new_n725_), .Y(new_new_n727_));
  OR2        g705(.A(new_new_n727_), .B(new_new_n723_), .Y(new_new_n728_));
  NO2        g706(.A(new_new_n625_), .B(i_2_), .Y(new_new_n729_));
  NA2        g707(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n730_));
  OAI210     g708(.A0(new_new_n730_), .A1(new_new_n372_), .B0(new_new_n324_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n731_), .B(new_new_n729_), .Y(new_new_n732_));
  AO220      g710(.A0(new_new_n323_), .A1(new_new_n314_), .B0(new_new_n362_), .B1(i_8_), .Y(new_new_n733_));
  NA3        g711(.A(new_new_n733_), .B(new_new_n234_), .C(i_7_), .Y(new_new_n734_));
  OR2        g712(.A(new_new_n559_), .B(new_new_n400_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n735_), .B(new_new_n139_), .Y(new_new_n736_));
  OR2        g714(.A(new_new_n675_), .B(new_new_n36_), .Y(new_new_n737_));
  NA4        g715(.A(new_new_n737_), .B(new_new_n736_), .C(new_new_n734_), .D(new_new_n732_), .Y(new_new_n738_));
  OAI210     g716(.A0(i_6_), .A1(i_11_), .B0(new_new_n78_), .Y(new_new_n739_));
  NA2        g717(.A(new_new_n739_), .B(new_new_n508_), .Y(new_new_n740_));
  NA3        g718(.A(new_new_n338_), .B(new_new_n222_), .C(new_new_n139_), .Y(new_new_n741_));
  OAI210     g719(.A0(new_new_n362_), .A1(new_new_n193_), .B0(new_new_n62_), .Y(new_new_n742_));
  NA4        g720(.A(new_new_n742_), .B(new_new_n741_), .C(new_new_n740_), .D(new_new_n545_), .Y(new_new_n743_));
  AO210      g721(.A0(new_new_n464_), .A1(new_new_n46_), .B0(new_new_n79_), .Y(new_new_n744_));
  NA3        g722(.A(new_new_n744_), .B(new_new_n435_), .C(new_new_n205_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n400_), .A1(new_new_n398_), .B0(new_new_n507_), .Y(new_new_n746_));
  NA2        g724(.A(new_new_n103_), .B(new_new_n371_), .Y(new_new_n747_));
  NA3        g725(.A(new_new_n747_), .B(new_new_n746_), .C(new_new_n745_), .Y(new_new_n748_));
  NO4        g726(.A(new_new_n748_), .B(new_new_n743_), .C(new_new_n738_), .D(new_new_n728_), .Y(new_new_n749_));
  NA4        g727(.A(new_new_n749_), .B(new_new_n718_), .C(new_new_n712_), .D(new_new_n346_), .Y(mai3));
  NA2        g728(.A(i_6_), .B(i_7_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n751_), .B(i_0_), .Y(new_new_n752_));
  NO2        g730(.A(i_11_), .B(new_new_n221_), .Y(new_new_n753_));
  OAI210     g731(.A0(new_new_n752_), .A1(new_new_n257_), .B0(new_new_n753_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n184_), .Y(new_new_n755_));
  NO3        g733(.A(new_new_n404_), .B(new_new_n81_), .C(new_new_n44_), .Y(new_new_n756_));
  OA210      g734(.A0(new_new_n756_), .A1(new_new_n755_), .B0(new_new_n165_), .Y(new_new_n757_));
  INV        g735(.A(new_new_n741_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n758_), .B(new_new_n40_), .Y(new_new_n759_));
  NO2        g737(.A(new_new_n567_), .B(new_new_n408_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n373_), .B(new_new_n45_), .Y(new_new_n761_));
  AOI210     g739(.A0(new_new_n934_), .A1(new_new_n759_), .B0(new_new_n48_), .Y(new_new_n762_));
  NO4        g740(.A(new_new_n342_), .B(new_new_n349_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n634_), .B(new_new_n604_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n299_), .B(i_5_), .Y(new_new_n765_));
  OAI220     g743(.A0(new_new_n765_), .A1(new_new_n764_), .B0(new_new_n938_), .B1(new_new_n57_), .Y(new_new_n766_));
  NOi21      g744(.An(i_5_), .B(i_9_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n767_), .B(new_new_n396_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n241_), .B(new_new_n428_), .Y(new_new_n769_));
  NO2        g747(.A(new_new_n166_), .B(new_new_n140_), .Y(new_new_n770_));
  INV        g748(.A(new_new_n770_), .Y(new_new_n771_));
  OAI220     g749(.A0(new_new_n771_), .A1(new_new_n172_), .B0(new_new_n769_), .B1(new_new_n768_), .Y(new_new_n772_));
  NO4        g750(.A(new_new_n772_), .B(new_new_n766_), .C(new_new_n762_), .D(new_new_n757_), .Y(new_new_n773_));
  NA2        g751(.A(new_new_n177_), .B(new_new_n24_), .Y(new_new_n774_));
  NO2        g752(.A(new_new_n37_), .B(new_new_n774_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n279_), .B(new_new_n121_), .Y(new_new_n776_));
  NAi21      g754(.An(new_new_n152_), .B(i_5_), .Y(new_new_n777_));
  NO2        g755(.A(new_new_n776_), .B(new_new_n364_), .Y(new_new_n778_));
  NO2        g756(.A(new_new_n778_), .B(new_new_n775_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n518_), .B(i_0_), .Y(new_new_n780_));
  NO3        g758(.A(new_new_n780_), .B(new_new_n351_), .C(new_new_n80_), .Y(new_new_n781_));
  INV        g759(.A(new_new_n781_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n673_), .B(new_new_n294_), .Y(new_new_n783_));
  OAI220     g761(.A0(i_6_), .A1(new_new_n783_), .B0(new_new_n592_), .B1(new_new_n482_), .Y(new_new_n784_));
  NA2        g762(.A(i_0_), .B(i_10_), .Y(new_new_n785_));
  NO4        g763(.A(new_new_n106_), .B(new_new_n53_), .C(new_new_n601_), .D(i_5_), .Y(new_new_n786_));
  AN2        g764(.A(new_new_n786_), .B(i_10_), .Y(new_new_n787_));
  NA2        g765(.A(new_new_n177_), .B(new_new_n76_), .Y(new_new_n788_));
  NA2        g766(.A(new_new_n512_), .B(i_4_), .Y(new_new_n789_));
  NA2        g767(.A(new_new_n180_), .B(new_new_n192_), .Y(new_new_n790_));
  OAI220     g768(.A0(new_new_n790_), .A1(new_new_n783_), .B0(new_new_n789_), .B1(new_new_n788_), .Y(new_new_n791_));
  NO3        g769(.A(new_new_n791_), .B(new_new_n787_), .C(new_new_n784_), .Y(new_new_n792_));
  NA3        g770(.A(new_new_n792_), .B(new_new_n782_), .C(new_new_n779_), .Y(new_new_n793_));
  NA2        g771(.A(i_11_), .B(i_9_), .Y(new_new_n794_));
  NO3        g772(.A(i_12_), .B(new_new_n794_), .C(new_new_n544_), .Y(new_new_n795_));
  AN2        g773(.A(new_new_n795_), .B(i_10_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n48_), .B(i_7_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n360_), .B(new_new_n170_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n798_), .B(new_new_n150_), .Y(new_new_n799_));
  NO2        g777(.A(new_new_n794_), .B(new_new_n65_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n166_), .B(i_0_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n426_), .B(new_new_n216_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n337_), .B(i_4_), .Y(new_new_n803_));
  OAI220     g781(.A0(new_new_n803_), .A1(new_new_n768_), .B0(new_new_n802_), .B1(new_new_n166_), .Y(new_new_n804_));
  NO3        g782(.A(new_new_n804_), .B(new_new_n799_), .C(new_new_n796_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n591_), .B(new_new_n113_), .Y(new_new_n806_));
  NO2        g784(.A(i_6_), .B(new_new_n806_), .Y(new_new_n807_));
  AOI210     g785(.A0(new_new_n399_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n808_));
  NA2        g786(.A(new_new_n162_), .B(new_new_n94_), .Y(new_new_n809_));
  NOi32      g787(.An(new_new_n808_), .Bn(new_new_n180_), .C(new_new_n809_), .Y(new_new_n810_));
  NA2        g788(.A(i_10_), .B(new_new_n294_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n811_), .B(new_new_n761_), .Y(new_new_n812_));
  NO3        g790(.A(new_new_n812_), .B(new_new_n810_), .C(new_new_n807_), .Y(new_new_n813_));
  NOi21      g791(.An(i_7_), .B(i_5_), .Y(new_new_n814_));
  NOi31      g792(.An(new_new_n814_), .B(i_0_), .C(new_new_n653_), .Y(new_new_n815_));
  NA3        g793(.A(new_new_n815_), .B(new_new_n350_), .C(i_6_), .Y(new_new_n816_));
  OA210      g794(.A0(new_new_n809_), .A1(new_new_n463_), .B0(new_new_n816_), .Y(new_new_n817_));
  NO3        g795(.A(new_new_n367_), .B(new_new_n326_), .C(new_new_n322_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n235_), .B(new_new_n284_), .Y(new_new_n819_));
  INV        g797(.A(new_new_n818_), .Y(new_new_n820_));
  NA4        g798(.A(new_new_n820_), .B(new_new_n817_), .C(new_new_n813_), .D(new_new_n805_), .Y(new_new_n821_));
  OA210      g799(.A0(new_new_n426_), .A1(new_new_n208_), .B0(new_new_n425_), .Y(new_new_n822_));
  NA3        g800(.A(new_new_n425_), .B(new_new_n373_), .C(new_new_n45_), .Y(new_new_n823_));
  OAI210     g801(.A0(new_new_n777_), .A1(i_6_), .B0(new_new_n823_), .Y(new_new_n824_));
  NA2        g802(.A(new_new_n800_), .B(new_new_n272_), .Y(new_new_n825_));
  NA2        g803(.A(new_new_n179_), .B(new_new_n825_), .Y(new_new_n826_));
  AOI220     g804(.A0(new_new_n826_), .A1(new_new_n426_), .B0(new_new_n824_), .B1(new_new_n65_), .Y(new_new_n827_));
  NO2        g805(.A(new_new_n67_), .B(new_new_n674_), .Y(new_new_n828_));
  AOI210     g806(.A0(new_new_n165_), .A1(i_10_), .B0(new_new_n828_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n829_), .B(new_new_n47_), .Y(new_new_n830_));
  NO3        g808(.A(i_5_), .B(new_new_n321_), .C(new_new_n24_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n492_), .B(new_new_n831_), .Y(new_new_n832_));
  NAi21      g810(.An(i_9_), .B(i_5_), .Y(new_new_n833_));
  NO2        g811(.A(new_new_n833_), .B(new_new_n367_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n541_), .B(new_new_n96_), .Y(new_new_n835_));
  AOI220     g813(.A0(new_new_n835_), .A1(i_0_), .B0(new_new_n834_), .B1(new_new_n559_), .Y(new_new_n836_));
  OAI220     g814(.A0(new_new_n836_), .A1(new_new_n77_), .B0(new_new_n832_), .B1(new_new_n163_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n830_), .Y(new_new_n838_));
  NA2        g816(.A(new_new_n838_), .B(new_new_n827_), .Y(new_new_n839_));
  NO3        g817(.A(new_new_n839_), .B(new_new_n821_), .C(new_new_n793_), .Y(new_new_n840_));
  NO2        g818(.A(i_0_), .B(new_new_n653_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n65_), .B(new_new_n44_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n785_), .B(new_new_n842_), .Y(new_new_n843_));
  NO2        g821(.A(i_5_), .B(new_new_n25_), .Y(new_new_n844_));
  AO220      g822(.A0(new_new_n844_), .A1(new_new_n843_), .B0(new_new_n841_), .B1(new_new_n165_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n714_), .B(new_new_n809_), .Y(new_new_n846_));
  AOI210     g824(.A0(new_new_n845_), .A1(new_new_n312_), .B0(new_new_n846_), .Y(new_new_n847_));
  NA3        g825(.A(new_new_n138_), .B(new_new_n604_), .C(new_new_n65_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n726_), .B(new_new_n367_), .Y(new_new_n849_));
  NA3        g827(.A(new_new_n752_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n753_), .B(i_9_), .Y(new_new_n851_));
  AOI210     g829(.A0(new_new_n850_), .A1(new_new_n446_), .B0(new_new_n851_), .Y(new_new_n852_));
  NA2        g830(.A(new_new_n227_), .B(new_new_n215_), .Y(new_new_n853_));
  AOI210     g831(.A0(new_new_n853_), .A1(new_new_n780_), .B0(new_new_n144_), .Y(new_new_n854_));
  NO3        g832(.A(new_new_n854_), .B(new_new_n852_), .C(new_new_n849_), .Y(new_new_n855_));
  NA3        g833(.A(new_new_n855_), .B(new_new_n848_), .C(new_new_n847_), .Y(new_new_n856_));
  NA3        g834(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n857_));
  NA2        g835(.A(new_new_n797_), .B(new_new_n438_), .Y(new_new_n858_));
  AOI210     g836(.A0(new_new_n857_), .A1(new_new_n152_), .B0(new_new_n858_), .Y(new_new_n859_));
  INV        g837(.A(new_new_n859_), .Y(new_new_n860_));
  NA2        g838(.A(new_new_n513_), .B(new_new_n67_), .Y(new_new_n861_));
  NO3        g839(.A(new_new_n197_), .B(new_new_n349_), .C(i_0_), .Y(new_new_n862_));
  OAI210     g840(.A0(new_new_n862_), .A1(new_new_n68_), .B0(i_13_), .Y(new_new_n863_));
  INV        g841(.A(new_new_n205_), .Y(new_new_n864_));
  OAI220     g842(.A0(new_new_n477_), .A1(new_new_n131_), .B0(new_new_n578_), .B1(new_new_n553_), .Y(new_new_n865_));
  NA3        g843(.A(new_new_n865_), .B(i_7_), .C(new_new_n864_), .Y(new_new_n866_));
  NA4        g844(.A(new_new_n866_), .B(new_new_n863_), .C(new_new_n861_), .D(new_new_n860_), .Y(new_new_n867_));
  NO2        g845(.A(new_new_n226_), .B(new_new_n84_), .Y(new_new_n868_));
  AOI210     g846(.A0(new_new_n868_), .A1(new_new_n841_), .B0(new_new_n100_), .Y(new_new_n869_));
  NA2        g847(.A(new_new_n814_), .B(new_new_n438_), .Y(new_new_n870_));
  INV        g848(.A(new_new_n167_), .Y(new_new_n871_));
  OA220      g849(.A0(new_new_n871_), .A1(new_new_n870_), .B0(new_new_n869_), .B1(i_5_), .Y(new_new_n872_));
  AOI210     g850(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n166_), .Y(new_new_n873_));
  NA2        g851(.A(new_new_n873_), .B(new_new_n822_), .Y(new_new_n874_));
  NA3        g852(.A(new_new_n797_), .B(new_new_n257_), .C(new_new_n215_), .Y(new_new_n875_));
  INV        g853(.A(new_new_n875_), .Y(new_new_n876_));
  NA3        g854(.A(new_new_n356_), .B(new_new_n300_), .C(new_new_n207_), .Y(new_new_n877_));
  INV        g855(.A(new_new_n877_), .Y(new_new_n878_));
  NOi31      g856(.An(new_new_n355_), .B(new_new_n842_), .C(new_new_n223_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n794_), .B(new_new_n205_), .C(new_new_n181_), .Y(new_new_n880_));
  NO4        g858(.A(new_new_n880_), .B(new_new_n879_), .C(new_new_n878_), .D(new_new_n876_), .Y(new_new_n881_));
  NA4        g859(.A(new_new_n881_), .B(new_new_n423_), .C(new_new_n874_), .D(new_new_n872_), .Y(new_new_n882_));
  NA3        g860(.A(new_new_n272_), .B(i_5_), .C(new_new_n184_), .Y(new_new_n883_));
  NA2        g861(.A(new_new_n883_), .B(new_new_n226_), .Y(new_new_n884_));
  NO4        g862(.A(new_new_n223_), .B(new_new_n197_), .C(i_0_), .D(i_12_), .Y(new_new_n885_));
  AOI220     g863(.A0(new_new_n885_), .A1(new_new_n884_), .B0(new_new_n709_), .B1(new_new_n167_), .Y(new_new_n886_));
  AN2        g864(.A(new_new_n785_), .B(new_new_n144_), .Y(new_new_n887_));
  NO3        g865(.A(new_new_n887_), .B(i_12_), .C(new_new_n580_), .Y(new_new_n888_));
  INV        g866(.A(new_new_n888_), .Y(new_new_n889_));
  NA3        g867(.A(new_new_n89_), .B(new_new_n517_), .C(i_11_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n814_), .B(new_new_n422_), .Y(new_new_n891_));
  OAI220     g869(.A0(i_7_), .A1(new_new_n883_), .B0(new_new_n891_), .B1(i_1_), .Y(new_new_n892_));
  NA2        g870(.A(new_new_n892_), .B(new_new_n801_), .Y(new_new_n893_));
  NA3        g871(.A(new_new_n893_), .B(new_new_n889_), .C(new_new_n886_), .Y(new_new_n894_));
  NO4        g872(.A(new_new_n894_), .B(new_new_n882_), .C(new_new_n867_), .D(new_new_n856_), .Y(new_new_n895_));
  OAI210     g873(.A0(new_new_n729_), .A1(new_new_n724_), .B0(new_new_n37_), .Y(new_new_n896_));
  NA3        g874(.A(new_new_n808_), .B(new_new_n334_), .C(i_5_), .Y(new_new_n897_));
  NA3        g875(.A(new_new_n897_), .B(new_new_n896_), .C(new_new_n937_), .Y(new_new_n898_));
  NA2        g876(.A(new_new_n898_), .B(new_new_n195_), .Y(new_new_n899_));
  NA2        g877(.A(new_new_n178_), .B(new_new_n180_), .Y(new_new_n900_));
  AO210      g878(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n900_), .Y(new_new_n901_));
  OAI210     g879(.A0(new_new_n552_), .A1(new_new_n550_), .B0(new_new_n283_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n902_), .B(new_new_n901_), .Y(new_new_n903_));
  NA2        g881(.A(new_new_n890_), .B(new_new_n413_), .Y(new_new_n904_));
  AOI210     g882(.A0(new_new_n903_), .A1(new_new_n48_), .B0(new_new_n904_), .Y(new_new_n905_));
  AOI210     g883(.A0(new_new_n905_), .A1(new_new_n899_), .B0(new_new_n65_), .Y(new_new_n906_));
  NO2        g884(.A(new_new_n510_), .B(new_new_n345_), .Y(new_new_n907_));
  NO2        g885(.A(new_new_n907_), .B(new_new_n679_), .Y(new_new_n908_));
  INV        g886(.A(new_new_n68_), .Y(new_new_n909_));
  AOI210     g887(.A0(new_new_n873_), .A1(new_new_n797_), .B0(new_new_n815_), .Y(new_new_n910_));
  AOI210     g888(.A0(new_new_n910_), .A1(new_new_n909_), .B0(new_new_n605_), .Y(new_new_n911_));
  NA2        g889(.A(i_8_), .B(new_new_n68_), .Y(new_new_n912_));
  NO2        g890(.A(new_new_n912_), .B(new_new_n221_), .Y(new_new_n913_));
  NO2        g891(.A(new_new_n913_), .B(new_new_n911_), .Y(new_new_n914_));
  OAI210     g892(.A0(new_new_n243_), .A1(new_new_n148_), .B0(new_new_n80_), .Y(new_new_n915_));
  NA3        g893(.A(new_new_n682_), .B(new_new_n257_), .C(new_new_n72_), .Y(new_new_n916_));
  AOI210     g894(.A0(new_new_n916_), .A1(new_new_n915_), .B0(i_11_), .Y(new_new_n917_));
  OAI210     g895(.A0(new_new_n935_), .A1(new_new_n808_), .B0(new_new_n195_), .Y(new_new_n918_));
  NA2        g896(.A(new_new_n154_), .B(i_5_), .Y(new_new_n919_));
  AOI210     g897(.A0(new_new_n918_), .A1(new_new_n690_), .B0(new_new_n919_), .Y(new_new_n920_));
  NA2        g898(.A(new_new_n819_), .B(new_new_n939_), .Y(new_new_n921_));
  NO2        g899(.A(new_new_n921_), .B(new_new_n653_), .Y(new_new_n922_));
  NO3        g900(.A(new_new_n833_), .B(new_new_n429_), .C(new_new_n233_), .Y(new_new_n923_));
  NO2        g901(.A(new_new_n923_), .B(new_new_n507_), .Y(new_new_n924_));
  INV        g902(.A(new_new_n327_), .Y(new_new_n925_));
  AOI210     g903(.A0(new_new_n925_), .A1(new_new_n924_), .B0(new_new_n41_), .Y(new_new_n926_));
  NO4        g904(.A(new_new_n926_), .B(new_new_n922_), .C(new_new_n920_), .D(new_new_n917_), .Y(new_new_n927_));
  OAI210     g905(.A0(new_new_n914_), .A1(i_4_), .B0(new_new_n927_), .Y(new_new_n928_));
  NO3        g906(.A(new_new_n928_), .B(new_new_n908_), .C(new_new_n906_), .Y(new_new_n929_));
  NA4        g907(.A(new_new_n929_), .B(new_new_n895_), .C(new_new_n840_), .D(new_new_n773_), .Y(mai4));
  INV        g908(.A(i_2_), .Y(new_new_n933_));
  INV        g909(.A(new_new_n760_), .Y(new_new_n934_));
  INV        g910(.A(i_12_), .Y(new_new_n935_));
  INV        g911(.A(new_new_n74_), .Y(new_new_n936_));
  INV        g912(.A(new_new_n151_), .Y(new_new_n937_));
  INV        g913(.A(new_new_n763_), .Y(new_new_n938_));
  INV        g914(.A(i_4_), .Y(new_new_n939_));
  INV        g915(.A(new_new_n229_), .Y(new_new_n940_));
  INV        g916(.A(new_new_n134_), .Y(new_new_n941_));
  INV        g917(.A(i_0_), .Y(new_new_n942_));
  INV        g918(.A(new_new_n378_), .Y(new_new_n943_));
  INV        g919(.A(i_3_), .Y(new_new_n944_));
  INV        g920(.A(i_6_), .Y(new_new_n945_));
  INV        g921(.A(new_new_n31_), .Y(new_new_n946_));
endmodule


