//Benchmark atmr_alu4_1266_0.125

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n123_, ori_ori_n124_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n504_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  OAI210     o027(.A0(ori_ori_n49_), .A1(i_3_), .B0(ori_ori_n47_), .Y(ori_ori_n50_));
  NO2        o028(.A(ori_ori_n50_), .B(ori_ori_n46_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n51_), .B(ori_ori_n45_), .Y(ori_ori_n53_));
  NO2        o031(.A(i_1_), .B(i_6_), .Y(ori_ori_n54_));
  NAi21      o032(.An(i_2_), .B(i_7_), .Y(ori_ori_n55_));
  INV        o033(.A(i_1_), .Y(ori_ori_n56_));
  NA2        o034(.A(ori_ori_n56_), .B(i_6_), .Y(ori_ori_n57_));
  NA3        o035(.A(ori_ori_n57_), .B(ori_ori_n55_), .C(ori_ori_n31_), .Y(ori_ori_n58_));
  NA2        o036(.A(i_1_), .B(i_10_), .Y(ori_ori_n59_));
  NO2        o037(.A(ori_ori_n59_), .B(i_6_), .Y(ori_ori_n60_));
  NAi21      o038(.An(ori_ori_n60_), .B(ori_ori_n58_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n62_));
  AOI210     o040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_1_), .B(i_6_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(ori_ori_n25_), .Y(ori_ori_n65_));
  INV        o043(.A(i_0_), .Y(ori_ori_n66_));
  NAi21      o044(.An(i_5_), .B(i_10_), .Y(ori_ori_n67_));
  NA2        o045(.A(i_5_), .B(i_9_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n67_), .B0(ori_ori_n66_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n65_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n63_), .A1(ori_ori_n62_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n61_), .B0(i_0_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_12_), .B(i_5_), .Y(ori_ori_n73_));
  INV        o051(.A(i_8_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n74_), .B(ori_ori_n54_), .Y(ori_ori_n75_));
  NO2        o053(.A(i_3_), .B(i_9_), .Y(ori_ori_n76_));
  NO2        o054(.A(i_3_), .B(i_7_), .Y(ori_ori_n77_));
  NO2        o055(.A(ori_ori_n76_), .B(ori_ori_n56_), .Y(ori_ori_n78_));
  INV        o056(.A(i_6_), .Y(ori_ori_n79_));
  NO2        o057(.A(i_2_), .B(i_7_), .Y(ori_ori_n80_));
  INV        o058(.A(ori_ori_n80_), .Y(ori_ori_n81_));
  OAI210     o059(.A0(ori_ori_n78_), .A1(ori_ori_n75_), .B0(ori_ori_n81_), .Y(ori_ori_n82_));
  NAi21      o060(.An(i_6_), .B(i_10_), .Y(ori_ori_n83_));
  NA2        o061(.A(i_6_), .B(i_9_), .Y(ori_ori_n84_));
  AOI210     o062(.A0(ori_ori_n84_), .A1(ori_ori_n83_), .B0(ori_ori_n56_), .Y(ori_ori_n85_));
  NA2        o063(.A(i_2_), .B(i_6_), .Y(ori_ori_n86_));
  NO2        o064(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n87_), .B(ori_ori_n85_), .Y(ori_ori_n88_));
  AOI210     o066(.A0(ori_ori_n88_), .A1(ori_ori_n82_), .B0(ori_ori_n73_), .Y(ori_ori_n89_));
  AN3        o067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n90_));
  NAi21      o068(.An(i_6_), .B(i_11_), .Y(ori_ori_n91_));
  NA2        o069(.A(ori_ori_n90_), .B(ori_ori_n32_), .Y(ori_ori_n92_));
  INV        o070(.A(i_7_), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n46_), .B(ori_ori_n93_), .Y(ori_ori_n94_));
  NO2        o072(.A(i_0_), .B(i_5_), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n95_), .B(ori_ori_n79_), .Y(ori_ori_n96_));
  NA2        o074(.A(i_12_), .B(i_3_), .Y(ori_ori_n97_));
  INV        o075(.A(ori_ori_n97_), .Y(ori_ori_n98_));
  NA3        o076(.A(ori_ori_n98_), .B(ori_ori_n96_), .C(ori_ori_n94_), .Y(ori_ori_n99_));
  NAi21      o077(.An(i_7_), .B(i_11_), .Y(ori_ori_n100_));
  AN2        o078(.A(i_2_), .B(i_10_), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n101_), .B(i_7_), .Y(ori_ori_n102_));
  OR2        o080(.A(ori_ori_n73_), .B(ori_ori_n54_), .Y(ori_ori_n103_));
  NA2        o081(.A(i_12_), .B(i_7_), .Y(ori_ori_n104_));
  NA2        o082(.A(i_11_), .B(i_12_), .Y(ori_ori_n105_));
  NA3        o083(.A(ori_ori_n105_), .B(ori_ori_n99_), .C(ori_ori_n92_), .Y(ori_ori_n106_));
  NOi21      o084(.An(i_1_), .B(i_5_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n107_), .B(i_11_), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n93_), .B(ori_ori_n37_), .Y(ori_ori_n109_));
  NA2        o087(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n110_), .B(ori_ori_n109_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(ori_ori_n46_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n84_), .B(ori_ori_n83_), .Y(ori_ori_n113_));
  NAi21      o091(.An(i_3_), .B(i_8_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(ori_ori_n55_), .Y(ori_ori_n115_));
  NOi31      o093(.An(ori_ori_n115_), .B(ori_ori_n113_), .C(ori_ori_n112_), .Y(ori_ori_n116_));
  NO2        o094(.A(i_1_), .B(ori_ori_n79_), .Y(ori_ori_n117_));
  NO2        o095(.A(i_6_), .B(i_5_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(i_3_), .Y(ori_ori_n119_));
  OAI220     o097(.A0(ori_ori_n119_), .A1(ori_ori_n100_), .B0(ori_ori_n116_), .B1(ori_ori_n108_), .Y(ori_ori_n120_));
  NO3        o098(.A(ori_ori_n120_), .B(ori_ori_n106_), .C(ori_ori_n89_), .Y(ori_ori_n121_));
  NA3        o099(.A(ori_ori_n121_), .B(ori_ori_n72_), .C(ori_ori_n53_), .Y(ori2));
  NO2        o100(.A(ori_ori_n56_), .B(ori_ori_n37_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n504_), .B(ori_ori_n123_), .Y(ori_ori_n124_));
  NA4        o102(.A(ori_ori_n124_), .B(ori_ori_n70_), .C(ori_ori_n62_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o103(.A(i_0_), .B(i_1_), .Y(ori_ori_n126_));
  NA2        o104(.A(i_2_), .B(i_3_), .Y(ori_ori_n127_));
  NO2        o105(.A(ori_ori_n127_), .B(i_4_), .Y(ori_ori_n128_));
  NA2        o106(.A(i_1_), .B(i_5_), .Y(ori_ori_n129_));
  OR2        o107(.A(i_0_), .B(i_1_), .Y(ori_ori_n130_));
  NO3        o108(.A(ori_ori_n130_), .B(ori_ori_n73_), .C(i_13_), .Y(ori_ori_n131_));
  NAi32      o109(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n132_));
  NAi21      o110(.An(ori_ori_n132_), .B(ori_ori_n131_), .Y(ori_ori_n133_));
  NOi21      o111(.An(i_4_), .B(i_10_), .Y(ori_ori_n134_));
  NOi21      o112(.An(i_4_), .B(i_9_), .Y(ori_ori_n135_));
  NOi21      o113(.An(i_11_), .B(i_13_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n66_), .B(ori_ori_n56_), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n66_), .B(i_5_), .Y(ori_ori_n139_));
  NO2        o117(.A(i_2_), .B(i_1_), .Y(ori_ori_n140_));
  NAi21      o118(.An(i_4_), .B(i_12_), .Y(ori_ori_n141_));
  INV        o119(.A(i_8_), .Y(ori_ori_n142_));
  NO2        o120(.A(i_3_), .B(i_8_), .Y(ori_ori_n143_));
  NO3        o121(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n95_), .B(ori_ori_n54_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_13_), .B(i_9_), .Y(ori_ori_n146_));
  NAi21      o124(.An(i_12_), .B(i_3_), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n148_));
  NA2        o126(.A(i_0_), .B(i_5_), .Y(ori_ori_n149_));
  INV        o127(.A(i_13_), .Y(ori_ori_n150_));
  NO2        o128(.A(i_12_), .B(ori_ori_n150_), .Y(ori_ori_n151_));
  NO2        o129(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n152_));
  OR2        o130(.A(i_8_), .B(i_7_), .Y(ori_ori_n153_));
  INV        o131(.A(i_12_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n44_), .B(ori_ori_n154_), .Y(ori_ori_n155_));
  NA2        o133(.A(i_2_), .B(i_1_), .Y(ori_ori_n156_));
  NO3        o134(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n157_));
  NAi21      o135(.An(i_4_), .B(i_3_), .Y(ori_ori_n158_));
  NO2        o136(.A(i_0_), .B(i_6_), .Y(ori_ori_n159_));
  NOi41      o137(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n160_));
  NO2        o138(.A(i_11_), .B(ori_ori_n150_), .Y(ori_ori_n161_));
  NOi21      o139(.An(i_1_), .B(i_6_), .Y(ori_ori_n162_));
  NAi21      o140(.An(i_3_), .B(i_7_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n154_), .B(i_9_), .Y(ori_ori_n164_));
  OR4        o142(.A(ori_ori_n164_), .B(ori_ori_n163_), .C(ori_ori_n162_), .D(ori_ori_n139_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n66_), .B(i_5_), .Y(ori_ori_n166_));
  NA2        o144(.A(i_3_), .B(i_9_), .Y(ori_ori_n167_));
  NAi21      o145(.An(i_7_), .B(i_10_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n168_), .B(ori_ori_n167_), .Y(ori_ori_n169_));
  NA3        o147(.A(ori_ori_n169_), .B(ori_ori_n166_), .C(ori_ori_n57_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n170_), .B(ori_ori_n165_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(ori_ori_n161_), .Y(ori_ori_n172_));
  NA2        o150(.A(i_12_), .B(i_6_), .Y(ori_ori_n173_));
  OR2        o151(.A(i_13_), .B(i_9_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n158_), .B(i_2_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n163_), .B(i_8_), .Y(ori_ori_n176_));
  NO3        o154(.A(i_12_), .B(ori_ori_n150_), .C(ori_ori_n37_), .Y(ori_ori_n177_));
  NO2        o155(.A(i_2_), .B(ori_ori_n93_), .Y(ori_ori_n178_));
  AN2        o156(.A(i_3_), .B(i_10_), .Y(ori_ori_n179_));
  NO2        o157(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n181_));
  NO2        o159(.A(i_2_), .B(i_3_), .Y(ori_ori_n182_));
  NO2        o160(.A(i_12_), .B(i_10_), .Y(ori_ori_n183_));
  NOi21      o161(.An(i_5_), .B(i_0_), .Y(ori_ori_n184_));
  NOi32      o162(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n185_));
  INV        o163(.A(ori_ori_n185_), .Y(ori_ori_n186_));
  NO2        o164(.A(ori_ori_n132_), .B(ori_ori_n130_), .Y(ori_ori_n187_));
  NOi32      o165(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n188_));
  NO2        o166(.A(i_1_), .B(ori_ori_n93_), .Y(ori_ori_n189_));
  NAi21      o167(.An(i_3_), .B(i_4_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n190_), .B(i_9_), .Y(ori_ori_n191_));
  AN2        o169(.A(i_6_), .B(i_7_), .Y(ori_ori_n192_));
  OAI210     o170(.A0(ori_ori_n192_), .A1(ori_ori_n189_), .B0(ori_ori_n191_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n190_), .B(i_10_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n193_), .B(ori_ori_n139_), .Y(ori_ori_n195_));
  AOI210     o173(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n196_));
  OAI210     o174(.A0(ori_ori_n196_), .A1(ori_ori_n140_), .B0(ori_ori_n194_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n197_), .B(i_5_), .Y(ori_ori_n198_));
  NO3        o176(.A(ori_ori_n198_), .B(ori_ori_n195_), .C(ori_ori_n187_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(ori_ori_n186_), .Y(ori_ori_n200_));
  AN2        o178(.A(i_12_), .B(i_5_), .Y(ori_ori_n201_));
  NO2        o179(.A(i_11_), .B(i_6_), .Y(ori_ori_n202_));
  NO2        o180(.A(i_5_), .B(i_10_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n79_), .B(ori_ori_n47_), .C(i_9_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_0_), .B(i_11_), .Y(ori_ori_n206_));
  NOi21      o184(.An(i_2_), .B(i_12_), .Y(ori_ori_n207_));
  NAi21      o185(.An(i_9_), .B(i_4_), .Y(ori_ori_n208_));
  OR2        o186(.A(i_13_), .B(i_10_), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n209_), .B(ori_ori_n105_), .C(ori_ori_n208_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n93_), .B(ori_ori_n25_), .Y(ori_ori_n211_));
  INV        o189(.A(ori_ori_n200_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n66_), .B(i_13_), .Y(ori_ori_n213_));
  NO2        o191(.A(i_10_), .B(i_9_), .Y(ori_ori_n214_));
  NAi21      o192(.An(i_12_), .B(i_8_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n215_), .B(i_3_), .Y(ori_ori_n216_));
  NO3        o194(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n173_), .B(ori_ori_n91_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  NA2        o197(.A(i_8_), .B(i_9_), .Y(ori_ori_n220_));
  NO2        o198(.A(i_7_), .B(i_2_), .Y(ori_ori_n221_));
  OR2        o199(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NA2        o200(.A(ori_ori_n177_), .B(ori_ori_n145_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n161_), .B(ori_ori_n180_), .Y(ori_ori_n225_));
  NO3        o203(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n226_));
  INV        o204(.A(ori_ori_n226_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n225_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n228_), .B(ori_ori_n224_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_11_), .B(i_1_), .Y(ori_ori_n230_));
  NOi21      o208(.An(i_2_), .B(i_7_), .Y(ori_ori_n231_));
  NA3        o209(.A(ori_ori_n160_), .B(ori_ori_n136_), .C(ori_ori_n118_), .Y(ori_ori_n232_));
  NA2        o210(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n130_), .B(i_3_), .Y(ori_ori_n234_));
  NAi31      o212(.An(ori_ori_n233_), .B(ori_ori_n234_), .C(ori_ori_n151_), .Y(ori_ori_n235_));
  NA3        o213(.A(ori_ori_n204_), .B(ori_ori_n138_), .C(ori_ori_n128_), .Y(ori_ori_n236_));
  NA3        o214(.A(ori_ori_n236_), .B(ori_ori_n235_), .C(ori_ori_n232_), .Y(ori_ori_n237_));
  INV        o215(.A(ori_ori_n237_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n217_), .B(ori_ori_n201_), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n226_), .B(ori_ori_n203_), .Y(ori_ori_n240_));
  NA2        o218(.A(ori_ori_n238_), .B(ori_ori_n229_), .Y(ori_ori_n241_));
  NA2        o219(.A(ori_ori_n201_), .B(ori_ori_n150_), .Y(ori_ori_n242_));
  NA2        o220(.A(ori_ori_n192_), .B(ori_ori_n188_), .Y(ori_ori_n243_));
  OR2        o221(.A(ori_ori_n242_), .B(ori_ori_n243_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n245_));
  AOI210     o223(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n210_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(ori_ori_n244_), .Y(ori_ori_n247_));
  NA3        o225(.A(ori_ori_n149_), .B(ori_ori_n64_), .C(ori_ori_n44_), .Y(ori_ori_n248_));
  NA2        o226(.A(ori_ori_n177_), .B(ori_ori_n77_), .Y(ori_ori_n249_));
  NO2        o227(.A(ori_ori_n248_), .B(ori_ori_n249_), .Y(ori_ori_n250_));
  NO3        o228(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n209_), .B(i_1_), .Y(ori_ori_n252_));
  NOi31      o230(.An(ori_ori_n252_), .B(ori_ori_n218_), .C(ori_ori_n66_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n79_), .B(ori_ori_n25_), .Y(ori_ori_n254_));
  NO2        o232(.A(ori_ori_n104_), .B(ori_ori_n23_), .Y(ori_ori_n255_));
  NO2        o233(.A(i_12_), .B(ori_ori_n79_), .Y(ori_ori_n256_));
  NO3        o234(.A(ori_ori_n250_), .B(ori_ori_n247_), .C(ori_ori_n241_), .Y(ori_ori_n257_));
  NA3        o235(.A(ori_ori_n257_), .B(ori_ori_n212_), .C(ori_ori_n172_), .Y(ori7));
  NO2        o236(.A(ori_ori_n86_), .B(ori_ori_n52_), .Y(ori_ori_n259_));
  NA2        o237(.A(i_11_), .B(ori_ori_n142_), .Y(ori_ori_n260_));
  NA3        o238(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n154_), .B(i_4_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n262_), .B(i_8_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n97_), .B(ori_ori_n261_), .Y(ori_ori_n264_));
  NA2        o242(.A(i_2_), .B(ori_ori_n79_), .Y(ori_ori_n265_));
  OAI210     o243(.A0(ori_ori_n80_), .A1(ori_ori_n143_), .B0(ori_ori_n144_), .Y(ori_ori_n266_));
  NO2        o244(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n267_));
  NA2        o245(.A(i_4_), .B(i_8_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n268_), .A1(ori_ori_n179_), .B0(ori_ori_n267_), .Y(ori_ori_n269_));
  OAI220     o247(.A0(ori_ori_n269_), .A1(ori_ori_n265_), .B0(ori_ori_n266_), .B1(i_13_), .Y(ori_ori_n270_));
  NO3        o248(.A(ori_ori_n270_), .B(ori_ori_n264_), .C(ori_ori_n259_), .Y(ori_ori_n271_));
  AOI210     o249(.A0(ori_ori_n114_), .A1(ori_ori_n55_), .B0(i_10_), .Y(ori_ori_n272_));
  AOI210     o250(.A0(ori_ori_n272_), .A1(ori_ori_n154_), .B0(ori_ori_n134_), .Y(ori_ori_n273_));
  OR2        o251(.A(i_6_), .B(i_10_), .Y(ori_ori_n274_));
  OR3        o252(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n275_));
  OR2        o253(.A(ori_ori_n273_), .B(ori_ori_n174_), .Y(ori_ori_n276_));
  AOI210     o254(.A0(ori_ori_n276_), .A1(ori_ori_n271_), .B0(ori_ori_n56_), .Y(ori_ori_n277_));
  NOi21      o255(.An(i_11_), .B(i_7_), .Y(ori_ori_n278_));
  AO210      o256(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n279_), .B(ori_ori_n278_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n146_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n281_), .B(ori_ori_n56_), .Y(ori_ori_n282_));
  NA2        o260(.A(ori_ori_n151_), .B(ori_ori_n56_), .Y(ori_ori_n283_));
  NO2        o261(.A(i_1_), .B(i_12_), .Y(ori_ori_n284_));
  INV        o262(.A(ori_ori_n283_), .Y(ori_ori_n285_));
  OAI210     o263(.A0(ori_ori_n285_), .A1(ori_ori_n282_), .B0(i_6_), .Y(ori_ori_n286_));
  NO2        o264(.A(i_6_), .B(i_11_), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n219_), .Y(ori_ori_n288_));
  NO3        o266(.A(ori_ori_n274_), .B(ori_ori_n153_), .C(ori_ori_n23_), .Y(ori_ori_n289_));
  AOI210     o267(.A0(i_1_), .A1(ori_ori_n169_), .B0(ori_ori_n289_), .Y(ori_ori_n290_));
  NO2        o268(.A(ori_ori_n290_), .B(ori_ori_n44_), .Y(ori_ori_n291_));
  INV        o269(.A(i_2_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n123_), .B(i_9_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n293_), .B(ori_ori_n292_), .Y(ori_ori_n295_));
  AOI210     o273(.A0(ori_ori_n230_), .A1(ori_ori_n211_), .B0(ori_ori_n157_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n296_), .B(ori_ori_n265_), .Y(ori_ori_n297_));
  NO2        o275(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n298_));
  OR2        o276(.A(ori_ori_n297_), .B(ori_ori_n295_), .Y(ori_ori_n299_));
  NO3        o277(.A(ori_ori_n299_), .B(ori_ori_n291_), .C(ori_ori_n288_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n154_), .B(ori_ori_n93_), .Y(ori_ori_n301_));
  NO2        o279(.A(ori_ori_n301_), .B(ori_ori_n278_), .Y(ori_ori_n302_));
  NA2        o280(.A(ori_ori_n302_), .B(i_1_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n303_), .B(ori_ori_n275_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n208_), .B(ori_ori_n79_), .Y(ori_ori_n305_));
  NA2        o283(.A(ori_ori_n304_), .B(ori_ori_n46_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n153_), .B(ori_ori_n44_), .Y(ori_ori_n307_));
  NO3        o285(.A(ori_ori_n307_), .B(ori_ori_n181_), .C(ori_ori_n155_), .Y(ori_ori_n308_));
  NO2        o286(.A(ori_ori_n105_), .B(ori_ori_n37_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n309_), .B(i_6_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n79_), .B(i_9_), .Y(ori_ori_n311_));
  NO2        o289(.A(ori_ori_n311_), .B(ori_ori_n56_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n312_), .B(ori_ori_n284_), .Y(ori_ori_n313_));
  NO4        o291(.A(ori_ori_n313_), .B(ori_ori_n310_), .C(ori_ori_n308_), .D(i_4_), .Y(ori_ori_n314_));
  INV        o292(.A(ori_ori_n314_), .Y(ori_ori_n315_));
  NA4        o293(.A(ori_ori_n315_), .B(ori_ori_n306_), .C(ori_ori_n300_), .D(ori_ori_n286_), .Y(ori_ori_n316_));
  AOI210     o294(.A0(ori_ori_n173_), .A1(ori_ori_n91_), .B0(i_1_), .Y(ori_ori_n317_));
  NO2        o295(.A(ori_ori_n190_), .B(i_2_), .Y(ori_ori_n318_));
  NA2        o296(.A(ori_ori_n318_), .B(ori_ori_n317_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n319_), .B(i_13_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n321_));
  INV        o299(.A(ori_ori_n321_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n231_), .B(ori_ori_n24_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n323_), .B(ori_ori_n305_), .Y(ori_ori_n324_));
  OAI220     o302(.A0(ori_ori_n324_), .A1(ori_ori_n41_), .B0(ori_ori_n322_), .B1(ori_ori_n86_), .Y(ori_ori_n325_));
  INV        o303(.A(ori_ori_n325_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n202_), .B(ori_ori_n294_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n327_), .B(ori_ori_n158_), .Y(ori_ori_n328_));
  NA2        o306(.A(ori_ori_n113_), .B(i_13_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n329_), .B(ori_ori_n317_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n26_), .B(ori_ori_n142_), .Y(ori_ori_n331_));
  AOI220     o309(.A0(ori_ori_n202_), .A1(ori_ori_n294_), .B0(ori_ori_n85_), .B1(ori_ori_n94_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n332_), .B(ori_ori_n263_), .Y(ori_ori_n333_));
  NO3        o311(.A(ori_ori_n333_), .B(ori_ori_n330_), .C(ori_ori_n328_), .Y(ori_ori_n334_));
  OR2        o312(.A(i_11_), .B(i_6_), .Y(ori_ori_n335_));
  NA3        o313(.A(ori_ori_n262_), .B(ori_ori_n331_), .C(i_7_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n336_), .B(ori_ori_n335_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n207_), .B(ori_ori_n267_), .C(ori_ori_n91_), .Y(ori_ori_n338_));
  NA2        o316(.A(ori_ori_n287_), .B(i_13_), .Y(ori_ori_n339_));
  NAi21      o317(.An(i_11_), .B(i_12_), .Y(ori_ori_n340_));
  NOi41      o318(.An(ori_ori_n102_), .B(ori_ori_n340_), .C(i_13_), .D(ori_ori_n79_), .Y(ori_ori_n341_));
  NA2        o319(.A(ori_ori_n341_), .B(ori_ori_n46_), .Y(ori_ori_n342_));
  NA3        o320(.A(ori_ori_n342_), .B(ori_ori_n339_), .C(ori_ori_n338_), .Y(ori_ori_n343_));
  OAI210     o321(.A0(ori_ori_n343_), .A1(ori_ori_n337_), .B0(ori_ori_n56_), .Y(ori_ori_n344_));
  NO2        o322(.A(i_2_), .B(i_12_), .Y(ori_ori_n345_));
  NA2        o323(.A(ori_ori_n189_), .B(ori_ori_n345_), .Y(ori_ori_n346_));
  INV        o324(.A(ori_ori_n346_), .Y(ori_ori_n347_));
  NA3        o325(.A(ori_ori_n347_), .B(ori_ori_n45_), .C(ori_ori_n150_), .Y(ori_ori_n348_));
  NA4        o326(.A(ori_ori_n348_), .B(ori_ori_n344_), .C(ori_ori_n334_), .D(ori_ori_n326_), .Y(ori_ori_n349_));
  OR4        o327(.A(ori_ori_n349_), .B(ori_ori_n320_), .C(ori_ori_n316_), .D(ori_ori_n277_), .Y(ori5));
  NA2        o328(.A(ori_ori_n302_), .B(ori_ori_n175_), .Y(ori_ori_n351_));
  AN2        o329(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n352_));
  NA3        o330(.A(ori_ori_n352_), .B(ori_ori_n345_), .C(ori_ori_n100_), .Y(ori_ori_n353_));
  NO2        o331(.A(ori_ori_n263_), .B(i_11_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n80_), .B(ori_ori_n354_), .Y(ori_ori_n355_));
  NA3        o333(.A(ori_ori_n355_), .B(ori_ori_n353_), .C(ori_ori_n351_), .Y(ori_ori_n356_));
  NO3        o334(.A(i_11_), .B(ori_ori_n154_), .C(i_13_), .Y(ori_ori_n357_));
  NO2        o335(.A(ori_ori_n110_), .B(ori_ori_n23_), .Y(ori_ori_n358_));
  NA2        o336(.A(i_12_), .B(i_8_), .Y(ori_ori_n359_));
  OAI210     o337(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n359_), .Y(ori_ori_n360_));
  INV        o338(.A(ori_ori_n214_), .Y(ori_ori_n361_));
  AOI220     o339(.A0(ori_ori_n182_), .A1(ori_ori_n255_), .B0(ori_ori_n360_), .B1(ori_ori_n358_), .Y(ori_ori_n362_));
  INV        o340(.A(ori_ori_n362_), .Y(ori_ori_n363_));
  NO2        o341(.A(ori_ori_n363_), .B(ori_ori_n356_), .Y(ori_ori_n364_));
  INV        o342(.A(ori_ori_n136_), .Y(ori_ori_n365_));
  INV        o343(.A(ori_ori_n160_), .Y(ori_ori_n366_));
  OAI210     o344(.A0(ori_ori_n318_), .A1(ori_ori_n216_), .B0(ori_ori_n102_), .Y(ori_ori_n367_));
  AOI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n366_), .B0(ori_ori_n365_), .Y(ori_ori_n368_));
  NO2        o346(.A(ori_ori_n220_), .B(ori_ori_n26_), .Y(ori_ori_n369_));
  NO2        o347(.A(ori_ori_n369_), .B(ori_ori_n211_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n370_), .B(i_2_), .Y(ori_ori_n371_));
  INV        o349(.A(ori_ori_n371_), .Y(ori_ori_n372_));
  AOI210     o350(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n209_), .Y(ori_ori_n373_));
  AOI210     o351(.A0(ori_ori_n373_), .A1(ori_ori_n372_), .B0(ori_ori_n368_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n141_), .B(ori_ori_n111_), .Y(ori_ori_n375_));
  OAI210     o353(.A0(ori_ori_n375_), .A1(ori_ori_n358_), .B0(i_2_), .Y(ori_ori_n376_));
  INV        o354(.A(ori_ori_n137_), .Y(ori_ori_n377_));
  NO3        o355(.A(ori_ori_n279_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n378_));
  AOI210     o356(.A0(ori_ori_n377_), .A1(ori_ori_n80_), .B0(ori_ori_n378_), .Y(ori_ori_n379_));
  AOI210     o357(.A0(ori_ori_n379_), .A1(ori_ori_n376_), .B0(ori_ori_n142_), .Y(ori_ori_n380_));
  OA210      o358(.A0(ori_ori_n280_), .A1(ori_ori_n112_), .B0(i_13_), .Y(ori_ori_n381_));
  AOI210     o359(.A0(ori_ori_n147_), .A1(ori_ori_n127_), .B0(ori_ori_n245_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n382_), .B(ori_ori_n211_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n94_), .B(ori_ori_n44_), .Y(ori_ori_n384_));
  INV        o362(.A(ori_ori_n178_), .Y(ori_ori_n385_));
  NA4        o363(.A(ori_ori_n385_), .B(ori_ori_n179_), .C(ori_ori_n110_), .D(ori_ori_n42_), .Y(ori_ori_n386_));
  OAI210     o364(.A0(ori_ori_n386_), .A1(ori_ori_n384_), .B0(ori_ori_n383_), .Y(ori_ori_n387_));
  NO3        o365(.A(ori_ori_n387_), .B(ori_ori_n381_), .C(ori_ori_n380_), .Y(ori_ori_n388_));
  NA2        o366(.A(ori_ori_n255_), .B(ori_ori_n28_), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n357_), .B(ori_ori_n176_), .Y(ori_ori_n390_));
  NA2        o368(.A(ori_ori_n390_), .B(ori_ori_n389_), .Y(ori_ori_n391_));
  NO2        o369(.A(ori_ori_n55_), .B(i_12_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n392_), .B(ori_ori_n112_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n393_), .B(ori_ori_n260_), .Y(ori_ori_n394_));
  AOI220     o372(.A0(ori_ori_n394_), .A1(ori_ori_n36_), .B0(ori_ori_n391_), .B1(ori_ori_n46_), .Y(ori_ori_n395_));
  NA4        o373(.A(ori_ori_n395_), .B(ori_ori_n388_), .C(ori_ori_n374_), .D(ori_ori_n364_), .Y(ori6));
  INV        o374(.A(ori_ori_n184_), .Y(ori_ori_n397_));
  OR2        o375(.A(ori_ori_n397_), .B(i_12_), .Y(ori_ori_n398_));
  NA2        o376(.A(ori_ori_n256_), .B(ori_ori_n56_), .Y(ori_ori_n399_));
  INV        o377(.A(ori_ori_n399_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n400_), .B(ori_ori_n66_), .Y(ori_ori_n401_));
  INV        o379(.A(ori_ori_n183_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n68_), .B(ori_ori_n117_), .Y(ori_ori_n403_));
  INV        o381(.A(ori_ori_n110_), .Y(ori_ori_n404_));
  NA2        o382(.A(ori_ori_n404_), .B(ori_ori_n46_), .Y(ori_ori_n405_));
  AOI210     o383(.A0(ori_ori_n405_), .A1(ori_ori_n403_), .B0(ori_ori_n402_), .Y(ori_ori_n406_));
  NO2        o384(.A(ori_ori_n162_), .B(i_9_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n407_), .B(ori_ori_n392_), .Y(ori_ori_n408_));
  AOI210     o386(.A0(ori_ori_n408_), .A1(ori_ori_n243_), .B0(ori_ori_n139_), .Y(ori_ori_n409_));
  NAi32      o387(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n335_), .B(ori_ori_n410_), .Y(ori_ori_n411_));
  OR3        o389(.A(ori_ori_n411_), .B(ori_ori_n409_), .C(ori_ori_n406_), .Y(ori_ori_n412_));
  BUFFER     o390(.A(ori_ori_n280_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n413_), .B(ori_ori_n126_), .Y(ori_ori_n414_));
  AO210      o392(.A0(ori_ori_n240_), .A1(ori_ori_n361_), .B0(ori_ori_n36_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(ori_ori_n414_), .Y(ori_ori_n416_));
  NO2        o394(.A(i_6_), .B(i_11_), .Y(ori_ori_n417_));
  NA2        o395(.A(ori_ori_n417_), .B(ori_ori_n251_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n205_), .B(ori_ori_n63_), .Y(ori_ori_n419_));
  NA3        o397(.A(ori_ori_n419_), .B(ori_ori_n418_), .C(ori_ori_n266_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n216_), .B(ori_ori_n214_), .Y(ori_ori_n421_));
  NA2        o399(.A(ori_ori_n103_), .B(ori_ori_n206_), .Y(ori_ori_n422_));
  NA2        o400(.A(ori_ori_n422_), .B(ori_ori_n421_), .Y(ori_ori_n423_));
  NO4        o401(.A(ori_ori_n423_), .B(ori_ori_n420_), .C(ori_ori_n416_), .D(ori_ori_n412_), .Y(ori_ori_n424_));
  NA4        o402(.A(ori_ori_n424_), .B(ori_ori_n401_), .C(ori_ori_n398_), .D(ori_ori_n199_), .Y(ori3));
  NA2        o403(.A(i_12_), .B(i_10_), .Y(ori_ori_n426_));
  NO2        o404(.A(i_11_), .B(ori_ori_n154_), .Y(ori_ori_n427_));
  NA2        o405(.A(ori_ori_n266_), .B(ori_ori_n193_), .Y(ori_ori_n428_));
  NA2        o406(.A(ori_ori_n428_), .B(ori_ori_n40_), .Y(ori_ori_n429_));
  NOi21      o407(.An(ori_ori_n90_), .B(ori_ori_n370_), .Y(ori_ori_n430_));
  INV        o408(.A(ori_ori_n430_), .Y(ori_ori_n431_));
  AOI210     o409(.A0(ori_ori_n431_), .A1(ori_ori_n429_), .B0(ori_ori_n47_), .Y(ori_ori_n432_));
  NO4        o410(.A(ori_ori_n196_), .B(ori_ori_n201_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n139_), .B(i_10_), .Y(ori_ori_n434_));
  NOi21      o412(.An(ori_ori_n434_), .B(ori_ori_n433_), .Y(ori_ori_n435_));
  NO2        o413(.A(ori_ori_n435_), .B(ori_ori_n56_), .Y(ori_ori_n436_));
  NOi21      o414(.An(i_5_), .B(i_9_), .Y(ori_ori_n437_));
  NA2        o415(.A(ori_ori_n437_), .B(ori_ori_n213_), .Y(ori_ori_n438_));
  BUFFER     o416(.A(ori_ori_n173_), .Y(ori_ori_n439_));
  NA2        o417(.A(ori_ori_n439_), .B(ori_ori_n230_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n440_), .B(ori_ori_n438_), .Y(ori_ori_n441_));
  NO3        o419(.A(ori_ori_n441_), .B(ori_ori_n436_), .C(ori_ori_n432_), .Y(ori_ori_n442_));
  NA2        o420(.A(ori_ori_n254_), .B(i_0_), .Y(ori_ori_n443_));
  NA2        o421(.A(ori_ori_n357_), .B(ori_ori_n184_), .Y(ori_ori_n444_));
  INV        o422(.A(ori_ori_n54_), .Y(ori_ori_n445_));
  NO2        o423(.A(ori_ori_n445_), .B(ori_ori_n444_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n164_), .B(ori_ori_n129_), .Y(ori_ori_n447_));
  NA2        o425(.A(i_0_), .B(i_10_), .Y(ori_ori_n448_));
  AN2        o426(.A(ori_ori_n447_), .B(i_6_), .Y(ori_ori_n449_));
  NO2        o427(.A(ori_ori_n449_), .B(ori_ori_n446_), .Y(ori_ori_n450_));
  INV        o428(.A(ori_ori_n450_), .Y(ori_ori_n451_));
  NA2        o429(.A(i_11_), .B(i_9_), .Y(ori_ori_n452_));
  NO3        o430(.A(i_12_), .B(ori_ori_n452_), .C(ori_ori_n265_), .Y(ori_ori_n453_));
  AN2        o431(.A(ori_ori_n453_), .B(i_5_), .Y(ori_ori_n454_));
  NA2        o432(.A(ori_ori_n204_), .B(ori_ori_n138_), .Y(ori_ori_n455_));
  NA2        o433(.A(ori_ori_n455_), .B(ori_ori_n133_), .Y(ori_ori_n456_));
  NO2        o434(.A(ori_ori_n452_), .B(ori_ori_n66_), .Y(ori_ori_n457_));
  NO2        o435(.A(ori_ori_n456_), .B(ori_ori_n454_), .Y(ori_ori_n458_));
  NA2        o436(.A(ori_ori_n298_), .B(ori_ori_n107_), .Y(ori_ori_n459_));
  NO2        o437(.A(i_6_), .B(ori_ori_n459_), .Y(ori_ori_n460_));
  NA2        o438(.A(ori_ori_n136_), .B(ori_ori_n95_), .Y(ori_ori_n461_));
  INV        o439(.A(ori_ori_n460_), .Y(ori_ori_n462_));
  NA2        o440(.A(ori_ori_n462_), .B(ori_ori_n458_), .Y(ori_ori_n463_));
  NO2        o441(.A(ori_ori_n426_), .B(ori_ori_n182_), .Y(ori_ori_n464_));
  NA2        o442(.A(ori_ori_n464_), .B(ori_ori_n457_), .Y(ori_ori_n465_));
  NA2        o443(.A(ori_ori_n244_), .B(ori_ori_n465_), .Y(ori_ori_n466_));
  NO3        o444(.A(ori_ori_n466_), .B(ori_ori_n463_), .C(ori_ori_n451_), .Y(ori_ori_n467_));
  NO2        o445(.A(ori_ori_n399_), .B(ori_ori_n461_), .Y(ori_ori_n468_));
  INV        o446(.A(ori_ori_n468_), .Y(ori_ori_n469_));
  NA2        o447(.A(ori_ori_n159_), .B(ori_ori_n152_), .Y(ori_ori_n470_));
  AOI210     o448(.A0(ori_ori_n470_), .A1(ori_ori_n443_), .B0(ori_ori_n129_), .Y(ori_ori_n471_));
  INV        o449(.A(ori_ori_n471_), .Y(ori_ori_n472_));
  NA2        o450(.A(ori_ori_n472_), .B(ori_ori_n469_), .Y(ori_ori_n473_));
  NO3        o451(.A(ori_ori_n448_), .B(ori_ori_n437_), .C(ori_ori_n141_), .Y(ori_ori_n474_));
  AOI220     o452(.A0(ori_ori_n474_), .A1(i_11_), .B0(ori_ori_n253_), .B1(ori_ori_n68_), .Y(ori_ori_n475_));
  NO3        o453(.A(ori_ori_n148_), .B(ori_ori_n201_), .C(i_0_), .Y(ori_ori_n476_));
  OAI210     o454(.A0(ori_ori_n476_), .A1(ori_ori_n69_), .B0(i_13_), .Y(ori_ori_n477_));
  NA2        o455(.A(ori_ori_n477_), .B(ori_ori_n475_), .Y(ori_ori_n478_));
  NA2        o456(.A(ori_ori_n239_), .B(ori_ori_n232_), .Y(ori_ori_n479_));
  INV        o457(.A(ori_ori_n479_), .Y(ori_ori_n480_));
  NA3        o458(.A(ori_ori_n203_), .B(ori_ori_n136_), .C(ori_ori_n135_), .Y(ori_ori_n481_));
  INV        o459(.A(ori_ori_n481_), .Y(ori_ori_n482_));
  NO3        o460(.A(ori_ori_n452_), .B(ori_ori_n149_), .C(ori_ori_n141_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n483_), .B(ori_ori_n482_), .Y(ori_ori_n484_));
  NA2        o462(.A(ori_ori_n484_), .B(ori_ori_n480_), .Y(ori_ori_n485_));
  NO2        o463(.A(ori_ori_n79_), .B(i_5_), .Y(ori_ori_n486_));
  NA3        o464(.A(ori_ori_n427_), .B(ori_ori_n101_), .C(ori_ori_n110_), .Y(ori_ori_n487_));
  INV        o465(.A(ori_ori_n487_), .Y(ori_ori_n488_));
  NA2        o466(.A(ori_ori_n488_), .B(ori_ori_n486_), .Y(ori_ori_n489_));
  NAi21      o467(.An(ori_ori_n157_), .B(ori_ori_n158_), .Y(ori_ori_n490_));
  NO4        o468(.A(ori_ori_n156_), .B(ori_ori_n148_), .C(i_0_), .D(i_12_), .Y(ori_ori_n491_));
  NA2        o469(.A(ori_ori_n491_), .B(ori_ori_n490_), .Y(ori_ori_n492_));
  NA2        o470(.A(ori_ori_n492_), .B(ori_ori_n489_), .Y(ori_ori_n493_));
  NO4        o471(.A(ori_ori_n493_), .B(ori_ori_n485_), .C(ori_ori_n478_), .D(ori_ori_n473_), .Y(ori_ori_n494_));
  INV        o472(.A(ori_ori_n273_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n495_), .B(ori_ori_n146_), .Y(ori_ori_n496_));
  NO2        o474(.A(ori_ori_n496_), .B(ori_ori_n66_), .Y(ori_ori_n497_));
  INV        o475(.A(ori_ori_n198_), .Y(ori_ori_n498_));
  NO2        o476(.A(ori_ori_n498_), .B(ori_ori_n365_), .Y(ori_ori_n499_));
  NO2        o477(.A(ori_ori_n499_), .B(ori_ori_n497_), .Y(ori_ori_n500_));
  NA4        o478(.A(ori_ori_n500_), .B(ori_ori_n494_), .C(ori_ori_n467_), .D(ori_ori_n442_), .Y(ori4));
  INV        o479(.A(i_6_), .Y(ori_ori_n504_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NO2        m028(.A(mai_mai_n47_), .B(mai_mai_n46_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_0_), .B(i_2_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_7_), .B(i_9_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  NA2        m032(.A(mai_mai_n51_), .B(mai_mai_n45_), .Y(mai_mai_n55_));
  NA3        m033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n56_));
  NO2        m034(.A(i_1_), .B(i_6_), .Y(mai_mai_n57_));
  NA2        m035(.A(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  OAI210     m036(.A0(mai_mai_n58_), .A1(mai_mai_n57_), .B0(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n60_));
  NAi21      m038(.An(i_2_), .B(i_7_), .Y(mai_mai_n61_));
  INV        m039(.A(i_1_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n62_), .B(i_6_), .Y(mai_mai_n63_));
  NA3        m041(.A(mai_mai_n63_), .B(mai_mai_n61_), .C(mai_mai_n31_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n60_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n67_));
  NA2        m045(.A(i_1_), .B(i_6_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n25_), .Y(mai_mai_n69_));
  INV        m047(.A(i_0_), .Y(mai_mai_n70_));
  NAi21      m048(.An(i_5_), .B(i_10_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_5_), .B(i_9_), .Y(mai_mai_n72_));
  AOI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n71_), .B0(mai_mai_n70_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n69_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n74_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n65_), .B0(i_0_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_12_), .B(i_5_), .Y(mai_mai_n77_));
  NO2        m055(.A(i_3_), .B(i_9_), .Y(mai_mai_n78_));
  NO2        m056(.A(i_3_), .B(i_7_), .Y(mai_mai_n79_));
  INV        m057(.A(i_6_), .Y(mai_mai_n80_));
  OR4        m058(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n81_));
  INV        m059(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m060(.A(i_2_), .B(i_7_), .Y(mai_mai_n83_));
  NAi21      m061(.An(i_6_), .B(i_10_), .Y(mai_mai_n84_));
  NA2        m062(.A(i_6_), .B(i_9_), .Y(mai_mai_n85_));
  AOI210     m063(.A0(mai_mai_n85_), .A1(mai_mai_n84_), .B0(mai_mai_n62_), .Y(mai_mai_n86_));
  NA2        m064(.A(i_2_), .B(i_6_), .Y(mai_mai_n87_));
  INV        m065(.A(mai_mai_n86_), .Y(mai_mai_n88_));
  NO2        m066(.A(mai_mai_n88_), .B(mai_mai_n77_), .Y(mai_mai_n89_));
  AN3        m067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n90_));
  NAi21      m068(.An(i_6_), .B(i_11_), .Y(mai_mai_n91_));
  NO2        m069(.A(i_5_), .B(i_8_), .Y(mai_mai_n92_));
  NOi21      m070(.An(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n93_));
  AOI220     m071(.A0(mai_mai_n93_), .A1(mai_mai_n61_), .B0(mai_mai_n90_), .B1(mai_mai_n32_), .Y(mai_mai_n94_));
  INV        m072(.A(i_7_), .Y(mai_mai_n95_));
  NA2        m073(.A(mai_mai_n46_), .B(mai_mai_n95_), .Y(mai_mai_n96_));
  NO2        m074(.A(i_0_), .B(i_5_), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n97_), .B(mai_mai_n80_), .Y(mai_mai_n98_));
  NA2        m076(.A(i_12_), .B(i_3_), .Y(mai_mai_n99_));
  INV        m077(.A(mai_mai_n99_), .Y(mai_mai_n100_));
  NA3        m078(.A(mai_mai_n100_), .B(mai_mai_n98_), .C(mai_mai_n96_), .Y(mai_mai_n101_));
  NAi21      m079(.An(i_7_), .B(i_11_), .Y(mai_mai_n102_));
  NO3        m080(.A(mai_mai_n102_), .B(mai_mai_n84_), .C(mai_mai_n52_), .Y(mai_mai_n103_));
  AN2        m081(.A(i_2_), .B(i_10_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n104_), .B(i_7_), .Y(mai_mai_n105_));
  OR2        m083(.A(mai_mai_n77_), .B(mai_mai_n57_), .Y(mai_mai_n106_));
  NO2        m084(.A(i_8_), .B(mai_mai_n95_), .Y(mai_mai_n107_));
  NO3        m085(.A(mai_mai_n107_), .B(mai_mai_n106_), .C(mai_mai_n105_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_12_), .B(i_7_), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n62_), .B(mai_mai_n26_), .Y(mai_mai_n110_));
  NA2        m088(.A(mai_mai_n110_), .B(i_0_), .Y(mai_mai_n111_));
  NA2        m089(.A(i_11_), .B(i_12_), .Y(mai_mai_n112_));
  OAI210     m090(.A0(mai_mai_n111_), .A1(mai_mai_n109_), .B0(mai_mai_n112_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n113_), .B(mai_mai_n108_), .Y(mai_mai_n114_));
  NAi41      m092(.An(mai_mai_n103_), .B(mai_mai_n114_), .C(mai_mai_n101_), .D(mai_mai_n94_), .Y(mai_mai_n115_));
  NOi21      m093(.An(i_1_), .B(i_5_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(i_11_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n95_), .B(mai_mai_n37_), .Y(mai_mai_n118_));
  NA2        m096(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(mai_mai_n46_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n122_));
  NAi21      m100(.An(i_3_), .B(i_8_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(mai_mai_n61_), .Y(mai_mai_n124_));
  NOi21      m102(.An(mai_mai_n124_), .B(mai_mai_n122_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_1_), .B(mai_mai_n80_), .Y(mai_mai_n126_));
  NO2        m104(.A(i_6_), .B(i_5_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(i_3_), .Y(mai_mai_n128_));
  AO210      m106(.A0(mai_mai_n128_), .A1(mai_mai_n47_), .B0(mai_mai_n126_), .Y(mai_mai_n129_));
  OAI220     m107(.A0(mai_mai_n129_), .A1(mai_mai_n102_), .B0(mai_mai_n125_), .B1(mai_mai_n117_), .Y(mai_mai_n130_));
  NO3        m108(.A(mai_mai_n130_), .B(mai_mai_n115_), .C(mai_mai_n89_), .Y(mai_mai_n131_));
  NA3        m109(.A(mai_mai_n131_), .B(mai_mai_n76_), .C(mai_mai_n55_), .Y(mai2));
  NO2        m110(.A(mai_mai_n62_), .B(mai_mai_n37_), .Y(mai_mai_n133_));
  NA2        m111(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .Y(mai_mai_n135_));
  NA4        m113(.A(mai_mai_n135_), .B(mai_mai_n74_), .C(mai_mai_n66_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m114(.A(i_8_), .B(i_7_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n137_), .B(i_6_), .Y(mai_mai_n138_));
  NO2        m116(.A(i_12_), .B(i_13_), .Y(mai_mai_n139_));
  NAi21      m117(.An(i_5_), .B(i_11_), .Y(mai_mai_n140_));
  NOi21      m118(.An(mai_mai_n139_), .B(mai_mai_n140_), .Y(mai_mai_n141_));
  NO2        m119(.A(i_0_), .B(i_1_), .Y(mai_mai_n142_));
  NA2        m120(.A(i_2_), .B(i_3_), .Y(mai_mai_n143_));
  NO2        m121(.A(mai_mai_n143_), .B(i_4_), .Y(mai_mai_n144_));
  NA2        m122(.A(mai_mai_n144_), .B(mai_mai_n141_), .Y(mai_mai_n145_));
  AN2        m123(.A(mai_mai_n139_), .B(mai_mai_n78_), .Y(mai_mai_n146_));
  NA2        m124(.A(i_1_), .B(i_5_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n70_), .B(mai_mai_n46_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(i_13_), .Y(mai_mai_n150_));
  OR2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n77_), .C(i_13_), .Y(mai_mai_n152_));
  NAi32      m130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n153_));
  NAi21      m131(.An(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m132(.An(i_4_), .B(i_10_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NO2        m134(.A(i_3_), .B(i_5_), .Y(mai_mai_n157_));
  NO3        m135(.A(mai_mai_n70_), .B(i_2_), .C(i_1_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n154_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(mai_mai_n150_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(mai_mai_n161_), .A1(mai_mai_n145_), .B0(mai_mai_n138_), .Y(mai_mai_n162_));
  NA3        m140(.A(mai_mai_n70_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n163_));
  NOi21      m141(.An(i_4_), .B(i_9_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_11_), .B(i_13_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  BUFFER     m144(.A(mai_mai_n166_), .Y(mai_mai_n167_));
  NO2        m145(.A(i_4_), .B(i_5_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_12_), .B(i_11_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(i_13_), .Y(mai_mai_n170_));
  NA2        m148(.A(mai_mai_n170_), .B(mai_mai_n78_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n167_), .B0(mai_mai_n163_), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n70_), .B(mai_mai_n62_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n173_), .B(mai_mai_n46_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n175_));
  NAi31      m153(.An(mai_mai_n175_), .B(mai_mai_n146_), .C(i_11_), .Y(mai_mai_n176_));
  NA2        m154(.A(i_3_), .B(i_5_), .Y(mai_mai_n177_));
  BUFFER     m155(.A(mai_mai_n166_), .Y(mai_mai_n178_));
  AOI210     m156(.A0(mai_mai_n178_), .A1(mai_mai_n176_), .B0(mai_mai_n174_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n180_));
  NO2        m158(.A(i_13_), .B(i_10_), .Y(mai_mai_n181_));
  NA3        m159(.A(mai_mai_n181_), .B(mai_mai_n180_), .C(mai_mai_n44_), .Y(mai_mai_n182_));
  NO2        m160(.A(i_2_), .B(i_1_), .Y(mai_mai_n183_));
  NA2        m161(.A(mai_mai_n183_), .B(i_3_), .Y(mai_mai_n184_));
  NAi21      m162(.An(i_4_), .B(i_12_), .Y(mai_mai_n185_));
  NO3        m163(.A(mai_mai_n185_), .B(mai_mai_n184_), .C(mai_mai_n182_), .Y(mai_mai_n186_));
  NO3        m164(.A(mai_mai_n186_), .B(mai_mai_n179_), .C(mai_mai_n172_), .Y(mai_mai_n187_));
  INV        m165(.A(i_8_), .Y(mai_mai_n188_));
  NA2        m166(.A(i_8_), .B(i_6_), .Y(mai_mai_n189_));
  NO3        m167(.A(i_3_), .B(mai_mai_n80_), .C(mai_mai_n48_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n190_), .B(mai_mai_n107_), .Y(mai_mai_n191_));
  NO3        m169(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n192_));
  NA3        m170(.A(mai_mai_n192_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n193_));
  NO3        m171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n194_));
  OAI210     m172(.A0(mai_mai_n90_), .A1(i_12_), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  AOI210     m173(.A0(mai_mai_n195_), .A1(mai_mai_n193_), .B0(mai_mai_n191_), .Y(mai_mai_n196_));
  NO2        m174(.A(i_3_), .B(i_8_), .Y(mai_mai_n197_));
  NO3        m175(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n198_));
  NA3        m176(.A(mai_mai_n198_), .B(mai_mai_n197_), .C(mai_mai_n40_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n97_), .B(mai_mai_n57_), .Y(mai_mai_n200_));
  NO2        m178(.A(i_13_), .B(i_9_), .Y(mai_mai_n201_));
  NA3        m179(.A(mai_mai_n201_), .B(i_6_), .C(mai_mai_n188_), .Y(mai_mai_n202_));
  NAi21      m180(.An(i_12_), .B(i_3_), .Y(mai_mai_n203_));
  NO2        m181(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n204_));
  NO3        m182(.A(i_0_), .B(i_2_), .C(mai_mai_n62_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n205_), .B(i_10_), .Y(mai_mai_n206_));
  OAI220     m184(.A0(mai_mai_n206_), .A1(mai_mai_n202_), .B0(mai_mai_n57_), .B1(mai_mai_n199_), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n207_), .A1(i_7_), .B0(mai_mai_n196_), .Y(mai_mai_n208_));
  OAI220     m186(.A0(mai_mai_n208_), .A1(i_4_), .B0(mai_mai_n189_), .B1(mai_mai_n187_), .Y(mai_mai_n209_));
  NAi21      m187(.An(i_12_), .B(i_7_), .Y(mai_mai_n210_));
  NA3        m188(.A(i_13_), .B(mai_mai_n188_), .C(i_10_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n211_), .B(mai_mai_n210_), .Y(mai_mai_n212_));
  NA2        m190(.A(i_0_), .B(i_5_), .Y(mai_mai_n213_));
  OAI220     m191(.A0(mai_mai_n80_), .A1(mai_mai_n184_), .B0(mai_mai_n174_), .B1(mai_mai_n128_), .Y(mai_mai_n214_));
  NAi31      m192(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n46_), .B(mai_mai_n62_), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n218_));
  INV        m196(.A(i_13_), .Y(mai_mai_n219_));
  NO2        m197(.A(i_12_), .B(mai_mai_n219_), .Y(mai_mai_n220_));
  NA3        m198(.A(mai_mai_n220_), .B(mai_mai_n192_), .C(mai_mai_n190_), .Y(mai_mai_n221_));
  OAI210     m199(.A0(mai_mai_n218_), .A1(mai_mai_n215_), .B0(mai_mai_n221_), .Y(mai_mai_n222_));
  AOI220     m200(.A0(mai_mai_n222_), .A1(mai_mai_n137_), .B0(mai_mai_n214_), .B1(mai_mai_n212_), .Y(mai_mai_n223_));
  NO2        m201(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  OR2        m204(.A(i_8_), .B(i_7_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n227_), .B(mai_mai_n80_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n52_), .B(i_1_), .Y(mai_mai_n229_));
  INV        m207(.A(i_12_), .Y(mai_mai_n230_));
  NO3        m208(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n231_));
  NA2        m209(.A(i_2_), .B(i_1_), .Y(mai_mai_n232_));
  NO3        m210(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n233_));
  NAi21      m211(.An(i_4_), .B(i_3_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n234_), .B(mai_mai_n72_), .Y(mai_mai_n235_));
  NO2        m213(.A(i_0_), .B(i_6_), .Y(mai_mai_n236_));
  NOi41      m214(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n232_), .B(mai_mai_n177_), .Y(mai_mai_n239_));
  NAi21      m217(.An(mai_mai_n238_), .B(mai_mai_n239_), .Y(mai_mai_n240_));
  NO2        m218(.A(i_11_), .B(mai_mai_n219_), .Y(mai_mai_n241_));
  NOi21      m219(.An(i_1_), .B(i_6_), .Y(mai_mai_n242_));
  NAi21      m220(.An(i_3_), .B(i_7_), .Y(mai_mai_n243_));
  NO2        m221(.A(mai_mai_n48_), .B(mai_mai_n25_), .Y(mai_mai_n244_));
  NO2        m222(.A(i_12_), .B(i_3_), .Y(mai_mai_n245_));
  NA3        m223(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n246_));
  INV        m224(.A(mai_mai_n138_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n230_), .B(i_13_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n248_), .B(mai_mai_n72_), .Y(mai_mai_n249_));
  NA2        m227(.A(mai_mai_n249_), .B(mai_mai_n247_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n227_), .B(mai_mai_n37_), .Y(mai_mai_n251_));
  NA2        m229(.A(i_12_), .B(i_6_), .Y(mai_mai_n252_));
  OR2        m230(.A(i_13_), .B(i_9_), .Y(mai_mai_n253_));
  NO3        m231(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n48_), .Y(mai_mai_n254_));
  NO2        m232(.A(mai_mai_n234_), .B(i_2_), .Y(mai_mai_n255_));
  NA3        m233(.A(mai_mai_n255_), .B(mai_mai_n254_), .C(mai_mai_n44_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n241_), .B(i_9_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n62_), .A1(mai_mai_n257_), .B0(mai_mai_n256_), .Y(mai_mai_n258_));
  NO3        m236(.A(i_11_), .B(mai_mai_n219_), .C(mai_mai_n25_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n243_), .B(i_8_), .Y(mai_mai_n260_));
  NO2        m238(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n261_));
  NA3        m239(.A(mai_mai_n261_), .B(mai_mai_n260_), .C(mai_mai_n259_), .Y(mai_mai_n262_));
  NO3        m240(.A(mai_mai_n26_), .B(mai_mai_n80_), .C(i_5_), .Y(mai_mai_n263_));
  NA3        m241(.A(mai_mai_n263_), .B(mai_mai_n251_), .C(mai_mai_n220_), .Y(mai_mai_n264_));
  AOI210     m242(.A0(mai_mai_n264_), .A1(mai_mai_n262_), .B0(i_1_), .Y(mai_mai_n265_));
  AOI210     m243(.A0(mai_mai_n258_), .A1(mai_mai_n251_), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  NA4        m244(.A(mai_mai_n266_), .B(mai_mai_n250_), .C(mai_mai_n240_), .D(mai_mai_n223_), .Y(mai_mai_n267_));
  NO3        m245(.A(i_12_), .B(mai_mai_n219_), .C(mai_mai_n37_), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n268_), .Y(mai_mai_n269_));
  NA2        m247(.A(i_8_), .B(mai_mai_n95_), .Y(mai_mai_n270_));
  NO3        m248(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n271_));
  AOI220     m249(.A0(mai_mai_n271_), .A1(mai_mai_n190_), .B0(mai_mai_n157_), .B1(mai_mai_n229_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n272_), .B(mai_mai_n270_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n232_), .B(i_0_), .Y(mai_mai_n274_));
  AOI220     m252(.A0(mai_mai_n274_), .A1(i_8_), .B0(i_1_), .B1(mai_mai_n137_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n261_), .B(mai_mai_n26_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(mai_mai_n275_), .Y(mai_mai_n277_));
  NA2        m255(.A(i_0_), .B(i_1_), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n278_), .B(i_2_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n58_), .B(i_6_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n280_), .B(mai_mai_n279_), .Y(mai_mai_n281_));
  OAI210     m259(.A0(mai_mai_n159_), .A1(mai_mai_n138_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  NO3        m260(.A(mai_mai_n282_), .B(mai_mai_n277_), .C(mai_mai_n273_), .Y(mai_mai_n283_));
  NO2        m261(.A(i_3_), .B(i_10_), .Y(mai_mai_n284_));
  NA3        m262(.A(mai_mai_n284_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n285_));
  NO2        m263(.A(i_2_), .B(mai_mai_n95_), .Y(mai_mai_n286_));
  NA2        m264(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n287_));
  NO2        m265(.A(mai_mai_n287_), .B(i_8_), .Y(mai_mai_n288_));
  INV        m266(.A(mai_mai_n288_), .Y(mai_mai_n289_));
  AN2        m267(.A(i_3_), .B(i_10_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n290_), .B(mai_mai_n192_), .C(mai_mai_n170_), .Y(mai_mai_n291_));
  NO2        m269(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n292_));
  NO2        m270(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n293_));
  OR2        m271(.A(mai_mai_n289_), .B(mai_mai_n285_), .Y(mai_mai_n294_));
  OAI220     m272(.A0(mai_mai_n294_), .A1(i_6_), .B0(mai_mai_n283_), .B1(mai_mai_n269_), .Y(mai_mai_n295_));
  NO4        m273(.A(mai_mai_n295_), .B(mai_mai_n267_), .C(mai_mai_n209_), .D(mai_mai_n162_), .Y(mai_mai_n296_));
  NO3        m274(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n297_));
  NO2        m275(.A(mai_mai_n58_), .B(mai_mai_n80_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n274_), .B(mai_mai_n298_), .Y(mai_mai_n299_));
  NO3        m277(.A(i_6_), .B(mai_mai_n188_), .C(i_7_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n300_), .B(mai_mai_n192_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n301_), .B(mai_mai_n299_), .Y(mai_mai_n302_));
  NO2        m280(.A(i_2_), .B(i_3_), .Y(mai_mai_n303_));
  OR2        m281(.A(i_0_), .B(i_5_), .Y(mai_mai_n304_));
  NA3        m282(.A(mai_mai_n228_), .B(mai_mai_n303_), .C(i_1_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n274_), .B(mai_mai_n157_), .C(mai_mai_n107_), .Y(mai_mai_n306_));
  NAi21      m284(.An(i_8_), .B(i_7_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n307_), .B(i_6_), .Y(mai_mai_n308_));
  NO2        m286(.A(mai_mai_n151_), .B(mai_mai_n46_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n309_), .B(mai_mai_n308_), .Y(mai_mai_n310_));
  NA3        m288(.A(mai_mai_n310_), .B(mai_mai_n306_), .C(mai_mai_n305_), .Y(mai_mai_n311_));
  OAI210     m289(.A0(mai_mai_n311_), .A1(mai_mai_n302_), .B0(i_4_), .Y(mai_mai_n312_));
  NO2        m290(.A(i_12_), .B(i_10_), .Y(mai_mai_n313_));
  NOi21      m291(.An(i_5_), .B(i_0_), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n287_), .B(mai_mai_n123_), .Y(mai_mai_n315_));
  NA4        m293(.A(mai_mai_n79_), .B(mai_mai_n36_), .C(mai_mai_n80_), .D(i_8_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n315_), .B(mai_mai_n313_), .Y(mai_mai_n317_));
  NO2        m295(.A(i_6_), .B(i_8_), .Y(mai_mai_n318_));
  NOi21      m296(.An(i_0_), .B(i_2_), .Y(mai_mai_n319_));
  AN2        m297(.A(mai_mai_n319_), .B(mai_mai_n318_), .Y(mai_mai_n320_));
  NO2        m298(.A(i_1_), .B(i_7_), .Y(mai_mai_n321_));
  AO220      m299(.A0(mai_mai_n321_), .A1(mai_mai_n320_), .B0(mai_mai_n308_), .B1(mai_mai_n229_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n322_), .B(i_4_), .Y(mai_mai_n323_));
  NA3        m301(.A(mai_mai_n323_), .B(mai_mai_n317_), .C(mai_mai_n312_), .Y(mai_mai_n324_));
  NO3        m302(.A(mai_mai_n227_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n325_));
  NO3        m303(.A(mai_mai_n307_), .B(i_2_), .C(i_1_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n326_), .A1(mai_mai_n325_), .B0(i_6_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n242_), .B(mai_mai_n286_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n328_), .B(mai_mai_n327_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(i_3_), .Y(mai_mai_n330_));
  INV        m308(.A(mai_mai_n79_), .Y(mai_mai_n331_));
  INV        m309(.A(mai_mai_n278_), .Y(mai_mai_n332_));
  NA2        m310(.A(mai_mai_n332_), .B(mai_mai_n127_), .Y(mai_mai_n333_));
  AOI210     m311(.A0(mai_mai_n87_), .A1(mai_mai_n333_), .B0(mai_mai_n331_), .Y(mai_mai_n334_));
  INV        m312(.A(i_9_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n335_), .B(mai_mai_n200_), .Y(mai_mai_n336_));
  NO2        m314(.A(mai_mai_n336_), .B(mai_mai_n46_), .Y(mai_mai_n337_));
  NO3        m315(.A(mai_mai_n337_), .B(mai_mai_n334_), .C(mai_mai_n277_), .Y(mai_mai_n338_));
  AOI210     m316(.A0(mai_mai_n338_), .A1(mai_mai_n330_), .B0(mai_mai_n156_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n324_), .A1(mai_mai_n297_), .B0(mai_mai_n339_), .Y(mai_mai_n340_));
  NOi32      m318(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n341_));
  INV        m319(.A(mai_mai_n341_), .Y(mai_mai_n342_));
  NAi21      m320(.An(i_0_), .B(i_6_), .Y(mai_mai_n343_));
  NAi21      m321(.An(i_1_), .B(i_5_), .Y(mai_mai_n344_));
  NA2        m322(.A(mai_mai_n344_), .B(mai_mai_n343_), .Y(mai_mai_n345_));
  NA2        m323(.A(mai_mai_n345_), .B(mai_mai_n25_), .Y(mai_mai_n346_));
  OAI210     m324(.A0(mai_mai_n346_), .A1(mai_mai_n153_), .B0(mai_mai_n238_), .Y(mai_mai_n347_));
  NAi41      m325(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n348_));
  OAI220     m326(.A0(mai_mai_n348_), .A1(mai_mai_n344_), .B0(mai_mai_n215_), .B1(mai_mai_n153_), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n348_), .A1(mai_mai_n153_), .B0(mai_mai_n151_), .Y(mai_mai_n350_));
  NOi32      m328(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n351_));
  NAi21      m329(.An(i_6_), .B(i_1_), .Y(mai_mai_n352_));
  NA3        m330(.A(mai_mai_n352_), .B(mai_mai_n351_), .C(mai_mai_n46_), .Y(mai_mai_n353_));
  NO2        m331(.A(mai_mai_n353_), .B(i_0_), .Y(mai_mai_n354_));
  OR3        m332(.A(mai_mai_n354_), .B(mai_mai_n350_), .C(mai_mai_n349_), .Y(mai_mai_n355_));
  NO2        m333(.A(i_1_), .B(mai_mai_n95_), .Y(mai_mai_n356_));
  NAi21      m334(.An(i_3_), .B(i_4_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n357_), .B(i_9_), .Y(mai_mai_n358_));
  AN2        m336(.A(i_6_), .B(i_7_), .Y(mai_mai_n359_));
  NA2        m337(.A(i_2_), .B(i_7_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n357_), .B(i_10_), .Y(mai_mai_n361_));
  NA3        m339(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n236_), .Y(mai_mai_n362_));
  INV        m340(.A(mai_mai_n362_), .Y(mai_mai_n363_));
  AOI210     m341(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n364_));
  AOI220     m342(.A0(mai_mai_n361_), .A1(mai_mai_n321_), .B0(mai_mai_n231_), .B1(mai_mai_n183_), .Y(mai_mai_n365_));
  NO2        m343(.A(mai_mai_n365_), .B(i_5_), .Y(mai_mai_n366_));
  NO4        m344(.A(mai_mai_n366_), .B(mai_mai_n363_), .C(mai_mai_n355_), .D(mai_mai_n347_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n367_), .B(mai_mai_n342_), .Y(mai_mai_n368_));
  NO2        m346(.A(mai_mai_n58_), .B(mai_mai_n25_), .Y(mai_mai_n369_));
  AN2        m347(.A(i_12_), .B(i_5_), .Y(mai_mai_n370_));
  NA2        m348(.A(i_3_), .B(mai_mai_n370_), .Y(mai_mai_n371_));
  NO2        m349(.A(i_11_), .B(i_6_), .Y(mai_mai_n372_));
  NA3        m350(.A(mai_mai_n372_), .B(mai_mai_n309_), .C(mai_mai_n219_), .Y(mai_mai_n373_));
  NO2        m351(.A(mai_mai_n373_), .B(mai_mai_n371_), .Y(mai_mai_n374_));
  NO2        m352(.A(mai_mai_n234_), .B(i_5_), .Y(mai_mai_n375_));
  NO2        m353(.A(i_5_), .B(i_10_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n139_), .B(mai_mai_n45_), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n377_), .B(mai_mai_n234_), .Y(mai_mai_n378_));
  OAI210     m356(.A0(mai_mai_n378_), .A1(mai_mai_n374_), .B0(mai_mai_n369_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n380_));
  NA2        m358(.A(mai_mai_n374_), .B(mai_mai_n380_), .Y(mai_mai_n381_));
  NO3        m359(.A(mai_mai_n80_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n382_));
  INV        m360(.A(mai_mai_n284_), .Y(mai_mai_n383_));
  NO2        m361(.A(i_11_), .B(i_12_), .Y(mai_mai_n384_));
  NA2        m362(.A(mai_mai_n384_), .B(mai_mai_n36_), .Y(mai_mai_n385_));
  NO2        m363(.A(mai_mai_n383_), .B(mai_mai_n385_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n376_), .B(mai_mai_n230_), .Y(mai_mai_n387_));
  NA2        m365(.A(i_4_), .B(i_11_), .Y(mai_mai_n388_));
  NO2        m366(.A(mai_mai_n388_), .B(mai_mai_n215_), .Y(mai_mai_n389_));
  NAi21      m367(.An(i_13_), .B(i_0_), .Y(mai_mai_n390_));
  NO2        m368(.A(mai_mai_n390_), .B(mai_mai_n232_), .Y(mai_mai_n391_));
  OAI210     m369(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n391_), .Y(mai_mai_n392_));
  NA3        m370(.A(mai_mai_n392_), .B(mai_mai_n381_), .C(mai_mai_n379_), .Y(mai_mai_n393_));
  NO3        m371(.A(i_1_), .B(i_12_), .C(mai_mai_n80_), .Y(mai_mai_n394_));
  NO2        m372(.A(i_0_), .B(i_11_), .Y(mai_mai_n395_));
  AN2        m373(.A(i_1_), .B(i_6_), .Y(mai_mai_n396_));
  NOi21      m374(.An(i_2_), .B(i_12_), .Y(mai_mai_n397_));
  NA2        m375(.A(mai_mai_n397_), .B(mai_mai_n396_), .Y(mai_mai_n398_));
  INV        m376(.A(mai_mai_n398_), .Y(mai_mai_n399_));
  NA2        m377(.A(mai_mai_n137_), .B(i_9_), .Y(mai_mai_n400_));
  NO2        m378(.A(mai_mai_n400_), .B(i_4_), .Y(mai_mai_n401_));
  NA2        m379(.A(mai_mai_n399_), .B(mai_mai_n401_), .Y(mai_mai_n402_));
  OR2        m380(.A(i_13_), .B(i_10_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n166_), .B(mai_mai_n118_), .Y(mai_mai_n404_));
  BUFFER     m382(.A(mai_mai_n211_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n95_), .B(mai_mai_n25_), .Y(mai_mai_n406_));
  NA2        m384(.A(mai_mai_n268_), .B(mai_mai_n406_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n261_), .B(mai_mai_n205_), .Y(mai_mai_n408_));
  OAI220     m386(.A0(mai_mai_n408_), .A1(mai_mai_n405_), .B0(mai_mai_n407_), .B1(mai_mai_n97_), .Y(mai_mai_n409_));
  INV        m387(.A(mai_mai_n409_), .Y(mai_mai_n410_));
  AOI210     m388(.A0(mai_mai_n410_), .A1(mai_mai_n402_), .B0(mai_mai_n26_), .Y(mai_mai_n411_));
  NA2        m389(.A(mai_mai_n306_), .B(mai_mai_n305_), .Y(mai_mai_n412_));
  AOI220     m390(.A0(mai_mai_n280_), .A1(mai_mai_n271_), .B0(mai_mai_n274_), .B1(mai_mai_n298_), .Y(mai_mai_n413_));
  NO2        m391(.A(mai_mai_n413_), .B(i_5_), .Y(mai_mai_n414_));
  NO2        m392(.A(mai_mai_n177_), .B(mai_mai_n80_), .Y(mai_mai_n415_));
  AOI220     m393(.A0(mai_mai_n415_), .A1(mai_mai_n279_), .B0(mai_mai_n263_), .B1(mai_mai_n205_), .Y(mai_mai_n416_));
  NO2        m394(.A(mai_mai_n416_), .B(mai_mai_n270_), .Y(mai_mai_n417_));
  NO3        m395(.A(mai_mai_n417_), .B(mai_mai_n414_), .C(mai_mai_n412_), .Y(mai_mai_n418_));
  NA2        m396(.A(mai_mai_n190_), .B(mai_mai_n90_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n309_), .B(mai_mai_n80_), .Y(mai_mai_n420_));
  AOI210     m398(.A0(mai_mai_n420_), .A1(mai_mai_n419_), .B0(mai_mai_n307_), .Y(mai_mai_n421_));
  NA2        m399(.A(mai_mai_n188_), .B(i_10_), .Y(mai_mai_n422_));
  NA2        m400(.A(mai_mai_n63_), .B(i_2_), .Y(mai_mai_n423_));
  NA2        m401(.A(mai_mai_n280_), .B(mai_mai_n229_), .Y(mai_mai_n424_));
  OAI220     m402(.A0(mai_mai_n424_), .A1(mai_mai_n177_), .B0(mai_mai_n423_), .B1(mai_mai_n422_), .Y(mai_mai_n425_));
  NA3        m403(.A(mai_mai_n321_), .B(mai_mai_n320_), .C(i_5_), .Y(mai_mai_n426_));
  INV        m404(.A(mai_mai_n300_), .Y(mai_mai_n427_));
  OAI210     m405(.A0(mai_mai_n427_), .A1(mai_mai_n184_), .B0(mai_mai_n426_), .Y(mai_mai_n428_));
  NO3        m406(.A(mai_mai_n428_), .B(mai_mai_n425_), .C(mai_mai_n421_), .Y(mai_mai_n429_));
  AOI210     m407(.A0(mai_mai_n429_), .A1(mai_mai_n418_), .B0(mai_mai_n257_), .Y(mai_mai_n430_));
  NO4        m408(.A(mai_mai_n430_), .B(mai_mai_n411_), .C(mai_mai_n393_), .D(mai_mai_n368_), .Y(mai_mai_n431_));
  NO2        m409(.A(mai_mai_n70_), .B(i_13_), .Y(mai_mai_n432_));
  NO2        m410(.A(i_10_), .B(i_9_), .Y(mai_mai_n433_));
  NAi21      m411(.An(i_12_), .B(i_8_), .Y(mai_mai_n434_));
  NO2        m412(.A(mai_mai_n434_), .B(i_3_), .Y(mai_mai_n435_));
  NA2        m413(.A(i_2_), .B(mai_mai_n98_), .Y(mai_mai_n436_));
  NO2        m414(.A(mai_mai_n436_), .B(mai_mai_n199_), .Y(mai_mai_n437_));
  NA2        m415(.A(mai_mai_n293_), .B(i_0_), .Y(mai_mai_n438_));
  NO3        m416(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n439_));
  NA2        m417(.A(mai_mai_n252_), .B(mai_mai_n91_), .Y(mai_mai_n440_));
  NA2        m418(.A(mai_mai_n440_), .B(mai_mai_n439_), .Y(mai_mai_n441_));
  NA2        m419(.A(i_8_), .B(i_9_), .Y(mai_mai_n442_));
  NO3        m420(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n443_));
  NA3        m421(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n444_));
  NA4        m422(.A(mai_mai_n140_), .B(mai_mai_n110_), .C(mai_mai_n77_), .D(mai_mai_n23_), .Y(mai_mai_n445_));
  NO2        m423(.A(mai_mai_n445_), .B(mai_mai_n444_), .Y(mai_mai_n446_));
  NO2        m424(.A(mai_mai_n446_), .B(mai_mai_n437_), .Y(mai_mai_n447_));
  OA210      m425(.A0(mai_mai_n336_), .A1(mai_mai_n95_), .B0(mai_mai_n281_), .Y(mai_mai_n448_));
  OA220      m426(.A0(mai_mai_n448_), .A1(mai_mai_n156_), .B0(mai_mai_n202_), .B1(mai_mai_n226_), .Y(mai_mai_n449_));
  NA2        m427(.A(mai_mai_n90_), .B(i_13_), .Y(mai_mai_n450_));
  NA2        m428(.A(mai_mai_n415_), .B(mai_mai_n369_), .Y(mai_mai_n451_));
  NO2        m429(.A(i_2_), .B(i_13_), .Y(mai_mai_n452_));
  NO2        m430(.A(mai_mai_n451_), .B(mai_mai_n450_), .Y(mai_mai_n453_));
  NO3        m431(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n454_));
  NO2        m432(.A(i_6_), .B(i_7_), .Y(mai_mai_n455_));
  NA2        m433(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n456_));
  NO2        m434(.A(i_11_), .B(i_1_), .Y(mai_mai_n457_));
  OR2        m435(.A(i_11_), .B(i_8_), .Y(mai_mai_n458_));
  NOi21      m436(.An(i_2_), .B(i_7_), .Y(mai_mai_n459_));
  NAi31      m437(.An(mai_mai_n458_), .B(mai_mai_n459_), .C(i_0_), .Y(mai_mai_n460_));
  NO2        m438(.A(mai_mai_n403_), .B(i_6_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n461_), .B(i_1_), .Y(mai_mai_n462_));
  NO2        m440(.A(mai_mai_n462_), .B(mai_mai_n460_), .Y(mai_mai_n463_));
  NO2        m441(.A(i_3_), .B(mai_mai_n188_), .Y(mai_mai_n464_));
  NO2        m442(.A(i_6_), .B(i_10_), .Y(mai_mai_n465_));
  NA3        m443(.A(mai_mai_n465_), .B(mai_mai_n297_), .C(mai_mai_n464_), .Y(mai_mai_n466_));
  NO2        m444(.A(mai_mai_n466_), .B(mai_mai_n149_), .Y(mai_mai_n467_));
  NA2        m445(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n468_));
  NO2        m446(.A(mai_mai_n151_), .B(i_3_), .Y(mai_mai_n469_));
  NO3        m447(.A(mai_mai_n467_), .B(mai_mai_n463_), .C(mai_mai_n453_), .Y(mai_mai_n470_));
  NAi21      m448(.An(mai_mai_n211_), .B(mai_mai_n384_), .Y(mai_mai_n471_));
  NA2        m449(.A(mai_mai_n321_), .B(mai_mai_n213_), .Y(mai_mai_n472_));
  NO2        m450(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n473_));
  NA3        m451(.A(i_6_), .B(mai_mai_n473_), .C(mai_mai_n137_), .Y(mai_mai_n474_));
  OR3        m452(.A(mai_mai_n287_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n475_));
  OAI220     m453(.A0(mai_mai_n475_), .A1(mai_mai_n474_), .B0(mai_mai_n472_), .B1(mai_mai_n471_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n477_));
  NA2        m455(.A(mai_mai_n297_), .B(mai_mai_n231_), .Y(mai_mai_n478_));
  OAI220     m456(.A0(mai_mai_n478_), .A1(mai_mai_n423_), .B0(mai_mai_n477_), .B1(mai_mai_n450_), .Y(mai_mai_n479_));
  NA3        m457(.A(mai_mai_n290_), .B(mai_mai_n217_), .C(mai_mai_n70_), .Y(mai_mai_n480_));
  NO2        m458(.A(mai_mai_n480_), .B(mai_mai_n456_), .Y(mai_mai_n481_));
  NO3        m459(.A(mai_mai_n481_), .B(mai_mai_n479_), .C(mai_mai_n476_), .Y(mai_mai_n482_));
  NA4        m460(.A(mai_mai_n482_), .B(mai_mai_n470_), .C(mai_mai_n449_), .D(mai_mai_n447_), .Y(mai_mai_n483_));
  NA3        m461(.A(mai_mai_n290_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n484_));
  INV        m462(.A(mai_mai_n484_), .Y(mai_mai_n485_));
  BUFFER     m463(.A(mai_mai_n271_), .Y(mai_mai_n486_));
  NA2        m464(.A(mai_mai_n486_), .B(mai_mai_n485_), .Y(mai_mai_n487_));
  AN2        m465(.A(i_11_), .B(mai_mai_n439_), .Y(mai_mai_n488_));
  INV        m466(.A(mai_mai_n158_), .Y(mai_mai_n489_));
  OAI210     m467(.A0(mai_mai_n489_), .A1(mai_mai_n226_), .B0(mai_mai_n291_), .Y(mai_mai_n490_));
  AOI220     m468(.A0(mai_mai_n490_), .A1(mai_mai_n308_), .B0(mai_mai_n488_), .B1(mai_mai_n293_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n341_), .B(mai_mai_n70_), .Y(mai_mai_n492_));
  INV        m470(.A(mai_mai_n351_), .Y(mai_mai_n493_));
  NO2        m471(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n494_));
  NAi41      m472(.An(mai_mai_n492_), .B(mai_mai_n465_), .C(mai_mai_n494_), .D(mai_mai_n46_), .Y(mai_mai_n495_));
  NA2        m473(.A(mai_mai_n39_), .B(i_13_), .Y(mai_mai_n496_));
  INV        m474(.A(mai_mai_n495_), .Y(mai_mai_n497_));
  NO2        m475(.A(i_7_), .B(mai_mai_n193_), .Y(mai_mai_n498_));
  OR2        m476(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n499_));
  INV        m477(.A(mai_mai_n499_), .Y(mai_mai_n500_));
  AOI220     m478(.A0(mai_mai_n500_), .A1(mai_mai_n498_), .B0(i_1_), .B1(mai_mai_n404_), .Y(mai_mai_n501_));
  NA4        m479(.A(mai_mai_n501_), .B(mai_mai_n496_), .C(mai_mai_n491_), .D(mai_mai_n487_), .Y(mai_mai_n502_));
  NA2        m480(.A(mai_mai_n375_), .B(mai_mai_n279_), .Y(mai_mai_n503_));
  NA2        m481(.A(mai_mai_n371_), .B(mai_mai_n503_), .Y(mai_mai_n504_));
  NO2        m482(.A(i_12_), .B(mai_mai_n188_), .Y(mai_mai_n505_));
  NA2        m483(.A(mai_mai_n505_), .B(mai_mai_n219_), .Y(mai_mai_n506_));
  NO2        m484(.A(i_10_), .B(mai_mai_n506_), .Y(mai_mai_n507_));
  NOi31      m485(.An(mai_mai_n300_), .B(mai_mai_n403_), .C(mai_mai_n38_), .Y(mai_mai_n508_));
  OAI210     m486(.A0(mai_mai_n508_), .A1(mai_mai_n507_), .B0(mai_mai_n504_), .Y(mai_mai_n509_));
  NO2        m487(.A(i_8_), .B(i_7_), .Y(mai_mai_n510_));
  OAI210     m488(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(mai_mai_n511_));
  NA2        m489(.A(mai_mai_n511_), .B(mai_mai_n217_), .Y(mai_mai_n512_));
  OAI220     m490(.A0(mai_mai_n46_), .A1(mai_mai_n499_), .B0(mai_mai_n512_), .B1(mai_mai_n234_), .Y(mai_mai_n513_));
  NA2        m491(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n514_));
  NO2        m492(.A(mai_mai_n514_), .B(i_6_), .Y(mai_mai_n515_));
  NA3        m493(.A(mai_mai_n515_), .B(mai_mai_n513_), .C(mai_mai_n510_), .Y(mai_mai_n516_));
  AOI220     m494(.A0(mai_mai_n415_), .A1(mai_mai_n309_), .B0(mai_mai_n239_), .B1(mai_mai_n236_), .Y(mai_mai_n517_));
  OAI220     m495(.A0(mai_mai_n517_), .A1(mai_mai_n248_), .B0(mai_mai_n450_), .B1(mai_mai_n128_), .Y(mai_mai_n518_));
  NA2        m496(.A(mai_mai_n518_), .B(mai_mai_n251_), .Y(mai_mai_n519_));
  NA3        m497(.A(mai_mai_n290_), .B(mai_mai_n168_), .C(mai_mai_n90_), .Y(mai_mai_n520_));
  NO2        m498(.A(mai_mai_n151_), .B(i_5_), .Y(mai_mai_n521_));
  NA2        m499(.A(mai_mai_n521_), .B(mai_mai_n303_), .Y(mai_mai_n522_));
  NA2        m500(.A(mai_mai_n522_), .B(mai_mai_n520_), .Y(mai_mai_n523_));
  NA2        m501(.A(mai_mai_n523_), .B(mai_mai_n443_), .Y(mai_mai_n524_));
  NA4        m502(.A(mai_mai_n524_), .B(mai_mai_n519_), .C(mai_mai_n516_), .D(mai_mai_n509_), .Y(mai_mai_n525_));
  NA2        m503(.A(mai_mai_n268_), .B(mai_mai_n79_), .Y(mai_mai_n526_));
  NO2        m504(.A(mai_mai_n333_), .B(mai_mai_n526_), .Y(mai_mai_n527_));
  NA2        m505(.A(mai_mai_n280_), .B(mai_mai_n271_), .Y(mai_mai_n528_));
  NO2        m506(.A(mai_mai_n528_), .B(mai_mai_n167_), .Y(mai_mai_n529_));
  NA2        m507(.A(mai_mai_n217_), .B(i_0_), .Y(mai_mai_n530_));
  NA2        m508(.A(mai_mai_n433_), .B(mai_mai_n216_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n530_), .B(mai_mai_n531_), .Y(mai_mai_n532_));
  AOI210     m510(.A0(mai_mai_n352_), .A1(mai_mai_n46_), .B0(mai_mai_n356_), .Y(mai_mai_n533_));
  NA2        m511(.A(i_0_), .B(mai_mai_n48_), .Y(mai_mai_n534_));
  NA3        m512(.A(mai_mai_n505_), .B(mai_mai_n259_), .C(mai_mai_n534_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n533_), .B(mai_mai_n535_), .Y(mai_mai_n536_));
  NO4        m514(.A(mai_mai_n536_), .B(mai_mai_n532_), .C(mai_mai_n529_), .D(mai_mai_n527_), .Y(mai_mai_n537_));
  NO4        m515(.A(mai_mai_n242_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n538_));
  NO3        m516(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n539_));
  NO2        m517(.A(mai_mai_n227_), .B(mai_mai_n36_), .Y(mai_mai_n540_));
  AN2        m518(.A(mai_mai_n540_), .B(mai_mai_n539_), .Y(mai_mai_n541_));
  OA210      m519(.A0(mai_mai_n541_), .A1(mai_mai_n538_), .B0(mai_mai_n341_), .Y(mai_mai_n542_));
  NO2        m520(.A(mai_mai_n403_), .B(i_1_), .Y(mai_mai_n543_));
  NOi31      m521(.An(mai_mai_n543_), .B(mai_mai_n440_), .C(mai_mai_n70_), .Y(mai_mai_n544_));
  AN3        m522(.A(mai_mai_n544_), .B(mai_mai_n401_), .C(mai_mai_n473_), .Y(mai_mai_n545_));
  NO2        m523(.A(mai_mai_n413_), .B(mai_mai_n171_), .Y(mai_mai_n546_));
  NO3        m524(.A(mai_mai_n546_), .B(mai_mai_n545_), .C(mai_mai_n542_), .Y(mai_mai_n547_));
  NOi21      m525(.An(i_10_), .B(i_6_), .Y(mai_mai_n548_));
  NO2        m526(.A(mai_mai_n80_), .B(mai_mai_n25_), .Y(mai_mai_n549_));
  AOI220     m527(.A0(mai_mai_n268_), .A1(mai_mai_n549_), .B0(mai_mai_n259_), .B1(mai_mai_n548_), .Y(mai_mai_n550_));
  NO2        m528(.A(mai_mai_n550_), .B(mai_mai_n438_), .Y(mai_mai_n551_));
  NO2        m529(.A(mai_mai_n109_), .B(mai_mai_n23_), .Y(mai_mai_n552_));
  NA2        m530(.A(mai_mai_n300_), .B(mai_mai_n158_), .Y(mai_mai_n553_));
  AOI220     m531(.A0(mai_mai_n553_), .A1(mai_mai_n424_), .B0(mai_mai_n178_), .B1(mai_mai_n176_), .Y(mai_mai_n554_));
  NOi21      m532(.An(mai_mai_n141_), .B(mai_mai_n316_), .Y(mai_mai_n555_));
  NO3        m533(.A(mai_mai_n555_), .B(mai_mai_n554_), .C(mai_mai_n551_), .Y(mai_mai_n556_));
  NO2        m534(.A(mai_mai_n492_), .B(mai_mai_n365_), .Y(mai_mai_n557_));
  INV        m535(.A(mai_mai_n303_), .Y(mai_mai_n558_));
  NO2        m536(.A(i_12_), .B(mai_mai_n80_), .Y(mai_mai_n559_));
  NA3        m537(.A(mai_mai_n559_), .B(mai_mai_n259_), .C(mai_mai_n534_), .Y(mai_mai_n560_));
  NA2        m538(.A(mai_mai_n372_), .B(mai_mai_n268_), .Y(mai_mai_n561_));
  AOI210     m539(.A0(mai_mai_n561_), .A1(mai_mai_n560_), .B0(mai_mai_n558_), .Y(mai_mai_n562_));
  NO3        m540(.A(i_4_), .B(mai_mai_n327_), .C(mai_mai_n285_), .Y(mai_mai_n563_));
  OR2        m541(.A(i_2_), .B(i_5_), .Y(mai_mai_n564_));
  OR2        m542(.A(mai_mai_n564_), .B(mai_mai_n396_), .Y(mai_mai_n565_));
  NA2        m543(.A(mai_mai_n360_), .B(mai_mai_n236_), .Y(mai_mai_n566_));
  AOI210     m544(.A0(mai_mai_n566_), .A1(mai_mai_n565_), .B0(mai_mai_n471_), .Y(mai_mai_n567_));
  NO4        m545(.A(mai_mai_n567_), .B(mai_mai_n563_), .C(mai_mai_n562_), .D(mai_mai_n557_), .Y(mai_mai_n568_));
  NA4        m546(.A(mai_mai_n568_), .B(mai_mai_n556_), .C(mai_mai_n547_), .D(mai_mai_n537_), .Y(mai_mai_n569_));
  NO4        m547(.A(mai_mai_n569_), .B(mai_mai_n525_), .C(mai_mai_n502_), .D(mai_mai_n483_), .Y(mai_mai_n570_));
  NA4        m548(.A(mai_mai_n570_), .B(mai_mai_n431_), .C(mai_mai_n340_), .D(mai_mai_n296_), .Y(mai7));
  NO2        m549(.A(mai_mai_n87_), .B(mai_mai_n53_), .Y(mai_mai_n572_));
  NO2        m550(.A(mai_mai_n102_), .B(mai_mai_n84_), .Y(mai_mai_n573_));
  NA2        m551(.A(i_3_), .B(mai_mai_n573_), .Y(mai_mai_n574_));
  NA2        m552(.A(mai_mai_n465_), .B(mai_mai_n79_), .Y(mai_mai_n575_));
  NA2        m553(.A(i_11_), .B(mai_mai_n188_), .Y(mai_mai_n576_));
  NA2        m554(.A(mai_mai_n139_), .B(mai_mai_n576_), .Y(mai_mai_n577_));
  OAI210     m555(.A0(mai_mai_n577_), .A1(mai_mai_n575_), .B0(mai_mai_n574_), .Y(mai_mai_n578_));
  NO2        m556(.A(mai_mai_n230_), .B(i_4_), .Y(mai_mai_n579_));
  NA2        m557(.A(mai_mai_n579_), .B(i_8_), .Y(mai_mai_n580_));
  NA2        m558(.A(i_2_), .B(mai_mai_n80_), .Y(mai_mai_n581_));
  OAI210     m559(.A0(mai_mai_n83_), .A1(mai_mai_n197_), .B0(mai_mai_n198_), .Y(mai_mai_n582_));
  NO2        m560(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n583_));
  NA2        m561(.A(i_4_), .B(i_8_), .Y(mai_mai_n584_));
  NO2        m562(.A(mai_mai_n578_), .B(mai_mai_n572_), .Y(mai_mai_n585_));
  INV        m563(.A(mai_mai_n155_), .Y(mai_mai_n586_));
  OR2        m564(.A(i_6_), .B(i_10_), .Y(mai_mai_n587_));
  NO2        m565(.A(mai_mai_n587_), .B(mai_mai_n23_), .Y(mai_mai_n588_));
  OR3        m566(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n589_));
  NO3        m567(.A(mai_mai_n589_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n590_));
  INV        m568(.A(mai_mai_n194_), .Y(mai_mai_n591_));
  NO2        m569(.A(mai_mai_n590_), .B(mai_mai_n588_), .Y(mai_mai_n592_));
  OA220      m570(.A0(mai_mai_n592_), .A1(mai_mai_n558_), .B0(mai_mai_n586_), .B1(mai_mai_n253_), .Y(mai_mai_n593_));
  AOI210     m571(.A0(mai_mai_n593_), .A1(mai_mai_n585_), .B0(mai_mai_n62_), .Y(mai_mai_n594_));
  NOi21      m572(.An(i_11_), .B(i_7_), .Y(mai_mai_n595_));
  AO210      m573(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n596_));
  NO2        m574(.A(mai_mai_n596_), .B(mai_mai_n595_), .Y(mai_mai_n597_));
  NA2        m575(.A(mai_mai_n597_), .B(mai_mai_n201_), .Y(mai_mai_n598_));
  NA3        m576(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n599_));
  NAi31      m577(.An(mai_mai_n599_), .B(mai_mai_n210_), .C(i_11_), .Y(mai_mai_n600_));
  AOI210     m578(.A0(mai_mai_n600_), .A1(mai_mai_n598_), .B0(mai_mai_n62_), .Y(mai_mai_n601_));
  NA2        m579(.A(mai_mai_n82_), .B(mai_mai_n62_), .Y(mai_mai_n602_));
  AO210      m580(.A0(mai_mai_n602_), .A1(mai_mai_n365_), .B0(mai_mai_n41_), .Y(mai_mai_n603_));
  NO3        m581(.A(i_7_), .B(mai_mai_n203_), .C(mai_mai_n576_), .Y(mai_mai_n604_));
  OAI210     m582(.A0(mai_mai_n604_), .A1(mai_mai_n220_), .B0(mai_mai_n62_), .Y(mai_mai_n605_));
  NA2        m583(.A(mai_mai_n397_), .B(mai_mai_n31_), .Y(mai_mai_n606_));
  OR2        m584(.A(mai_mai_n203_), .B(mai_mai_n102_), .Y(mai_mai_n607_));
  NA2        m585(.A(mai_mai_n607_), .B(mai_mai_n606_), .Y(mai_mai_n608_));
  NO2        m586(.A(mai_mai_n62_), .B(i_9_), .Y(mai_mai_n609_));
  NO2        m587(.A(mai_mai_n609_), .B(i_4_), .Y(mai_mai_n610_));
  NA2        m588(.A(mai_mai_n610_), .B(mai_mai_n608_), .Y(mai_mai_n611_));
  NO2        m589(.A(i_1_), .B(i_12_), .Y(mai_mai_n612_));
  NA3        m590(.A(mai_mai_n612_), .B(mai_mai_n104_), .C(mai_mai_n24_), .Y(mai_mai_n613_));
  NA4        m591(.A(mai_mai_n613_), .B(mai_mai_n611_), .C(mai_mai_n605_), .D(mai_mai_n603_), .Y(mai_mai_n614_));
  OAI210     m592(.A0(mai_mai_n614_), .A1(mai_mai_n601_), .B0(i_6_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n599_), .B(mai_mai_n102_), .Y(mai_mai_n616_));
  NA2        m594(.A(mai_mai_n616_), .B(mai_mai_n559_), .Y(mai_mai_n617_));
  NO2        m595(.A(i_6_), .B(i_11_), .Y(mai_mai_n618_));
  NA2        m596(.A(mai_mai_n617_), .B(mai_mai_n441_), .Y(mai_mai_n619_));
  NO4        m597(.A(mai_mai_n210_), .B(mai_mai_n123_), .C(i_13_), .D(mai_mai_n80_), .Y(mai_mai_n620_));
  NA2        m598(.A(mai_mai_n620_), .B(mai_mai_n609_), .Y(mai_mai_n621_));
  INV        m599(.A(mai_mai_n621_), .Y(mai_mai_n622_));
  NA3        m600(.A(mai_mai_n510_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n623_));
  NA2        m601(.A(mai_mai_n133_), .B(i_9_), .Y(mai_mai_n624_));
  NA3        m602(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n626_));
  NA3        m604(.A(mai_mai_n626_), .B(mai_mai_n252_), .C(mai_mai_n44_), .Y(mai_mai_n627_));
  OAI220     m605(.A0(mai_mai_n627_), .A1(mai_mai_n625_), .B0(mai_mai_n624_), .B1(mai_mai_n1003_), .Y(mai_mai_n628_));
  NA3        m606(.A(mai_mai_n609_), .B(mai_mai_n303_), .C(i_6_), .Y(mai_mai_n629_));
  NO2        m607(.A(mai_mai_n629_), .B(mai_mai_n23_), .Y(mai_mai_n630_));
  AOI210     m608(.A0(mai_mai_n457_), .A1(mai_mai_n406_), .B0(mai_mai_n233_), .Y(mai_mai_n631_));
  NO2        m609(.A(mai_mai_n631_), .B(mai_mai_n581_), .Y(mai_mai_n632_));
  NAi21      m610(.An(mai_mai_n623_), .B(mai_mai_n86_), .Y(mai_mai_n633_));
  NA2        m611(.A(mai_mai_n626_), .B(mai_mai_n252_), .Y(mai_mai_n634_));
  NO2        m612(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n635_));
  NA2        m613(.A(mai_mai_n635_), .B(mai_mai_n24_), .Y(mai_mai_n636_));
  OAI210     m614(.A0(mai_mai_n636_), .A1(mai_mai_n634_), .B0(mai_mai_n633_), .Y(mai_mai_n637_));
  OR4        m615(.A(mai_mai_n637_), .B(mai_mai_n632_), .C(mai_mai_n630_), .D(mai_mai_n628_), .Y(mai_mai_n638_));
  NO3        m616(.A(mai_mai_n638_), .B(mai_mai_n622_), .C(mai_mai_n619_), .Y(mai_mai_n639_));
  NO2        m617(.A(mai_mai_n230_), .B(mai_mai_n95_), .Y(mai_mai_n640_));
  NO2        m618(.A(mai_mai_n640_), .B(mai_mai_n595_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n641_), .B(i_1_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n642_), .B(mai_mai_n589_), .Y(mai_mai_n643_));
  NA2        m621(.A(mai_mai_n643_), .B(mai_mai_n46_), .Y(mai_mai_n644_));
  NA2        m622(.A(i_3_), .B(mai_mai_n188_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n645_), .B(mai_mai_n109_), .Y(mai_mai_n646_));
  AN2        m624(.A(mai_mai_n646_), .B(mai_mai_n515_), .Y(mai_mai_n647_));
  NO2        m625(.A(mai_mai_n112_), .B(mai_mai_n37_), .Y(mai_mai_n648_));
  NO2        m626(.A(mai_mai_n80_), .B(i_9_), .Y(mai_mai_n649_));
  NA2        m627(.A(i_1_), .B(i_3_), .Y(mai_mai_n650_));
  NO2        m628(.A(mai_mai_n442_), .B(mai_mai_n87_), .Y(mai_mai_n651_));
  INV        m629(.A(mai_mai_n651_), .Y(mai_mai_n652_));
  NO2        m630(.A(mai_mai_n652_), .B(mai_mai_n650_), .Y(mai_mai_n653_));
  NO2        m631(.A(mai_mai_n653_), .B(mai_mai_n647_), .Y(mai_mai_n654_));
  NA4        m632(.A(mai_mai_n654_), .B(mai_mai_n644_), .C(mai_mai_n639_), .D(mai_mai_n615_), .Y(mai_mai_n655_));
  NO3        m633(.A(mai_mai_n458_), .B(i_3_), .C(i_7_), .Y(mai_mai_n656_));
  NOi21      m634(.An(mai_mai_n656_), .B(i_10_), .Y(mai_mai_n657_));
  OA210      m635(.A0(mai_mai_n657_), .A1(mai_mai_n237_), .B0(mai_mai_n80_), .Y(mai_mai_n658_));
  NA2        m636(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n659_));
  NA3        m637(.A(mai_mai_n465_), .B(mai_mai_n494_), .C(mai_mai_n46_), .Y(mai_mai_n660_));
  NO3        m638(.A(mai_mai_n459_), .B(mai_mai_n584_), .C(mai_mai_n80_), .Y(mai_mai_n661_));
  NA2        m639(.A(mai_mai_n661_), .B(mai_mai_n25_), .Y(mai_mai_n662_));
  NA3        m640(.A(mai_mai_n155_), .B(mai_mai_n79_), .C(mai_mai_n80_), .Y(mai_mai_n663_));
  NA4        m641(.A(mai_mai_n663_), .B(mai_mai_n662_), .C(mai_mai_n660_), .D(mai_mai_n659_), .Y(mai_mai_n664_));
  OAI210     m642(.A0(mai_mai_n664_), .A1(mai_mai_n658_), .B0(i_1_), .Y(mai_mai_n665_));
  AOI210     m643(.A0(mai_mai_n252_), .A1(mai_mai_n91_), .B0(i_1_), .Y(mai_mai_n666_));
  NO2        m644(.A(mai_mai_n357_), .B(i_2_), .Y(mai_mai_n667_));
  NA2        m645(.A(mai_mai_n667_), .B(mai_mai_n666_), .Y(mai_mai_n668_));
  OAI210     m646(.A0(mai_mai_n629_), .A1(mai_mai_n434_), .B0(mai_mai_n668_), .Y(mai_mai_n669_));
  INV        m647(.A(mai_mai_n669_), .Y(mai_mai_n670_));
  AOI210     m648(.A0(mai_mai_n670_), .A1(mai_mai_n665_), .B0(i_13_), .Y(mai_mai_n671_));
  OR2        m649(.A(i_11_), .B(i_7_), .Y(mai_mai_n672_));
  NA3        m650(.A(mai_mai_n672_), .B(mai_mai_n100_), .C(mai_mai_n133_), .Y(mai_mai_n673_));
  AOI220     m651(.A0(mai_mai_n452_), .A1(mai_mai_n155_), .B0(i_2_), .B1(mai_mai_n133_), .Y(mai_mai_n674_));
  OAI210     m652(.A0(mai_mai_n674_), .A1(mai_mai_n44_), .B0(mai_mai_n673_), .Y(mai_mai_n675_));
  AOI210     m653(.A0(mai_mai_n625_), .A1(mai_mai_n53_), .B0(i_12_), .Y(mai_mai_n676_));
  NA2        m654(.A(mai_mai_n237_), .B(mai_mai_n126_), .Y(mai_mai_n677_));
  OAI220     m655(.A0(mai_mai_n677_), .A1(mai_mai_n41_), .B0(mai_mai_n1002_), .B1(mai_mai_n87_), .Y(mai_mai_n678_));
  AOI210     m656(.A0(mai_mai_n675_), .A1(mai_mai_n318_), .B0(mai_mai_n678_), .Y(mai_mai_n679_));
  AOI220     m657(.A0(i_12_), .A1(mai_mai_n69_), .B0(mai_mai_n372_), .B1(mai_mai_n626_), .Y(mai_mai_n680_));
  NO2        m658(.A(mai_mai_n680_), .B(mai_mai_n234_), .Y(mai_mai_n681_));
  AOI210     m659(.A0(mai_mai_n434_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n682_));
  NOi31      m660(.An(mai_mai_n682_), .B(mai_mai_n575_), .C(mai_mai_n44_), .Y(mai_mai_n683_));
  NA2        m661(.A(mai_mai_n122_), .B(i_13_), .Y(mai_mai_n684_));
  NO2        m662(.A(mai_mai_n625_), .B(mai_mai_n109_), .Y(mai_mai_n685_));
  INV        m663(.A(mai_mai_n685_), .Y(mai_mai_n686_));
  OAI220     m664(.A0(mai_mai_n686_), .A1(mai_mai_n68_), .B0(mai_mai_n684_), .B1(mai_mai_n666_), .Y(mai_mai_n687_));
  NO3        m665(.A(mai_mai_n68_), .B(mai_mai_n32_), .C(mai_mai_n95_), .Y(mai_mai_n688_));
  NA2        m666(.A(mai_mai_n26_), .B(mai_mai_n188_), .Y(mai_mai_n689_));
  NA2        m667(.A(mai_mai_n689_), .B(i_7_), .Y(mai_mai_n690_));
  NO3        m668(.A(mai_mai_n459_), .B(mai_mai_n230_), .C(mai_mai_n80_), .Y(mai_mai_n691_));
  AOI210     m669(.A0(mai_mai_n691_), .A1(mai_mai_n690_), .B0(mai_mai_n688_), .Y(mai_mai_n692_));
  NA2        m670(.A(mai_mai_n86_), .B(mai_mai_n96_), .Y(mai_mai_n693_));
  OAI220     m671(.A0(mai_mai_n693_), .A1(mai_mai_n580_), .B0(mai_mai_n692_), .B1(mai_mai_n591_), .Y(mai_mai_n694_));
  NO4        m672(.A(mai_mai_n694_), .B(mai_mai_n687_), .C(mai_mai_n683_), .D(mai_mai_n681_), .Y(mai_mai_n695_));
  OR2        m673(.A(i_11_), .B(i_6_), .Y(mai_mai_n696_));
  NA3        m674(.A(mai_mai_n579_), .B(mai_mai_n689_), .C(i_7_), .Y(mai_mai_n697_));
  AOI210     m675(.A0(mai_mai_n697_), .A1(mai_mai_n686_), .B0(mai_mai_n696_), .Y(mai_mai_n698_));
  NA3        m676(.A(mai_mai_n397_), .B(mai_mai_n583_), .C(mai_mai_n91_), .Y(mai_mai_n699_));
  NA2        m677(.A(mai_mai_n618_), .B(i_13_), .Y(mai_mai_n700_));
  NAi21      m678(.An(i_11_), .B(i_12_), .Y(mai_mai_n701_));
  NOi41      m679(.An(mai_mai_n105_), .B(mai_mai_n701_), .C(i_13_), .D(mai_mai_n80_), .Y(mai_mai_n702_));
  NO3        m680(.A(mai_mai_n459_), .B(mai_mai_n559_), .C(mai_mai_n584_), .Y(mai_mai_n703_));
  AOI210     m681(.A0(mai_mai_n703_), .A1(mai_mai_n297_), .B0(mai_mai_n702_), .Y(mai_mai_n704_));
  NA3        m682(.A(mai_mai_n704_), .B(mai_mai_n700_), .C(mai_mai_n699_), .Y(mai_mai_n705_));
  OAI210     m683(.A0(mai_mai_n705_), .A1(mai_mai_n698_), .B0(mai_mai_n62_), .Y(mai_mai_n706_));
  OAI210     m684(.A0(mai_mai_n230_), .A1(mai_mai_n358_), .B0(mai_mai_n356_), .Y(mai_mai_n707_));
  NO2        m685(.A(mai_mai_n123_), .B(i_2_), .Y(mai_mai_n708_));
  NA2        m686(.A(mai_mai_n708_), .B(mai_mai_n612_), .Y(mai_mai_n709_));
  NA2        m687(.A(mai_mai_n709_), .B(mai_mai_n707_), .Y(mai_mai_n710_));
  NA3        m688(.A(mai_mai_n710_), .B(mai_mai_n45_), .C(mai_mai_n219_), .Y(mai_mai_n711_));
  NA4        m689(.A(mai_mai_n711_), .B(mai_mai_n706_), .C(mai_mai_n695_), .D(mai_mai_n679_), .Y(mai_mai_n712_));
  OR4        m690(.A(mai_mai_n712_), .B(mai_mai_n671_), .C(mai_mai_n655_), .D(mai_mai_n594_), .Y(mai5));
  AOI210     m691(.A0(mai_mai_n641_), .A1(mai_mai_n255_), .B0(mai_mai_n404_), .Y(mai_mai_n714_));
  NO2        m692(.A(mai_mai_n580_), .B(i_11_), .Y(mai_mai_n715_));
  NA2        m693(.A(mai_mai_n83_), .B(mai_mai_n715_), .Y(mai_mai_n716_));
  NA2        m694(.A(mai_mai_n716_), .B(mai_mai_n714_), .Y(mai_mai_n717_));
  NO3        m695(.A(i_11_), .B(mai_mai_n230_), .C(i_13_), .Y(mai_mai_n718_));
  NO2        m696(.A(mai_mai_n119_), .B(mai_mai_n23_), .Y(mai_mai_n719_));
  NA2        m697(.A(i_12_), .B(i_8_), .Y(mai_mai_n720_));
  OAI210     m698(.A0(mai_mai_n46_), .A1(i_3_), .B0(mai_mai_n720_), .Y(mai_mai_n721_));
  INV        m699(.A(mai_mai_n433_), .Y(mai_mai_n722_));
  AOI220     m700(.A0(mai_mai_n303_), .A1(mai_mai_n552_), .B0(mai_mai_n721_), .B1(mai_mai_n719_), .Y(mai_mai_n723_));
  INV        m701(.A(mai_mai_n723_), .Y(mai_mai_n724_));
  NO2        m702(.A(mai_mai_n724_), .B(mai_mai_n717_), .Y(mai_mai_n725_));
  INV        m703(.A(mai_mai_n165_), .Y(mai_mai_n726_));
  INV        m704(.A(mai_mai_n237_), .Y(mai_mai_n727_));
  OAI210     m705(.A0(mai_mai_n667_), .A1(mai_mai_n435_), .B0(mai_mai_n105_), .Y(mai_mai_n728_));
  AOI210     m706(.A0(mai_mai_n728_), .A1(mai_mai_n727_), .B0(mai_mai_n726_), .Y(mai_mai_n729_));
  NO2        m707(.A(mai_mai_n442_), .B(mai_mai_n26_), .Y(mai_mai_n730_));
  NO2        m708(.A(mai_mai_n730_), .B(mai_mai_n406_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n731_), .B(i_2_), .Y(mai_mai_n732_));
  INV        m710(.A(mai_mai_n732_), .Y(mai_mai_n733_));
  AOI210     m711(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n403_), .Y(mai_mai_n734_));
  AOI210     m712(.A0(mai_mai_n734_), .A1(mai_mai_n733_), .B0(mai_mai_n729_), .Y(mai_mai_n735_));
  NO2        m713(.A(mai_mai_n185_), .B(mai_mai_n120_), .Y(mai_mai_n736_));
  OAI210     m714(.A0(mai_mai_n736_), .A1(mai_mai_n719_), .B0(i_2_), .Y(mai_mai_n737_));
  NO2        m715(.A(mai_mai_n737_), .B(mai_mai_n188_), .Y(mai_mai_n738_));
  OA210      m716(.A0(mai_mai_n597_), .A1(mai_mai_n121_), .B0(i_13_), .Y(mai_mai_n739_));
  NA2        m717(.A(mai_mai_n194_), .B(mai_mai_n197_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n146_), .B(mai_mai_n576_), .Y(mai_mai_n741_));
  AOI210     m719(.A0(mai_mai_n741_), .A1(mai_mai_n740_), .B0(mai_mai_n360_), .Y(mai_mai_n742_));
  AOI210     m720(.A0(mai_mai_n203_), .A1(mai_mai_n143_), .B0(mai_mai_n494_), .Y(mai_mai_n743_));
  NA2        m721(.A(mai_mai_n743_), .B(mai_mai_n406_), .Y(mai_mai_n744_));
  NO2        m722(.A(mai_mai_n96_), .B(mai_mai_n44_), .Y(mai_mai_n745_));
  INV        m723(.A(mai_mai_n286_), .Y(mai_mai_n746_));
  NA4        m724(.A(mai_mai_n746_), .B(mai_mai_n290_), .C(mai_mai_n119_), .D(mai_mai_n42_), .Y(mai_mai_n747_));
  OAI210     m725(.A0(mai_mai_n747_), .A1(mai_mai_n745_), .B0(mai_mai_n744_), .Y(mai_mai_n748_));
  NO4        m726(.A(mai_mai_n748_), .B(mai_mai_n742_), .C(mai_mai_n739_), .D(mai_mai_n738_), .Y(mai_mai_n749_));
  NA2        m727(.A(mai_mai_n552_), .B(mai_mai_n28_), .Y(mai_mai_n750_));
  NA2        m728(.A(mai_mai_n718_), .B(mai_mai_n260_), .Y(mai_mai_n751_));
  NA2        m729(.A(mai_mai_n751_), .B(mai_mai_n750_), .Y(mai_mai_n752_));
  NO2        m730(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n753_));
  NO2        m731(.A(mai_mai_n753_), .B(mai_mai_n121_), .Y(mai_mai_n754_));
  NO2        m732(.A(mai_mai_n754_), .B(mai_mai_n576_), .Y(mai_mai_n755_));
  AOI220     m733(.A0(mai_mai_n755_), .A1(mai_mai_n36_), .B0(mai_mai_n752_), .B1(mai_mai_n46_), .Y(mai_mai_n756_));
  NA4        m734(.A(mai_mai_n756_), .B(mai_mai_n749_), .C(mai_mai_n735_), .D(mai_mai_n725_), .Y(mai6));
  NO3        m735(.A(mai_mai_n244_), .B(mai_mai_n292_), .C(i_1_), .Y(mai_mai_n758_));
  NO2        m736(.A(mai_mai_n180_), .B(mai_mai_n134_), .Y(mai_mai_n759_));
  OAI210     m737(.A0(mai_mai_n759_), .A1(mai_mai_n758_), .B0(mai_mai_n708_), .Y(mai_mai_n760_));
  NA4        m738(.A(mai_mai_n376_), .B(mai_mai_n464_), .C(mai_mai_n68_), .D(mai_mai_n95_), .Y(mai_mai_n761_));
  INV        m739(.A(mai_mai_n761_), .Y(mai_mai_n762_));
  NO2        m740(.A(mai_mai_n215_), .B(mai_mai_n468_), .Y(mai_mai_n763_));
  NO2        m741(.A(i_11_), .B(i_9_), .Y(mai_mai_n764_));
  NO2        m742(.A(mai_mai_n762_), .B(mai_mai_n314_), .Y(mai_mai_n765_));
  AO210      m743(.A0(mai_mai_n765_), .A1(mai_mai_n760_), .B0(i_12_), .Y(mai_mai_n766_));
  NA2        m744(.A(mai_mai_n361_), .B(mai_mai_n321_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n559_), .B(mai_mai_n62_), .Y(mai_mai_n768_));
  NA2        m746(.A(mai_mai_n657_), .B(mai_mai_n68_), .Y(mai_mai_n769_));
  NA4        m747(.A(mai_mai_n602_), .B(mai_mai_n769_), .C(mai_mai_n768_), .D(mai_mai_n767_), .Y(mai_mai_n770_));
  INV        m748(.A(mai_mai_n191_), .Y(mai_mai_n771_));
  AOI220     m749(.A0(mai_mai_n771_), .A1(mai_mai_n764_), .B0(mai_mai_n770_), .B1(mai_mai_n70_), .Y(mai_mai_n772_));
  INV        m750(.A(mai_mai_n313_), .Y(mai_mai_n773_));
  NA2        m751(.A(mai_mai_n72_), .B(mai_mai_n126_), .Y(mai_mai_n774_));
  NO2        m752(.A(mai_mai_n774_), .B(mai_mai_n773_), .Y(mai_mai_n775_));
  NO2        m753(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n776_));
  NA3        m754(.A(mai_mai_n776_), .B(mai_mai_n455_), .C(mai_mai_n376_), .Y(mai_mai_n777_));
  NAi32      m755(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n778_));
  AOI210     m756(.A0(mai_mai_n696_), .A1(mai_mai_n81_), .B0(mai_mai_n778_), .Y(mai_mai_n779_));
  OAI210     m757(.A0(mai_mai_n656_), .A1(mai_mai_n540_), .B0(mai_mai_n539_), .Y(mai_mai_n780_));
  NAi31      m758(.An(mai_mai_n779_), .B(mai_mai_n780_), .C(mai_mai_n777_), .Y(mai_mai_n781_));
  OR2        m759(.A(mai_mai_n781_), .B(mai_mai_n775_), .Y(mai_mai_n782_));
  NO2        m760(.A(mai_mai_n672_), .B(i_2_), .Y(mai_mai_n783_));
  NA2        m761(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n784_));
  OAI210     m762(.A0(mai_mai_n784_), .A1(mai_mai_n396_), .B0(mai_mai_n346_), .Y(mai_mai_n785_));
  NA2        m763(.A(mai_mai_n785_), .B(mai_mai_n783_), .Y(mai_mai_n786_));
  AO220      m764(.A0(mai_mai_n345_), .A1(mai_mai_n335_), .B0(mai_mai_n382_), .B1(mai_mai_n576_), .Y(mai_mai_n787_));
  NA3        m765(.A(mai_mai_n787_), .B(mai_mai_n245_), .C(i_7_), .Y(mai_mai_n788_));
  OR2        m766(.A(mai_mai_n597_), .B(mai_mai_n435_), .Y(mai_mai_n789_));
  NA3        m767(.A(mai_mai_n789_), .B(mai_mai_n142_), .C(mai_mai_n66_), .Y(mai_mai_n790_));
  OR2        m768(.A(mai_mai_n722_), .B(mai_mai_n36_), .Y(mai_mai_n791_));
  NA4        m769(.A(mai_mai_n791_), .B(mai_mai_n790_), .C(mai_mai_n788_), .D(mai_mai_n786_), .Y(mai_mai_n792_));
  OAI210     m770(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n81_), .Y(mai_mai_n793_));
  AOI220     m771(.A0(mai_mai_n793_), .A1(mai_mai_n539_), .B0(mai_mai_n763_), .B1(mai_mai_n690_), .Y(mai_mai_n794_));
  NA3        m772(.A(mai_mai_n360_), .B(mai_mai_n231_), .C(mai_mai_n142_), .Y(mai_mai_n795_));
  NA2        m773(.A(mai_mai_n382_), .B(mai_mai_n67_), .Y(mai_mai_n796_));
  NA4        m774(.A(mai_mai_n796_), .B(mai_mai_n795_), .C(mai_mai_n794_), .D(mai_mai_n582_), .Y(mai_mai_n797_));
  AO210      m775(.A0(mai_mai_n494_), .A1(mai_mai_n46_), .B0(mai_mai_n82_), .Y(mai_mai_n798_));
  NA3        m776(.A(mai_mai_n798_), .B(mai_mai_n465_), .C(mai_mai_n213_), .Y(mai_mai_n799_));
  AOI210     m777(.A0(mai_mai_n435_), .A1(mai_mai_n433_), .B0(mai_mai_n538_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n587_), .B(mai_mai_n96_), .Y(mai_mai_n801_));
  OAI210     m779(.A0(mai_mai_n801_), .A1(mai_mai_n106_), .B0(mai_mai_n395_), .Y(mai_mai_n802_));
  INV        m780(.A(mai_mai_n565_), .Y(mai_mai_n803_));
  NA3        m781(.A(mai_mai_n803_), .B(mai_mai_n313_), .C(i_7_), .Y(mai_mai_n804_));
  NA4        m782(.A(mai_mai_n804_), .B(mai_mai_n802_), .C(mai_mai_n800_), .D(mai_mai_n799_), .Y(mai_mai_n805_));
  NO4        m783(.A(mai_mai_n805_), .B(mai_mai_n797_), .C(mai_mai_n792_), .D(mai_mai_n782_), .Y(mai_mai_n806_));
  NA4        m784(.A(mai_mai_n806_), .B(mai_mai_n772_), .C(mai_mai_n766_), .D(mai_mai_n367_), .Y(mai3));
  NA2        m785(.A(i_6_), .B(i_7_), .Y(mai_mai_n808_));
  NO2        m786(.A(mai_mai_n808_), .B(i_0_), .Y(mai_mai_n809_));
  NO2        m787(.A(i_11_), .B(mai_mai_n230_), .Y(mai_mai_n810_));
  OAI210     m788(.A0(mai_mai_n809_), .A1(mai_mai_n274_), .B0(mai_mai_n810_), .Y(mai_mai_n811_));
  INV        m789(.A(mai_mai_n811_), .Y(mai_mai_n812_));
  NO3        m790(.A(mai_mai_n438_), .B(mai_mai_n84_), .C(mai_mai_n44_), .Y(mai_mai_n813_));
  OA210      m791(.A0(mai_mai_n813_), .A1(mai_mai_n812_), .B0(mai_mai_n168_), .Y(mai_mai_n814_));
  INV        m792(.A(mai_mai_n795_), .Y(mai_mai_n815_));
  NA2        m793(.A(mai_mai_n815_), .B(mai_mai_n40_), .Y(mai_mai_n816_));
  NO3        m794(.A(mai_mai_n607_), .B(mai_mai_n442_), .C(mai_mai_n126_), .Y(mai_mai_n817_));
  NA2        m795(.A(mai_mai_n397_), .B(mai_mai_n45_), .Y(mai_mai_n818_));
  AN2        m796(.A(mai_mai_n440_), .B(mai_mai_n54_), .Y(mai_mai_n819_));
  NO2        m797(.A(mai_mai_n819_), .B(mai_mai_n817_), .Y(mai_mai_n820_));
  AOI210     m798(.A0(mai_mai_n820_), .A1(mai_mai_n816_), .B0(mai_mai_n48_), .Y(mai_mai_n821_));
  NO4        m799(.A(mai_mai_n364_), .B(mai_mai_n370_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n822_));
  NA2        m800(.A(mai_mai_n180_), .B(mai_mai_n548_), .Y(mai_mai_n823_));
  NOi21      m801(.An(mai_mai_n823_), .B(mai_mai_n822_), .Y(mai_mai_n824_));
  NA2        m802(.A(mai_mai_n682_), .B(mai_mai_n649_), .Y(mai_mai_n825_));
  NA2        m803(.A(mai_mai_n319_), .B(i_5_), .Y(mai_mai_n826_));
  OAI220     m804(.A0(mai_mai_n826_), .A1(mai_mai_n825_), .B0(mai_mai_n824_), .B1(mai_mai_n62_), .Y(mai_mai_n827_));
  NOi21      m805(.An(i_5_), .B(i_9_), .Y(mai_mai_n828_));
  NA2        m806(.A(mai_mai_n828_), .B(mai_mai_n432_), .Y(mai_mai_n829_));
  AOI210     m807(.A0(mai_mai_n252_), .A1(mai_mai_n457_), .B0(mai_mai_n661_), .Y(mai_mai_n830_));
  NO3        m808(.A(mai_mai_n400_), .B(mai_mai_n252_), .C(mai_mai_n70_), .Y(mai_mai_n831_));
  NO2        m809(.A(mai_mai_n169_), .B(mai_mai_n143_), .Y(mai_mai_n832_));
  AOI210     m810(.A0(mai_mai_n832_), .A1(mai_mai_n236_), .B0(mai_mai_n831_), .Y(mai_mai_n833_));
  OAI220     m811(.A0(mai_mai_n833_), .A1(mai_mai_n175_), .B0(mai_mai_n830_), .B1(mai_mai_n829_), .Y(mai_mai_n834_));
  NO4        m812(.A(mai_mai_n834_), .B(mai_mai_n827_), .C(mai_mai_n821_), .D(mai_mai_n814_), .Y(mai_mai_n835_));
  NA2        m813(.A(mai_mai_n180_), .B(mai_mai_n24_), .Y(mai_mai_n836_));
  NO2        m814(.A(mai_mai_n648_), .B(mai_mai_n573_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n837_), .B(mai_mai_n836_), .Y(mai_mai_n838_));
  NA2        m816(.A(mai_mai_n297_), .B(mai_mai_n124_), .Y(mai_mai_n839_));
  NAi21      m817(.An(mai_mai_n156_), .B(i_5_), .Y(mai_mai_n840_));
  NO2        m818(.A(mai_mai_n839_), .B(mai_mai_n387_), .Y(mai_mai_n841_));
  NO2        m819(.A(mai_mai_n841_), .B(mai_mai_n838_), .Y(mai_mai_n842_));
  NA2        m820(.A(mai_mai_n549_), .B(i_0_), .Y(mai_mai_n843_));
  NO3        m821(.A(mai_mai_n843_), .B(mai_mai_n371_), .C(mai_mai_n83_), .Y(mai_mai_n844_));
  NO4        m822(.A(mai_mai_n564_), .B(mai_mai_n210_), .C(mai_mai_n403_), .D(mai_mai_n396_), .Y(mai_mai_n845_));
  AOI210     m823(.A0(mai_mai_n845_), .A1(i_11_), .B0(mai_mai_n844_), .Y(mai_mai_n846_));
  AN2        m824(.A(mai_mai_n90_), .B(mai_mai_n235_), .Y(mai_mai_n847_));
  NA2        m825(.A(mai_mai_n718_), .B(mai_mai_n314_), .Y(mai_mai_n848_));
  AOI210     m826(.A0(mai_mai_n465_), .A1(mai_mai_n83_), .B0(mai_mai_n57_), .Y(mai_mai_n849_));
  OAI220     m827(.A0(mai_mai_n849_), .A1(mai_mai_n848_), .B0(mai_mai_n636_), .B1(mai_mai_n512_), .Y(mai_mai_n850_));
  INV        m828(.A(mai_mai_n514_), .Y(mai_mai_n851_));
  NO4        m829(.A(mai_mai_n109_), .B(mai_mai_n57_), .C(mai_mai_n645_), .D(i_5_), .Y(mai_mai_n852_));
  AN2        m830(.A(mai_mai_n852_), .B(mai_mai_n851_), .Y(mai_mai_n853_));
  NA2        m831(.A(mai_mai_n180_), .B(mai_mai_n79_), .Y(mai_mai_n854_));
  NA2        m832(.A(mai_mai_n543_), .B(i_4_), .Y(mai_mai_n855_));
  NA2        m833(.A(mai_mai_n183_), .B(mai_mai_n197_), .Y(mai_mai_n856_));
  OAI220     m834(.A0(mai_mai_n856_), .A1(mai_mai_n848_), .B0(mai_mai_n855_), .B1(mai_mai_n854_), .Y(mai_mai_n857_));
  NO4        m835(.A(mai_mai_n857_), .B(mai_mai_n853_), .C(mai_mai_n850_), .D(mai_mai_n847_), .Y(mai_mai_n858_));
  NA3        m836(.A(mai_mai_n858_), .B(mai_mai_n846_), .C(mai_mai_n842_), .Y(mai_mai_n859_));
  NO2        m837(.A(mai_mai_n97_), .B(mai_mai_n37_), .Y(mai_mai_n860_));
  NA2        m838(.A(i_11_), .B(i_9_), .Y(mai_mai_n861_));
  NO3        m839(.A(i_12_), .B(mai_mai_n861_), .C(mai_mai_n581_), .Y(mai_mai_n862_));
  AN2        m840(.A(mai_mai_n862_), .B(mai_mai_n860_), .Y(mai_mai_n863_));
  NA2        m841(.A(mai_mai_n380_), .B(mai_mai_n173_), .Y(mai_mai_n864_));
  NA2        m842(.A(mai_mai_n864_), .B(mai_mai_n154_), .Y(mai_mai_n865_));
  NO2        m843(.A(mai_mai_n861_), .B(mai_mai_n70_), .Y(mai_mai_n866_));
  NO2        m844(.A(mai_mai_n169_), .B(i_0_), .Y(mai_mai_n867_));
  INV        m845(.A(mai_mai_n867_), .Y(mai_mai_n868_));
  NA2        m846(.A(mai_mai_n455_), .B(mai_mai_n225_), .Y(mai_mai_n869_));
  AOI210     m847(.A0(mai_mai_n359_), .A1(i_4_), .B0(mai_mai_n394_), .Y(mai_mai_n870_));
  OAI220     m848(.A0(mai_mai_n870_), .A1(mai_mai_n829_), .B0(mai_mai_n869_), .B1(mai_mai_n868_), .Y(mai_mai_n871_));
  NO3        m849(.A(mai_mai_n871_), .B(mai_mai_n865_), .C(mai_mai_n863_), .Y(mai_mai_n872_));
  NA2        m850(.A(mai_mai_n635_), .B(mai_mai_n116_), .Y(mai_mai_n873_));
  NO2        m851(.A(i_6_), .B(mai_mai_n873_), .Y(mai_mai_n874_));
  AOI210     m852(.A0(mai_mai_n434_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n875_));
  NA2        m853(.A(mai_mai_n165_), .B(mai_mai_n97_), .Y(mai_mai_n876_));
  NOi32      m854(.An(mai_mai_n875_), .Bn(mai_mai_n183_), .C(mai_mai_n876_), .Y(mai_mai_n877_));
  NA2        m855(.A(mai_mai_n583_), .B(mai_mai_n314_), .Y(mai_mai_n878_));
  NO2        m856(.A(mai_mai_n878_), .B(mai_mai_n818_), .Y(mai_mai_n879_));
  NO3        m857(.A(mai_mai_n879_), .B(mai_mai_n877_), .C(mai_mai_n874_), .Y(mai_mai_n880_));
  NOi21      m858(.An(i_7_), .B(i_5_), .Y(mai_mai_n881_));
  NOi31      m859(.An(mai_mai_n881_), .B(i_0_), .C(mai_mai_n701_), .Y(mai_mai_n882_));
  OR2        m860(.A(mai_mai_n876_), .B(mai_mai_n493_), .Y(mai_mai_n883_));
  NO3        m861(.A(mai_mai_n390_), .B(mai_mai_n348_), .C(mai_mai_n344_), .Y(mai_mai_n884_));
  NO2        m862(.A(mai_mai_n246_), .B(mai_mai_n304_), .Y(mai_mai_n885_));
  INV        m863(.A(mai_mai_n701_), .Y(mai_mai_n886_));
  AOI210     m864(.A0(mai_mai_n886_), .A1(mai_mai_n885_), .B0(mai_mai_n884_), .Y(mai_mai_n887_));
  NA4        m865(.A(mai_mai_n887_), .B(mai_mai_n883_), .C(mai_mai_n880_), .D(mai_mai_n872_), .Y(mai_mai_n888_));
  AN2        m866(.A(mai_mai_n318_), .B(mai_mai_n314_), .Y(mai_mai_n889_));
  AN2        m867(.A(mai_mai_n889_), .B(mai_mai_n832_), .Y(mai_mai_n890_));
  NA2        m868(.A(mai_mai_n890_), .B(i_10_), .Y(mai_mai_n891_));
  OA210      m869(.A0(mai_mai_n455_), .A1(mai_mai_n217_), .B0(mai_mai_n454_), .Y(mai_mai_n892_));
  NA3        m870(.A(mai_mai_n454_), .B(mai_mai_n397_), .C(mai_mai_n45_), .Y(mai_mai_n893_));
  OAI210     m871(.A0(mai_mai_n840_), .A1(i_6_), .B0(mai_mai_n893_), .Y(mai_mai_n894_));
  NA2        m872(.A(mai_mai_n866_), .B(mai_mai_n290_), .Y(mai_mai_n895_));
  NA2        m873(.A(mai_mai_n182_), .B(mai_mai_n895_), .Y(mai_mai_n896_));
  AOI220     m874(.A0(mai_mai_n896_), .A1(mai_mai_n455_), .B0(mai_mai_n894_), .B1(mai_mai_n70_), .Y(mai_mai_n897_));
  NO2        m875(.A(mai_mai_n72_), .B(mai_mai_n720_), .Y(mai_mai_n898_));
  AOI210     m876(.A0(mai_mai_n168_), .A1(mai_mai_n573_), .B0(mai_mai_n898_), .Y(mai_mai_n899_));
  NO2        m877(.A(mai_mai_n899_), .B(mai_mai_n47_), .Y(mai_mai_n900_));
  NO3        m878(.A(mai_mai_n564_), .B(mai_mai_n343_), .C(mai_mai_n24_), .Y(mai_mai_n901_));
  NO2        m879(.A(mai_mai_n521_), .B(mai_mai_n901_), .Y(mai_mai_n902_));
  NAi21      m880(.An(i_9_), .B(i_5_), .Y(mai_mai_n903_));
  NO2        m881(.A(mai_mai_n903_), .B(mai_mai_n390_), .Y(mai_mai_n904_));
  NA2        m882(.A(mai_mai_n904_), .B(mai_mai_n597_), .Y(mai_mai_n905_));
  OAI220     m883(.A0(mai_mai_n905_), .A1(mai_mai_n80_), .B0(mai_mai_n902_), .B1(mai_mai_n166_), .Y(mai_mai_n906_));
  NO3        m884(.A(mai_mai_n906_), .B(mai_mai_n900_), .C(mai_mai_n497_), .Y(mai_mai_n907_));
  NA3        m885(.A(mai_mai_n907_), .B(mai_mai_n897_), .C(mai_mai_n891_), .Y(mai_mai_n908_));
  NO3        m886(.A(mai_mai_n908_), .B(mai_mai_n888_), .C(mai_mai_n859_), .Y(mai_mai_n909_));
  NO2        m887(.A(i_0_), .B(mai_mai_n701_), .Y(mai_mai_n910_));
  AOI210     m888(.A0(mai_mai_n768_), .A1(mai_mai_n659_), .B0(mai_mai_n876_), .Y(mai_mai_n911_));
  INV        m889(.A(mai_mai_n911_), .Y(mai_mai_n912_));
  NA3        m890(.A(mai_mai_n141_), .B(mai_mai_n649_), .C(mai_mai_n70_), .Y(mai_mai_n913_));
  NO2        m891(.A(mai_mai_n780_), .B(mai_mai_n390_), .Y(mai_mai_n914_));
  NA2        m892(.A(mai_mai_n810_), .B(i_9_), .Y(mai_mai_n915_));
  NO2        m893(.A(mai_mai_n474_), .B(mai_mai_n915_), .Y(mai_mai_n916_));
  NA2        m894(.A(mai_mai_n236_), .B(mai_mai_n224_), .Y(mai_mai_n917_));
  AOI210     m895(.A0(mai_mai_n917_), .A1(mai_mai_n843_), .B0(mai_mai_n147_), .Y(mai_mai_n918_));
  NO3        m896(.A(mai_mai_n918_), .B(mai_mai_n916_), .C(mai_mai_n914_), .Y(mai_mai_n919_));
  NA3        m897(.A(mai_mai_n919_), .B(mai_mai_n913_), .C(mai_mai_n912_), .Y(mai_mai_n920_));
  NA2        m898(.A(mai_mai_n889_), .B(mai_mai_n360_), .Y(mai_mai_n921_));
  AOI210     m899(.A0(mai_mai_n285_), .A1(mai_mai_n156_), .B0(mai_mai_n921_), .Y(mai_mai_n922_));
  NA3        m900(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n923_));
  NA2        m901(.A(i_5_), .B(mai_mai_n469_), .Y(mai_mai_n924_));
  AOI210     m902(.A0(mai_mai_n923_), .A1(mai_mai_n156_), .B0(mai_mai_n924_), .Y(mai_mai_n925_));
  NO2        m903(.A(mai_mai_n925_), .B(mai_mai_n922_), .Y(mai_mai_n926_));
  NA2        m904(.A(mai_mai_n544_), .B(mai_mai_n72_), .Y(mai_mai_n927_));
  NO3        m905(.A(mai_mai_n204_), .B(mai_mai_n370_), .C(i_0_), .Y(mai_mai_n928_));
  OAI210     m906(.A0(mai_mai_n928_), .A1(mai_mai_n73_), .B0(i_13_), .Y(mai_mai_n929_));
  INV        m907(.A(mai_mai_n213_), .Y(mai_mai_n930_));
  OAI220     m908(.A0(mai_mai_n506_), .A1(mai_mai_n134_), .B0(i_12_), .B1(mai_mai_n591_), .Y(mai_mai_n931_));
  NA3        m909(.A(mai_mai_n931_), .B(i_7_), .C(mai_mai_n930_), .Y(mai_mai_n932_));
  NA4        m910(.A(mai_mai_n932_), .B(mai_mai_n929_), .C(mai_mai_n927_), .D(mai_mai_n926_), .Y(mai_mai_n933_));
  INV        m911(.A(mai_mai_n87_), .Y(mai_mai_n934_));
  AOI210     m912(.A0(mai_mai_n934_), .A1(mai_mai_n910_), .B0(mai_mai_n103_), .Y(mai_mai_n935_));
  NA2        m913(.A(mai_mai_n881_), .B(mai_mai_n469_), .Y(mai_mai_n936_));
  NA2        m914(.A(mai_mai_n335_), .B(mai_mai_n170_), .Y(mai_mai_n937_));
  OA220      m915(.A0(mai_mai_n937_), .A1(mai_mai_n936_), .B0(mai_mai_n935_), .B1(i_5_), .Y(mai_mai_n938_));
  AOI210     m916(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n169_), .Y(mai_mai_n939_));
  NA2        m917(.A(mai_mai_n939_), .B(mai_mai_n892_), .Y(mai_mai_n940_));
  NA3        m918(.A(i_5_), .B(mai_mai_n274_), .C(mai_mai_n224_), .Y(mai_mai_n941_));
  INV        m919(.A(mai_mai_n941_), .Y(mai_mai_n942_));
  NA3        m920(.A(mai_mai_n376_), .B(mai_mai_n320_), .C(mai_mai_n216_), .Y(mai_mai_n943_));
  OAI210     m921(.A0(mai_mai_n823_), .A1(mai_mai_n623_), .B0(mai_mai_n943_), .Y(mai_mai_n944_));
  NO2        m922(.A(mai_mai_n944_), .B(mai_mai_n942_), .Y(mai_mai_n945_));
  NA3        m923(.A(mai_mai_n945_), .B(mai_mai_n940_), .C(mai_mai_n938_), .Y(mai_mai_n946_));
  NA2        m924(.A(mai_mai_n290_), .B(i_5_), .Y(mai_mai_n947_));
  NA2        m925(.A(mai_mai_n762_), .B(mai_mai_n170_), .Y(mai_mai_n948_));
  BUFFER     m926(.A(mai_mai_n147_), .Y(mai_mai_n949_));
  NO3        m927(.A(mai_mai_n949_), .B(i_12_), .C(mai_mai_n623_), .Y(mai_mai_n950_));
  NA2        m928(.A(mai_mai_n950_), .B(mai_mai_n213_), .Y(mai_mai_n951_));
  NA3        m929(.A(mai_mai_n92_), .B(mai_mai_n548_), .C(i_11_), .Y(mai_mai_n952_));
  NO2        m930(.A(mai_mai_n952_), .B(mai_mai_n149_), .Y(mai_mai_n953_));
  NA2        m931(.A(mai_mai_n881_), .B(mai_mai_n452_), .Y(mai_mai_n954_));
  OAI220     m932(.A0(i_7_), .A1(mai_mai_n947_), .B0(mai_mai_n954_), .B1(i_1_), .Y(mai_mai_n955_));
  AOI210     m933(.A0(mai_mai_n955_), .A1(mai_mai_n867_), .B0(mai_mai_n953_), .Y(mai_mai_n956_));
  NA3        m934(.A(mai_mai_n956_), .B(mai_mai_n951_), .C(mai_mai_n948_), .Y(mai_mai_n957_));
  NO4        m935(.A(mai_mai_n957_), .B(mai_mai_n946_), .C(mai_mai_n933_), .D(mai_mai_n920_), .Y(mai_mai_n958_));
  OAI210     m936(.A0(mai_mai_n783_), .A1(mai_mai_n776_), .B0(mai_mai_n37_), .Y(mai_mai_n959_));
  NA3        m937(.A(mai_mai_n875_), .B(mai_mai_n356_), .C(i_5_), .Y(mai_mai_n960_));
  NA3        m938(.A(mai_mai_n960_), .B(mai_mai_n959_), .C(mai_mai_n586_), .Y(mai_mai_n961_));
  NA2        m939(.A(mai_mai_n961_), .B(mai_mai_n201_), .Y(mai_mai_n962_));
  NA2        m940(.A(mai_mai_n181_), .B(mai_mai_n183_), .Y(mai_mai_n963_));
  AO210      m941(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n963_), .Y(mai_mai_n964_));
  OAI210     m942(.A0(mai_mai_n590_), .A1(mai_mai_n588_), .B0(mai_mai_n303_), .Y(mai_mai_n965_));
  NAi31      m943(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n966_));
  NO2        m944(.A(mai_mai_n67_), .B(mai_mai_n966_), .Y(mai_mai_n967_));
  INV        m945(.A(mai_mai_n967_), .Y(mai_mai_n968_));
  NA3        m946(.A(mai_mai_n968_), .B(mai_mai_n965_), .C(mai_mai_n964_), .Y(mai_mai_n969_));
  NO2        m947(.A(mai_mai_n444_), .B(mai_mai_n252_), .Y(mai_mai_n970_));
  NO2        m948(.A(mai_mai_n970_), .B(mai_mai_n845_), .Y(mai_mai_n971_));
  OAI210     m949(.A0(mai_mai_n952_), .A1(mai_mai_n143_), .B0(mai_mai_n971_), .Y(mai_mai_n972_));
  AOI210     m950(.A0(mai_mai_n969_), .A1(mai_mai_n48_), .B0(mai_mai_n972_), .Y(mai_mai_n973_));
  AOI210     m951(.A0(mai_mai_n973_), .A1(mai_mai_n962_), .B0(mai_mai_n70_), .Y(mai_mai_n974_));
  NO2        m952(.A(mai_mai_n541_), .B(mai_mai_n366_), .Y(mai_mai_n975_));
  NO2        m953(.A(mai_mai_n975_), .B(mai_mai_n726_), .Y(mai_mai_n976_));
  AOI210     m954(.A0(mai_mai_n939_), .A1(i_5_), .B0(mai_mai_n882_), .Y(mai_mai_n977_));
  NO2        m955(.A(mai_mai_n977_), .B(mai_mai_n650_), .Y(mai_mai_n978_));
  INV        m956(.A(mai_mai_n56_), .Y(mai_mai_n979_));
  AOI220     m957(.A0(mai_mai_n979_), .A1(mai_mai_n73_), .B0(mai_mai_n332_), .B1(mai_mai_n244_), .Y(mai_mai_n980_));
  NO2        m958(.A(mai_mai_n980_), .B(mai_mai_n230_), .Y(mai_mai_n981_));
  NO2        m959(.A(mai_mai_n981_), .B(mai_mai_n978_), .Y(mai_mai_n982_));
  OAI210     m960(.A0(mai_mai_n254_), .A1(mai_mai_n152_), .B0(mai_mai_n83_), .Y(mai_mai_n983_));
  NA3        m961(.A(mai_mai_n730_), .B(mai_mai_n274_), .C(mai_mai_n77_), .Y(mai_mai_n984_));
  AOI210     m962(.A0(mai_mai_n984_), .A1(mai_mai_n983_), .B0(i_11_), .Y(mai_mai_n985_));
  OAI210     m963(.A0(mai_mai_n1004_), .A1(mai_mai_n875_), .B0(mai_mai_n201_), .Y(mai_mai_n986_));
  NA2        m964(.A(mai_mai_n158_), .B(i_5_), .Y(mai_mai_n987_));
  AOI210     m965(.A0(mai_mai_n986_), .A1(mai_mai_n740_), .B0(mai_mai_n987_), .Y(mai_mai_n988_));
  NO3        m966(.A(mai_mai_n58_), .B(mai_mai_n57_), .C(i_4_), .Y(mai_mai_n989_));
  NA2        m967(.A(mai_mai_n292_), .B(mai_mai_n989_), .Y(mai_mai_n990_));
  NO2        m968(.A(mai_mai_n990_), .B(mai_mai_n701_), .Y(mai_mai_n991_));
  NO3        m969(.A(mai_mai_n903_), .B(mai_mai_n458_), .C(mai_mai_n243_), .Y(mai_mai_n992_));
  NO2        m970(.A(mai_mai_n992_), .B(mai_mai_n538_), .Y(mai_mai_n993_));
  INV        m971(.A(mai_mai_n349_), .Y(mai_mai_n994_));
  AOI210     m972(.A0(mai_mai_n994_), .A1(mai_mai_n993_), .B0(mai_mai_n41_), .Y(mai_mai_n995_));
  NO4        m973(.A(mai_mai_n995_), .B(mai_mai_n991_), .C(mai_mai_n988_), .D(mai_mai_n985_), .Y(mai_mai_n996_));
  OAI210     m974(.A0(mai_mai_n982_), .A1(i_4_), .B0(mai_mai_n996_), .Y(mai_mai_n997_));
  NO3        m975(.A(mai_mai_n997_), .B(mai_mai_n976_), .C(mai_mai_n974_), .Y(mai_mai_n998_));
  NA4        m976(.A(mai_mai_n998_), .B(mai_mai_n958_), .C(mai_mai_n909_), .D(mai_mai_n835_), .Y(mai4));
  INV        m977(.A(mai_mai_n676_), .Y(mai_mai_n1002_));
  INV        m978(.A(i_2_), .Y(mai_mai_n1003_));
  INV        m979(.A(i_12_), .Y(mai_mai_n1004_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  OAI210     u0028(.A0(men_men_n50_), .A1(i_3_), .B0(men_men_n48_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA2        u0042(.A(i_1_), .B(i_10_), .Y(men_men_n65_));
  NO2        u0043(.A(men_men_n65_), .B(i_6_), .Y(men_men_n66_));
  NAi21      u0044(.An(men_men_n66_), .B(men_men_n61_), .Y(men_men_n67_));
  NA2        u0045(.A(men_men_n50_), .B(i_2_), .Y(men_men_n68_));
  NA2        u0046(.A(i_1_), .B(i_6_), .Y(men_men_n69_));
  NO2        u0047(.A(men_men_n69_), .B(men_men_n25_), .Y(men_men_n70_));
  INV        u0048(.A(i_0_), .Y(men_men_n71_));
  NAi21      u0049(.An(i_5_), .B(i_10_), .Y(men_men_n72_));
  NA2        u0050(.A(i_5_), .B(i_9_), .Y(men_men_n73_));
  AOI210     u0051(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n71_), .Y(men_men_n74_));
  NO2        u0052(.A(men_men_n74_), .B(men_men_n70_), .Y(men_men_n75_));
  INV        u0053(.A(men_men_n75_), .Y(men_men_n76_));
  OAI210     u0054(.A0(men_men_n76_), .A1(men_men_n67_), .B0(i_0_), .Y(men_men_n77_));
  NA2        u0055(.A(i_12_), .B(i_5_), .Y(men_men_n78_));
  NA2        u0056(.A(i_2_), .B(i_8_), .Y(men_men_n79_));
  NO2        u0057(.A(men_men_n79_), .B(men_men_n58_), .Y(men_men_n80_));
  NO2        u0058(.A(i_3_), .B(i_9_), .Y(men_men_n81_));
  NO2        u0059(.A(i_3_), .B(i_7_), .Y(men_men_n82_));
  NO3        u0060(.A(men_men_n82_), .B(men_men_n81_), .C(men_men_n63_), .Y(men_men_n83_));
  INV        u0061(.A(i_6_), .Y(men_men_n84_));
  OR4        u0062(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n85_));
  INV        u0063(.A(men_men_n85_), .Y(men_men_n86_));
  NO2        u0064(.A(i_2_), .B(i_7_), .Y(men_men_n87_));
  NO2        u0065(.A(men_men_n86_), .B(men_men_n87_), .Y(men_men_n88_));
  OAI210     u0066(.A0(men_men_n83_), .A1(men_men_n80_), .B0(men_men_n88_), .Y(men_men_n89_));
  NAi21      u0067(.An(i_6_), .B(i_10_), .Y(men_men_n90_));
  NA2        u0068(.A(i_6_), .B(i_9_), .Y(men_men_n91_));
  AOI210     u0069(.A0(men_men_n91_), .A1(men_men_n90_), .B0(men_men_n63_), .Y(men_men_n92_));
  NA2        u0070(.A(i_2_), .B(i_6_), .Y(men_men_n93_));
  NO3        u0071(.A(men_men_n93_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n94_));
  NO2        u0072(.A(men_men_n94_), .B(men_men_n92_), .Y(men_men_n95_));
  AOI210     u0073(.A0(men_men_n95_), .A1(men_men_n89_), .B0(men_men_n78_), .Y(men_men_n96_));
  AN3        u0074(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n97_));
  NAi21      u0075(.An(i_6_), .B(i_11_), .Y(men_men_n98_));
  NO2        u0076(.A(i_5_), .B(i_8_), .Y(men_men_n99_));
  NOi21      u0077(.An(men_men_n99_), .B(men_men_n98_), .Y(men_men_n100_));
  AOI220     u0078(.A0(men_men_n100_), .A1(men_men_n62_), .B0(men_men_n97_), .B1(men_men_n32_), .Y(men_men_n101_));
  INV        u0079(.A(i_7_), .Y(men_men_n102_));
  NA2        u0080(.A(men_men_n46_), .B(men_men_n102_), .Y(men_men_n103_));
  NO2        u0081(.A(i_0_), .B(i_5_), .Y(men_men_n104_));
  NO2        u0082(.A(men_men_n104_), .B(men_men_n84_), .Y(men_men_n105_));
  NA2        u0083(.A(i_12_), .B(i_3_), .Y(men_men_n106_));
  INV        u0084(.A(men_men_n106_), .Y(men_men_n107_));
  NA3        u0085(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n103_), .Y(men_men_n108_));
  NAi21      u0086(.An(i_7_), .B(i_11_), .Y(men_men_n109_));
  NO3        u0087(.A(men_men_n109_), .B(men_men_n90_), .C(men_men_n53_), .Y(men_men_n110_));
  AN2        u0088(.A(i_2_), .B(i_10_), .Y(men_men_n111_));
  NO2        u0089(.A(men_men_n111_), .B(i_7_), .Y(men_men_n112_));
  OR2        u0090(.A(men_men_n78_), .B(men_men_n58_), .Y(men_men_n113_));
  NO2        u0091(.A(i_8_), .B(men_men_n102_), .Y(men_men_n114_));
  NO3        u0092(.A(men_men_n114_), .B(men_men_n113_), .C(men_men_n112_), .Y(men_men_n115_));
  NA2        u0093(.A(i_12_), .B(i_7_), .Y(men_men_n116_));
  NO2        u0094(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n117_));
  NA2        u0095(.A(men_men_n117_), .B(i_0_), .Y(men_men_n118_));
  NA2        u0096(.A(i_11_), .B(i_12_), .Y(men_men_n119_));
  OAI210     u0097(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n119_), .Y(men_men_n120_));
  NO2        u0098(.A(men_men_n120_), .B(men_men_n115_), .Y(men_men_n121_));
  NAi41      u0099(.An(men_men_n110_), .B(men_men_n121_), .C(men_men_n108_), .D(men_men_n101_), .Y(men_men_n122_));
  NOi21      u0100(.An(i_1_), .B(i_5_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n123_), .B(i_11_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n102_), .B(men_men_n37_), .Y(men_men_n125_));
  NA2        u0103(.A(i_7_), .B(men_men_n25_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n126_), .B(men_men_n125_), .Y(men_men_n127_));
  NO2        u0105(.A(men_men_n127_), .B(men_men_n46_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n129_));
  NAi21      u0107(.An(i_3_), .B(i_8_), .Y(men_men_n130_));
  NA2        u0108(.A(men_men_n130_), .B(men_men_n62_), .Y(men_men_n131_));
  NOi31      u0109(.An(men_men_n131_), .B(men_men_n129_), .C(men_men_n128_), .Y(men_men_n132_));
  NO2        u0110(.A(i_1_), .B(men_men_n84_), .Y(men_men_n133_));
  NO2        u0111(.A(i_6_), .B(i_5_), .Y(men_men_n134_));
  NA2        u0112(.A(men_men_n134_), .B(i_3_), .Y(men_men_n135_));
  AO210      u0113(.A0(men_men_n135_), .A1(men_men_n47_), .B0(men_men_n133_), .Y(men_men_n136_));
  OAI220     u0114(.A0(men_men_n136_), .A1(men_men_n109_), .B0(men_men_n132_), .B1(men_men_n124_), .Y(men_men_n137_));
  NO3        u0115(.A(men_men_n137_), .B(men_men_n122_), .C(men_men_n96_), .Y(men_men_n138_));
  NA3        u0116(.A(men_men_n138_), .B(men_men_n77_), .C(men_men_n56_), .Y(men2));
  NO2        u0117(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n140_));
  INV        u0118(.A(i_6_), .Y(men_men_n141_));
  NA2        u0119(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n142_));
  NA4        u0120(.A(men_men_n142_), .B(men_men_n75_), .C(men_men_n68_), .D(men_men_n30_), .Y(men0));
  AN2        u0121(.A(i_8_), .B(i_7_), .Y(men_men_n144_));
  NA2        u0122(.A(men_men_n144_), .B(i_6_), .Y(men_men_n145_));
  NO2        u0123(.A(i_12_), .B(i_13_), .Y(men_men_n146_));
  NAi21      u0124(.An(i_5_), .B(i_11_), .Y(men_men_n147_));
  NOi21      u0125(.An(men_men_n146_), .B(men_men_n147_), .Y(men_men_n148_));
  NO2        u0126(.A(i_0_), .B(i_1_), .Y(men_men_n149_));
  NA2        u0127(.A(i_2_), .B(i_3_), .Y(men_men_n150_));
  NO2        u0128(.A(men_men_n150_), .B(i_4_), .Y(men_men_n151_));
  NA3        u0129(.A(men_men_n151_), .B(men_men_n149_), .C(men_men_n148_), .Y(men_men_n152_));
  OR2        u0130(.A(men_men_n152_), .B(men_men_n25_), .Y(men_men_n153_));
  AN2        u0131(.A(men_men_n146_), .B(men_men_n81_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n154_), .B(men_men_n27_), .Y(men_men_n155_));
  NA2        u0133(.A(i_1_), .B(i_5_), .Y(men_men_n156_));
  NO2        u0134(.A(men_men_n71_), .B(men_men_n46_), .Y(men_men_n157_));
  NA2        u0135(.A(men_men_n157_), .B(men_men_n36_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n156_), .C(men_men_n155_), .Y(men_men_n159_));
  OR2        u0137(.A(i_0_), .B(i_1_), .Y(men_men_n160_));
  NO3        u0138(.A(men_men_n160_), .B(men_men_n78_), .C(i_13_), .Y(men_men_n161_));
  NAi32      u0139(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n162_));
  NAi21      u0140(.An(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  NOi21      u0141(.An(i_4_), .B(i_10_), .Y(men_men_n164_));
  NA2        u0142(.A(men_men_n164_), .B(men_men_n39_), .Y(men_men_n165_));
  NO2        u0143(.A(i_3_), .B(i_5_), .Y(men_men_n166_));
  NO3        u0144(.A(men_men_n71_), .B(i_2_), .C(i_1_), .Y(men_men_n167_));
  NA2        u0145(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  OAI210     u0146(.A0(men_men_n168_), .A1(men_men_n165_), .B0(men_men_n163_), .Y(men_men_n169_));
  NO2        u0147(.A(men_men_n169_), .B(men_men_n159_), .Y(men_men_n170_));
  AOI210     u0148(.A0(men_men_n170_), .A1(men_men_n153_), .B0(men_men_n145_), .Y(men_men_n171_));
  NA3        u0149(.A(men_men_n71_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n172_));
  NA2        u0150(.A(i_3_), .B(men_men_n48_), .Y(men_men_n173_));
  NOi21      u0151(.An(i_4_), .B(i_9_), .Y(men_men_n174_));
  NOi21      u0152(.An(i_11_), .B(i_13_), .Y(men_men_n175_));
  NA2        u0153(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  OR2        u0154(.A(men_men_n176_), .B(men_men_n173_), .Y(men_men_n177_));
  NO2        u0155(.A(i_4_), .B(i_5_), .Y(men_men_n178_));
  NAi21      u0156(.An(i_12_), .B(i_11_), .Y(men_men_n179_));
  NO2        u0157(.A(men_men_n179_), .B(i_13_), .Y(men_men_n180_));
  NA3        u0158(.A(men_men_n180_), .B(men_men_n178_), .C(men_men_n81_), .Y(men_men_n181_));
  AOI210     u0159(.A0(men_men_n181_), .A1(men_men_n177_), .B0(men_men_n172_), .Y(men_men_n182_));
  NO2        u0160(.A(men_men_n71_), .B(men_men_n63_), .Y(men_men_n183_));
  NA2        u0161(.A(men_men_n183_), .B(men_men_n46_), .Y(men_men_n184_));
  NA2        u0162(.A(men_men_n36_), .B(i_5_), .Y(men_men_n185_));
  NAi31      u0163(.An(men_men_n185_), .B(men_men_n154_), .C(i_11_), .Y(men_men_n186_));
  NA2        u0164(.A(i_3_), .B(i_5_), .Y(men_men_n187_));
  OR2        u0165(.A(men_men_n187_), .B(men_men_n176_), .Y(men_men_n188_));
  AOI210     u0166(.A0(men_men_n188_), .A1(men_men_n186_), .B0(men_men_n184_), .Y(men_men_n189_));
  NO2        u0167(.A(men_men_n71_), .B(i_5_), .Y(men_men_n190_));
  NO2        u0168(.A(i_13_), .B(i_10_), .Y(men_men_n191_));
  NA3        u0169(.A(men_men_n191_), .B(men_men_n190_), .C(men_men_n44_), .Y(men_men_n192_));
  NO2        u0170(.A(i_2_), .B(i_1_), .Y(men_men_n193_));
  NA2        u0171(.A(men_men_n193_), .B(i_3_), .Y(men_men_n194_));
  NAi21      u0172(.An(i_4_), .B(i_12_), .Y(men_men_n195_));
  NO4        u0173(.A(men_men_n195_), .B(men_men_n194_), .C(men_men_n192_), .D(men_men_n25_), .Y(men_men_n196_));
  NO3        u0174(.A(men_men_n196_), .B(men_men_n189_), .C(men_men_n182_), .Y(men_men_n197_));
  INV        u0175(.A(i_8_), .Y(men_men_n198_));
  NO2        u0176(.A(men_men_n198_), .B(i_7_), .Y(men_men_n199_));
  NA2        u0177(.A(men_men_n199_), .B(i_6_), .Y(men_men_n200_));
  NO3        u0178(.A(i_3_), .B(men_men_n84_), .C(men_men_n48_), .Y(men_men_n201_));
  NA2        u0179(.A(men_men_n201_), .B(men_men_n114_), .Y(men_men_n202_));
  NO3        u0180(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n203_));
  NA3        u0181(.A(men_men_n203_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n204_));
  NO3        u0182(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n205_));
  OAI210     u0183(.A0(men_men_n97_), .A1(i_12_), .B0(men_men_n205_), .Y(men_men_n206_));
  AOI210     u0184(.A0(men_men_n206_), .A1(men_men_n204_), .B0(men_men_n202_), .Y(men_men_n207_));
  NO2        u0185(.A(i_3_), .B(i_8_), .Y(men_men_n208_));
  NO3        u0186(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n209_));
  NA3        u0187(.A(men_men_n209_), .B(men_men_n208_), .C(men_men_n39_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n104_), .B(men_men_n58_), .Y(men_men_n211_));
  NO2        u0189(.A(i_13_), .B(i_9_), .Y(men_men_n212_));
  NAi21      u0190(.An(i_12_), .B(i_3_), .Y(men_men_n213_));
  OR2        u0191(.A(men_men_n213_), .B(i_8_), .Y(men_men_n214_));
  NO2        u0192(.A(men_men_n44_), .B(i_5_), .Y(men_men_n215_));
  NO3        u0193(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n216_));
  NA3        u0194(.A(men_men_n216_), .B(men_men_n215_), .C(i_10_), .Y(men_men_n217_));
  OAI220     u0195(.A0(men_men_n217_), .A1(men_men_n214_), .B0(men_men_n104_), .B1(men_men_n210_), .Y(men_men_n218_));
  AOI210     u0196(.A0(men_men_n218_), .A1(i_7_), .B0(men_men_n207_), .Y(men_men_n219_));
  OAI220     u0197(.A0(men_men_n219_), .A1(i_4_), .B0(men_men_n200_), .B1(men_men_n197_), .Y(men_men_n220_));
  NAi21      u0198(.An(i_12_), .B(i_7_), .Y(men_men_n221_));
  NA3        u0199(.A(i_13_), .B(men_men_n198_), .C(i_10_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n222_), .B(men_men_n221_), .Y(men_men_n223_));
  NA2        u0201(.A(i_0_), .B(i_5_), .Y(men_men_n224_));
  NA2        u0202(.A(men_men_n224_), .B(men_men_n105_), .Y(men_men_n225_));
  OAI220     u0203(.A0(men_men_n225_), .A1(men_men_n194_), .B0(men_men_n184_), .B1(men_men_n135_), .Y(men_men_n226_));
  NAi31      u0204(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n227_));
  NO2        u0205(.A(men_men_n36_), .B(i_13_), .Y(men_men_n228_));
  NO2        u0206(.A(men_men_n71_), .B(men_men_n26_), .Y(men_men_n229_));
  NO2        u0207(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n230_));
  NA3        u0208(.A(men_men_n230_), .B(men_men_n229_), .C(men_men_n228_), .Y(men_men_n231_));
  INV        u0209(.A(i_13_), .Y(men_men_n232_));
  NO2        u0210(.A(i_12_), .B(men_men_n232_), .Y(men_men_n233_));
  NA3        u0211(.A(men_men_n233_), .B(men_men_n203_), .C(men_men_n201_), .Y(men_men_n234_));
  OAI210     u0212(.A0(men_men_n231_), .A1(men_men_n227_), .B0(men_men_n234_), .Y(men_men_n235_));
  AOI220     u0213(.A0(men_men_n235_), .A1(men_men_n144_), .B0(men_men_n226_), .B1(men_men_n223_), .Y(men_men_n236_));
  NO2        u0214(.A(i_12_), .B(men_men_n37_), .Y(men_men_n237_));
  NO2        u0215(.A(men_men_n187_), .B(i_4_), .Y(men_men_n238_));
  NA2        u0216(.A(men_men_n238_), .B(men_men_n237_), .Y(men_men_n239_));
  OR2        u0217(.A(i_8_), .B(i_7_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n240_), .B(men_men_n84_), .Y(men_men_n241_));
  NO2        u0219(.A(men_men_n53_), .B(i_1_), .Y(men_men_n242_));
  NA2        u0220(.A(men_men_n242_), .B(men_men_n241_), .Y(men_men_n243_));
  INV        u0221(.A(i_12_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n44_), .B(men_men_n244_), .Y(men_men_n245_));
  NO3        u0223(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n246_));
  NA2        u0224(.A(i_2_), .B(i_1_), .Y(men_men_n247_));
  NO2        u0225(.A(men_men_n243_), .B(men_men_n239_), .Y(men_men_n248_));
  NO3        u0226(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n249_));
  NAi21      u0227(.An(i_4_), .B(i_3_), .Y(men_men_n250_));
  NO2        u0228(.A(men_men_n250_), .B(men_men_n73_), .Y(men_men_n251_));
  NO2        u0229(.A(i_0_), .B(i_6_), .Y(men_men_n252_));
  NOi41      u0230(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n253_));
  NA2        u0231(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NO2        u0232(.A(men_men_n247_), .B(men_men_n187_), .Y(men_men_n255_));
  INV        u0233(.A(men_men_n248_), .Y(men_men_n256_));
  NO2        u0234(.A(i_11_), .B(men_men_n232_), .Y(men_men_n257_));
  NOi21      u0235(.An(i_1_), .B(i_6_), .Y(men_men_n258_));
  NA2        u0236(.A(men_men_n244_), .B(i_9_), .Y(men_men_n259_));
  OR4        u0237(.A(men_men_n259_), .B(i_3_), .C(men_men_n258_), .D(men_men_n190_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n261_));
  NO2        u0239(.A(i_12_), .B(i_3_), .Y(men_men_n262_));
  NA2        u0240(.A(men_men_n71_), .B(i_5_), .Y(men_men_n263_));
  NA2        u0241(.A(i_3_), .B(i_9_), .Y(men_men_n264_));
  NAi21      u0242(.An(i_7_), .B(i_10_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n265_), .B(men_men_n264_), .Y(men_men_n266_));
  NA3        u0244(.A(men_men_n266_), .B(men_men_n263_), .C(men_men_n64_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n267_), .B(men_men_n260_), .Y(men_men_n268_));
  NA3        u0246(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n269_));
  INV        u0247(.A(men_men_n145_), .Y(men_men_n270_));
  NA2        u0248(.A(men_men_n244_), .B(i_13_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n271_), .B(men_men_n73_), .Y(men_men_n272_));
  AOI220     u0250(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n268_), .B1(men_men_n257_), .Y(men_men_n273_));
  NO2        u0251(.A(men_men_n240_), .B(men_men_n37_), .Y(men_men_n274_));
  NA2        u0252(.A(i_12_), .B(i_6_), .Y(men_men_n275_));
  OR2        u0253(.A(i_13_), .B(i_9_), .Y(men_men_n276_));
  NO3        u0254(.A(men_men_n276_), .B(men_men_n275_), .C(men_men_n48_), .Y(men_men_n277_));
  NO2        u0255(.A(men_men_n250_), .B(i_2_), .Y(men_men_n278_));
  NA3        u0256(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n44_), .Y(men_men_n279_));
  NA2        u0257(.A(men_men_n257_), .B(i_9_), .Y(men_men_n280_));
  OAI210     u0258(.A0(men_men_n71_), .A1(men_men_n280_), .B0(men_men_n279_), .Y(men_men_n281_));
  NA2        u0259(.A(men_men_n157_), .B(men_men_n63_), .Y(men_men_n282_));
  NO3        u0260(.A(i_11_), .B(men_men_n232_), .C(men_men_n25_), .Y(men_men_n283_));
  NO2        u0261(.A(i_6_), .B(men_men_n48_), .Y(men_men_n284_));
  NA3        u0262(.A(men_men_n284_), .B(i_7_), .C(men_men_n283_), .Y(men_men_n285_));
  NA3        u0263(.A(men_men_n1084_), .B(men_men_n274_), .C(men_men_n233_), .Y(men_men_n286_));
  AOI210     u0264(.A0(men_men_n286_), .A1(men_men_n285_), .B0(men_men_n282_), .Y(men_men_n287_));
  AOI210     u0265(.A0(men_men_n281_), .A1(men_men_n274_), .B0(men_men_n287_), .Y(men_men_n288_));
  NA4        u0266(.A(men_men_n288_), .B(men_men_n273_), .C(men_men_n256_), .D(men_men_n236_), .Y(men_men_n289_));
  NO3        u0267(.A(i_12_), .B(men_men_n232_), .C(men_men_n37_), .Y(men_men_n290_));
  INV        u0268(.A(men_men_n290_), .Y(men_men_n291_));
  NOi21      u0269(.An(men_men_n166_), .B(men_men_n84_), .Y(men_men_n292_));
  NO3        u0270(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n293_));
  AOI220     u0271(.A0(men_men_n293_), .A1(men_men_n201_), .B0(men_men_n292_), .B1(men_men_n242_), .Y(men_men_n294_));
  NO2        u0272(.A(men_men_n294_), .B(i_7_), .Y(men_men_n295_));
  NO3        u0273(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n296_));
  NO2        u0274(.A(men_men_n247_), .B(i_0_), .Y(men_men_n297_));
  AOI220     u0275(.A0(men_men_n297_), .A1(men_men_n199_), .B0(men_men_n296_), .B1(men_men_n144_), .Y(men_men_n298_));
  NA2        u0276(.A(men_men_n284_), .B(men_men_n26_), .Y(men_men_n299_));
  NO2        u0277(.A(men_men_n299_), .B(men_men_n298_), .Y(men_men_n300_));
  NA2        u0278(.A(i_0_), .B(i_1_), .Y(men_men_n301_));
  NO2        u0279(.A(men_men_n301_), .B(i_2_), .Y(men_men_n302_));
  NO2        u0280(.A(men_men_n59_), .B(i_6_), .Y(men_men_n303_));
  NA3        u0281(.A(men_men_n303_), .B(men_men_n302_), .C(men_men_n166_), .Y(men_men_n304_));
  OAI210     u0282(.A0(men_men_n168_), .A1(men_men_n145_), .B0(men_men_n304_), .Y(men_men_n305_));
  NO3        u0283(.A(men_men_n305_), .B(men_men_n300_), .C(men_men_n295_), .Y(men_men_n306_));
  NO2        u0284(.A(i_3_), .B(i_10_), .Y(men_men_n307_));
  NA3        u0285(.A(men_men_n307_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n308_));
  NO2        u0286(.A(i_2_), .B(men_men_n102_), .Y(men_men_n309_));
  NOi21      u0287(.An(men_men_n224_), .B(men_men_n104_), .Y(men_men_n310_));
  NA3        u0288(.A(men_men_n310_), .B(men_men_n36_), .C(men_men_n309_), .Y(men_men_n311_));
  AN2        u0289(.A(i_3_), .B(i_10_), .Y(men_men_n312_));
  NA4        u0290(.A(men_men_n312_), .B(men_men_n203_), .C(men_men_n180_), .D(men_men_n178_), .Y(men_men_n313_));
  NO2        u0291(.A(i_5_), .B(men_men_n37_), .Y(men_men_n314_));
  NO2        u0292(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n315_));
  OR2        u0293(.A(men_men_n311_), .B(men_men_n308_), .Y(men_men_n316_));
  OAI220     u0294(.A0(men_men_n316_), .A1(i_6_), .B0(men_men_n306_), .B1(men_men_n291_), .Y(men_men_n317_));
  NO4        u0295(.A(men_men_n317_), .B(men_men_n289_), .C(men_men_n220_), .D(men_men_n171_), .Y(men_men_n318_));
  NO3        u0296(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n319_));
  NO3        u0297(.A(i_6_), .B(men_men_n198_), .C(i_7_), .Y(men_men_n320_));
  NA2        u0298(.A(men_men_n320_), .B(men_men_n203_), .Y(men_men_n321_));
  AOI210     u0299(.A0(men_men_n321_), .A1(men_men_n247_), .B0(men_men_n173_), .Y(men_men_n322_));
  NO2        u0300(.A(i_2_), .B(i_3_), .Y(men_men_n323_));
  OR2        u0301(.A(i_0_), .B(i_5_), .Y(men_men_n324_));
  NA2        u0302(.A(men_men_n224_), .B(men_men_n324_), .Y(men_men_n325_));
  NA3        u0303(.A(men_men_n325_), .B(men_men_n241_), .C(men_men_n323_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n297_), .B(men_men_n292_), .C(men_men_n114_), .Y(men_men_n327_));
  NO2        u0305(.A(i_8_), .B(i_6_), .Y(men_men_n328_));
  NO2        u0306(.A(men_men_n160_), .B(men_men_n46_), .Y(men_men_n329_));
  NA3        u0307(.A(men_men_n329_), .B(men_men_n328_), .C(men_men_n166_), .Y(men_men_n330_));
  NA3        u0308(.A(men_men_n330_), .B(men_men_n327_), .C(men_men_n326_), .Y(men_men_n331_));
  OAI210     u0309(.A0(men_men_n331_), .A1(men_men_n322_), .B0(i_4_), .Y(men_men_n332_));
  NO2        u0310(.A(i_12_), .B(i_10_), .Y(men_men_n333_));
  NOi21      u0311(.An(i_5_), .B(i_0_), .Y(men_men_n334_));
  AOI210     u0312(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n102_), .Y(men_men_n335_));
  NO4        u0313(.A(men_men_n335_), .B(i_4_), .C(men_men_n334_), .D(men_men_n130_), .Y(men_men_n336_));
  NA4        u0314(.A(men_men_n82_), .B(men_men_n36_), .C(men_men_n84_), .D(i_8_), .Y(men_men_n337_));
  NA2        u0315(.A(men_men_n336_), .B(men_men_n333_), .Y(men_men_n338_));
  NO2        u0316(.A(i_6_), .B(i_8_), .Y(men_men_n339_));
  AN2        u0317(.A(i_0_), .B(men_men_n339_), .Y(men_men_n340_));
  NO2        u0318(.A(i_1_), .B(i_7_), .Y(men_men_n341_));
  NA3        u0319(.A(men_men_n340_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n342_));
  NA3        u0320(.A(men_men_n342_), .B(men_men_n338_), .C(men_men_n332_), .Y(men_men_n343_));
  NO2        u0321(.A(i_8_), .B(men_men_n325_), .Y(men_men_n344_));
  NOi21      u0322(.An(men_men_n156_), .B(men_men_n105_), .Y(men_men_n345_));
  NO2        u0323(.A(men_men_n345_), .B(men_men_n126_), .Y(men_men_n346_));
  OAI210     u0324(.A0(men_men_n346_), .A1(men_men_n344_), .B0(i_3_), .Y(men_men_n347_));
  NO2        u0325(.A(men_men_n301_), .B(men_men_n79_), .Y(men_men_n348_));
  NA2        u0326(.A(men_men_n348_), .B(men_men_n134_), .Y(men_men_n349_));
  NO2        u0327(.A(men_men_n93_), .B(men_men_n198_), .Y(men_men_n350_));
  NA3        u0328(.A(men_men_n310_), .B(men_men_n350_), .C(men_men_n63_), .Y(men_men_n351_));
  AOI210     u0329(.A0(men_men_n351_), .A1(men_men_n349_), .B0(i_3_), .Y(men_men_n352_));
  NO2        u0330(.A(men_men_n198_), .B(i_9_), .Y(men_men_n353_));
  NA2        u0331(.A(men_men_n353_), .B(men_men_n211_), .Y(men_men_n354_));
  NO2        u0332(.A(men_men_n354_), .B(men_men_n46_), .Y(men_men_n355_));
  NO3        u0333(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n300_), .Y(men_men_n356_));
  AOI210     u0334(.A0(men_men_n356_), .A1(men_men_n347_), .B0(men_men_n165_), .Y(men_men_n357_));
  AOI210     u0335(.A0(men_men_n343_), .A1(men_men_n319_), .B0(men_men_n357_), .Y(men_men_n358_));
  NOi32      u0336(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n359_));
  INV        u0337(.A(men_men_n359_), .Y(men_men_n360_));
  NAi21      u0338(.An(i_0_), .B(i_6_), .Y(men_men_n361_));
  NAi21      u0339(.An(i_1_), .B(i_5_), .Y(men_men_n362_));
  NA2        u0340(.A(men_men_n362_), .B(men_men_n361_), .Y(men_men_n363_));
  NA2        u0341(.A(men_men_n363_), .B(men_men_n25_), .Y(men_men_n364_));
  OAI210     u0342(.A0(men_men_n364_), .A1(men_men_n162_), .B0(men_men_n254_), .Y(men_men_n365_));
  NAi41      u0343(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n366_));
  OAI220     u0344(.A0(men_men_n366_), .A1(men_men_n362_), .B0(men_men_n227_), .B1(men_men_n162_), .Y(men_men_n367_));
  AOI210     u0345(.A0(men_men_n366_), .A1(men_men_n162_), .B0(men_men_n160_), .Y(men_men_n368_));
  NOi32      u0346(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n369_));
  NA2        u0347(.A(men_men_n369_), .B(men_men_n46_), .Y(men_men_n370_));
  NO2        u0348(.A(men_men_n370_), .B(i_0_), .Y(men_men_n371_));
  OR3        u0349(.A(men_men_n371_), .B(men_men_n368_), .C(men_men_n367_), .Y(men_men_n372_));
  NO2        u0350(.A(i_1_), .B(men_men_n102_), .Y(men_men_n373_));
  NAi21      u0351(.An(i_3_), .B(i_4_), .Y(men_men_n374_));
  NO2        u0352(.A(men_men_n374_), .B(i_9_), .Y(men_men_n375_));
  AN2        u0353(.A(i_6_), .B(i_7_), .Y(men_men_n376_));
  OAI210     u0354(.A0(men_men_n376_), .A1(men_men_n373_), .B0(men_men_n375_), .Y(men_men_n377_));
  NA2        u0355(.A(i_2_), .B(i_7_), .Y(men_men_n378_));
  NO2        u0356(.A(men_men_n374_), .B(i_10_), .Y(men_men_n379_));
  NA3        u0357(.A(men_men_n379_), .B(men_men_n378_), .C(men_men_n252_), .Y(men_men_n380_));
  AOI210     u0358(.A0(men_men_n380_), .A1(men_men_n377_), .B0(men_men_n190_), .Y(men_men_n381_));
  AOI210     u0359(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n382_));
  OAI210     u0360(.A0(men_men_n382_), .A1(men_men_n193_), .B0(men_men_n379_), .Y(men_men_n383_));
  AOI220     u0361(.A0(men_men_n379_), .A1(men_men_n341_), .B0(men_men_n246_), .B1(men_men_n193_), .Y(men_men_n384_));
  AOI210     u0362(.A0(men_men_n384_), .A1(men_men_n383_), .B0(i_5_), .Y(men_men_n385_));
  NO4        u0363(.A(men_men_n385_), .B(men_men_n381_), .C(men_men_n372_), .D(men_men_n365_), .Y(men_men_n386_));
  NO2        u0364(.A(men_men_n386_), .B(men_men_n360_), .Y(men_men_n387_));
  NO2        u0365(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n388_));
  AN2        u0366(.A(i_12_), .B(i_5_), .Y(men_men_n389_));
  NO2        u0367(.A(i_4_), .B(men_men_n26_), .Y(men_men_n390_));
  NA2        u0368(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n391_));
  NO2        u0369(.A(i_11_), .B(i_6_), .Y(men_men_n392_));
  NA3        u0370(.A(men_men_n392_), .B(men_men_n329_), .C(men_men_n232_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n393_), .B(men_men_n391_), .Y(men_men_n394_));
  NO2        u0372(.A(men_men_n250_), .B(i_5_), .Y(men_men_n395_));
  NO2        u0373(.A(i_5_), .B(i_10_), .Y(men_men_n396_));
  AOI220     u0374(.A0(men_men_n396_), .A1(men_men_n278_), .B0(men_men_n395_), .B1(men_men_n203_), .Y(men_men_n397_));
  NA2        u0375(.A(men_men_n146_), .B(men_men_n45_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n398_), .B(men_men_n397_), .Y(men_men_n399_));
  OAI210     u0377(.A0(men_men_n399_), .A1(men_men_n394_), .B0(men_men_n388_), .Y(men_men_n400_));
  NO2        u0378(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n401_));
  NO2        u0379(.A(men_men_n152_), .B(men_men_n84_), .Y(men_men_n402_));
  OAI210     u0380(.A0(men_men_n402_), .A1(men_men_n394_), .B0(men_men_n401_), .Y(men_men_n403_));
  NO2        u0381(.A(i_11_), .B(i_12_), .Y(men_men_n404_));
  NA2        u0382(.A(men_men_n396_), .B(men_men_n244_), .Y(men_men_n405_));
  NA3        u0383(.A(men_men_n114_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n406_));
  NO2        u0384(.A(men_men_n406_), .B(men_men_n227_), .Y(men_men_n407_));
  NAi21      u0385(.An(i_13_), .B(i_0_), .Y(men_men_n408_));
  NA2        u0386(.A(men_men_n407_), .B(i_0_), .Y(men_men_n409_));
  NA3        u0387(.A(men_men_n409_), .B(men_men_n403_), .C(men_men_n400_), .Y(men_men_n410_));
  NA2        u0388(.A(men_men_n44_), .B(men_men_n232_), .Y(men_men_n411_));
  NO3        u0389(.A(i_1_), .B(i_12_), .C(men_men_n84_), .Y(men_men_n412_));
  NO2        u0390(.A(i_0_), .B(i_11_), .Y(men_men_n413_));
  AN2        u0391(.A(i_1_), .B(i_6_), .Y(men_men_n414_));
  NOi21      u0392(.An(i_2_), .B(i_12_), .Y(men_men_n415_));
  NA2        u0393(.A(men_men_n415_), .B(men_men_n414_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n416_), .B(men_men_n1079_), .Y(men_men_n417_));
  NA2        u0395(.A(men_men_n144_), .B(i_9_), .Y(men_men_n418_));
  NO2        u0396(.A(men_men_n418_), .B(i_4_), .Y(men_men_n419_));
  NA2        u0397(.A(men_men_n417_), .B(men_men_n419_), .Y(men_men_n420_));
  NAi21      u0398(.An(i_9_), .B(i_4_), .Y(men_men_n421_));
  OR2        u0399(.A(i_13_), .B(i_10_), .Y(men_men_n422_));
  NO3        u0400(.A(men_men_n422_), .B(men_men_n119_), .C(men_men_n421_), .Y(men_men_n423_));
  NO2        u0401(.A(men_men_n176_), .B(men_men_n125_), .Y(men_men_n424_));
  OR2        u0402(.A(men_men_n222_), .B(men_men_n221_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n102_), .B(men_men_n25_), .Y(men_men_n426_));
  NA2        u0404(.A(men_men_n290_), .B(men_men_n426_), .Y(men_men_n427_));
  INV        u0405(.A(men_men_n216_), .Y(men_men_n428_));
  OAI220     u0406(.A0(men_men_n428_), .A1(men_men_n425_), .B0(men_men_n427_), .B1(men_men_n345_), .Y(men_men_n429_));
  INV        u0407(.A(men_men_n429_), .Y(men_men_n430_));
  AOI210     u0408(.A0(men_men_n430_), .A1(men_men_n420_), .B0(men_men_n26_), .Y(men_men_n431_));
  NA2        u0409(.A(men_men_n327_), .B(men_men_n326_), .Y(men_men_n432_));
  AOI220     u0410(.A0(men_men_n303_), .A1(men_men_n293_), .B0(men_men_n297_), .B1(i_7_), .Y(men_men_n433_));
  NO2        u0411(.A(men_men_n433_), .B(men_men_n173_), .Y(men_men_n434_));
  NO2        u0412(.A(men_men_n187_), .B(men_men_n84_), .Y(men_men_n435_));
  AOI220     u0413(.A0(men_men_n435_), .A1(men_men_n302_), .B0(men_men_n1084_), .B1(men_men_n216_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n436_), .B(i_7_), .Y(men_men_n437_));
  NO3        u0415(.A(men_men_n437_), .B(men_men_n434_), .C(men_men_n432_), .Y(men_men_n438_));
  NA2        u0416(.A(men_men_n201_), .B(men_men_n97_), .Y(men_men_n439_));
  NA3        u0417(.A(men_men_n329_), .B(men_men_n166_), .C(men_men_n84_), .Y(men_men_n440_));
  AOI210     u0418(.A0(men_men_n440_), .A1(men_men_n439_), .B0(i_8_), .Y(men_men_n441_));
  NA2        u0419(.A(men_men_n198_), .B(i_10_), .Y(men_men_n442_));
  NA3        u0420(.A(men_men_n263_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n303_), .B(men_men_n242_), .Y(men_men_n444_));
  OAI220     u0422(.A0(men_men_n444_), .A1(men_men_n187_), .B0(men_men_n443_), .B1(men_men_n442_), .Y(men_men_n445_));
  NO2        u0423(.A(i_3_), .B(men_men_n48_), .Y(men_men_n446_));
  NA3        u0424(.A(men_men_n341_), .B(men_men_n340_), .C(men_men_n446_), .Y(men_men_n447_));
  NA2        u0425(.A(men_men_n320_), .B(men_men_n325_), .Y(men_men_n448_));
  OAI210     u0426(.A0(men_men_n448_), .A1(men_men_n194_), .B0(men_men_n447_), .Y(men_men_n449_));
  NO3        u0427(.A(men_men_n449_), .B(men_men_n445_), .C(men_men_n441_), .Y(men_men_n450_));
  AOI210     u0428(.A0(men_men_n450_), .A1(men_men_n438_), .B0(men_men_n280_), .Y(men_men_n451_));
  NO4        u0429(.A(men_men_n451_), .B(men_men_n431_), .C(men_men_n410_), .D(men_men_n387_), .Y(men_men_n452_));
  NO2        u0430(.A(men_men_n63_), .B(i_4_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n71_), .B(i_13_), .Y(men_men_n454_));
  NA3        u0432(.A(men_men_n454_), .B(men_men_n453_), .C(i_2_), .Y(men_men_n455_));
  NO2        u0433(.A(i_10_), .B(i_9_), .Y(men_men_n456_));
  NAi21      u0434(.An(i_12_), .B(i_8_), .Y(men_men_n457_));
  NO2        u0435(.A(men_men_n457_), .B(i_3_), .Y(men_men_n458_));
  NA2        u0436(.A(men_men_n458_), .B(men_men_n456_), .Y(men_men_n459_));
  NO2        u0437(.A(men_men_n46_), .B(i_4_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n460_), .B(men_men_n105_), .Y(men_men_n461_));
  OAI220     u0439(.A0(men_men_n461_), .A1(men_men_n210_), .B0(men_men_n459_), .B1(men_men_n455_), .Y(men_men_n462_));
  NA2        u0440(.A(men_men_n315_), .B(i_0_), .Y(men_men_n463_));
  NO3        u0441(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n464_));
  NA2        u0442(.A(men_men_n275_), .B(men_men_n98_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n465_), .B(men_men_n464_), .Y(men_men_n466_));
  NA2        u0444(.A(i_8_), .B(i_9_), .Y(men_men_n467_));
  AOI210     u0445(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n468_));
  OR2        u0446(.A(men_men_n468_), .B(men_men_n467_), .Y(men_men_n469_));
  NA2        u0447(.A(men_men_n290_), .B(men_men_n211_), .Y(men_men_n470_));
  OAI220     u0448(.A0(men_men_n470_), .A1(men_men_n469_), .B0(men_men_n466_), .B1(men_men_n463_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n257_), .B(men_men_n314_), .Y(men_men_n472_));
  NO3        u0450(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n473_));
  INV        u0451(.A(men_men_n473_), .Y(men_men_n474_));
  NA3        u0452(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n475_));
  NA4        u0453(.A(men_men_n147_), .B(men_men_n117_), .C(men_men_n78_), .D(men_men_n23_), .Y(men_men_n476_));
  OAI220     u0454(.A0(men_men_n476_), .A1(men_men_n475_), .B0(men_men_n474_), .B1(men_men_n472_), .Y(men_men_n477_));
  NO3        u0455(.A(men_men_n477_), .B(men_men_n471_), .C(men_men_n462_), .Y(men_men_n478_));
  NA2        u0456(.A(men_men_n302_), .B(men_men_n109_), .Y(men_men_n479_));
  OR2        u0457(.A(men_men_n479_), .B(i_8_), .Y(men_men_n480_));
  OA210      u0458(.A0(men_men_n354_), .A1(men_men_n102_), .B0(men_men_n304_), .Y(men_men_n481_));
  OA220      u0459(.A0(men_men_n481_), .A1(men_men_n165_), .B0(men_men_n480_), .B1(men_men_n239_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n97_), .B(i_13_), .Y(men_men_n483_));
  NA2        u0461(.A(men_men_n435_), .B(men_men_n388_), .Y(men_men_n484_));
  NO2        u0462(.A(i_2_), .B(i_13_), .Y(men_men_n485_));
  NA3        u0463(.A(men_men_n485_), .B(men_men_n164_), .C(men_men_n100_), .Y(men_men_n486_));
  OAI220     u0464(.A0(men_men_n486_), .A1(men_men_n244_), .B0(men_men_n484_), .B1(men_men_n483_), .Y(men_men_n487_));
  NO3        u0465(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n488_));
  NO2        u0466(.A(i_6_), .B(i_7_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n490_));
  NO2        u0468(.A(men_men_n71_), .B(i_3_), .Y(men_men_n491_));
  NOi21      u0469(.An(i_2_), .B(i_7_), .Y(men_men_n492_));
  NAi31      u0470(.An(i_11_), .B(men_men_n492_), .C(men_men_n491_), .Y(men_men_n493_));
  NO2        u0471(.A(men_men_n422_), .B(i_6_), .Y(men_men_n494_));
  NA3        u0472(.A(men_men_n494_), .B(men_men_n453_), .C(men_men_n73_), .Y(men_men_n495_));
  NO2        u0473(.A(men_men_n495_), .B(men_men_n493_), .Y(men_men_n496_));
  NO2        u0474(.A(i_3_), .B(men_men_n198_), .Y(men_men_n497_));
  NO2        u0475(.A(i_6_), .B(i_10_), .Y(men_men_n498_));
  NA3        u0476(.A(men_men_n253_), .B(men_men_n175_), .C(men_men_n134_), .Y(men_men_n499_));
  NA2        u0477(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n500_));
  NO2        u0478(.A(men_men_n160_), .B(i_3_), .Y(men_men_n501_));
  NAi31      u0479(.An(men_men_n500_), .B(men_men_n501_), .C(men_men_n233_), .Y(men_men_n502_));
  NA3        u0480(.A(men_men_n401_), .B(men_men_n183_), .C(men_men_n151_), .Y(men_men_n503_));
  NA3        u0481(.A(men_men_n503_), .B(men_men_n502_), .C(men_men_n499_), .Y(men_men_n504_));
  NO3        u0482(.A(men_men_n504_), .B(men_men_n496_), .C(men_men_n487_), .Y(men_men_n505_));
  NA2        u0483(.A(men_men_n464_), .B(men_men_n389_), .Y(men_men_n506_));
  NA2        u0484(.A(men_men_n473_), .B(men_men_n396_), .Y(men_men_n507_));
  NO2        u0485(.A(men_men_n507_), .B(men_men_n231_), .Y(men_men_n508_));
  NAi21      u0486(.An(men_men_n222_), .B(men_men_n404_), .Y(men_men_n509_));
  NA2        u0487(.A(men_men_n341_), .B(men_men_n224_), .Y(men_men_n510_));
  NO2        u0488(.A(men_men_n26_), .B(i_5_), .Y(men_men_n511_));
  NO2        u0489(.A(i_0_), .B(men_men_n84_), .Y(men_men_n512_));
  NA3        u0490(.A(men_men_n512_), .B(men_men_n511_), .C(men_men_n144_), .Y(men_men_n513_));
  OAI220     u0491(.A0(men_men_n38_), .A1(men_men_n513_), .B0(men_men_n510_), .B1(men_men_n509_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n27_), .B(i_10_), .Y(men_men_n515_));
  NA2        u0493(.A(men_men_n319_), .B(men_men_n246_), .Y(men_men_n516_));
  OAI220     u0494(.A0(men_men_n516_), .A1(men_men_n443_), .B0(men_men_n515_), .B1(men_men_n483_), .Y(men_men_n517_));
  NA4        u0495(.A(men_men_n312_), .B(men_men_n230_), .C(men_men_n71_), .D(men_men_n244_), .Y(men_men_n518_));
  NO2        u0496(.A(men_men_n518_), .B(men_men_n490_), .Y(men_men_n519_));
  NO4        u0497(.A(men_men_n519_), .B(men_men_n517_), .C(men_men_n514_), .D(men_men_n508_), .Y(men_men_n520_));
  NA4        u0498(.A(men_men_n520_), .B(men_men_n505_), .C(men_men_n482_), .D(men_men_n478_), .Y(men_men_n521_));
  NA3        u0499(.A(men_men_n312_), .B(men_men_n180_), .C(men_men_n178_), .Y(men_men_n522_));
  OAI210     u0500(.A0(men_men_n308_), .A1(men_men_n185_), .B0(men_men_n522_), .Y(men_men_n523_));
  AN2        u0501(.A(men_men_n293_), .B(men_men_n241_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n524_), .B(men_men_n523_), .Y(men_men_n525_));
  NA2        u0503(.A(men_men_n319_), .B(men_men_n167_), .Y(men_men_n526_));
  OAI210     u0504(.A0(men_men_n526_), .A1(men_men_n239_), .B0(men_men_n313_), .Y(men_men_n527_));
  NA2        u0505(.A(men_men_n527_), .B(men_men_n328_), .Y(men_men_n528_));
  NA4        u0506(.A(men_men_n454_), .B(men_men_n453_), .C(men_men_n208_), .D(i_2_), .Y(men_men_n529_));
  INV        u0507(.A(men_men_n529_), .Y(men_men_n530_));
  NA2        u0508(.A(men_men_n389_), .B(men_men_n232_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n359_), .B(men_men_n71_), .Y(men_men_n532_));
  NA2        u0510(.A(men_men_n376_), .B(men_men_n369_), .Y(men_men_n533_));
  AO210      u0511(.A0(men_men_n532_), .A1(men_men_n531_), .B0(men_men_n533_), .Y(men_men_n534_));
  NO2        u0512(.A(men_men_n36_), .B(i_8_), .Y(men_men_n535_));
  INV        u0513(.A(men_men_n423_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n536_), .B(men_men_n534_), .Y(men_men_n537_));
  AOI210     u0515(.A0(men_men_n530_), .A1(men_men_n209_), .B0(men_men_n537_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n263_), .B(men_men_n64_), .Y(men_men_n539_));
  OAI210     u0517(.A0(i_8_), .A1(men_men_n539_), .B0(men_men_n136_), .Y(men_men_n540_));
  AOI210     u0518(.A0(men_men_n199_), .A1(i_9_), .B0(men_men_n274_), .Y(men_men_n541_));
  NO2        u0519(.A(men_men_n541_), .B(men_men_n204_), .Y(men_men_n542_));
  AOI220     u0520(.A0(i_6_), .A1(men_men_n542_), .B0(men_men_n540_), .B1(men_men_n424_), .Y(men_men_n543_));
  NA4        u0521(.A(men_men_n543_), .B(men_men_n538_), .C(men_men_n528_), .D(men_men_n525_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n395_), .B(men_men_n302_), .Y(men_men_n545_));
  OAI210     u0523(.A0(men_men_n391_), .A1(men_men_n172_), .B0(men_men_n545_), .Y(men_men_n546_));
  NO2        u0524(.A(i_12_), .B(men_men_n198_), .Y(men_men_n547_));
  NA3        u0525(.A(men_men_n498_), .B(men_men_n178_), .C(men_men_n27_), .Y(men_men_n548_));
  NO3        u0526(.A(men_men_n548_), .B(i_13_), .C(men_men_n479_), .Y(men_men_n549_));
  NOi21      u0527(.An(men_men_n320_), .B(men_men_n38_), .Y(men_men_n550_));
  OAI210     u0528(.A0(men_men_n550_), .A1(men_men_n549_), .B0(men_men_n546_), .Y(men_men_n551_));
  NO2        u0529(.A(i_8_), .B(i_7_), .Y(men_men_n552_));
  OAI210     u0530(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n553_), .B(men_men_n230_), .Y(men_men_n554_));
  AOI220     u0532(.A0(men_men_n329_), .A1(men_men_n39_), .B0(men_men_n242_), .B1(men_men_n212_), .Y(men_men_n555_));
  OAI220     u0533(.A0(men_men_n555_), .A1(i_4_), .B0(men_men_n554_), .B1(men_men_n250_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n44_), .B(i_10_), .Y(men_men_n557_));
  NO2        u0535(.A(men_men_n557_), .B(i_6_), .Y(men_men_n558_));
  NA3        u0536(.A(men_men_n558_), .B(men_men_n556_), .C(men_men_n552_), .Y(men_men_n559_));
  AOI220     u0537(.A0(men_men_n435_), .A1(men_men_n329_), .B0(men_men_n255_), .B1(men_men_n252_), .Y(men_men_n560_));
  OAI220     u0538(.A0(men_men_n560_), .A1(men_men_n271_), .B0(men_men_n483_), .B1(men_men_n135_), .Y(men_men_n561_));
  NA2        u0539(.A(men_men_n561_), .B(men_men_n274_), .Y(men_men_n562_));
  NOi31      u0540(.An(men_men_n297_), .B(men_men_n308_), .C(men_men_n185_), .Y(men_men_n563_));
  NA3        u0541(.A(men_men_n312_), .B(men_men_n178_), .C(men_men_n97_), .Y(men_men_n564_));
  NO2        u0542(.A(men_men_n228_), .B(men_men_n44_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n160_), .B(i_5_), .Y(men_men_n566_));
  NA3        u0544(.A(men_men_n566_), .B(men_men_n411_), .C(men_men_n323_), .Y(men_men_n567_));
  OAI210     u0545(.A0(men_men_n567_), .A1(men_men_n565_), .B0(men_men_n564_), .Y(men_men_n568_));
  OAI210     u0546(.A0(men_men_n568_), .A1(men_men_n563_), .B0(men_men_n473_), .Y(men_men_n569_));
  NA4        u0547(.A(men_men_n569_), .B(men_men_n562_), .C(men_men_n559_), .D(men_men_n551_), .Y(men_men_n570_));
  NA3        u0548(.A(men_men_n224_), .B(men_men_n69_), .C(men_men_n44_), .Y(men_men_n571_));
  NA2        u0549(.A(men_men_n290_), .B(men_men_n82_), .Y(men_men_n572_));
  AOI210     u0550(.A0(men_men_n571_), .A1(men_men_n349_), .B0(men_men_n572_), .Y(men_men_n573_));
  NA2        u0551(.A(men_men_n303_), .B(men_men_n293_), .Y(men_men_n574_));
  NO2        u0552(.A(men_men_n574_), .B(men_men_n177_), .Y(men_men_n575_));
  NA2        u0553(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n576_));
  NA2        u0554(.A(men_men_n456_), .B(men_men_n228_), .Y(men_men_n577_));
  NO2        u0555(.A(men_men_n576_), .B(men_men_n577_), .Y(men_men_n578_));
  NA2        u0556(.A(i_0_), .B(men_men_n48_), .Y(men_men_n579_));
  NA3        u0557(.A(men_men_n547_), .B(men_men_n283_), .C(men_men_n579_), .Y(men_men_n580_));
  INV        u0558(.A(men_men_n580_), .Y(men_men_n581_));
  NO4        u0559(.A(men_men_n581_), .B(men_men_n578_), .C(men_men_n575_), .D(men_men_n573_), .Y(men_men_n582_));
  NO4        u0560(.A(men_men_n258_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n583_));
  NO3        u0561(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n584_));
  NO2        u0562(.A(men_men_n240_), .B(men_men_n36_), .Y(men_men_n585_));
  AN2        u0563(.A(men_men_n585_), .B(men_men_n584_), .Y(men_men_n586_));
  OA210      u0564(.A0(men_men_n586_), .A1(men_men_n583_), .B0(men_men_n359_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n422_), .B(i_1_), .Y(men_men_n588_));
  NOi31      u0566(.An(men_men_n588_), .B(men_men_n465_), .C(men_men_n71_), .Y(men_men_n589_));
  AN3        u0567(.A(men_men_n589_), .B(men_men_n419_), .C(i_2_), .Y(men_men_n590_));
  NO2        u0568(.A(men_men_n433_), .B(men_men_n181_), .Y(men_men_n591_));
  NO3        u0569(.A(men_men_n591_), .B(men_men_n590_), .C(men_men_n587_), .Y(men_men_n592_));
  NOi21      u0570(.An(i_10_), .B(i_6_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n84_), .B(men_men_n25_), .Y(men_men_n594_));
  AOI220     u0572(.A0(men_men_n290_), .A1(men_men_n594_), .B0(men_men_n283_), .B1(men_men_n593_), .Y(men_men_n595_));
  NO2        u0573(.A(men_men_n595_), .B(men_men_n463_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n116_), .B(men_men_n23_), .Y(men_men_n597_));
  NA2        u0575(.A(men_men_n320_), .B(men_men_n167_), .Y(men_men_n598_));
  AOI220     u0576(.A0(men_men_n598_), .A1(men_men_n444_), .B0(men_men_n188_), .B1(men_men_n186_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n203_), .B(men_men_n37_), .Y(men_men_n600_));
  NOi31      u0578(.An(men_men_n148_), .B(men_men_n600_), .C(men_men_n337_), .Y(men_men_n601_));
  NO3        u0579(.A(men_men_n601_), .B(men_men_n599_), .C(men_men_n596_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n532_), .B(men_men_n384_), .Y(men_men_n603_));
  INV        u0581(.A(men_men_n323_), .Y(men_men_n604_));
  NO2        u0582(.A(i_12_), .B(men_men_n84_), .Y(men_men_n605_));
  NA3        u0583(.A(men_men_n392_), .B(men_men_n290_), .C(men_men_n224_), .Y(men_men_n606_));
  NO2        u0584(.A(men_men_n606_), .B(men_men_n604_), .Y(men_men_n607_));
  NA2        u0585(.A(men_men_n178_), .B(i_0_), .Y(men_men_n608_));
  NO3        u0586(.A(men_men_n608_), .B(men_men_n1081_), .C(men_men_n308_), .Y(men_men_n609_));
  OR2        u0587(.A(i_2_), .B(i_5_), .Y(men_men_n610_));
  OR2        u0588(.A(men_men_n610_), .B(men_men_n414_), .Y(men_men_n611_));
  NO2        u0589(.A(men_men_n252_), .B(men_men_n203_), .Y(men_men_n612_));
  AOI210     u0590(.A0(men_men_n612_), .A1(men_men_n611_), .B0(men_men_n509_), .Y(men_men_n613_));
  NO4        u0591(.A(men_men_n613_), .B(men_men_n609_), .C(men_men_n607_), .D(men_men_n603_), .Y(men_men_n614_));
  NA4        u0592(.A(men_men_n614_), .B(men_men_n602_), .C(men_men_n592_), .D(men_men_n582_), .Y(men_men_n615_));
  NO4        u0593(.A(men_men_n615_), .B(men_men_n570_), .C(men_men_n544_), .D(men_men_n521_), .Y(men_men_n616_));
  NA4        u0594(.A(men_men_n616_), .B(men_men_n452_), .C(men_men_n358_), .D(men_men_n318_), .Y(men7));
  NO2        u0595(.A(men_men_n93_), .B(men_men_n54_), .Y(men_men_n618_));
  NO2        u0596(.A(men_men_n109_), .B(men_men_n90_), .Y(men_men_n619_));
  NA2        u0597(.A(men_men_n390_), .B(men_men_n619_), .Y(men_men_n620_));
  NA2        u0598(.A(men_men_n498_), .B(men_men_n82_), .Y(men_men_n621_));
  NA2        u0599(.A(i_11_), .B(men_men_n198_), .Y(men_men_n622_));
  INV        u0600(.A(men_men_n620_), .Y(men_men_n623_));
  NA3        u0601(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n624_));
  NO2        u0602(.A(men_men_n244_), .B(i_4_), .Y(men_men_n625_));
  NA2        u0603(.A(men_men_n625_), .B(i_8_), .Y(men_men_n626_));
  AOI210     u0604(.A0(men_men_n626_), .A1(men_men_n106_), .B0(men_men_n624_), .Y(men_men_n627_));
  NA2        u0605(.A(i_2_), .B(men_men_n84_), .Y(men_men_n628_));
  OAI210     u0606(.A0(men_men_n87_), .A1(men_men_n208_), .B0(men_men_n209_), .Y(men_men_n629_));
  NO2        u0607(.A(i_7_), .B(men_men_n37_), .Y(men_men_n630_));
  NA2        u0608(.A(i_4_), .B(i_8_), .Y(men_men_n631_));
  NO2        u0609(.A(men_men_n312_), .B(men_men_n630_), .Y(men_men_n632_));
  OAI220     u0610(.A0(men_men_n632_), .A1(men_men_n628_), .B0(men_men_n629_), .B1(i_13_), .Y(men_men_n633_));
  NO4        u0611(.A(men_men_n633_), .B(men_men_n627_), .C(men_men_n623_), .D(men_men_n618_), .Y(men_men_n634_));
  AOI210     u0612(.A0(men_men_n130_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n635_));
  AOI210     u0613(.A0(men_men_n635_), .A1(men_men_n244_), .B0(men_men_n164_), .Y(men_men_n636_));
  OR2        u0614(.A(i_6_), .B(i_10_), .Y(men_men_n637_));
  NO2        u0615(.A(men_men_n637_), .B(men_men_n23_), .Y(men_men_n638_));
  OR3        u0616(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n639_));
  NO3        u0617(.A(men_men_n639_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n640_));
  INV        u0618(.A(men_men_n205_), .Y(men_men_n641_));
  NO2        u0619(.A(men_men_n640_), .B(men_men_n638_), .Y(men_men_n642_));
  OA220      u0620(.A0(men_men_n642_), .A1(men_men_n604_), .B0(men_men_n636_), .B1(men_men_n276_), .Y(men_men_n643_));
  AOI210     u0621(.A0(men_men_n643_), .A1(men_men_n634_), .B0(men_men_n63_), .Y(men_men_n644_));
  NOi21      u0622(.An(i_11_), .B(i_7_), .Y(men_men_n645_));
  AO210      u0623(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n646_), .B(men_men_n645_), .Y(men_men_n647_));
  NA2        u0625(.A(men_men_n647_), .B(men_men_n212_), .Y(men_men_n648_));
  NA3        u0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n649_));
  NAi21      u0627(.An(men_men_n649_), .B(i_11_), .Y(men_men_n650_));
  AOI210     u0628(.A0(men_men_n650_), .A1(men_men_n648_), .B0(men_men_n63_), .Y(men_men_n651_));
  NA2        u0629(.A(men_men_n86_), .B(men_men_n63_), .Y(men_men_n652_));
  AO210      u0630(.A0(men_men_n652_), .A1(men_men_n384_), .B0(men_men_n40_), .Y(men_men_n653_));
  NO3        u0631(.A(men_men_n265_), .B(men_men_n213_), .C(men_men_n622_), .Y(men_men_n654_));
  OAI210     u0632(.A0(men_men_n654_), .A1(men_men_n233_), .B0(men_men_n63_), .Y(men_men_n655_));
  NA2        u0633(.A(men_men_n415_), .B(men_men_n31_), .Y(men_men_n656_));
  OR2        u0634(.A(men_men_n213_), .B(men_men_n109_), .Y(men_men_n657_));
  NA2        u0635(.A(men_men_n657_), .B(men_men_n656_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n63_), .B(i_9_), .Y(men_men_n659_));
  NO2        u0637(.A(men_men_n659_), .B(i_4_), .Y(men_men_n660_));
  NA2        u0638(.A(men_men_n660_), .B(men_men_n658_), .Y(men_men_n661_));
  NO2        u0639(.A(i_1_), .B(i_12_), .Y(men_men_n662_));
  NA3        u0640(.A(men_men_n662_), .B(men_men_n111_), .C(men_men_n24_), .Y(men_men_n663_));
  NA4        u0641(.A(men_men_n663_), .B(men_men_n661_), .C(men_men_n655_), .D(men_men_n653_), .Y(men_men_n664_));
  OAI210     u0642(.A0(men_men_n664_), .A1(men_men_n651_), .B0(i_6_), .Y(men_men_n665_));
  OAI210     u0643(.A0(men_men_n649_), .A1(men_men_n109_), .B0(men_men_n475_), .Y(men_men_n666_));
  NA2        u0644(.A(men_men_n666_), .B(men_men_n605_), .Y(men_men_n667_));
  NO2        u0645(.A(i_6_), .B(i_11_), .Y(men_men_n668_));
  NA2        u0646(.A(men_men_n667_), .B(men_men_n466_), .Y(men_men_n669_));
  NO4        u0647(.A(men_men_n221_), .B(men_men_n130_), .C(i_13_), .D(men_men_n84_), .Y(men_men_n670_));
  NA2        u0648(.A(men_men_n670_), .B(men_men_n659_), .Y(men_men_n671_));
  NO3        u0649(.A(men_men_n637_), .B(men_men_n240_), .C(men_men_n23_), .Y(men_men_n672_));
  AOI210     u0650(.A0(i_1_), .A1(men_men_n266_), .B0(men_men_n672_), .Y(men_men_n673_));
  OAI210     u0651(.A0(men_men_n673_), .A1(men_men_n44_), .B0(men_men_n671_), .Y(men_men_n674_));
  NA3        u0652(.A(men_men_n552_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n675_));
  NA2        u0653(.A(men_men_n140_), .B(i_9_), .Y(men_men_n676_));
  NA3        u0654(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n677_));
  NO2        u0655(.A(men_men_n46_), .B(i_1_), .Y(men_men_n678_));
  NA3        u0656(.A(men_men_n678_), .B(men_men_n275_), .C(men_men_n44_), .Y(men_men_n679_));
  OAI220     u0657(.A0(men_men_n679_), .A1(men_men_n677_), .B0(men_men_n676_), .B1(men_men_n1078_), .Y(men_men_n680_));
  NA3        u0658(.A(men_men_n659_), .B(men_men_n323_), .C(i_6_), .Y(men_men_n681_));
  NAi21      u0659(.An(men_men_n675_), .B(men_men_n92_), .Y(men_men_n682_));
  NA2        u0660(.A(men_men_n678_), .B(men_men_n275_), .Y(men_men_n683_));
  NO2        u0661(.A(i_11_), .B(men_men_n37_), .Y(men_men_n684_));
  NA2        u0662(.A(men_men_n684_), .B(men_men_n24_), .Y(men_men_n685_));
  OAI210     u0663(.A0(men_men_n685_), .A1(men_men_n683_), .B0(men_men_n682_), .Y(men_men_n686_));
  OR2        u0664(.A(men_men_n686_), .B(men_men_n680_), .Y(men_men_n687_));
  NO3        u0665(.A(men_men_n687_), .B(men_men_n674_), .C(men_men_n669_), .Y(men_men_n688_));
  NO2        u0666(.A(men_men_n244_), .B(men_men_n102_), .Y(men_men_n689_));
  NO2        u0667(.A(men_men_n689_), .B(men_men_n645_), .Y(men_men_n690_));
  NO2        u0668(.A(men_men_n421_), .B(men_men_n84_), .Y(men_men_n691_));
  NA2        u0669(.A(i_3_), .B(men_men_n198_), .Y(men_men_n692_));
  NO2        u0670(.A(men_men_n692_), .B(men_men_n116_), .Y(men_men_n693_));
  AN2        u0671(.A(men_men_n693_), .B(men_men_n558_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n240_), .B(men_men_n44_), .Y(men_men_n695_));
  NO3        u0673(.A(men_men_n695_), .B(men_men_n315_), .C(men_men_n245_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n119_), .B(men_men_n37_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n697_), .B(i_6_), .Y(men_men_n698_));
  NO2        u0676(.A(men_men_n84_), .B(i_9_), .Y(men_men_n699_));
  NO2        u0677(.A(men_men_n699_), .B(men_men_n63_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n700_), .B(men_men_n662_), .Y(men_men_n701_));
  NO4        u0679(.A(men_men_n701_), .B(men_men_n698_), .C(men_men_n696_), .D(i_4_), .Y(men_men_n702_));
  NA2        u0680(.A(i_1_), .B(i_3_), .Y(men_men_n703_));
  NO2        u0681(.A(men_men_n467_), .B(men_men_n93_), .Y(men_men_n704_));
  AOI210     u0682(.A0(men_men_n695_), .A1(men_men_n593_), .B0(men_men_n704_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(men_men_n703_), .Y(men_men_n706_));
  NO3        u0684(.A(men_men_n706_), .B(men_men_n702_), .C(men_men_n694_), .Y(men_men_n707_));
  NA3        u0685(.A(men_men_n707_), .B(men_men_n688_), .C(men_men_n665_), .Y(men_men_n708_));
  NO3        u0686(.A(i_11_), .B(i_3_), .C(i_7_), .Y(men_men_n709_));
  NOi21      u0687(.An(men_men_n709_), .B(i_10_), .Y(men_men_n710_));
  OA210      u0688(.A0(men_men_n710_), .A1(men_men_n253_), .B0(men_men_n84_), .Y(men_men_n711_));
  NA2        u0689(.A(men_men_n376_), .B(men_men_n375_), .Y(men_men_n712_));
  NA3        u0690(.A(men_men_n498_), .B(men_men_n535_), .C(men_men_n46_), .Y(men_men_n713_));
  NO3        u0691(.A(men_men_n492_), .B(men_men_n631_), .C(men_men_n84_), .Y(men_men_n714_));
  NA2        u0692(.A(men_men_n714_), .B(men_men_n25_), .Y(men_men_n715_));
  NA3        u0693(.A(men_men_n715_), .B(men_men_n713_), .C(men_men_n712_), .Y(men_men_n716_));
  OAI210     u0694(.A0(men_men_n716_), .A1(men_men_n711_), .B0(i_1_), .Y(men_men_n717_));
  INV        u0695(.A(i_1_), .Y(men_men_n718_));
  NO2        u0696(.A(men_men_n374_), .B(i_2_), .Y(men_men_n719_));
  AOI210     u0697(.A0(men_men_n681_), .A1(men_men_n717_), .B0(i_13_), .Y(men_men_n720_));
  OR2        u0698(.A(i_11_), .B(i_7_), .Y(men_men_n721_));
  NA2        u0699(.A(men_men_n107_), .B(men_men_n140_), .Y(men_men_n722_));
  AOI220     u0700(.A0(men_men_n485_), .A1(men_men_n164_), .B0(men_men_n460_), .B1(men_men_n140_), .Y(men_men_n723_));
  OAI210     u0701(.A0(men_men_n723_), .A1(men_men_n44_), .B0(men_men_n722_), .Y(men_men_n724_));
  NO2        u0702(.A(men_men_n492_), .B(men_men_n24_), .Y(men_men_n725_));
  AOI220     u0703(.A0(men_men_n725_), .A1(men_men_n691_), .B0(men_men_n253_), .B1(men_men_n133_), .Y(men_men_n726_));
  NO2        u0704(.A(men_men_n726_), .B(men_men_n40_), .Y(men_men_n727_));
  AOI210     u0705(.A0(men_men_n724_), .A1(men_men_n339_), .B0(men_men_n727_), .Y(men_men_n728_));
  AOI220     u0706(.A0(i_7_), .A1(men_men_n70_), .B0(men_men_n392_), .B1(men_men_n678_), .Y(men_men_n729_));
  NO2        u0707(.A(men_men_n729_), .B(men_men_n250_), .Y(men_men_n730_));
  AOI210     u0708(.A0(men_men_n457_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n731_));
  NOi31      u0709(.An(men_men_n731_), .B(men_men_n621_), .C(men_men_n44_), .Y(men_men_n732_));
  NA2        u0710(.A(men_men_n129_), .B(i_13_), .Y(men_men_n733_));
  NO2        u0711(.A(men_men_n677_), .B(men_men_n116_), .Y(men_men_n734_));
  INV        u0712(.A(men_men_n734_), .Y(men_men_n735_));
  OAI220     u0713(.A0(men_men_n735_), .A1(men_men_n69_), .B0(men_men_n733_), .B1(men_men_n718_), .Y(men_men_n736_));
  NO3        u0714(.A(men_men_n69_), .B(men_men_n32_), .C(men_men_n102_), .Y(men_men_n737_));
  NA2        u0715(.A(men_men_n26_), .B(men_men_n198_), .Y(men_men_n738_));
  INV        u0716(.A(i_7_), .Y(men_men_n739_));
  INV        u0717(.A(men_men_n737_), .Y(men_men_n740_));
  AOI220     u0718(.A0(men_men_n392_), .A1(men_men_n678_), .B0(men_men_n92_), .B1(men_men_n103_), .Y(men_men_n741_));
  OAI220     u0719(.A0(men_men_n741_), .A1(men_men_n626_), .B0(men_men_n740_), .B1(men_men_n641_), .Y(men_men_n742_));
  NO4        u0720(.A(men_men_n742_), .B(men_men_n736_), .C(men_men_n732_), .D(men_men_n730_), .Y(men_men_n743_));
  OR2        u0721(.A(i_11_), .B(i_6_), .Y(men_men_n744_));
  NO2        u0722(.A(men_men_n735_), .B(men_men_n744_), .Y(men_men_n745_));
  NA2        u0723(.A(men_men_n668_), .B(i_13_), .Y(men_men_n746_));
  NA2        u0724(.A(men_men_n103_), .B(men_men_n738_), .Y(men_men_n747_));
  NAi21      u0725(.An(i_11_), .B(i_12_), .Y(men_men_n748_));
  NO3        u0726(.A(men_men_n748_), .B(i_13_), .C(men_men_n84_), .Y(men_men_n749_));
  NO3        u0727(.A(men_men_n492_), .B(men_men_n605_), .C(men_men_n631_), .Y(men_men_n750_));
  AOI220     u0728(.A0(men_men_n750_), .A1(men_men_n319_), .B0(men_men_n749_), .B1(men_men_n747_), .Y(men_men_n751_));
  NA2        u0729(.A(men_men_n751_), .B(men_men_n746_), .Y(men_men_n752_));
  OAI210     u0730(.A0(men_men_n752_), .A1(men_men_n745_), .B0(men_men_n63_), .Y(men_men_n753_));
  NO2        u0731(.A(i_2_), .B(i_12_), .Y(men_men_n754_));
  OAI210     u0732(.A0(men_men_n635_), .A1(men_men_n373_), .B0(men_men_n754_), .Y(men_men_n755_));
  NA2        u0733(.A(i_8_), .B(men_men_n25_), .Y(men_men_n756_));
  NO3        u0734(.A(men_men_n756_), .B(men_men_n390_), .C(men_men_n625_), .Y(men_men_n757_));
  OAI210     u0735(.A0(men_men_n757_), .A1(men_men_n375_), .B0(men_men_n373_), .Y(men_men_n758_));
  NO2        u0736(.A(men_men_n130_), .B(i_2_), .Y(men_men_n759_));
  NA2        u0737(.A(men_men_n759_), .B(men_men_n662_), .Y(men_men_n760_));
  NA3        u0738(.A(men_men_n760_), .B(men_men_n758_), .C(men_men_n755_), .Y(men_men_n761_));
  NA3        u0739(.A(men_men_n761_), .B(men_men_n45_), .C(men_men_n232_), .Y(men_men_n762_));
  NA4        u0740(.A(men_men_n762_), .B(men_men_n753_), .C(men_men_n743_), .D(men_men_n728_), .Y(men_men_n763_));
  OR4        u0741(.A(men_men_n763_), .B(men_men_n720_), .C(men_men_n708_), .D(men_men_n644_), .Y(men5));
  AOI210     u0742(.A0(men_men_n690_), .A1(men_men_n278_), .B0(men_men_n424_), .Y(men_men_n765_));
  AO210      u0743(.A0(men_men_n24_), .A1(i_10_), .B0(men_men_n257_), .Y(men_men_n766_));
  NA3        u0744(.A(men_men_n766_), .B(men_men_n754_), .C(men_men_n109_), .Y(men_men_n767_));
  NA2        u0745(.A(men_men_n767_), .B(men_men_n765_), .Y(men_men_n768_));
  NO3        u0746(.A(i_11_), .B(men_men_n244_), .C(i_13_), .Y(men_men_n769_));
  NO2        u0747(.A(men_men_n126_), .B(men_men_n23_), .Y(men_men_n770_));
  NA2        u0748(.A(i_12_), .B(i_8_), .Y(men_men_n771_));
  INV        u0749(.A(men_men_n456_), .Y(men_men_n772_));
  AOI220     u0750(.A0(men_men_n323_), .A1(men_men_n597_), .B0(i_12_), .B1(men_men_n770_), .Y(men_men_n773_));
  INV        u0751(.A(men_men_n773_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n774_), .B(men_men_n768_), .Y(men_men_n775_));
  INV        u0753(.A(men_men_n175_), .Y(men_men_n776_));
  INV        u0754(.A(men_men_n253_), .Y(men_men_n777_));
  OAI210     u0755(.A0(men_men_n719_), .A1(men_men_n458_), .B0(men_men_n112_), .Y(men_men_n778_));
  AOI210     u0756(.A0(men_men_n778_), .A1(men_men_n777_), .B0(men_men_n776_), .Y(men_men_n779_));
  NO2        u0757(.A(men_men_n467_), .B(men_men_n26_), .Y(men_men_n780_));
  NO2        u0758(.A(men_men_n780_), .B(men_men_n426_), .Y(men_men_n781_));
  NA2        u0759(.A(men_men_n781_), .B(i_2_), .Y(men_men_n782_));
  INV        u0760(.A(men_men_n782_), .Y(men_men_n783_));
  AOI210     u0761(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n422_), .Y(men_men_n784_));
  AOI210     u0762(.A0(men_men_n784_), .A1(men_men_n783_), .B0(men_men_n779_), .Y(men_men_n785_));
  NO2        u0763(.A(men_men_n195_), .B(men_men_n127_), .Y(men_men_n786_));
  OAI210     u0764(.A0(men_men_n786_), .A1(men_men_n770_), .B0(i_2_), .Y(men_men_n787_));
  INV        u0765(.A(men_men_n176_), .Y(men_men_n788_));
  NO3        u0766(.A(men_men_n646_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n789_));
  AOI210     u0767(.A0(men_men_n788_), .A1(men_men_n87_), .B0(men_men_n789_), .Y(men_men_n790_));
  AOI210     u0768(.A0(men_men_n790_), .A1(men_men_n787_), .B0(men_men_n198_), .Y(men_men_n791_));
  OA210      u0769(.A0(men_men_n647_), .A1(men_men_n128_), .B0(i_13_), .Y(men_men_n792_));
  NA2        u0770(.A(men_men_n205_), .B(men_men_n208_), .Y(men_men_n793_));
  INV        u0771(.A(men_men_n154_), .Y(men_men_n794_));
  AOI210     u0772(.A0(men_men_n794_), .A1(men_men_n793_), .B0(men_men_n378_), .Y(men_men_n795_));
  AOI210     u0773(.A0(men_men_n213_), .A1(men_men_n150_), .B0(men_men_n535_), .Y(men_men_n796_));
  NA2        u0774(.A(men_men_n796_), .B(men_men_n426_), .Y(men_men_n797_));
  NA3        u0775(.A(men_men_n312_), .B(men_men_n126_), .C(men_men_n42_), .Y(men_men_n798_));
  OAI210     u0776(.A0(men_men_n798_), .A1(men_men_n46_), .B0(men_men_n797_), .Y(men_men_n799_));
  NO4        u0777(.A(men_men_n799_), .B(men_men_n795_), .C(men_men_n792_), .D(men_men_n791_), .Y(men_men_n800_));
  NO2        u0778(.A(men_men_n62_), .B(i_12_), .Y(men_men_n801_));
  NO2        u0779(.A(men_men_n801_), .B(men_men_n128_), .Y(men_men_n802_));
  NO2        u0780(.A(men_men_n802_), .B(men_men_n622_), .Y(men_men_n803_));
  NA2        u0781(.A(men_men_n803_), .B(men_men_n36_), .Y(men_men_n804_));
  NA4        u0782(.A(men_men_n804_), .B(men_men_n800_), .C(men_men_n785_), .D(men_men_n775_), .Y(men6));
  NA2        u0783(.A(men_men_n25_), .B(men_men_n759_), .Y(men_men_n806_));
  NA4        u0784(.A(men_men_n396_), .B(men_men_n497_), .C(men_men_n69_), .D(men_men_n102_), .Y(men_men_n807_));
  INV        u0785(.A(men_men_n807_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n227_), .B(men_men_n500_), .Y(men_men_n809_));
  NO2        u0787(.A(i_11_), .B(i_9_), .Y(men_men_n810_));
  NO2        u0788(.A(men_men_n808_), .B(men_men_n334_), .Y(men_men_n811_));
  AO210      u0789(.A0(men_men_n811_), .A1(men_men_n806_), .B0(i_12_), .Y(men_men_n812_));
  NA2        u0790(.A(men_men_n379_), .B(men_men_n341_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n605_), .B(men_men_n63_), .Y(men_men_n814_));
  NA2        u0792(.A(men_men_n710_), .B(men_men_n69_), .Y(men_men_n815_));
  NA4        u0793(.A(men_men_n652_), .B(men_men_n815_), .C(men_men_n814_), .D(men_men_n813_), .Y(men_men_n816_));
  INV        u0794(.A(men_men_n202_), .Y(men_men_n817_));
  AOI220     u0795(.A0(men_men_n817_), .A1(men_men_n810_), .B0(men_men_n816_), .B1(men_men_n71_), .Y(men_men_n818_));
  INV        u0796(.A(men_men_n333_), .Y(men_men_n819_));
  NA2        u0797(.A(men_men_n73_), .B(men_men_n133_), .Y(men_men_n820_));
  INV        u0798(.A(men_men_n126_), .Y(men_men_n821_));
  NA2        u0799(.A(men_men_n821_), .B(men_men_n46_), .Y(men_men_n822_));
  AOI210     u0800(.A0(men_men_n822_), .A1(men_men_n820_), .B0(men_men_n819_), .Y(men_men_n823_));
  NA2        u0801(.A(men_men_n1083_), .B(men_men_n801_), .Y(men_men_n824_));
  AOI210     u0802(.A0(men_men_n824_), .A1(men_men_n533_), .B0(men_men_n190_), .Y(men_men_n825_));
  NO2        u0803(.A(men_men_n32_), .B(i_11_), .Y(men_men_n826_));
  NA3        u0804(.A(men_men_n826_), .B(men_men_n489_), .C(men_men_n396_), .Y(men_men_n827_));
  OAI210     u0805(.A0(men_men_n709_), .A1(men_men_n585_), .B0(men_men_n584_), .Y(men_men_n828_));
  NA2        u0806(.A(men_men_n828_), .B(men_men_n827_), .Y(men_men_n829_));
  OR3        u0807(.A(men_men_n829_), .B(men_men_n825_), .C(men_men_n823_), .Y(men_men_n830_));
  NO2        u0808(.A(men_men_n721_), .B(i_2_), .Y(men_men_n831_));
  NA2        u0809(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n832_));
  OAI210     u0810(.A0(men_men_n832_), .A1(men_men_n414_), .B0(men_men_n364_), .Y(men_men_n833_));
  NA2        u0811(.A(men_men_n833_), .B(men_men_n831_), .Y(men_men_n834_));
  NA3        u0812(.A(men_men_n353_), .B(men_men_n262_), .C(i_7_), .Y(men_men_n835_));
  BUFFER     u0813(.A(men_men_n458_), .Y(men_men_n836_));
  NA3        u0814(.A(men_men_n836_), .B(men_men_n149_), .C(men_men_n68_), .Y(men_men_n837_));
  AO210      u0815(.A0(men_men_n507_), .A1(men_men_n772_), .B0(men_men_n36_), .Y(men_men_n838_));
  NA4        u0816(.A(men_men_n838_), .B(men_men_n837_), .C(men_men_n835_), .D(men_men_n834_), .Y(men_men_n839_));
  OAI210     u0817(.A0(i_6_), .A1(i_11_), .B0(men_men_n85_), .Y(men_men_n840_));
  AOI220     u0818(.A0(men_men_n840_), .A1(men_men_n584_), .B0(men_men_n809_), .B1(men_men_n739_), .Y(men_men_n841_));
  NA3        u0819(.A(men_men_n378_), .B(men_men_n246_), .C(men_men_n149_), .Y(men_men_n842_));
  NA3        u0820(.A(men_men_n842_), .B(men_men_n841_), .C(men_men_n629_), .Y(men_men_n843_));
  AO210      u0821(.A0(men_men_n535_), .A1(men_men_n46_), .B0(men_men_n86_), .Y(men_men_n844_));
  NA3        u0822(.A(men_men_n844_), .B(men_men_n498_), .C(men_men_n224_), .Y(men_men_n845_));
  INV        u0823(.A(men_men_n583_), .Y(men_men_n846_));
  NO2        u0824(.A(men_men_n637_), .B(men_men_n103_), .Y(men_men_n847_));
  OAI210     u0825(.A0(men_men_n847_), .A1(men_men_n113_), .B0(men_men_n413_), .Y(men_men_n848_));
  INV        u0826(.A(men_men_n611_), .Y(men_men_n849_));
  NA3        u0827(.A(men_men_n849_), .B(men_men_n333_), .C(i_7_), .Y(men_men_n850_));
  NA4        u0828(.A(men_men_n850_), .B(men_men_n848_), .C(men_men_n846_), .D(men_men_n845_), .Y(men_men_n851_));
  NO4        u0829(.A(men_men_n851_), .B(men_men_n843_), .C(men_men_n839_), .D(men_men_n830_), .Y(men_men_n852_));
  NA4        u0830(.A(men_men_n852_), .B(men_men_n818_), .C(men_men_n812_), .D(men_men_n386_), .Y(men3));
  NA2        u0831(.A(i_6_), .B(i_7_), .Y(men_men_n854_));
  NO2        u0832(.A(men_men_n854_), .B(i_0_), .Y(men_men_n855_));
  NO2        u0833(.A(i_11_), .B(men_men_n244_), .Y(men_men_n856_));
  OAI210     u0834(.A0(men_men_n855_), .A1(men_men_n297_), .B0(men_men_n856_), .Y(men_men_n857_));
  NO2        u0835(.A(men_men_n857_), .B(men_men_n198_), .Y(men_men_n858_));
  NO3        u0836(.A(men_men_n463_), .B(men_men_n90_), .C(men_men_n44_), .Y(men_men_n859_));
  OA210      u0837(.A0(men_men_n859_), .A1(men_men_n858_), .B0(men_men_n178_), .Y(men_men_n860_));
  NA3        u0838(.A(men_men_n842_), .B(men_men_n629_), .C(men_men_n377_), .Y(men_men_n861_));
  NA2        u0839(.A(men_men_n861_), .B(men_men_n39_), .Y(men_men_n862_));
  NOi21      u0840(.An(men_men_n97_), .B(men_men_n781_), .Y(men_men_n863_));
  NO3        u0841(.A(men_men_n657_), .B(men_men_n467_), .C(men_men_n133_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n415_), .B(men_men_n45_), .Y(men_men_n865_));
  AN2        u0843(.A(men_men_n465_), .B(men_men_n55_), .Y(men_men_n866_));
  NO3        u0844(.A(men_men_n866_), .B(men_men_n864_), .C(men_men_n863_), .Y(men_men_n867_));
  AOI210     u0845(.A0(men_men_n867_), .A1(men_men_n862_), .B0(men_men_n48_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n731_), .B(men_men_n699_), .Y(men_men_n869_));
  NA2        u0847(.A(i_0_), .B(men_men_n446_), .Y(men_men_n870_));
  NO2        u0848(.A(men_men_n870_), .B(men_men_n869_), .Y(men_men_n871_));
  NOi21      u0849(.An(i_5_), .B(i_9_), .Y(men_men_n872_));
  NA2        u0850(.A(men_men_n872_), .B(men_men_n454_), .Y(men_men_n873_));
  INV        u0851(.A(men_men_n714_), .Y(men_men_n874_));
  NO3        u0852(.A(men_men_n418_), .B(men_men_n275_), .C(men_men_n71_), .Y(men_men_n875_));
  NO2        u0853(.A(men_men_n179_), .B(men_men_n150_), .Y(men_men_n876_));
  AOI210     u0854(.A0(men_men_n876_), .A1(men_men_n252_), .B0(men_men_n875_), .Y(men_men_n877_));
  OAI220     u0855(.A0(men_men_n877_), .A1(men_men_n185_), .B0(men_men_n874_), .B1(men_men_n873_), .Y(men_men_n878_));
  NO4        u0856(.A(men_men_n878_), .B(men_men_n871_), .C(men_men_n868_), .D(men_men_n860_), .Y(men_men_n879_));
  NA2        u0857(.A(men_men_n190_), .B(men_men_n24_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n697_), .B(men_men_n619_), .Y(men_men_n881_));
  NO2        u0859(.A(men_men_n881_), .B(men_men_n880_), .Y(men_men_n882_));
  NA2        u0860(.A(men_men_n319_), .B(men_men_n131_), .Y(men_men_n883_));
  NAi21      u0861(.An(men_men_n165_), .B(men_men_n446_), .Y(men_men_n884_));
  OAI220     u0862(.A0(men_men_n884_), .A1(i_2_), .B0(men_men_n883_), .B1(men_men_n405_), .Y(men_men_n885_));
  NO2        u0863(.A(men_men_n885_), .B(men_men_n882_), .Y(men_men_n886_));
  NO2        u0864(.A(men_men_n396_), .B(men_men_n301_), .Y(men_men_n887_));
  NA2        u0865(.A(men_men_n887_), .B(men_men_n734_), .Y(men_men_n888_));
  NA2        u0866(.A(men_men_n594_), .B(i_0_), .Y(men_men_n889_));
  NO3        u0867(.A(men_men_n889_), .B(men_men_n391_), .C(men_men_n87_), .Y(men_men_n890_));
  NO4        u0868(.A(men_men_n610_), .B(men_men_n221_), .C(men_men_n422_), .D(men_men_n414_), .Y(men_men_n891_));
  AOI210     u0869(.A0(men_men_n891_), .A1(i_11_), .B0(men_men_n890_), .Y(men_men_n892_));
  AN2        u0870(.A(men_men_n97_), .B(men_men_n251_), .Y(men_men_n893_));
  NA2        u0871(.A(men_men_n769_), .B(men_men_n334_), .Y(men_men_n894_));
  AOI210     u0872(.A0(men_men_n498_), .A1(men_men_n87_), .B0(men_men_n58_), .Y(men_men_n895_));
  OAI220     u0873(.A0(men_men_n895_), .A1(men_men_n894_), .B0(men_men_n685_), .B1(men_men_n554_), .Y(men_men_n896_));
  NO2        u0874(.A(men_men_n259_), .B(men_men_n156_), .Y(men_men_n897_));
  NA2        u0875(.A(i_0_), .B(i_10_), .Y(men_men_n898_));
  INV        u0876(.A(men_men_n557_), .Y(men_men_n899_));
  NO4        u0877(.A(men_men_n116_), .B(men_men_n58_), .C(men_men_n692_), .D(i_5_), .Y(men_men_n900_));
  AO220      u0878(.A0(men_men_n900_), .A1(men_men_n899_), .B0(men_men_n897_), .B1(i_6_), .Y(men_men_n901_));
  AOI220     u0879(.A0(i_0_), .A1(men_men_n99_), .B0(men_men_n190_), .B1(men_men_n82_), .Y(men_men_n902_));
  NA2        u0880(.A(men_men_n588_), .B(i_4_), .Y(men_men_n903_));
  NA2        u0881(.A(men_men_n193_), .B(men_men_n208_), .Y(men_men_n904_));
  OAI220     u0882(.A0(men_men_n904_), .A1(men_men_n894_), .B0(men_men_n903_), .B1(men_men_n902_), .Y(men_men_n905_));
  NO4        u0883(.A(men_men_n905_), .B(men_men_n901_), .C(men_men_n896_), .D(men_men_n893_), .Y(men_men_n906_));
  NA4        u0884(.A(men_men_n906_), .B(men_men_n892_), .C(men_men_n888_), .D(men_men_n886_), .Y(men_men_n907_));
  NA2        u0885(.A(i_11_), .B(i_9_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n48_), .B(i_7_), .Y(men_men_n909_));
  NO2        u0887(.A(men_men_n908_), .B(men_men_n71_), .Y(men_men_n910_));
  NO2        u0888(.A(men_men_n179_), .B(i_0_), .Y(men_men_n911_));
  INV        u0889(.A(men_men_n911_), .Y(men_men_n912_));
  NA2        u0890(.A(men_men_n489_), .B(men_men_n238_), .Y(men_men_n913_));
  INV        u0891(.A(men_men_n412_), .Y(men_men_n914_));
  OAI220     u0892(.A0(men_men_n914_), .A1(men_men_n873_), .B0(men_men_n913_), .B1(men_men_n912_), .Y(men_men_n915_));
  INV        u0893(.A(men_men_n915_), .Y(men_men_n916_));
  NA2        u0894(.A(men_men_n684_), .B(men_men_n123_), .Y(men_men_n917_));
  NO2        u0895(.A(i_6_), .B(men_men_n917_), .Y(men_men_n918_));
  AOI210     u0896(.A0(men_men_n457_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n919_));
  NA2        u0897(.A(men_men_n175_), .B(men_men_n104_), .Y(men_men_n920_));
  NOi32      u0898(.An(men_men_n919_), .Bn(men_men_n193_), .C(men_men_n920_), .Y(men_men_n921_));
  AOI210     u0899(.A0(men_men_n630_), .A1(men_men_n334_), .B0(men_men_n251_), .Y(men_men_n922_));
  NO2        u0900(.A(men_men_n922_), .B(men_men_n865_), .Y(men_men_n923_));
  NO3        u0901(.A(men_men_n923_), .B(men_men_n921_), .C(men_men_n918_), .Y(men_men_n924_));
  NOi21      u0902(.An(i_7_), .B(i_5_), .Y(men_men_n925_));
  NOi31      u0903(.An(men_men_n925_), .B(i_0_), .C(men_men_n748_), .Y(men_men_n926_));
  NA3        u0904(.A(men_men_n926_), .B(men_men_n390_), .C(i_6_), .Y(men_men_n927_));
  OA210      u0905(.A0(men_men_n920_), .A1(men_men_n533_), .B0(men_men_n927_), .Y(men_men_n928_));
  NO3        u0906(.A(men_men_n408_), .B(men_men_n366_), .C(men_men_n362_), .Y(men_men_n929_));
  NO2        u0907(.A(men_men_n269_), .B(men_men_n324_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n748_), .B(men_men_n264_), .Y(men_men_n931_));
  AOI210     u0909(.A0(men_men_n931_), .A1(men_men_n930_), .B0(men_men_n929_), .Y(men_men_n932_));
  NA4        u0910(.A(men_men_n932_), .B(men_men_n928_), .C(men_men_n924_), .D(men_men_n916_), .Y(men_men_n933_));
  NO2        u0911(.A(men_men_n880_), .B(men_men_n247_), .Y(men_men_n934_));
  AN2        u0912(.A(men_men_n339_), .B(men_men_n334_), .Y(men_men_n935_));
  AN2        u0913(.A(men_men_n935_), .B(men_men_n876_), .Y(men_men_n936_));
  OAI210     u0914(.A0(men_men_n936_), .A1(men_men_n934_), .B0(i_10_), .Y(men_men_n937_));
  OA210      u0915(.A0(men_men_n489_), .A1(men_men_n230_), .B0(men_men_n488_), .Y(men_men_n938_));
  NA2        u0916(.A(i_10_), .B(men_men_n910_), .Y(men_men_n939_));
  NA3        u0917(.A(men_men_n488_), .B(men_men_n415_), .C(men_men_n45_), .Y(men_men_n940_));
  OAI210     u0918(.A0(men_men_n884_), .A1(i_7_), .B0(men_men_n940_), .Y(men_men_n941_));
  NO2        u0919(.A(men_men_n262_), .B(men_men_n46_), .Y(men_men_n942_));
  NO2        u0920(.A(men_men_n942_), .B(men_men_n192_), .Y(men_men_n943_));
  AOI220     u0921(.A0(men_men_n943_), .A1(men_men_n489_), .B0(men_men_n941_), .B1(men_men_n71_), .Y(men_men_n944_));
  NA3        u0922(.A(men_men_n832_), .B(men_men_n388_), .C(i_6_), .Y(men_men_n945_));
  NA2        u0923(.A(men_men_n93_), .B(men_men_n44_), .Y(men_men_n946_));
  NO2        u0924(.A(men_men_n73_), .B(men_men_n771_), .Y(men_men_n947_));
  AOI220     u0925(.A0(men_men_n947_), .A1(men_men_n946_), .B0(men_men_n178_), .B1(men_men_n619_), .Y(men_men_n948_));
  AOI210     u0926(.A0(men_men_n948_), .A1(men_men_n945_), .B0(men_men_n47_), .Y(men_men_n949_));
  NO3        u0927(.A(men_men_n610_), .B(men_men_n361_), .C(men_men_n24_), .Y(men_men_n950_));
  AOI210     u0928(.A0(men_men_n725_), .A1(men_men_n566_), .B0(men_men_n950_), .Y(men_men_n951_));
  NAi21      u0929(.An(i_9_), .B(i_5_), .Y(men_men_n952_));
  NO2        u0930(.A(men_men_n952_), .B(men_men_n408_), .Y(men_men_n953_));
  NO2        u0931(.A(men_men_n624_), .B(men_men_n106_), .Y(men_men_n954_));
  AOI220     u0932(.A0(men_men_n954_), .A1(i_0_), .B0(men_men_n953_), .B1(men_men_n647_), .Y(men_men_n955_));
  OAI220     u0933(.A0(men_men_n955_), .A1(men_men_n84_), .B0(men_men_n951_), .B1(men_men_n176_), .Y(men_men_n956_));
  NO3        u0934(.A(men_men_n956_), .B(men_men_n949_), .C(men_men_n537_), .Y(men_men_n957_));
  NA4        u0935(.A(men_men_n957_), .B(men_men_n944_), .C(men_men_n939_), .D(men_men_n937_), .Y(men_men_n958_));
  NO3        u0936(.A(men_men_n958_), .B(men_men_n933_), .C(men_men_n907_), .Y(men_men_n959_));
  NO2        u0937(.A(i_0_), .B(men_men_n748_), .Y(men_men_n960_));
  NA2        u0938(.A(men_men_n71_), .B(men_men_n44_), .Y(men_men_n961_));
  NA2        u0939(.A(men_men_n898_), .B(men_men_n961_), .Y(men_men_n962_));
  NO3        u0940(.A(men_men_n106_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n963_));
  AO220      u0941(.A0(men_men_n963_), .A1(men_men_n962_), .B0(men_men_n960_), .B1(men_men_n178_), .Y(men_men_n964_));
  AOI210     u0942(.A0(men_men_n814_), .A1(men_men_n712_), .B0(men_men_n920_), .Y(men_men_n965_));
  AOI210     u0943(.A0(men_men_n964_), .A1(men_men_n350_), .B0(men_men_n965_), .Y(men_men_n966_));
  NA2        u0944(.A(men_men_n759_), .B(men_men_n148_), .Y(men_men_n967_));
  INV        u0945(.A(men_men_n967_), .Y(men_men_n968_));
  NA3        u0946(.A(men_men_n968_), .B(men_men_n699_), .C(men_men_n71_), .Y(men_men_n969_));
  NO2        u0947(.A(men_men_n828_), .B(men_men_n408_), .Y(men_men_n970_));
  NA3        u0948(.A(men_men_n855_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n971_));
  NA2        u0949(.A(men_men_n856_), .B(i_9_), .Y(men_men_n972_));
  AOI210     u0950(.A0(men_men_n971_), .A1(men_men_n513_), .B0(men_men_n972_), .Y(men_men_n973_));
  NA2        u0951(.A(men_men_n252_), .B(men_men_n237_), .Y(men_men_n974_));
  AOI210     u0952(.A0(men_men_n974_), .A1(men_men_n889_), .B0(men_men_n156_), .Y(men_men_n975_));
  NO3        u0953(.A(men_men_n975_), .B(men_men_n973_), .C(men_men_n970_), .Y(men_men_n976_));
  NA3        u0954(.A(men_men_n976_), .B(men_men_n969_), .C(men_men_n966_), .Y(men_men_n977_));
  NA2        u0955(.A(men_men_n935_), .B(men_men_n378_), .Y(men_men_n978_));
  AOI210     u0956(.A0(men_men_n308_), .A1(men_men_n165_), .B0(men_men_n978_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n39_), .B(men_men_n44_), .Y(men_men_n980_));
  NA2        u0958(.A(men_men_n909_), .B(men_men_n501_), .Y(men_men_n981_));
  AOI210     u0959(.A0(men_men_n980_), .A1(men_men_n165_), .B0(men_men_n981_), .Y(men_men_n982_));
  NO2        u0960(.A(men_men_n982_), .B(men_men_n979_), .Y(men_men_n983_));
  NO3        u0961(.A(men_men_n898_), .B(men_men_n872_), .C(men_men_n195_), .Y(men_men_n984_));
  AOI220     u0962(.A0(men_men_n984_), .A1(i_11_), .B0(men_men_n589_), .B1(men_men_n73_), .Y(men_men_n985_));
  NO3        u0963(.A(men_men_n215_), .B(men_men_n389_), .C(i_0_), .Y(men_men_n986_));
  OAI210     u0964(.A0(men_men_n986_), .A1(men_men_n74_), .B0(i_13_), .Y(men_men_n987_));
  INV        u0965(.A(men_men_n224_), .Y(men_men_n988_));
  NO2        u0966(.A(men_men_n1082_), .B(men_men_n641_), .Y(men_men_n989_));
  NA3        u0967(.A(men_men_n989_), .B(men_men_n1080_), .C(men_men_n988_), .Y(men_men_n990_));
  NA4        u0968(.A(men_men_n990_), .B(men_men_n987_), .C(men_men_n985_), .D(men_men_n983_), .Y(men_men_n991_));
  NO2        u0969(.A(men_men_n250_), .B(men_men_n93_), .Y(men_men_n992_));
  AOI210     u0970(.A0(men_men_n992_), .A1(men_men_n960_), .B0(men_men_n110_), .Y(men_men_n993_));
  AOI220     u0971(.A0(men_men_n925_), .A1(men_men_n501_), .B0(men_men_n855_), .B1(men_men_n166_), .Y(men_men_n994_));
  NA2        u0972(.A(men_men_n353_), .B(men_men_n180_), .Y(men_men_n995_));
  OA220      u0973(.A0(men_men_n995_), .A1(men_men_n994_), .B0(men_men_n993_), .B1(i_5_), .Y(men_men_n996_));
  AOI210     u0974(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n179_), .Y(men_men_n997_));
  NA2        u0975(.A(men_men_n997_), .B(men_men_n938_), .Y(men_men_n998_));
  NA3        u0976(.A(men_men_n638_), .B(men_men_n190_), .C(men_men_n82_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n999_), .B(men_men_n564_), .Y(men_men_n1000_));
  NO3        u0978(.A(men_men_n865_), .B(men_men_n54_), .C(men_men_n48_), .Y(men_men_n1001_));
  NA3        u0979(.A(men_men_n506_), .B(men_men_n499_), .C(men_men_n486_), .Y(men_men_n1002_));
  NO3        u0980(.A(men_men_n1002_), .B(men_men_n1001_), .C(men_men_n1000_), .Y(men_men_n1003_));
  NA3        u0981(.A(men_men_n396_), .B(men_men_n175_), .C(men_men_n174_), .Y(men_men_n1004_));
  NA3        u0982(.A(men_men_n909_), .B(men_men_n297_), .C(men_men_n237_), .Y(men_men_n1005_));
  NA2        u0983(.A(men_men_n1005_), .B(men_men_n1004_), .Y(men_men_n1006_));
  NA3        u0984(.A(men_men_n396_), .B(men_men_n340_), .C(men_men_n228_), .Y(men_men_n1007_));
  INV        u0985(.A(men_men_n1007_), .Y(men_men_n1008_));
  NOi31      u0986(.An(men_men_n395_), .B(men_men_n961_), .C(men_men_n247_), .Y(men_men_n1009_));
  NO3        u0987(.A(men_men_n908_), .B(men_men_n224_), .C(men_men_n195_), .Y(men_men_n1010_));
  NO4        u0988(.A(men_men_n1010_), .B(men_men_n1009_), .C(men_men_n1008_), .D(men_men_n1006_), .Y(men_men_n1011_));
  NA4        u0989(.A(men_men_n1011_), .B(men_men_n1003_), .C(men_men_n998_), .D(men_men_n996_), .Y(men_men_n1012_));
  INV        u0990(.A(men_men_n640_), .Y(men_men_n1013_));
  NO3        u0991(.A(men_men_n1013_), .B(men_men_n579_), .C(i_3_), .Y(men_men_n1014_));
  INV        u0992(.A(men_men_n1014_), .Y(men_men_n1015_));
  NA3        u0993(.A(men_men_n312_), .B(i_5_), .C(men_men_n198_), .Y(men_men_n1016_));
  NAi31      u0994(.An(men_men_n249_), .B(men_men_n1016_), .C(men_men_n250_), .Y(men_men_n1017_));
  NO4        u0995(.A(men_men_n247_), .B(men_men_n215_), .C(i_0_), .D(i_12_), .Y(men_men_n1018_));
  AOI220     u0996(.A0(men_men_n1018_), .A1(men_men_n1017_), .B0(men_men_n808_), .B1(men_men_n180_), .Y(men_men_n1019_));
  AN2        u0997(.A(men_men_n898_), .B(men_men_n156_), .Y(men_men_n1020_));
  NO4        u0998(.A(men_men_n1020_), .B(i_12_), .C(men_men_n675_), .D(men_men_n133_), .Y(men_men_n1021_));
  NA2        u0999(.A(men_men_n1021_), .B(men_men_n224_), .Y(men_men_n1022_));
  NA3        u1000(.A(men_men_n99_), .B(men_men_n593_), .C(i_11_), .Y(men_men_n1023_));
  NA2        u1001(.A(men_men_n925_), .B(men_men_n485_), .Y(men_men_n1024_));
  NA2        u1002(.A(men_men_n64_), .B(men_men_n102_), .Y(men_men_n1025_));
  OAI220     u1003(.A0(men_men_n1025_), .A1(men_men_n1016_), .B0(men_men_n1024_), .B1(men_men_n700_), .Y(men_men_n1026_));
  NA2        u1004(.A(men_men_n1026_), .B(men_men_n911_), .Y(men_men_n1027_));
  NA4        u1005(.A(men_men_n1027_), .B(men_men_n1022_), .C(men_men_n1019_), .D(men_men_n1015_), .Y(men_men_n1028_));
  NO4        u1006(.A(men_men_n1028_), .B(men_men_n1012_), .C(men_men_n991_), .D(men_men_n977_), .Y(men_men_n1029_));
  OAI210     u1007(.A0(men_men_n831_), .A1(men_men_n826_), .B0(men_men_n37_), .Y(men_men_n1030_));
  NA3        u1008(.A(men_men_n919_), .B(men_men_n373_), .C(i_5_), .Y(men_men_n1031_));
  NA3        u1009(.A(men_men_n1031_), .B(men_men_n1030_), .C(men_men_n636_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n1032_), .B(men_men_n212_), .Y(men_men_n1033_));
  AN2        u1011(.A(men_men_n721_), .B(men_men_n374_), .Y(men_men_n1034_));
  NA2        u1012(.A(men_men_n191_), .B(men_men_n193_), .Y(men_men_n1035_));
  AO210      u1013(.A0(men_men_n1034_), .A1(men_men_n33_), .B0(men_men_n1035_), .Y(men_men_n1036_));
  NA2        u1014(.A(men_men_n638_), .B(men_men_n323_), .Y(men_men_n1037_));
  NAi31      u1015(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1038_));
  NA3        u1016(.A(men_men_n1038_), .B(men_men_n1037_), .C(men_men_n1036_), .Y(men_men_n1039_));
  NO2        u1017(.A(men_men_n475_), .B(men_men_n275_), .Y(men_men_n1040_));
  NO4        u1018(.A(men_men_n240_), .B(men_men_n147_), .C(men_men_n703_), .D(men_men_n37_), .Y(men_men_n1041_));
  NO3        u1019(.A(men_men_n1041_), .B(men_men_n1040_), .C(men_men_n891_), .Y(men_men_n1042_));
  NA2        u1020(.A(men_men_n1023_), .B(men_men_n1042_), .Y(men_men_n1043_));
  AOI210     u1021(.A0(men_men_n1039_), .A1(men_men_n48_), .B0(men_men_n1043_), .Y(men_men_n1044_));
  AOI210     u1022(.A0(men_men_n1044_), .A1(men_men_n1033_), .B0(men_men_n71_), .Y(men_men_n1045_));
  NO2        u1023(.A(men_men_n586_), .B(men_men_n385_), .Y(men_men_n1046_));
  NO2        u1024(.A(men_men_n1046_), .B(men_men_n776_), .Y(men_men_n1047_));
  OAI210     u1025(.A0(men_men_n78_), .A1(men_men_n54_), .B0(men_men_n109_), .Y(men_men_n1048_));
  NA2        u1026(.A(men_men_n1048_), .B(men_men_n74_), .Y(men_men_n1049_));
  AOI210     u1027(.A0(men_men_n997_), .A1(men_men_n909_), .B0(men_men_n926_), .Y(men_men_n1050_));
  AOI210     u1028(.A0(men_men_n1050_), .A1(men_men_n1049_), .B0(men_men_n703_), .Y(men_men_n1051_));
  NA2        u1029(.A(men_men_n269_), .B(men_men_n57_), .Y(men_men_n1052_));
  AOI220     u1030(.A0(men_men_n1052_), .A1(men_men_n74_), .B0(men_men_n348_), .B1(men_men_n261_), .Y(men_men_n1053_));
  NO2        u1031(.A(men_men_n1053_), .B(men_men_n244_), .Y(men_men_n1054_));
  NA3        u1032(.A(men_men_n97_), .B(men_men_n314_), .C(men_men_n31_), .Y(men_men_n1055_));
  INV        u1033(.A(men_men_n1055_), .Y(men_men_n1056_));
  NO3        u1034(.A(men_men_n1056_), .B(men_men_n1054_), .C(men_men_n1051_), .Y(men_men_n1057_));
  OAI210     u1035(.A0(men_men_n277_), .A1(men_men_n161_), .B0(men_men_n87_), .Y(men_men_n1058_));
  NA3        u1036(.A(men_men_n780_), .B(men_men_n297_), .C(men_men_n78_), .Y(men_men_n1059_));
  AOI210     u1037(.A0(men_men_n1059_), .A1(men_men_n1058_), .B0(i_11_), .Y(men_men_n1060_));
  NA2        u1038(.A(men_men_n631_), .B(men_men_n221_), .Y(men_men_n1061_));
  OAI210     u1039(.A0(men_men_n1061_), .A1(men_men_n919_), .B0(men_men_n212_), .Y(men_men_n1062_));
  NA2        u1040(.A(men_men_n167_), .B(i_5_), .Y(men_men_n1063_));
  AOI210     u1041(.A0(men_men_n1062_), .A1(men_men_n793_), .B0(men_men_n1063_), .Y(men_men_n1064_));
  NO3        u1042(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1065_));
  OAI210     u1043(.A0(men_men_n930_), .A1(men_men_n314_), .B0(men_men_n1065_), .Y(men_men_n1066_));
  NO2        u1044(.A(men_men_n1066_), .B(men_men_n748_), .Y(men_men_n1067_));
  NO4        u1045(.A(men_men_n952_), .B(i_11_), .C(i_3_), .D(men_men_n258_), .Y(men_men_n1068_));
  NO2        u1046(.A(men_men_n1068_), .B(men_men_n583_), .Y(men_men_n1069_));
  INV        u1047(.A(men_men_n367_), .Y(men_men_n1070_));
  AOI210     u1048(.A0(men_men_n1070_), .A1(men_men_n1069_), .B0(men_men_n40_), .Y(men_men_n1071_));
  NO4        u1049(.A(men_men_n1071_), .B(men_men_n1067_), .C(men_men_n1064_), .D(men_men_n1060_), .Y(men_men_n1072_));
  OAI210     u1050(.A0(men_men_n1057_), .A1(i_4_), .B0(men_men_n1072_), .Y(men_men_n1073_));
  NO3        u1051(.A(men_men_n1073_), .B(men_men_n1047_), .C(men_men_n1045_), .Y(men_men_n1074_));
  NA4        u1052(.A(men_men_n1074_), .B(men_men_n1029_), .C(men_men_n959_), .D(men_men_n879_), .Y(men4));
  INV        u1053(.A(i_2_), .Y(men_men_n1078_));
  INV        u1054(.A(i_5_), .Y(men_men_n1079_));
  INV        u1055(.A(i_3_), .Y(men_men_n1080_));
  INV        u1056(.A(i_6_), .Y(men_men_n1081_));
  INV        u1057(.A(i_6_), .Y(men_men_n1082_));
  INV        u1058(.A(i_9_), .Y(men_men_n1083_));
  INV        u1059(.A(i_5_), .Y(men_men_n1084_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule