typedef uvm_sequencer #(spi_beat) empty_sequencer;

// //  Class: empty_sequencer
// //
// class empty_sequencer extends uvm_sequencer #(empty_tx);
//   `uvm_component_utils(empty_sequencer);

//   //  Group: Configuration Object(s)


//   //  Group: Components


//   //  Group: Variables


//   //  Group: Functions

//   //  Constructor: new
//   function new(string name = "empty_sequencer", uvm_component parent);
//     super.new(name, parent);
//   endfunction: new


// endclass: empty_sequencer





