//Benchmark atmr_misex3_1774_0.125

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  INV        o0001(.A(d), .Y(ori_ori_n30_));
  BUFFER     o0002(.A(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  INV        o0010(.A(h), .Y(ori_ori_n39_));
  NAi21      o0011(.An(j), .B(l), .Y(ori_ori_n40_));
  NAi32      o0012(.An(n), .Bn(g), .C(m), .Y(ori_ori_n41_));
  NO3        o0013(.A(ori_ori_n41_), .B(ori_ori_n40_), .C(ori_ori_n39_), .Y(ori_ori_n42_));
  NAi31      o0014(.An(n), .B(m), .C(l), .Y(ori_ori_n43_));
  INV        o0015(.A(i), .Y(ori_ori_n44_));
  AN2        o0016(.A(h), .B(g), .Y(ori_ori_n45_));
  NA2        o0017(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori_ori_n46_));
  NO2        o0018(.A(ori_ori_n46_), .B(ori_ori_n43_), .Y(ori_ori_n47_));
  NAi21      o0019(.An(n), .B(m), .Y(ori_ori_n48_));
  NOi32      o0020(.An(k), .Bn(h), .C(l), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(g), .Y(ori_ori_n50_));
  INV        o0022(.A(ori_ori_n50_), .Y(ori_ori_n51_));
  NO2        o0023(.A(ori_ori_n51_), .B(ori_ori_n48_), .Y(ori_ori_n52_));
  NO3        o0024(.A(ori_ori_n52_), .B(ori_ori_n47_), .C(ori_ori_n42_), .Y(ori_ori_n53_));
  AOI210     o0025(.A0(ori_ori_n53_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n54_));
  INV        o0026(.A(c), .Y(ori_ori_n55_));
  NA2        o0027(.A(e), .B(b), .Y(ori_ori_n56_));
  INV        o0028(.A(d), .Y(ori_ori_n57_));
  NAi21      o0029(.An(i), .B(h), .Y(ori_ori_n58_));
  NAi41      o0030(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n59_));
  NA2        o0031(.A(g), .B(f), .Y(ori_ori_n60_));
  NO2        o0032(.A(ori_ori_n60_), .B(ori_ori_n59_), .Y(ori_ori_n61_));
  NAi31      o0033(.An(l), .B(m), .C(k), .Y(ori_ori_n62_));
  NAi41      o0034(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n63_));
  INV        o0035(.A(m), .Y(ori_ori_n64_));
  NOi21      o0036(.An(k), .B(l), .Y(ori_ori_n65_));
  NA2        o0037(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  AN4        o0038(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n67_));
  NOi31      o0039(.An(h), .B(g), .C(f), .Y(ori_ori_n68_));
  NA2        o0040(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  NAi32      o0041(.An(m), .Bn(k), .C(j), .Y(ori_ori_n70_));
  NOi32      o0042(.An(h), .Bn(g), .C(f), .Y(ori_ori_n71_));
  NA2        o0043(.A(ori_ori_n71_), .B(ori_ori_n67_), .Y(ori_ori_n72_));
  OA220      o0044(.A0(ori_ori_n72_), .A1(ori_ori_n70_), .B0(ori_ori_n69_), .B1(ori_ori_n66_), .Y(ori_ori_n73_));
  INV        o0045(.A(ori_ori_n73_), .Y(ori_ori_n74_));
  INV        o0046(.A(n), .Y(ori_ori_n75_));
  BUFFER     o0047(.A(b), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  INV        o0049(.A(j), .Y(ori_ori_n78_));
  AN3        o0050(.A(m), .B(k), .C(i), .Y(ori_ori_n79_));
  NA3        o0051(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .Y(ori_ori_n80_));
  NAi32      o0052(.An(g), .Bn(f), .C(h), .Y(ori_ori_n81_));
  NAi31      o0053(.An(j), .B(m), .C(l), .Y(ori_ori_n82_));
  NO2        o0054(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n83_));
  NA2        o0055(.A(m), .B(l), .Y(ori_ori_n84_));
  NAi31      o0056(.An(k), .B(j), .C(g), .Y(ori_ori_n85_));
  NO3        o0057(.A(ori_ori_n85_), .B(ori_ori_n84_), .C(f), .Y(ori_ori_n86_));
  NOi32      o0058(.An(m), .Bn(l), .C(i), .Y(ori_ori_n87_));
  NOi32      o0059(.An(m), .Bn(j), .C(k), .Y(ori_ori_n88_));
  AOI220     o0060(.A0(ori_ori_n88_), .A1(g), .B0(ori_ori_n87_), .B1(g), .Y(ori_ori_n89_));
  NO2        o0061(.A(ori_ori_n89_), .B(f), .Y(ori_ori_n90_));
  NAi41      o0062(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n91_));
  AN2        o0063(.A(e), .B(b), .Y(ori_ori_n92_));
  NOi21      o0064(.An(i), .B(h), .Y(ori_ori_n93_));
  INV        o0065(.A(a), .Y(ori_ori_n94_));
  NA2        o0066(.A(ori_ori_n92_), .B(ori_ori_n94_), .Y(ori_ori_n95_));
  INV        o0067(.A(l), .Y(ori_ori_n96_));
  NOi21      o0068(.An(m), .B(n), .Y(ori_ori_n97_));
  AN2        o0069(.A(k), .B(h), .Y(ori_ori_n98_));
  INV        o0070(.A(b), .Y(ori_ori_n99_));
  NA2        o0071(.A(l), .B(j), .Y(ori_ori_n100_));
  AN2        o0072(.A(k), .B(i), .Y(ori_ori_n101_));
  NA2        o0073(.A(ori_ori_n101_), .B(ori_ori_n100_), .Y(ori_ori_n102_));
  NA2        o0074(.A(g), .B(e), .Y(ori_ori_n103_));
  NOi32      o0075(.An(c), .Bn(a), .C(d), .Y(ori_ori_n104_));
  NA2        o0076(.A(ori_ori_n104_), .B(ori_ori_n97_), .Y(ori_ori_n105_));
  NO2        o0077(.A(ori_ori_n1119_), .B(ori_ori_n77_), .Y(ori_ori_n106_));
  NOi31      o0078(.An(k), .B(m), .C(j), .Y(ori_ori_n107_));
  NA3        o0079(.A(ori_ori_n107_), .B(ori_ori_n68_), .C(ori_ori_n67_), .Y(ori_ori_n108_));
  NOi31      o0080(.An(k), .B(m), .C(i), .Y(ori_ori_n109_));
  INV        o0081(.A(ori_ori_n108_), .Y(ori_ori_n110_));
  NAi21      o0082(.An(g), .B(h), .Y(ori_ori_n111_));
  NAi21      o0083(.An(m), .B(n), .Y(ori_ori_n112_));
  NAi31      o0084(.An(e), .B(f), .C(b), .Y(ori_ori_n113_));
  NAi31      o0085(.An(j), .B(k), .C(h), .Y(ori_ori_n114_));
  NO2        o0086(.A(k), .B(j), .Y(ori_ori_n115_));
  AN2        o0087(.A(k), .B(j), .Y(ori_ori_n116_));
  NAi21      o0088(.An(c), .B(b), .Y(ori_ori_n117_));
  NA2        o0089(.A(f), .B(d), .Y(ori_ori_n118_));
  NA2        o0090(.A(h), .B(c), .Y(ori_ori_n119_));
  NAi31      o0091(.An(f), .B(e), .C(b), .Y(ori_ori_n120_));
  NA2        o0092(.A(d), .B(b), .Y(ori_ori_n121_));
  NAi21      o0093(.An(e), .B(f), .Y(ori_ori_n122_));
  NO2        o0094(.A(ori_ori_n122_), .B(ori_ori_n121_), .Y(ori_ori_n123_));
  NA2        o0095(.A(b), .B(a), .Y(ori_ori_n124_));
  NAi21      o0096(.An(c), .B(d), .Y(ori_ori_n125_));
  NAi31      o0097(.An(l), .B(k), .C(h), .Y(ori_ori_n126_));
  NO2        o0098(.A(ori_ori_n112_), .B(ori_ori_n126_), .Y(ori_ori_n127_));
  NA2        o0099(.A(ori_ori_n127_), .B(ori_ori_n123_), .Y(ori_ori_n128_));
  NAi21      o0100(.An(ori_ori_n110_), .B(ori_ori_n128_), .Y(ori_ori_n129_));
  NAi31      o0101(.An(e), .B(f), .C(b), .Y(ori_ori_n130_));
  INV        o0102(.A(ori_ori_n130_), .Y(ori_ori_n131_));
  NOi21      o0103(.An(h), .B(i), .Y(ori_ori_n132_));
  NOi21      o0104(.An(k), .B(m), .Y(ori_ori_n133_));
  NA3        o0105(.A(ori_ori_n133_), .B(ori_ori_n132_), .C(n), .Y(ori_ori_n134_));
  NOi21      o0106(.An(ori_ori_n131_), .B(ori_ori_n134_), .Y(ori_ori_n135_));
  NOi21      o0107(.An(h), .B(g), .Y(ori_ori_n136_));
  NO2        o0108(.A(ori_ori_n118_), .B(ori_ori_n117_), .Y(ori_ori_n137_));
  NAi31      o0109(.An(l), .B(j), .C(h), .Y(ori_ori_n138_));
  NO2        o0110(.A(ori_ori_n138_), .B(ori_ori_n48_), .Y(ori_ori_n139_));
  NA2        o0111(.A(ori_ori_n139_), .B(ori_ori_n61_), .Y(ori_ori_n140_));
  NOi32      o0112(.An(n), .Bn(k), .C(m), .Y(ori_ori_n141_));
  INV        o0113(.A(ori_ori_n140_), .Y(ori_ori_n142_));
  NAi31      o0114(.An(d), .B(f), .C(c), .Y(ori_ori_n143_));
  NAi31      o0115(.An(e), .B(f), .C(c), .Y(ori_ori_n144_));
  NA2        o0116(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n145_));
  NA2        o0117(.A(j), .B(h), .Y(ori_ori_n146_));
  OR3        o0118(.A(n), .B(m), .C(k), .Y(ori_ori_n147_));
  NO2        o0119(.A(ori_ori_n147_), .B(ori_ori_n146_), .Y(ori_ori_n148_));
  NAi32      o0120(.An(m), .Bn(k), .C(n), .Y(ori_ori_n149_));
  NO2        o0121(.A(ori_ori_n149_), .B(ori_ori_n146_), .Y(ori_ori_n150_));
  AOI220     o0122(.A0(ori_ori_n150_), .A1(ori_ori_n131_), .B0(ori_ori_n148_), .B1(ori_ori_n145_), .Y(ori_ori_n151_));
  NO2        o0123(.A(n), .B(m), .Y(ori_ori_n152_));
  NA2        o0124(.A(ori_ori_n152_), .B(ori_ori_n49_), .Y(ori_ori_n153_));
  NAi21      o0125(.An(f), .B(e), .Y(ori_ori_n154_));
  NA2        o0126(.A(d), .B(c), .Y(ori_ori_n155_));
  NO2        o0127(.A(ori_ori_n155_), .B(ori_ori_n154_), .Y(ori_ori_n156_));
  NOi21      o0128(.An(ori_ori_n156_), .B(ori_ori_n153_), .Y(ori_ori_n157_));
  NAi21      o0129(.An(h), .B(f), .Y(ori_ori_n158_));
  NOi32      o0130(.An(f), .Bn(c), .C(d), .Y(ori_ori_n159_));
  NOi32      o0131(.An(f), .Bn(c), .C(e), .Y(ori_ori_n160_));
  NO2        o0132(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NO3        o0133(.A(n), .B(m), .C(j), .Y(ori_ori_n162_));
  NA2        o0134(.A(ori_ori_n162_), .B(ori_ori_n98_), .Y(ori_ori_n163_));
  AO210      o0135(.A0(ori_ori_n163_), .A1(ori_ori_n153_), .B0(ori_ori_n161_), .Y(ori_ori_n164_));
  NAi31      o0136(.An(ori_ori_n157_), .B(ori_ori_n164_), .C(ori_ori_n151_), .Y(ori_ori_n165_));
  OR4        o0137(.A(ori_ori_n165_), .B(ori_ori_n142_), .C(ori_ori_n135_), .D(ori_ori_n129_), .Y(ori_ori_n166_));
  NO4        o0138(.A(ori_ori_n166_), .B(ori_ori_n106_), .C(ori_ori_n74_), .D(ori_ori_n54_), .Y(ori_ori_n167_));
  NA3        o0139(.A(m), .B(ori_ori_n96_), .C(j), .Y(ori_ori_n168_));
  NAi31      o0140(.An(n), .B(h), .C(g), .Y(ori_ori_n169_));
  NO2        o0141(.A(ori_ori_n169_), .B(ori_ori_n168_), .Y(ori_ori_n170_));
  NOi32      o0142(.An(m), .Bn(k), .C(l), .Y(ori_ori_n171_));
  NA3        o0143(.A(ori_ori_n171_), .B(ori_ori_n78_), .C(g), .Y(ori_ori_n172_));
  NO2        o0144(.A(ori_ori_n172_), .B(n), .Y(ori_ori_n173_));
  NOi21      o0145(.An(k), .B(j), .Y(ori_ori_n174_));
  NA4        o0146(.A(ori_ori_n174_), .B(ori_ori_n97_), .C(i), .D(g), .Y(ori_ori_n175_));
  AN2        o0147(.A(i), .B(g), .Y(ori_ori_n176_));
  INV        o0148(.A(ori_ori_n175_), .Y(ori_ori_n177_));
  NO2        o0149(.A(ori_ori_n177_), .B(ori_ori_n170_), .Y(ori_ori_n178_));
  NAi41      o0150(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n179_));
  INV        o0151(.A(ori_ori_n179_), .Y(ori_ori_n180_));
  INV        o0152(.A(f), .Y(ori_ori_n181_));
  INV        o0153(.A(g), .Y(ori_ori_n182_));
  NOi31      o0154(.An(i), .B(j), .C(h), .Y(ori_ori_n183_));
  NOi21      o0155(.An(l), .B(m), .Y(ori_ori_n184_));
  NA2        o0156(.A(ori_ori_n184_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NO3        o0157(.A(ori_ori_n185_), .B(ori_ori_n182_), .C(ori_ori_n181_), .Y(ori_ori_n186_));
  NA2        o0158(.A(ori_ori_n186_), .B(ori_ori_n180_), .Y(ori_ori_n187_));
  OAI210     o0159(.A0(ori_ori_n178_), .A1(ori_ori_n32_), .B0(ori_ori_n187_), .Y(ori_ori_n188_));
  NOi21      o0160(.An(n), .B(m), .Y(ori_ori_n189_));
  NAi21      o0161(.An(j), .B(h), .Y(ori_ori_n190_));
  XN2        o0162(.A(i), .B(h), .Y(ori_ori_n191_));
  NOi31      o0163(.An(k), .B(n), .C(m), .Y(ori_ori_n192_));
  NAi31      o0164(.An(f), .B(e), .C(c), .Y(ori_ori_n193_));
  NAi32      o0165(.An(m), .Bn(i), .C(k), .Y(ori_ori_n194_));
  INV        o0166(.A(k), .Y(ori_ori_n195_));
  NAi21      o0167(.An(n), .B(a), .Y(ori_ori_n196_));
  NO2        o0168(.A(ori_ori_n196_), .B(ori_ori_n121_), .Y(ori_ori_n197_));
  NAi41      o0169(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n198_));
  NO2        o0170(.A(ori_ori_n198_), .B(e), .Y(ori_ori_n199_));
  NAi41      o0171(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n200_));
  NO2        o0172(.A(ori_ori_n200_), .B(ori_ori_n181_), .Y(ori_ori_n201_));
  NA2        o0173(.A(ori_ori_n133_), .B(ori_ori_n93_), .Y(ori_ori_n202_));
  NAi21      o0174(.An(ori_ori_n202_), .B(ori_ori_n201_), .Y(ori_ori_n203_));
  NO2        o0175(.A(n), .B(a), .Y(ori_ori_n204_));
  NAi21      o0176(.An(h), .B(i), .Y(ori_ori_n205_));
  NA2        o0177(.A(ori_ori_n152_), .B(k), .Y(ori_ori_n206_));
  NO2        o0178(.A(ori_ori_n206_), .B(ori_ori_n205_), .Y(ori_ori_n207_));
  NA2        o0179(.A(ori_ori_n207_), .B(ori_ori_n159_), .Y(ori_ori_n208_));
  NA2        o0180(.A(ori_ori_n208_), .B(ori_ori_n203_), .Y(ori_ori_n209_));
  NOi21      o0181(.An(g), .B(e), .Y(ori_ori_n210_));
  NO2        o0182(.A(ori_ori_n63_), .B(ori_ori_n64_), .Y(ori_ori_n211_));
  NA2        o0183(.A(ori_ori_n211_), .B(ori_ori_n210_), .Y(ori_ori_n212_));
  NOi32      o0184(.An(l), .Bn(j), .C(i), .Y(ori_ori_n213_));
  AOI210     o0185(.A0(ori_ori_n65_), .A1(ori_ori_n78_), .B0(ori_ori_n213_), .Y(ori_ori_n214_));
  NAi21      o0186(.An(f), .B(g), .Y(ori_ori_n215_));
  NO2        o0187(.A(ori_ori_n215_), .B(ori_ori_n59_), .Y(ori_ori_n216_));
  NO2        o0188(.A(ori_ori_n214_), .B(ori_ori_n212_), .Y(ori_ori_n217_));
  NO3        o0189(.A(ori_ori_n217_), .B(ori_ori_n209_), .C(ori_ori_n188_), .Y(ori_ori_n218_));
  NO3        o0190(.A(ori_ori_n170_), .B(ori_ori_n47_), .C(ori_ori_n42_), .Y(ori_ori_n219_));
  NO2        o0191(.A(ori_ori_n219_), .B(ori_ori_n95_), .Y(ori_ori_n220_));
  NA3        o0192(.A(ori_ori_n57_), .B(c), .C(b), .Y(ori_ori_n221_));
  NAi21      o0193(.An(h), .B(g), .Y(ori_ori_n222_));
  NO2        o0194(.A(ori_ori_n202_), .B(ori_ori_n215_), .Y(ori_ori_n223_));
  NAi31      o0195(.An(e), .B(d), .C(a), .Y(ori_ori_n224_));
  NA3        o0196(.A(ori_ori_n133_), .B(ori_ori_n71_), .C(ori_ori_n67_), .Y(ori_ori_n225_));
  NA3        o0197(.A(ori_ori_n133_), .B(ori_ori_n132_), .C(ori_ori_n75_), .Y(ori_ori_n226_));
  NA3        o0198(.A(e), .B(c), .C(b), .Y(ori_ori_n227_));
  NAi32      o0199(.An(k), .Bn(i), .C(j), .Y(ori_ori_n228_));
  NAi31      o0200(.An(h), .B(l), .C(i), .Y(ori_ori_n229_));
  NA3        o0201(.A(ori_ori_n229_), .B(ori_ori_n228_), .C(ori_ori_n138_), .Y(ori_ori_n230_));
  NA2        o0202(.A(ori_ori_n216_), .B(ori_ori_n1120_), .Y(ori_ori_n231_));
  NAi21      o0203(.An(l), .B(k), .Y(ori_ori_n232_));
  NA2        o0204(.A(ori_ori_n136_), .B(l), .Y(ori_ori_n233_));
  NA2        o0205(.A(ori_ori_n101_), .B(g), .Y(ori_ori_n234_));
  OR3        o0206(.A(ori_ori_n63_), .B(ori_ori_n64_), .C(e), .Y(ori_ori_n235_));
  AOI210     o0207(.A0(ori_ori_n234_), .A1(ori_ori_n233_), .B0(ori_ori_n235_), .Y(ori_ori_n236_));
  INV        o0208(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NAi32      o0209(.An(j), .Bn(h), .C(i), .Y(ori_ori_n238_));
  NAi21      o0210(.An(m), .B(l), .Y(ori_ori_n239_));
  NA2        o0211(.A(h), .B(g), .Y(ori_ori_n240_));
  NA2        o0212(.A(ori_ori_n141_), .B(ori_ori_n44_), .Y(ori_ori_n241_));
  NO2        o0213(.A(ori_ori_n241_), .B(ori_ori_n240_), .Y(ori_ori_n242_));
  NA2        o0214(.A(ori_ori_n242_), .B(ori_ori_n137_), .Y(ori_ori_n243_));
  NA4        o0215(.A(ori_ori_n243_), .B(ori_ori_n237_), .C(ori_ori_n231_), .D(ori_ori_n225_), .Y(ori_ori_n244_));
  NAi32      o0216(.An(n), .Bn(m), .C(l), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n245_), .B(ori_ori_n238_), .Y(ori_ori_n246_));
  NA2        o0218(.A(ori_ori_n246_), .B(ori_ori_n156_), .Y(ori_ori_n247_));
  NAi31      o0219(.An(k), .B(l), .C(j), .Y(ori_ori_n248_));
  OAI210     o0220(.A0(ori_ori_n232_), .A1(j), .B0(ori_ori_n248_), .Y(ori_ori_n249_));
  INV        o0221(.A(ori_ori_n247_), .Y(ori_ori_n250_));
  NO3        o0222(.A(ori_ori_n250_), .B(ori_ori_n244_), .C(ori_ori_n220_), .Y(ori_ori_n251_));
  NAi41      o0223(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n252_));
  NAi31      o0224(.An(i), .B(l), .C(h), .Y(ori_ori_n253_));
  NO4        o0225(.A(ori_ori_n253_), .B(e), .C(ori_ori_n63_), .D(ori_ori_n64_), .Y(ori_ori_n254_));
  NA2        o0226(.A(e), .B(c), .Y(ori_ori_n255_));
  NO3        o0227(.A(ori_ori_n255_), .B(n), .C(d), .Y(ori_ori_n256_));
  NOi21      o0228(.An(f), .B(h), .Y(ori_ori_n257_));
  NA2        o0229(.A(ori_ori_n257_), .B(ori_ori_n101_), .Y(ori_ori_n258_));
  NO2        o0230(.A(ori_ori_n258_), .B(ori_ori_n182_), .Y(ori_ori_n259_));
  NAi31      o0231(.An(d), .B(e), .C(b), .Y(ori_ori_n260_));
  NA2        o0232(.A(ori_ori_n204_), .B(ori_ori_n92_), .Y(ori_ori_n261_));
  NOi31      o0233(.An(l), .B(n), .C(m), .Y(ori_ori_n262_));
  NA2        o0234(.A(ori_ori_n262_), .B(ori_ori_n183_), .Y(ori_ori_n263_));
  NO2        o0235(.A(ori_ori_n263_), .B(ori_ori_n161_), .Y(ori_ori_n264_));
  NAi32      o0236(.An(m), .Bn(j), .C(k), .Y(ori_ori_n265_));
  NAi41      o0237(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n266_));
  NOi31      o0238(.An(j), .B(m), .C(k), .Y(ori_ori_n267_));
  NO2        o0239(.A(ori_ori_n107_), .B(ori_ori_n267_), .Y(ori_ori_n268_));
  AN3        o0240(.A(h), .B(g), .C(f), .Y(ori_ori_n269_));
  NOi32      o0241(.An(m), .Bn(j), .C(l), .Y(ori_ori_n270_));
  NO2        o0242(.A(ori_ori_n239_), .B(ori_ori_n238_), .Y(ori_ori_n271_));
  NO2        o0243(.A(ori_ori_n185_), .B(g), .Y(ori_ori_n272_));
  NO2        o0244(.A(ori_ori_n130_), .B(ori_ori_n75_), .Y(ori_ori_n273_));
  AOI220     o0245(.A0(ori_ori_n273_), .A1(ori_ori_n272_), .B0(ori_ori_n201_), .B1(ori_ori_n271_), .Y(ori_ori_n274_));
  INV        o0246(.A(ori_ori_n194_), .Y(ori_ori_n275_));
  NA3        o0247(.A(ori_ori_n275_), .B(ori_ori_n269_), .C(ori_ori_n180_), .Y(ori_ori_n276_));
  NA2        o0248(.A(ori_ori_n276_), .B(ori_ori_n274_), .Y(ori_ori_n277_));
  NA3        o0249(.A(h), .B(g), .C(f), .Y(ori_ori_n278_));
  NO2        o0250(.A(ori_ori_n278_), .B(ori_ori_n66_), .Y(ori_ori_n279_));
  NA2        o0251(.A(ori_ori_n266_), .B(ori_ori_n179_), .Y(ori_ori_n280_));
  NA2        o0252(.A(ori_ori_n136_), .B(e), .Y(ori_ori_n281_));
  NA2        o0253(.A(ori_ori_n280_), .B(ori_ori_n279_), .Y(ori_ori_n282_));
  NOi32      o0254(.An(j), .Bn(g), .C(i), .Y(ori_ori_n283_));
  NA2        o0255(.A(ori_ori_n283_), .B(ori_ori_n97_), .Y(ori_ori_n284_));
  AO210      o0256(.A0(ori_ori_n95_), .A1(ori_ori_n32_), .B0(ori_ori_n284_), .Y(ori_ori_n285_));
  NOi32      o0257(.An(e), .Bn(b), .C(a), .Y(ori_ori_n286_));
  INV        o0258(.A(m), .Y(ori_ori_n287_));
  NO3        o0259(.A(ori_ori_n252_), .B(e), .C(ori_ori_n182_), .Y(ori_ori_n288_));
  NA2        o0260(.A(ori_ori_n175_), .B(ori_ori_n35_), .Y(ori_ori_n289_));
  AOI220     o0261(.A0(ori_ori_n289_), .A1(ori_ori_n286_), .B0(ori_ori_n288_), .B1(ori_ori_n287_), .Y(ori_ori_n290_));
  NO2        o0262(.A(ori_ori_n260_), .B(n), .Y(ori_ori_n291_));
  NA2        o0263(.A(ori_ori_n176_), .B(k), .Y(ori_ori_n292_));
  NA2        o0264(.A(m), .B(ori_ori_n181_), .Y(ori_ori_n293_));
  NA4        o0265(.A(ori_ori_n171_), .B(ori_ori_n78_), .C(g), .D(ori_ori_n181_), .Y(ori_ori_n294_));
  NAi41      o0266(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n295_));
  NA2        o0267(.A(ori_ori_n50_), .B(ori_ori_n97_), .Y(ori_ori_n296_));
  NO2        o0268(.A(ori_ori_n296_), .B(ori_ori_n295_), .Y(ori_ori_n297_));
  NA2        o0269(.A(ori_ori_n171_), .B(ori_ori_n291_), .Y(ori_ori_n298_));
  NA4        o0270(.A(ori_ori_n298_), .B(ori_ori_n290_), .C(ori_ori_n285_), .D(ori_ori_n282_), .Y(ori_ori_n299_));
  NO4        o0271(.A(ori_ori_n299_), .B(ori_ori_n277_), .C(ori_ori_n264_), .D(ori_ori_n254_), .Y(ori_ori_n300_));
  NA4        o0272(.A(ori_ori_n300_), .B(ori_ori_n251_), .C(ori_ori_n218_), .D(ori_ori_n167_), .Y(ori10));
  NA3        o0273(.A(m), .B(k), .C(i), .Y(ori_ori_n302_));
  NOi21      o0274(.An(e), .B(f), .Y(ori_ori_n303_));
  NAi31      o0275(.An(b), .B(f), .C(c), .Y(ori_ori_n304_));
  INV        o0276(.A(ori_ori_n304_), .Y(ori_ori_n305_));
  NOi32      o0277(.An(k), .Bn(h), .C(j), .Y(ori_ori_n306_));
  AN2        o0278(.A(j), .B(h), .Y(ori_ori_n307_));
  NO3        o0279(.A(n), .B(m), .C(k), .Y(ori_ori_n308_));
  NA2        o0280(.A(ori_ori_n308_), .B(ori_ori_n307_), .Y(ori_ori_n309_));
  NO3        o0281(.A(ori_ori_n309_), .B(ori_ori_n125_), .C(ori_ori_n181_), .Y(ori_ori_n310_));
  OR2        o0282(.A(m), .B(k), .Y(ori_ori_n311_));
  NO2        o0283(.A(ori_ori_n146_), .B(ori_ori_n311_), .Y(ori_ori_n312_));
  NA4        o0284(.A(n), .B(f), .C(c), .D(ori_ori_n99_), .Y(ori_ori_n313_));
  NOi21      o0285(.An(ori_ori_n312_), .B(ori_ori_n313_), .Y(ori_ori_n314_));
  NOi32      o0286(.An(d), .Bn(a), .C(c), .Y(ori_ori_n315_));
  NA2        o0287(.A(ori_ori_n315_), .B(ori_ori_n154_), .Y(ori_ori_n316_));
  NAi21      o0288(.An(i), .B(g), .Y(ori_ori_n317_));
  NAi31      o0289(.An(k), .B(m), .C(j), .Y(ori_ori_n318_));
  NO3        o0290(.A(ori_ori_n318_), .B(ori_ori_n317_), .C(n), .Y(ori_ori_n319_));
  NOi21      o0291(.An(ori_ori_n319_), .B(ori_ori_n316_), .Y(ori_ori_n320_));
  NO3        o0292(.A(ori_ori_n320_), .B(ori_ori_n314_), .C(ori_ori_n310_), .Y(ori_ori_n321_));
  NO2        o0293(.A(ori_ori_n313_), .B(ori_ori_n239_), .Y(ori_ori_n322_));
  NOi32      o0294(.An(f), .Bn(d), .C(c), .Y(ori_ori_n323_));
  NA2        o0295(.A(ori_ori_n323_), .B(ori_ori_n246_), .Y(ori_ori_n324_));
  NA2        o0296(.A(ori_ori_n324_), .B(ori_ori_n321_), .Y(ori_ori_n325_));
  NO2        o0297(.A(ori_ori_n57_), .B(ori_ori_n99_), .Y(ori_ori_n326_));
  NA2        o0298(.A(ori_ori_n204_), .B(ori_ori_n326_), .Y(ori_ori_n327_));
  INV        o0299(.A(e), .Y(ori_ori_n328_));
  NA2        o0300(.A(ori_ori_n45_), .B(e), .Y(ori_ori_n329_));
  OAI220     o0301(.A0(ori_ori_n329_), .A1(ori_ori_n168_), .B0(ori_ori_n172_), .B1(ori_ori_n328_), .Y(ori_ori_n330_));
  NO2        o0302(.A(ori_ori_n80_), .B(ori_ori_n328_), .Y(ori_ori_n331_));
  NO2        o0303(.A(ori_ori_n331_), .B(ori_ori_n330_), .Y(ori_ori_n332_));
  NOi32      o0304(.An(h), .Bn(e), .C(g), .Y(ori_ori_n333_));
  NA3        o0305(.A(ori_ori_n333_), .B(l), .C(m), .Y(ori_ori_n334_));
  NOi21      o0306(.An(g), .B(h), .Y(ori_ori_n335_));
  AN3        o0307(.A(m), .B(l), .C(i), .Y(ori_ori_n336_));
  NA3        o0308(.A(ori_ori_n336_), .B(ori_ori_n335_), .C(e), .Y(ori_ori_n337_));
  AN3        o0309(.A(h), .B(g), .C(e), .Y(ori_ori_n338_));
  NA2        o0310(.A(ori_ori_n338_), .B(ori_ori_n87_), .Y(ori_ori_n339_));
  AN3        o0311(.A(ori_ori_n339_), .B(ori_ori_n337_), .C(ori_ori_n334_), .Y(ori_ori_n340_));
  AOI210     o0312(.A0(ori_ori_n340_), .A1(ori_ori_n332_), .B0(ori_ori_n327_), .Y(ori_ori_n341_));
  NA3        o0313(.A(ori_ori_n315_), .B(ori_ori_n154_), .C(ori_ori_n75_), .Y(ori_ori_n342_));
  NAi31      o0314(.An(b), .B(c), .C(a), .Y(ori_ori_n343_));
  NO2        o0315(.A(ori_ori_n343_), .B(n), .Y(ori_ori_n344_));
  NA2        o0316(.A(ori_ori_n50_), .B(m), .Y(ori_ori_n345_));
  NO2        o0317(.A(ori_ori_n345_), .B(ori_ori_n122_), .Y(ori_ori_n346_));
  NA2        o0318(.A(ori_ori_n346_), .B(ori_ori_n344_), .Y(ori_ori_n347_));
  INV        o0319(.A(ori_ori_n347_), .Y(ori_ori_n348_));
  NO3        o0320(.A(ori_ori_n348_), .B(ori_ori_n341_), .C(ori_ori_n325_), .Y(ori_ori_n349_));
  NA2        o0321(.A(i), .B(g), .Y(ori_ori_n350_));
  NOi21      o0322(.An(a), .B(n), .Y(ori_ori_n351_));
  NOi21      o0323(.An(d), .B(c), .Y(ori_ori_n352_));
  NA2        o0324(.A(ori_ori_n352_), .B(ori_ori_n351_), .Y(ori_ori_n353_));
  NA3        o0325(.A(i), .B(g), .C(f), .Y(ori_ori_n354_));
  OR2        o0326(.A(ori_ori_n354_), .B(ori_ori_n62_), .Y(ori_ori_n355_));
  NA3        o0327(.A(ori_ori_n336_), .B(ori_ori_n335_), .C(ori_ori_n154_), .Y(ori_ori_n356_));
  AOI210     o0328(.A0(ori_ori_n356_), .A1(ori_ori_n355_), .B0(ori_ori_n353_), .Y(ori_ori_n357_));
  INV        o0329(.A(ori_ori_n357_), .Y(ori_ori_n358_));
  OR2        o0330(.A(n), .B(m), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n359_), .B(ori_ori_n126_), .Y(ori_ori_n360_));
  NO2        o0332(.A(ori_ori_n155_), .B(ori_ori_n122_), .Y(ori_ori_n361_));
  OAI210     o0333(.A0(ori_ori_n360_), .A1(ori_ori_n148_), .B0(ori_ori_n361_), .Y(ori_ori_n362_));
  INV        o0334(.A(ori_ori_n296_), .Y(ori_ori_n363_));
  NO2        o0335(.A(ori_ori_n343_), .B(ori_ori_n48_), .Y(ori_ori_n364_));
  NO2        o0336(.A(ori_ori_n60_), .B(ori_ori_n96_), .Y(ori_ori_n365_));
  NAi21      o0337(.An(k), .B(j), .Y(ori_ori_n366_));
  NA2        o0338(.A(ori_ori_n205_), .B(ori_ori_n366_), .Y(ori_ori_n367_));
  NA3        o0339(.A(ori_ori_n367_), .B(ori_ori_n365_), .C(ori_ori_n364_), .Y(ori_ori_n368_));
  NAi21      o0340(.An(e), .B(d), .Y(ori_ori_n369_));
  INV        o0341(.A(ori_ori_n369_), .Y(ori_ori_n370_));
  NO2        o0342(.A(ori_ori_n206_), .B(ori_ori_n181_), .Y(ori_ori_n371_));
  NA2        o0343(.A(ori_ori_n368_), .B(ori_ori_n362_), .Y(ori_ori_n372_));
  NO2        o0344(.A(ori_ori_n263_), .B(ori_ori_n181_), .Y(ori_ori_n373_));
  NA2        o0345(.A(ori_ori_n373_), .B(ori_ori_n370_), .Y(ori_ori_n374_));
  NOi31      o0346(.An(n), .B(m), .C(k), .Y(ori_ori_n375_));
  AOI220     o0347(.A0(ori_ori_n375_), .A1(ori_ori_n307_), .B0(ori_ori_n189_), .B1(ori_ori_n49_), .Y(ori_ori_n376_));
  NAi31      o0348(.An(g), .B(f), .C(c), .Y(ori_ori_n377_));
  NA2        o0349(.A(ori_ori_n374_), .B(ori_ori_n247_), .Y(ori_ori_n378_));
  NOi41      o0350(.An(ori_ori_n358_), .B(ori_ori_n378_), .C(ori_ori_n372_), .D(ori_ori_n217_), .Y(ori_ori_n379_));
  NOi32      o0351(.An(c), .Bn(a), .C(b), .Y(ori_ori_n380_));
  NA2        o0352(.A(ori_ori_n380_), .B(ori_ori_n97_), .Y(ori_ori_n381_));
  AN2        o0353(.A(e), .B(d), .Y(ori_ori_n382_));
  NO2        o0354(.A(ori_ori_n111_), .B(ori_ori_n40_), .Y(ori_ori_n383_));
  NO2        o0355(.A(ori_ori_n60_), .B(e), .Y(ori_ori_n384_));
  NOi31      o0356(.An(j), .B(k), .C(i), .Y(ori_ori_n385_));
  NOi21      o0357(.An(ori_ori_n138_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  NA3        o0358(.A(ori_ori_n386_), .B(ori_ori_n214_), .C(ori_ori_n102_), .Y(ori_ori_n387_));
  NA2        o0359(.A(ori_ori_n387_), .B(ori_ori_n384_), .Y(ori_ori_n388_));
  NO2        o0360(.A(ori_ori_n388_), .B(ori_ori_n381_), .Y(ori_ori_n389_));
  NO2        o0361(.A(ori_ori_n177_), .B(ori_ori_n173_), .Y(ori_ori_n390_));
  NOi21      o0362(.An(a), .B(b), .Y(ori_ori_n391_));
  NA3        o0363(.A(e), .B(d), .C(c), .Y(ori_ori_n392_));
  NAi21      o0364(.An(ori_ori_n392_), .B(ori_ori_n391_), .Y(ori_ori_n393_));
  NO2        o0365(.A(ori_ori_n342_), .B(ori_ori_n172_), .Y(ori_ori_n394_));
  NOi21      o0366(.An(ori_ori_n393_), .B(ori_ori_n394_), .Y(ori_ori_n395_));
  AOI210     o0367(.A0(ori_ori_n219_), .A1(ori_ori_n390_), .B0(ori_ori_n395_), .Y(ori_ori_n396_));
  NA2        o0368(.A(ori_ori_n305_), .B(ori_ori_n127_), .Y(ori_ori_n397_));
  OR2        o0369(.A(k), .B(j), .Y(ori_ori_n398_));
  NA2        o0370(.A(l), .B(k), .Y(ori_ori_n399_));
  NA3        o0371(.A(ori_ori_n399_), .B(ori_ori_n398_), .C(ori_ori_n189_), .Y(ori_ori_n400_));
  AOI210     o0372(.A0(ori_ori_n194_), .A1(ori_ori_n265_), .B0(ori_ori_n75_), .Y(ori_ori_n401_));
  NOi21      o0373(.An(ori_ori_n400_), .B(ori_ori_n401_), .Y(ori_ori_n402_));
  OR3        o0374(.A(ori_ori_n402_), .B(ori_ori_n119_), .C(ori_ori_n113_), .Y(ori_ori_n403_));
  NA2        o0375(.A(ori_ori_n225_), .B(ori_ori_n108_), .Y(ori_ori_n404_));
  NO3        o0376(.A(ori_ori_n342_), .B(ori_ori_n82_), .C(ori_ori_n111_), .Y(ori_ori_n405_));
  NO3        o0377(.A(ori_ori_n405_), .B(ori_ori_n404_), .C(ori_ori_n254_), .Y(ori_ori_n406_));
  NA3        o0378(.A(ori_ori_n406_), .B(ori_ori_n403_), .C(ori_ori_n397_), .Y(ori_ori_n407_));
  NO3        o0379(.A(ori_ori_n407_), .B(ori_ori_n396_), .C(ori_ori_n389_), .Y(ori_ori_n408_));
  NO2        o0380(.A(ori_ori_n158_), .B(ori_ori_n55_), .Y(ori_ori_n409_));
  NAi31      o0381(.An(j), .B(l), .C(i), .Y(ori_ori_n410_));
  OAI210     o0382(.A0(ori_ori_n410_), .A1(ori_ori_n112_), .B0(ori_ori_n91_), .Y(ori_ori_n411_));
  NA2        o0383(.A(ori_ori_n411_), .B(ori_ori_n409_), .Y(ori_ori_n412_));
  INV        o0384(.A(ori_ori_n157_), .Y(ori_ori_n413_));
  NA2        o0385(.A(ori_ori_n413_), .B(ori_ori_n412_), .Y(ori_ori_n414_));
  OAI210     o0386(.A0(ori_ori_n109_), .A1(ori_ori_n107_), .B0(n), .Y(ori_ori_n415_));
  XO2        o0387(.A(i), .B(h), .Y(ori_ori_n416_));
  NAi31      o0388(.An(c), .B(f), .C(d), .Y(ori_ori_n417_));
  AOI210     o0389(.A0(ori_ori_n226_), .A1(ori_ori_n163_), .B0(ori_ori_n417_), .Y(ori_ori_n418_));
  BUFFER     o0390(.A(ori_ori_n73_), .Y(ori_ori_n419_));
  NA2        o0391(.A(ori_ori_n192_), .B(ori_ori_n93_), .Y(ori_ori_n420_));
  AOI210     o0392(.A0(ori_ori_n420_), .A1(ori_ori_n153_), .B0(ori_ori_n417_), .Y(ori_ori_n421_));
  AOI210     o0393(.A0(ori_ori_n284_), .A1(ori_ori_n35_), .B0(ori_ori_n393_), .Y(ori_ori_n422_));
  NO2        o0394(.A(ori_ori_n422_), .B(ori_ori_n421_), .Y(ori_ori_n423_));
  AO220      o0395(.A0(ori_ori_n1120_), .A1(ori_ori_n216_), .B0(ori_ori_n139_), .B1(ori_ori_n61_), .Y(ori_ori_n424_));
  INV        o0396(.A(ori_ori_n236_), .Y(ori_ori_n425_));
  NAi41      o0397(.An(ori_ori_n424_), .B(ori_ori_n425_), .C(ori_ori_n423_), .D(ori_ori_n419_), .Y(ori_ori_n426_));
  NO2        o0398(.A(ori_ori_n426_), .B(ori_ori_n414_), .Y(ori_ori_n427_));
  NA4        o0399(.A(ori_ori_n427_), .B(ori_ori_n408_), .C(ori_ori_n379_), .D(ori_ori_n349_), .Y(ori11));
  NO2        o0400(.A(ori_ori_n63_), .B(f), .Y(ori_ori_n429_));
  NA2        o0401(.A(j), .B(g), .Y(ori_ori_n430_));
  NAi31      o0402(.An(i), .B(m), .C(l), .Y(ori_ori_n431_));
  NA3        o0403(.A(m), .B(k), .C(j), .Y(ori_ori_n432_));
  OAI220     o0404(.A0(ori_ori_n432_), .A1(ori_ori_n111_), .B0(ori_ori_n431_), .B1(ori_ori_n430_), .Y(ori_ori_n433_));
  NA2        o0405(.A(ori_ori_n433_), .B(ori_ori_n429_), .Y(ori_ori_n434_));
  NOi32      o0406(.An(e), .Bn(b), .C(f), .Y(ori_ori_n435_));
  NA2        o0407(.A(ori_ori_n45_), .B(j), .Y(ori_ori_n436_));
  NO2        o0408(.A(ori_ori_n436_), .B(ori_ori_n241_), .Y(ori_ori_n437_));
  NAi31      o0409(.An(d), .B(e), .C(a), .Y(ori_ori_n438_));
  NO2        o0410(.A(ori_ori_n438_), .B(n), .Y(ori_ori_n439_));
  AOI220     o0411(.A0(ori_ori_n439_), .A1(ori_ori_n90_), .B0(ori_ori_n437_), .B1(ori_ori_n435_), .Y(ori_ori_n440_));
  NAi41      o0412(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n441_));
  AN2        o0413(.A(ori_ori_n441_), .B(ori_ori_n295_), .Y(ori_ori_n442_));
  AOI210     o0414(.A0(ori_ori_n442_), .A1(ori_ori_n316_), .B0(ori_ori_n222_), .Y(ori_ori_n443_));
  NA2        o0415(.A(j), .B(i), .Y(ori_ori_n444_));
  NAi31      o0416(.An(n), .B(m), .C(k), .Y(ori_ori_n445_));
  NO3        o0417(.A(ori_ori_n445_), .B(ori_ori_n444_), .C(ori_ori_n96_), .Y(ori_ori_n446_));
  NO4        o0418(.A(n), .B(d), .C(ori_ori_n99_), .D(a), .Y(ori_ori_n447_));
  OR2        o0419(.A(n), .B(c), .Y(ori_ori_n448_));
  NO2        o0420(.A(ori_ori_n448_), .B(ori_ori_n124_), .Y(ori_ori_n449_));
  NO2        o0421(.A(ori_ori_n449_), .B(ori_ori_n447_), .Y(ori_ori_n450_));
  NOi32      o0422(.An(g), .Bn(f), .C(i), .Y(ori_ori_n451_));
  AOI220     o0423(.A0(ori_ori_n451_), .A1(ori_ori_n88_), .B0(ori_ori_n433_), .B1(f), .Y(ori_ori_n452_));
  NO2        o0424(.A(ori_ori_n452_), .B(ori_ori_n450_), .Y(ori_ori_n453_));
  INV        o0425(.A(ori_ori_n453_), .Y(ori_ori_n454_));
  NA2        o0426(.A(ori_ori_n116_), .B(ori_ori_n34_), .Y(ori_ori_n455_));
  OAI220     o0427(.A0(ori_ori_n455_), .A1(m), .B0(ori_ori_n436_), .B1(ori_ori_n194_), .Y(ori_ori_n456_));
  NOi41      o0428(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n457_));
  NAi32      o0429(.An(e), .Bn(b), .C(c), .Y(ori_ori_n458_));
  OR2        o0430(.A(ori_ori_n458_), .B(ori_ori_n75_), .Y(ori_ori_n459_));
  AN2        o0431(.A(ori_ori_n266_), .B(ori_ori_n252_), .Y(ori_ori_n460_));
  NA2        o0432(.A(ori_ori_n460_), .B(ori_ori_n459_), .Y(ori_ori_n461_));
  OA210      o0433(.A0(ori_ori_n461_), .A1(ori_ori_n457_), .B0(ori_ori_n456_), .Y(ori_ori_n462_));
  OAI220     o0434(.A0(ori_ori_n318_), .A1(ori_ori_n317_), .B0(ori_ori_n431_), .B1(ori_ori_n430_), .Y(ori_ori_n463_));
  NAi31      o0435(.An(d), .B(c), .C(a), .Y(ori_ori_n464_));
  NO2        o0436(.A(ori_ori_n464_), .B(n), .Y(ori_ori_n465_));
  NO2        o0437(.A(ori_ori_n224_), .B(n), .Y(ori_ori_n466_));
  NO2        o0438(.A(ori_ori_n344_), .B(ori_ori_n466_), .Y(ori_ori_n467_));
  NA2        o0439(.A(ori_ori_n463_), .B(f), .Y(ori_ori_n468_));
  NAi32      o0440(.An(d), .Bn(a), .C(b), .Y(ori_ori_n469_));
  NA2        o0441(.A(h), .B(f), .Y(ori_ori_n470_));
  NO2        o0442(.A(ori_ori_n470_), .B(ori_ori_n85_), .Y(ori_ori_n471_));
  NO2        o0443(.A(ori_ori_n468_), .B(ori_ori_n467_), .Y(ori_ori_n472_));
  AN3        o0444(.A(j), .B(h), .C(g), .Y(ori_ori_n473_));
  NO2        o0445(.A(ori_ori_n121_), .B(c), .Y(ori_ori_n474_));
  NA3        o0446(.A(ori_ori_n474_), .B(ori_ori_n473_), .C(ori_ori_n375_), .Y(ori_ori_n475_));
  INV        o0447(.A(ori_ori_n475_), .Y(ori_ori_n476_));
  NO3        o0448(.A(ori_ori_n476_), .B(ori_ori_n472_), .C(ori_ori_n462_), .Y(ori_ori_n477_));
  AN4        o0449(.A(ori_ori_n477_), .B(ori_ori_n454_), .C(ori_ori_n440_), .D(ori_ori_n434_), .Y(ori_ori_n478_));
  INV        o0450(.A(k), .Y(ori_ori_n479_));
  NA3        o0451(.A(l), .B(ori_ori_n479_), .C(i), .Y(ori_ori_n480_));
  INV        o0452(.A(ori_ori_n480_), .Y(ori_ori_n481_));
  NA4        o0453(.A(ori_ori_n315_), .B(ori_ori_n335_), .C(ori_ori_n154_), .D(ori_ori_n97_), .Y(ori_ori_n482_));
  NAi32      o0454(.An(h), .Bn(f), .C(g), .Y(ori_ori_n483_));
  NAi41      o0455(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n484_));
  OAI210     o0456(.A0(ori_ori_n438_), .A1(n), .B0(ori_ori_n484_), .Y(ori_ori_n485_));
  NA2        o0457(.A(ori_ori_n485_), .B(m), .Y(ori_ori_n486_));
  NAi31      o0458(.An(h), .B(g), .C(f), .Y(ori_ori_n487_));
  OR2        o0459(.A(ori_ori_n486_), .B(ori_ori_n483_), .Y(ori_ori_n488_));
  NO3        o0460(.A(ori_ori_n483_), .B(ori_ori_n63_), .C(ori_ori_n64_), .Y(ori_ori_n489_));
  NO4        o0461(.A(ori_ori_n487_), .B(ori_ori_n448_), .C(ori_ori_n124_), .D(ori_ori_n64_), .Y(ori_ori_n490_));
  OR2        o0462(.A(ori_ori_n490_), .B(ori_ori_n489_), .Y(ori_ori_n491_));
  NAi31      o0463(.An(ori_ori_n491_), .B(ori_ori_n488_), .C(ori_ori_n482_), .Y(ori_ori_n492_));
  NAi31      o0464(.An(f), .B(h), .C(g), .Y(ori_ori_n493_));
  NOi32      o0465(.An(b), .Bn(a), .C(c), .Y(ori_ori_n494_));
  NOi32      o0466(.An(d), .Bn(a), .C(e), .Y(ori_ori_n495_));
  NA2        o0467(.A(ori_ori_n495_), .B(ori_ori_n97_), .Y(ori_ori_n496_));
  NO2        o0468(.A(n), .B(c), .Y(ori_ori_n497_));
  NA3        o0469(.A(ori_ori_n497_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n498_));
  NA2        o0470(.A(ori_ori_n498_), .B(ori_ori_n496_), .Y(ori_ori_n499_));
  NOi32      o0471(.An(e), .Bn(a), .C(d), .Y(ori_ori_n500_));
  AOI210     o0472(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n500_), .Y(ori_ori_n501_));
  INV        o0473(.A(ori_ori_n455_), .Y(ori_ori_n502_));
  NA2        o0474(.A(ori_ori_n502_), .B(ori_ori_n499_), .Y(ori_ori_n503_));
  OAI210     o0475(.A0(ori_ori_n203_), .A1(ori_ori_n78_), .B0(ori_ori_n503_), .Y(ori_ori_n504_));
  AOI210     o0476(.A0(ori_ori_n492_), .A1(ori_ori_n481_), .B0(ori_ori_n504_), .Y(ori_ori_n505_));
  NO3        o0477(.A(m), .B(ori_ori_n58_), .C(n), .Y(ori_ori_n506_));
  NA3        o0478(.A(ori_ori_n417_), .B(ori_ori_n144_), .C(ori_ori_n143_), .Y(ori_ori_n507_));
  NA2        o0479(.A(ori_ori_n377_), .B(ori_ori_n193_), .Y(ori_ori_n508_));
  BUFFER     o0480(.A(ori_ori_n507_), .Y(ori_ori_n509_));
  AOI220     o0481(.A0(ori_ori_n97_), .A1(ori_ori_n443_), .B0(ori_ori_n509_), .B1(ori_ori_n506_), .Y(ori_ori_n510_));
  NO2        o0482(.A(ori_ori_n510_), .B(ori_ori_n78_), .Y(ori_ori_n511_));
  NA3        o0483(.A(ori_ori_n457_), .B(ori_ori_n267_), .C(ori_ori_n45_), .Y(ori_ori_n512_));
  NOi32      o0484(.An(e), .Bn(c), .C(f), .Y(ori_ori_n513_));
  INV        o0485(.A(ori_ori_n179_), .Y(ori_ori_n514_));
  NA2        o0486(.A(ori_ori_n513_), .B(ori_ori_n148_), .Y(ori_ori_n515_));
  NA3        o0487(.A(ori_ori_n515_), .B(ori_ori_n512_), .C(ori_ori_n151_), .Y(ori_ori_n516_));
  AOI210     o0488(.A0(ori_ori_n442_), .A1(ori_ori_n316_), .B0(ori_ori_n240_), .Y(ori_ori_n517_));
  NAi21      o0489(.An(k), .B(h), .Y(ori_ori_n518_));
  NO2        o0490(.A(ori_ori_n518_), .B(ori_ori_n215_), .Y(ori_ori_n519_));
  NA2        o0491(.A(ori_ori_n519_), .B(j), .Y(ori_ori_n520_));
  OR2        o0492(.A(ori_ori_n520_), .B(ori_ori_n486_), .Y(ori_ori_n521_));
  NOi31      o0493(.An(m), .B(n), .C(k), .Y(ori_ori_n522_));
  NA2        o0494(.A(j), .B(ori_ori_n522_), .Y(ori_ori_n523_));
  AOI210     o0495(.A0(ori_ori_n316_), .A1(ori_ori_n295_), .B0(ori_ori_n240_), .Y(ori_ori_n524_));
  NAi21      o0496(.An(ori_ori_n523_), .B(ori_ori_n524_), .Y(ori_ori_n525_));
  NO2        o0497(.A(ori_ori_n224_), .B(ori_ori_n48_), .Y(ori_ori_n526_));
  NA2        o0498(.A(ori_ori_n526_), .B(ori_ori_n471_), .Y(ori_ori_n527_));
  NA3        o0499(.A(ori_ori_n527_), .B(ori_ori_n525_), .C(ori_ori_n521_), .Y(ori_ori_n528_));
  NA2        o0500(.A(ori_ori_n93_), .B(ori_ori_n36_), .Y(ori_ori_n529_));
  INV        o0501(.A(ori_ori_n286_), .Y(ori_ori_n530_));
  NO2        o0502(.A(ori_ori_n530_), .B(n), .Y(ori_ori_n531_));
  NAi31      o0503(.An(ori_ori_n529_), .B(ori_ori_n531_), .C(g), .Y(ori_ori_n532_));
  NO2        o0504(.A(ori_ori_n436_), .B(ori_ori_n149_), .Y(ori_ori_n533_));
  NA3        o0505(.A(ori_ori_n458_), .B(ori_ori_n221_), .C(ori_ori_n120_), .Y(ori_ori_n534_));
  NA2        o0506(.A(ori_ori_n416_), .B(ori_ori_n133_), .Y(ori_ori_n535_));
  NA2        o0507(.A(ori_ori_n534_), .B(ori_ori_n533_), .Y(ori_ori_n536_));
  AN3        o0508(.A(f), .B(d), .C(b), .Y(ori_ori_n537_));
  NAi31      o0509(.An(m), .B(n), .C(k), .Y(ori_ori_n538_));
  OR2        o0510(.A(ori_ori_n113_), .B(ori_ori_n58_), .Y(ori_ori_n539_));
  NO2        o0511(.A(ori_ori_n539_), .B(ori_ori_n538_), .Y(ori_ori_n540_));
  NA2        o0512(.A(ori_ori_n540_), .B(j), .Y(ori_ori_n541_));
  NA3        o0513(.A(ori_ori_n541_), .B(ori_ori_n536_), .C(ori_ori_n532_), .Y(ori_ori_n542_));
  NO4        o0514(.A(ori_ori_n542_), .B(ori_ori_n528_), .C(ori_ori_n516_), .D(ori_ori_n511_), .Y(ori_ori_n543_));
  NAi31      o0515(.An(g), .B(h), .C(f), .Y(ori_ori_n544_));
  OR3        o0516(.A(ori_ori_n544_), .B(ori_ori_n224_), .C(n), .Y(ori_ori_n545_));
  OA210      o0517(.A0(ori_ori_n438_), .A1(n), .B0(ori_ori_n484_), .Y(ori_ori_n546_));
  NA3        o0518(.A(ori_ori_n333_), .B(ori_ori_n104_), .C(ori_ori_n75_), .Y(ori_ori_n547_));
  OAI210     o0519(.A0(ori_ori_n546_), .A1(ori_ori_n81_), .B0(ori_ori_n547_), .Y(ori_ori_n548_));
  NOi21      o0520(.An(ori_ori_n545_), .B(ori_ori_n548_), .Y(ori_ori_n549_));
  NO2        o0521(.A(ori_ori_n549_), .B(ori_ori_n432_), .Y(ori_ori_n550_));
  NO3        o0522(.A(g), .B(ori_ori_n181_), .C(ori_ori_n55_), .Y(ori_ori_n551_));
  OR2        o0523(.A(ori_ori_n63_), .B(ori_ori_n64_), .Y(ori_ori_n552_));
  NA2        o0524(.A(ori_ori_n494_), .B(ori_ori_n269_), .Y(ori_ori_n553_));
  OA220      o0525(.A0(ori_ori_n523_), .A1(ori_ori_n553_), .B0(ori_ori_n520_), .B1(ori_ori_n552_), .Y(ori_ori_n554_));
  NA2        o0526(.A(h), .B(ori_ori_n37_), .Y(ori_ori_n555_));
  NA2        o0527(.A(ori_ori_n88_), .B(ori_ori_n45_), .Y(ori_ori_n556_));
  NO2        o0528(.A(ori_ori_n556_), .B(ori_ori_n261_), .Y(ori_ori_n557_));
  AOI210     o0529(.A0(ori_ori_n469_), .A1(ori_ori_n343_), .B0(ori_ori_n48_), .Y(ori_ori_n558_));
  OAI220     o0530(.A0(ori_ori_n487_), .A1(ori_ori_n480_), .B0(ori_ori_n258_), .B1(ori_ori_n430_), .Y(ori_ori_n559_));
  AOI210     o0531(.A0(ori_ori_n559_), .A1(ori_ori_n558_), .B0(ori_ori_n557_), .Y(ori_ori_n560_));
  NA2        o0532(.A(ori_ori_n560_), .B(ori_ori_n554_), .Y(ori_ori_n561_));
  INV        o0533(.A(ori_ori_n112_), .Y(ori_ori_n562_));
  AOI220     o0534(.A0(ori_ori_n562_), .A1(ori_ori_n435_), .B0(ori_ori_n286_), .B1(ori_ori_n97_), .Y(ori_ori_n563_));
  OR2        o0535(.A(ori_ori_n563_), .B(ori_ori_n455_), .Y(ori_ori_n564_));
  INV        o0536(.A(ori_ori_n564_), .Y(ori_ori_n565_));
  NO3        o0537(.A(ori_ori_n323_), .B(ori_ori_n160_), .C(ori_ori_n159_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n193_), .Y(ori_ori_n567_));
  NA3        o0539(.A(ori_ori_n567_), .B(ori_ori_n207_), .C(j), .Y(ori_ori_n568_));
  NO3        o0540(.A(ori_ori_n377_), .B(ori_ori_n146_), .C(i), .Y(ori_ori_n569_));
  NA2        o0541(.A(ori_ori_n380_), .B(ori_ori_n75_), .Y(ori_ori_n570_));
  NA2        o0542(.A(ori_ori_n568_), .B(ori_ori_n321_), .Y(ori_ori_n571_));
  NO4        o0543(.A(ori_ori_n571_), .B(ori_ori_n565_), .C(ori_ori_n561_), .D(ori_ori_n550_), .Y(ori_ori_n572_));
  NA4        o0544(.A(ori_ori_n572_), .B(ori_ori_n543_), .C(ori_ori_n505_), .D(ori_ori_n478_), .Y(ori08));
  NO2        o0545(.A(k), .B(h), .Y(ori_ori_n574_));
  AO210      o0546(.A0(ori_ori_n205_), .A1(ori_ori_n366_), .B0(ori_ori_n574_), .Y(ori_ori_n575_));
  NO2        o0547(.A(ori_ori_n575_), .B(ori_ori_n239_), .Y(ori_ori_n576_));
  NA2        o0548(.A(ori_ori_n513_), .B(ori_ori_n75_), .Y(ori_ori_n577_));
  INV        o0549(.A(ori_ori_n577_), .Y(ori_ori_n578_));
  AOI210     o0550(.A0(ori_ori_n578_), .A1(ori_ori_n576_), .B0(ori_ori_n405_), .Y(ori_ori_n579_));
  NA2        o0551(.A(ori_ori_n75_), .B(ori_ori_n94_), .Y(ori_ori_n580_));
  NO2        o0552(.A(ori_ori_n580_), .B(ori_ori_n56_), .Y(ori_ori_n581_));
  NO4        o0553(.A(ori_ori_n302_), .B(ori_ori_n96_), .C(j), .D(ori_ori_n182_), .Y(ori_ori_n582_));
  NA2        o0554(.A(ori_ori_n582_), .B(ori_ori_n581_), .Y(ori_ori_n583_));
  AN2        o0555(.A(l), .B(k), .Y(ori_ori_n584_));
  NA3        o0556(.A(ori_ori_n584_), .B(ori_ori_n93_), .C(ori_ori_n64_), .Y(ori_ori_n585_));
  NA3        o0557(.A(ori_ori_n583_), .B(ori_ori_n579_), .C(ori_ori_n274_), .Y(ori_ori_n586_));
  NO4        o0558(.A(ori_ori_n146_), .B(ori_ori_n311_), .C(ori_ori_n96_), .D(g), .Y(ori_ori_n587_));
  INV        o0559(.A(ori_ori_n38_), .Y(ori_ori_n588_));
  AOI220     o0560(.A0(ori_ori_n514_), .A1(ori_ori_n271_), .B0(ori_ori_n588_), .B1(ori_ori_n466_), .Y(ori_ori_n589_));
  INV        o0561(.A(ori_ori_n589_), .Y(ori_ori_n590_));
  NO2        o0562(.A(ori_ori_n442_), .B(ori_ori_n35_), .Y(ori_ori_n591_));
  OAI210     o0563(.A0(ori_ori_n458_), .A1(ori_ori_n46_), .B0(ori_ori_n539_), .Y(ori_ori_n592_));
  NO2        o0564(.A(ori_ori_n399_), .B(ori_ori_n112_), .Y(ori_ori_n593_));
  AOI210     o0565(.A0(ori_ori_n593_), .A1(ori_ori_n592_), .B0(ori_ori_n591_), .Y(ori_ori_n594_));
  INV        o0566(.A(ori_ori_n585_), .Y(ori_ori_n595_));
  NA2        o0567(.A(ori_ori_n575_), .B(ori_ori_n114_), .Y(ori_ori_n596_));
  AOI220     o0568(.A0(ori_ori_n596_), .A1(ori_ori_n322_), .B0(ori_ori_n595_), .B1(ori_ori_n67_), .Y(ori_ori_n597_));
  NA2        o0569(.A(ori_ori_n594_), .B(ori_ori_n597_), .Y(ori_ori_n598_));
  NA2        o0570(.A(ori_ori_n286_), .B(ori_ori_n42_), .Y(ori_ori_n599_));
  NA3        o0571(.A(m), .B(l), .C(k), .Y(ori_ori_n600_));
  AOI210     o0572(.A0(ori_ori_n547_), .A1(ori_ori_n545_), .B0(ori_ori_n600_), .Y(ori_ori_n601_));
  INV        o0573(.A(ori_ori_n601_), .Y(ori_ori_n602_));
  NA2        o0574(.A(ori_ori_n602_), .B(ori_ori_n599_), .Y(ori_ori_n603_));
  NO4        o0575(.A(ori_ori_n603_), .B(ori_ori_n598_), .C(ori_ori_n590_), .D(ori_ori_n586_), .Y(ori_ori_n604_));
  NO3        o0576(.A(ori_ori_n316_), .B(ori_ori_n430_), .C(h), .Y(ori_ori_n605_));
  NA2        o0577(.A(ori_ori_n605_), .B(ori_ori_n97_), .Y(ori_ori_n606_));
  NA2        o0578(.A(ori_ori_n606_), .B(ori_ori_n203_), .Y(ori_ori_n607_));
  NA2        o0579(.A(ori_ori_n584_), .B(ori_ori_n64_), .Y(ori_ori_n608_));
  NOi21      o0580(.An(h), .B(j), .Y(ori_ori_n609_));
  NA2        o0581(.A(ori_ori_n609_), .B(f), .Y(ori_ori_n610_));
  NO2        o0582(.A(ori_ori_n610_), .B(ori_ori_n200_), .Y(ori_ori_n611_));
  NO2        o0583(.A(ori_ori_n611_), .B(ori_ori_n569_), .Y(ori_ori_n612_));
  NO2        o0584(.A(ori_ori_n612_), .B(ori_ori_n608_), .Y(ori_ori_n613_));
  AOI210     o0585(.A0(ori_ori_n607_), .A1(l), .B0(ori_ori_n613_), .Y(ori_ori_n614_));
  NA2        o0586(.A(ori_ori_n71_), .B(l), .Y(ori_ori_n615_));
  OR2        o0587(.A(ori_ori_n615_), .B(ori_ori_n486_), .Y(ori_ori_n616_));
  NO3        o0588(.A(ori_ori_n125_), .B(ori_ori_n48_), .C(ori_ori_n94_), .Y(ori_ori_n617_));
  NO3        o0589(.A(ori_ori_n399_), .B(ori_ori_n354_), .C(j), .Y(ori_ori_n618_));
  INV        o0590(.A(j), .Y(ori_ori_n619_));
  NO3        o0591(.A(ori_ori_n239_), .B(ori_ori_n619_), .C(ori_ori_n39_), .Y(ori_ori_n620_));
  AOI210     o0592(.A0(ori_ori_n435_), .A1(n), .B0(ori_ori_n457_), .Y(ori_ori_n621_));
  NA2        o0593(.A(ori_ori_n621_), .B(ori_ori_n460_), .Y(ori_ori_n622_));
  AN3        o0594(.A(ori_ori_n622_), .B(ori_ori_n620_), .C(g), .Y(ori_ori_n623_));
  NO3        o0595(.A(ori_ori_n146_), .B(ori_ori_n311_), .C(ori_ori_n96_), .Y(ori_ori_n624_));
  AOI220     o0596(.A0(ori_ori_n624_), .A1(ori_ori_n201_), .B0(ori_ori_n508_), .B1(ori_ori_n246_), .Y(ori_ori_n625_));
  NAi31      o0597(.An(ori_ori_n501_), .B(ori_ori_n83_), .C(ori_ori_n75_), .Y(ori_ori_n626_));
  NA2        o0598(.A(ori_ori_n626_), .B(ori_ori_n625_), .Y(ori_ori_n627_));
  NO2        o0599(.A(ori_ori_n239_), .B(ori_ori_n114_), .Y(ori_ori_n628_));
  NA2        o0600(.A(ori_ori_n628_), .B(ori_ori_n514_), .Y(ori_ori_n629_));
  NO2        o0601(.A(ori_ori_n600_), .B(ori_ori_n81_), .Y(ori_ori_n630_));
  NO2        o0602(.A(ori_ori_n487_), .B(ori_ori_n100_), .Y(ori_ori_n631_));
  OAI210     o0603(.A0(ori_ori_n631_), .A1(ori_ori_n618_), .B0(ori_ori_n558_), .Y(ori_ori_n632_));
  NA2        o0604(.A(ori_ori_n632_), .B(ori_ori_n629_), .Y(ori_ori_n633_));
  OR3        o0605(.A(ori_ori_n633_), .B(ori_ori_n627_), .C(ori_ori_n623_), .Y(ori_ori_n634_));
  NA3        o0606(.A(ori_ori_n621_), .B(ori_ori_n460_), .C(ori_ori_n459_), .Y(ori_ori_n635_));
  NA4        o0607(.A(ori_ori_n635_), .B(ori_ori_n184_), .C(ori_ori_n366_), .D(ori_ori_n34_), .Y(ori_ori_n636_));
  NO3        o0608(.A(ori_ori_n399_), .B(ori_ori_n350_), .C(f), .Y(ori_ori_n637_));
  NO2        o0609(.A(ori_ori_n261_), .B(ori_ori_n38_), .Y(ori_ori_n638_));
  AOI210     o0610(.A0(ori_ori_n637_), .A1(ori_ori_n211_), .B0(ori_ori_n638_), .Y(ori_ori_n639_));
  NA3        o0611(.A(ori_ori_n451_), .B(l), .C(h), .Y(ori_ori_n640_));
  NO2        o0612(.A(ori_ori_n82_), .B(ori_ori_n46_), .Y(ori_ori_n641_));
  OAI220     o0613(.A0(ori_ori_n640_), .A1(ori_ori_n498_), .B0(ori_ori_n615_), .B1(ori_ori_n552_), .Y(ori_ori_n642_));
  AOI210     o0614(.A0(ori_ori_n641_), .A1(ori_ori_n531_), .B0(ori_ori_n642_), .Y(ori_ori_n643_));
  NA3        o0615(.A(ori_ori_n643_), .B(ori_ori_n639_), .C(ori_ori_n636_), .Y(ori_ori_n644_));
  BUFFER     o0616(.A(ori_ori_n630_), .Y(ori_ori_n645_));
  AOI220     o0617(.A0(ori_ori_n645_), .A1(ori_ori_n197_), .B0(ori_ori_n618_), .B1(ori_ori_n526_), .Y(ori_ori_n646_));
  NO2        o0618(.A(ori_ori_n546_), .B(ori_ori_n64_), .Y(ori_ori_n647_));
  AOI210     o0619(.A0(ori_ori_n637_), .A1(ori_ori_n647_), .B0(ori_ori_n264_), .Y(ori_ori_n648_));
  NO2        o0620(.A(ori_ori_n600_), .B(ori_ori_n544_), .Y(ori_ori_n649_));
  NA3        o0621(.A(ori_ori_n204_), .B(ori_ori_n57_), .C(b), .Y(ori_ori_n650_));
  AOI220     o0622(.A0(ori_ori_n497_), .A1(ori_ori_n29_), .B0(ori_ori_n380_), .B1(ori_ori_n75_), .Y(ori_ori_n651_));
  NA2        o0623(.A(ori_ori_n651_), .B(ori_ori_n650_), .Y(ori_ori_n652_));
  NA2        o0624(.A(ori_ori_n652_), .B(ori_ori_n649_), .Y(ori_ori_n653_));
  NA3        o0625(.A(ori_ori_n653_), .B(ori_ori_n648_), .C(ori_ori_n646_), .Y(ori_ori_n654_));
  NOi41      o0626(.An(ori_ori_n616_), .B(ori_ori_n654_), .C(ori_ori_n644_), .D(ori_ori_n634_), .Y(ori_ori_n655_));
  NO3        o0627(.A(ori_ori_n268_), .B(ori_ori_n240_), .C(ori_ori_n96_), .Y(ori_ori_n656_));
  NA2        o0628(.A(ori_ori_n656_), .B(ori_ori_n622_), .Y(ori_ori_n657_));
  NA2        o0629(.A(ori_ori_n657_), .B(ori_ori_n324_), .Y(ori_ori_n658_));
  NOi31      o0630(.An(b), .B(d), .C(a), .Y(ori_ori_n659_));
  NO2        o0631(.A(ori_ori_n659_), .B(ori_ori_n495_), .Y(ori_ori_n660_));
  NO2        o0632(.A(ori_ori_n660_), .B(n), .Y(ori_ori_n661_));
  NO2        o0633(.A(ori_ori_n640_), .B(ori_ori_n496_), .Y(ori_ori_n662_));
  NO2        o0634(.A(ori_ori_n458_), .B(ori_ori_n75_), .Y(ori_ori_n663_));
  NA2        o0635(.A(ori_ori_n656_), .B(ori_ori_n663_), .Y(ori_ori_n664_));
  INV        o0636(.A(ori_ori_n664_), .Y(ori_ori_n665_));
  NO2        o0637(.A(ori_ori_n566_), .B(n), .Y(ori_ori_n666_));
  BUFFER     o0638(.A(ori_ori_n628_), .Y(ori_ori_n667_));
  AOI220     o0639(.A0(ori_ori_n667_), .A1(ori_ori_n551_), .B0(ori_ori_n666_), .B1(ori_ori_n576_), .Y(ori_ori_n668_));
  NO2        o0640(.A(ori_ori_n255_), .B(ori_ori_n196_), .Y(ori_ori_n669_));
  NA2        o0641(.A(ori_ori_n83_), .B(ori_ori_n669_), .Y(ori_ori_n670_));
  INV        o0642(.A(ori_ori_n670_), .Y(ori_ori_n671_));
  NA2        o0643(.A(ori_ori_n587_), .B(ori_ori_n273_), .Y(ori_ori_n672_));
  OAI210     o0644(.A0(ori_ori_n490_), .A1(ori_ori_n489_), .B0(l), .Y(ori_ori_n673_));
  AN2        o0645(.A(ori_ori_n673_), .B(ori_ori_n672_), .Y(ori_ori_n674_));
  NAi31      o0646(.An(ori_ori_n671_), .B(ori_ori_n674_), .C(ori_ori_n668_), .Y(ori_ori_n675_));
  NO4        o0647(.A(ori_ori_n675_), .B(ori_ori_n665_), .C(ori_ori_n662_), .D(ori_ori_n658_), .Y(ori_ori_n676_));
  NA4        o0648(.A(ori_ori_n676_), .B(ori_ori_n655_), .C(ori_ori_n614_), .D(ori_ori_n604_), .Y(ori09));
  INV        o0649(.A(ori_ori_n105_), .Y(ori_ori_n678_));
  NA2        o0650(.A(f), .B(e), .Y(ori_ori_n679_));
  NO2        o0651(.A(ori_ori_n191_), .B(ori_ori_n96_), .Y(ori_ori_n680_));
  NA4        o0652(.A(ori_ori_n248_), .B(ori_ori_n386_), .C(ori_ori_n214_), .D(ori_ori_n102_), .Y(ori_ori_n681_));
  NA2        o0653(.A(ori_ori_n681_), .B(g), .Y(ori_ori_n682_));
  NO2        o0654(.A(ori_ori_n682_), .B(ori_ori_n679_), .Y(ori_ori_n683_));
  NA2        o0655(.A(ori_ori_n360_), .B(e), .Y(ori_ori_n684_));
  NO2        o0656(.A(ori_ori_n684_), .B(ori_ori_n417_), .Y(ori_ori_n685_));
  AOI210     o0657(.A0(ori_ori_n683_), .A1(ori_ori_n678_), .B0(ori_ori_n685_), .Y(ori_ori_n686_));
  NO2        o0658(.A(ori_ori_n172_), .B(ori_ori_n181_), .Y(ori_ori_n687_));
  NA3        o0659(.A(m), .B(l), .C(i), .Y(ori_ori_n688_));
  OAI220     o0660(.A0(ori_ori_n487_), .A1(ori_ori_n688_), .B0(ori_ori_n278_), .B1(ori_ori_n431_), .Y(ori_ori_n689_));
  NA4        o0661(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .D(f), .Y(ori_ori_n690_));
  NAi31      o0662(.An(ori_ori_n689_), .B(ori_ori_n690_), .C(ori_ori_n355_), .Y(ori_ori_n691_));
  OR2        o0663(.A(ori_ori_n691_), .B(ori_ori_n687_), .Y(ori_ori_n692_));
  INV        o0664(.A(ori_ori_n468_), .Y(ori_ori_n693_));
  OA210      o0665(.A0(ori_ori_n693_), .A1(ori_ori_n692_), .B0(ori_ori_n661_), .Y(ori_ori_n694_));
  INV        o0666(.A(ori_ori_n266_), .Y(ori_ori_n695_));
  NO2        o0667(.A(ori_ori_n109_), .B(ori_ori_n107_), .Y(ori_ori_n696_));
  NOi31      o0668(.An(k), .B(m), .C(l), .Y(ori_ori_n697_));
  NO2        o0669(.A(ori_ori_n267_), .B(ori_ori_n697_), .Y(ori_ori_n698_));
  AOI210     o0670(.A0(ori_ori_n698_), .A1(ori_ori_n696_), .B0(ori_ori_n493_), .Y(ori_ori_n699_));
  NA2        o0671(.A(ori_ori_n650_), .B(ori_ori_n261_), .Y(ori_ori_n700_));
  NA2        o0672(.A(ori_ori_n269_), .B(ori_ori_n270_), .Y(ori_ori_n701_));
  OAI210     o0673(.A0(ori_ori_n172_), .A1(ori_ori_n181_), .B0(ori_ori_n701_), .Y(ori_ori_n702_));
  AOI220     o0674(.A0(ori_ori_n702_), .A1(ori_ori_n700_), .B0(ori_ori_n699_), .B1(ori_ori_n695_), .Y(ori_ori_n703_));
  NA3        o0675(.A(ori_ori_n703_), .B(ori_ori_n515_), .C(ori_ori_n73_), .Y(ori_ori_n704_));
  NOi21      o0676(.An(f), .B(d), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n705_), .B(m), .Y(ori_ori_n706_));
  NO2        o0678(.A(ori_ori_n706_), .B(ori_ori_n51_), .Y(ori_ori_n707_));
  NOi32      o0679(.An(g), .Bn(f), .C(d), .Y(ori_ori_n708_));
  NA4        o0680(.A(ori_ori_n708_), .B(ori_ori_n497_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n709_));
  NOi21      o0681(.An(ori_ori_n249_), .B(ori_ori_n709_), .Y(ori_ori_n710_));
  AOI210     o0682(.A0(ori_ori_n707_), .A1(ori_ori_n449_), .B0(ori_ori_n710_), .Y(ori_ori_n711_));
  NA2        o0683(.A(ori_ori_n214_), .B(ori_ori_n102_), .Y(ori_ori_n712_));
  AN2        o0684(.A(f), .B(d), .Y(ori_ori_n713_));
  NA3        o0685(.A(ori_ori_n391_), .B(ori_ori_n713_), .C(ori_ori_n75_), .Y(ori_ori_n714_));
  NO3        o0686(.A(ori_ori_n714_), .B(ori_ori_n64_), .C(ori_ori_n182_), .Y(ori_ori_n715_));
  NA2        o0687(.A(ori_ori_n712_), .B(ori_ori_n715_), .Y(ori_ori_n716_));
  NAi31      o0688(.An(ori_ori_n404_), .B(ori_ori_n716_), .C(ori_ori_n711_), .Y(ori_ori_n717_));
  NO3        o0689(.A(ori_ori_n112_), .B(ori_ori_n260_), .C(ori_ori_n126_), .Y(ori_ori_n718_));
  INV        o0690(.A(ori_ori_n718_), .Y(ori_ori_n719_));
  NA2        o0691(.A(ori_ori_n495_), .B(ori_ori_n75_), .Y(ori_ori_n720_));
  NO2        o0692(.A(ori_ori_n701_), .B(ori_ori_n720_), .Y(ori_ori_n721_));
  INV        o0693(.A(ori_ori_n721_), .Y(ori_ori_n722_));
  NA2        o0694(.A(c), .B(ori_ori_n99_), .Y(ori_ori_n723_));
  OR2        o0695(.A(ori_ori_n544_), .B(ori_ori_n445_), .Y(ori_ori_n724_));
  INV        o0696(.A(ori_ori_n724_), .Y(ori_ori_n725_));
  INV        o0697(.A(ori_ori_n660_), .Y(ori_ori_n726_));
  NA2        o0698(.A(ori_ori_n726_), .B(ori_ori_n725_), .Y(ori_ori_n727_));
  NA3        o0699(.A(ori_ori_n727_), .B(ori_ori_n722_), .C(ori_ori_n719_), .Y(ori_ori_n728_));
  NO4        o0700(.A(ori_ori_n728_), .B(ori_ori_n717_), .C(ori_ori_n704_), .D(ori_ori_n694_), .Y(ori_ori_n729_));
  NO2        o0701(.A(ori_ori_n261_), .B(ori_ori_n690_), .Y(ori_ori_n730_));
  NO2        o0702(.A(ori_ori_n345_), .B(ori_ori_n679_), .Y(ori_ori_n731_));
  NA2        o0703(.A(ori_ori_n731_), .B(ori_ori_n465_), .Y(ori_ori_n732_));
  INV        o0704(.A(ori_ori_n732_), .Y(ori_ori_n733_));
  NA2        o0705(.A(e), .B(d), .Y(ori_ori_n734_));
  OAI220     o0706(.A0(ori_ori_n734_), .A1(c), .B0(ori_ori_n255_), .B1(d), .Y(ori_ori_n735_));
  NA3        o0707(.A(ori_ori_n735_), .B(ori_ori_n371_), .C(ori_ori_n416_), .Y(ori_ori_n736_));
  AOI210     o0708(.A0(ori_ori_n420_), .A1(ori_ori_n153_), .B0(ori_ori_n193_), .Y(ori_ori_n737_));
  AOI210     o0709(.A0(ori_ori_n514_), .A1(ori_ori_n271_), .B0(ori_ori_n737_), .Y(ori_ori_n738_));
  NA2        o0710(.A(ori_ori_n228_), .B(ori_ori_n138_), .Y(ori_ori_n739_));
  NA2        o0711(.A(ori_ori_n715_), .B(ori_ori_n739_), .Y(ori_ori_n740_));
  NA3        o0712(.A(ori_ori_n740_), .B(ori_ori_n738_), .C(ori_ori_n736_), .Y(ori_ori_n741_));
  NO3        o0713(.A(ori_ori_n741_), .B(ori_ori_n733_), .C(ori_ori_n730_), .Y(ori_ori_n742_));
  OR2        o0714(.A(ori_ori_n577_), .B(ori_ori_n185_), .Y(ori_ori_n743_));
  NO2        o0715(.A(ori_ori_n684_), .B(ori_ori_n143_), .Y(ori_ori_n744_));
  OAI210     o0716(.A0(ori_ori_n680_), .A1(ori_ori_n739_), .B0(ori_ori_n708_), .Y(ori_ori_n745_));
  NO2        o0717(.A(ori_ori_n745_), .B(ori_ori_n498_), .Y(ori_ori_n746_));
  AOI210     o0718(.A0(ori_ori_n101_), .A1(ori_ori_n100_), .B0(ori_ori_n213_), .Y(ori_ori_n747_));
  NO2        o0719(.A(ori_ori_n747_), .B(ori_ori_n709_), .Y(ori_ori_n748_));
  AO210      o0720(.A0(ori_ori_n700_), .A1(ori_ori_n689_), .B0(ori_ori_n748_), .Y(ori_ori_n749_));
  NOi31      o0721(.An(ori_ori_n449_), .B(ori_ori_n706_), .C(ori_ori_n233_), .Y(ori_ori_n750_));
  NO4        o0722(.A(ori_ori_n750_), .B(ori_ori_n749_), .C(ori_ori_n746_), .D(ori_ori_n744_), .Y(ori_ori_n751_));
  AN2        o0723(.A(ori_ori_n148_), .B(f), .Y(ori_ori_n752_));
  OAI210     o0724(.A0(ori_ori_n752_), .A1(ori_ori_n373_), .B0(ori_ori_n735_), .Y(ori_ori_n753_));
  NO2        o0725(.A(ori_ori_n354_), .B(ori_ori_n62_), .Y(ori_ori_n754_));
  OAI210     o0726(.A0(ori_ori_n693_), .A1(ori_ori_n754_), .B0(ori_ori_n581_), .Y(ori_ori_n755_));
  AN4        o0727(.A(ori_ori_n755_), .B(ori_ori_n753_), .C(ori_ori_n751_), .D(ori_ori_n743_), .Y(ori_ori_n756_));
  NA4        o0728(.A(ori_ori_n756_), .B(ori_ori_n742_), .C(ori_ori_n729_), .D(ori_ori_n686_), .Y(ori12));
  NO2        o0729(.A(ori_ori_n369_), .B(c), .Y(ori_ori_n758_));
  NO4        o0730(.A(ori_ori_n359_), .B(ori_ori_n205_), .C(ori_ori_n479_), .D(ori_ori_n182_), .Y(ori_ori_n759_));
  NA2        o0731(.A(ori_ori_n759_), .B(ori_ori_n758_), .Y(ori_ori_n760_));
  NA2        o0732(.A(ori_ori_n449_), .B(ori_ori_n754_), .Y(ori_ori_n761_));
  NO2        o0733(.A(ori_ori_n369_), .B(ori_ori_n99_), .Y(ori_ori_n762_));
  NO2        o0734(.A(ori_ori_n696_), .B(ori_ori_n278_), .Y(ori_ori_n763_));
  NO2        o0735(.A(ori_ori_n544_), .B(ori_ori_n302_), .Y(ori_ori_n764_));
  AOI220     o0736(.A0(ori_ori_n764_), .A1(ori_ori_n447_), .B0(ori_ori_n763_), .B1(ori_ori_n762_), .Y(ori_ori_n765_));
  NA4        o0737(.A(ori_ori_n765_), .B(ori_ori_n761_), .C(ori_ori_n760_), .D(ori_ori_n358_), .Y(ori_ori_n766_));
  AOI210     o0738(.A0(ori_ori_n194_), .A1(ori_ori_n265_), .B0(ori_ori_n169_), .Y(ori_ori_n767_));
  BUFFER     o0739(.A(ori_ori_n759_), .Y(ori_ori_n768_));
  AOI210     o0740(.A0(ori_ori_n263_), .A1(ori_ori_n309_), .B0(ori_ori_n182_), .Y(ori_ori_n769_));
  OAI210     o0741(.A0(ori_ori_n769_), .A1(ori_ori_n768_), .B0(ori_ori_n323_), .Y(ori_ori_n770_));
  NO2        o0742(.A(ori_ori_n529_), .B(ori_ori_n215_), .Y(ori_ori_n771_));
  NO2        o0743(.A(ori_ori_n487_), .B(ori_ori_n688_), .Y(ori_ori_n772_));
  NA2        o0744(.A(ori_ori_n669_), .B(ori_ori_n771_), .Y(ori_ori_n773_));
  NO2        o0745(.A(ori_ori_n125_), .B(ori_ori_n196_), .Y(ori_ori_n774_));
  NA2        o0746(.A(ori_ori_n774_), .B(ori_ori_n199_), .Y(ori_ori_n775_));
  NA3        o0747(.A(ori_ori_n775_), .B(ori_ori_n773_), .C(ori_ori_n770_), .Y(ori_ori_n776_));
  OR2        o0748(.A(ori_ori_n256_), .B(ori_ori_n762_), .Y(ori_ori_n777_));
  NA2        o0749(.A(ori_ori_n777_), .B(ori_ori_n279_), .Y(ori_ori_n778_));
  NO3        o0750(.A(ori_ori_n112_), .B(ori_ori_n126_), .C(ori_ori_n182_), .Y(ori_ori_n779_));
  NA2        o0751(.A(ori_ori_n779_), .B(ori_ori_n435_), .Y(ori_ori_n780_));
  NA4        o0752(.A(ori_ori_n360_), .B(ori_ori_n352_), .C(ori_ori_n154_), .D(g), .Y(ori_ori_n781_));
  NA3        o0753(.A(ori_ori_n781_), .B(ori_ori_n780_), .C(ori_ori_n778_), .Y(ori_ori_n782_));
  NO3        o0754(.A(ori_ori_n549_), .B(ori_ori_n82_), .C(ori_ori_n44_), .Y(ori_ori_n783_));
  NO4        o0755(.A(ori_ori_n783_), .B(ori_ori_n782_), .C(ori_ori_n776_), .D(ori_ori_n766_), .Y(ori_ori_n784_));
  NO2        o0756(.A(ori_ori_n293_), .B(ori_ori_n292_), .Y(ori_ori_n785_));
  NA2        o0757(.A(ori_ori_n484_), .B(ori_ori_n63_), .Y(ori_ori_n786_));
  INV        o0758(.A(ori_ori_n458_), .Y(ori_ori_n787_));
  NOi21      o0759(.An(ori_ori_n34_), .B(ori_ori_n538_), .Y(ori_ori_n788_));
  AOI220     o0760(.A0(ori_ori_n788_), .A1(ori_ori_n787_), .B0(ori_ori_n786_), .B1(ori_ori_n785_), .Y(ori_ori_n789_));
  INV        o0761(.A(ori_ori_n789_), .Y(ori_ori_n790_));
  NO2        o0762(.A(ori_ori_n48_), .B(ori_ori_n44_), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n415_), .B(ori_ori_n240_), .Y(ori_ori_n792_));
  INV        o0764(.A(ori_ori_n792_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n793_), .B(ori_ori_n120_), .Y(ori_ori_n794_));
  INV        o0766(.A(ori_ori_n290_), .Y(ori_ori_n795_));
  NO3        o0767(.A(ori_ori_n795_), .B(ori_ori_n794_), .C(ori_ori_n790_), .Y(ori_ori_n796_));
  NA2        o0768(.A(ori_ori_n271_), .B(g), .Y(ori_ori_n797_));
  NA2        o0769(.A(ori_ori_n136_), .B(i), .Y(ori_ori_n798_));
  NA2        o0770(.A(ori_ori_n45_), .B(i), .Y(ori_ori_n799_));
  OAI220     o0771(.A0(ori_ori_n799_), .A1(ori_ori_n168_), .B0(ori_ori_n798_), .B1(ori_ori_n82_), .Y(ori_ori_n800_));
  INV        o0772(.A(ori_ori_n800_), .Y(ori_ori_n801_));
  NO2        o0773(.A(ori_ori_n120_), .B(ori_ori_n75_), .Y(ori_ori_n802_));
  OR2        o0774(.A(ori_ori_n802_), .B(ori_ori_n457_), .Y(ori_ori_n803_));
  NA2        o0775(.A(ori_ori_n458_), .B(ori_ori_n304_), .Y(ori_ori_n804_));
  AOI210     o0776(.A0(ori_ori_n804_), .A1(n), .B0(ori_ori_n803_), .Y(ori_ori_n805_));
  OAI220     o0777(.A0(ori_ori_n805_), .A1(ori_ori_n797_), .B0(ori_ori_n801_), .B1(ori_ori_n261_), .Y(ori_ori_n806_));
  NA2        o0778(.A(ori_ori_n500_), .B(ori_ori_n97_), .Y(ori_ori_n807_));
  OR3        o0779(.A(ori_ori_n248_), .B(ori_ori_n350_), .C(f), .Y(ori_ori_n808_));
  NA3        o0780(.A(j), .B(ori_ori_n71_), .C(i), .Y(ori_ori_n809_));
  OA220      o0781(.A0(ori_ori_n809_), .A1(ori_ori_n807_), .B0(ori_ori_n808_), .B1(ori_ori_n486_), .Y(ori_ori_n810_));
  NA3        o0782(.A(ori_ori_n257_), .B(ori_ori_n101_), .C(g), .Y(ori_ori_n811_));
  AOI210     o0783(.A0(ori_ori_n555_), .A1(ori_ori_n811_), .B0(m), .Y(ori_ori_n812_));
  OAI210     o0784(.A0(ori_ori_n812_), .A1(ori_ori_n763_), .B0(ori_ori_n256_), .Y(ori_ori_n813_));
  NA2        o0785(.A(ori_ori_n570_), .B(ori_ori_n720_), .Y(ori_ori_n814_));
  NA2        o0786(.A(ori_ori_n690_), .B(ori_ori_n355_), .Y(ori_ori_n815_));
  NA2        o0787(.A(i), .B(ori_ori_n68_), .Y(ori_ori_n816_));
  NA2        o0788(.A(ori_ori_n816_), .B(ori_ori_n809_), .Y(ori_ori_n817_));
  AOI220     o0789(.A0(ori_ori_n817_), .A1(ori_ori_n211_), .B0(ori_ori_n815_), .B1(ori_ori_n814_), .Y(ori_ori_n818_));
  NA3        o0790(.A(ori_ori_n818_), .B(ori_ori_n813_), .C(ori_ori_n810_), .Y(ori_ori_n819_));
  NA2        o0791(.A(ori_ori_n771_), .B(ori_ori_n197_), .Y(ori_ori_n820_));
  NA2        o0792(.A(ori_ori_n548_), .B(ori_ori_n79_), .Y(ori_ori_n821_));
  NO2        o0793(.A(ori_ori_n376_), .B(ori_ori_n182_), .Y(ori_ori_n822_));
  AOI220     o0794(.A0(ori_ori_n822_), .A1(ori_ori_n305_), .B0(ori_ori_n777_), .B1(ori_ori_n186_), .Y(ori_ori_n823_));
  NA3        o0795(.A(ori_ori_n823_), .B(ori_ori_n821_), .C(ori_ori_n820_), .Y(ori_ori_n824_));
  OAI210     o0796(.A0(ori_ori_n815_), .A1(ori_ori_n772_), .B0(ori_ori_n447_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n293_), .B(ori_ori_n292_), .Y(ori_ori_n826_));
  NA2        o0798(.A(ori_ori_n826_), .B(ori_ori_n439_), .Y(ori_ori_n827_));
  NA2        o0799(.A(ori_ori_n812_), .B(ori_ori_n762_), .Y(ori_ori_n828_));
  NO3        o0800(.A(l), .B(ori_ori_n48_), .C(ori_ori_n44_), .Y(ori_ori_n829_));
  AOI220     o0801(.A0(ori_ori_n829_), .A1(ori_ori_n517_), .B0(ori_ori_n533_), .B1(ori_ori_n435_), .Y(ori_ori_n830_));
  NA4        o0802(.A(ori_ori_n830_), .B(ori_ori_n828_), .C(ori_ori_n827_), .D(ori_ori_n825_), .Y(ori_ori_n831_));
  NO4        o0803(.A(ori_ori_n831_), .B(ori_ori_n824_), .C(ori_ori_n819_), .D(ori_ori_n806_), .Y(ori_ori_n832_));
  NAi31      o0804(.An(ori_ori_n117_), .B(ori_ori_n338_), .C(n), .Y(ori_ori_n833_));
  NO3        o0805(.A(ori_ori_n107_), .B(ori_ori_n267_), .C(ori_ori_n697_), .Y(ori_ori_n834_));
  NO2        o0806(.A(ori_ori_n834_), .B(ori_ori_n833_), .Y(ori_ori_n835_));
  INV        o0807(.A(ori_ori_n835_), .Y(ori_ori_n836_));
  INV        o0808(.A(ori_ori_n405_), .Y(ori_ori_n837_));
  NA2        o0809(.A(ori_ori_n837_), .B(ori_ori_n836_), .Y(ori_ori_n838_));
  NA2        o0810(.A(ori_ori_n193_), .B(ori_ori_n144_), .Y(ori_ori_n839_));
  NO3        o0811(.A(ori_ori_n246_), .B(ori_ori_n360_), .C(ori_ori_n148_), .Y(ori_ori_n840_));
  NOi31      o0812(.An(ori_ori_n839_), .B(ori_ori_n840_), .C(ori_ori_n182_), .Y(ori_ori_n841_));
  NAi21      o0813(.An(ori_ori_n458_), .B(ori_ori_n822_), .Y(ori_ori_n842_));
  INV        o0814(.A(ori_ori_n842_), .Y(ori_ori_n843_));
  NO2        o0815(.A(ori_ori_n545_), .B(ori_ori_n302_), .Y(ori_ori_n844_));
  NA2        o0816(.A(ori_ori_n767_), .B(ori_ori_n758_), .Y(ori_ori_n845_));
  OAI220     o0817(.A0(ori_ori_n764_), .A1(ori_ori_n772_), .B0(ori_ori_n449_), .B1(ori_ori_n344_), .Y(ori_ori_n846_));
  NA3        o0818(.A(ori_ori_n846_), .B(ori_ori_n845_), .C(ori_ori_n512_), .Y(ori_ori_n847_));
  NA2        o0819(.A(ori_ori_n759_), .B(ori_ori_n839_), .Y(ori_ori_n848_));
  NA3        o0820(.A(ori_ori_n804_), .B(ori_ori_n401_), .C(ori_ori_n45_), .Y(ori_ori_n849_));
  NA2        o0821(.A(ori_ori_n849_), .B(ori_ori_n848_), .Y(ori_ori_n850_));
  OR3        o0822(.A(ori_ori_n850_), .B(ori_ori_n847_), .C(ori_ori_n844_), .Y(ori_ori_n851_));
  NO4        o0823(.A(ori_ori_n851_), .B(ori_ori_n843_), .C(ori_ori_n841_), .D(ori_ori_n838_), .Y(ori_ori_n852_));
  NA4        o0824(.A(ori_ori_n852_), .B(ori_ori_n832_), .C(ori_ori_n796_), .D(ori_ori_n784_), .Y(ori13));
  AN2        o0825(.A(d), .B(c), .Y(ori_ori_n854_));
  INV        o0826(.A(ori_ori_n854_), .Y(ori_ori_n855_));
  NAi32      o0827(.An(f), .Bn(e), .C(c), .Y(ori_ori_n856_));
  NO3        o0828(.A(m), .B(i), .C(h), .Y(ori_ori_n857_));
  NA3        o0829(.A(k), .B(j), .C(i), .Y(ori_ori_n858_));
  NO2        o0830(.A(f), .B(c), .Y(ori_ori_n859_));
  NOi21      o0831(.An(ori_ori_n859_), .B(ori_ori_n359_), .Y(ori_ori_n860_));
  AN3        o0832(.A(g), .B(f), .C(c), .Y(ori_ori_n861_));
  NA3        o0833(.A(l), .B(k), .C(j), .Y(ori_ori_n862_));
  NA2        o0834(.A(i), .B(h), .Y(ori_ori_n863_));
  NO3        o0835(.A(ori_ori_n863_), .B(ori_ori_n862_), .C(ori_ori_n112_), .Y(ori_ori_n864_));
  NO3        o0836(.A(ori_ori_n118_), .B(ori_ori_n227_), .C(ori_ori_n182_), .Y(ori_ori_n865_));
  NA3        o0837(.A(c), .B(b), .C(a), .Y(ori_ori_n866_));
  NO2        o0838(.A(ori_ori_n431_), .B(ori_ori_n493_), .Y(ori_ori_n867_));
  NA3        o0839(.A(ori_ori_n473_), .B(m), .C(ori_ori_n181_), .Y(ori_ori_n868_));
  NA2        o0840(.A(ori_ori_n868_), .B(ori_ori_n294_), .Y(ori_ori_n869_));
  NO3        o0841(.A(ori_ori_n869_), .B(ori_ori_n867_), .C(ori_ori_n826_), .Y(ori_ori_n870_));
  NO3        o0842(.A(ori_ori_n702_), .B(ori_ori_n691_), .C(ori_ori_n588_), .Y(ori_ori_n871_));
  OAI220     o0843(.A0(ori_ori_n871_), .A1(ori_ori_n570_), .B0(ori_ori_n870_), .B1(ori_ori_n484_), .Y(ori_ori_n872_));
  NOi31      o0844(.An(m), .B(n), .C(f), .Y(ori_ori_n873_));
  NA2        o0845(.A(ori_ori_n873_), .B(ori_ori_n50_), .Y(ori_ori_n874_));
  NO2        o0846(.A(ori_ori_n78_), .B(g), .Y(ori_ori_n875_));
  INV        o0847(.A(ori_ori_n872_), .Y(ori_ori_n876_));
  NA2        o0848(.A(c), .B(b), .Y(ori_ori_n877_));
  NO2        o0849(.A(ori_ori_n580_), .B(ori_ori_n877_), .Y(ori_ori_n878_));
  OAI210     o0850(.A0(ori_ori_n706_), .A1(ori_ori_n682_), .B0(ori_ori_n332_), .Y(ori_ori_n879_));
  OAI210     o0851(.A0(ori_ori_n879_), .A1(ori_ori_n707_), .B0(ori_ori_n878_), .Y(ori_ori_n880_));
  NAi21      o0852(.An(ori_ori_n340_), .B(ori_ori_n878_), .Y(ori_ori_n881_));
  NA2        o0853(.A(ori_ori_n344_), .B(ori_ori_n463_), .Y(ori_ori_n882_));
  NA2        o0854(.A(ori_ori_n882_), .B(ori_ori_n881_), .Y(ori_ori_n883_));
  OAI210     o0855(.A0(k), .A1(ori_ori_n230_), .B0(g), .Y(ori_ori_n884_));
  NAi21      o0856(.An(f), .B(d), .Y(ori_ori_n885_));
  NO2        o0857(.A(ori_ori_n885_), .B(ori_ori_n866_), .Y(ori_ori_n886_));
  INV        o0858(.A(ori_ori_n886_), .Y(ori_ori_n887_));
  NO2        o0859(.A(ori_ori_n884_), .B(ori_ori_n887_), .Y(ori_ori_n888_));
  AOI210     o0860(.A0(ori_ori_n888_), .A1(ori_ori_n97_), .B0(ori_ori_n883_), .Y(ori_ori_n889_));
  INV        o0861(.A(ori_ori_n383_), .Y(ori_ori_n890_));
  NO2        o0862(.A(ori_ori_n155_), .B(ori_ori_n196_), .Y(ori_ori_n891_));
  NA2        o0863(.A(ori_ori_n891_), .B(m), .Y(ori_ori_n892_));
  NA2        o0864(.A(ori_ori_n747_), .B(ori_ori_n386_), .Y(ori_ori_n893_));
  OAI210     o0865(.A0(ori_ori_n893_), .A1(ori_ori_n249_), .B0(ori_ori_n384_), .Y(ori_ori_n894_));
  AOI210     o0866(.A0(ori_ori_n894_), .A1(ori_ori_n890_), .B0(ori_ori_n892_), .Y(ori_ori_n895_));
  NA2        o0867(.A(ori_ori_n465_), .B(ori_ori_n330_), .Y(ori_ori_n896_));
  NA2        o0868(.A(ori_ori_n363_), .B(ori_ori_n886_), .Y(ori_ori_n897_));
  NO2        o0869(.A(ori_ori_n296_), .B(ori_ori_n295_), .Y(ori_ori_n898_));
  NA2        o0870(.A(ori_ori_n891_), .B(ori_ori_n346_), .Y(ori_ori_n899_));
  NAi41      o0871(.An(ori_ori_n898_), .B(ori_ori_n899_), .C(ori_ori_n897_), .D(ori_ori_n896_), .Y(ori_ori_n900_));
  NO2        o0872(.A(ori_ori_n900_), .B(ori_ori_n895_), .Y(ori_ori_n901_));
  NA4        o0873(.A(ori_ori_n901_), .B(ori_ori_n889_), .C(ori_ori_n880_), .D(ori_ori_n876_), .Y(ori00));
  INV        o0874(.A(ori_ori_n827_), .Y(ori_ori_n903_));
  OAI210     o0875(.A0(ori_ori_n834_), .A1(ori_ori_n39_), .B0(ori_ori_n535_), .Y(ori_ori_n904_));
  NA3        o0876(.A(ori_ori_n904_), .B(ori_ori_n210_), .C(n), .Y(ori_ori_n905_));
  NO2        o0877(.A(ori_ori_n905_), .B(ori_ori_n855_), .Y(ori_ori_n906_));
  NO2        o0878(.A(ori_ori_n906_), .B(ori_ori_n903_), .Y(ori_ori_n907_));
  NA3        o0879(.A(d), .B(ori_ori_n55_), .C(b), .Y(ori_ori_n908_));
  INV        o0880(.A(ori_ori_n475_), .Y(ori_ori_n909_));
  NO3        o0881(.A(ori_ori_n909_), .B(ori_ori_n898_), .C(ori_ori_n750_), .Y(ori_ori_n910_));
  NO3        o0882(.A(ori_ori_n402_), .B(ori_ori_n281_), .C(ori_ori_n877_), .Y(ori_ori_n911_));
  NA3        o0883(.A(ori_ori_n306_), .B(ori_ori_n189_), .C(g), .Y(ori_ori_n912_));
  OR2        o0884(.A(ori_ori_n912_), .B(ori_ori_n908_), .Y(ori_ori_n913_));
  NO2        o0885(.A(h), .B(g), .Y(ori_ori_n914_));
  NO2        o0886(.A(ori_ori_n82_), .B(ori_ori_n81_), .Y(ori_ori_n915_));
  AOI220     o0887(.A0(ori_ori_n915_), .A1(ori_ori_n439_), .B0(ori_ori_n779_), .B1(ori_ori_n474_), .Y(ori_ori_n916_));
  NA2        o0888(.A(ori_ori_n916_), .B(ori_ori_n913_), .Y(ori_ori_n917_));
  NO3        o0889(.A(ori_ori_n917_), .B(ori_ori_n911_), .C(ori_ori_n217_), .Y(ori_ori_n918_));
  INV        o0890(.A(ori_ori_n254_), .Y(ori_ori_n919_));
  NA2        o0891(.A(ori_ori_n201_), .B(ori_ori_n271_), .Y(ori_ori_n920_));
  NA3        o0892(.A(ori_ori_n920_), .B(ori_ori_n919_), .C(ori_ori_n128_), .Y(ori_ori_n921_));
  NO2        o0893(.A(ori_ori_n921_), .B(ori_ori_n424_), .Y(ori_ori_n922_));
  AN3        o0894(.A(ori_ori_n922_), .B(ori_ori_n918_), .C(ori_ori_n910_), .Y(ori_ori_n923_));
  NA2        o0895(.A(ori_ori_n439_), .B(ori_ori_n90_), .Y(ori_ori_n924_));
  INV        o0896(.A(ori_ori_n924_), .Y(ori_ori_n925_));
  NA2        o0897(.A(ori_ori_n869_), .B(ori_ori_n439_), .Y(ori_ori_n926_));
  NA4        o0898(.A(ori_ori_n537_), .B(ori_ori_n174_), .C(ori_ori_n189_), .D(ori_ori_n136_), .Y(ori_ori_n927_));
  NA3        o0899(.A(ori_ori_n927_), .B(ori_ori_n926_), .C(ori_ori_n237_), .Y(ori_ori_n928_));
  OAI210     o0900(.A0(ori_ori_n381_), .A1(ori_ori_n103_), .B0(ori_ori_n709_), .Y(ori_ori_n929_));
  AOI220     o0901(.A0(ori_ori_n929_), .A1(ori_ori_n893_), .B0(ori_ori_n465_), .B1(ori_ori_n330_), .Y(ori_ori_n930_));
  NA2        o0902(.A(n), .B(e), .Y(ori_ori_n931_));
  NO2        o0903(.A(ori_ori_n931_), .B(ori_ori_n121_), .Y(ori_ori_n932_));
  NA2        o0904(.A(ori_ori_n932_), .B(ori_ori_n223_), .Y(ori_ori_n933_));
  NA2        o0905(.A(ori_ori_n933_), .B(ori_ori_n930_), .Y(ori_ori_n934_));
  NA2        o0906(.A(ori_ori_n932_), .B(ori_ori_n699_), .Y(ori_ori_n935_));
  NA2        o0907(.A(ori_ori_n935_), .B(ori_ori_n711_), .Y(ori_ori_n936_));
  NO4        o0908(.A(ori_ori_n936_), .B(ori_ori_n934_), .C(ori_ori_n928_), .D(ori_ori_n925_), .Y(ori_ori_n937_));
  NA2        o0909(.A(ori_ori_n683_), .B(ori_ori_n617_), .Y(ori_ori_n938_));
  NA4        o0910(.A(ori_ori_n938_), .B(ori_ori_n937_), .C(ori_ori_n923_), .D(ori_ori_n907_), .Y(ori01));
  INV        o0911(.A(ori_ori_n394_), .Y(ori_ori_n940_));
  NA2        o0912(.A(ori_ori_n314_), .B(i), .Y(ori_ori_n941_));
  NA3        o0913(.A(ori_ori_n941_), .B(ori_ori_n940_), .C(ori_ori_n845_), .Y(ori_ori_n942_));
  NA2        o0914(.A(ori_ori_n458_), .B(ori_ori_n221_), .Y(ori_ori_n943_));
  NA2        o0915(.A(ori_ori_n792_), .B(ori_ori_n943_), .Y(ori_ori_n944_));
  INV        o0916(.A(ori_ori_n944_), .Y(ori_ori_n945_));
  NA2        o0917(.A(ori_ori_n44_), .B(f), .Y(ori_ori_n946_));
  NA2        o0918(.A(ori_ori_n584_), .B(g), .Y(ori_ori_n947_));
  NO2        o0919(.A(ori_ori_n947_), .B(ori_ori_n946_), .Y(ori_ori_n948_));
  OAI210     o0920(.A0(ori_ori_n640_), .A1(ori_ori_n496_), .B0(ori_ori_n927_), .Y(ori_ori_n949_));
  AOI210     o0921(.A0(ori_ori_n948_), .A1(ori_ori_n526_), .B0(ori_ori_n949_), .Y(ori_ori_n950_));
  INV        o0922(.A(ori_ori_n101_), .Y(ori_ori_n951_));
  OA220      o0923(.A0(ori_ori_n951_), .A1(ori_ori_n482_), .B0(ori_ori_n546_), .B1(ori_ori_n294_), .Y(ori_ori_n952_));
  NAi31      o0924(.An(ori_ori_n135_), .B(ori_ori_n952_), .C(ori_ori_n950_), .Y(ori_ori_n953_));
  NO2        o0925(.A(ori_ori_n557_), .B(ori_ori_n418_), .Y(ori_ori_n954_));
  NA3        o0926(.A(ori_ori_n584_), .B(g), .C(ori_ori_n181_), .Y(ori_ori_n955_));
  OA220      o0927(.A0(ori_ori_n955_), .A1(ori_ori_n552_), .B0(ori_ori_n163_), .B1(ori_ori_n161_), .Y(ori_ori_n956_));
  NA2        o0928(.A(ori_ori_n956_), .B(ori_ori_n954_), .Y(ori_ori_n957_));
  NO4        o0929(.A(ori_ori_n957_), .B(ori_ori_n953_), .C(ori_ori_n945_), .D(ori_ori_n942_), .Y(ori_ori_n958_));
  INV        o0930(.A(ori_ori_n912_), .Y(ori_ori_n959_));
  OAI210     o0931(.A0(ori_ori_n959_), .A1(ori_ori_n242_), .B0(ori_ori_n435_), .Y(ori_ori_n960_));
  AOI210     o0932(.A0(ori_ori_n172_), .A1(ori_ori_n80_), .B0(ori_ori_n181_), .Y(ori_ori_n961_));
  OAI210     o0933(.A0(ori_ori_n661_), .A1(ori_ori_n344_), .B0(ori_ori_n961_), .Y(ori_ori_n962_));
  NA2        o0934(.A(ori_ori_n962_), .B(ori_ori_n960_), .Y(ori_ori_n963_));
  NA2        o0935(.A(ori_ori_n491_), .B(ori_ori_n101_), .Y(ori_ori_n964_));
  OAI210     o0936(.A0(ori_ori_n951_), .A1(ori_ori_n488_), .B0(ori_ori_n964_), .Y(ori_ori_n965_));
  NA2        o0937(.A(ori_ori_n226_), .B(ori_ori_n163_), .Y(ori_ori_n966_));
  NA2        o0938(.A(ori_ori_n966_), .B(ori_ori_n551_), .Y(ori_ori_n967_));
  OAI210     o0939(.A0(ori_ori_n948_), .A1(ori_ori_n259_), .B0(ori_ori_n558_), .Y(ori_ori_n968_));
  NA3        o0940(.A(ori_ori_n968_), .B(ori_ori_n967_), .C(ori_ori_n643_), .Y(ori_ori_n969_));
  NO3        o0941(.A(ori_ori_n969_), .B(ori_ori_n965_), .C(ori_ori_n963_), .Y(ori_ori_n970_));
  NA3        o0942(.A(ori_ori_n497_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n971_));
  NO2        o0943(.A(ori_ori_n971_), .B(ori_ori_n172_), .Y(ori_ori_n972_));
  INV        o0944(.A(ori_ori_n972_), .Y(ori_ori_n973_));
  OR3        o0945(.A(ori_ori_n947_), .B(ori_ori_n498_), .C(ori_ori_n946_), .Y(ori_ori_n974_));
  NO2        o0946(.A(ori_ori_n955_), .B(ori_ori_n807_), .Y(ori_ori_n975_));
  NO2        o0947(.A(ori_ori_n175_), .B(ori_ori_n95_), .Y(ori_ori_n976_));
  NO2        o0948(.A(ori_ori_n976_), .B(ori_ori_n975_), .Y(ori_ori_n977_));
  NA4        o0949(.A(ori_ori_n977_), .B(ori_ori_n974_), .C(ori_ori_n973_), .D(ori_ori_n616_), .Y(ori_ori_n978_));
  NO3        o0950(.A(ori_ori_n70_), .B(ori_ori_n240_), .C(ori_ori_n44_), .Y(ori_ori_n979_));
  NA2        o0951(.A(ori_ori_n979_), .B(ori_ori_n457_), .Y(ori_ori_n980_));
  NA2        o0952(.A(ori_ori_n980_), .B(ori_ori_n554_), .Y(ori_ori_n981_));
  OR2        o0953(.A(ori_ori_n912_), .B(ori_ori_n908_), .Y(ori_ori_n982_));
  NO2        o0954(.A(ori_ori_n294_), .B(ori_ori_n63_), .Y(ori_ori_n983_));
  INV        o0955(.A(ori_ori_n983_), .Y(ori_ori_n984_));
  NA2        o0956(.A(ori_ori_n979_), .B(ori_ori_n663_), .Y(ori_ori_n985_));
  NA3        o0957(.A(ori_ori_n985_), .B(ori_ori_n984_), .C(ori_ori_n982_), .Y(ori_ori_n986_));
  NO3        o0958(.A(ori_ori_n986_), .B(ori_ori_n981_), .C(ori_ori_n978_), .Y(ori_ori_n987_));
  INV        o0959(.A(ori_ori_n113_), .Y(ori_ori_n988_));
  NO3        o0960(.A(ori_ori_n863_), .B(ori_ori_n149_), .C(ori_ori_n78_), .Y(ori_ori_n989_));
  AOI220     o0961(.A0(ori_ori_n989_), .A1(ori_ori_n988_), .B0(ori_ori_n979_), .B1(ori_ori_n802_), .Y(ori_ori_n990_));
  INV        o0962(.A(ori_ori_n990_), .Y(ori_ori_n991_));
  NO2        o0963(.A(ori_ori_n508_), .B(ori_ori_n507_), .Y(ori_ori_n992_));
  NO4        o0964(.A(ori_ori_n863_), .B(ori_ori_n992_), .C(ori_ori_n147_), .D(ori_ori_n78_), .Y(ori_ori_n993_));
  NO3        o0965(.A(ori_ori_n993_), .B(ori_ori_n991_), .C(ori_ori_n528_), .Y(ori_ori_n994_));
  NA4        o0966(.A(ori_ori_n994_), .B(ori_ori_n987_), .C(ori_ori_n970_), .D(ori_ori_n958_), .Y(ori06));
  NO2        o0967(.A(ori_ori_n190_), .B(ori_ori_n91_), .Y(ori_ori_n996_));
  OAI210     o0968(.A0(ori_ori_n996_), .A1(ori_ori_n989_), .B0(ori_ori_n305_), .Y(ori_ori_n997_));
  NO3        o0969(.A(ori_ori_n494_), .B(ori_ori_n659_), .C(ori_ori_n495_), .Y(ori_ori_n998_));
  OR2        o0970(.A(ori_ori_n998_), .B(ori_ori_n724_), .Y(ori_ori_n999_));
  NA2        o0971(.A(ori_ori_n999_), .B(ori_ori_n997_), .Y(ori_ori_n1000_));
  NO3        o0972(.A(ori_ori_n1000_), .B(ori_ori_n981_), .C(ori_ori_n209_), .Y(ori_ori_n1001_));
  NO2        o0973(.A(ori_ori_n240_), .B(ori_ori_n44_), .Y(ori_ori_n1002_));
  NA2        o0974(.A(ori_ori_n1002_), .B(ori_ori_n803_), .Y(ori_ori_n1003_));
  NA2        o0975(.A(ori_ori_n1002_), .B(ori_ori_n461_), .Y(ori_ori_n1004_));
  AOI210     o0976(.A0(ori_ori_n1004_), .A1(ori_ori_n1003_), .B0(ori_ori_n265_), .Y(ori_ori_n1005_));
  OAI210     o0977(.A0(ori_ori_n80_), .A1(ori_ori_n39_), .B0(ori_ori_n556_), .Y(ori_ori_n1006_));
  NA2        o0978(.A(ori_ori_n1006_), .B(ori_ori_n531_), .Y(ori_ori_n1007_));
  NO2        o0979(.A(ori_ori_n420_), .B(ori_ori_n144_), .Y(ori_ori_n1008_));
  NO2        o0980(.A(ori_ori_n501_), .B(ori_ori_n874_), .Y(ori_ori_n1009_));
  NO2        o0981(.A(ori_ori_n1009_), .B(ori_ori_n1008_), .Y(ori_ori_n1010_));
  NA2        o0982(.A(ori_ori_n1010_), .B(ori_ori_n1007_), .Y(ori_ori_n1011_));
  NO2        o0983(.A(ori_ori_n610_), .B(ori_ori_n292_), .Y(ori_ori_n1012_));
  NO2        o0984(.A(ori_ori_n558_), .B(ori_ori_n526_), .Y(ori_ori_n1013_));
  NOi21      o0985(.An(ori_ori_n1012_), .B(ori_ori_n1013_), .Y(ori_ori_n1014_));
  AN2        o0986(.A(ori_ori_n788_), .B(ori_ori_n534_), .Y(ori_ori_n1015_));
  NO4        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1014_), .C(ori_ori_n1011_), .D(ori_ori_n1005_), .Y(ori_ori_n1016_));
  NO3        o0988(.A(g), .B(ori_ori_n91_), .C(ori_ori_n227_), .Y(ori_ori_n1017_));
  OAI220     o0989(.A0(ori_ori_n577_), .A1(ori_ori_n202_), .B0(ori_ori_n417_), .B1(ori_ori_n420_), .Y(ori_ori_n1018_));
  NO2        o0990(.A(ori_ori_n493_), .B(j), .Y(ori_ori_n1019_));
  NOi21      o0991(.An(ori_ori_n1019_), .B(ori_ori_n552_), .Y(ori_ori_n1020_));
  NO3        o0992(.A(ori_ori_n1020_), .B(ori_ori_n1018_), .C(ori_ori_n1017_), .Y(ori_ori_n1021_));
  NA4        o0993(.A(ori_ori_n651_), .B(ori_ori_n650_), .C(ori_ori_n353_), .D(ori_ori_n720_), .Y(ori_ori_n1022_));
  NAi31      o0994(.An(ori_ori_n610_), .B(ori_ori_n1022_), .C(ori_ori_n171_), .Y(ori_ori_n1023_));
  NA2        o0995(.A(ori_ori_n1023_), .B(ori_ori_n1021_), .Y(ori_ori_n1024_));
  OR3        o0996(.A(ori_ori_n998_), .B(ori_ori_n640_), .C(ori_ori_n445_), .Y(ori_ori_n1025_));
  INV        o0997(.A(ori_ori_n297_), .Y(ori_ori_n1026_));
  NA2        o0998(.A(ori_ori_n1019_), .B(ori_ori_n647_), .Y(ori_ori_n1027_));
  NA3        o0999(.A(ori_ori_n1027_), .B(ori_ori_n1026_), .C(ori_ori_n1025_), .Y(ori_ori_n1028_));
  AN2        o1000(.A(ori_ori_n759_), .B(ori_ori_n758_), .Y(ori_ori_n1029_));
  INV        o1001(.A(ori_ori_n1029_), .Y(ori_ori_n1030_));
  NA2        o1002(.A(ori_ori_n1030_), .B(ori_ori_n985_), .Y(ori_ori_n1031_));
  NAi21      o1003(.An(j), .B(i), .Y(ori_ori_n1032_));
  NO4        o1004(.A(ori_ori_n992_), .B(ori_ori_n1032_), .C(ori_ori_n359_), .D(ori_ori_n195_), .Y(ori_ori_n1033_));
  NO4        o1005(.A(ori_ori_n1033_), .B(ori_ori_n1031_), .C(ori_ori_n1028_), .D(ori_ori_n1024_), .Y(ori_ori_n1034_));
  NA4        o1006(.A(ori_ori_n1034_), .B(ori_ori_n1016_), .C(ori_ori_n1001_), .D(ori_ori_n994_), .Y(ori07));
  NAi32      o1007(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1036_));
  NO3        o1008(.A(ori_ori_n1036_), .B(g), .C(f), .Y(ori_ori_n1037_));
  NOi31      o1009(.An(n), .B(m), .C(b), .Y(ori_ori_n1038_));
  NO3        o1010(.A(ori_ori_n112_), .B(ori_ori_n366_), .C(h), .Y(ori_ori_n1039_));
  NOi31      o1011(.An(i), .B(n), .C(h), .Y(ori_ori_n1040_));
  NO2        o1012(.A(ori_ori_n856_), .B(ori_ori_n359_), .Y(ori_ori_n1041_));
  NO2        o1013(.A(ori_ori_n858_), .B(ori_ori_n245_), .Y(ori_ori_n1042_));
  NO2        o1014(.A(ori_ori_n1041_), .B(ori_ori_n1037_), .Y(ori_ori_n1043_));
  NA3        o1015(.A(ori_ori_n574_), .B(ori_ori_n562_), .C(ori_ori_n96_), .Y(ori_ori_n1044_));
  NO2        o1016(.A(l), .B(k), .Y(ori_ori_n1045_));
  NO3        o1017(.A(ori_ori_n359_), .B(d), .C(c), .Y(ori_ori_n1046_));
  NO2        o1018(.A(g), .B(c), .Y(ori_ori_n1047_));
  NO2        o1019(.A(ori_ori_n369_), .B(a), .Y(ori_ori_n1048_));
  NA2        o1020(.A(ori_ori_n1048_), .B(ori_ori_n97_), .Y(ori_ori_n1049_));
  NOi31      o1021(.An(m), .B(n), .C(b), .Y(ori_ori_n1050_));
  NOi31      o1022(.An(f), .B(d), .C(c), .Y(ori_ori_n1051_));
  NA2        o1023(.A(ori_ori_n1051_), .B(ori_ori_n1050_), .Y(ori_ori_n1052_));
  NA2        o1024(.A(ori_ori_n861_), .B(ori_ori_n382_), .Y(ori_ori_n1053_));
  NO2        o1025(.A(ori_ori_n1053_), .B(ori_ori_n359_), .Y(ori_ori_n1054_));
  NO3        o1026(.A(ori_ori_n40_), .B(i), .C(h), .Y(ori_ori_n1055_));
  NO2        o1027(.A(ori_ori_n857_), .B(ori_ori_n1054_), .Y(ori_ori_n1056_));
  AN3        o1028(.A(ori_ori_n1056_), .B(ori_ori_n1052_), .C(ori_ori_n1049_), .Y(ori_ori_n1057_));
  NA2        o1029(.A(ori_ori_n1038_), .B(ori_ori_n303_), .Y(ori_ori_n1058_));
  INV        o1030(.A(ori_ori_n1058_), .Y(ori_ori_n1059_));
  INV        o1031(.A(ori_ori_n864_), .Y(ori_ori_n1060_));
  NAi21      o1032(.An(ori_ori_n1059_), .B(ori_ori_n1060_), .Y(ori_ori_n1061_));
  NO4        o1033(.A(ori_ori_n112_), .B(g), .C(f), .D(e), .Y(ori_ori_n1062_));
  NA2        o1034(.A(ori_ori_n1040_), .B(ori_ori_n1045_), .Y(ori_ori_n1063_));
  INV        o1035(.A(ori_ori_n1063_), .Y(ori_ori_n1064_));
  NA2        o1036(.A(ori_ori_n873_), .B(ori_ori_n328_), .Y(ori_ori_n1065_));
  NO2        o1037(.A(ori_ori_n1064_), .B(ori_ori_n1061_), .Y(ori_ori_n1066_));
  NA4        o1038(.A(ori_ori_n1066_), .B(ori_ori_n1057_), .C(ori_ori_n1044_), .D(ori_ori_n1043_), .Y(ori_ori_n1067_));
  NO2        o1039(.A(ori_ori_n877_), .B(ori_ori_n94_), .Y(ori_ori_n1068_));
  NO2        o1040(.A(ori_ori_n311_), .B(j), .Y(ori_ori_n1069_));
  NA2        o1041(.A(ori_ori_n1055_), .B(ori_ori_n873_), .Y(ori_ori_n1070_));
  NA2        o1042(.A(ori_ori_n860_), .B(e), .Y(ori_ori_n1071_));
  NA2        o1043(.A(ori_ori_n1071_), .B(ori_ori_n1070_), .Y(ori_ori_n1072_));
  NA2        o1044(.A(ori_ori_n1069_), .B(ori_ori_n132_), .Y(ori_ori_n1073_));
  INV        o1045(.A(ori_ori_n1073_), .Y(ori_ori_n1074_));
  NO2        o1046(.A(ori_ori_n1074_), .B(ori_ori_n1072_), .Y(ori_ori_n1075_));
  INV        o1047(.A(ori_ori_n48_), .Y(ori_ori_n1076_));
  NA2        o1048(.A(ori_ori_n1076_), .B(ori_ori_n914_), .Y(ori_ori_n1077_));
  INV        o1049(.A(ori_ori_n1077_), .Y(ori_ori_n1078_));
  NO2        o1050(.A(ori_ori_n190_), .B(ori_ori_n149_), .Y(ori_ori_n1079_));
  NO2        o1051(.A(ori_ori_n1079_), .B(ori_ori_n1078_), .Y(ori_ori_n1080_));
  NA2        o1052(.A(ori_ori_n1068_), .B(f), .Y(ori_ori_n1081_));
  NO2        o1053(.A(ori_ori_n1117_), .B(ori_ori_n1081_), .Y(ori_ori_n1082_));
  NO2        o1054(.A(ori_ori_n1032_), .B(ori_ori_n147_), .Y(ori_ori_n1083_));
  NOi21      o1055(.An(d), .B(f), .Y(ori_ori_n1084_));
  NA2        o1056(.A(h), .B(ori_ori_n1083_), .Y(ori_ori_n1085_));
  INV        o1057(.A(ori_ori_n240_), .Y(ori_ori_n1086_));
  NA2        o1058(.A(ori_ori_n1086_), .B(ori_ori_n446_), .Y(ori_ori_n1087_));
  NA2        o1059(.A(ori_ori_n1087_), .B(ori_ori_n1085_), .Y(ori_ori_n1088_));
  NO2        o1060(.A(ori_ori_n1088_), .B(ori_ori_n1082_), .Y(ori_ori_n1089_));
  NA3        o1061(.A(ori_ori_n1089_), .B(ori_ori_n1080_), .C(ori_ori_n1075_), .Y(ori_ori_n1090_));
  NA2        o1062(.A(h), .B(ori_ori_n1042_), .Y(ori_ori_n1091_));
  OAI210     o1063(.A0(ori_ori_n1062_), .A1(ori_ori_n1038_), .B0(ori_ori_n723_), .Y(ori_ori_n1092_));
  NA2        o1064(.A(ori_ori_n1092_), .B(ori_ori_n1091_), .Y(ori_ori_n1093_));
  NA2        o1065(.A(ori_ori_n1047_), .B(ori_ori_n1084_), .Y(ori_ori_n1094_));
  NO2        o1066(.A(ori_ori_n1094_), .B(m), .Y(ori_ori_n1095_));
  NO2        o1067(.A(ori_ori_n125_), .B(ori_ori_n154_), .Y(ori_ori_n1096_));
  OAI210     o1068(.A0(ori_ori_n1096_), .A1(ori_ori_n94_), .B0(ori_ori_n1050_), .Y(ori_ori_n1097_));
  INV        o1069(.A(ori_ori_n1097_), .Y(ori_ori_n1098_));
  NO3        o1070(.A(ori_ori_n1098_), .B(ori_ori_n1095_), .C(ori_ori_n1093_), .Y(ori_ori_n1099_));
  NA2        o1071(.A(ori_ori_n875_), .B(ori_ori_n522_), .Y(ori_ori_n1100_));
  OR2        o1072(.A(h), .B(ori_ori_n444_), .Y(ori_ori_n1101_));
  NO2        o1073(.A(ori_ori_n1101_), .B(ori_ori_n147_), .Y(ori_ori_n1102_));
  NA2        o1074(.A(ori_ori_n865_), .B(ori_ori_n189_), .Y(ori_ori_n1103_));
  NO2        o1075(.A(ori_ori_n48_), .B(l), .Y(ori_ori_n1104_));
  INV        o1076(.A(ori_ori_n398_), .Y(ori_ori_n1105_));
  NA2        o1077(.A(ori_ori_n1105_), .B(ori_ori_n1104_), .Y(ori_ori_n1106_));
  NA2        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1103_), .Y(ori_ori_n1107_));
  NO3        o1079(.A(ori_ori_n1107_), .B(ori_ori_n1102_), .C(ori_ori_n1046_), .Y(ori_ori_n1108_));
  NA3        o1080(.A(ori_ori_n1108_), .B(ori_ori_n1100_), .C(ori_ori_n1099_), .Y(ori_ori_n1109_));
  NA3        o1081(.A(ori_ori_n791_), .B(ori_ori_n115_), .C(ori_ori_n45_), .Y(ori_ori_n1110_));
  NO2        o1082(.A(ori_ori_n1065_), .B(d), .Y(ori_ori_n1111_));
  INV        o1083(.A(ori_ori_n1111_), .Y(ori_ori_n1112_));
  NA3        o1084(.A(ori_ori_n1112_), .B(ori_ori_n1118_), .C(ori_ori_n1110_), .Y(ori_ori_n1113_));
  OR4        o1085(.A(ori_ori_n1113_), .B(ori_ori_n1109_), .C(ori_ori_n1090_), .D(ori_ori_n1067_), .Y(ori04));
  INV        o1086(.A(ori_ori_n97_), .Y(ori_ori_n1117_));
  INV        o1087(.A(ori_ori_n1039_), .Y(ori_ori_n1118_));
  INV        o1088(.A(ori_ori_n86_), .Y(ori_ori_n1119_));
  INV        o1089(.A(ori_ori_n48_), .Y(ori_ori_n1120_));
  ZERO       o1090(.Y(ori02));
  ZERO       o1091(.Y(ori03));
  ZERO       o1092(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  INV        m0014(.A(i), .Y(mai_mai_n43_));
  AN2        m0015(.A(h), .B(g), .Y(mai_mai_n44_));
  NAi21      m0016(.An(n), .B(m), .Y(mai_mai_n45_));
  NOi32      m0017(.An(k), .Bn(h), .C(l), .Y(mai_mai_n46_));
  NOi32      m0018(.An(k), .Bn(h), .C(g), .Y(mai_mai_n47_));
  INV        m0019(.A(mai_mai_n47_), .Y(mai_mai_n48_));
  NO2        m0020(.A(mai_mai_n48_), .B(mai_mai_n45_), .Y(mai_mai_n49_));
  NO2        m0021(.A(mai_mai_n49_), .B(mai_mai_n39_), .Y(mai_mai_n50_));
  AOI210     m0022(.A0(mai_mai_n50_), .A1(mai_mai_n35_), .B0(mai_mai_n32_), .Y(mai_mai_n51_));
  INV        m0023(.A(c), .Y(mai_mai_n52_));
  NA2        m0024(.A(e), .B(b), .Y(mai_mai_n53_));
  NO2        m0025(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  INV        m0026(.A(d), .Y(mai_mai_n55_));
  NAi21      m0027(.An(i), .B(h), .Y(mai_mai_n56_));
  NAi31      m0028(.An(i), .B(l), .C(j), .Y(mai_mai_n57_));
  NAi41      m0029(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n58_));
  NA2        m0030(.A(g), .B(f), .Y(mai_mai_n59_));
  NO2        m0031(.A(mai_mai_n59_), .B(mai_mai_n58_), .Y(mai_mai_n60_));
  NAi21      m0032(.An(i), .B(j), .Y(mai_mai_n61_));
  NAi32      m0033(.An(n), .Bn(k), .C(m), .Y(mai_mai_n62_));
  NO2        m0034(.A(mai_mai_n62_), .B(mai_mai_n61_), .Y(mai_mai_n63_));
  NAi21      m0035(.An(e), .B(h), .Y(mai_mai_n64_));
  NAi41      m0036(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n65_));
  NA2        m0037(.A(mai_mai_n63_), .B(mai_mai_n60_), .Y(mai_mai_n66_));
  INV        m0038(.A(m), .Y(mai_mai_n67_));
  NOi21      m0039(.An(k), .B(l), .Y(mai_mai_n68_));
  NA2        m0040(.A(mai_mai_n68_), .B(mai_mai_n67_), .Y(mai_mai_n69_));
  AN4        m0041(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n70_));
  NOi31      m0042(.An(h), .B(g), .C(f), .Y(mai_mai_n71_));
  NA2        m0043(.A(mai_mai_n71_), .B(mai_mai_n70_), .Y(mai_mai_n72_));
  NAi32      m0044(.An(m), .Bn(k), .C(j), .Y(mai_mai_n73_));
  NOi32      m0045(.An(h), .Bn(g), .C(f), .Y(mai_mai_n74_));
  INV        m0046(.A(mai_mai_n66_), .Y(mai_mai_n75_));
  INV        m0047(.A(n), .Y(mai_mai_n76_));
  NOi32      m0048(.An(e), .Bn(b), .C(d), .Y(mai_mai_n77_));
  NA2        m0049(.A(mai_mai_n77_), .B(mai_mai_n76_), .Y(mai_mai_n78_));
  INV        m0050(.A(j), .Y(mai_mai_n79_));
  AN3        m0051(.A(m), .B(k), .C(i), .Y(mai_mai_n80_));
  NA3        m0052(.A(mai_mai_n80_), .B(mai_mai_n79_), .C(g), .Y(mai_mai_n81_));
  NAi32      m0053(.An(g), .Bn(f), .C(h), .Y(mai_mai_n82_));
  NAi31      m0054(.An(j), .B(m), .C(l), .Y(mai_mai_n83_));
  NO2        m0055(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  NA2        m0056(.A(m), .B(l), .Y(mai_mai_n85_));
  NAi31      m0057(.An(k), .B(j), .C(g), .Y(mai_mai_n86_));
  NO3        m0058(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(f), .Y(mai_mai_n87_));
  AN2        m0059(.A(j), .B(g), .Y(mai_mai_n88_));
  NOi32      m0060(.An(m), .Bn(l), .C(i), .Y(mai_mai_n89_));
  NOi21      m0061(.An(g), .B(i), .Y(mai_mai_n90_));
  NOi32      m0062(.An(m), .Bn(j), .C(k), .Y(mai_mai_n91_));
  AOI220     m0063(.A0(mai_mai_n91_), .A1(mai_mai_n90_), .B0(mai_mai_n89_), .B1(mai_mai_n88_), .Y(mai_mai_n92_));
  NAi41      m0064(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n93_));
  AN2        m0065(.A(e), .B(b), .Y(mai_mai_n94_));
  NOi31      m0066(.An(c), .B(h), .C(f), .Y(mai_mai_n95_));
  NA2        m0067(.A(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  NO3        m0068(.A(mai_mai_n96_), .B(mai_mai_n93_), .C(g), .Y(mai_mai_n97_));
  NOi21      m0069(.An(g), .B(f), .Y(mai_mai_n98_));
  NOi21      m0070(.An(i), .B(h), .Y(mai_mai_n99_));
  NA3        m0071(.A(mai_mai_n99_), .B(mai_mai_n98_), .C(mai_mai_n36_), .Y(mai_mai_n100_));
  INV        m0072(.A(a), .Y(mai_mai_n101_));
  NA2        m0073(.A(mai_mai_n94_), .B(mai_mai_n101_), .Y(mai_mai_n102_));
  INV        m0074(.A(l), .Y(mai_mai_n103_));
  NOi21      m0075(.An(m), .B(n), .Y(mai_mai_n104_));
  AN2        m0076(.A(k), .B(h), .Y(mai_mai_n105_));
  NO2        m0077(.A(mai_mai_n100_), .B(mai_mai_n78_), .Y(mai_mai_n106_));
  INV        m0078(.A(b), .Y(mai_mai_n107_));
  NA2        m0079(.A(l), .B(j), .Y(mai_mai_n108_));
  AN2        m0080(.A(k), .B(i), .Y(mai_mai_n109_));
  NA2        m0081(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NA2        m0082(.A(g), .B(e), .Y(mai_mai_n111_));
  NOi32      m0083(.An(c), .Bn(a), .C(d), .Y(mai_mai_n112_));
  NA2        m0084(.A(mai_mai_n112_), .B(mai_mai_n104_), .Y(mai_mai_n113_));
  NO4        m0085(.A(mai_mai_n113_), .B(mai_mai_n111_), .C(mai_mai_n110_), .D(mai_mai_n107_), .Y(mai_mai_n114_));
  NO3        m0086(.A(mai_mai_n114_), .B(mai_mai_n106_), .C(mai_mai_n97_), .Y(mai_mai_n115_));
  OAI210     m0087(.A0(mai_mai_n92_), .A1(mai_mai_n78_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  NOi31      m0088(.An(k), .B(m), .C(j), .Y(mai_mai_n117_));
  NOi31      m0089(.An(k), .B(m), .C(i), .Y(mai_mai_n118_));
  NOi32      m0090(.An(f), .Bn(b), .C(e), .Y(mai_mai_n119_));
  NAi21      m0091(.An(g), .B(h), .Y(mai_mai_n120_));
  NAi21      m0092(.An(m), .B(n), .Y(mai_mai_n121_));
  NAi21      m0093(.An(j), .B(k), .Y(mai_mai_n122_));
  NO3        m0094(.A(mai_mai_n122_), .B(mai_mai_n121_), .C(mai_mai_n120_), .Y(mai_mai_n123_));
  NAi41      m0095(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n124_));
  NAi31      m0096(.An(j), .B(k), .C(h), .Y(mai_mai_n125_));
  NO3        m0097(.A(mai_mai_n125_), .B(mai_mai_n124_), .C(mai_mai_n121_), .Y(mai_mai_n126_));
  AOI210     m0098(.A0(mai_mai_n123_), .A1(mai_mai_n119_), .B0(mai_mai_n126_), .Y(mai_mai_n127_));
  NO2        m0099(.A(k), .B(j), .Y(mai_mai_n128_));
  NO2        m0100(.A(mai_mai_n128_), .B(mai_mai_n121_), .Y(mai_mai_n129_));
  AN2        m0101(.A(k), .B(j), .Y(mai_mai_n130_));
  NAi21      m0102(.An(c), .B(b), .Y(mai_mai_n131_));
  NA2        m0103(.A(f), .B(d), .Y(mai_mai_n132_));
  NO4        m0104(.A(mai_mai_n132_), .B(mai_mai_n131_), .C(mai_mai_n130_), .D(mai_mai_n120_), .Y(mai_mai_n133_));
  NAi31      m0105(.An(f), .B(e), .C(b), .Y(mai_mai_n134_));
  NA2        m0106(.A(mai_mai_n133_), .B(mai_mai_n129_), .Y(mai_mai_n135_));
  NA2        m0107(.A(d), .B(b), .Y(mai_mai_n136_));
  NAi21      m0108(.An(e), .B(f), .Y(mai_mai_n137_));
  NA2        m0109(.A(b), .B(a), .Y(mai_mai_n138_));
  NAi21      m0110(.An(c), .B(d), .Y(mai_mai_n139_));
  NAi31      m0111(.An(l), .B(k), .C(h), .Y(mai_mai_n140_));
  NA2        m0112(.A(mai_mai_n135_), .B(mai_mai_n127_), .Y(mai_mai_n141_));
  NAi31      m0113(.An(e), .B(f), .C(b), .Y(mai_mai_n142_));
  NOi21      m0114(.An(g), .B(d), .Y(mai_mai_n143_));
  NO2        m0115(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NOi21      m0116(.An(h), .B(i), .Y(mai_mai_n145_));
  NOi21      m0117(.An(k), .B(m), .Y(mai_mai_n146_));
  NA3        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .C(n), .Y(mai_mai_n147_));
  NOi21      m0119(.An(h), .B(g), .Y(mai_mai_n148_));
  NO2        m0120(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n149_));
  NA2        m0121(.A(mai_mai_n149_), .B(mai_mai_n148_), .Y(mai_mai_n150_));
  NOi32      m0122(.An(n), .Bn(k), .C(m), .Y(mai_mai_n151_));
  NA2        m0123(.A(l), .B(i), .Y(mai_mai_n152_));
  NA2        m0124(.A(mai_mai_n152_), .B(mai_mai_n151_), .Y(mai_mai_n153_));
  NO2        m0125(.A(mai_mai_n153_), .B(mai_mai_n150_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(c), .Y(mai_mai_n155_));
  INV        m0127(.A(mai_mai_n155_), .Y(mai_mai_n156_));
  NA2        m0128(.A(j), .B(h), .Y(mai_mai_n157_));
  OR3        m0129(.A(n), .B(m), .C(k), .Y(mai_mai_n158_));
  NO2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NAi32      m0131(.An(m), .Bn(k), .C(n), .Y(mai_mai_n160_));
  NO2        m0132(.A(mai_mai_n160_), .B(mai_mai_n157_), .Y(mai_mai_n161_));
  AOI220     m0133(.A0(mai_mai_n161_), .A1(mai_mai_n144_), .B0(mai_mai_n159_), .B1(mai_mai_n156_), .Y(mai_mai_n162_));
  NO2        m0134(.A(n), .B(m), .Y(mai_mai_n163_));
  NAi21      m0135(.An(f), .B(e), .Y(mai_mai_n164_));
  NA2        m0136(.A(d), .B(c), .Y(mai_mai_n165_));
  NAi21      m0137(.An(d), .B(c), .Y(mai_mai_n166_));
  NAi31      m0138(.An(m), .B(n), .C(b), .Y(mai_mai_n167_));
  NA2        m0139(.A(k), .B(i), .Y(mai_mai_n168_));
  NAi21      m0140(.An(h), .B(f), .Y(mai_mai_n169_));
  NO2        m0141(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NO2        m0142(.A(mai_mai_n167_), .B(mai_mai_n139_), .Y(mai_mai_n171_));
  NA2        m0143(.A(mai_mai_n171_), .B(mai_mai_n170_), .Y(mai_mai_n172_));
  NOi32      m0144(.An(f), .Bn(c), .C(d), .Y(mai_mai_n173_));
  NOi32      m0145(.An(f), .Bn(c), .C(e), .Y(mai_mai_n174_));
  NO2        m0146(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NO3        m0147(.A(n), .B(m), .C(j), .Y(mai_mai_n176_));
  NA2        m0148(.A(mai_mai_n176_), .B(mai_mai_n105_), .Y(mai_mai_n177_));
  NA2        m0149(.A(mai_mai_n172_), .B(mai_mai_n162_), .Y(mai_mai_n178_));
  OR3        m0150(.A(mai_mai_n178_), .B(mai_mai_n154_), .C(mai_mai_n141_), .Y(mai_mai_n179_));
  NO4        m0151(.A(mai_mai_n179_), .B(mai_mai_n116_), .C(mai_mai_n75_), .D(mai_mai_n51_), .Y(mai_mai_n180_));
  NAi31      m0152(.An(n), .B(h), .C(g), .Y(mai_mai_n181_));
  NOi32      m0153(.An(m), .Bn(k), .C(l), .Y(mai_mai_n182_));
  NA3        m0154(.A(mai_mai_n182_), .B(mai_mai_n79_), .C(g), .Y(mai_mai_n183_));
  INV        m0155(.A(mai_mai_n183_), .Y(mai_mai_n184_));
  NOi21      m0156(.An(k), .B(j), .Y(mai_mai_n185_));
  NA4        m0157(.A(mai_mai_n185_), .B(mai_mai_n104_), .C(i), .D(g), .Y(mai_mai_n186_));
  AN2        m0158(.A(i), .B(g), .Y(mai_mai_n187_));
  NA3        m0159(.A(mai_mai_n68_), .B(mai_mai_n187_), .C(mai_mai_n104_), .Y(mai_mai_n188_));
  NA2        m0160(.A(mai_mai_n188_), .B(mai_mai_n186_), .Y(mai_mai_n189_));
  NAi41      m0161(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n190_));
  INV        m0162(.A(mai_mai_n190_), .Y(mai_mai_n191_));
  INV        m0163(.A(f), .Y(mai_mai_n192_));
  INV        m0164(.A(g), .Y(mai_mai_n193_));
  NOi31      m0165(.An(i), .B(j), .C(h), .Y(mai_mai_n194_));
  NOi21      m0166(.An(l), .B(m), .Y(mai_mai_n195_));
  NA2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NO3        m0168(.A(mai_mai_n196_), .B(mai_mai_n193_), .C(mai_mai_n192_), .Y(mai_mai_n197_));
  NA2        m0169(.A(mai_mai_n197_), .B(mai_mai_n191_), .Y(mai_mai_n198_));
  OAI210     m0170(.A0(mai_mai_n188_), .A1(mai_mai_n32_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  NOi21      m0171(.An(n), .B(m), .Y(mai_mai_n200_));
  NOi32      m0172(.An(l), .Bn(i), .C(j), .Y(mai_mai_n201_));
  NA2        m0173(.A(mai_mai_n201_), .B(mai_mai_n200_), .Y(mai_mai_n202_));
  OA220      m0174(.A0(mai_mai_n202_), .A1(mai_mai_n96_), .B0(mai_mai_n73_), .B1(mai_mai_n72_), .Y(mai_mai_n203_));
  NAi21      m0175(.An(j), .B(h), .Y(mai_mai_n204_));
  XN2        m0176(.A(i), .B(h), .Y(mai_mai_n205_));
  NA2        m0177(.A(mai_mai_n205_), .B(mai_mai_n204_), .Y(mai_mai_n206_));
  NOi31      m0178(.An(k), .B(n), .C(m), .Y(mai_mai_n207_));
  NOi31      m0179(.An(mai_mai_n207_), .B(mai_mai_n165_), .C(mai_mai_n164_), .Y(mai_mai_n208_));
  NA2        m0180(.A(mai_mai_n208_), .B(mai_mai_n206_), .Y(mai_mai_n209_));
  NAi31      m0181(.An(f), .B(e), .C(c), .Y(mai_mai_n210_));
  NO4        m0182(.A(mai_mai_n210_), .B(mai_mai_n158_), .C(mai_mai_n157_), .D(mai_mai_n55_), .Y(mai_mai_n211_));
  NA4        m0183(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n212_));
  NAi32      m0184(.An(m), .Bn(i), .C(k), .Y(mai_mai_n213_));
  NO3        m0185(.A(mai_mai_n213_), .B(mai_mai_n82_), .C(mai_mai_n212_), .Y(mai_mai_n214_));
  NO2        m0186(.A(mai_mai_n214_), .B(mai_mai_n211_), .Y(mai_mai_n215_));
  NAi21      m0187(.An(n), .B(a), .Y(mai_mai_n216_));
  NO2        m0188(.A(mai_mai_n216_), .B(mai_mai_n136_), .Y(mai_mai_n217_));
  NAi41      m0189(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n218_));
  NO2        m0190(.A(mai_mai_n218_), .B(e), .Y(mai_mai_n219_));
  NO3        m0191(.A(mai_mai_n137_), .B(mai_mai_n86_), .C(mai_mai_n85_), .Y(mai_mai_n220_));
  OAI210     m0192(.A0(mai_mai_n220_), .A1(mai_mai_n219_), .B0(mai_mai_n217_), .Y(mai_mai_n221_));
  AN4        m0193(.A(mai_mai_n221_), .B(mai_mai_n215_), .C(mai_mai_n209_), .D(mai_mai_n203_), .Y(mai_mai_n222_));
  OR2        m0194(.A(h), .B(g), .Y(mai_mai_n223_));
  NO2        m0195(.A(mai_mai_n223_), .B(mai_mai_n93_), .Y(mai_mai_n224_));
  NA2        m0196(.A(mai_mai_n224_), .B(mai_mai_n119_), .Y(mai_mai_n225_));
  NA2        m0197(.A(mai_mai_n146_), .B(mai_mai_n99_), .Y(mai_mai_n226_));
  NO2        m0198(.A(n), .B(a), .Y(mai_mai_n227_));
  NAi31      m0199(.An(mai_mai_n218_), .B(mai_mai_n227_), .C(mai_mai_n94_), .Y(mai_mai_n228_));
  NAi21      m0200(.An(h), .B(i), .Y(mai_mai_n229_));
  NA2        m0201(.A(mai_mai_n163_), .B(k), .Y(mai_mai_n230_));
  NO2        m0202(.A(mai_mai_n230_), .B(mai_mai_n229_), .Y(mai_mai_n231_));
  NA2        m0203(.A(mai_mai_n228_), .B(mai_mai_n225_), .Y(mai_mai_n232_));
  NOi21      m0204(.An(g), .B(e), .Y(mai_mai_n233_));
  NO2        m0205(.A(mai_mai_n65_), .B(mai_mai_n67_), .Y(mai_mai_n234_));
  NA2        m0206(.A(mai_mai_n234_), .B(mai_mai_n233_), .Y(mai_mai_n235_));
  NOi32      m0207(.An(l), .Bn(j), .C(i), .Y(mai_mai_n236_));
  AOI210     m0208(.A0(mai_mai_n68_), .A1(mai_mai_n79_), .B0(mai_mai_n236_), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n229_), .B(n), .Y(mai_mai_n238_));
  NAi21      m0210(.An(f), .B(g), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(mai_mai_n58_), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n62_), .B(mai_mai_n108_), .Y(mai_mai_n241_));
  AOI220     m0213(.A0(mai_mai_n241_), .A1(mai_mai_n240_), .B0(mai_mai_n238_), .B1(mai_mai_n60_), .Y(mai_mai_n242_));
  OAI210     m0214(.A0(mai_mai_n237_), .A1(mai_mai_n235_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  NOi41      m0215(.An(mai_mai_n222_), .B(mai_mai_n243_), .C(mai_mai_n232_), .D(mai_mai_n199_), .Y(mai_mai_n244_));
  INV        m0216(.A(mai_mai_n39_), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n245_), .B(mai_mai_n102_), .Y(mai_mai_n246_));
  NAi21      m0218(.An(h), .B(g), .Y(mai_mai_n247_));
  NO2        m0219(.A(mai_mai_n226_), .B(mai_mai_n239_), .Y(mai_mai_n248_));
  NA2        m0220(.A(mai_mai_n248_), .B(mai_mai_n70_), .Y(mai_mai_n249_));
  NAi31      m0221(.An(g), .B(k), .C(h), .Y(mai_mai_n250_));
  NO3        m0222(.A(mai_mai_n121_), .B(mai_mai_n250_), .C(l), .Y(mai_mai_n251_));
  NAi31      m0223(.An(e), .B(d), .C(a), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n251_), .B(mai_mai_n119_), .Y(mai_mai_n253_));
  NA2        m0225(.A(mai_mai_n253_), .B(mai_mai_n249_), .Y(mai_mai_n254_));
  NA4        m0226(.A(mai_mai_n146_), .B(mai_mai_n74_), .C(mai_mai_n70_), .D(mai_mai_n108_), .Y(mai_mai_n255_));
  NA3        m0227(.A(mai_mai_n146_), .B(mai_mai_n145_), .C(mai_mai_n76_), .Y(mai_mai_n256_));
  NO2        m0228(.A(mai_mai_n256_), .B(mai_mai_n175_), .Y(mai_mai_n257_));
  NOi21      m0229(.An(mai_mai_n255_), .B(mai_mai_n257_), .Y(mai_mai_n258_));
  NA3        m0230(.A(e), .B(c), .C(b), .Y(mai_mai_n259_));
  NAi21      m0231(.An(l), .B(k), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n260_), .B(mai_mai_n45_), .Y(mai_mai_n261_));
  NOi21      m0233(.An(l), .B(j), .Y(mai_mai_n262_));
  NA2        m0234(.A(mai_mai_n148_), .B(mai_mai_n262_), .Y(mai_mai_n263_));
  NA3        m0235(.A(mai_mai_n109_), .B(mai_mai_n108_), .C(g), .Y(mai_mai_n264_));
  OR3        m0236(.A(mai_mai_n65_), .B(mai_mai_n67_), .C(e), .Y(mai_mai_n265_));
  AOI210     m0237(.A0(mai_mai_n264_), .A1(mai_mai_n263_), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  INV        m0238(.A(mai_mai_n266_), .Y(mai_mai_n267_));
  NAi32      m0239(.An(j), .Bn(h), .C(i), .Y(mai_mai_n268_));
  NAi21      m0240(.An(m), .B(l), .Y(mai_mai_n269_));
  NO3        m0241(.A(mai_mai_n269_), .B(mai_mai_n268_), .C(mai_mai_n76_), .Y(mai_mai_n270_));
  NA2        m0242(.A(h), .B(g), .Y(mai_mai_n271_));
  NA2        m0243(.A(mai_mai_n270_), .B(mai_mai_n149_), .Y(mai_mai_n272_));
  NA3        m0244(.A(mai_mai_n272_), .B(mai_mai_n267_), .C(mai_mai_n258_), .Y(mai_mai_n273_));
  NO2        m0245(.A(mai_mai_n134_), .B(d), .Y(mai_mai_n274_));
  NA2        m0246(.A(mai_mai_n274_), .B(mai_mai_n49_), .Y(mai_mai_n275_));
  NO2        m0247(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n276_));
  NAi32      m0248(.An(n), .Bn(m), .C(l), .Y(mai_mai_n277_));
  NO2        m0249(.A(mai_mai_n277_), .B(mai_mai_n268_), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n113_), .B(mai_mai_n107_), .Y(mai_mai_n279_));
  NAi31      m0251(.An(k), .B(l), .C(j), .Y(mai_mai_n280_));
  OAI210     m0252(.A0(mai_mai_n260_), .A1(j), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  NOi21      m0253(.An(mai_mai_n281_), .B(mai_mai_n111_), .Y(mai_mai_n282_));
  NA2        m0254(.A(mai_mai_n282_), .B(mai_mai_n279_), .Y(mai_mai_n283_));
  NA2        m0255(.A(mai_mai_n283_), .B(mai_mai_n275_), .Y(mai_mai_n284_));
  NO4        m0256(.A(mai_mai_n284_), .B(mai_mai_n273_), .C(mai_mai_n254_), .D(mai_mai_n246_), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n231_), .B(mai_mai_n174_), .Y(mai_mai_n286_));
  NAi21      m0258(.An(m), .B(k), .Y(mai_mai_n287_));
  NAi41      m0259(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n288_));
  NA2        m0260(.A(e), .B(c), .Y(mai_mai_n289_));
  NA2        m0261(.A(f), .B(mai_mai_n109_), .Y(mai_mai_n290_));
  NO2        m0262(.A(mai_mai_n290_), .B(mai_mai_n193_), .Y(mai_mai_n291_));
  NAi31      m0263(.An(d), .B(e), .C(b), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n121_), .B(mai_mai_n292_), .Y(mai_mai_n293_));
  NA2        m0265(.A(mai_mai_n293_), .B(mai_mai_n291_), .Y(mai_mai_n294_));
  NA2        m0266(.A(mai_mai_n294_), .B(mai_mai_n286_), .Y(mai_mai_n295_));
  NO4        m0267(.A(mai_mai_n288_), .B(mai_mai_n73_), .C(mai_mai_n64_), .D(mai_mai_n193_), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n227_), .B(mai_mai_n94_), .Y(mai_mai_n297_));
  OR2        m0269(.A(mai_mai_n297_), .B(mai_mai_n183_), .Y(mai_mai_n298_));
  NOi31      m0270(.An(l), .B(n), .C(m), .Y(mai_mai_n299_));
  NA2        m0271(.A(mai_mai_n299_), .B(mai_mai_n194_), .Y(mai_mai_n300_));
  NO2        m0272(.A(mai_mai_n300_), .B(mai_mai_n175_), .Y(mai_mai_n301_));
  NAi32      m0273(.An(mai_mai_n301_), .Bn(mai_mai_n296_), .C(mai_mai_n298_), .Y(mai_mai_n302_));
  NAi32      m0274(.An(m), .Bn(j), .C(k), .Y(mai_mai_n303_));
  NAi41      m0275(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n190_), .B(mai_mai_n304_), .Y(mai_mai_n305_));
  NOi31      m0277(.An(j), .B(m), .C(k), .Y(mai_mai_n306_));
  NO2        m0278(.A(mai_mai_n117_), .B(mai_mai_n306_), .Y(mai_mai_n307_));
  AN3        m0279(.A(h), .B(g), .C(f), .Y(mai_mai_n308_));
  NAi31      m0280(.An(mai_mai_n307_), .B(mai_mai_n308_), .C(mai_mai_n305_), .Y(mai_mai_n309_));
  NOi32      m0281(.An(m), .Bn(j), .C(l), .Y(mai_mai_n310_));
  NO2        m0282(.A(mai_mai_n310_), .B(mai_mai_n89_), .Y(mai_mai_n311_));
  NAi32      m0283(.An(mai_mai_n311_), .Bn(mai_mai_n181_), .C(mai_mai_n274_), .Y(mai_mai_n312_));
  NO2        m0284(.A(mai_mai_n269_), .B(mai_mai_n268_), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n196_), .B(g), .Y(mai_mai_n314_));
  INV        m0286(.A(mai_mai_n142_), .Y(mai_mai_n315_));
  INV        m0287(.A(mai_mai_n213_), .Y(mai_mai_n316_));
  NA3        m0288(.A(mai_mai_n316_), .B(mai_mai_n308_), .C(mai_mai_n191_), .Y(mai_mai_n317_));
  NA3        m0289(.A(mai_mai_n317_), .B(mai_mai_n312_), .C(mai_mai_n309_), .Y(mai_mai_n318_));
  NA3        m0290(.A(h), .B(g), .C(f), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n319_), .B(mai_mai_n69_), .Y(mai_mai_n320_));
  INV        m0292(.A(mai_mai_n304_), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n148_), .B(e), .Y(mai_mai_n322_));
  NO2        m0294(.A(mai_mai_n322_), .B(mai_mai_n41_), .Y(mai_mai_n323_));
  AOI220     m0295(.A0(mai_mai_n323_), .A1(mai_mai_n279_), .B0(mai_mai_n321_), .B1(mai_mai_n320_), .Y(mai_mai_n324_));
  NOi32      m0296(.An(j), .Bn(g), .C(i), .Y(mai_mai_n325_));
  NA3        m0297(.A(mai_mai_n325_), .B(mai_mai_n260_), .C(mai_mai_n104_), .Y(mai_mai_n326_));
  OR2        m0298(.A(mai_mai_n102_), .B(mai_mai_n326_), .Y(mai_mai_n327_));
  NOi32      m0299(.An(e), .Bn(b), .C(a), .Y(mai_mai_n328_));
  AN2        m0300(.A(l), .B(j), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n287_), .B(mai_mai_n329_), .Y(mai_mai_n330_));
  NO3        m0302(.A(mai_mai_n288_), .B(mai_mai_n64_), .C(mai_mai_n193_), .Y(mai_mai_n331_));
  NA3        m0303(.A(mai_mai_n188_), .B(mai_mai_n186_), .C(mai_mai_n35_), .Y(mai_mai_n332_));
  AOI220     m0304(.A0(mai_mai_n332_), .A1(mai_mai_n328_), .B0(mai_mai_n331_), .B1(mai_mai_n330_), .Y(mai_mai_n333_));
  NO2        m0305(.A(mai_mai_n292_), .B(n), .Y(mai_mai_n334_));
  NA2        m0306(.A(mai_mai_n187_), .B(k), .Y(mai_mai_n335_));
  NA3        m0307(.A(m), .B(mai_mai_n103_), .C(mai_mai_n192_), .Y(mai_mai_n336_));
  NA4        m0308(.A(mai_mai_n182_), .B(mai_mai_n79_), .C(g), .D(mai_mai_n192_), .Y(mai_mai_n337_));
  INV        m0309(.A(mai_mai_n337_), .Y(mai_mai_n338_));
  NAi41      m0310(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n339_));
  NA2        m0311(.A(mai_mai_n47_), .B(mai_mai_n104_), .Y(mai_mai_n340_));
  NO2        m0312(.A(mai_mai_n340_), .B(mai_mai_n339_), .Y(mai_mai_n341_));
  AOI220     m0313(.A0(mai_mai_n341_), .A1(b), .B0(mai_mai_n338_), .B1(mai_mai_n334_), .Y(mai_mai_n342_));
  NA4        m0314(.A(mai_mai_n342_), .B(mai_mai_n333_), .C(mai_mai_n327_), .D(mai_mai_n324_), .Y(mai_mai_n343_));
  NO4        m0315(.A(mai_mai_n343_), .B(mai_mai_n318_), .C(mai_mai_n302_), .D(mai_mai_n295_), .Y(mai_mai_n344_));
  NA4        m0316(.A(mai_mai_n344_), .B(mai_mai_n285_), .C(mai_mai_n244_), .D(mai_mai_n180_), .Y(mai10));
  NA3        m0317(.A(m), .B(k), .C(i), .Y(mai_mai_n346_));
  NO3        m0318(.A(mai_mai_n346_), .B(j), .C(mai_mai_n193_), .Y(mai_mai_n347_));
  NOi21      m0319(.An(e), .B(f), .Y(mai_mai_n348_));
  NO4        m0320(.A(mai_mai_n139_), .B(mai_mai_n348_), .C(n), .D(mai_mai_n101_), .Y(mai_mai_n349_));
  NAi31      m0321(.An(b), .B(f), .C(c), .Y(mai_mai_n350_));
  INV        m0322(.A(mai_mai_n350_), .Y(mai_mai_n351_));
  NOi32      m0323(.An(k), .Bn(h), .C(j), .Y(mai_mai_n352_));
  NA2        m0324(.A(mai_mai_n352_), .B(mai_mai_n200_), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n147_), .B(mai_mai_n353_), .Y(mai_mai_n354_));
  AOI220     m0326(.A0(mai_mai_n354_), .A1(mai_mai_n351_), .B0(mai_mai_n349_), .B1(mai_mai_n347_), .Y(mai_mai_n355_));
  AN2        m0327(.A(j), .B(h), .Y(mai_mai_n356_));
  NO3        m0328(.A(n), .B(m), .C(k), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n357_), .B(mai_mai_n356_), .Y(mai_mai_n358_));
  NO3        m0330(.A(mai_mai_n358_), .B(mai_mai_n139_), .C(mai_mai_n192_), .Y(mai_mai_n359_));
  OR2        m0331(.A(m), .B(k), .Y(mai_mai_n360_));
  NO2        m0332(.A(mai_mai_n157_), .B(mai_mai_n360_), .Y(mai_mai_n361_));
  NA4        m0333(.A(n), .B(f), .C(c), .D(mai_mai_n107_), .Y(mai_mai_n362_));
  NOi21      m0334(.An(mai_mai_n361_), .B(mai_mai_n362_), .Y(mai_mai_n363_));
  NOi32      m0335(.An(d), .Bn(a), .C(c), .Y(mai_mai_n364_));
  NA2        m0336(.A(mai_mai_n364_), .B(mai_mai_n164_), .Y(mai_mai_n365_));
  NAi21      m0337(.An(i), .B(g), .Y(mai_mai_n366_));
  NAi31      m0338(.An(k), .B(m), .C(j), .Y(mai_mai_n367_));
  NO3        m0339(.A(mai_mai_n367_), .B(mai_mai_n366_), .C(n), .Y(mai_mai_n368_));
  NOi21      m0340(.An(mai_mai_n368_), .B(mai_mai_n365_), .Y(mai_mai_n369_));
  NO3        m0341(.A(mai_mai_n369_), .B(mai_mai_n363_), .C(mai_mai_n359_), .Y(mai_mai_n370_));
  NO2        m0342(.A(mai_mai_n362_), .B(mai_mai_n269_), .Y(mai_mai_n371_));
  NOi32      m0343(.An(f), .Bn(d), .C(c), .Y(mai_mai_n372_));
  AOI220     m0344(.A0(mai_mai_n372_), .A1(mai_mai_n278_), .B0(mai_mai_n371_), .B1(mai_mai_n194_), .Y(mai_mai_n373_));
  NA3        m0345(.A(mai_mai_n373_), .B(mai_mai_n370_), .C(mai_mai_n355_), .Y(mai_mai_n374_));
  NO2        m0346(.A(mai_mai_n55_), .B(mai_mai_n107_), .Y(mai_mai_n375_));
  NA2        m0347(.A(mai_mai_n227_), .B(mai_mai_n375_), .Y(mai_mai_n376_));
  INV        m0348(.A(e), .Y(mai_mai_n377_));
  NA2        m0349(.A(mai_mai_n44_), .B(e), .Y(mai_mai_n378_));
  AN2        m0350(.A(g), .B(e), .Y(mai_mai_n379_));
  NA3        m0351(.A(mai_mai_n379_), .B(mai_mai_n182_), .C(i), .Y(mai_mai_n380_));
  OAI210     m0352(.A0(mai_mai_n81_), .A1(mai_mai_n377_), .B0(mai_mai_n380_), .Y(mai_mai_n381_));
  NO2        m0353(.A(mai_mai_n92_), .B(mai_mai_n377_), .Y(mai_mai_n382_));
  NO2        m0354(.A(mai_mai_n382_), .B(mai_mai_n381_), .Y(mai_mai_n383_));
  NOi32      m0355(.An(h), .Bn(e), .C(g), .Y(mai_mai_n384_));
  NA3        m0356(.A(mai_mai_n384_), .B(mai_mai_n262_), .C(m), .Y(mai_mai_n385_));
  NOi21      m0357(.An(g), .B(h), .Y(mai_mai_n386_));
  AN3        m0358(.A(m), .B(l), .C(i), .Y(mai_mai_n387_));
  NA3        m0359(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(e), .Y(mai_mai_n388_));
  AN3        m0360(.A(h), .B(g), .C(e), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n389_), .B(mai_mai_n89_), .Y(mai_mai_n390_));
  NO2        m0362(.A(mai_mai_n383_), .B(mai_mai_n376_), .Y(mai_mai_n391_));
  NA3        m0363(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n392_));
  NO2        m0364(.A(mai_mai_n392_), .B(mai_mai_n376_), .Y(mai_mai_n393_));
  NA3        m0365(.A(mai_mai_n364_), .B(mai_mai_n164_), .C(mai_mai_n76_), .Y(mai_mai_n394_));
  NAi31      m0366(.An(b), .B(c), .C(a), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n395_), .B(n), .Y(mai_mai_n396_));
  NA2        m0368(.A(mai_mai_n47_), .B(m), .Y(mai_mai_n397_));
  NO2        m0369(.A(mai_mai_n397_), .B(mai_mai_n137_), .Y(mai_mai_n398_));
  NA2        m0370(.A(mai_mai_n398_), .B(mai_mai_n396_), .Y(mai_mai_n399_));
  INV        m0371(.A(mai_mai_n399_), .Y(mai_mai_n400_));
  NO4        m0372(.A(mai_mai_n400_), .B(mai_mai_n393_), .C(mai_mai_n391_), .D(mai_mai_n374_), .Y(mai_mai_n401_));
  NA2        m0373(.A(i), .B(g), .Y(mai_mai_n402_));
  NO3        m0374(.A(mai_mai_n252_), .B(mai_mai_n402_), .C(c), .Y(mai_mai_n403_));
  NOi21      m0375(.An(a), .B(n), .Y(mai_mai_n404_));
  NOi21      m0376(.An(d), .B(c), .Y(mai_mai_n405_));
  NA2        m0377(.A(mai_mai_n405_), .B(mai_mai_n404_), .Y(mai_mai_n406_));
  NA3        m0378(.A(i), .B(g), .C(f), .Y(mai_mai_n407_));
  NA2        m0379(.A(mai_mai_n403_), .B(mai_mai_n261_), .Y(mai_mai_n408_));
  OR2        m0380(.A(n), .B(m), .Y(mai_mai_n409_));
  NO2        m0381(.A(mai_mai_n165_), .B(mai_mai_n137_), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n159_), .B(mai_mai_n410_), .Y(mai_mai_n411_));
  INV        m0383(.A(mai_mai_n340_), .Y(mai_mai_n412_));
  NA3        m0384(.A(mai_mai_n412_), .B(mai_mai_n328_), .C(d), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n395_), .B(mai_mai_n45_), .Y(mai_mai_n414_));
  NAi21      m0386(.An(k), .B(j), .Y(mai_mai_n415_));
  NAi21      m0387(.An(e), .B(d), .Y(mai_mai_n416_));
  INV        m0388(.A(mai_mai_n416_), .Y(mai_mai_n417_));
  NO2        m0389(.A(mai_mai_n230_), .B(mai_mai_n192_), .Y(mai_mai_n418_));
  NA3        m0390(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(mai_mai_n206_), .Y(mai_mai_n419_));
  NA3        m0391(.A(mai_mai_n419_), .B(mai_mai_n413_), .C(mai_mai_n411_), .Y(mai_mai_n420_));
  NO2        m0392(.A(mai_mai_n300_), .B(mai_mai_n192_), .Y(mai_mai_n421_));
  NA2        m0393(.A(mai_mai_n421_), .B(mai_mai_n417_), .Y(mai_mai_n422_));
  NOi31      m0394(.An(n), .B(m), .C(k), .Y(mai_mai_n423_));
  AOI220     m0395(.A0(mai_mai_n423_), .A1(mai_mai_n356_), .B0(mai_mai_n200_), .B1(mai_mai_n46_), .Y(mai_mai_n424_));
  NAi31      m0396(.An(g), .B(f), .C(c), .Y(mai_mai_n425_));
  OR3        m0397(.A(mai_mai_n425_), .B(mai_mai_n424_), .C(e), .Y(mai_mai_n426_));
  NA2        m0398(.A(mai_mai_n426_), .B(mai_mai_n422_), .Y(mai_mai_n427_));
  NOi41      m0399(.An(mai_mai_n408_), .B(mai_mai_n427_), .C(mai_mai_n420_), .D(mai_mai_n243_), .Y(mai_mai_n428_));
  NOi32      m0400(.An(c), .Bn(a), .C(b), .Y(mai_mai_n429_));
  NA2        m0401(.A(mai_mai_n429_), .B(mai_mai_n104_), .Y(mai_mai_n430_));
  INV        m0402(.A(mai_mai_n250_), .Y(mai_mai_n431_));
  AN2        m0403(.A(e), .B(d), .Y(mai_mai_n432_));
  NA2        m0404(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  NO2        m0405(.A(mai_mai_n120_), .B(mai_mai_n41_), .Y(mai_mai_n434_));
  NO2        m0406(.A(mai_mai_n59_), .B(e), .Y(mai_mai_n435_));
  NOi31      m0407(.An(j), .B(k), .C(i), .Y(mai_mai_n436_));
  INV        m0408(.A(mai_mai_n436_), .Y(mai_mai_n437_));
  AOI210     m0409(.A0(mai_mai_n434_), .A1(f), .B0(mai_mai_n435_), .Y(mai_mai_n438_));
  AOI210     m0410(.A0(mai_mai_n438_), .A1(mai_mai_n433_), .B0(mai_mai_n430_), .Y(mai_mai_n439_));
  NO2        m0411(.A(mai_mai_n189_), .B(mai_mai_n184_), .Y(mai_mai_n440_));
  NOi21      m0412(.An(a), .B(b), .Y(mai_mai_n441_));
  NA3        m0413(.A(e), .B(d), .C(c), .Y(mai_mai_n442_));
  NAi21      m0414(.An(mai_mai_n442_), .B(mai_mai_n441_), .Y(mai_mai_n443_));
  NO2        m0415(.A(mai_mai_n394_), .B(mai_mai_n183_), .Y(mai_mai_n444_));
  NOi21      m0416(.An(mai_mai_n443_), .B(mai_mai_n444_), .Y(mai_mai_n445_));
  AOI210     m0417(.A0(mai_mai_n245_), .A1(mai_mai_n440_), .B0(mai_mai_n445_), .Y(mai_mai_n446_));
  NO4        m0418(.A(mai_mai_n169_), .B(mai_mai_n93_), .C(mai_mai_n52_), .D(b), .Y(mai_mai_n447_));
  OR2        m0419(.A(k), .B(j), .Y(mai_mai_n448_));
  NA2        m0420(.A(l), .B(k), .Y(mai_mai_n449_));
  INV        m0421(.A(mai_mai_n255_), .Y(mai_mai_n450_));
  NA2        m0422(.A(mai_mai_n364_), .B(mai_mai_n104_), .Y(mai_mai_n451_));
  NO4        m0423(.A(mai_mai_n451_), .B(mai_mai_n86_), .C(mai_mai_n103_), .D(e), .Y(mai_mai_n452_));
  NO3        m0424(.A(mai_mai_n394_), .B(mai_mai_n83_), .C(mai_mai_n120_), .Y(mai_mai_n453_));
  NO3        m0425(.A(mai_mai_n453_), .B(mai_mai_n452_), .C(mai_mai_n450_), .Y(mai_mai_n454_));
  INV        m0426(.A(mai_mai_n454_), .Y(mai_mai_n455_));
  NO4        m0427(.A(mai_mai_n455_), .B(mai_mai_n447_), .C(mai_mai_n446_), .D(mai_mai_n439_), .Y(mai_mai_n456_));
  NA2        m0428(.A(mai_mai_n63_), .B(mai_mai_n60_), .Y(mai_mai_n457_));
  NAi31      m0429(.An(j), .B(l), .C(i), .Y(mai_mai_n458_));
  OAI210     m0430(.A0(mai_mai_n458_), .A1(mai_mai_n121_), .B0(mai_mai_n93_), .Y(mai_mai_n459_));
  NO3        m0431(.A(mai_mai_n365_), .B(mai_mai_n311_), .C(mai_mai_n181_), .Y(mai_mai_n460_));
  NO2        m0432(.A(mai_mai_n365_), .B(mai_mai_n340_), .Y(mai_mai_n461_));
  NO3        m0433(.A(mai_mai_n461_), .B(mai_mai_n460_), .C(mai_mai_n276_), .Y(mai_mai_n462_));
  NA3        m0434(.A(mai_mai_n462_), .B(mai_mai_n457_), .C(mai_mai_n222_), .Y(mai_mai_n463_));
  OAI210     m0435(.A0(mai_mai_n118_), .A1(mai_mai_n117_), .B0(n), .Y(mai_mai_n464_));
  NO2        m0436(.A(mai_mai_n464_), .B(mai_mai_n120_), .Y(mai_mai_n465_));
  OA210      m0437(.A0(mai_mai_n224_), .A1(mai_mai_n465_), .B0(mai_mai_n174_), .Y(mai_mai_n466_));
  XO2        m0438(.A(i), .B(h), .Y(mai_mai_n467_));
  NA3        m0439(.A(mai_mai_n467_), .B(mai_mai_n146_), .C(n), .Y(mai_mai_n468_));
  NAi41      m0440(.An(mai_mai_n270_), .B(mai_mai_n468_), .C(mai_mai_n424_), .D(mai_mai_n353_), .Y(mai_mai_n469_));
  NAi31      m0441(.An(c), .B(f), .C(d), .Y(mai_mai_n470_));
  AOI210     m0442(.A0(mai_mai_n256_), .A1(mai_mai_n177_), .B0(mai_mai_n470_), .Y(mai_mai_n471_));
  INV        m0443(.A(mai_mai_n471_), .Y(mai_mai_n472_));
  NA3        m0444(.A(mai_mai_n349_), .B(mai_mai_n89_), .C(mai_mai_n88_), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n207_), .B(mai_mai_n99_), .Y(mai_mai_n474_));
  NA3        m0446(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n475_));
  NO2        m0447(.A(mai_mai_n475_), .B(mai_mai_n406_), .Y(mai_mai_n476_));
  NO2        m0448(.A(mai_mai_n476_), .B(mai_mai_n266_), .Y(mai_mai_n477_));
  NA3        m0449(.A(mai_mai_n477_), .B(mai_mai_n473_), .C(mai_mai_n472_), .Y(mai_mai_n478_));
  NO3        m0450(.A(mai_mai_n478_), .B(mai_mai_n466_), .C(mai_mai_n463_), .Y(mai_mai_n479_));
  NA4        m0451(.A(mai_mai_n479_), .B(mai_mai_n456_), .C(mai_mai_n428_), .D(mai_mai_n401_), .Y(mai11));
  NO2        m0452(.A(mai_mai_n65_), .B(f), .Y(mai_mai_n481_));
  NA2        m0453(.A(j), .B(g), .Y(mai_mai_n482_));
  NAi31      m0454(.An(i), .B(m), .C(l), .Y(mai_mai_n483_));
  NA3        m0455(.A(m), .B(k), .C(j), .Y(mai_mai_n484_));
  OAI220     m0456(.A0(mai_mai_n484_), .A1(mai_mai_n120_), .B0(mai_mai_n483_), .B1(mai_mai_n482_), .Y(mai_mai_n485_));
  NOi32      m0457(.An(e), .Bn(b), .C(f), .Y(mai_mai_n486_));
  NA2        m0458(.A(mai_mai_n236_), .B(mai_mai_n104_), .Y(mai_mai_n487_));
  NA2        m0459(.A(mai_mai_n44_), .B(j), .Y(mai_mai_n488_));
  NAi31      m0460(.An(d), .B(e), .C(a), .Y(mai_mai_n489_));
  NO2        m0461(.A(mai_mai_n489_), .B(n), .Y(mai_mai_n490_));
  NAi41      m0462(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n491_));
  AN2        m0463(.A(mai_mai_n491_), .B(mai_mai_n339_), .Y(mai_mai_n492_));
  NA2        m0464(.A(j), .B(i), .Y(mai_mai_n493_));
  NAi31      m0465(.An(n), .B(m), .C(k), .Y(mai_mai_n494_));
  NO3        m0466(.A(mai_mai_n494_), .B(mai_mai_n493_), .C(mai_mai_n103_), .Y(mai_mai_n495_));
  NO4        m0467(.A(n), .B(d), .C(mai_mai_n107_), .D(a), .Y(mai_mai_n496_));
  OR2        m0468(.A(n), .B(c), .Y(mai_mai_n497_));
  NO2        m0469(.A(mai_mai_n497_), .B(mai_mai_n138_), .Y(mai_mai_n498_));
  NO2        m0470(.A(mai_mai_n498_), .B(mai_mai_n496_), .Y(mai_mai_n499_));
  NOi32      m0471(.An(g), .Bn(f), .C(i), .Y(mai_mai_n500_));
  NA2        m0472(.A(mai_mai_n485_), .B(f), .Y(mai_mai_n501_));
  NO2        m0473(.A(mai_mai_n250_), .B(mai_mai_n45_), .Y(mai_mai_n502_));
  NO2        m0474(.A(mai_mai_n501_), .B(mai_mai_n499_), .Y(mai_mai_n503_));
  INV        m0475(.A(mai_mai_n503_), .Y(mai_mai_n504_));
  NA2        m0476(.A(mai_mai_n130_), .B(mai_mai_n34_), .Y(mai_mai_n505_));
  OAI220     m0477(.A0(mai_mai_n505_), .A1(m), .B0(mai_mai_n488_), .B1(mai_mai_n213_), .Y(mai_mai_n506_));
  NOi41      m0478(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n507_));
  AN2        m0479(.A(mai_mai_n304_), .B(mai_mai_n288_), .Y(mai_mai_n508_));
  AN2        m0480(.A(mai_mai_n507_), .B(mai_mai_n506_), .Y(mai_mai_n509_));
  OAI220     m0481(.A0(mai_mai_n367_), .A1(mai_mai_n366_), .B0(mai_mai_n483_), .B1(mai_mai_n482_), .Y(mai_mai_n510_));
  NAi31      m0482(.An(d), .B(c), .C(a), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n511_), .B(n), .Y(mai_mai_n512_));
  NA3        m0484(.A(mai_mai_n512_), .B(mai_mai_n510_), .C(e), .Y(mai_mai_n513_));
  NO3        m0485(.A(mai_mai_n57_), .B(mai_mai_n45_), .C(mai_mai_n193_), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n210_), .B(mai_mai_n101_), .Y(mai_mai_n515_));
  OAI210     m0487(.A0(mai_mai_n514_), .A1(mai_mai_n368_), .B0(mai_mai_n515_), .Y(mai_mai_n516_));
  NA2        m0488(.A(mai_mai_n516_), .B(mai_mai_n513_), .Y(mai_mai_n517_));
  NO2        m0489(.A(mai_mai_n252_), .B(n), .Y(mai_mai_n518_));
  NO2        m0490(.A(mai_mai_n396_), .B(mai_mai_n518_), .Y(mai_mai_n519_));
  NA2        m0491(.A(mai_mai_n510_), .B(f), .Y(mai_mai_n520_));
  NAi32      m0492(.An(d), .Bn(a), .C(b), .Y(mai_mai_n521_));
  NO2        m0493(.A(mai_mai_n521_), .B(mai_mai_n45_), .Y(mai_mai_n522_));
  NA2        m0494(.A(h), .B(f), .Y(mai_mai_n523_));
  NO2        m0495(.A(mai_mai_n523_), .B(mai_mai_n86_), .Y(mai_mai_n524_));
  NO3        m0496(.A(mai_mai_n160_), .B(mai_mai_n157_), .C(g), .Y(mai_mai_n525_));
  AOI220     m0497(.A0(mai_mai_n525_), .A1(mai_mai_n54_), .B0(mai_mai_n524_), .B1(mai_mai_n522_), .Y(mai_mai_n526_));
  OAI210     m0498(.A0(mai_mai_n520_), .A1(mai_mai_n519_), .B0(mai_mai_n526_), .Y(mai_mai_n527_));
  AN3        m0499(.A(j), .B(h), .C(g), .Y(mai_mai_n528_));
  NO2        m0500(.A(mai_mai_n136_), .B(c), .Y(mai_mai_n529_));
  NA3        m0501(.A(mai_mai_n529_), .B(mai_mai_n528_), .C(mai_mai_n423_), .Y(mai_mai_n530_));
  NA3        m0502(.A(f), .B(d), .C(b), .Y(mai_mai_n531_));
  NO4        m0503(.A(mai_mai_n531_), .B(mai_mai_n160_), .C(mai_mai_n157_), .D(g), .Y(mai_mai_n532_));
  NAi21      m0504(.An(mai_mai_n532_), .B(mai_mai_n530_), .Y(mai_mai_n533_));
  NO4        m0505(.A(mai_mai_n533_), .B(mai_mai_n527_), .C(mai_mai_n517_), .D(mai_mai_n509_), .Y(mai_mai_n534_));
  AN2        m0506(.A(mai_mai_n534_), .B(mai_mai_n504_), .Y(mai_mai_n535_));
  INV        m0507(.A(k), .Y(mai_mai_n536_));
  NA3        m0508(.A(l), .B(mai_mai_n536_), .C(i), .Y(mai_mai_n537_));
  INV        m0509(.A(mai_mai_n537_), .Y(mai_mai_n538_));
  NAi32      m0510(.An(h), .Bn(f), .C(g), .Y(mai_mai_n539_));
  NAi41      m0511(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n540_));
  OAI210     m0512(.A0(mai_mai_n489_), .A1(n), .B0(mai_mai_n540_), .Y(mai_mai_n541_));
  NAi31      m0513(.An(h), .B(g), .C(f), .Y(mai_mai_n542_));
  OR3        m0514(.A(mai_mai_n542_), .B(mai_mai_n252_), .C(mai_mai_n45_), .Y(mai_mai_n543_));
  NA4        m0515(.A(mai_mai_n386_), .B(mai_mai_n112_), .C(mai_mai_n104_), .D(e), .Y(mai_mai_n544_));
  AN2        m0516(.A(mai_mai_n544_), .B(mai_mai_n543_), .Y(mai_mai_n545_));
  NO3        m0517(.A(mai_mai_n539_), .B(mai_mai_n65_), .C(mai_mai_n67_), .Y(mai_mai_n546_));
  NO4        m0518(.A(mai_mai_n542_), .B(mai_mai_n497_), .C(mai_mai_n138_), .D(mai_mai_n67_), .Y(mai_mai_n547_));
  OR2        m0519(.A(mai_mai_n547_), .B(mai_mai_n546_), .Y(mai_mai_n548_));
  NAi21      m0520(.An(mai_mai_n548_), .B(mai_mai_n545_), .Y(mai_mai_n549_));
  NAi31      m0521(.An(f), .B(h), .C(g), .Y(mai_mai_n550_));
  NO4        m0522(.A(mai_mai_n280_), .B(mai_mai_n550_), .C(mai_mai_n65_), .D(mai_mai_n67_), .Y(mai_mai_n551_));
  NOi32      m0523(.An(b), .Bn(a), .C(c), .Y(mai_mai_n552_));
  NOi41      m0524(.An(mai_mai_n552_), .B(mai_mai_n319_), .C(mai_mai_n62_), .D(mai_mai_n108_), .Y(mai_mai_n553_));
  OR2        m0525(.A(mai_mai_n553_), .B(mai_mai_n551_), .Y(mai_mai_n554_));
  NOi32      m0526(.An(d), .Bn(a), .C(e), .Y(mai_mai_n555_));
  NA2        m0527(.A(mai_mai_n555_), .B(mai_mai_n104_), .Y(mai_mai_n556_));
  NO2        m0528(.A(n), .B(c), .Y(mai_mai_n557_));
  NA3        m0529(.A(mai_mai_n557_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n558_));
  NOi32      m0530(.An(e), .Bn(a), .C(d), .Y(mai_mai_n559_));
  AOI210     m0531(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n559_), .Y(mai_mai_n560_));
  AOI210     m0532(.A0(mai_mai_n560_), .A1(mai_mai_n192_), .B0(mai_mai_n505_), .Y(mai_mai_n561_));
  AOI210     m0533(.A0(mai_mai_n561_), .A1(mai_mai_n104_), .B0(mai_mai_n554_), .Y(mai_mai_n562_));
  INV        m0534(.A(mai_mai_n562_), .Y(mai_mai_n563_));
  AOI210     m0535(.A0(mai_mai_n549_), .A1(mai_mai_n538_), .B0(mai_mai_n563_), .Y(mai_mai_n564_));
  NO3        m0536(.A(mai_mai_n287_), .B(mai_mai_n56_), .C(n), .Y(mai_mai_n565_));
  NA2        m0537(.A(mai_mai_n470_), .B(mai_mai_n155_), .Y(mai_mai_n566_));
  NA2        m0538(.A(mai_mai_n425_), .B(mai_mai_n210_), .Y(mai_mai_n567_));
  NA2        m0539(.A(mai_mai_n68_), .B(mai_mai_n104_), .Y(mai_mai_n568_));
  NA2        m0540(.A(mai_mai_n567_), .B(mai_mai_n565_), .Y(mai_mai_n569_));
  NO2        m0541(.A(mai_mai_n569_), .B(mai_mai_n79_), .Y(mai_mai_n570_));
  NOi32      m0542(.An(e), .Bn(c), .C(f), .Y(mai_mai_n571_));
  NOi21      m0543(.An(f), .B(g), .Y(mai_mai_n572_));
  NO2        m0544(.A(mai_mai_n572_), .B(mai_mai_n190_), .Y(mai_mai_n573_));
  AOI220     m0545(.A0(mai_mai_n573_), .A1(mai_mai_n361_), .B0(mai_mai_n571_), .B1(mai_mai_n159_), .Y(mai_mai_n574_));
  NA2        m0546(.A(mai_mai_n574_), .B(mai_mai_n162_), .Y(mai_mai_n575_));
  AOI210     m0547(.A0(mai_mai_n492_), .A1(mai_mai_n365_), .B0(mai_mai_n271_), .Y(mai_mai_n576_));
  NA2        m0548(.A(mai_mai_n576_), .B(mai_mai_n241_), .Y(mai_mai_n577_));
  NAi21      m0549(.An(k), .B(h), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n578_), .B(mai_mai_n239_), .Y(mai_mai_n579_));
  NOi31      m0551(.An(m), .B(n), .C(k), .Y(mai_mai_n580_));
  NA2        m0552(.A(j), .B(mai_mai_n580_), .Y(mai_mai_n581_));
  AOI210     m0553(.A0(mai_mai_n365_), .A1(mai_mai_n339_), .B0(mai_mai_n271_), .Y(mai_mai_n582_));
  NAi21      m0554(.An(mai_mai_n581_), .B(mai_mai_n582_), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n489_), .B(mai_mai_n45_), .Y(mai_mai_n584_));
  NA2        m0556(.A(mai_mai_n583_), .B(mai_mai_n577_), .Y(mai_mai_n585_));
  INV        m0557(.A(mai_mai_n328_), .Y(mai_mai_n586_));
  NO2        m0558(.A(mai_mai_n586_), .B(n), .Y(mai_mai_n587_));
  NA2        m0559(.A(mai_mai_n467_), .B(mai_mai_n146_), .Y(mai_mai_n588_));
  NO3        m0560(.A(mai_mai_n362_), .B(mai_mai_n588_), .C(mai_mai_n79_), .Y(mai_mai_n589_));
  INV        m0561(.A(mai_mai_n589_), .Y(mai_mai_n590_));
  AN3        m0562(.A(f), .B(d), .C(b), .Y(mai_mai_n591_));
  NO2        m0563(.A(mai_mai_n591_), .B(mai_mai_n119_), .Y(mai_mai_n592_));
  NA3        m0564(.A(mai_mai_n467_), .B(mai_mai_n146_), .C(mai_mai_n193_), .Y(mai_mai_n593_));
  AOI210     m0565(.A0(mai_mai_n592_), .A1(mai_mai_n212_), .B0(mai_mai_n593_), .Y(mai_mai_n594_));
  NAi31      m0566(.An(m), .B(n), .C(k), .Y(mai_mai_n595_));
  INV        m0567(.A(mai_mai_n228_), .Y(mai_mai_n596_));
  OAI210     m0568(.A0(mai_mai_n596_), .A1(mai_mai_n594_), .B0(j), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n597_), .B(mai_mai_n590_), .Y(mai_mai_n598_));
  NO4        m0570(.A(mai_mai_n598_), .B(mai_mai_n585_), .C(mai_mai_n575_), .D(mai_mai_n570_), .Y(mai_mai_n599_));
  NA2        m0571(.A(mai_mai_n349_), .B(mai_mai_n148_), .Y(mai_mai_n600_));
  NAi31      m0572(.An(g), .B(h), .C(f), .Y(mai_mai_n601_));
  OR3        m0573(.A(mai_mai_n601_), .B(mai_mai_n252_), .C(n), .Y(mai_mai_n602_));
  OA210      m0574(.A0(mai_mai_n489_), .A1(n), .B0(mai_mai_n540_), .Y(mai_mai_n603_));
  NA3        m0575(.A(mai_mai_n384_), .B(mai_mai_n112_), .C(mai_mai_n76_), .Y(mai_mai_n604_));
  OAI210     m0576(.A0(mai_mai_n603_), .A1(mai_mai_n82_), .B0(mai_mai_n604_), .Y(mai_mai_n605_));
  NOi21      m0577(.An(mai_mai_n602_), .B(mai_mai_n605_), .Y(mai_mai_n606_));
  AOI210     m0578(.A0(mai_mai_n606_), .A1(mai_mai_n600_), .B0(mai_mai_n484_), .Y(mai_mai_n607_));
  NO3        m0579(.A(g), .B(mai_mai_n192_), .C(mai_mai_n52_), .Y(mai_mai_n608_));
  NAi21      m0580(.An(h), .B(j), .Y(mai_mai_n609_));
  NO2        m0581(.A(mai_mai_n474_), .B(mai_mai_n79_), .Y(mai_mai_n610_));
  OAI210     m0582(.A0(mai_mai_n610_), .A1(mai_mai_n361_), .B0(mai_mai_n608_), .Y(mai_mai_n611_));
  NA3        m0583(.A(mai_mai_n481_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n612_));
  NA2        m0584(.A(h), .B(mai_mai_n37_), .Y(mai_mai_n613_));
  NA2        m0585(.A(mai_mai_n91_), .B(mai_mai_n44_), .Y(mai_mai_n614_));
  OAI220     m0586(.A0(mai_mai_n614_), .A1(mai_mai_n297_), .B0(mai_mai_n613_), .B1(mai_mai_n430_), .Y(mai_mai_n615_));
  AOI210     m0587(.A0(mai_mai_n521_), .A1(mai_mai_n395_), .B0(mai_mai_n45_), .Y(mai_mai_n616_));
  NO2        m0588(.A(mai_mai_n542_), .B(mai_mai_n537_), .Y(mai_mai_n617_));
  AOI210     m0589(.A0(mai_mai_n617_), .A1(mai_mai_n616_), .B0(mai_mai_n615_), .Y(mai_mai_n618_));
  NA3        m0590(.A(mai_mai_n618_), .B(mai_mai_n612_), .C(mai_mai_n611_), .Y(mai_mai_n619_));
  NO2        m0591(.A(mai_mai_n229_), .B(f), .Y(mai_mai_n620_));
  NO2        m0592(.A(mai_mai_n572_), .B(mai_mai_n56_), .Y(mai_mai_n621_));
  NO3        m0593(.A(mai_mai_n621_), .B(mai_mai_n620_), .C(mai_mai_n34_), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n293_), .B(mai_mai_n130_), .Y(mai_mai_n623_));
  AOI220     m0595(.A0(mai_mai_n1372_), .A1(mai_mai_n486_), .B0(mai_mai_n328_), .B1(mai_mai_n104_), .Y(mai_mai_n624_));
  OA220      m0596(.A0(mai_mai_n624_), .A1(mai_mai_n505_), .B0(mai_mai_n326_), .B1(mai_mai_n102_), .Y(mai_mai_n625_));
  OAI210     m0597(.A0(mai_mai_n623_), .A1(mai_mai_n622_), .B0(mai_mai_n625_), .Y(mai_mai_n626_));
  NO3        m0598(.A(mai_mai_n372_), .B(mai_mai_n174_), .C(mai_mai_n173_), .Y(mai_mai_n627_));
  NA2        m0599(.A(mai_mai_n627_), .B(mai_mai_n210_), .Y(mai_mai_n628_));
  NA3        m0600(.A(mai_mai_n628_), .B(mai_mai_n231_), .C(j), .Y(mai_mai_n629_));
  NO3        m0601(.A(mai_mai_n425_), .B(mai_mai_n157_), .C(i), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n429_), .B(mai_mai_n76_), .Y(mai_mai_n631_));
  NO4        m0603(.A(mai_mai_n484_), .B(mai_mai_n631_), .C(mai_mai_n120_), .D(mai_mai_n192_), .Y(mai_mai_n632_));
  INV        m0604(.A(mai_mai_n632_), .Y(mai_mai_n633_));
  NA4        m0605(.A(mai_mai_n633_), .B(mai_mai_n629_), .C(mai_mai_n473_), .D(mai_mai_n370_), .Y(mai_mai_n634_));
  NO4        m0606(.A(mai_mai_n634_), .B(mai_mai_n626_), .C(mai_mai_n619_), .D(mai_mai_n607_), .Y(mai_mai_n635_));
  NA4        m0607(.A(mai_mai_n635_), .B(mai_mai_n599_), .C(mai_mai_n564_), .D(mai_mai_n535_), .Y(mai08));
  NO2        m0608(.A(k), .B(h), .Y(mai_mai_n637_));
  AO210      m0609(.A0(mai_mai_n229_), .A1(mai_mai_n415_), .B0(mai_mai_n637_), .Y(mai_mai_n638_));
  NO2        m0610(.A(mai_mai_n638_), .B(mai_mai_n269_), .Y(mai_mai_n639_));
  NA2        m0611(.A(mai_mai_n571_), .B(mai_mai_n76_), .Y(mai_mai_n640_));
  NA2        m0612(.A(mai_mai_n640_), .B(mai_mai_n425_), .Y(mai_mai_n641_));
  AOI210     m0613(.A0(mai_mai_n641_), .A1(mai_mai_n639_), .B0(mai_mai_n453_), .Y(mai_mai_n642_));
  NA2        m0614(.A(mai_mai_n76_), .B(mai_mai_n101_), .Y(mai_mai_n643_));
  NO2        m0615(.A(mai_mai_n643_), .B(mai_mai_n53_), .Y(mai_mai_n644_));
  NO3        m0616(.A(mai_mai_n346_), .B(mai_mai_n103_), .C(mai_mai_n193_), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n531_), .B(mai_mai_n212_), .Y(mai_mai_n646_));
  AOI220     m0618(.A0(mai_mai_n646_), .A1(mai_mai_n314_), .B0(mai_mai_n645_), .B1(mai_mai_n644_), .Y(mai_mai_n647_));
  AOI210     m0619(.A0(mai_mai_n531_), .A1(mai_mai_n142_), .B0(mai_mai_n76_), .Y(mai_mai_n648_));
  NA4        m0620(.A(mai_mai_n195_), .B(mai_mai_n130_), .C(mai_mai_n43_), .D(h), .Y(mai_mai_n649_));
  AN2        m0621(.A(l), .B(k), .Y(mai_mai_n650_));
  NA4        m0622(.A(mai_mai_n650_), .B(mai_mai_n99_), .C(mai_mai_n67_), .D(mai_mai_n193_), .Y(mai_mai_n651_));
  OAI210     m0623(.A0(mai_mai_n649_), .A1(g), .B0(mai_mai_n651_), .Y(mai_mai_n652_));
  NA2        m0624(.A(mai_mai_n652_), .B(mai_mai_n648_), .Y(mai_mai_n653_));
  NA3        m0625(.A(mai_mai_n653_), .B(mai_mai_n647_), .C(mai_mai_n642_), .Y(mai_mai_n654_));
  NO4        m0626(.A(mai_mai_n157_), .B(mai_mai_n360_), .C(mai_mai_n103_), .D(g), .Y(mai_mai_n655_));
  AOI210     m0627(.A0(mai_mai_n655_), .A1(mai_mai_n646_), .B0(mai_mai_n476_), .Y(mai_mai_n656_));
  INV        m0628(.A(mai_mai_n656_), .Y(mai_mai_n657_));
  NO3        m0629(.A(mai_mai_n287_), .B(mai_mai_n120_), .C(mai_mai_n41_), .Y(mai_mai_n658_));
  BUFFER     m0630(.A(mai_mai_n658_), .Y(mai_mai_n659_));
  INV        m0631(.A(mai_mai_n638_), .Y(mai_mai_n660_));
  AOI220     m0632(.A0(mai_mai_n660_), .A1(mai_mai_n371_), .B0(mai_mai_n659_), .B1(mai_mai_n70_), .Y(mai_mai_n661_));
  INV        m0633(.A(mai_mai_n661_), .Y(mai_mai_n662_));
  NA3        m0634(.A(mai_mai_n628_), .B(mai_mai_n299_), .C(mai_mai_n352_), .Y(mai_mai_n663_));
  NA2        m0635(.A(mai_mai_n650_), .B(mai_mai_n200_), .Y(mai_mai_n664_));
  NO2        m0636(.A(mai_mai_n664_), .B(mai_mai_n292_), .Y(mai_mai_n665_));
  AOI210     m0637(.A0(mai_mai_n665_), .A1(mai_mai_n620_), .B0(mai_mai_n452_), .Y(mai_mai_n666_));
  NA3        m0638(.A(m), .B(l), .C(k), .Y(mai_mai_n667_));
  AOI210     m0639(.A0(mai_mai_n604_), .A1(mai_mai_n602_), .B0(mai_mai_n667_), .Y(mai_mai_n668_));
  NO2        m0640(.A(mai_mai_n491_), .B(mai_mai_n247_), .Y(mai_mai_n669_));
  NOi21      m0641(.An(mai_mai_n669_), .B(mai_mai_n487_), .Y(mai_mai_n670_));
  NA4        m0642(.A(mai_mai_n104_), .B(l), .C(k), .D(mai_mai_n79_), .Y(mai_mai_n671_));
  NA3        m0643(.A(mai_mai_n112_), .B(mai_mai_n379_), .C(i), .Y(mai_mai_n672_));
  NO2        m0644(.A(mai_mai_n672_), .B(mai_mai_n671_), .Y(mai_mai_n673_));
  NO3        m0645(.A(mai_mai_n673_), .B(mai_mai_n670_), .C(mai_mai_n668_), .Y(mai_mai_n674_));
  NA3        m0646(.A(mai_mai_n674_), .B(mai_mai_n666_), .C(mai_mai_n663_), .Y(mai_mai_n675_));
  NO4        m0647(.A(mai_mai_n675_), .B(mai_mai_n662_), .C(mai_mai_n657_), .D(mai_mai_n654_), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n573_), .B(mai_mai_n361_), .Y(mai_mai_n677_));
  NOi31      m0649(.An(g), .B(h), .C(f), .Y(mai_mai_n678_));
  NA2        m0650(.A(mai_mai_n584_), .B(mai_mai_n678_), .Y(mai_mai_n679_));
  AO210      m0651(.A0(mai_mai_n679_), .A1(mai_mai_n543_), .B0(mai_mai_n493_), .Y(mai_mai_n680_));
  INV        m0652(.A(mai_mai_n461_), .Y(mai_mai_n681_));
  NA4        m0653(.A(mai_mai_n681_), .B(mai_mai_n680_), .C(mai_mai_n677_), .D(mai_mai_n228_), .Y(mai_mai_n682_));
  NA2        m0654(.A(mai_mai_n650_), .B(mai_mai_n67_), .Y(mai_mai_n683_));
  NO3        m0655(.A(mai_mai_n627_), .B(mai_mai_n157_), .C(i), .Y(mai_mai_n684_));
  NOi21      m0656(.An(h), .B(j), .Y(mai_mai_n685_));
  NA2        m0657(.A(mai_mai_n685_), .B(f), .Y(mai_mai_n686_));
  NO2        m0658(.A(mai_mai_n684_), .B(mai_mai_n630_), .Y(mai_mai_n687_));
  OAI220     m0659(.A0(mai_mai_n687_), .A1(mai_mai_n683_), .B0(mai_mai_n545_), .B1(mai_mai_n57_), .Y(mai_mai_n688_));
  AOI210     m0660(.A0(mai_mai_n682_), .A1(l), .B0(mai_mai_n688_), .Y(mai_mai_n689_));
  NO2        m0661(.A(j), .B(i), .Y(mai_mai_n690_));
  NA2        m0662(.A(mai_mai_n690_), .B(mai_mai_n33_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n389_), .B(mai_mai_n112_), .Y(mai_mai_n692_));
  OR2        m0664(.A(mai_mai_n692_), .B(mai_mai_n691_), .Y(mai_mai_n693_));
  NO3        m0665(.A(mai_mai_n139_), .B(mai_mai_n45_), .C(mai_mai_n101_), .Y(mai_mai_n694_));
  NO3        m0666(.A(mai_mai_n497_), .B(mai_mai_n138_), .C(mai_mai_n67_), .Y(mai_mai_n695_));
  NO2        m0667(.A(mai_mai_n449_), .B(mai_mai_n407_), .Y(mai_mai_n696_));
  OAI210     m0668(.A0(mai_mai_n695_), .A1(mai_mai_n694_), .B0(mai_mai_n696_), .Y(mai_mai_n697_));
  OAI210     m0669(.A0(mai_mai_n679_), .A1(mai_mai_n57_), .B0(mai_mai_n697_), .Y(mai_mai_n698_));
  NA2        m0670(.A(k), .B(j), .Y(mai_mai_n699_));
  NAi31      m0671(.An(mai_mai_n560_), .B(mai_mai_n84_), .C(mai_mai_n76_), .Y(mai_mai_n700_));
  INV        m0672(.A(mai_mai_n700_), .Y(mai_mai_n701_));
  NO2        m0673(.A(mai_mai_n269_), .B(mai_mai_n125_), .Y(mai_mai_n702_));
  AOI220     m0674(.A0(mai_mai_n702_), .A1(mai_mai_n573_), .B0(mai_mai_n658_), .B1(mai_mai_n648_), .Y(mai_mai_n703_));
  NO2        m0675(.A(mai_mai_n667_), .B(mai_mai_n82_), .Y(mai_mai_n704_));
  NA2        m0676(.A(mai_mai_n704_), .B(mai_mai_n541_), .Y(mai_mai_n705_));
  NA2        m0677(.A(mai_mai_n705_), .B(mai_mai_n703_), .Y(mai_mai_n706_));
  OR3        m0678(.A(mai_mai_n706_), .B(mai_mai_n701_), .C(mai_mai_n698_), .Y(mai_mai_n707_));
  OAI220     m0679(.A0(mai_mai_n649_), .A1(mai_mai_n640_), .B0(mai_mai_n297_), .B1(mai_mai_n38_), .Y(mai_mai_n708_));
  INV        m0680(.A(mai_mai_n708_), .Y(mai_mai_n709_));
  NA3        m0681(.A(mai_mai_n500_), .B(mai_mai_n262_), .C(h), .Y(mai_mai_n710_));
  NOi21      m0682(.An(mai_mai_n616_), .B(mai_mai_n710_), .Y(mai_mai_n711_));
  NAi21      m0683(.An(mai_mai_n711_), .B(mai_mai_n709_), .Y(mai_mai_n712_));
  BUFFER     m0684(.A(mai_mai_n87_), .Y(mai_mai_n713_));
  NA2        m0685(.A(mai_mai_n713_), .B(mai_mai_n217_), .Y(mai_mai_n714_));
  INV        m0686(.A(mai_mai_n301_), .Y(mai_mai_n715_));
  OAI210     m0687(.A0(mai_mai_n667_), .A1(mai_mai_n601_), .B0(mai_mai_n475_), .Y(mai_mai_n716_));
  NA3        m0688(.A(mai_mai_n227_), .B(mai_mai_n55_), .C(b), .Y(mai_mai_n717_));
  AOI220     m0689(.A0(mai_mai_n557_), .A1(mai_mai_n29_), .B0(mai_mai_n429_), .B1(mai_mai_n76_), .Y(mai_mai_n718_));
  NA2        m0690(.A(mai_mai_n718_), .B(mai_mai_n717_), .Y(mai_mai_n719_));
  NO2        m0691(.A(mai_mai_n710_), .B(mai_mai_n451_), .Y(mai_mai_n720_));
  AOI210     m0692(.A0(mai_mai_n719_), .A1(mai_mai_n716_), .B0(mai_mai_n720_), .Y(mai_mai_n721_));
  NA3        m0693(.A(mai_mai_n721_), .B(mai_mai_n715_), .C(mai_mai_n714_), .Y(mai_mai_n722_));
  NOi41      m0694(.An(mai_mai_n693_), .B(mai_mai_n722_), .C(mai_mai_n712_), .D(mai_mai_n707_), .Y(mai_mai_n723_));
  OR3        m0695(.A(mai_mai_n649_), .B(mai_mai_n212_), .C(g), .Y(mai_mai_n724_));
  INV        m0696(.A(mai_mai_n44_), .Y(mai_mai_n725_));
  NO3        m0697(.A(mai_mai_n725_), .B(mai_mai_n691_), .C(mai_mai_n252_), .Y(mai_mai_n726_));
  NO3        m0698(.A(mai_mai_n482_), .B(mai_mai_n85_), .C(h), .Y(mai_mai_n727_));
  AOI210     m0699(.A0(mai_mai_n727_), .A1(mai_mai_n644_), .B0(mai_mai_n726_), .Y(mai_mai_n728_));
  NA3        m0700(.A(mai_mai_n728_), .B(mai_mai_n724_), .C(mai_mai_n373_), .Y(mai_mai_n729_));
  OR2        m0701(.A(mai_mai_n601_), .B(mai_mai_n83_), .Y(mai_mai_n730_));
  NOi31      m0702(.An(b), .B(d), .C(a), .Y(mai_mai_n731_));
  NO2        m0703(.A(mai_mai_n731_), .B(mai_mai_n555_), .Y(mai_mai_n732_));
  NO2        m0704(.A(mai_mai_n732_), .B(n), .Y(mai_mai_n733_));
  NOi21      m0705(.An(mai_mai_n718_), .B(mai_mai_n733_), .Y(mai_mai_n734_));
  NO2        m0706(.A(mai_mai_n734_), .B(mai_mai_n730_), .Y(mai_mai_n735_));
  NO3        m0707(.A(mai_mai_n572_), .B(mai_mai_n292_), .C(mai_mai_n108_), .Y(mai_mai_n736_));
  NOi21      m0708(.An(mai_mai_n736_), .B(mai_mai_n147_), .Y(mai_mai_n737_));
  INV        m0709(.A(mai_mai_n737_), .Y(mai_mai_n738_));
  OAI210     m0710(.A0(mai_mai_n649_), .A1(mai_mai_n362_), .B0(mai_mai_n738_), .Y(mai_mai_n739_));
  NO2        m0711(.A(mai_mai_n627_), .B(n), .Y(mai_mai_n740_));
  AOI220     m0712(.A0(mai_mai_n702_), .A1(mai_mai_n608_), .B0(mai_mai_n740_), .B1(mai_mai_n639_), .Y(mai_mai_n741_));
  NA2        m0713(.A(mai_mai_n112_), .B(mai_mai_n76_), .Y(mai_mai_n742_));
  AOI210     m0714(.A0(mai_mai_n392_), .A1(mai_mai_n385_), .B0(mai_mai_n742_), .Y(mai_mai_n743_));
  NA2        m0715(.A(mai_mai_n665_), .B(mai_mai_n34_), .Y(mai_mai_n744_));
  NAi21      m0716(.An(mai_mai_n671_), .B(mai_mai_n403_), .Y(mai_mai_n745_));
  NO2        m0717(.A(mai_mai_n247_), .B(i), .Y(mai_mai_n746_));
  NA2        m0718(.A(mai_mai_n655_), .B(mai_mai_n315_), .Y(mai_mai_n747_));
  OAI210     m0719(.A0(mai_mai_n547_), .A1(mai_mai_n546_), .B0(mai_mai_n329_), .Y(mai_mai_n748_));
  AN3        m0720(.A(mai_mai_n748_), .B(mai_mai_n747_), .C(mai_mai_n745_), .Y(mai_mai_n749_));
  NAi41      m0721(.An(mai_mai_n743_), .B(mai_mai_n749_), .C(mai_mai_n744_), .D(mai_mai_n741_), .Y(mai_mai_n750_));
  NO4        m0722(.A(mai_mai_n750_), .B(mai_mai_n739_), .C(mai_mai_n735_), .D(mai_mai_n729_), .Y(mai_mai_n751_));
  NA4        m0723(.A(mai_mai_n751_), .B(mai_mai_n723_), .C(mai_mai_n689_), .D(mai_mai_n676_), .Y(mai09));
  INV        m0724(.A(mai_mai_n113_), .Y(mai_mai_n753_));
  NA2        m0725(.A(f), .B(e), .Y(mai_mai_n754_));
  NO2        m0726(.A(g), .B(mai_mai_n434_), .Y(mai_mai_n755_));
  NO2        m0727(.A(mai_mai_n755_), .B(mai_mai_n754_), .Y(mai_mai_n756_));
  NA2        m0728(.A(mai_mai_n756_), .B(mai_mai_n753_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n183_), .B(mai_mai_n192_), .Y(mai_mai_n758_));
  NA3        m0730(.A(m), .B(l), .C(i), .Y(mai_mai_n759_));
  NA3        m0731(.A(mai_mai_n80_), .B(g), .C(f), .Y(mai_mai_n760_));
  INV        m0732(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  OR2        m0733(.A(mai_mai_n761_), .B(mai_mai_n758_), .Y(mai_mai_n762_));
  NA3        m0734(.A(mai_mai_n730_), .B(mai_mai_n520_), .C(mai_mai_n475_), .Y(mai_mai_n763_));
  OA210      m0735(.A0(mai_mai_n763_), .A1(mai_mai_n762_), .B0(mai_mai_n733_), .Y(mai_mai_n764_));
  INV        m0736(.A(mai_mai_n304_), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n766_));
  NOi31      m0738(.An(k), .B(m), .C(l), .Y(mai_mai_n767_));
  NO2        m0739(.A(mai_mai_n306_), .B(mai_mai_n767_), .Y(mai_mai_n768_));
  AOI210     m0740(.A0(mai_mai_n768_), .A1(mai_mai_n766_), .B0(mai_mai_n550_), .Y(mai_mai_n769_));
  NA2        m0741(.A(mai_mai_n769_), .B(mai_mai_n765_), .Y(mai_mai_n770_));
  NA2        m0742(.A(mai_mai_n152_), .B(mai_mai_n105_), .Y(mai_mai_n771_));
  NA3        m0743(.A(mai_mai_n771_), .B(mai_mai_n638_), .C(mai_mai_n125_), .Y(mai_mai_n772_));
  NA3        m0744(.A(mai_mai_n772_), .B(mai_mai_n171_), .C(mai_mai_n31_), .Y(mai_mai_n773_));
  NA3        m0745(.A(mai_mai_n773_), .B(mai_mai_n770_), .C(mai_mai_n574_), .Y(mai_mai_n774_));
  NO2        m0746(.A(mai_mai_n539_), .B(mai_mai_n458_), .Y(mai_mai_n775_));
  NA2        m0747(.A(mai_mai_n775_), .B(mai_mai_n171_), .Y(mai_mai_n776_));
  NOi21      m0748(.An(f), .B(d), .Y(mai_mai_n777_));
  NA2        m0749(.A(mai_mai_n777_), .B(m), .Y(mai_mai_n778_));
  NO2        m0750(.A(mai_mai_n778_), .B(mai_mai_n48_), .Y(mai_mai_n779_));
  NOi32      m0751(.An(g), .Bn(f), .C(d), .Y(mai_mai_n780_));
  NA4        m0752(.A(mai_mai_n780_), .B(mai_mai_n557_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n781_));
  NA2        m0753(.A(mai_mai_n779_), .B(mai_mai_n498_), .Y(mai_mai_n782_));
  AN2        m0754(.A(f), .B(d), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n441_), .B(mai_mai_n783_), .C(mai_mai_n76_), .Y(mai_mai_n784_));
  NO3        m0756(.A(mai_mai_n784_), .B(mai_mai_n67_), .C(mai_mai_n193_), .Y(mai_mai_n785_));
  NO2        m0757(.A(k), .B(mai_mai_n52_), .Y(mai_mai_n786_));
  INV        m0758(.A(mai_mai_n785_), .Y(mai_mai_n787_));
  NAi41      m0759(.An(mai_mai_n450_), .B(mai_mai_n787_), .C(mai_mai_n782_), .D(mai_mai_n776_), .Y(mai_mai_n788_));
  NO4        m0760(.A(mai_mai_n572_), .B(mai_mai_n121_), .C(mai_mai_n292_), .D(mai_mai_n140_), .Y(mai_mai_n789_));
  NO2        m0761(.A(mai_mai_n595_), .B(mai_mai_n292_), .Y(mai_mai_n790_));
  AN2        m0762(.A(mai_mai_n790_), .B(mai_mai_n620_), .Y(mai_mai_n791_));
  NO3        m0763(.A(mai_mai_n791_), .B(mai_mai_n789_), .C(mai_mai_n214_), .Y(mai_mai_n792_));
  NA2        m0764(.A(mai_mai_n555_), .B(mai_mai_n76_), .Y(mai_mai_n793_));
  NA3        m0765(.A(mai_mai_n146_), .B(mai_mai_n99_), .C(mai_mai_n98_), .Y(mai_mai_n794_));
  OAI220     m0766(.A0(mai_mai_n784_), .A1(mai_mai_n397_), .B0(mai_mai_n304_), .B1(mai_mai_n794_), .Y(mai_mai_n795_));
  NOi31      m0767(.An(mai_mai_n203_), .B(mai_mai_n795_), .C(mai_mai_n276_), .Y(mai_mai_n796_));
  NA2        m0768(.A(c), .B(mai_mai_n107_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n797_), .B(mai_mai_n377_), .Y(mai_mai_n798_));
  NA3        m0770(.A(mai_mai_n798_), .B(mai_mai_n469_), .C(f), .Y(mai_mai_n799_));
  OR2        m0771(.A(mai_mai_n601_), .B(mai_mai_n494_), .Y(mai_mai_n800_));
  INV        m0772(.A(mai_mai_n800_), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n732_), .B(mai_mai_n102_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n801_), .Y(mai_mai_n803_));
  NA4        m0775(.A(mai_mai_n803_), .B(mai_mai_n799_), .C(mai_mai_n796_), .D(mai_mai_n792_), .Y(mai_mai_n804_));
  NO4        m0776(.A(mai_mai_n804_), .B(mai_mai_n788_), .C(mai_mai_n774_), .D(mai_mai_n764_), .Y(mai_mai_n805_));
  BUFFER     m0777(.A(mai_mai_n784_), .Y(mai_mai_n806_));
  NA2        m0778(.A(mai_mai_n103_), .B(j), .Y(mai_mai_n807_));
  NO2        m0779(.A(mai_mai_n263_), .B(mai_mai_n806_), .Y(mai_mai_n808_));
  NO2        m0780(.A(mai_mai_n297_), .B(mai_mai_n760_), .Y(mai_mai_n809_));
  NO2        m0781(.A(mai_mai_n125_), .B(mai_mai_n121_), .Y(mai_mai_n810_));
  NO2        m0782(.A(mai_mai_n210_), .B(mai_mai_n204_), .Y(mai_mai_n811_));
  AOI220     m0783(.A0(mai_mai_n811_), .A1(mai_mai_n207_), .B0(mai_mai_n274_), .B1(mai_mai_n810_), .Y(mai_mai_n812_));
  NO2        m0784(.A(mai_mai_n397_), .B(mai_mai_n754_), .Y(mai_mai_n813_));
  NA2        m0785(.A(mai_mai_n813_), .B(mai_mai_n512_), .Y(mai_mai_n814_));
  NA2        m0786(.A(mai_mai_n814_), .B(mai_mai_n812_), .Y(mai_mai_n815_));
  NA2        m0787(.A(e), .B(d), .Y(mai_mai_n816_));
  OAI220     m0788(.A0(mai_mai_n816_), .A1(c), .B0(mai_mai_n289_), .B1(d), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n474_), .B(mai_mai_n210_), .Y(mai_mai_n818_));
  INV        m0790(.A(mai_mai_n818_), .Y(mai_mai_n819_));
  NA3        m0791(.A(mai_mai_n151_), .B(mai_mai_n77_), .C(mai_mai_n34_), .Y(mai_mai_n820_));
  NA2        m0792(.A(mai_mai_n820_), .B(mai_mai_n819_), .Y(mai_mai_n821_));
  NO4        m0793(.A(mai_mai_n821_), .B(mai_mai_n815_), .C(mai_mai_n809_), .D(mai_mai_n808_), .Y(mai_mai_n822_));
  NA2        m0794(.A(mai_mai_n765_), .B(mai_mai_n31_), .Y(mai_mai_n823_));
  OR2        m0795(.A(mai_mai_n823_), .B(mai_mai_n196_), .Y(mai_mai_n824_));
  OAI220     m0796(.A0(mai_mai_n572_), .A1(mai_mai_n56_), .B0(mai_mai_n271_), .B1(j), .Y(mai_mai_n825_));
  AOI220     m0797(.A0(mai_mai_n825_), .A1(mai_mai_n790_), .B0(mai_mai_n565_), .B1(mai_mai_n571_), .Y(mai_mai_n826_));
  INV        m0798(.A(mai_mai_n826_), .Y(mai_mai_n827_));
  AOI210     m0799(.A0(mai_mai_n109_), .A1(mai_mai_n108_), .B0(mai_mai_n236_), .Y(mai_mai_n828_));
  NO2        m0800(.A(mai_mai_n828_), .B(mai_mai_n781_), .Y(mai_mai_n829_));
  BUFFER     m0801(.A(mai_mai_n829_), .Y(mai_mai_n830_));
  NO2        m0802(.A(mai_mai_n830_), .B(mai_mai_n827_), .Y(mai_mai_n831_));
  AO220      m0803(.A0(mai_mai_n418_), .A1(mai_mai_n685_), .B0(mai_mai_n159_), .B1(f), .Y(mai_mai_n832_));
  OAI210     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n421_), .B0(mai_mai_n817_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n763_), .B(mai_mai_n644_), .Y(mai_mai_n834_));
  AN4        m0806(.A(mai_mai_n834_), .B(mai_mai_n833_), .C(mai_mai_n831_), .D(mai_mai_n824_), .Y(mai_mai_n835_));
  NA4        m0807(.A(mai_mai_n835_), .B(mai_mai_n822_), .C(mai_mai_n805_), .D(mai_mai_n757_), .Y(mai12));
  NO2        m0808(.A(mai_mai_n416_), .B(c), .Y(mai_mai_n837_));
  NO4        m0809(.A(mai_mai_n409_), .B(mai_mai_n229_), .C(mai_mai_n536_), .D(mai_mai_n193_), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n838_), .B(mai_mai_n837_), .Y(mai_mai_n839_));
  NO2        m0811(.A(mai_mai_n601_), .B(mai_mai_n346_), .Y(mai_mai_n840_));
  NA2        m0812(.A(mai_mai_n840_), .B(mai_mai_n496_), .Y(mai_mai_n841_));
  NA3        m0813(.A(mai_mai_n841_), .B(mai_mai_n839_), .C(mai_mai_n408_), .Y(mai_mai_n842_));
  AOI210     m0814(.A0(mai_mai_n213_), .A1(mai_mai_n303_), .B0(mai_mai_n181_), .Y(mai_mai_n843_));
  BUFFER     m0815(.A(mai_mai_n843_), .Y(mai_mai_n844_));
  AOI210     m0816(.A0(mai_mai_n300_), .A1(mai_mai_n358_), .B0(mai_mai_n193_), .Y(mai_mai_n845_));
  OAI210     m0817(.A0(mai_mai_n845_), .A1(mai_mai_n844_), .B0(mai_mai_n372_), .Y(mai_mai_n846_));
  NO2        m0818(.A(mai_mai_n542_), .B(mai_mai_n759_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n847_), .B(mai_mai_n518_), .Y(mai_mai_n848_));
  NO2        m0820(.A(mai_mai_n139_), .B(mai_mai_n216_), .Y(mai_mai_n849_));
  NA3        m0821(.A(mai_mai_n849_), .B(mai_mai_n219_), .C(i), .Y(mai_mai_n850_));
  NA3        m0822(.A(mai_mai_n850_), .B(mai_mai_n848_), .C(mai_mai_n846_), .Y(mai_mai_n851_));
  NO3        m0823(.A(mai_mai_n121_), .B(mai_mai_n140_), .C(mai_mai_n193_), .Y(mai_mai_n852_));
  NA2        m0824(.A(mai_mai_n852_), .B(mai_mai_n486_), .Y(mai_mai_n853_));
  INV        m0825(.A(mai_mai_n853_), .Y(mai_mai_n854_));
  NO3        m0826(.A(mai_mai_n606_), .B(mai_mai_n83_), .C(mai_mai_n43_), .Y(mai_mai_n855_));
  NO4        m0827(.A(mai_mai_n855_), .B(mai_mai_n854_), .C(mai_mai_n851_), .D(mai_mai_n842_), .Y(mai_mai_n856_));
  NO2        m0828(.A(mai_mai_n336_), .B(mai_mai_n335_), .Y(mai_mai_n857_));
  NA2        m0829(.A(mai_mai_n540_), .B(mai_mai_n65_), .Y(mai_mai_n858_));
  INV        m0830(.A(mai_mai_n134_), .Y(mai_mai_n859_));
  NOi21      m0831(.An(mai_mai_n34_), .B(mai_mai_n595_), .Y(mai_mai_n860_));
  AOI220     m0832(.A0(mai_mai_n860_), .A1(mai_mai_n859_), .B0(mai_mai_n858_), .B1(mai_mai_n857_), .Y(mai_mai_n861_));
  OAI210     m0833(.A0(mai_mai_n228_), .A1(mai_mai_n43_), .B0(mai_mai_n861_), .Y(mai_mai_n862_));
  NA2        m0834(.A(mai_mai_n403_), .B(mai_mai_n241_), .Y(mai_mai_n863_));
  NO3        m0835(.A(mai_mai_n742_), .B(mai_mai_n81_), .C(mai_mai_n377_), .Y(mai_mai_n864_));
  NAi21      m0836(.An(mai_mai_n864_), .B(mai_mai_n863_), .Y(mai_mai_n865_));
  NO2        m0837(.A(mai_mai_n45_), .B(mai_mai_n43_), .Y(mai_mai_n866_));
  NA2        m0838(.A(mai_mai_n580_), .B(mai_mai_n329_), .Y(mai_mai_n867_));
  OAI210     m0839(.A0(mai_mai_n672_), .A1(mai_mai_n867_), .B0(mai_mai_n333_), .Y(mai_mai_n868_));
  NO3        m0840(.A(mai_mai_n868_), .B(mai_mai_n865_), .C(mai_mai_n862_), .Y(mai_mai_n869_));
  NA2        m0841(.A(mai_mai_n313_), .B(g), .Y(mai_mai_n870_));
  NA2        m0842(.A(mai_mai_n148_), .B(i), .Y(mai_mai_n871_));
  NA2        m0843(.A(mai_mai_n44_), .B(i), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n387_), .B(mai_mai_n37_), .Y(mai_mai_n873_));
  NO2        m0845(.A(mai_mai_n134_), .B(mai_mai_n76_), .Y(mai_mai_n874_));
  OR2        m0846(.A(mai_mai_n874_), .B(mai_mai_n507_), .Y(mai_mai_n875_));
  INV        m0847(.A(mai_mai_n875_), .Y(mai_mai_n876_));
  OAI220     m0848(.A0(mai_mai_n876_), .A1(mai_mai_n870_), .B0(mai_mai_n873_), .B1(mai_mai_n297_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n601_), .B(mai_mai_n458_), .Y(mai_mai_n878_));
  NA3        m0850(.A(mai_mai_n308_), .B(j), .C(i), .Y(mai_mai_n879_));
  INV        m0851(.A(mai_mai_n879_), .Y(mai_mai_n880_));
  OAI220     m0852(.A0(mai_mai_n880_), .A1(mai_mai_n878_), .B0(mai_mai_n616_), .B1(mai_mai_n695_), .Y(mai_mai_n881_));
  OR3        m0853(.A(mai_mai_n280_), .B(mai_mai_n402_), .C(f), .Y(mai_mai_n882_));
  NA2        m0854(.A(mai_mai_n631_), .B(mai_mai_n793_), .Y(mai_mai_n883_));
  INV        m0855(.A(mai_mai_n760_), .Y(mai_mai_n884_));
  NA2        m0856(.A(mai_mai_n201_), .B(mai_mai_n71_), .Y(mai_mai_n885_));
  NA2        m0857(.A(mai_mai_n885_), .B(mai_mai_n882_), .Y(mai_mai_n886_));
  AOI220     m0858(.A0(mai_mai_n886_), .A1(mai_mai_n234_), .B0(mai_mai_n884_), .B1(mai_mai_n883_), .Y(mai_mai_n887_));
  NA2        m0859(.A(mai_mai_n887_), .B(mai_mai_n881_), .Y(mai_mai_n888_));
  NA2        m0860(.A(mai_mai_n605_), .B(mai_mai_n80_), .Y(mai_mai_n889_));
  NO2        m0861(.A(mai_mai_n424_), .B(mai_mai_n193_), .Y(mai_mai_n890_));
  NA2        m0862(.A(mai_mai_n890_), .B(mai_mai_n351_), .Y(mai_mai_n891_));
  NA2        m0863(.A(mai_mai_n840_), .B(mai_mai_n849_), .Y(mai_mai_n892_));
  NA3        m0864(.A(mai_mai_n892_), .B(mai_mai_n891_), .C(mai_mai_n889_), .Y(mai_mai_n893_));
  OAI210     m0865(.A0(mai_mai_n884_), .A1(mai_mai_n847_), .B0(mai_mai_n496_), .Y(mai_mai_n894_));
  AOI210     m0866(.A0(mai_mai_n388_), .A1(mai_mai_n380_), .B0(mai_mai_n742_), .Y(mai_mai_n895_));
  OAI210     m0867(.A0(mai_mai_n336_), .A1(mai_mai_n335_), .B0(mai_mai_n100_), .Y(mai_mai_n896_));
  AOI210     m0868(.A0(mai_mai_n896_), .A1(mai_mai_n490_), .B0(mai_mai_n895_), .Y(mai_mai_n897_));
  NO3        m0869(.A(mai_mai_n807_), .B(mai_mai_n45_), .C(mai_mai_n43_), .Y(mai_mai_n898_));
  NA2        m0870(.A(mai_mai_n898_), .B(mai_mai_n576_), .Y(mai_mai_n899_));
  NA3        m0871(.A(mai_mai_n899_), .B(mai_mai_n897_), .C(mai_mai_n894_), .Y(mai_mai_n900_));
  NO4        m0872(.A(mai_mai_n900_), .B(mai_mai_n893_), .C(mai_mai_n888_), .D(mai_mai_n877_), .Y(mai_mai_n901_));
  NAi31      m0873(.An(mai_mai_n131_), .B(mai_mai_n389_), .C(n), .Y(mai_mai_n902_));
  NO3        m0874(.A(mai_mai_n117_), .B(mai_mai_n306_), .C(mai_mai_n767_), .Y(mai_mai_n903_));
  NO2        m0875(.A(mai_mai_n903_), .B(mai_mai_n902_), .Y(mai_mai_n904_));
  NO3        m0876(.A(mai_mai_n247_), .B(mai_mai_n131_), .C(mai_mai_n377_), .Y(mai_mai_n905_));
  AOI210     m0877(.A0(mai_mai_n905_), .A1(mai_mai_n459_), .B0(mai_mai_n904_), .Y(mai_mai_n906_));
  NA2        m0878(.A(mai_mai_n453_), .B(i), .Y(mai_mai_n907_));
  NA2        m0879(.A(mai_mai_n907_), .B(mai_mai_n906_), .Y(mai_mai_n908_));
  NA2        m0880(.A(mai_mai_n210_), .B(mai_mai_n155_), .Y(mai_mai_n909_));
  NO2        m0881(.A(mai_mai_n278_), .B(mai_mai_n159_), .Y(mai_mai_n910_));
  NOi31      m0882(.An(mai_mai_n909_), .B(mai_mai_n910_), .C(mai_mai_n193_), .Y(mai_mai_n911_));
  NA2        m0883(.A(mai_mai_n406_), .B(mai_mai_n793_), .Y(mai_mai_n912_));
  NO2        m0884(.A(mai_mai_n407_), .B(mai_mai_n280_), .Y(mai_mai_n913_));
  AOI220     m0885(.A0(mai_mai_n913_), .A1(mai_mai_n912_), .B0(mai_mai_n447_), .B1(g), .Y(mai_mai_n914_));
  INV        m0886(.A(mai_mai_n914_), .Y(mai_mai_n915_));
  OAI220     m0887(.A0(mai_mai_n902_), .A1(mai_mai_n213_), .B0(mai_mai_n879_), .B1(mai_mai_n556_), .Y(mai_mai_n916_));
  NO2        m0888(.A(mai_mai_n602_), .B(mai_mai_n346_), .Y(mai_mai_n917_));
  NA2        m0889(.A(mai_mai_n843_), .B(mai_mai_n837_), .Y(mai_mai_n918_));
  NO3        m0890(.A(mai_mai_n497_), .B(mai_mai_n138_), .C(mai_mai_n192_), .Y(mai_mai_n919_));
  OAI210     m0891(.A0(mai_mai_n919_), .A1(mai_mai_n481_), .B0(mai_mai_n347_), .Y(mai_mai_n920_));
  OAI220     m0892(.A0(mai_mai_n840_), .A1(mai_mai_n847_), .B0(mai_mai_n498_), .B1(mai_mai_n396_), .Y(mai_mai_n921_));
  NA3        m0893(.A(mai_mai_n921_), .B(mai_mai_n920_), .C(mai_mai_n918_), .Y(mai_mai_n922_));
  OAI210     m0894(.A0(mai_mai_n843_), .A1(mai_mai_n838_), .B0(mai_mai_n909_), .Y(mai_mai_n923_));
  AOI210     m0895(.A0(mai_mai_n349_), .A1(mai_mai_n347_), .B0(mai_mai_n296_), .Y(mai_mai_n924_));
  NA2        m0896(.A(mai_mai_n924_), .B(mai_mai_n923_), .Y(mai_mai_n925_));
  OR4        m0897(.A(mai_mai_n925_), .B(mai_mai_n922_), .C(mai_mai_n917_), .D(mai_mai_n916_), .Y(mai_mai_n926_));
  NO4        m0898(.A(mai_mai_n926_), .B(mai_mai_n915_), .C(mai_mai_n911_), .D(mai_mai_n908_), .Y(mai_mai_n927_));
  NA4        m0899(.A(mai_mai_n927_), .B(mai_mai_n901_), .C(mai_mai_n869_), .D(mai_mai_n856_), .Y(mai13));
  INV        m0900(.A(mai_mai_n44_), .Y(mai_mai_n929_));
  AN2        m0901(.A(c), .B(b), .Y(mai_mai_n930_));
  NA3        m0902(.A(mai_mai_n227_), .B(mai_mai_n930_), .C(m), .Y(mai_mai_n931_));
  NO4        m0903(.A(e), .B(mai_mai_n931_), .C(mai_mai_n929_), .D(mai_mai_n537_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n241_), .B(mai_mai_n930_), .Y(mai_mai_n933_));
  NO3        m0905(.A(mai_mai_n933_), .B(e), .C(mai_mai_n871_), .Y(mai_mai_n934_));
  NAi32      m0906(.An(d), .Bn(c), .C(e), .Y(mai_mai_n935_));
  NA2        m0907(.A(mai_mai_n130_), .B(mai_mai_n43_), .Y(mai_mai_n936_));
  NO4        m0908(.A(mai_mai_n936_), .B(mai_mai_n935_), .C(mai_mai_n542_), .D(mai_mai_n277_), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n609_), .B(mai_mai_n204_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n379_), .B(mai_mai_n192_), .Y(mai_mai_n939_));
  AN2        m0911(.A(d), .B(c), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n940_), .B(mai_mai_n107_), .Y(mai_mai_n941_));
  NO4        m0913(.A(mai_mai_n941_), .B(mai_mai_n939_), .C(mai_mai_n160_), .D(mai_mai_n152_), .Y(mai_mai_n942_));
  NA2        m0914(.A(d), .B(c), .Y(mai_mai_n943_));
  NO4        m0915(.A(mai_mai_n936_), .B(mai_mai_n539_), .C(mai_mai_n943_), .D(mai_mai_n277_), .Y(mai_mai_n944_));
  AO210      m0916(.A0(mai_mai_n942_), .A1(mai_mai_n938_), .B0(mai_mai_n944_), .Y(mai_mai_n945_));
  OR4        m0917(.A(mai_mai_n945_), .B(mai_mai_n937_), .C(mai_mai_n934_), .D(mai_mai_n932_), .Y(mai_mai_n946_));
  NO2        m0918(.A(f), .B(mai_mai_n136_), .Y(mai_mai_n947_));
  NA2        m0919(.A(mai_mai_n947_), .B(g), .Y(mai_mai_n948_));
  OR3        m0920(.A(mai_mai_n204_), .B(mai_mai_n160_), .C(mai_mai_n152_), .Y(mai_mai_n949_));
  NO2        m0921(.A(mai_mai_n949_), .B(mai_mai_n948_), .Y(mai_mai_n950_));
  NO2        m0922(.A(mai_mai_n943_), .B(mai_mai_n277_), .Y(mai_mai_n951_));
  NA2        m0923(.A(mai_mai_n579_), .B(mai_mai_n1371_), .Y(mai_mai_n952_));
  NOi21      m0924(.An(mai_mai_n951_), .B(mai_mai_n952_), .Y(mai_mai_n953_));
  NO2        m0925(.A(mai_mai_n699_), .B(mai_mai_n103_), .Y(mai_mai_n954_));
  NOi41      m0926(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n955_));
  NA2        m0927(.A(mai_mai_n955_), .B(mai_mai_n954_), .Y(mai_mai_n956_));
  NO2        m0928(.A(mai_mai_n956_), .B(mai_mai_n948_), .Y(mai_mai_n957_));
  OR3        m0929(.A(e), .B(d), .C(c), .Y(mai_mai_n958_));
  NA3        m0930(.A(k), .B(j), .C(i), .Y(mai_mai_n959_));
  NO3        m0931(.A(mai_mai_n959_), .B(mai_mai_n277_), .C(mai_mai_n82_), .Y(mai_mai_n960_));
  NOi21      m0932(.An(mai_mai_n960_), .B(mai_mai_n958_), .Y(mai_mai_n961_));
  OR4        m0933(.A(mai_mai_n961_), .B(mai_mai_n957_), .C(mai_mai_n953_), .D(mai_mai_n950_), .Y(mai_mai_n962_));
  NA3        m0934(.A(mai_mai_n432_), .B(mai_mai_n299_), .C(mai_mai_n52_), .Y(mai_mai_n963_));
  NO2        m0935(.A(mai_mai_n963_), .B(mai_mai_n952_), .Y(mai_mai_n964_));
  NO3        m0936(.A(mai_mai_n963_), .B(mai_mai_n539_), .C(mai_mai_n415_), .Y(mai_mai_n965_));
  NO2        m0937(.A(f), .B(c), .Y(mai_mai_n966_));
  NOi21      m0938(.An(mai_mai_n966_), .B(mai_mai_n409_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n967_), .B(mai_mai_n55_), .Y(mai_mai_n968_));
  NO3        m0940(.A(k), .B(mai_mai_n223_), .C(l), .Y(mai_mai_n969_));
  NOi21      m0941(.An(mai_mai_n969_), .B(mai_mai_n968_), .Y(mai_mai_n970_));
  OR3        m0942(.A(mai_mai_n970_), .B(mai_mai_n965_), .C(mai_mai_n964_), .Y(mai_mai_n971_));
  OR3        m0943(.A(mai_mai_n971_), .B(mai_mai_n962_), .C(mai_mai_n946_), .Y(mai02));
  OR2        m0944(.A(l), .B(k), .Y(mai_mai_n973_));
  OR3        m0945(.A(n), .B(m), .C(i), .Y(mai_mai_n974_));
  NO4        m0946(.A(mai_mai_n974_), .B(h), .C(mai_mai_n973_), .D(mai_mai_n958_), .Y(mai_mai_n975_));
  NOi31      m0947(.An(e), .B(d), .C(c), .Y(mai_mai_n976_));
  AOI210     m0948(.A0(mai_mai_n960_), .A1(mai_mai_n976_), .B0(mai_mai_n937_), .Y(mai_mai_n977_));
  AN3        m0949(.A(g), .B(f), .C(c), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n978_), .B(mai_mai_n432_), .Y(mai_mai_n979_));
  OR2        m0951(.A(mai_mai_n959_), .B(mai_mai_n277_), .Y(mai_mai_n980_));
  OR2        m0952(.A(mai_mai_n980_), .B(mai_mai_n979_), .Y(mai_mai_n981_));
  NO3        m0953(.A(mai_mai_n963_), .B(mai_mai_n936_), .C(mai_mai_n539_), .Y(mai_mai_n982_));
  NO2        m0954(.A(mai_mai_n982_), .B(mai_mai_n950_), .Y(mai_mai_n983_));
  NA3        m0955(.A(l), .B(k), .C(j), .Y(mai_mai_n984_));
  NA2        m0956(.A(i), .B(h), .Y(mai_mai_n985_));
  NO3        m0957(.A(mai_mai_n985_), .B(mai_mai_n984_), .C(mai_mai_n121_), .Y(mai_mai_n986_));
  NO3        m0958(.A(mai_mai_n132_), .B(mai_mai_n259_), .C(mai_mai_n193_), .Y(mai_mai_n987_));
  AOI210     m0959(.A0(mai_mai_n987_), .A1(mai_mai_n986_), .B0(mai_mai_n953_), .Y(mai_mai_n988_));
  NA3        m0960(.A(c), .B(b), .C(a), .Y(mai_mai_n989_));
  NO3        m0961(.A(mai_mai_n989_), .B(mai_mai_n816_), .C(mai_mai_n192_), .Y(mai_mai_n990_));
  NO3        m0962(.A(mai_mai_n959_), .B(mai_mai_n271_), .C(mai_mai_n45_), .Y(mai_mai_n991_));
  AOI210     m0963(.A0(mai_mai_n991_), .A1(mai_mai_n990_), .B0(mai_mai_n964_), .Y(mai_mai_n992_));
  AN4        m0964(.A(mai_mai_n992_), .B(mai_mai_n988_), .C(mai_mai_n983_), .D(mai_mai_n981_), .Y(mai_mai_n993_));
  NO2        m0965(.A(mai_mai_n941_), .B(mai_mai_n939_), .Y(mai_mai_n994_));
  NA2        m0966(.A(mai_mai_n956_), .B(mai_mai_n949_), .Y(mai_mai_n995_));
  AOI210     m0967(.A0(mai_mai_n995_), .A1(mai_mai_n994_), .B0(mai_mai_n932_), .Y(mai_mai_n996_));
  NAi41      m0968(.An(mai_mai_n975_), .B(mai_mai_n996_), .C(mai_mai_n993_), .D(mai_mai_n977_), .Y(mai03));
  NA4        m0969(.A(mai_mai_n528_), .B(m), .C(mai_mai_n103_), .D(mai_mai_n192_), .Y(mai_mai_n998_));
  NA2        m0970(.A(mai_mai_n998_), .B(mai_mai_n337_), .Y(mai_mai_n999_));
  NO2        m0971(.A(mai_mai_n999_), .B(mai_mai_n896_), .Y(mai_mai_n1000_));
  NOi21      m0972(.An(mai_mai_n730_), .B(mai_mai_n761_), .Y(mai_mai_n1001_));
  OAI220     m0973(.A0(mai_mai_n1001_), .A1(mai_mai_n631_), .B0(mai_mai_n1000_), .B1(mai_mai_n540_), .Y(mai_mai_n1002_));
  NA3        m0974(.A(mai_mai_n976_), .B(mai_mai_n308_), .C(mai_mai_n299_), .Y(mai_mai_n1003_));
  OAI210     m0975(.A0(mai_mai_n742_), .A1(mai_mai_n390_), .B0(mai_mai_n1003_), .Y(mai_mai_n1004_));
  NOi31      m0976(.An(m), .B(n), .C(f), .Y(mai_mai_n1005_));
  NA2        m0977(.A(mai_mai_n1005_), .B(mai_mai_n47_), .Y(mai_mai_n1006_));
  AN2        m0978(.A(e), .B(c), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n1007_), .B(a), .Y(mai_mai_n1008_));
  OAI220     m0980(.A0(mai_mai_n1008_), .A1(mai_mai_n1006_), .B0(mai_mai_n800_), .B1(mai_mai_n395_), .Y(mai_mai_n1009_));
  NA2        m0981(.A(mai_mai_n467_), .B(l), .Y(mai_mai_n1010_));
  NOi31      m0982(.An(mai_mai_n780_), .B(mai_mai_n931_), .C(mai_mai_n1010_), .Y(mai_mai_n1011_));
  NO4        m0983(.A(mai_mai_n1011_), .B(mai_mai_n1009_), .C(mai_mai_n1004_), .D(mai_mai_n895_), .Y(mai_mai_n1012_));
  NO2        m0984(.A(mai_mai_n259_), .B(a), .Y(mai_mai_n1013_));
  INV        m0985(.A(mai_mai_n937_), .Y(mai_mai_n1014_));
  NO2        m0986(.A(mai_mai_n985_), .B(mai_mai_n449_), .Y(mai_mai_n1015_));
  NO2        m0987(.A(mai_mai_n79_), .B(g), .Y(mai_mai_n1016_));
  AOI210     m0988(.A0(mai_mai_n1016_), .A1(mai_mai_n1015_), .B0(mai_mai_n969_), .Y(mai_mai_n1017_));
  OR2        m0989(.A(mai_mai_n1017_), .B(mai_mai_n968_), .Y(mai_mai_n1018_));
  NA3        m0990(.A(mai_mai_n1018_), .B(mai_mai_n1014_), .C(mai_mai_n1012_), .Y(mai_mai_n1019_));
  NO4        m0991(.A(mai_mai_n1019_), .B(mai_mai_n1002_), .C(mai_mai_n743_), .D(mai_mai_n517_), .Y(mai_mai_n1020_));
  NA2        m0992(.A(c), .B(b), .Y(mai_mai_n1021_));
  NO2        m0993(.A(mai_mai_n643_), .B(mai_mai_n1021_), .Y(mai_mai_n1022_));
  OAI210     m0994(.A0(mai_mai_n778_), .A1(mai_mai_n755_), .B0(mai_mai_n383_), .Y(mai_mai_n1023_));
  OAI210     m0995(.A0(mai_mai_n1023_), .A1(mai_mai_n779_), .B0(mai_mai_n1022_), .Y(mai_mai_n1024_));
  NA3        m0996(.A(mai_mai_n396_), .B(mai_mai_n510_), .C(f), .Y(mai_mai_n1025_));
  OAI210     m0997(.A0(mai_mai_n502_), .A1(mai_mai_n39_), .B0(mai_mai_n1013_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n1026_), .B(mai_mai_n1025_), .Y(mai_mai_n1027_));
  NA2        m0999(.A(mai_mai_n237_), .B(mai_mai_n110_), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n1028_), .B(g), .Y(mai_mai_n1029_));
  NAi21      m1001(.An(f), .B(d), .Y(mai_mai_n1030_));
  NO2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n989_), .Y(mai_mai_n1031_));
  INV        m1003(.A(mai_mai_n1031_), .Y(mai_mai_n1032_));
  AOI210     m1004(.A0(mai_mai_n1029_), .A1(mai_mai_n263_), .B0(mai_mai_n1032_), .Y(mai_mai_n1033_));
  AOI210     m1005(.A0(mai_mai_n1033_), .A1(mai_mai_n104_), .B0(mai_mai_n1027_), .Y(mai_mai_n1034_));
  NO2        m1006(.A(mai_mai_n165_), .B(mai_mai_n216_), .Y(mai_mai_n1035_));
  NA2        m1007(.A(mai_mai_n1035_), .B(m), .Y(mai_mai_n1036_));
  NA3        m1008(.A(mai_mai_n828_), .B(mai_mai_n1010_), .C(mai_mai_n437_), .Y(mai_mai_n1037_));
  INV        m1009(.A(mai_mai_n435_), .Y(mai_mai_n1038_));
  NO2        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n145_), .B(mai_mai_n33_), .Y(mai_mai_n1040_));
  AOI210     m1012(.A0(mai_mai_n867_), .A1(mai_mai_n1040_), .B0(mai_mai_n193_), .Y(mai_mai_n1041_));
  NA2        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1031_), .Y(mai_mai_n1042_));
  NO2        m1014(.A(mai_mai_n340_), .B(mai_mai_n339_), .Y(mai_mai_n1043_));
  AOI210     m1015(.A0(mai_mai_n1035_), .A1(mai_mai_n398_), .B0(mai_mai_n864_), .Y(mai_mai_n1044_));
  NAi31      m1016(.An(mai_mai_n1043_), .B(mai_mai_n1044_), .C(mai_mai_n1042_), .Y(mai_mai_n1045_));
  NO2        m1017(.A(mai_mai_n1045_), .B(mai_mai_n1039_), .Y(mai_mai_n1046_));
  NA4        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1034_), .C(mai_mai_n1024_), .D(mai_mai_n1020_), .Y(mai00));
  AOI210     m1019(.A0(mai_mai_n270_), .A1(mai_mai_n193_), .B0(mai_mai_n251_), .Y(mai_mai_n1048_));
  NO2        m1020(.A(mai_mai_n1048_), .B(mai_mai_n531_), .Y(mai_mai_n1049_));
  AOI210     m1021(.A0(mai_mai_n813_), .A1(mai_mai_n849_), .B0(mai_mai_n1004_), .Y(mai_mai_n1050_));
  NO2        m1022(.A(mai_mai_n982_), .B(mai_mai_n864_), .Y(mai_mai_n1051_));
  NA3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1050_), .C(mai_mai_n897_), .Y(mai_mai_n1052_));
  NA2        m1024(.A(mai_mai_n469_), .B(f), .Y(mai_mai_n1053_));
  NO2        m1025(.A(mai_mai_n903_), .B(mai_mai_n40_), .Y(mai_mai_n1054_));
  NA3        m1026(.A(mai_mai_n1054_), .B(mai_mai_n233_), .C(n), .Y(mai_mai_n1055_));
  AOI210     m1027(.A0(mai_mai_n1055_), .A1(mai_mai_n1053_), .B0(mai_mai_n941_), .Y(mai_mai_n1056_));
  NO4        m1028(.A(mai_mai_n1056_), .B(mai_mai_n1052_), .C(mai_mai_n1049_), .D(mai_mai_n962_), .Y(mai_mai_n1057_));
  NA3        m1029(.A(mai_mai_n151_), .B(mai_mai_n44_), .C(mai_mai_n43_), .Y(mai_mai_n1058_));
  NA3        m1030(.A(d), .B(mai_mai_n52_), .C(b), .Y(mai_mai_n1059_));
  NOi31      m1031(.An(n), .B(m), .C(i), .Y(mai_mai_n1060_));
  NA3        m1032(.A(mai_mai_n1060_), .B(mai_mai_n591_), .C(mai_mai_n47_), .Y(mai_mai_n1061_));
  OAI210     m1033(.A0(mai_mai_n1059_), .A1(mai_mai_n1058_), .B0(mai_mai_n1061_), .Y(mai_mai_n1062_));
  INV        m1034(.A(mai_mai_n530_), .Y(mai_mai_n1063_));
  NO3        m1035(.A(mai_mai_n1063_), .B(mai_mai_n1062_), .C(mai_mai_n1043_), .Y(mai_mai_n1064_));
  NA3        m1036(.A(mai_mai_n352_), .B(mai_mai_n200_), .C(g), .Y(mai_mai_n1065_));
  OA220      m1037(.A0(mai_mai_n1065_), .A1(mai_mai_n1059_), .B0(mai_mai_n353_), .B1(mai_mai_n124_), .Y(mai_mai_n1066_));
  NO2        m1038(.A(h), .B(g), .Y(mai_mai_n1067_));
  NA4        m1039(.A(mai_mai_n459_), .B(mai_mai_n432_), .C(mai_mai_n1067_), .D(mai_mai_n930_), .Y(mai_mai_n1068_));
  NA2        m1040(.A(mai_mai_n852_), .B(mai_mai_n529_), .Y(mai_mai_n1069_));
  NA3        m1041(.A(mai_mai_n1069_), .B(mai_mai_n1068_), .C(mai_mai_n1066_), .Y(mai_mai_n1070_));
  NO2        m1042(.A(mai_mai_n1070_), .B(mai_mai_n243_), .Y(mai_mai_n1071_));
  NO2        m1043(.A(mai_mai_n218_), .B(mai_mai_n164_), .Y(mai_mai_n1072_));
  NA2        m1044(.A(mai_mai_n1072_), .B(mai_mai_n396_), .Y(mai_mai_n1073_));
  NA3        m1045(.A(mai_mai_n163_), .B(mai_mai_n103_), .C(g), .Y(mai_mai_n1074_));
  NA3        m1046(.A(mai_mai_n432_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1075_));
  NOi31      m1047(.An(mai_mai_n786_), .B(mai_mai_n1075_), .C(mai_mai_n1074_), .Y(mai_mai_n1076_));
  NAi31      m1048(.An(mai_mai_n167_), .B(mai_mai_n775_), .C(mai_mai_n432_), .Y(mai_mai_n1077_));
  NAi31      m1049(.An(mai_mai_n1076_), .B(mai_mai_n1077_), .C(mai_mai_n1073_), .Y(mai_mai_n1078_));
  NO2        m1050(.A(mai_mai_n250_), .B(mai_mai_n67_), .Y(mai_mai_n1079_));
  NO3        m1051(.A(mai_mai_n395_), .B(mai_mai_n754_), .C(n), .Y(mai_mai_n1080_));
  AOI210     m1052(.A0(mai_mai_n1080_), .A1(mai_mai_n1079_), .B0(mai_mai_n975_), .Y(mai_mai_n1081_));
  NAi31      m1053(.An(mai_mai_n944_), .B(mai_mai_n1081_), .C(mai_mai_n66_), .Y(mai_mai_n1082_));
  NO3        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1078_), .C(mai_mai_n532_), .Y(mai_mai_n1083_));
  AN3        m1055(.A(mai_mai_n1083_), .B(mai_mai_n1071_), .C(mai_mai_n1064_), .Y(mai_mai_n1084_));
  NA3        m1056(.A(mai_mai_n1005_), .B(mai_mai_n559_), .C(mai_mai_n431_), .Y(mai_mai_n1085_));
  NA3        m1057(.A(mai_mai_n1085_), .B(mai_mai_n513_), .C(mai_mai_n221_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n999_), .B(mai_mai_n490_), .Y(mai_mai_n1087_));
  NA2        m1059(.A(mai_mai_n1087_), .B(mai_mai_n267_), .Y(mai_mai_n1088_));
  OAI210     m1060(.A0(mai_mai_n430_), .A1(mai_mai_n111_), .B0(mai_mai_n781_), .Y(mai_mai_n1089_));
  NA2        m1061(.A(mai_mai_n1089_), .B(mai_mai_n1037_), .Y(mai_mai_n1090_));
  OR3        m1062(.A(mai_mai_n941_), .B(mai_mai_n202_), .C(e), .Y(mai_mai_n1091_));
  NO2        m1063(.A(mai_mai_n196_), .B(mai_mai_n193_), .Y(mai_mai_n1092_));
  NA2        m1064(.A(n), .B(e), .Y(mai_mai_n1093_));
  NO2        m1065(.A(mai_mai_n1093_), .B(mai_mai_n136_), .Y(mai_mai_n1094_));
  AOI220     m1066(.A0(mai_mai_n1094_), .A1(mai_mai_n248_), .B0(mai_mai_n765_), .B1(mai_mai_n1092_), .Y(mai_mai_n1095_));
  OAI210     m1067(.A0(mai_mai_n323_), .A1(mai_mai_n282_), .B0(mai_mai_n414_), .Y(mai_mai_n1096_));
  NA4        m1068(.A(mai_mai_n1096_), .B(mai_mai_n1095_), .C(mai_mai_n1091_), .D(mai_mai_n1090_), .Y(mai_mai_n1097_));
  AOI210     m1069(.A0(mai_mai_n1094_), .A1(mai_mai_n769_), .B0(mai_mai_n743_), .Y(mai_mai_n1098_));
  AOI220     m1070(.A0(mai_mai_n860_), .A1(mai_mai_n529_), .B0(mai_mai_n591_), .B1(mai_mai_n224_), .Y(mai_mai_n1099_));
  NO2        m1071(.A(mai_mai_n61_), .B(h), .Y(mai_mai_n1100_));
  NO3        m1072(.A(mai_mai_n941_), .B(mai_mai_n939_), .C(mai_mai_n664_), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n973_), .B(mai_mai_n121_), .Y(mai_mai_n1102_));
  AN2        m1074(.A(mai_mai_n1102_), .B(mai_mai_n987_), .Y(mai_mai_n1103_));
  OAI210     m1075(.A0(mai_mai_n1103_), .A1(mai_mai_n1101_), .B0(mai_mai_n1100_), .Y(mai_mai_n1104_));
  NA4        m1076(.A(mai_mai_n1104_), .B(mai_mai_n1099_), .C(mai_mai_n1098_), .D(mai_mai_n782_), .Y(mai_mai_n1105_));
  NO4        m1077(.A(mai_mai_n1105_), .B(mai_mai_n1097_), .C(mai_mai_n1088_), .D(mai_mai_n1086_), .Y(mai_mai_n1106_));
  NA2        m1078(.A(mai_mai_n756_), .B(mai_mai_n694_), .Y(mai_mai_n1107_));
  NA4        m1079(.A(mai_mai_n1107_), .B(mai_mai_n1106_), .C(mai_mai_n1084_), .D(mai_mai_n1057_), .Y(mai01));
  AN2        m1080(.A(mai_mai_n920_), .B(mai_mai_n918_), .Y(mai_mai_n1109_));
  NO4        m1081(.A(mai_mai_n726_), .B(mai_mai_n720_), .C(mai_mai_n444_), .D(mai_mai_n257_), .Y(mai_mai_n1110_));
  NA2        m1082(.A(mai_mai_n363_), .B(i), .Y(mai_mai_n1111_));
  NA3        m1083(.A(mai_mai_n1111_), .B(mai_mai_n1110_), .C(mai_mai_n1109_), .Y(mai_mai_n1112_));
  NA2        m1084(.A(mai_mai_n826_), .B(mai_mai_n298_), .Y(mai_mai_n1113_));
  NA2        m1085(.A(mai_mai_n650_), .B(mai_mai_n88_), .Y(mai_mai_n1114_));
  NO2        m1086(.A(mai_mai_n1114_), .B(mai_mai_n1367_), .Y(mai_mai_n1115_));
  INV        m1087(.A(mai_mai_n109_), .Y(mai_mai_n1116_));
  OR2        m1088(.A(mai_mai_n603_), .B(mai_mai_n337_), .Y(mai_mai_n1117_));
  NA2        m1089(.A(mai_mai_n1117_), .B(mai_mai_n812_), .Y(mai_mai_n1118_));
  NO3        m1090(.A(mai_mai_n711_), .B(mai_mai_n615_), .C(mai_mai_n471_), .Y(mai_mai_n1119_));
  NA2        m1091(.A(mai_mai_n1119_), .B(mai_mai_n127_), .Y(mai_mai_n1120_));
  NO4        m1092(.A(mai_mai_n1120_), .B(mai_mai_n1118_), .C(mai_mai_n1113_), .D(mai_mai_n1112_), .Y(mai_mai_n1121_));
  INV        m1093(.A(mai_mai_n1065_), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n1122_), .B(mai_mai_n486_), .Y(mai_mai_n1123_));
  NA2        m1095(.A(mai_mai_n492_), .B(mai_mai_n365_), .Y(mai_mai_n1124_));
  NOi21      m1096(.An(mai_mai_n514_), .B(mai_mai_n536_), .Y(mai_mai_n1125_));
  NA2        m1097(.A(mai_mai_n1125_), .B(mai_mai_n1124_), .Y(mai_mai_n1126_));
  AOI210     m1098(.A0(mai_mai_n183_), .A1(mai_mai_n81_), .B0(mai_mai_n192_), .Y(mai_mai_n1127_));
  OAI210     m1099(.A0(mai_mai_n733_), .A1(mai_mai_n396_), .B0(mai_mai_n1127_), .Y(mai_mai_n1128_));
  AN3        m1100(.A(m), .B(l), .C(k), .Y(mai_mai_n1129_));
  OAI210     m1101(.A0(mai_mai_n325_), .A1(mai_mai_n34_), .B0(mai_mai_n1129_), .Y(mai_mai_n1130_));
  NA2        m1102(.A(mai_mai_n182_), .B(mai_mai_n34_), .Y(mai_mai_n1131_));
  AO210      m1103(.A0(mai_mai_n1131_), .A1(mai_mai_n1130_), .B0(mai_mai_n297_), .Y(mai_mai_n1132_));
  NA4        m1104(.A(mai_mai_n1132_), .B(mai_mai_n1128_), .C(mai_mai_n1126_), .D(mai_mai_n1123_), .Y(mai_mai_n1133_));
  AOI210     m1105(.A0(mai_mai_n548_), .A1(mai_mai_n109_), .B0(mai_mai_n554_), .Y(mai_mai_n1134_));
  OAI210     m1106(.A0(mai_mai_n1116_), .A1(mai_mai_n545_), .B0(mai_mai_n1134_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n256_), .B(mai_mai_n177_), .Y(mai_mai_n1136_));
  NA2        m1108(.A(mai_mai_n1136_), .B(mai_mai_n608_), .Y(mai_mai_n1137_));
  NO3        m1109(.A(mai_mai_n742_), .B(mai_mai_n183_), .C(mai_mai_n377_), .Y(mai_mai_n1138_));
  NO2        m1110(.A(mai_mai_n1138_), .B(mai_mai_n864_), .Y(mai_mai_n1139_));
  OAI210     m1111(.A0(mai_mai_n1115_), .A1(mai_mai_n291_), .B0(mai_mai_n616_), .Y(mai_mai_n1140_));
  NA3        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1139_), .C(mai_mai_n1137_), .Y(mai_mai_n1141_));
  NO3        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1135_), .C(mai_mai_n1133_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n465_), .B(mai_mai_n54_), .Y(mai_mai_n1143_));
  OR3        m1115(.A(mai_mai_n1114_), .B(mai_mai_n558_), .C(mai_mai_n1367_), .Y(mai_mai_n1144_));
  NO2        m1116(.A(mai_mai_n186_), .B(mai_mai_n102_), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n1145_), .B(mai_mai_n1062_), .Y(mai_mai_n1146_));
  NA4        m1118(.A(mai_mai_n1146_), .B(mai_mai_n1144_), .C(mai_mai_n1143_), .D(mai_mai_n693_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n871_), .B(mai_mai_n212_), .Y(mai_mai_n1148_));
  NO2        m1120(.A(mai_mai_n872_), .B(mai_mai_n508_), .Y(mai_mai_n1149_));
  OAI210     m1121(.A0(mai_mai_n1149_), .A1(mai_mai_n1148_), .B0(mai_mai_n306_), .Y(mai_mai_n1150_));
  NA2        m1122(.A(mai_mai_n524_), .B(mai_mai_n522_), .Y(mai_mai_n1151_));
  INV        m1123(.A(mai_mai_n1151_), .Y(mai_mai_n1152_));
  OR2        m1124(.A(mai_mai_n1065_), .B(mai_mai_n1059_), .Y(mai_mai_n1153_));
  NO2        m1125(.A(mai_mai_n337_), .B(mai_mai_n65_), .Y(mai_mai_n1154_));
  INV        m1126(.A(mai_mai_n1154_), .Y(mai_mai_n1155_));
  NA3        m1127(.A(mai_mai_n1155_), .B(mai_mai_n1153_), .C(mai_mai_n355_), .Y(mai_mai_n1156_));
  NOi41      m1128(.An(mai_mai_n1150_), .B(mai_mai_n1156_), .C(mai_mai_n1152_), .D(mai_mai_n1147_), .Y(mai_mai_n1157_));
  NO2        m1129(.A(mai_mai_n120_), .B(mai_mai_n43_), .Y(mai_mai_n1158_));
  AO220      m1130(.A0(i), .A1(mai_mai_n573_), .B0(mai_mai_n1158_), .B1(mai_mai_n648_), .Y(mai_mai_n1159_));
  NA2        m1131(.A(mai_mai_n1159_), .B(mai_mai_n306_), .Y(mai_mai_n1160_));
  NO3        m1132(.A(mai_mai_n985_), .B(mai_mai_n160_), .C(mai_mai_n79_), .Y(mai_mai_n1161_));
  INV        m1133(.A(mai_mai_n1160_), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n567_), .B(mai_mai_n566_), .Y(mai_mai_n1163_));
  NO4        m1135(.A(mai_mai_n985_), .B(mai_mai_n1163_), .C(mai_mai_n158_), .D(mai_mai_n79_), .Y(mai_mai_n1164_));
  NO3        m1136(.A(mai_mai_n1164_), .B(mai_mai_n1162_), .C(mai_mai_n585_), .Y(mai_mai_n1165_));
  NA4        m1137(.A(mai_mai_n1165_), .B(mai_mai_n1157_), .C(mai_mai_n1142_), .D(mai_mai_n1121_), .Y(mai06));
  NO2        m1138(.A(mai_mai_n378_), .B(mai_mai_n511_), .Y(mai_mai_n1167_));
  INV        m1139(.A(mai_mai_n671_), .Y(mai_mai_n1168_));
  NA2        m1140(.A(mai_mai_n1168_), .B(mai_mai_n1167_), .Y(mai_mai_n1169_));
  NO2        m1141(.A(mai_mai_n204_), .B(mai_mai_n93_), .Y(mai_mai_n1170_));
  OAI210     m1142(.A0(mai_mai_n1170_), .A1(mai_mai_n1161_), .B0(mai_mai_n351_), .Y(mai_mai_n1171_));
  NO3        m1143(.A(mai_mai_n552_), .B(mai_mai_n731_), .C(mai_mai_n555_), .Y(mai_mai_n1172_));
  OR2        m1144(.A(mai_mai_n1172_), .B(mai_mai_n800_), .Y(mai_mai_n1173_));
  NA4        m1145(.A(mai_mai_n1173_), .B(mai_mai_n1171_), .C(mai_mai_n1169_), .D(mai_mai_n1150_), .Y(mai_mai_n1174_));
  NO3        m1146(.A(mai_mai_n1174_), .B(mai_mai_n1152_), .C(mai_mai_n232_), .Y(mai_mai_n1175_));
  AOI210     m1147(.A0(i), .A1(mai_mai_n875_), .B0(mai_mai_n1148_), .Y(mai_mai_n1176_));
  INV        m1148(.A(mai_mai_n1159_), .Y(mai_mai_n1177_));
  AOI210     m1149(.A0(mai_mai_n1177_), .A1(mai_mai_n1176_), .B0(mai_mai_n303_), .Y(mai_mai_n1178_));
  OAI210     m1150(.A0(mai_mai_n81_), .A1(mai_mai_n40_), .B0(mai_mai_n614_), .Y(mai_mai_n1179_));
  NA2        m1151(.A(mai_mai_n1179_), .B(mai_mai_n587_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n474_), .B(mai_mai_n155_), .Y(mai_mai_n1181_));
  NO2        m1153(.A(mai_mai_n560_), .B(mai_mai_n1006_), .Y(mai_mai_n1182_));
  OAI210     m1154(.A0(mai_mai_n425_), .A1(mai_mai_n226_), .B0(mai_mai_n820_), .Y(mai_mai_n1183_));
  NO4        m1155(.A(mai_mai_n1183_), .B(mai_mai_n1182_), .C(mai_mai_n126_), .D(mai_mai_n1181_), .Y(mai_mai_n1184_));
  OR2        m1156(.A(mai_mai_n553_), .B(mai_mai_n551_), .Y(mai_mai_n1185_));
  NO2        m1157(.A(mai_mai_n336_), .B(mai_mai_n125_), .Y(mai_mai_n1186_));
  AOI210     m1158(.A0(mai_mai_n1186_), .A1(mai_mai_n541_), .B0(mai_mai_n1185_), .Y(mai_mai_n1187_));
  NA3        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1184_), .C(mai_mai_n1180_), .Y(mai_mai_n1188_));
  NO2        m1160(.A(mai_mai_n686_), .B(mai_mai_n335_), .Y(mai_mai_n1189_));
  NO2        m1161(.A(mai_mai_n616_), .B(mai_mai_n695_), .Y(mai_mai_n1190_));
  NOi21      m1162(.An(mai_mai_n1189_), .B(mai_mai_n1190_), .Y(mai_mai_n1191_));
  NO3        m1163(.A(mai_mai_n1191_), .B(mai_mai_n1188_), .C(mai_mai_n1178_), .Y(mai_mai_n1192_));
  OAI220     m1164(.A0(mai_mai_n671_), .A1(mai_mai_n1370_), .B0(mai_mai_n204_), .B1(mai_mai_n568_), .Y(mai_mai_n1193_));
  OAI210     m1165(.A0(mai_mai_n252_), .A1(c), .B0(mai_mai_n586_), .Y(mai_mai_n1194_));
  NA2        m1166(.A(mai_mai_n1194_), .B(mai_mai_n1193_), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n640_), .B(mai_mai_n226_), .Y(mai_mai_n1196_));
  NO2        m1168(.A(mai_mai_n1196_), .B(mai_mai_n1009_), .Y(mai_mai_n1197_));
  NA4        m1169(.A(mai_mai_n718_), .B(mai_mai_n717_), .C(mai_mai_n406_), .D(mai_mai_n793_), .Y(mai_mai_n1198_));
  NAi31      m1170(.An(mai_mai_n686_), .B(mai_mai_n1198_), .C(mai_mai_n182_), .Y(mai_mai_n1199_));
  NA4        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1197_), .C(mai_mai_n1195_), .D(mai_mai_n1099_), .Y(mai_mai_n1200_));
  NO2        m1172(.A(mai_mai_n429_), .B(mai_mai_n364_), .Y(mai_mai_n1201_));
  OR3        m1173(.A(mai_mai_n1201_), .B(mai_mai_n710_), .C(mai_mai_n494_), .Y(mai_mai_n1202_));
  OR3        m1174(.A(mai_mai_n339_), .B(mai_mai_n204_), .C(mai_mai_n568_), .Y(mai_mai_n1203_));
  AOI210     m1175(.A0(mai_mai_n524_), .A1(mai_mai_n414_), .B0(mai_mai_n341_), .Y(mai_mai_n1204_));
  NA3        m1176(.A(mai_mai_n1204_), .B(mai_mai_n1203_), .C(mai_mai_n1202_), .Y(mai_mai_n1205_));
  AOI220     m1177(.A0(mai_mai_n1189_), .A1(mai_mai_n694_), .B0(mai_mai_n1186_), .B1(mai_mai_n217_), .Y(mai_mai_n1206_));
  AN2        m1178(.A(mai_mai_n838_), .B(mai_mai_n837_), .Y(mai_mai_n1207_));
  NO4        m1179(.A(mai_mai_n1207_), .B(mai_mai_n791_), .C(mai_mai_n461_), .D(mai_mai_n447_), .Y(mai_mai_n1208_));
  NA2        m1180(.A(mai_mai_n1208_), .B(mai_mai_n1206_), .Y(mai_mai_n1209_));
  NO3        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1205_), .C(mai_mai_n1200_), .Y(mai_mai_n1210_));
  NA4        m1182(.A(mai_mai_n1210_), .B(mai_mai_n1192_), .C(mai_mai_n1175_), .D(mai_mai_n1165_), .Y(mai07));
  NOi21      m1183(.An(j), .B(k), .Y(mai_mai_n1212_));
  NA4        m1184(.A(mai_mai_n163_), .B(mai_mai_n99_), .C(mai_mai_n1212_), .D(f), .Y(mai_mai_n1213_));
  NAi21      m1185(.An(f), .B(c), .Y(mai_mai_n1214_));
  OR2        m1186(.A(e), .B(d), .Y(mai_mai_n1215_));
  OAI220     m1187(.A0(mai_mai_n1215_), .A1(mai_mai_n1214_), .B0(mai_mai_n578_), .B1(mai_mai_n289_), .Y(mai_mai_n1216_));
  NA3        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1371_), .C(mai_mai_n163_), .Y(mai_mai_n1217_));
  NOi31      m1189(.An(n), .B(m), .C(b), .Y(mai_mai_n1218_));
  NA2        m1190(.A(mai_mai_n1217_), .B(mai_mai_n1213_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(k), .B(i), .Y(mai_mai_n1220_));
  NA2        m1192(.A(mai_mai_n79_), .B(mai_mai_n43_), .Y(mai_mai_n1221_));
  NO2        m1193(.A(mai_mai_n959_), .B(mai_mai_n277_), .Y(mai_mai_n1222_));
  NA2        m1194(.A(mai_mai_n495_), .B(mai_mai_n74_), .Y(mai_mai_n1223_));
  NA2        m1195(.A(mai_mai_n1100_), .B(mai_mai_n261_), .Y(mai_mai_n1224_));
  NA2        m1196(.A(mai_mai_n1224_), .B(mai_mai_n1223_), .Y(mai_mai_n1225_));
  NO2        m1197(.A(mai_mai_n1225_), .B(mai_mai_n1219_), .Y(mai_mai_n1226_));
  NO3        m1198(.A(e), .B(d), .C(c), .Y(mai_mai_n1227_));
  NA2        m1199(.A(mai_mai_n1366_), .B(mai_mai_n1227_), .Y(mai_mai_n1228_));
  NO2        m1200(.A(mai_mai_n1228_), .B(mai_mai_n193_), .Y(mai_mai_n1229_));
  NA3        m1201(.A(mai_mai_n637_), .B(mai_mai_n1372_), .C(mai_mai_n103_), .Y(mai_mai_n1230_));
  NO2        m1202(.A(mai_mai_n1230_), .B(mai_mai_n43_), .Y(mai_mai_n1231_));
  NO2        m1203(.A(l), .B(k), .Y(mai_mai_n1232_));
  NOi41      m1204(.An(mai_mai_n500_), .B(mai_mai_n1232_), .C(mai_mai_n442_), .D(mai_mai_n409_), .Y(mai_mai_n1233_));
  NO3        m1205(.A(mai_mai_n409_), .B(d), .C(c), .Y(mai_mai_n1234_));
  NO3        m1206(.A(mai_mai_n1233_), .B(mai_mai_n1231_), .C(mai_mai_n1229_), .Y(mai_mai_n1235_));
  NO2        m1207(.A(k), .B(l), .Y(mai_mai_n1236_));
  NO2        m1208(.A(g), .B(c), .Y(mai_mai_n1237_));
  NA3        m1209(.A(mai_mai_n1237_), .B(mai_mai_n132_), .C(mai_mai_n168_), .Y(mai_mai_n1238_));
  NO2        m1210(.A(mai_mai_n1238_), .B(mai_mai_n1236_), .Y(mai_mai_n1239_));
  NA2        m1211(.A(mai_mai_n1239_), .B(mai_mai_n163_), .Y(mai_mai_n1240_));
  NO2        m1212(.A(mai_mai_n416_), .B(a), .Y(mai_mai_n1241_));
  NA3        m1213(.A(mai_mai_n1241_), .B(mai_mai_n1369_), .C(mai_mai_n104_), .Y(mai_mai_n1242_));
  NO2        m1214(.A(i), .B(h), .Y(mai_mai_n1243_));
  NA2        m1215(.A(mai_mai_n1030_), .B(h), .Y(mai_mai_n1244_));
  NA2        m1216(.A(mai_mai_n128_), .B(mai_mai_n200_), .Y(mai_mai_n1245_));
  NO2        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1244_), .Y(mai_mai_n1246_));
  NO2        m1218(.A(mai_mai_n691_), .B(mai_mai_n169_), .Y(mai_mai_n1247_));
  NOi31      m1219(.An(m), .B(n), .C(b), .Y(mai_mai_n1248_));
  NO2        m1220(.A(mai_mai_n1247_), .B(mai_mai_n1246_), .Y(mai_mai_n1249_));
  NA2        m1221(.A(mai_mai_n978_), .B(mai_mai_n432_), .Y(mai_mai_n1250_));
  NO4        m1222(.A(mai_mai_n1250_), .B(mai_mai_n954_), .C(mai_mai_n409_), .D(mai_mai_n43_), .Y(mai_mai_n1251_));
  OAI210     m1223(.A0(mai_mai_n165_), .A1(mai_mai_n482_), .B0(mai_mai_n955_), .Y(mai_mai_n1252_));
  NO3        m1224(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1253_));
  INV        m1225(.A(mai_mai_n1252_), .Y(mai_mai_n1254_));
  NO2        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1251_), .Y(mai_mai_n1255_));
  AN4        m1227(.A(mai_mai_n1255_), .B(mai_mai_n1249_), .C(mai_mai_n1242_), .D(mai_mai_n1240_), .Y(mai_mai_n1256_));
  NA2        m1228(.A(mai_mai_n1218_), .B(mai_mai_n348_), .Y(mai_mai_n1257_));
  NO2        m1229(.A(mai_mai_n1257_), .B(mai_mai_n938_), .Y(mai_mai_n1258_));
  NA2        m1230(.A(mai_mai_n1234_), .B(mai_mai_n194_), .Y(mai_mai_n1259_));
  NO2        m1231(.A(mai_mai_n169_), .B(b), .Y(mai_mai_n1260_));
  AOI220     m1232(.A0(mai_mai_n1060_), .A1(mai_mai_n1260_), .B0(mai_mai_n986_), .B1(mai_mai_n1250_), .Y(mai_mai_n1261_));
  NAi31      m1233(.An(mai_mai_n1258_), .B(mai_mai_n1261_), .C(mai_mai_n1259_), .Y(mai_mai_n1262_));
  NO4        m1234(.A(mai_mai_n121_), .B(g), .C(f), .D(e), .Y(mai_mai_n1263_));
  NA2        m1235(.A(mai_mai_n1220_), .B(mai_mai_n262_), .Y(mai_mai_n1264_));
  OR2        m1236(.A(e), .B(a), .Y(mai_mai_n1265_));
  NOi41      m1237(.An(h), .B(f), .C(e), .D(a), .Y(mai_mai_n1266_));
  NA2        m1238(.A(mai_mai_n1266_), .B(mai_mai_n104_), .Y(mai_mai_n1267_));
  INV        m1239(.A(mai_mai_n1267_), .Y(mai_mai_n1268_));
  OR3        m1240(.A(mai_mai_n494_), .B(mai_mai_n493_), .C(mai_mai_n103_), .Y(mai_mai_n1269_));
  NA2        m1241(.A(mai_mai_n1005_), .B(mai_mai_n377_), .Y(mai_mai_n1270_));
  NO2        m1242(.A(mai_mai_n1270_), .B(mai_mai_n405_), .Y(mai_mai_n1271_));
  AO210      m1243(.A0(mai_mai_n1271_), .A1(mai_mai_n107_), .B0(mai_mai_n1268_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n1272_), .B(mai_mai_n1262_), .Y(mai_mai_n1273_));
  NA4        m1245(.A(mai_mai_n1273_), .B(mai_mai_n1256_), .C(mai_mai_n1235_), .D(mai_mai_n1226_), .Y(mai_mai_n1274_));
  NO2        m1246(.A(mai_mai_n1021_), .B(mai_mai_n101_), .Y(mai_mai_n1275_));
  NA3        m1247(.A(mai_mai_n1253_), .B(mai_mai_n1215_), .C(mai_mai_n1005_), .Y(mai_mai_n1276_));
  NAi31      m1248(.An(mai_mai_n1243_), .B(mai_mai_n967_), .C(mai_mai_n152_), .Y(mai_mai_n1277_));
  NA2        m1249(.A(mai_mai_n1277_), .B(mai_mai_n1276_), .Y(mai_mai_n1278_));
  NO3        m1250(.A(mai_mai_n686_), .B(mai_mai_n158_), .C(mai_mai_n379_), .Y(mai_mai_n1279_));
  NO2        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1278_), .Y(mai_mai_n1280_));
  OR2        m1252(.A(n), .B(i), .Y(mai_mai_n1281_));
  OAI210     m1253(.A0(mai_mai_n1281_), .A1(mai_mai_n966_), .B0(mai_mai_n45_), .Y(mai_mai_n1282_));
  AOI220     m1254(.A0(mai_mai_n1282_), .A1(mai_mai_n1067_), .B0(mai_mai_n746_), .B1(mai_mai_n176_), .Y(mai_mai_n1283_));
  INV        m1255(.A(mai_mai_n1283_), .Y(mai_mai_n1284_));
  OAI220     m1256(.A0(mai_mai_n609_), .A1(g), .B0(mai_mai_n204_), .B1(c), .Y(mai_mai_n1285_));
  AOI210     m1257(.A0(mai_mai_n1260_), .A1(mai_mai_n41_), .B0(mai_mai_n1285_), .Y(mai_mai_n1286_));
  NO2        m1258(.A(mai_mai_n121_), .B(l), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n204_), .B(k), .Y(mai_mai_n1288_));
  OAI210     m1260(.A0(mai_mai_n1288_), .A1(mai_mai_n1243_), .B0(mai_mai_n1287_), .Y(mai_mai_n1289_));
  OAI220     m1261(.A0(mai_mai_n1289_), .A1(mai_mai_n31_), .B0(mai_mai_n1286_), .B1(mai_mai_n160_), .Y(mai_mai_n1290_));
  NO3        m1262(.A(mai_mai_n1269_), .B(mai_mai_n432_), .C(mai_mai_n319_), .Y(mai_mai_n1291_));
  NO3        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1290_), .C(mai_mai_n1284_), .Y(mai_mai_n1292_));
  NO3        m1264(.A(mai_mai_n989_), .B(mai_mai_n1215_), .C(mai_mai_n45_), .Y(mai_mai_n1293_));
  NO2        m1265(.A(mai_mai_n974_), .B(h), .Y(mai_mai_n1294_));
  NA3        m1266(.A(mai_mai_n1294_), .B(d), .C(mai_mai_n939_), .Y(mai_mai_n1295_));
  NO2        m1267(.A(mai_mai_n1295_), .B(c), .Y(mai_mai_n1296_));
  NA3        m1268(.A(mai_mai_n1275_), .B(mai_mai_n432_), .C(f), .Y(mai_mai_n1297_));
  NA2        m1269(.A(mai_mai_n163_), .B(mai_mai_n103_), .Y(mai_mai_n1298_));
  NO2        m1270(.A(mai_mai_n1212_), .B(mai_mai_n42_), .Y(mai_mai_n1299_));
  AOI210     m1271(.A0(mai_mai_n104_), .A1(mai_mai_n40_), .B0(mai_mai_n1299_), .Y(mai_mai_n1300_));
  NO2        m1272(.A(mai_mai_n1300_), .B(mai_mai_n1297_), .Y(mai_mai_n1301_));
  NO2        m1273(.A(mai_mai_n1215_), .B(f), .Y(mai_mai_n1302_));
  NA2        m1274(.A(mai_mai_n1241_), .B(mai_mai_n1299_), .Y(mai_mai_n1303_));
  INV        m1275(.A(mai_mai_n1303_), .Y(mai_mai_n1304_));
  NO3        m1276(.A(mai_mai_n1304_), .B(mai_mai_n1301_), .C(mai_mai_n1296_), .Y(mai_mai_n1305_));
  NA3        m1277(.A(mai_mai_n1305_), .B(mai_mai_n1292_), .C(mai_mai_n1280_), .Y(mai_mai_n1306_));
  NO3        m1278(.A(mai_mai_n978_), .B(mai_mai_n966_), .C(mai_mai_n40_), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n432_), .B(mai_mai_n271_), .Y(mai_mai_n1308_));
  OAI210     m1280(.A0(mai_mai_n1308_), .A1(mai_mai_n1307_), .B0(mai_mai_n1222_), .Y(mai_mai_n1309_));
  OAI210     m1281(.A0(mai_mai_n1263_), .A1(mai_mai_n1218_), .B0(mai_mai_n797_), .Y(mai_mai_n1310_));
  NO2        m1282(.A(mai_mai_n935_), .B(mai_mai_n121_), .Y(mai_mai_n1311_));
  NA2        m1283(.A(mai_mai_n1311_), .B(mai_mai_n572_), .Y(mai_mai_n1312_));
  NA3        m1284(.A(mai_mai_n1312_), .B(mai_mai_n1310_), .C(mai_mai_n1309_), .Y(mai_mai_n1313_));
  NO2        m1285(.A(mai_mai_n139_), .B(mai_mai_n164_), .Y(mai_mai_n1314_));
  OAI210     m1286(.A0(mai_mai_n1314_), .A1(mai_mai_n101_), .B0(mai_mai_n1248_), .Y(mai_mai_n1315_));
  INV        m1287(.A(mai_mai_n1315_), .Y(mai_mai_n1316_));
  NO2        m1288(.A(mai_mai_n1316_), .B(mai_mai_n1313_), .Y(mai_mai_n1317_));
  NO2        m1289(.A(mai_mai_n1214_), .B(e), .Y(mai_mai_n1318_));
  INV        m1290(.A(mai_mai_n1318_), .Y(mai_mai_n1319_));
  NA2        m1291(.A(mai_mai_n1016_), .B(mai_mai_n580_), .Y(mai_mai_n1320_));
  OR3        m1292(.A(mai_mai_n1288_), .B(mai_mai_n1100_), .C(mai_mai_n121_), .Y(mai_mai_n1321_));
  OAI220     m1293(.A0(mai_mai_n1321_), .A1(mai_mai_n1319_), .B0(mai_mai_n1320_), .B1(mai_mai_n410_), .Y(mai_mai_n1322_));
  INV        m1294(.A(mai_mai_n1322_), .Y(mai_mai_n1323_));
  INV        m1295(.A(g), .Y(mai_mai_n1324_));
  AOI210     m1296(.A0(mai_mai_n1324_), .A1(mai_mai_n1234_), .B0(mai_mai_n1293_), .Y(mai_mai_n1325_));
  NO2        m1297(.A(mai_mai_n1265_), .B(f), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n1325_), .B(mai_mai_n192_), .Y(mai_mai_n1327_));
  NA2        m1299(.A(mai_mai_n1326_), .B(mai_mai_n1221_), .Y(mai_mai_n1328_));
  OAI220     m1300(.A0(mai_mai_n1328_), .A1(mai_mai_n45_), .B0(mai_mai_n1368_), .B1(mai_mai_n158_), .Y(mai_mai_n1329_));
  NA4        m1301(.A(mai_mai_n987_), .B(mai_mai_n984_), .C(mai_mai_n200_), .D(mai_mai_n61_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n45_), .B(l), .Y(mai_mai_n1331_));
  INV        m1303(.A(mai_mai_n448_), .Y(mai_mai_n1332_));
  OAI210     m1304(.A0(mai_mai_n1332_), .A1(mai_mai_n990_), .B0(mai_mai_n1331_), .Y(mai_mai_n1333_));
  NA2        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1330_), .Y(mai_mai_n1334_));
  NO3        m1306(.A(mai_mai_n1334_), .B(mai_mai_n1329_), .C(mai_mai_n1327_), .Y(mai_mai_n1335_));
  NA3        m1307(.A(mai_mai_n1335_), .B(mai_mai_n1323_), .C(mai_mai_n1317_), .Y(mai_mai_n1336_));
  NA2        m1308(.A(mai_mai_n866_), .B(mai_mai_n128_), .Y(mai_mai_n1337_));
  AOI210     m1309(.A0(f), .A1(c), .B0(mai_mai_n1337_), .Y(mai_mai_n1338_));
  INV        m1310(.A(mai_mai_n166_), .Y(mai_mai_n1339_));
  NA2        m1311(.A(mai_mai_n1339_), .B(mai_mai_n1294_), .Y(mai_mai_n1340_));
  INV        m1312(.A(mai_mai_n1340_), .Y(mai_mai_n1341_));
  NO2        m1313(.A(mai_mai_n1341_), .B(mai_mai_n1338_), .Y(mai_mai_n1342_));
  AOI210     m1314(.A0(mai_mai_n143_), .A1(mai_mai_n52_), .B0(mai_mai_n1318_), .Y(mai_mai_n1343_));
  NO2        m1315(.A(mai_mai_n1343_), .B(mai_mai_n1298_), .Y(mai_mai_n1344_));
  INV        m1316(.A(mai_mai_n1344_), .Y(mai_mai_n1345_));
  AN2        m1317(.A(mai_mai_n987_), .B(mai_mai_n973_), .Y(mai_mai_n1346_));
  NA2        m1318(.A(mai_mai_n1346_), .B(mai_mai_n1060_), .Y(mai_mai_n1347_));
  NO2        m1319(.A(mai_mai_n1297_), .B(mai_mai_n62_), .Y(mai_mai_n1348_));
  NA2        m1320(.A(mai_mai_n55_), .B(a), .Y(mai_mai_n1349_));
  NO2        m1321(.A(mai_mai_n1220_), .B(mai_mai_n109_), .Y(mai_mai_n1350_));
  OAI220     m1322(.A0(mai_mai_n1350_), .A1(mai_mai_n1257_), .B0(mai_mai_n1270_), .B1(mai_mai_n1349_), .Y(mai_mai_n1351_));
  NO2        m1323(.A(mai_mai_n1351_), .B(mai_mai_n1348_), .Y(mai_mai_n1352_));
  NA4        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1347_), .C(mai_mai_n1345_), .D(mai_mai_n1342_), .Y(mai_mai_n1353_));
  OR4        m1325(.A(mai_mai_n1353_), .B(mai_mai_n1336_), .C(mai_mai_n1306_), .D(mai_mai_n1274_), .Y(mai04));
  NOi31      m1326(.An(mai_mai_n1263_), .B(mai_mai_n1264_), .C(mai_mai_n941_), .Y(mai_mai_n1355_));
  NA2        m1327(.A(mai_mai_n1302_), .B(mai_mai_n746_), .Y(mai_mai_n1356_));
  NO2        m1328(.A(mai_mai_n1356_), .B(mai_mai_n931_), .Y(mai_mai_n1357_));
  OR3        m1329(.A(mai_mai_n1357_), .B(mai_mai_n1355_), .C(mai_mai_n957_), .Y(mai_mai_n1358_));
  NO2        m1330(.A(mai_mai_n1221_), .B(mai_mai_n82_), .Y(mai_mai_n1359_));
  AOI210     m1331(.A0(mai_mai_n1359_), .A1(mai_mai_n951_), .B0(mai_mai_n1076_), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n1360_), .B(mai_mai_n1104_), .Y(mai_mai_n1361_));
  NO4        m1333(.A(mai_mai_n1361_), .B(mai_mai_n1358_), .C(mai_mai_n965_), .D(mai_mai_n946_), .Y(mai_mai_n1362_));
  NA4        m1334(.A(mai_mai_n1362_), .B(mai_mai_n1018_), .C(mai_mai_n1003_), .D(mai_mai_n993_), .Y(mai05));
  INV        m1335(.A(m), .Y(mai_mai_n1366_));
  INV        m1336(.A(f), .Y(mai_mai_n1367_));
  INV        m1337(.A(mai_mai_n95_), .Y(mai_mai_n1368_));
  INV        m1338(.A(i), .Y(mai_mai_n1369_));
  INV        m1339(.A(h), .Y(mai_mai_n1370_));
  INV        m1340(.A(j), .Y(mai_mai_n1371_));
  INV        m1341(.A(m), .Y(mai_mai_n1372_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n44_), .B(men_men_n32_), .Y(men_men_n52_));
  INV        u0024(.A(c), .Y(men_men_n53_));
  NA2        u0025(.A(e), .B(b), .Y(men_men_n54_));
  NO2        u0026(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  INV        u0027(.A(d), .Y(men_men_n56_));
  NAi21      u0028(.An(i), .B(h), .Y(men_men_n57_));
  NAi31      u0029(.An(i), .B(l), .C(j), .Y(men_men_n58_));
  NO2        u0030(.A(men_men_n57_), .B(men_men_n44_), .Y(men_men_n59_));
  NAi31      u0031(.An(d), .B(men_men_n59_), .C(men_men_n55_), .Y(men_men_n60_));
  NAi41      u0032(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n61_));
  NA2        u0033(.A(g), .B(f), .Y(men_men_n62_));
  NO2        u0034(.A(men_men_n62_), .B(men_men_n61_), .Y(men_men_n63_));
  NAi21      u0035(.An(i), .B(j), .Y(men_men_n64_));
  NAi32      u0036(.An(n), .Bn(k), .C(m), .Y(men_men_n65_));
  NO2        u0037(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NAi31      u0038(.An(l), .B(m), .C(k), .Y(men_men_n67_));
  NAi21      u0039(.An(e), .B(h), .Y(men_men_n68_));
  NAi41      u0040(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n69_));
  NA2        u0041(.A(men_men_n66_), .B(men_men_n63_), .Y(men_men_n70_));
  INV        u0042(.A(m), .Y(men_men_n71_));
  NOi21      u0043(.An(k), .B(l), .Y(men_men_n72_));
  NA2        u0044(.A(men_men_n72_), .B(men_men_n71_), .Y(men_men_n73_));
  AN4        u0045(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n74_));
  NOi31      u0046(.An(h), .B(g), .C(f), .Y(men_men_n75_));
  NA2        u0047(.A(men_men_n75_), .B(men_men_n74_), .Y(men_men_n76_));
  NAi32      u0048(.An(m), .Bn(k), .C(j), .Y(men_men_n77_));
  NOi32      u0049(.An(h), .Bn(g), .C(f), .Y(men_men_n78_));
  NA2        u0050(.A(men_men_n78_), .B(men_men_n74_), .Y(men_men_n79_));
  OA220      u0051(.A0(men_men_n79_), .A1(men_men_n77_), .B0(men_men_n76_), .B1(men_men_n73_), .Y(men_men_n80_));
  NA3        u0052(.A(men_men_n80_), .B(men_men_n70_), .C(men_men_n60_), .Y(men_men_n81_));
  INV        u0053(.A(n), .Y(men_men_n82_));
  NOi32      u0054(.An(e), .Bn(b), .C(d), .Y(men_men_n83_));
  NA2        u0055(.A(men_men_n83_), .B(men_men_n82_), .Y(men_men_n84_));
  INV        u0056(.A(j), .Y(men_men_n85_));
  AN3        u0057(.A(m), .B(k), .C(i), .Y(men_men_n86_));
  NA3        u0058(.A(men_men_n86_), .B(men_men_n85_), .C(g), .Y(men_men_n87_));
  NO2        u0059(.A(men_men_n87_), .B(f), .Y(men_men_n88_));
  NAi32      u0060(.An(g), .Bn(f), .C(h), .Y(men_men_n89_));
  NAi31      u0061(.An(j), .B(m), .C(l), .Y(men_men_n90_));
  NO2        u0062(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n91_));
  NA2        u0063(.A(m), .B(l), .Y(men_men_n92_));
  NAi31      u0064(.An(k), .B(j), .C(g), .Y(men_men_n93_));
  NO3        u0065(.A(men_men_n93_), .B(men_men_n92_), .C(f), .Y(men_men_n94_));
  AN2        u0066(.A(j), .B(g), .Y(men_men_n95_));
  NOi32      u0067(.An(m), .Bn(l), .C(i), .Y(men_men_n96_));
  NOi21      u0068(.An(g), .B(i), .Y(men_men_n97_));
  NOi32      u0069(.An(m), .Bn(j), .C(k), .Y(men_men_n98_));
  AOI220     u0070(.A0(men_men_n98_), .A1(men_men_n97_), .B0(men_men_n96_), .B1(men_men_n95_), .Y(men_men_n99_));
  NO2        u0071(.A(men_men_n99_), .B(f), .Y(men_men_n100_));
  NO4        u0072(.A(men_men_n100_), .B(men_men_n94_), .C(men_men_n91_), .D(men_men_n88_), .Y(men_men_n101_));
  NAi41      u0073(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n102_));
  AN2        u0074(.A(e), .B(b), .Y(men_men_n103_));
  NOi31      u0075(.An(c), .B(h), .C(f), .Y(men_men_n104_));
  NA2        u0076(.A(men_men_n104_), .B(men_men_n103_), .Y(men_men_n105_));
  NO2        u0077(.A(men_men_n105_), .B(men_men_n102_), .Y(men_men_n106_));
  NOi21      u0078(.An(i), .B(h), .Y(men_men_n107_));
  NA3        u0079(.A(men_men_n107_), .B(g), .C(men_men_n36_), .Y(men_men_n108_));
  INV        u0080(.A(a), .Y(men_men_n109_));
  NA2        u0081(.A(men_men_n103_), .B(men_men_n109_), .Y(men_men_n110_));
  INV        u0082(.A(l), .Y(men_men_n111_));
  NOi21      u0083(.An(m), .B(n), .Y(men_men_n112_));
  AN2        u0084(.A(k), .B(h), .Y(men_men_n113_));
  NO2        u0085(.A(men_men_n108_), .B(men_men_n84_), .Y(men_men_n114_));
  INV        u0086(.A(b), .Y(men_men_n115_));
  NA2        u0087(.A(l), .B(j), .Y(men_men_n116_));
  AN2        u0088(.A(k), .B(i), .Y(men_men_n117_));
  NA2        u0089(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u0090(.A(g), .B(e), .Y(men_men_n119_));
  NOi32      u0091(.An(c), .Bn(a), .C(d), .Y(men_men_n120_));
  NA2        u0092(.A(men_men_n120_), .B(men_men_n112_), .Y(men_men_n121_));
  NO2        u0093(.A(men_men_n114_), .B(men_men_n106_), .Y(men_men_n122_));
  OAI210     u0094(.A0(men_men_n101_), .A1(men_men_n84_), .B0(men_men_n122_), .Y(men_men_n123_));
  NOi31      u0095(.An(k), .B(m), .C(j), .Y(men_men_n124_));
  NA3        u0096(.A(men_men_n124_), .B(men_men_n75_), .C(men_men_n74_), .Y(men_men_n125_));
  NOi31      u0097(.An(k), .B(m), .C(i), .Y(men_men_n126_));
  NA3        u0098(.A(men_men_n126_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n127_));
  NA2        u0099(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n128_));
  NOi32      u0100(.An(f), .Bn(b), .C(e), .Y(men_men_n129_));
  NAi21      u0101(.An(g), .B(h), .Y(men_men_n130_));
  NAi21      u0102(.An(m), .B(n), .Y(men_men_n131_));
  NAi21      u0103(.An(j), .B(k), .Y(men_men_n132_));
  NO3        u0104(.A(men_men_n132_), .B(men_men_n131_), .C(men_men_n130_), .Y(men_men_n133_));
  NAi41      u0105(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n134_));
  NAi31      u0106(.An(j), .B(k), .C(h), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n131_), .Y(men_men_n136_));
  AOI210     u0108(.A0(men_men_n133_), .A1(men_men_n129_), .B0(men_men_n136_), .Y(men_men_n137_));
  NO2        u0109(.A(k), .B(j), .Y(men_men_n138_));
  NO2        u0110(.A(men_men_n138_), .B(men_men_n131_), .Y(men_men_n139_));
  AN2        u0111(.A(k), .B(j), .Y(men_men_n140_));
  NAi21      u0112(.An(c), .B(b), .Y(men_men_n141_));
  NA2        u0113(.A(f), .B(d), .Y(men_men_n142_));
  NO3        u0114(.A(men_men_n142_), .B(men_men_n141_), .C(men_men_n130_), .Y(men_men_n143_));
  NA2        u0115(.A(h), .B(c), .Y(men_men_n144_));
  NAi31      u0116(.An(f), .B(e), .C(b), .Y(men_men_n145_));
  NA2        u0117(.A(men_men_n143_), .B(men_men_n139_), .Y(men_men_n146_));
  NA2        u0118(.A(d), .B(b), .Y(men_men_n147_));
  NAi21      u0119(.An(e), .B(f), .Y(men_men_n148_));
  NO2        u0120(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n149_));
  NA2        u0121(.A(b), .B(a), .Y(men_men_n150_));
  NAi21      u0122(.An(e), .B(g), .Y(men_men_n151_));
  NAi21      u0123(.An(c), .B(d), .Y(men_men_n152_));
  NAi31      u0124(.An(l), .B(k), .C(h), .Y(men_men_n153_));
  NO2        u0125(.A(men_men_n131_), .B(men_men_n153_), .Y(men_men_n154_));
  NA2        u0126(.A(men_men_n154_), .B(men_men_n149_), .Y(men_men_n155_));
  NAi41      u0127(.An(men_men_n128_), .B(men_men_n155_), .C(men_men_n146_), .D(men_men_n137_), .Y(men_men_n156_));
  NAi31      u0128(.An(e), .B(f), .C(b), .Y(men_men_n157_));
  NOi21      u0129(.An(g), .B(d), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n158_), .B(men_men_n157_), .Y(men_men_n159_));
  NOi21      u0131(.An(h), .B(i), .Y(men_men_n160_));
  NOi21      u0132(.An(k), .B(m), .Y(men_men_n161_));
  NA3        u0133(.A(men_men_n161_), .B(men_men_n160_), .C(n), .Y(men_men_n162_));
  NOi21      u0134(.An(men_men_n159_), .B(men_men_n162_), .Y(men_men_n163_));
  NOi21      u0135(.An(h), .B(g), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n142_), .B(men_men_n141_), .Y(men_men_n165_));
  NAi31      u0137(.An(l), .B(j), .C(h), .Y(men_men_n166_));
  NO2        u0138(.A(men_men_n166_), .B(men_men_n49_), .Y(men_men_n167_));
  NA2        u0139(.A(men_men_n167_), .B(men_men_n63_), .Y(men_men_n168_));
  NOi32      u0140(.An(n), .Bn(k), .C(m), .Y(men_men_n169_));
  INV        u0141(.A(men_men_n168_), .Y(men_men_n170_));
  NAi31      u0142(.An(d), .B(f), .C(c), .Y(men_men_n171_));
  NAi31      u0143(.An(e), .B(f), .C(c), .Y(men_men_n172_));
  NA2        u0144(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  NA2        u0145(.A(j), .B(h), .Y(men_men_n174_));
  OR3        u0146(.A(n), .B(m), .C(k), .Y(men_men_n175_));
  NO2        u0147(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  NAi32      u0148(.An(m), .Bn(k), .C(n), .Y(men_men_n177_));
  NA2        u0149(.A(men_men_n176_), .B(men_men_n173_), .Y(men_men_n178_));
  NO2        u0150(.A(n), .B(m), .Y(men_men_n179_));
  NA2        u0151(.A(men_men_n179_), .B(men_men_n50_), .Y(men_men_n180_));
  NAi21      u0152(.An(f), .B(e), .Y(men_men_n181_));
  NA2        u0153(.A(d), .B(c), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n181_), .Y(men_men_n183_));
  NOi21      u0155(.An(men_men_n183_), .B(men_men_n180_), .Y(men_men_n184_));
  NAi31      u0156(.An(m), .B(n), .C(b), .Y(men_men_n185_));
  NA2        u0157(.A(k), .B(i), .Y(men_men_n186_));
  NAi21      u0158(.An(h), .B(f), .Y(men_men_n187_));
  NO2        u0159(.A(men_men_n187_), .B(men_men_n186_), .Y(men_men_n188_));
  NO2        u0160(.A(men_men_n185_), .B(men_men_n152_), .Y(men_men_n189_));
  NA2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NOi32      u0162(.An(f), .Bn(c), .C(d), .Y(men_men_n191_));
  NOi32      u0163(.An(f), .Bn(c), .C(e), .Y(men_men_n192_));
  NO2        u0164(.A(men_men_n192_), .B(men_men_n191_), .Y(men_men_n193_));
  NO3        u0165(.A(n), .B(m), .C(j), .Y(men_men_n194_));
  NA2        u0166(.A(men_men_n194_), .B(men_men_n113_), .Y(men_men_n195_));
  AO210      u0167(.A0(men_men_n195_), .A1(men_men_n180_), .B0(men_men_n193_), .Y(men_men_n196_));
  NAi41      u0168(.An(men_men_n184_), .B(men_men_n196_), .C(men_men_n190_), .D(men_men_n178_), .Y(men_men_n197_));
  OR4        u0169(.A(men_men_n197_), .B(men_men_n170_), .C(men_men_n163_), .D(men_men_n156_), .Y(men_men_n198_));
  NO4        u0170(.A(men_men_n198_), .B(men_men_n123_), .C(men_men_n81_), .D(men_men_n52_), .Y(men_men_n199_));
  NA3        u0171(.A(m), .B(men_men_n111_), .C(j), .Y(men_men_n200_));
  NAi31      u0172(.An(n), .B(h), .C(g), .Y(men_men_n201_));
  NO2        u0173(.A(men_men_n201_), .B(men_men_n200_), .Y(men_men_n202_));
  NOi32      u0174(.An(m), .Bn(k), .C(l), .Y(men_men_n203_));
  NA3        u0175(.A(men_men_n203_), .B(men_men_n85_), .C(g), .Y(men_men_n204_));
  INV        u0176(.A(men_men_n204_), .Y(men_men_n205_));
  NA3        u0177(.A(men_men_n112_), .B(i), .C(g), .Y(men_men_n206_));
  AN2        u0178(.A(i), .B(g), .Y(men_men_n207_));
  NA3        u0179(.A(men_men_n72_), .B(men_men_n207_), .C(men_men_n112_), .Y(men_men_n208_));
  INV        u0180(.A(men_men_n206_), .Y(men_men_n209_));
  NO3        u0181(.A(men_men_n209_), .B(men_men_n205_), .C(men_men_n202_), .Y(men_men_n210_));
  NAi41      u0182(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n211_));
  INV        u0183(.A(f), .Y(men_men_n212_));
  INV        u0184(.A(g), .Y(men_men_n213_));
  NOi31      u0185(.An(i), .B(j), .C(h), .Y(men_men_n214_));
  NOi21      u0186(.An(l), .B(m), .Y(men_men_n215_));
  NA2        u0187(.A(men_men_n215_), .B(men_men_n214_), .Y(men_men_n216_));
  NO3        u0188(.A(men_men_n216_), .B(men_men_n213_), .C(men_men_n212_), .Y(men_men_n217_));
  NO2        u0189(.A(men_men_n210_), .B(men_men_n32_), .Y(men_men_n218_));
  NOi21      u0190(.An(n), .B(m), .Y(men_men_n219_));
  NOi32      u0191(.An(l), .Bn(i), .C(j), .Y(men_men_n220_));
  NA2        u0192(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n221_));
  OA220      u0193(.A0(men_men_n221_), .A1(men_men_n105_), .B0(men_men_n77_), .B1(men_men_n76_), .Y(men_men_n222_));
  NAi21      u0194(.An(j), .B(h), .Y(men_men_n223_));
  XN2        u0195(.A(i), .B(h), .Y(men_men_n224_));
  NA2        u0196(.A(men_men_n224_), .B(men_men_n223_), .Y(men_men_n225_));
  NOi31      u0197(.An(k), .B(n), .C(m), .Y(men_men_n226_));
  NOi31      u0198(.An(men_men_n226_), .B(men_men_n182_), .C(men_men_n181_), .Y(men_men_n227_));
  NA2        u0199(.A(men_men_n227_), .B(men_men_n225_), .Y(men_men_n228_));
  NAi31      u0200(.An(f), .B(e), .C(c), .Y(men_men_n229_));
  NO4        u0201(.A(men_men_n229_), .B(men_men_n175_), .C(men_men_n174_), .D(men_men_n56_), .Y(men_men_n230_));
  NA4        u0202(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n231_));
  NAi32      u0203(.An(m), .Bn(i), .C(k), .Y(men_men_n232_));
  NO3        u0204(.A(men_men_n232_), .B(men_men_n89_), .C(men_men_n231_), .Y(men_men_n233_));
  INV        u0205(.A(k), .Y(men_men_n234_));
  NO2        u0206(.A(men_men_n233_), .B(men_men_n230_), .Y(men_men_n235_));
  NAi21      u0207(.An(n), .B(a), .Y(men_men_n236_));
  NO2        u0208(.A(men_men_n236_), .B(men_men_n147_), .Y(men_men_n237_));
  NAi41      u0209(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n238_));
  NO2        u0210(.A(men_men_n238_), .B(e), .Y(men_men_n239_));
  NO3        u0211(.A(men_men_n148_), .B(men_men_n93_), .C(men_men_n92_), .Y(men_men_n240_));
  OAI210     u0212(.A0(men_men_n240_), .A1(men_men_n239_), .B0(men_men_n237_), .Y(men_men_n241_));
  AN4        u0213(.A(men_men_n241_), .B(men_men_n235_), .C(men_men_n228_), .D(men_men_n222_), .Y(men_men_n242_));
  OR2        u0214(.A(h), .B(g), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n243_), .B(men_men_n102_), .Y(men_men_n244_));
  NA2        u0216(.A(men_men_n244_), .B(men_men_n129_), .Y(men_men_n245_));
  NAi41      u0217(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n246_));
  NO2        u0218(.A(men_men_n246_), .B(men_men_n212_), .Y(men_men_n247_));
  NA2        u0219(.A(men_men_n161_), .B(men_men_n107_), .Y(men_men_n248_));
  NAi21      u0220(.An(men_men_n248_), .B(men_men_n247_), .Y(men_men_n249_));
  NO2        u0221(.A(n), .B(a), .Y(men_men_n250_));
  NAi31      u0222(.An(men_men_n238_), .B(men_men_n250_), .C(men_men_n103_), .Y(men_men_n251_));
  AN2        u0223(.A(men_men_n251_), .B(men_men_n249_), .Y(men_men_n252_));
  NAi21      u0224(.An(h), .B(i), .Y(men_men_n253_));
  NA2        u0225(.A(men_men_n179_), .B(k), .Y(men_men_n254_));
  NO2        u0226(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n255_), .B(men_men_n191_), .Y(men_men_n256_));
  NA3        u0228(.A(men_men_n256_), .B(men_men_n252_), .C(men_men_n245_), .Y(men_men_n257_));
  NOi21      u0229(.An(g), .B(e), .Y(men_men_n258_));
  NO2        u0230(.A(men_men_n69_), .B(men_men_n71_), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n253_), .B(men_men_n44_), .Y(men_men_n260_));
  NAi21      u0232(.An(f), .B(g), .Y(men_men_n261_));
  NO2        u0233(.A(men_men_n261_), .B(men_men_n61_), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n65_), .B(men_men_n116_), .Y(men_men_n263_));
  AOI220     u0235(.A0(men_men_n263_), .A1(men_men_n262_), .B0(men_men_n260_), .B1(men_men_n63_), .Y(men_men_n264_));
  INV        u0236(.A(men_men_n264_), .Y(men_men_n265_));
  NO3        u0237(.A(men_men_n132_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n266_));
  NOi41      u0238(.An(men_men_n242_), .B(men_men_n265_), .C(men_men_n257_), .D(men_men_n218_), .Y(men_men_n267_));
  NO4        u0239(.A(men_men_n202_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n268_), .B(men_men_n110_), .Y(men_men_n269_));
  NA3        u0241(.A(men_men_n56_), .B(c), .C(b), .Y(men_men_n270_));
  NAi21      u0242(.An(h), .B(g), .Y(men_men_n271_));
  OR4        u0243(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n221_), .D(e), .Y(men_men_n272_));
  NAi31      u0244(.An(g), .B(k), .C(h), .Y(men_men_n273_));
  NO3        u0245(.A(men_men_n131_), .B(men_men_n273_), .C(l), .Y(men_men_n274_));
  NAi31      u0246(.An(e), .B(d), .C(a), .Y(men_men_n275_));
  NA2        u0247(.A(men_men_n274_), .B(men_men_n129_), .Y(men_men_n276_));
  NA2        u0248(.A(men_men_n276_), .B(men_men_n272_), .Y(men_men_n277_));
  NA3        u0249(.A(men_men_n161_), .B(men_men_n160_), .C(men_men_n82_), .Y(men_men_n278_));
  NO2        u0250(.A(men_men_n278_), .B(men_men_n193_), .Y(men_men_n279_));
  INV        u0251(.A(men_men_n279_), .Y(men_men_n280_));
  NA3        u0252(.A(e), .B(c), .C(b), .Y(men_men_n281_));
  NO2        u0253(.A(d), .B(men_men_n281_), .Y(men_men_n282_));
  NAi32      u0254(.An(k), .Bn(i), .C(j), .Y(men_men_n283_));
  NAi31      u0255(.An(h), .B(l), .C(i), .Y(men_men_n284_));
  NA3        u0256(.A(men_men_n284_), .B(men_men_n283_), .C(men_men_n166_), .Y(men_men_n285_));
  NOi21      u0257(.An(men_men_n285_), .B(men_men_n49_), .Y(men_men_n286_));
  OAI210     u0258(.A0(men_men_n262_), .A1(men_men_n282_), .B0(men_men_n286_), .Y(men_men_n287_));
  NAi21      u0259(.An(l), .B(k), .Y(men_men_n288_));
  NO2        u0260(.A(men_men_n288_), .B(men_men_n49_), .Y(men_men_n289_));
  NOi21      u0261(.An(l), .B(j), .Y(men_men_n290_));
  NA2        u0262(.A(men_men_n164_), .B(men_men_n290_), .Y(men_men_n291_));
  NAi32      u0263(.An(j), .Bn(h), .C(i), .Y(men_men_n292_));
  NAi21      u0264(.An(m), .B(l), .Y(men_men_n293_));
  NO3        u0265(.A(men_men_n293_), .B(men_men_n292_), .C(men_men_n82_), .Y(men_men_n294_));
  NA2        u0266(.A(h), .B(g), .Y(men_men_n295_));
  NA2        u0267(.A(men_men_n169_), .B(men_men_n45_), .Y(men_men_n296_));
  NO2        u0268(.A(men_men_n296_), .B(men_men_n295_), .Y(men_men_n297_));
  OAI210     u0269(.A0(men_men_n297_), .A1(men_men_n294_), .B0(men_men_n165_), .Y(men_men_n298_));
  NA3        u0270(.A(men_men_n298_), .B(men_men_n287_), .C(men_men_n280_), .Y(men_men_n299_));
  NO2        u0271(.A(men_men_n145_), .B(d), .Y(men_men_n300_));
  NO2        u0272(.A(men_men_n105_), .B(men_men_n102_), .Y(men_men_n301_));
  NAi32      u0273(.An(n), .Bn(m), .C(l), .Y(men_men_n302_));
  NO2        u0274(.A(men_men_n302_), .B(men_men_n292_), .Y(men_men_n303_));
  NA2        u0275(.A(men_men_n303_), .B(men_men_n183_), .Y(men_men_n304_));
  NO2        u0276(.A(men_men_n121_), .B(men_men_n115_), .Y(men_men_n305_));
  NAi31      u0277(.An(k), .B(l), .C(j), .Y(men_men_n306_));
  OAI210     u0278(.A0(men_men_n288_), .A1(j), .B0(men_men_n306_), .Y(men_men_n307_));
  NOi21      u0279(.An(men_men_n307_), .B(men_men_n119_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n308_), .B(men_men_n305_), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n309_), .B(men_men_n304_), .Y(men_men_n310_));
  NO4        u0282(.A(men_men_n310_), .B(men_men_n299_), .C(men_men_n277_), .D(men_men_n269_), .Y(men_men_n311_));
  NA2        u0283(.A(men_men_n255_), .B(men_men_n192_), .Y(men_men_n312_));
  NAi21      u0284(.An(m), .B(k), .Y(men_men_n313_));
  NO2        u0285(.A(men_men_n224_), .B(men_men_n313_), .Y(men_men_n314_));
  NAi41      u0286(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n315_));
  NO2        u0287(.A(men_men_n315_), .B(men_men_n151_), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n316_), .B(men_men_n314_), .Y(men_men_n317_));
  NAi31      u0289(.An(i), .B(l), .C(h), .Y(men_men_n318_));
  NO4        u0290(.A(men_men_n318_), .B(men_men_n151_), .C(men_men_n69_), .D(men_men_n71_), .Y(men_men_n319_));
  NA2        u0291(.A(e), .B(c), .Y(men_men_n320_));
  NO3        u0292(.A(men_men_n320_), .B(n), .C(d), .Y(men_men_n321_));
  NOi21      u0293(.An(f), .B(h), .Y(men_men_n322_));
  NA2        u0294(.A(men_men_n322_), .B(men_men_n117_), .Y(men_men_n323_));
  NO2        u0295(.A(men_men_n323_), .B(men_men_n213_), .Y(men_men_n324_));
  NAi31      u0296(.An(d), .B(e), .C(b), .Y(men_men_n325_));
  NO2        u0297(.A(men_men_n131_), .B(men_men_n325_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n324_), .Y(men_men_n327_));
  NAi41      u0299(.An(men_men_n319_), .B(men_men_n327_), .C(men_men_n317_), .D(men_men_n312_), .Y(men_men_n328_));
  NO4        u0300(.A(men_men_n315_), .B(men_men_n77_), .C(men_men_n68_), .D(men_men_n213_), .Y(men_men_n329_));
  NA2        u0301(.A(men_men_n250_), .B(men_men_n103_), .Y(men_men_n330_));
  OR2        u0302(.A(men_men_n330_), .B(men_men_n204_), .Y(men_men_n331_));
  NOi31      u0303(.An(l), .B(n), .C(m), .Y(men_men_n332_));
  NAi21      u0304(.An(men_men_n329_), .B(men_men_n331_), .Y(men_men_n333_));
  NAi32      u0305(.An(m), .Bn(j), .C(k), .Y(men_men_n334_));
  NAi41      u0306(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n335_));
  NA2        u0307(.A(men_men_n211_), .B(men_men_n335_), .Y(men_men_n336_));
  NOi31      u0308(.An(j), .B(m), .C(k), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n124_), .B(men_men_n337_), .Y(men_men_n338_));
  AN3        u0310(.A(h), .B(g), .C(f), .Y(men_men_n339_));
  NAi31      u0311(.An(men_men_n338_), .B(men_men_n339_), .C(men_men_n336_), .Y(men_men_n340_));
  NOi32      u0312(.An(m), .Bn(j), .C(l), .Y(men_men_n341_));
  NO2        u0313(.A(men_men_n341_), .B(men_men_n96_), .Y(men_men_n342_));
  NO2        u0314(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n343_));
  NO2        u0315(.A(men_men_n216_), .B(g), .Y(men_men_n344_));
  INV        u0316(.A(men_men_n157_), .Y(men_men_n345_));
  AOI220     u0317(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n247_), .B1(men_men_n343_), .Y(men_men_n346_));
  NA2        u0318(.A(men_men_n346_), .B(men_men_n340_), .Y(men_men_n347_));
  NA3        u0319(.A(h), .B(g), .C(f), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n73_), .Y(men_men_n349_));
  NA2        u0321(.A(men_men_n164_), .B(e), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n350_), .B(men_men_n41_), .Y(men_men_n351_));
  NOi32      u0323(.An(j), .Bn(g), .C(i), .Y(men_men_n352_));
  NA3        u0324(.A(men_men_n352_), .B(men_men_n288_), .C(men_men_n112_), .Y(men_men_n353_));
  NOi32      u0325(.An(e), .Bn(b), .C(a), .Y(men_men_n354_));
  NA2        u0326(.A(men_men_n208_), .B(men_men_n35_), .Y(men_men_n355_));
  NA2        u0327(.A(men_men_n355_), .B(men_men_n354_), .Y(men_men_n356_));
  NO2        u0328(.A(men_men_n325_), .B(n), .Y(men_men_n357_));
  NA2        u0329(.A(men_men_n207_), .B(k), .Y(men_men_n358_));
  NA2        u0330(.A(m), .B(men_men_n111_), .Y(men_men_n359_));
  NO2        u0331(.A(men_men_n359_), .B(men_men_n358_), .Y(men_men_n360_));
  NAi41      u0332(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n361_));
  NA2        u0333(.A(men_men_n51_), .B(men_men_n112_), .Y(men_men_n362_));
  NA2        u0334(.A(men_men_n360_), .B(men_men_n357_), .Y(men_men_n363_));
  NA2        u0335(.A(men_men_n363_), .B(men_men_n356_), .Y(men_men_n364_));
  NO4        u0336(.A(men_men_n364_), .B(men_men_n347_), .C(men_men_n333_), .D(men_men_n328_), .Y(men_men_n365_));
  NA4        u0337(.A(men_men_n365_), .B(men_men_n311_), .C(men_men_n267_), .D(men_men_n199_), .Y(men10));
  NA3        u0338(.A(m), .B(k), .C(i), .Y(men_men_n367_));
  NO3        u0339(.A(men_men_n367_), .B(j), .C(men_men_n213_), .Y(men_men_n368_));
  NOi21      u0340(.An(e), .B(f), .Y(men_men_n369_));
  NO4        u0341(.A(men_men_n152_), .B(men_men_n369_), .C(n), .D(men_men_n109_), .Y(men_men_n370_));
  NAi31      u0342(.An(b), .B(f), .C(c), .Y(men_men_n371_));
  INV        u0343(.A(men_men_n371_), .Y(men_men_n372_));
  NOi32      u0344(.An(k), .Bn(h), .C(j), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n373_), .B(men_men_n219_), .Y(men_men_n374_));
  NA2        u0346(.A(men_men_n162_), .B(men_men_n374_), .Y(men_men_n375_));
  AOI220     u0347(.A0(men_men_n375_), .A1(men_men_n372_), .B0(men_men_n370_), .B1(men_men_n368_), .Y(men_men_n376_));
  AN2        u0348(.A(j), .B(h), .Y(men_men_n377_));
  OR2        u0349(.A(m), .B(k), .Y(men_men_n378_));
  NO2        u0350(.A(men_men_n174_), .B(men_men_n378_), .Y(men_men_n379_));
  NA4        u0351(.A(n), .B(f), .C(c), .D(men_men_n115_), .Y(men_men_n380_));
  NOi32      u0352(.An(d), .Bn(a), .C(c), .Y(men_men_n381_));
  NA2        u0353(.A(men_men_n381_), .B(men_men_n181_), .Y(men_men_n382_));
  NAi31      u0354(.An(k), .B(m), .C(j), .Y(men_men_n383_));
  NO2        u0355(.A(men_men_n380_), .B(men_men_n293_), .Y(men_men_n384_));
  NOi32      u0356(.An(f), .Bn(d), .C(c), .Y(men_men_n385_));
  NA2        u0357(.A(men_men_n384_), .B(men_men_n214_), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n386_), .B(men_men_n376_), .Y(men_men_n387_));
  NO2        u0359(.A(men_men_n56_), .B(men_men_n115_), .Y(men_men_n388_));
  NA2        u0360(.A(men_men_n250_), .B(men_men_n388_), .Y(men_men_n389_));
  INV        u0361(.A(e), .Y(men_men_n390_));
  NA2        u0362(.A(men_men_n46_), .B(e), .Y(men_men_n391_));
  OAI220     u0363(.A0(men_men_n391_), .A1(men_men_n200_), .B0(men_men_n204_), .B1(men_men_n390_), .Y(men_men_n392_));
  AN2        u0364(.A(g), .B(e), .Y(men_men_n393_));
  NA3        u0365(.A(men_men_n393_), .B(men_men_n203_), .C(i), .Y(men_men_n394_));
  INV        u0366(.A(men_men_n394_), .Y(men_men_n395_));
  NO2        u0367(.A(men_men_n99_), .B(men_men_n390_), .Y(men_men_n396_));
  NO3        u0368(.A(men_men_n396_), .B(men_men_n395_), .C(men_men_n392_), .Y(men_men_n397_));
  NOi32      u0369(.An(h), .Bn(e), .C(g), .Y(men_men_n398_));
  NA3        u0370(.A(men_men_n398_), .B(men_men_n290_), .C(m), .Y(men_men_n399_));
  NOi21      u0371(.An(g), .B(h), .Y(men_men_n400_));
  AN3        u0372(.A(m), .B(l), .C(i), .Y(men_men_n401_));
  NA3        u0373(.A(men_men_n401_), .B(men_men_n400_), .C(e), .Y(men_men_n402_));
  AN3        u0374(.A(h), .B(g), .C(e), .Y(men_men_n403_));
  NA2        u0375(.A(men_men_n403_), .B(men_men_n96_), .Y(men_men_n404_));
  AN3        u0376(.A(men_men_n404_), .B(men_men_n402_), .C(men_men_n399_), .Y(men_men_n405_));
  AOI210     u0377(.A0(men_men_n405_), .A1(men_men_n397_), .B0(men_men_n389_), .Y(men_men_n406_));
  NA3        u0378(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n407_));
  NO2        u0379(.A(men_men_n407_), .B(men_men_n389_), .Y(men_men_n408_));
  NAi31      u0380(.An(b), .B(c), .C(a), .Y(men_men_n409_));
  NO2        u0381(.A(men_men_n409_), .B(n), .Y(men_men_n410_));
  NA2        u0382(.A(men_men_n51_), .B(m), .Y(men_men_n411_));
  NO3        u0383(.A(men_men_n408_), .B(men_men_n406_), .C(men_men_n387_), .Y(men_men_n412_));
  NA2        u0384(.A(i), .B(g), .Y(men_men_n413_));
  NO3        u0385(.A(men_men_n275_), .B(men_men_n413_), .C(c), .Y(men_men_n414_));
  NOi21      u0386(.An(a), .B(n), .Y(men_men_n415_));
  NOi21      u0387(.An(d), .B(c), .Y(men_men_n416_));
  NA2        u0388(.A(men_men_n416_), .B(men_men_n415_), .Y(men_men_n417_));
  NA3        u0389(.A(i), .B(g), .C(f), .Y(men_men_n418_));
  OR2        u0390(.A(men_men_n418_), .B(men_men_n67_), .Y(men_men_n419_));
  NA3        u0391(.A(men_men_n401_), .B(men_men_n400_), .C(men_men_n181_), .Y(men_men_n420_));
  AOI210     u0392(.A0(men_men_n420_), .A1(men_men_n419_), .B0(men_men_n417_), .Y(men_men_n421_));
  AOI210     u0393(.A0(men_men_n414_), .A1(men_men_n289_), .B0(men_men_n421_), .Y(men_men_n422_));
  OR2        u0394(.A(n), .B(m), .Y(men_men_n423_));
  NO2        u0395(.A(men_men_n423_), .B(men_men_n153_), .Y(men_men_n424_));
  NO2        u0396(.A(men_men_n182_), .B(men_men_n148_), .Y(men_men_n425_));
  OAI210     u0397(.A0(men_men_n424_), .A1(men_men_n176_), .B0(men_men_n425_), .Y(men_men_n426_));
  INV        u0398(.A(men_men_n362_), .Y(men_men_n427_));
  NA3        u0399(.A(men_men_n427_), .B(men_men_n354_), .C(d), .Y(men_men_n428_));
  NO2        u0400(.A(men_men_n409_), .B(men_men_n49_), .Y(men_men_n429_));
  NAi21      u0401(.An(k), .B(j), .Y(men_men_n430_));
  NAi21      u0402(.An(e), .B(d), .Y(men_men_n431_));
  INV        u0403(.A(men_men_n431_), .Y(men_men_n432_));
  NO2        u0404(.A(men_men_n254_), .B(men_men_n212_), .Y(men_men_n433_));
  NA3        u0405(.A(men_men_n433_), .B(men_men_n432_), .C(men_men_n225_), .Y(men_men_n434_));
  NA3        u0406(.A(men_men_n434_), .B(men_men_n428_), .C(men_men_n426_), .Y(men_men_n435_));
  NOi31      u0407(.An(n), .B(m), .C(k), .Y(men_men_n436_));
  AOI220     u0408(.A0(men_men_n436_), .A1(men_men_n377_), .B0(men_men_n219_), .B1(men_men_n50_), .Y(men_men_n437_));
  NAi31      u0409(.An(g), .B(f), .C(c), .Y(men_men_n438_));
  INV        u0410(.A(men_men_n304_), .Y(men_men_n439_));
  NOi41      u0411(.An(men_men_n422_), .B(men_men_n439_), .C(men_men_n435_), .D(men_men_n265_), .Y(men_men_n440_));
  NOi32      u0412(.An(c), .Bn(a), .C(b), .Y(men_men_n441_));
  NA2        u0413(.A(men_men_n441_), .B(men_men_n112_), .Y(men_men_n442_));
  INV        u0414(.A(men_men_n273_), .Y(men_men_n443_));
  AN2        u0415(.A(e), .B(d), .Y(men_men_n444_));
  NA2        u0416(.A(men_men_n444_), .B(men_men_n443_), .Y(men_men_n445_));
  INV        u0417(.A(men_men_n148_), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n130_), .B(men_men_n41_), .Y(men_men_n447_));
  NO2        u0419(.A(men_men_n62_), .B(e), .Y(men_men_n448_));
  NA2        u0420(.A(men_men_n318_), .B(men_men_n166_), .Y(men_men_n449_));
  AOI220     u0421(.A0(men_men_n449_), .A1(men_men_n448_), .B0(men_men_n447_), .B1(men_men_n446_), .Y(men_men_n450_));
  AOI210     u0422(.A0(men_men_n450_), .A1(men_men_n445_), .B0(men_men_n442_), .Y(men_men_n451_));
  NOi21      u0423(.An(a), .B(b), .Y(men_men_n452_));
  NA3        u0424(.A(e), .B(d), .C(c), .Y(men_men_n453_));
  NAi21      u0425(.An(men_men_n453_), .B(men_men_n452_), .Y(men_men_n454_));
  AOI210     u0426(.A0(men_men_n268_), .A1(men_men_n208_), .B0(men_men_n454_), .Y(men_men_n455_));
  NO4        u0427(.A(men_men_n187_), .B(men_men_n102_), .C(men_men_n53_), .D(b), .Y(men_men_n456_));
  NA2        u0428(.A(men_men_n372_), .B(men_men_n154_), .Y(men_men_n457_));
  OR2        u0429(.A(k), .B(j), .Y(men_men_n458_));
  NA2        u0430(.A(l), .B(k), .Y(men_men_n459_));
  AOI210     u0431(.A0(men_men_n232_), .A1(men_men_n334_), .B0(men_men_n82_), .Y(men_men_n460_));
  OR3        u0432(.A(men_men_n1419_), .B(men_men_n144_), .C(men_men_n134_), .Y(men_men_n461_));
  NA2        u0433(.A(men_men_n127_), .B(men_men_n125_), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n381_), .B(men_men_n112_), .Y(men_men_n463_));
  NO4        u0435(.A(men_men_n463_), .B(men_men_n93_), .C(men_men_n111_), .D(e), .Y(men_men_n464_));
  NO3        u0436(.A(men_men_n464_), .B(men_men_n462_), .C(men_men_n319_), .Y(men_men_n465_));
  NA3        u0437(.A(men_men_n465_), .B(men_men_n461_), .C(men_men_n457_), .Y(men_men_n466_));
  NO4        u0438(.A(men_men_n466_), .B(men_men_n456_), .C(men_men_n455_), .D(men_men_n451_), .Y(men_men_n467_));
  NA2        u0439(.A(men_men_n66_), .B(men_men_n63_), .Y(men_men_n468_));
  NOi21      u0440(.An(d), .B(e), .Y(men_men_n469_));
  NO2        u0441(.A(men_men_n187_), .B(men_men_n53_), .Y(men_men_n470_));
  NAi31      u0442(.An(j), .B(l), .C(i), .Y(men_men_n471_));
  OAI210     u0443(.A0(men_men_n471_), .A1(men_men_n131_), .B0(men_men_n102_), .Y(men_men_n472_));
  NA3        u0444(.A(men_men_n472_), .B(men_men_n470_), .C(men_men_n469_), .Y(men_men_n473_));
  NO3        u0445(.A(men_men_n382_), .B(men_men_n342_), .C(men_men_n201_), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n382_), .B(men_men_n362_), .Y(men_men_n475_));
  NO4        u0447(.A(men_men_n475_), .B(men_men_n474_), .C(men_men_n184_), .D(men_men_n301_), .Y(men_men_n476_));
  NA4        u0448(.A(men_men_n476_), .B(men_men_n473_), .C(men_men_n468_), .D(men_men_n242_), .Y(men_men_n477_));
  OAI210     u0449(.A0(men_men_n126_), .A1(men_men_n124_), .B0(n), .Y(men_men_n478_));
  NO2        u0450(.A(men_men_n478_), .B(men_men_n130_), .Y(men_men_n479_));
  BUFFER     u0451(.A(men_men_n294_), .Y(men_men_n480_));
  OA210      u0452(.A0(men_men_n480_), .A1(men_men_n479_), .B0(men_men_n192_), .Y(men_men_n481_));
  XO2        u0453(.A(i), .B(h), .Y(men_men_n482_));
  NA3        u0454(.A(men_men_n482_), .B(men_men_n161_), .C(n), .Y(men_men_n483_));
  NAi41      u0455(.An(men_men_n294_), .B(men_men_n483_), .C(men_men_n437_), .D(men_men_n374_), .Y(men_men_n484_));
  NOi32      u0456(.An(men_men_n484_), .Bn(men_men_n448_), .C(men_men_n270_), .Y(men_men_n485_));
  NAi31      u0457(.An(c), .B(f), .C(d), .Y(men_men_n486_));
  AOI210     u0458(.A0(men_men_n278_), .A1(men_men_n195_), .B0(men_men_n486_), .Y(men_men_n487_));
  NOi21      u0459(.An(men_men_n80_), .B(men_men_n487_), .Y(men_men_n488_));
  NA3        u0460(.A(men_men_n370_), .B(men_men_n96_), .C(men_men_n95_), .Y(men_men_n489_));
  NA2        u0461(.A(men_men_n226_), .B(men_men_n107_), .Y(men_men_n490_));
  AOI210     u0462(.A0(men_men_n490_), .A1(men_men_n180_), .B0(men_men_n486_), .Y(men_men_n491_));
  AOI210     u0463(.A0(men_men_n353_), .A1(men_men_n35_), .B0(men_men_n454_), .Y(men_men_n492_));
  NOi31      u0464(.An(men_men_n489_), .B(men_men_n492_), .C(men_men_n491_), .Y(men_men_n493_));
  AO220      u0465(.A0(men_men_n286_), .A1(men_men_n262_), .B0(men_men_n167_), .B1(men_men_n63_), .Y(men_men_n494_));
  NA3        u0466(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n495_));
  NO2        u0467(.A(men_men_n495_), .B(men_men_n417_), .Y(men_men_n496_));
  INV        u0468(.A(men_men_n496_), .Y(men_men_n497_));
  NAi41      u0469(.An(men_men_n494_), .B(men_men_n497_), .C(men_men_n493_), .D(men_men_n488_), .Y(men_men_n498_));
  NO4        u0470(.A(men_men_n498_), .B(men_men_n485_), .C(men_men_n481_), .D(men_men_n477_), .Y(men_men_n499_));
  NA4        u0471(.A(men_men_n499_), .B(men_men_n467_), .C(men_men_n440_), .D(men_men_n412_), .Y(men11));
  NO2        u0472(.A(men_men_n69_), .B(f), .Y(men_men_n501_));
  NA2        u0473(.A(j), .B(g), .Y(men_men_n502_));
  NAi31      u0474(.An(i), .B(m), .C(l), .Y(men_men_n503_));
  NA3        u0475(.A(m), .B(k), .C(j), .Y(men_men_n504_));
  OAI220     u0476(.A0(men_men_n504_), .A1(men_men_n130_), .B0(men_men_n503_), .B1(men_men_n502_), .Y(men_men_n505_));
  NA2        u0477(.A(men_men_n505_), .B(men_men_n501_), .Y(men_men_n506_));
  NOi32      u0478(.An(e), .Bn(b), .C(f), .Y(men_men_n507_));
  NA2        u0479(.A(j), .B(men_men_n112_), .Y(men_men_n508_));
  NA2        u0480(.A(men_men_n46_), .B(j), .Y(men_men_n509_));
  NO2        u0481(.A(men_men_n509_), .B(men_men_n296_), .Y(men_men_n510_));
  NAi31      u0482(.An(d), .B(e), .C(a), .Y(men_men_n511_));
  NO2        u0483(.A(men_men_n511_), .B(n), .Y(men_men_n512_));
  AOI220     u0484(.A0(men_men_n512_), .A1(men_men_n100_), .B0(men_men_n510_), .B1(men_men_n507_), .Y(men_men_n513_));
  NAi41      u0485(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n514_));
  AN2        u0486(.A(men_men_n514_), .B(men_men_n361_), .Y(men_men_n515_));
  AOI210     u0487(.A0(men_men_n515_), .A1(men_men_n382_), .B0(men_men_n271_), .Y(men_men_n516_));
  NA2        u0488(.A(j), .B(i), .Y(men_men_n517_));
  NAi31      u0489(.An(n), .B(m), .C(k), .Y(men_men_n518_));
  NO3        u0490(.A(men_men_n518_), .B(men_men_n517_), .C(men_men_n111_), .Y(men_men_n519_));
  NO2        u0491(.A(n), .B(men_men_n150_), .Y(men_men_n520_));
  NOi32      u0492(.An(g), .Bn(f), .C(i), .Y(men_men_n521_));
  NA2        u0493(.A(men_men_n521_), .B(men_men_n98_), .Y(men_men_n522_));
  NO2        u0494(.A(men_men_n273_), .B(men_men_n49_), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n522_), .B(n), .Y(men_men_n524_));
  AOI210     u0496(.A0(men_men_n519_), .A1(men_men_n516_), .B0(men_men_n524_), .Y(men_men_n525_));
  NA2        u0497(.A(men_men_n140_), .B(men_men_n34_), .Y(men_men_n526_));
  OAI220     u0498(.A0(men_men_n526_), .A1(m), .B0(men_men_n509_), .B1(men_men_n232_), .Y(men_men_n527_));
  NOi41      u0499(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n528_));
  NAi32      u0500(.An(e), .Bn(b), .C(c), .Y(men_men_n529_));
  OR2        u0501(.A(men_men_n529_), .B(men_men_n82_), .Y(men_men_n530_));
  AN2        u0502(.A(men_men_n335_), .B(men_men_n315_), .Y(men_men_n531_));
  NA2        u0503(.A(men_men_n531_), .B(men_men_n530_), .Y(men_men_n532_));
  AN2        u0504(.A(men_men_n532_), .B(men_men_n527_), .Y(men_men_n533_));
  OAI220     u0505(.A0(men_men_n383_), .A1(i), .B0(men_men_n503_), .B1(men_men_n502_), .Y(men_men_n534_));
  NAi31      u0506(.An(d), .B(c), .C(a), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n535_), .B(n), .Y(men_men_n536_));
  NA3        u0508(.A(men_men_n536_), .B(men_men_n534_), .C(e), .Y(men_men_n537_));
  NO3        u0509(.A(men_men_n58_), .B(men_men_n49_), .C(men_men_n213_), .Y(men_men_n538_));
  NO2        u0510(.A(men_men_n229_), .B(men_men_n109_), .Y(men_men_n539_));
  NA2        u0511(.A(men_men_n538_), .B(men_men_n539_), .Y(men_men_n540_));
  NA2        u0512(.A(men_men_n540_), .B(men_men_n537_), .Y(men_men_n541_));
  NO2        u0513(.A(men_men_n275_), .B(n), .Y(men_men_n542_));
  NAi32      u0514(.An(d), .Bn(a), .C(b), .Y(men_men_n543_));
  NO2        u0515(.A(men_men_n543_), .B(men_men_n49_), .Y(men_men_n544_));
  NA2        u0516(.A(h), .B(f), .Y(men_men_n545_));
  NO2        u0517(.A(men_men_n545_), .B(men_men_n93_), .Y(men_men_n546_));
  NO2        u0518(.A(men_men_n177_), .B(men_men_n174_), .Y(men_men_n547_));
  AOI220     u0519(.A0(men_men_n547_), .A1(men_men_n55_), .B0(men_men_n546_), .B1(men_men_n544_), .Y(men_men_n548_));
  INV        u0520(.A(men_men_n548_), .Y(men_men_n549_));
  NO2        u0521(.A(men_men_n147_), .B(c), .Y(men_men_n550_));
  NA3        u0522(.A(f), .B(d), .C(b), .Y(men_men_n551_));
  NO3        u0523(.A(men_men_n551_), .B(men_men_n177_), .C(men_men_n174_), .Y(men_men_n552_));
  NO4        u0524(.A(men_men_n552_), .B(men_men_n549_), .C(men_men_n541_), .D(men_men_n533_), .Y(men_men_n553_));
  AN4        u0525(.A(men_men_n553_), .B(men_men_n525_), .C(men_men_n513_), .D(men_men_n506_), .Y(men_men_n554_));
  INV        u0526(.A(k), .Y(men_men_n555_));
  NA3        u0527(.A(l), .B(men_men_n555_), .C(i), .Y(men_men_n556_));
  INV        u0528(.A(men_men_n556_), .Y(men_men_n557_));
  NA4        u0529(.A(men_men_n381_), .B(men_men_n400_), .C(men_men_n181_), .D(men_men_n112_), .Y(men_men_n558_));
  NAi32      u0530(.An(h), .Bn(f), .C(g), .Y(men_men_n559_));
  NAi41      u0531(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n560_));
  OAI210     u0532(.A0(men_men_n511_), .A1(n), .B0(men_men_n560_), .Y(men_men_n561_));
  NA2        u0533(.A(men_men_n561_), .B(m), .Y(men_men_n562_));
  NAi31      u0534(.An(h), .B(g), .C(f), .Y(men_men_n563_));
  OR3        u0535(.A(men_men_n563_), .B(men_men_n275_), .C(men_men_n49_), .Y(men_men_n564_));
  NA4        u0536(.A(men_men_n400_), .B(men_men_n120_), .C(men_men_n112_), .D(e), .Y(men_men_n565_));
  AN2        u0537(.A(men_men_n565_), .B(men_men_n564_), .Y(men_men_n566_));
  OA210      u0538(.A0(men_men_n562_), .A1(men_men_n559_), .B0(men_men_n566_), .Y(men_men_n567_));
  NA2        u0539(.A(men_men_n567_), .B(men_men_n558_), .Y(men_men_n568_));
  NAi31      u0540(.An(f), .B(h), .C(g), .Y(men_men_n569_));
  NO4        u0541(.A(men_men_n306_), .B(men_men_n569_), .C(men_men_n69_), .D(men_men_n71_), .Y(men_men_n570_));
  NOi41      u0542(.An(a), .B(men_men_n348_), .C(men_men_n65_), .D(men_men_n116_), .Y(men_men_n571_));
  OR2        u0543(.A(men_men_n571_), .B(men_men_n570_), .Y(men_men_n572_));
  NOi32      u0544(.An(d), .Bn(a), .C(e), .Y(men_men_n573_));
  NA2        u0545(.A(men_men_n573_), .B(men_men_n112_), .Y(men_men_n574_));
  NO2        u0546(.A(n), .B(c), .Y(men_men_n575_));
  NA3        u0547(.A(men_men_n575_), .B(men_men_n29_), .C(m), .Y(men_men_n576_));
  NAi32      u0548(.An(n), .Bn(f), .C(m), .Y(men_men_n577_));
  NOi32      u0549(.An(e), .Bn(a), .C(d), .Y(men_men_n578_));
  INV        u0550(.A(men_men_n578_), .Y(men_men_n579_));
  NO2        u0551(.A(men_men_n579_), .B(men_men_n526_), .Y(men_men_n580_));
  AOI210     u0552(.A0(men_men_n580_), .A1(men_men_n1417_), .B0(men_men_n572_), .Y(men_men_n581_));
  OAI210     u0553(.A0(men_men_n249_), .A1(men_men_n85_), .B0(men_men_n581_), .Y(men_men_n582_));
  AOI210     u0554(.A0(men_men_n568_), .A1(men_men_n557_), .B0(men_men_n582_), .Y(men_men_n583_));
  NO3        u0555(.A(men_men_n313_), .B(men_men_n57_), .C(n), .Y(men_men_n584_));
  NA3        u0556(.A(men_men_n486_), .B(men_men_n172_), .C(men_men_n171_), .Y(men_men_n585_));
  NA2        u0557(.A(men_men_n438_), .B(men_men_n229_), .Y(men_men_n586_));
  OR2        u0558(.A(men_men_n586_), .B(men_men_n585_), .Y(men_men_n587_));
  NA2        u0559(.A(men_men_n72_), .B(men_men_n112_), .Y(men_men_n588_));
  NO2        u0560(.A(men_men_n588_), .B(men_men_n45_), .Y(men_men_n589_));
  AOI220     u0561(.A0(men_men_n589_), .A1(men_men_n516_), .B0(men_men_n587_), .B1(men_men_n584_), .Y(men_men_n590_));
  NO2        u0562(.A(men_men_n590_), .B(men_men_n85_), .Y(men_men_n591_));
  NA3        u0563(.A(men_men_n528_), .B(men_men_n337_), .C(men_men_n46_), .Y(men_men_n592_));
  NOi32      u0564(.An(e), .Bn(c), .C(f), .Y(men_men_n593_));
  NOi21      u0565(.An(f), .B(g), .Y(men_men_n594_));
  NO2        u0566(.A(men_men_n594_), .B(men_men_n211_), .Y(men_men_n595_));
  AOI220     u0567(.A0(men_men_n595_), .A1(men_men_n379_), .B0(men_men_n593_), .B1(men_men_n176_), .Y(men_men_n596_));
  NA3        u0568(.A(men_men_n596_), .B(men_men_n592_), .C(men_men_n178_), .Y(men_men_n597_));
  AOI210     u0569(.A0(men_men_n515_), .A1(men_men_n382_), .B0(men_men_n295_), .Y(men_men_n598_));
  NA2        u0570(.A(men_men_n598_), .B(men_men_n263_), .Y(men_men_n599_));
  NOi21      u0571(.An(j), .B(l), .Y(men_men_n600_));
  NAi21      u0572(.An(k), .B(h), .Y(men_men_n601_));
  NO2        u0573(.A(men_men_n601_), .B(men_men_n261_), .Y(men_men_n602_));
  NA2        u0574(.A(men_men_n602_), .B(men_men_n600_), .Y(men_men_n603_));
  OR2        u0575(.A(men_men_n603_), .B(men_men_n562_), .Y(men_men_n604_));
  NOi31      u0576(.An(m), .B(n), .C(k), .Y(men_men_n605_));
  NA2        u0577(.A(men_men_n600_), .B(men_men_n605_), .Y(men_men_n606_));
  NO2        u0578(.A(men_men_n275_), .B(men_men_n49_), .Y(men_men_n607_));
  NO2        u0579(.A(men_men_n306_), .B(men_men_n569_), .Y(men_men_n608_));
  NO2        u0580(.A(men_men_n511_), .B(men_men_n49_), .Y(men_men_n609_));
  NA2        u0581(.A(men_men_n609_), .B(men_men_n608_), .Y(men_men_n610_));
  NA3        u0582(.A(men_men_n610_), .B(men_men_n604_), .C(men_men_n599_), .Y(men_men_n611_));
  NA2        u0583(.A(men_men_n107_), .B(men_men_n36_), .Y(men_men_n612_));
  NO2        u0584(.A(k), .B(men_men_n213_), .Y(men_men_n613_));
  NO2        u0585(.A(men_men_n507_), .B(men_men_n354_), .Y(men_men_n614_));
  NO2        u0586(.A(men_men_n614_), .B(n), .Y(men_men_n615_));
  NAi31      u0587(.An(men_men_n612_), .B(men_men_n615_), .C(men_men_n613_), .Y(men_men_n616_));
  NO2        u0588(.A(men_men_n509_), .B(men_men_n177_), .Y(men_men_n617_));
  NA3        u0589(.A(men_men_n529_), .B(men_men_n270_), .C(men_men_n145_), .Y(men_men_n618_));
  NA2        u0590(.A(men_men_n482_), .B(men_men_n161_), .Y(men_men_n619_));
  NO3        u0591(.A(men_men_n380_), .B(men_men_n619_), .C(men_men_n85_), .Y(men_men_n620_));
  AOI210     u0592(.A0(men_men_n618_), .A1(men_men_n617_), .B0(men_men_n620_), .Y(men_men_n621_));
  AN3        u0593(.A(f), .B(d), .C(b), .Y(men_men_n622_));
  OAI210     u0594(.A0(men_men_n622_), .A1(men_men_n129_), .B0(n), .Y(men_men_n623_));
  NA3        u0595(.A(men_men_n482_), .B(men_men_n161_), .C(men_men_n213_), .Y(men_men_n624_));
  AOI210     u0596(.A0(men_men_n623_), .A1(men_men_n231_), .B0(men_men_n624_), .Y(men_men_n625_));
  NAi31      u0597(.An(m), .B(n), .C(k), .Y(men_men_n626_));
  OR2        u0598(.A(men_men_n134_), .B(men_men_n57_), .Y(men_men_n627_));
  OAI210     u0599(.A0(men_men_n627_), .A1(men_men_n626_), .B0(men_men_n251_), .Y(men_men_n628_));
  OAI210     u0600(.A0(men_men_n628_), .A1(men_men_n625_), .B0(j), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n629_), .B(men_men_n621_), .C(men_men_n616_), .Y(men_men_n630_));
  NO4        u0602(.A(men_men_n630_), .B(men_men_n611_), .C(men_men_n597_), .D(men_men_n591_), .Y(men_men_n631_));
  NA2        u0603(.A(men_men_n370_), .B(men_men_n164_), .Y(men_men_n632_));
  NAi31      u0604(.An(g), .B(h), .C(f), .Y(men_men_n633_));
  OA210      u0605(.A0(men_men_n511_), .A1(n), .B0(men_men_n560_), .Y(men_men_n634_));
  NO2        u0606(.A(men_men_n632_), .B(men_men_n504_), .Y(men_men_n635_));
  NO3        u0607(.A(g), .B(men_men_n212_), .C(men_men_n53_), .Y(men_men_n636_));
  NO2        u0608(.A(men_men_n490_), .B(men_men_n85_), .Y(men_men_n637_));
  OAI210     u0609(.A0(men_men_n637_), .A1(men_men_n379_), .B0(men_men_n636_), .Y(men_men_n638_));
  INV        u0610(.A(men_men_n339_), .Y(men_men_n639_));
  OA220      u0611(.A0(men_men_n606_), .A1(men_men_n639_), .B0(men_men_n603_), .B1(men_men_n69_), .Y(men_men_n640_));
  NA3        u0612(.A(men_men_n501_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n641_));
  AN2        u0613(.A(h), .B(f), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n642_), .B(men_men_n37_), .Y(men_men_n643_));
  AOI210     u0615(.A0(men_men_n543_), .A1(men_men_n409_), .B0(men_men_n49_), .Y(men_men_n644_));
  NA3        u0616(.A(men_men_n641_), .B(men_men_n640_), .C(men_men_n638_), .Y(men_men_n645_));
  NO2        u0617(.A(men_men_n253_), .B(f), .Y(men_men_n646_));
  NO3        u0618(.A(h), .B(men_men_n646_), .C(men_men_n34_), .Y(men_men_n647_));
  NA2        u0619(.A(men_men_n326_), .B(men_men_n140_), .Y(men_men_n648_));
  NA2        u0620(.A(men_men_n131_), .B(men_men_n49_), .Y(men_men_n649_));
  OR2        u0621(.A(men_men_n353_), .B(men_men_n110_), .Y(men_men_n650_));
  OAI210     u0622(.A0(men_men_n648_), .A1(men_men_n647_), .B0(men_men_n650_), .Y(men_men_n651_));
  NO3        u0623(.A(men_men_n385_), .B(men_men_n192_), .C(men_men_n191_), .Y(men_men_n652_));
  NA2        u0624(.A(men_men_n652_), .B(men_men_n229_), .Y(men_men_n653_));
  NA3        u0625(.A(men_men_n653_), .B(men_men_n255_), .C(j), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n441_), .B(men_men_n82_), .Y(men_men_n655_));
  NO4        u0627(.A(men_men_n504_), .B(men_men_n655_), .C(men_men_n130_), .D(men_men_n212_), .Y(men_men_n656_));
  INV        u0628(.A(men_men_n656_), .Y(men_men_n657_));
  NA3        u0629(.A(men_men_n657_), .B(men_men_n654_), .C(men_men_n489_), .Y(men_men_n658_));
  NO4        u0630(.A(men_men_n658_), .B(men_men_n651_), .C(men_men_n645_), .D(men_men_n635_), .Y(men_men_n659_));
  NA4        u0631(.A(men_men_n659_), .B(men_men_n631_), .C(men_men_n583_), .D(men_men_n554_), .Y(men08));
  NO2        u0632(.A(k), .B(h), .Y(men_men_n661_));
  AO210      u0633(.A0(men_men_n253_), .A1(men_men_n430_), .B0(men_men_n661_), .Y(men_men_n662_));
  NO2        u0634(.A(men_men_n662_), .B(men_men_n293_), .Y(men_men_n663_));
  NA2        u0635(.A(men_men_n593_), .B(men_men_n82_), .Y(men_men_n664_));
  NA2        u0636(.A(men_men_n664_), .B(men_men_n438_), .Y(men_men_n665_));
  NA2        u0637(.A(men_men_n665_), .B(men_men_n663_), .Y(men_men_n666_));
  NA2        u0638(.A(men_men_n82_), .B(men_men_n109_), .Y(men_men_n667_));
  NO2        u0639(.A(men_men_n667_), .B(men_men_n54_), .Y(men_men_n668_));
  NA2        u0640(.A(men_men_n551_), .B(men_men_n231_), .Y(men_men_n669_));
  NA2        u0641(.A(men_men_n669_), .B(men_men_n344_), .Y(men_men_n670_));
  AOI210     u0642(.A0(men_men_n551_), .A1(men_men_n157_), .B0(men_men_n82_), .Y(men_men_n671_));
  NA4        u0643(.A(men_men_n215_), .B(men_men_n140_), .C(men_men_n45_), .D(h), .Y(men_men_n672_));
  AN2        u0644(.A(l), .B(k), .Y(men_men_n673_));
  NA4        u0645(.A(men_men_n673_), .B(men_men_n107_), .C(men_men_n71_), .D(men_men_n213_), .Y(men_men_n674_));
  OAI210     u0646(.A0(men_men_n672_), .A1(g), .B0(men_men_n674_), .Y(men_men_n675_));
  NA2        u0647(.A(men_men_n675_), .B(men_men_n671_), .Y(men_men_n676_));
  NA4        u0648(.A(men_men_n676_), .B(men_men_n670_), .C(men_men_n666_), .D(men_men_n346_), .Y(men_men_n677_));
  AN2        u0649(.A(men_men_n512_), .B(men_men_n94_), .Y(men_men_n678_));
  NO4        u0650(.A(men_men_n174_), .B(men_men_n378_), .C(men_men_n111_), .D(g), .Y(men_men_n679_));
  AOI210     u0651(.A0(men_men_n679_), .A1(men_men_n669_), .B0(men_men_n496_), .Y(men_men_n680_));
  NO2        u0652(.A(men_men_n38_), .B(men_men_n212_), .Y(men_men_n681_));
  AOI220     u0653(.A0(men_men_n595_), .A1(men_men_n343_), .B0(men_men_n681_), .B1(men_men_n542_), .Y(men_men_n682_));
  NAi31      u0654(.An(men_men_n678_), .B(men_men_n682_), .C(men_men_n680_), .Y(men_men_n683_));
  NO2        u0655(.A(men_men_n515_), .B(men_men_n35_), .Y(men_men_n684_));
  OAI210     u0656(.A0(men_men_n529_), .A1(men_men_n47_), .B0(men_men_n627_), .Y(men_men_n685_));
  NO2        u0657(.A(men_men_n459_), .B(men_men_n131_), .Y(men_men_n686_));
  AOI210     u0658(.A0(men_men_n686_), .A1(men_men_n685_), .B0(men_men_n684_), .Y(men_men_n687_));
  NO3        u0659(.A(men_men_n313_), .B(men_men_n130_), .C(men_men_n41_), .Y(men_men_n688_));
  NAi21      u0660(.An(men_men_n688_), .B(men_men_n674_), .Y(men_men_n689_));
  AOI220     u0661(.A0(men_men_n1418_), .A1(men_men_n384_), .B0(men_men_n689_), .B1(men_men_n74_), .Y(men_men_n690_));
  OAI210     u0662(.A0(men_men_n687_), .A1(men_men_n85_), .B0(men_men_n690_), .Y(men_men_n691_));
  NA2        u0663(.A(men_men_n354_), .B(men_men_n43_), .Y(men_men_n692_));
  NA3        u0664(.A(men_men_n653_), .B(men_men_n332_), .C(men_men_n373_), .Y(men_men_n693_));
  NA2        u0665(.A(men_men_n673_), .B(men_men_n219_), .Y(men_men_n694_));
  NO2        u0666(.A(men_men_n694_), .B(men_men_n325_), .Y(men_men_n695_));
  AOI210     u0667(.A0(men_men_n695_), .A1(men_men_n646_), .B0(men_men_n464_), .Y(men_men_n696_));
  NA3        u0668(.A(m), .B(l), .C(k), .Y(men_men_n697_));
  NO2        u0669(.A(men_men_n514_), .B(men_men_n271_), .Y(men_men_n698_));
  NOi21      u0670(.An(men_men_n698_), .B(men_men_n508_), .Y(men_men_n699_));
  NA4        u0671(.A(men_men_n112_), .B(l), .C(k), .D(men_men_n85_), .Y(men_men_n700_));
  INV        u0672(.A(men_men_n699_), .Y(men_men_n701_));
  NA4        u0673(.A(men_men_n701_), .B(men_men_n696_), .C(men_men_n693_), .D(men_men_n692_), .Y(men_men_n702_));
  NO4        u0674(.A(men_men_n702_), .B(men_men_n691_), .C(men_men_n683_), .D(men_men_n677_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n595_), .B(men_men_n379_), .Y(men_men_n704_));
  NOi31      u0676(.An(g), .B(h), .C(f), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n609_), .B(men_men_n705_), .Y(men_men_n706_));
  AO210      u0678(.A0(men_men_n706_), .A1(men_men_n564_), .B0(men_men_n517_), .Y(men_men_n707_));
  NO3        u0679(.A(men_men_n382_), .B(men_men_n502_), .C(h), .Y(men_men_n708_));
  AOI210     u0680(.A0(men_men_n708_), .A1(men_men_n112_), .B0(men_men_n475_), .Y(men_men_n709_));
  NA4        u0681(.A(men_men_n709_), .B(men_men_n707_), .C(men_men_n704_), .D(men_men_n252_), .Y(men_men_n710_));
  NA2        u0682(.A(men_men_n673_), .B(men_men_n71_), .Y(men_men_n711_));
  NO4        u0683(.A(men_men_n652_), .B(men_men_n174_), .C(n), .D(i), .Y(men_men_n712_));
  NOi21      u0684(.An(h), .B(j), .Y(men_men_n713_));
  NA2        u0685(.A(men_men_n713_), .B(f), .Y(men_men_n714_));
  NO2        u0686(.A(men_men_n714_), .B(men_men_n246_), .Y(men_men_n715_));
  NO2        u0687(.A(men_men_n715_), .B(men_men_n712_), .Y(men_men_n716_));
  OAI220     u0688(.A0(men_men_n716_), .A1(men_men_n711_), .B0(men_men_n566_), .B1(men_men_n58_), .Y(men_men_n717_));
  AOI210     u0689(.A0(men_men_n710_), .A1(l), .B0(men_men_n717_), .Y(men_men_n718_));
  NO2        u0690(.A(j), .B(i), .Y(men_men_n719_));
  NA3        u0691(.A(men_men_n719_), .B(men_men_n78_), .C(l), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n719_), .B(men_men_n33_), .Y(men_men_n721_));
  NA2        u0693(.A(men_men_n403_), .B(men_men_n120_), .Y(men_men_n722_));
  OA220      u0694(.A0(men_men_n722_), .A1(men_men_n721_), .B0(men_men_n720_), .B1(men_men_n562_), .Y(men_men_n723_));
  NO3        u0695(.A(men_men_n152_), .B(men_men_n49_), .C(men_men_n109_), .Y(men_men_n724_));
  NO3        u0696(.A(n), .B(men_men_n150_), .C(men_men_n71_), .Y(men_men_n725_));
  NO3        u0697(.A(men_men_n459_), .B(men_men_n418_), .C(j), .Y(men_men_n726_));
  OAI210     u0698(.A0(men_men_n725_), .A1(men_men_n724_), .B0(men_men_n726_), .Y(men_men_n727_));
  OAI210     u0699(.A0(men_men_n706_), .A1(men_men_n58_), .B0(men_men_n727_), .Y(men_men_n728_));
  NO2        u0700(.A(men_men_n293_), .B(men_men_n40_), .Y(men_men_n729_));
  AOI210     u0701(.A0(men_men_n507_), .A1(n), .B0(men_men_n528_), .Y(men_men_n730_));
  NA2        u0702(.A(men_men_n730_), .B(men_men_n531_), .Y(men_men_n731_));
  AN3        u0703(.A(men_men_n731_), .B(men_men_n729_), .C(men_men_n97_), .Y(men_men_n732_));
  NO3        u0704(.A(men_men_n174_), .B(men_men_n378_), .C(men_men_n111_), .Y(men_men_n733_));
  AOI220     u0705(.A0(men_men_n733_), .A1(men_men_n247_), .B0(men_men_n586_), .B1(men_men_n303_), .Y(men_men_n734_));
  INV        u0706(.A(men_men_n734_), .Y(men_men_n735_));
  NA2        u0707(.A(men_men_n688_), .B(men_men_n671_), .Y(men_men_n736_));
  NO2        u0708(.A(men_men_n697_), .B(men_men_n89_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n737_), .B(men_men_n561_), .Y(men_men_n738_));
  NO2        u0710(.A(men_men_n563_), .B(men_men_n116_), .Y(men_men_n739_));
  OAI210     u0711(.A0(men_men_n739_), .A1(men_men_n726_), .B0(men_men_n644_), .Y(men_men_n740_));
  NA3        u0712(.A(men_men_n740_), .B(men_men_n738_), .C(men_men_n736_), .Y(men_men_n741_));
  OR4        u0713(.A(men_men_n741_), .B(men_men_n735_), .C(men_men_n732_), .D(men_men_n728_), .Y(men_men_n742_));
  NA3        u0714(.A(men_men_n730_), .B(men_men_n531_), .C(men_men_n530_), .Y(men_men_n743_));
  NA4        u0715(.A(men_men_n743_), .B(men_men_n215_), .C(men_men_n430_), .D(men_men_n34_), .Y(men_men_n744_));
  NO4        u0716(.A(men_men_n459_), .B(men_men_n413_), .C(j), .D(f), .Y(men_men_n745_));
  NO2        u0717(.A(men_men_n672_), .B(men_men_n664_), .Y(men_men_n746_));
  AOI210     u0718(.A0(men_men_n745_), .A1(men_men_n259_), .B0(men_men_n746_), .Y(men_men_n747_));
  NA3        u0719(.A(men_men_n521_), .B(men_men_n290_), .C(h), .Y(men_men_n748_));
  NOi21      u0720(.An(men_men_n644_), .B(men_men_n748_), .Y(men_men_n749_));
  NO2        u0721(.A(men_men_n90_), .B(men_men_n47_), .Y(men_men_n750_));
  OAI220     u0722(.A0(men_men_n748_), .A1(men_men_n576_), .B0(men_men_n720_), .B1(men_men_n69_), .Y(men_men_n751_));
  AOI210     u0723(.A0(men_men_n750_), .A1(men_men_n615_), .B0(men_men_n751_), .Y(men_men_n752_));
  NAi41      u0724(.An(men_men_n749_), .B(men_men_n752_), .C(men_men_n747_), .D(men_men_n744_), .Y(men_men_n753_));
  OR2        u0725(.A(men_men_n737_), .B(men_men_n94_), .Y(men_men_n754_));
  NA2        u0726(.A(men_men_n754_), .B(men_men_n237_), .Y(men_men_n755_));
  NO2        u0727(.A(men_men_n634_), .B(men_men_n71_), .Y(men_men_n756_));
  NA2        u0728(.A(men_men_n745_), .B(men_men_n756_), .Y(men_men_n757_));
  INV        u0729(.A(men_men_n495_), .Y(men_men_n758_));
  NA3        u0730(.A(men_men_n250_), .B(men_men_n56_), .C(b), .Y(men_men_n759_));
  AOI220     u0731(.A0(men_men_n575_), .A1(men_men_n29_), .B0(men_men_n441_), .B1(men_men_n82_), .Y(men_men_n760_));
  NA2        u0732(.A(men_men_n760_), .B(men_men_n759_), .Y(men_men_n761_));
  NO2        u0733(.A(men_men_n748_), .B(men_men_n463_), .Y(men_men_n762_));
  AOI210     u0734(.A0(men_men_n761_), .A1(men_men_n758_), .B0(men_men_n762_), .Y(men_men_n763_));
  NA3        u0735(.A(men_men_n763_), .B(men_men_n757_), .C(men_men_n755_), .Y(men_men_n764_));
  NOi41      u0736(.An(men_men_n723_), .B(men_men_n764_), .C(men_men_n753_), .D(men_men_n742_), .Y(men_men_n765_));
  OR2        u0737(.A(men_men_n672_), .B(men_men_n231_), .Y(men_men_n766_));
  NO3        u0738(.A(men_men_n338_), .B(men_men_n295_), .C(men_men_n111_), .Y(men_men_n767_));
  NA2        u0739(.A(men_men_n767_), .B(men_men_n731_), .Y(men_men_n768_));
  NA2        u0740(.A(men_men_n46_), .B(men_men_n53_), .Y(men_men_n769_));
  NO3        u0741(.A(men_men_n769_), .B(men_men_n721_), .C(men_men_n275_), .Y(men_men_n770_));
  NO3        u0742(.A(men_men_n502_), .B(men_men_n92_), .C(h), .Y(men_men_n771_));
  AOI210     u0743(.A0(men_men_n771_), .A1(men_men_n668_), .B0(men_men_n770_), .Y(men_men_n772_));
  NA4        u0744(.A(men_men_n772_), .B(men_men_n768_), .C(men_men_n766_), .D(men_men_n386_), .Y(men_men_n773_));
  OR2        u0745(.A(men_men_n633_), .B(men_men_n90_), .Y(men_men_n774_));
  NOi31      u0746(.An(b), .B(d), .C(a), .Y(men_men_n775_));
  NO2        u0747(.A(men_men_n775_), .B(men_men_n573_), .Y(men_men_n776_));
  NO2        u0748(.A(men_men_n776_), .B(n), .Y(men_men_n777_));
  NOi21      u0749(.An(men_men_n760_), .B(men_men_n777_), .Y(men_men_n778_));
  OAI220     u0750(.A0(men_men_n778_), .A1(men_men_n774_), .B0(men_men_n748_), .B1(men_men_n574_), .Y(men_men_n779_));
  NO2        u0751(.A(men_men_n529_), .B(men_men_n82_), .Y(men_men_n780_));
  NO2        u0752(.A(men_men_n325_), .B(men_men_n116_), .Y(men_men_n781_));
  NOi21      u0753(.An(men_men_n781_), .B(men_men_n162_), .Y(men_men_n782_));
  AOI210     u0754(.A0(men_men_n767_), .A1(men_men_n780_), .B0(men_men_n782_), .Y(men_men_n783_));
  OAI210     u0755(.A0(men_men_n672_), .A1(men_men_n380_), .B0(men_men_n783_), .Y(men_men_n784_));
  NO2        u0756(.A(men_men_n652_), .B(n), .Y(men_men_n785_));
  NA2        u0757(.A(men_men_n785_), .B(men_men_n663_), .Y(men_men_n786_));
  NO2        u0758(.A(men_men_n320_), .B(men_men_n236_), .Y(men_men_n787_));
  OAI210     u0759(.A0(men_men_n94_), .A1(men_men_n91_), .B0(men_men_n787_), .Y(men_men_n788_));
  NA2        u0760(.A(men_men_n120_), .B(men_men_n82_), .Y(men_men_n789_));
  AOI210     u0761(.A0(men_men_n407_), .A1(men_men_n399_), .B0(men_men_n789_), .Y(men_men_n790_));
  NAi21      u0762(.An(men_men_n790_), .B(men_men_n788_), .Y(men_men_n791_));
  NA2        u0763(.A(men_men_n695_), .B(men_men_n34_), .Y(men_men_n792_));
  NAi21      u0764(.An(men_men_n700_), .B(men_men_n414_), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n271_), .B(i), .Y(men_men_n794_));
  NAi41      u0766(.An(men_men_n791_), .B(men_men_n793_), .C(men_men_n792_), .D(men_men_n786_), .Y(men_men_n795_));
  NO4        u0767(.A(men_men_n795_), .B(men_men_n784_), .C(men_men_n779_), .D(men_men_n773_), .Y(men_men_n796_));
  NA4        u0768(.A(men_men_n796_), .B(men_men_n765_), .C(men_men_n718_), .D(men_men_n703_), .Y(men09));
  INV        u0769(.A(men_men_n121_), .Y(men_men_n798_));
  NA2        u0770(.A(f), .B(e), .Y(men_men_n799_));
  NO2        u0771(.A(men_men_n224_), .B(men_men_n111_), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n800_), .B(g), .Y(men_men_n801_));
  AOI210     u0773(.A0(men_men_n1420_), .A1(g), .B0(men_men_n447_), .Y(men_men_n802_));
  AOI210     u0774(.A0(men_men_n802_), .A1(men_men_n801_), .B0(men_men_n799_), .Y(men_men_n803_));
  NA2        u0775(.A(men_men_n424_), .B(e), .Y(men_men_n804_));
  NO2        u0776(.A(men_men_n804_), .B(men_men_n486_), .Y(men_men_n805_));
  AOI210     u0777(.A0(men_men_n803_), .A1(men_men_n798_), .B0(men_men_n805_), .Y(men_men_n806_));
  NA3        u0778(.A(m), .B(l), .C(i), .Y(men_men_n807_));
  OAI220     u0779(.A0(men_men_n563_), .A1(men_men_n807_), .B0(men_men_n348_), .B1(men_men_n503_), .Y(men_men_n808_));
  NA2        u0780(.A(men_men_n774_), .B(men_men_n495_), .Y(men_men_n809_));
  OA210      u0781(.A0(men_men_n809_), .A1(men_men_n808_), .B0(men_men_n777_), .Y(men_men_n810_));
  INV        u0782(.A(men_men_n335_), .Y(men_men_n811_));
  NO2        u0783(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n812_));
  NA2        u0784(.A(men_men_n759_), .B(men_men_n330_), .Y(men_men_n813_));
  NA2        u0785(.A(men_men_n339_), .B(men_men_n341_), .Y(men_men_n814_));
  OAI210     u0786(.A0(men_men_n204_), .A1(men_men_n212_), .B0(men_men_n814_), .Y(men_men_n815_));
  NA2        u0787(.A(men_men_n815_), .B(men_men_n813_), .Y(men_men_n816_));
  INV        u0788(.A(men_men_n113_), .Y(men_men_n817_));
  NA2        u0789(.A(men_men_n817_), .B(men_men_n662_), .Y(men_men_n818_));
  NA3        u0790(.A(men_men_n818_), .B(men_men_n189_), .C(men_men_n31_), .Y(men_men_n819_));
  NA4        u0791(.A(men_men_n819_), .B(men_men_n816_), .C(men_men_n596_), .D(men_men_n80_), .Y(men_men_n820_));
  NO2        u0792(.A(men_men_n559_), .B(men_men_n471_), .Y(men_men_n821_));
  NOi21      u0793(.An(f), .B(d), .Y(men_men_n822_));
  NA2        u0794(.A(men_men_n822_), .B(m), .Y(men_men_n823_));
  NOi32      u0795(.An(g), .Bn(f), .C(d), .Y(men_men_n824_));
  NA4        u0796(.A(men_men_n824_), .B(men_men_n575_), .C(men_men_n29_), .D(m), .Y(men_men_n825_));
  INV        u0797(.A(men_men_n306_), .Y(men_men_n826_));
  AN2        u0798(.A(f), .B(d), .Y(men_men_n827_));
  NA3        u0799(.A(men_men_n452_), .B(men_men_n827_), .C(men_men_n82_), .Y(men_men_n828_));
  NO3        u0800(.A(men_men_n828_), .B(men_men_n71_), .C(men_men_n213_), .Y(men_men_n829_));
  NO2        u0801(.A(men_men_n283_), .B(men_men_n53_), .Y(men_men_n830_));
  NA2        u0802(.A(men_men_n826_), .B(men_men_n829_), .Y(men_men_n831_));
  NAi31      u0803(.An(men_men_n462_), .B(men_men_n831_), .C(men_men_n825_), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n626_), .B(men_men_n325_), .Y(men_men_n833_));
  AN2        u0805(.A(men_men_n833_), .B(men_men_n646_), .Y(men_men_n834_));
  NO2        u0806(.A(men_men_n834_), .B(men_men_n233_), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n573_), .B(men_men_n82_), .Y(men_men_n836_));
  NO2        u0808(.A(men_men_n814_), .B(men_men_n836_), .Y(men_men_n837_));
  NA3        u0809(.A(men_men_n161_), .B(men_men_n107_), .C(g), .Y(men_men_n838_));
  OAI220     u0810(.A0(men_men_n828_), .A1(men_men_n411_), .B0(men_men_n335_), .B1(men_men_n838_), .Y(men_men_n839_));
  NOi41      u0811(.An(men_men_n222_), .B(men_men_n839_), .C(men_men_n837_), .D(men_men_n301_), .Y(men_men_n840_));
  NA2        u0812(.A(c), .B(men_men_n115_), .Y(men_men_n841_));
  NO2        u0813(.A(men_men_n841_), .B(men_men_n390_), .Y(men_men_n842_));
  NA3        u0814(.A(men_men_n842_), .B(men_men_n484_), .C(f), .Y(men_men_n843_));
  OR2        u0815(.A(men_men_n633_), .B(men_men_n518_), .Y(men_men_n844_));
  INV        u0816(.A(men_men_n844_), .Y(men_men_n845_));
  NA2        u0817(.A(men_men_n776_), .B(men_men_n110_), .Y(men_men_n846_));
  NA2        u0818(.A(men_men_n846_), .B(men_men_n845_), .Y(men_men_n847_));
  NA4        u0819(.A(men_men_n847_), .B(men_men_n843_), .C(men_men_n840_), .D(men_men_n835_), .Y(men_men_n848_));
  NO4        u0820(.A(men_men_n848_), .B(men_men_n832_), .C(men_men_n820_), .D(men_men_n810_), .Y(men_men_n849_));
  OR2        u0821(.A(men_men_n828_), .B(men_men_n71_), .Y(men_men_n850_));
  NA2        u0822(.A(men_men_n800_), .B(g), .Y(men_men_n851_));
  AOI210     u0823(.A0(men_men_n851_), .A1(men_men_n291_), .B0(men_men_n850_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n135_), .B(men_men_n131_), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n229_), .B(men_men_n223_), .Y(men_men_n854_));
  AOI220     u0826(.A0(men_men_n854_), .A1(men_men_n226_), .B0(men_men_n300_), .B1(men_men_n853_), .Y(men_men_n855_));
  NO2        u0827(.A(men_men_n411_), .B(men_men_n799_), .Y(men_men_n856_));
  INV        u0828(.A(men_men_n855_), .Y(men_men_n857_));
  NA2        u0829(.A(e), .B(d), .Y(men_men_n858_));
  OAI220     u0830(.A0(men_men_n858_), .A1(c), .B0(men_men_n320_), .B1(d), .Y(men_men_n859_));
  NA3        u0831(.A(men_men_n859_), .B(men_men_n433_), .C(men_men_n482_), .Y(men_men_n860_));
  AOI210     u0832(.A0(men_men_n490_), .A1(men_men_n180_), .B0(men_men_n229_), .Y(men_men_n861_));
  AOI210     u0833(.A0(men_men_n595_), .A1(men_men_n343_), .B0(men_men_n861_), .Y(men_men_n862_));
  NA2        u0834(.A(men_men_n283_), .B(men_men_n166_), .Y(men_men_n863_));
  NA2        u0835(.A(men_men_n829_), .B(men_men_n863_), .Y(men_men_n864_));
  NA3        u0836(.A(men_men_n169_), .B(men_men_n83_), .C(men_men_n34_), .Y(men_men_n865_));
  NA4        u0837(.A(men_men_n865_), .B(men_men_n864_), .C(men_men_n862_), .D(men_men_n860_), .Y(men_men_n866_));
  NO3        u0838(.A(men_men_n866_), .B(men_men_n857_), .C(men_men_n852_), .Y(men_men_n867_));
  AO210      u0839(.A0(men_men_n335_), .A1(men_men_n664_), .B0(men_men_n216_), .Y(men_men_n868_));
  OAI220     u0840(.A0(men_men_n594_), .A1(men_men_n57_), .B0(men_men_n295_), .B1(j), .Y(men_men_n869_));
  AOI220     u0841(.A0(men_men_n869_), .A1(men_men_n833_), .B0(men_men_n584_), .B1(men_men_n593_), .Y(men_men_n870_));
  OAI210     u0842(.A0(men_men_n804_), .A1(men_men_n171_), .B0(men_men_n870_), .Y(men_men_n871_));
  AN2        u0843(.A(men_men_n813_), .B(men_men_n808_), .Y(men_men_n872_));
  NOi31      u0844(.An(men_men_n520_), .B(men_men_n823_), .C(men_men_n291_), .Y(men_men_n873_));
  NO3        u0845(.A(men_men_n873_), .B(men_men_n872_), .C(men_men_n871_), .Y(men_men_n874_));
  AO220      u0846(.A0(men_men_n433_), .A1(men_men_n713_), .B0(men_men_n176_), .B1(f), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n875_), .B(men_men_n859_), .Y(men_men_n876_));
  NO2        u0848(.A(men_men_n418_), .B(men_men_n67_), .Y(men_men_n877_));
  OAI210     u0849(.A0(men_men_n809_), .A1(men_men_n877_), .B0(men_men_n668_), .Y(men_men_n878_));
  AN4        u0850(.A(men_men_n878_), .B(men_men_n876_), .C(men_men_n874_), .D(men_men_n868_), .Y(men_men_n879_));
  NA4        u0851(.A(men_men_n879_), .B(men_men_n867_), .C(men_men_n849_), .D(men_men_n806_), .Y(men12));
  NO4        u0852(.A(men_men_n423_), .B(men_men_n253_), .C(men_men_n555_), .D(men_men_n213_), .Y(men_men_n881_));
  NA2        u0853(.A(men_men_n520_), .B(men_men_n877_), .Y(men_men_n882_));
  NO2        u0854(.A(men_men_n431_), .B(men_men_n115_), .Y(men_men_n883_));
  NO2        u0855(.A(men_men_n812_), .B(men_men_n348_), .Y(men_men_n884_));
  NO2        u0856(.A(men_men_n633_), .B(men_men_n367_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n884_), .B(men_men_n883_), .Y(men_men_n886_));
  NA3        u0858(.A(men_men_n886_), .B(men_men_n882_), .C(men_men_n422_), .Y(men_men_n887_));
  AOI210     u0859(.A0(men_men_n232_), .A1(men_men_n334_), .B0(men_men_n201_), .Y(men_men_n888_));
  OR2        u0860(.A(men_men_n888_), .B(men_men_n881_), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n889_), .B(men_men_n385_), .Y(men_men_n890_));
  NO2        u0862(.A(men_men_n612_), .B(men_men_n261_), .Y(men_men_n891_));
  NO2        u0863(.A(men_men_n563_), .B(men_men_n807_), .Y(men_men_n892_));
  AOI220     u0864(.A0(men_men_n892_), .A1(men_men_n542_), .B0(men_men_n787_), .B1(men_men_n891_), .Y(men_men_n893_));
  NO2        u0865(.A(men_men_n152_), .B(men_men_n236_), .Y(men_men_n894_));
  NA2        u0866(.A(men_men_n893_), .B(men_men_n890_), .Y(men_men_n895_));
  OR2        u0867(.A(men_men_n321_), .B(men_men_n883_), .Y(men_men_n896_));
  NA2        u0868(.A(men_men_n896_), .B(men_men_n349_), .Y(men_men_n897_));
  NA4        u0869(.A(men_men_n424_), .B(men_men_n416_), .C(men_men_n181_), .D(g), .Y(men_men_n898_));
  NA2        u0870(.A(men_men_n898_), .B(men_men_n897_), .Y(men_men_n899_));
  NO3        u0871(.A(men_men_n899_), .B(men_men_n895_), .C(men_men_n887_), .Y(men_men_n900_));
  NA2        u0872(.A(men_men_n529_), .B(men_men_n145_), .Y(men_men_n901_));
  NOi21      u0873(.An(men_men_n34_), .B(men_men_n626_), .Y(men_men_n902_));
  NA2        u0874(.A(men_men_n902_), .B(men_men_n901_), .Y(men_men_n903_));
  OAI210     u0875(.A0(men_men_n251_), .A1(men_men_n45_), .B0(men_men_n903_), .Y(men_men_n904_));
  NA2        u0876(.A(men_men_n414_), .B(men_men_n263_), .Y(men_men_n905_));
  NO3        u0877(.A(men_men_n789_), .B(men_men_n87_), .C(men_men_n390_), .Y(men_men_n906_));
  NAi31      u0878(.An(men_men_n906_), .B(men_men_n905_), .C(men_men_n317_), .Y(men_men_n907_));
  NO2        u0879(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n908_));
  NO2        u0880(.A(men_men_n478_), .B(men_men_n295_), .Y(men_men_n909_));
  INV        u0881(.A(men_men_n909_), .Y(men_men_n910_));
  NO2        u0882(.A(men_men_n910_), .B(men_men_n145_), .Y(men_men_n911_));
  NA2        u0883(.A(men_men_n605_), .B(j), .Y(men_men_n912_));
  INV        u0884(.A(men_men_n356_), .Y(men_men_n913_));
  NO4        u0885(.A(men_men_n913_), .B(men_men_n911_), .C(men_men_n907_), .D(men_men_n904_), .Y(men_men_n914_));
  NA2        u0886(.A(men_men_n343_), .B(g), .Y(men_men_n915_));
  NA2        u0887(.A(men_men_n164_), .B(i), .Y(men_men_n916_));
  NA2        u0888(.A(men_men_n46_), .B(i), .Y(men_men_n917_));
  OAI220     u0889(.A0(men_men_n917_), .A1(men_men_n200_), .B0(men_men_n916_), .B1(men_men_n90_), .Y(men_men_n918_));
  AOI210     u0890(.A0(men_men_n401_), .A1(men_men_n37_), .B0(men_men_n918_), .Y(men_men_n919_));
  INV        u0891(.A(men_men_n145_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n529_), .B(men_men_n371_), .Y(men_men_n921_));
  NA2        u0893(.A(men_men_n921_), .B(n), .Y(men_men_n922_));
  OAI220     u0894(.A0(men_men_n922_), .A1(men_men_n915_), .B0(men_men_n919_), .B1(men_men_n330_), .Y(men_men_n923_));
  NO2        u0895(.A(men_men_n633_), .B(men_men_n471_), .Y(men_men_n924_));
  NA3        u0896(.A(men_men_n339_), .B(men_men_n600_), .C(i), .Y(men_men_n925_));
  OAI210     u0897(.A0(men_men_n418_), .A1(men_men_n306_), .B0(men_men_n925_), .Y(men_men_n926_));
  OAI220     u0898(.A0(men_men_n926_), .A1(men_men_n924_), .B0(men_men_n644_), .B1(men_men_n725_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n578_), .B(men_men_n112_), .Y(men_men_n928_));
  OR3        u0900(.A(men_men_n306_), .B(men_men_n413_), .C(f), .Y(men_men_n929_));
  NA3        u0901(.A(men_men_n600_), .B(men_men_n78_), .C(i), .Y(men_men_n930_));
  OA220      u0902(.A0(men_men_n930_), .A1(men_men_n928_), .B0(men_men_n929_), .B1(men_men_n562_), .Y(men_men_n931_));
  NA3        u0903(.A(men_men_n322_), .B(men_men_n117_), .C(g), .Y(men_men_n932_));
  AOI210     u0904(.A0(men_men_n643_), .A1(men_men_n932_), .B0(m), .Y(men_men_n933_));
  OAI210     u0905(.A0(men_men_n933_), .A1(men_men_n884_), .B0(men_men_n321_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n930_), .B(men_men_n929_), .Y(men_men_n935_));
  NA2        u0907(.A(men_men_n935_), .B(men_men_n259_), .Y(men_men_n936_));
  NA4        u0908(.A(men_men_n936_), .B(men_men_n934_), .C(men_men_n931_), .D(men_men_n927_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n367_), .B(men_men_n89_), .Y(men_men_n938_));
  OAI210     u0910(.A0(men_men_n938_), .A1(men_men_n891_), .B0(men_men_n237_), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n437_), .B(men_men_n213_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n896_), .B(men_men_n217_), .Y(men_men_n941_));
  AOI220     u0913(.A0(men_men_n885_), .A1(men_men_n894_), .B0(men_men_n561_), .B1(men_men_n88_), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n942_), .B(men_men_n941_), .C(men_men_n939_), .Y(men_men_n943_));
  AOI210     u0915(.A0(men_men_n402_), .A1(men_men_n394_), .B0(men_men_n789_), .Y(men_men_n944_));
  INV        u0916(.A(men_men_n108_), .Y(men_men_n945_));
  AOI210     u0917(.A0(men_men_n945_), .A1(men_men_n512_), .B0(men_men_n944_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n933_), .B(men_men_n883_), .Y(men_men_n947_));
  NA2        u0919(.A(men_men_n617_), .B(men_men_n507_), .Y(men_men_n948_));
  NA3        u0920(.A(men_men_n948_), .B(men_men_n947_), .C(men_men_n946_), .Y(men_men_n949_));
  NO4        u0921(.A(men_men_n949_), .B(men_men_n943_), .C(men_men_n937_), .D(men_men_n923_), .Y(men_men_n950_));
  NAi31      u0922(.An(men_men_n141_), .B(men_men_n403_), .C(n), .Y(men_men_n951_));
  NO3        u0923(.A(men_men_n271_), .B(men_men_n141_), .C(men_men_n390_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n472_), .Y(men_men_n953_));
  INV        u0925(.A(men_men_n953_), .Y(men_men_n954_));
  NA2        u0926(.A(men_men_n229_), .B(men_men_n172_), .Y(men_men_n955_));
  NO2        u0927(.A(men_men_n424_), .B(men_men_n176_), .Y(men_men_n956_));
  NOi31      u0928(.An(men_men_n955_), .B(men_men_n956_), .C(men_men_n213_), .Y(men_men_n957_));
  NAi21      u0929(.An(men_men_n529_), .B(men_men_n940_), .Y(men_men_n958_));
  NO3        u0930(.A(men_men_n418_), .B(men_men_n306_), .C(men_men_n71_), .Y(men_men_n959_));
  AOI220     u0931(.A0(men_men_n959_), .A1(men_men_n415_), .B0(men_men_n456_), .B1(g), .Y(men_men_n960_));
  NA2        u0932(.A(men_men_n960_), .B(men_men_n958_), .Y(men_men_n961_));
  NO2        u0933(.A(men_men_n951_), .B(men_men_n232_), .Y(men_men_n962_));
  NO3        u0934(.A(n), .B(men_men_n150_), .C(men_men_n212_), .Y(men_men_n963_));
  OAI210     u0935(.A0(men_men_n963_), .A1(men_men_n501_), .B0(men_men_n368_), .Y(men_men_n964_));
  NA2        u0936(.A(men_men_n964_), .B(men_men_n592_), .Y(men_men_n965_));
  OAI210     u0937(.A0(men_men_n888_), .A1(men_men_n881_), .B0(men_men_n955_), .Y(men_men_n966_));
  NA3        u0938(.A(men_men_n921_), .B(men_men_n460_), .C(men_men_n46_), .Y(men_men_n967_));
  AOI210     u0939(.A0(men_men_n370_), .A1(men_men_n368_), .B0(men_men_n329_), .Y(men_men_n968_));
  NA4        u0940(.A(men_men_n968_), .B(men_men_n967_), .C(men_men_n966_), .D(men_men_n272_), .Y(men_men_n969_));
  OR3        u0941(.A(men_men_n969_), .B(men_men_n965_), .C(men_men_n962_), .Y(men_men_n970_));
  NO4        u0942(.A(men_men_n970_), .B(men_men_n961_), .C(men_men_n957_), .D(men_men_n954_), .Y(men_men_n971_));
  NA4        u0943(.A(men_men_n971_), .B(men_men_n950_), .C(men_men_n914_), .D(men_men_n900_), .Y(men13));
  AN2        u0944(.A(c), .B(b), .Y(men_men_n973_));
  NA3        u0945(.A(men_men_n250_), .B(men_men_n973_), .C(m), .Y(men_men_n974_));
  NA2        u0946(.A(men_men_n469_), .B(f), .Y(men_men_n975_));
  NO4        u0947(.A(men_men_n975_), .B(men_men_n974_), .C(j), .D(men_men_n556_), .Y(men_men_n976_));
  INV        u0948(.A(men_men_n263_), .Y(men_men_n977_));
  NO4        u0949(.A(men_men_n977_), .B(men_men_n975_), .C(men_men_n916_), .D(a), .Y(men_men_n978_));
  NAi32      u0950(.An(d), .Bn(c), .C(e), .Y(men_men_n979_));
  NA2        u0951(.A(men_men_n140_), .B(men_men_n45_), .Y(men_men_n980_));
  NO4        u0952(.A(men_men_n980_), .B(men_men_n979_), .C(men_men_n563_), .D(men_men_n302_), .Y(men_men_n981_));
  NA2        u0953(.A(men_men_n393_), .B(men_men_n212_), .Y(men_men_n982_));
  AN2        u0954(.A(d), .B(c), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n983_), .B(men_men_n115_), .Y(men_men_n984_));
  NO3        u0956(.A(men_men_n984_), .B(men_men_n982_), .C(men_men_n177_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n469_), .B(c), .Y(men_men_n986_));
  NO4        u0958(.A(men_men_n980_), .B(men_men_n559_), .C(men_men_n986_), .D(men_men_n302_), .Y(men_men_n987_));
  OR2        u0959(.A(men_men_n985_), .B(men_men_n987_), .Y(men_men_n988_));
  OR4        u0960(.A(men_men_n988_), .B(men_men_n981_), .C(men_men_n978_), .D(men_men_n976_), .Y(men_men_n989_));
  NAi32      u0961(.An(f), .Bn(e), .C(c), .Y(men_men_n990_));
  NO2        u0962(.A(men_men_n990_), .B(men_men_n147_), .Y(men_men_n991_));
  NA2        u0963(.A(men_men_n991_), .B(g), .Y(men_men_n992_));
  OR2        u0964(.A(men_men_n223_), .B(men_men_n177_), .Y(men_men_n993_));
  NO2        u0965(.A(men_men_n993_), .B(men_men_n992_), .Y(men_men_n994_));
  NO2        u0966(.A(men_men_n986_), .B(men_men_n302_), .Y(men_men_n995_));
  NO2        u0967(.A(j), .B(men_men_n45_), .Y(men_men_n996_));
  NA2        u0968(.A(men_men_n602_), .B(men_men_n996_), .Y(men_men_n997_));
  NOi21      u0969(.An(men_men_n995_), .B(men_men_n997_), .Y(men_men_n998_));
  NOi41      u0970(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n999_));
  NA2        u0971(.A(men_men_n999_), .B(l), .Y(men_men_n1000_));
  NO2        u0972(.A(men_men_n1000_), .B(men_men_n992_), .Y(men_men_n1001_));
  OR3        u0973(.A(e), .B(d), .C(c), .Y(men_men_n1002_));
  NA3        u0974(.A(k), .B(j), .C(i), .Y(men_men_n1003_));
  NO3        u0975(.A(men_men_n1003_), .B(men_men_n302_), .C(men_men_n89_), .Y(men_men_n1004_));
  BUFFER     u0976(.A(men_men_n1004_), .Y(men_men_n1005_));
  OR4        u0977(.A(men_men_n1005_), .B(men_men_n1001_), .C(men_men_n998_), .D(men_men_n994_), .Y(men_men_n1006_));
  NA3        u0978(.A(men_men_n444_), .B(men_men_n332_), .C(men_men_n53_), .Y(men_men_n1007_));
  NO2        u0979(.A(men_men_n1007_), .B(men_men_n997_), .Y(men_men_n1008_));
  NO4        u0980(.A(men_men_n1007_), .B(men_men_n559_), .C(men_men_n430_), .D(men_men_n45_), .Y(men_men_n1009_));
  NO2        u0981(.A(f), .B(c), .Y(men_men_n1010_));
  NOi21      u0982(.An(men_men_n1010_), .B(men_men_n423_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n1011_), .B(men_men_n56_), .Y(men_men_n1012_));
  NO3        u0984(.A(i), .B(men_men_n243_), .C(l), .Y(men_men_n1013_));
  NOi31      u0985(.An(men_men_n1013_), .B(men_men_n1012_), .C(j), .Y(men_men_n1014_));
  OR3        u0986(.A(men_men_n1014_), .B(men_men_n1009_), .C(men_men_n1008_), .Y(men_men_n1015_));
  OR3        u0987(.A(men_men_n1015_), .B(men_men_n1006_), .C(men_men_n989_), .Y(men02));
  OR3        u0988(.A(h), .B(g), .C(f), .Y(men_men_n1017_));
  OR3        u0989(.A(n), .B(m), .C(i), .Y(men_men_n1018_));
  NO4        u0990(.A(men_men_n1018_), .B(men_men_n1017_), .C(l), .D(men_men_n1002_), .Y(men_men_n1019_));
  NO2        u0991(.A(men_men_n1004_), .B(men_men_n981_), .Y(men_men_n1020_));
  AN3        u0992(.A(g), .B(f), .C(c), .Y(men_men_n1021_));
  NA3        u0993(.A(men_men_n1021_), .B(men_men_n444_), .C(h), .Y(men_men_n1022_));
  BUFFER     u0994(.A(men_men_n302_), .Y(men_men_n1023_));
  OR2        u0995(.A(men_men_n1023_), .B(men_men_n1022_), .Y(men_men_n1024_));
  NO3        u0996(.A(men_men_n1007_), .B(men_men_n980_), .C(men_men_n559_), .Y(men_men_n1025_));
  NO2        u0997(.A(men_men_n1025_), .B(men_men_n994_), .Y(men_men_n1026_));
  NA2        u0998(.A(i), .B(h), .Y(men_men_n1027_));
  NO2        u0999(.A(men_men_n1027_), .B(men_men_n131_), .Y(men_men_n1028_));
  NO3        u1000(.A(men_men_n142_), .B(men_men_n281_), .C(men_men_n213_), .Y(men_men_n1029_));
  AOI210     u1001(.A0(men_men_n1029_), .A1(men_men_n1028_), .B0(men_men_n998_), .Y(men_men_n1030_));
  NA3        u1002(.A(c), .B(b), .C(a), .Y(men_men_n1031_));
  NO3        u1003(.A(men_men_n1031_), .B(men_men_n858_), .C(men_men_n212_), .Y(men_men_n1032_));
  NO3        u1004(.A(men_men_n1003_), .B(men_men_n49_), .C(men_men_n111_), .Y(men_men_n1033_));
  AOI210     u1005(.A0(men_men_n1033_), .A1(men_men_n1032_), .B0(men_men_n1008_), .Y(men_men_n1034_));
  AN4        u1006(.A(men_men_n1034_), .B(men_men_n1030_), .C(men_men_n1026_), .D(men_men_n1024_), .Y(men_men_n1035_));
  NO2        u1007(.A(men_men_n984_), .B(men_men_n982_), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n1000_), .B(men_men_n993_), .Y(men_men_n1037_));
  AOI210     u1009(.A0(men_men_n1037_), .A1(men_men_n1036_), .B0(men_men_n976_), .Y(men_men_n1038_));
  NAi41      u1010(.An(men_men_n1019_), .B(men_men_n1038_), .C(men_men_n1035_), .D(men_men_n1020_), .Y(men03));
  NO2        u1011(.A(men_men_n503_), .B(men_men_n569_), .Y(men_men_n1040_));
  NA4        u1012(.A(men_men_n86_), .B(men_men_n85_), .C(g), .D(men_men_n212_), .Y(men_men_n1041_));
  INV        u1013(.A(men_men_n1041_), .Y(men_men_n1042_));
  NO3        u1014(.A(men_men_n1042_), .B(men_men_n1040_), .C(men_men_n945_), .Y(men_men_n1043_));
  NOi41      u1015(.An(men_men_n774_), .B(men_men_n815_), .C(men_men_n808_), .D(men_men_n681_), .Y(men_men_n1044_));
  OAI220     u1016(.A0(men_men_n1044_), .A1(men_men_n655_), .B0(men_men_n1043_), .B1(men_men_n560_), .Y(men_men_n1045_));
  NOi31      u1017(.An(i), .B(k), .C(j), .Y(men_men_n1046_));
  NA4        u1018(.A(men_men_n1046_), .B(e), .C(men_men_n339_), .D(men_men_n332_), .Y(men_men_n1047_));
  OAI210     u1019(.A0(men_men_n789_), .A1(men_men_n404_), .B0(men_men_n1047_), .Y(men_men_n1048_));
  NOi31      u1020(.An(m), .B(n), .C(f), .Y(men_men_n1049_));
  NA2        u1021(.A(men_men_n1049_), .B(men_men_n51_), .Y(men_men_n1050_));
  AN2        u1022(.A(e), .B(c), .Y(men_men_n1051_));
  NA2        u1023(.A(men_men_n1051_), .B(a), .Y(men_men_n1052_));
  OAI220     u1024(.A0(men_men_n1052_), .A1(men_men_n1050_), .B0(men_men_n844_), .B1(men_men_n409_), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n482_), .B(l), .Y(men_men_n1054_));
  NOi31      u1026(.An(men_men_n824_), .B(men_men_n974_), .C(men_men_n1054_), .Y(men_men_n1055_));
  NO3        u1027(.A(men_men_n1055_), .B(men_men_n1053_), .C(men_men_n1048_), .Y(men_men_n1056_));
  NO2        u1028(.A(men_men_n281_), .B(a), .Y(men_men_n1057_));
  INV        u1029(.A(men_men_n981_), .Y(men_men_n1058_));
  NO2        u1030(.A(men_men_n1027_), .B(men_men_n459_), .Y(men_men_n1059_));
  NO2        u1031(.A(men_men_n85_), .B(g), .Y(men_men_n1060_));
  AOI210     u1032(.A0(men_men_n1060_), .A1(men_men_n1059_), .B0(men_men_n1013_), .Y(men_men_n1061_));
  OR2        u1033(.A(men_men_n1061_), .B(men_men_n1012_), .Y(men_men_n1062_));
  NA3        u1034(.A(men_men_n1062_), .B(men_men_n1058_), .C(men_men_n1056_), .Y(men_men_n1063_));
  NO4        u1035(.A(men_men_n1063_), .B(men_men_n1045_), .C(men_men_n791_), .D(men_men_n541_), .Y(men_men_n1064_));
  NA2        u1036(.A(c), .B(b), .Y(men_men_n1065_));
  NO2        u1037(.A(men_men_n667_), .B(men_men_n1065_), .Y(men_men_n1066_));
  OAI210     u1038(.A0(men_men_n823_), .A1(men_men_n802_), .B0(men_men_n397_), .Y(men_men_n1067_));
  NA2        u1039(.A(men_men_n1067_), .B(men_men_n1066_), .Y(men_men_n1068_));
  NAi21      u1040(.An(men_men_n405_), .B(men_men_n1066_), .Y(men_men_n1069_));
  OAI210     u1041(.A0(men_men_n523_), .A1(men_men_n39_), .B0(men_men_n1057_), .Y(men_men_n1070_));
  NA2        u1042(.A(men_men_n1070_), .B(men_men_n1069_), .Y(men_men_n1071_));
  INV        u1043(.A(men_men_n118_), .Y(men_men_n1072_));
  OAI210     u1044(.A0(men_men_n1072_), .A1(men_men_n285_), .B0(g), .Y(men_men_n1073_));
  NO2        u1045(.A(f), .B(men_men_n1031_), .Y(men_men_n1074_));
  NO2        u1046(.A(men_men_n1073_), .B(men_men_n1031_), .Y(men_men_n1075_));
  AOI210     u1047(.A0(men_men_n1075_), .A1(men_men_n112_), .B0(men_men_n1071_), .Y(men_men_n1076_));
  NA2        u1048(.A(men_men_n447_), .B(men_men_n446_), .Y(men_men_n1077_));
  NO2        u1049(.A(men_men_n182_), .B(men_men_n236_), .Y(men_men_n1078_));
  NA2        u1050(.A(men_men_n1078_), .B(m), .Y(men_men_n1079_));
  NA2        u1051(.A(men_men_n1054_), .B(men_men_n166_), .Y(men_men_n1080_));
  NA2        u1052(.A(men_men_n1080_), .B(men_men_n448_), .Y(men_men_n1081_));
  AOI210     u1053(.A0(men_men_n1081_), .A1(men_men_n1077_), .B0(men_men_n1079_), .Y(men_men_n1082_));
  NA2        u1054(.A(men_men_n536_), .B(men_men_n392_), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n160_), .B(men_men_n33_), .Y(men_men_n1084_));
  AOI210     u1056(.A0(men_men_n912_), .A1(men_men_n1084_), .B0(men_men_n213_), .Y(men_men_n1085_));
  OAI210     u1057(.A0(men_men_n1085_), .A1(men_men_n427_), .B0(men_men_n1074_), .Y(men_men_n1086_));
  INV        u1058(.A(men_men_n906_), .Y(men_men_n1087_));
  NA3        u1059(.A(men_men_n1087_), .B(men_men_n1086_), .C(men_men_n1083_), .Y(men_men_n1088_));
  NO2        u1060(.A(men_men_n1088_), .B(men_men_n1082_), .Y(men_men_n1089_));
  NA4        u1061(.A(men_men_n1089_), .B(men_men_n1076_), .C(men_men_n1068_), .D(men_men_n1064_), .Y(men00));
  AOI210     u1062(.A0(men_men_n856_), .A1(men_men_n894_), .B0(men_men_n1048_), .Y(men_men_n1091_));
  NO3        u1063(.A(men_men_n1025_), .B(men_men_n906_), .C(men_men_n678_), .Y(men_men_n1092_));
  NA3        u1064(.A(men_men_n1092_), .B(men_men_n1091_), .C(men_men_n946_), .Y(men_men_n1093_));
  NA2        u1065(.A(men_men_n484_), .B(f), .Y(men_men_n1094_));
  INV        u1066(.A(men_men_n619_), .Y(men_men_n1095_));
  NA3        u1067(.A(men_men_n1095_), .B(men_men_n258_), .C(n), .Y(men_men_n1096_));
  AOI210     u1068(.A0(men_men_n1096_), .A1(men_men_n1094_), .B0(men_men_n984_), .Y(men_men_n1097_));
  NO3        u1069(.A(men_men_n1097_), .B(men_men_n1093_), .C(men_men_n1006_), .Y(men_men_n1098_));
  NA3        u1070(.A(men_men_n169_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1099_));
  NA3        u1071(.A(d), .B(men_men_n53_), .C(b), .Y(men_men_n1100_));
  NO2        u1072(.A(men_men_n1100_), .B(men_men_n1099_), .Y(men_men_n1101_));
  NO2        u1073(.A(men_men_n1101_), .B(men_men_n873_), .Y(men_men_n1102_));
  NO4        u1074(.A(men_men_n1419_), .B(men_men_n350_), .C(men_men_n1065_), .D(men_men_n56_), .Y(men_men_n1103_));
  OR2        u1075(.A(men_men_n374_), .B(men_men_n134_), .Y(men_men_n1104_));
  NO2        u1076(.A(h), .B(g), .Y(men_men_n1105_));
  NA4        u1077(.A(men_men_n472_), .B(men_men_n444_), .C(men_men_n1105_), .D(men_men_n973_), .Y(men_men_n1106_));
  OAI220     u1078(.A0(men_men_n503_), .A1(men_men_n569_), .B0(men_men_n90_), .B1(men_men_n89_), .Y(men_men_n1107_));
  NA2        u1079(.A(men_men_n1107_), .B(men_men_n512_), .Y(men_men_n1108_));
  NA2        u1080(.A(men_men_n314_), .B(men_men_n247_), .Y(men_men_n1109_));
  NA4        u1081(.A(men_men_n1109_), .B(men_men_n1108_), .C(men_men_n1106_), .D(men_men_n1104_), .Y(men_men_n1110_));
  NO3        u1082(.A(men_men_n1110_), .B(men_men_n1103_), .C(men_men_n265_), .Y(men_men_n1111_));
  INV        u1083(.A(men_men_n319_), .Y(men_men_n1112_));
  AOI210     u1084(.A0(men_men_n247_), .A1(men_men_n343_), .B0(men_men_n552_), .Y(men_men_n1113_));
  NA3        u1085(.A(men_men_n1113_), .B(men_men_n1112_), .C(men_men_n155_), .Y(men_men_n1114_));
  NO2        u1086(.A(men_men_n238_), .B(men_men_n181_), .Y(men_men_n1115_));
  NA2        u1087(.A(men_men_n1115_), .B(men_men_n410_), .Y(men_men_n1116_));
  NA3        u1088(.A(men_men_n179_), .B(men_men_n111_), .C(g), .Y(men_men_n1117_));
  NA2        u1089(.A(men_men_n444_), .B(f), .Y(men_men_n1118_));
  NOi31      u1090(.An(men_men_n830_), .B(men_men_n1118_), .C(men_men_n1117_), .Y(men_men_n1119_));
  NAi31      u1091(.An(men_men_n185_), .B(men_men_n821_), .C(men_men_n444_), .Y(men_men_n1120_));
  NAi31      u1092(.An(men_men_n1119_), .B(men_men_n1120_), .C(men_men_n1116_), .Y(men_men_n1121_));
  NO2        u1093(.A(men_men_n273_), .B(men_men_n71_), .Y(men_men_n1122_));
  NO3        u1094(.A(men_men_n409_), .B(men_men_n799_), .C(n), .Y(men_men_n1123_));
  AOI210     u1095(.A0(men_men_n1123_), .A1(men_men_n1122_), .B0(men_men_n1019_), .Y(men_men_n1124_));
  NAi31      u1096(.An(men_men_n987_), .B(men_men_n1124_), .C(men_men_n70_), .Y(men_men_n1125_));
  NO4        u1097(.A(men_men_n1125_), .B(men_men_n1121_), .C(men_men_n1114_), .D(men_men_n494_), .Y(men_men_n1126_));
  AN3        u1098(.A(men_men_n1126_), .B(men_men_n1111_), .C(men_men_n1102_), .Y(men_men_n1127_));
  NA2        u1099(.A(men_men_n512_), .B(men_men_n100_), .Y(men_men_n1128_));
  NA3        u1100(.A(men_men_n1049_), .B(men_men_n578_), .C(men_men_n443_), .Y(men_men_n1129_));
  NA4        u1101(.A(men_men_n1129_), .B(men_men_n537_), .C(men_men_n1128_), .D(men_men_n241_), .Y(men_men_n1130_));
  NA2        u1102(.A(men_men_n1042_), .B(men_men_n512_), .Y(men_men_n1131_));
  NA4        u1103(.A(men_men_n622_), .B(k), .C(men_men_n219_), .D(men_men_n164_), .Y(men_men_n1132_));
  NA2        u1104(.A(men_men_n1132_), .B(men_men_n1131_), .Y(men_men_n1133_));
  OAI210     u1105(.A0(men_men_n442_), .A1(men_men_n119_), .B0(men_men_n825_), .Y(men_men_n1134_));
  AOI220     u1106(.A0(men_men_n1134_), .A1(men_men_n1080_), .B0(men_men_n536_), .B1(men_men_n392_), .Y(men_men_n1135_));
  OR3        u1107(.A(men_men_n984_), .B(men_men_n271_), .C(men_men_n221_), .Y(men_men_n1136_));
  INV        u1108(.A(men_men_n216_), .Y(men_men_n1137_));
  NA2        u1109(.A(men_men_n811_), .B(men_men_n1137_), .Y(men_men_n1138_));
  OAI210     u1110(.A0(men_men_n351_), .A1(men_men_n308_), .B0(men_men_n429_), .Y(men_men_n1139_));
  NA4        u1111(.A(men_men_n1139_), .B(men_men_n1138_), .C(men_men_n1136_), .D(men_men_n1135_), .Y(men_men_n1140_));
  INV        u1112(.A(men_men_n790_), .Y(men_men_n1141_));
  AOI220     u1113(.A0(men_men_n902_), .A1(men_men_n550_), .B0(men_men_n622_), .B1(men_men_n244_), .Y(men_men_n1142_));
  NO2        u1114(.A(men_men_n64_), .B(h), .Y(men_men_n1143_));
  NO3        u1115(.A(men_men_n984_), .B(men_men_n982_), .C(men_men_n694_), .Y(men_men_n1144_));
  OAI210     u1116(.A0(men_men_n1029_), .A1(men_men_n1144_), .B0(men_men_n1143_), .Y(men_men_n1145_));
  NA4        u1117(.A(men_men_n1145_), .B(men_men_n1142_), .C(men_men_n1141_), .D(men_men_n825_), .Y(men_men_n1146_));
  NO4        u1118(.A(men_men_n1146_), .B(men_men_n1140_), .C(men_men_n1133_), .D(men_men_n1130_), .Y(men_men_n1147_));
  NA2        u1119(.A(men_men_n803_), .B(men_men_n724_), .Y(men_men_n1148_));
  NA4        u1120(.A(men_men_n1148_), .B(men_men_n1147_), .C(men_men_n1127_), .D(men_men_n1098_), .Y(men01));
  NO3        u1121(.A(men_men_n770_), .B(men_men_n762_), .C(men_men_n279_), .Y(men_men_n1150_));
  NA2        u1122(.A(men_men_n1150_), .B(men_men_n964_), .Y(men_men_n1151_));
  NA2        u1123(.A(men_men_n561_), .B(men_men_n88_), .Y(men_men_n1152_));
  NA2        u1124(.A(men_men_n529_), .B(men_men_n270_), .Y(men_men_n1153_));
  NA2        u1125(.A(men_men_n909_), .B(men_men_n1153_), .Y(men_men_n1154_));
  NA4        u1126(.A(men_men_n1154_), .B(men_men_n1152_), .C(men_men_n870_), .D(men_men_n331_), .Y(men_men_n1155_));
  NA2        u1127(.A(men_men_n673_), .B(men_men_n95_), .Y(men_men_n1156_));
  NO2        u1128(.A(men_men_n1156_), .B(i), .Y(men_men_n1157_));
  OAI210     u1129(.A0(men_men_n748_), .A1(men_men_n574_), .B0(men_men_n1132_), .Y(men_men_n1158_));
  AOI210     u1130(.A0(men_men_n1157_), .A1(men_men_n607_), .B0(men_men_n1158_), .Y(men_men_n1159_));
  INV        u1131(.A(men_men_n117_), .Y(men_men_n1160_));
  OR2        u1132(.A(men_men_n1160_), .B(men_men_n558_), .Y(men_men_n1161_));
  NAi41      u1133(.An(men_men_n163_), .B(men_men_n1161_), .C(men_men_n1159_), .D(men_men_n855_), .Y(men_men_n1162_));
  NO2        u1134(.A(men_men_n749_), .B(men_men_n487_), .Y(men_men_n1163_));
  NA4        u1135(.A(men_men_n673_), .B(men_men_n95_), .C(men_men_n45_), .D(men_men_n212_), .Y(men_men_n1164_));
  OA220      u1136(.A0(men_men_n1164_), .A1(men_men_n69_), .B0(men_men_n195_), .B1(men_men_n193_), .Y(men_men_n1165_));
  NA3        u1137(.A(men_men_n1165_), .B(men_men_n1163_), .C(men_men_n137_), .Y(men_men_n1166_));
  NO4        u1138(.A(men_men_n1166_), .B(men_men_n1162_), .C(men_men_n1155_), .D(men_men_n1151_), .Y(men_men_n1167_));
  NA2        u1139(.A(men_men_n297_), .B(men_men_n507_), .Y(men_men_n1168_));
  NA2        u1140(.A(men_men_n515_), .B(men_men_n382_), .Y(men_men_n1169_));
  BUFFER     u1141(.A(men_men_n538_), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n1170_), .B(men_men_n1169_), .Y(men_men_n1171_));
  AN3        u1143(.A(m), .B(l), .C(k), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n352_), .A1(men_men_n34_), .B0(men_men_n1172_), .Y(men_men_n1173_));
  NA2        u1145(.A(men_men_n203_), .B(men_men_n34_), .Y(men_men_n1174_));
  AO210      u1146(.A0(men_men_n1174_), .A1(men_men_n1173_), .B0(men_men_n330_), .Y(men_men_n1175_));
  NA3        u1147(.A(men_men_n1175_), .B(men_men_n1171_), .C(men_men_n1168_), .Y(men_men_n1176_));
  INV        u1148(.A(men_men_n572_), .Y(men_men_n1177_));
  OAI210     u1149(.A0(men_men_n1160_), .A1(men_men_n567_), .B0(men_men_n1177_), .Y(men_men_n1178_));
  NO3        u1150(.A(men_men_n789_), .B(men_men_n204_), .C(men_men_n390_), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n1179_), .B(men_men_n906_), .Y(men_men_n1180_));
  NA2        u1152(.A(men_men_n1180_), .B(men_men_n752_), .Y(men_men_n1181_));
  NO3        u1153(.A(men_men_n1181_), .B(men_men_n1178_), .C(men_men_n1176_), .Y(men_men_n1182_));
  NA3        u1154(.A(men_men_n575_), .B(men_men_n29_), .C(f), .Y(men_men_n1183_));
  NO2        u1155(.A(men_men_n1183_), .B(men_men_n204_), .Y(men_men_n1184_));
  AOI210     u1156(.A0(men_men_n479_), .A1(men_men_n55_), .B0(men_men_n1184_), .Y(men_men_n1185_));
  NO2        u1157(.A(men_men_n1164_), .B(men_men_n928_), .Y(men_men_n1186_));
  NO2        u1158(.A(men_men_n1186_), .B(men_men_n1101_), .Y(men_men_n1187_));
  NA3        u1159(.A(men_men_n1187_), .B(men_men_n1185_), .C(men_men_n723_), .Y(men_men_n1188_));
  NO2        u1160(.A(men_men_n916_), .B(men_men_n231_), .Y(men_men_n1189_));
  NO2        u1161(.A(men_men_n917_), .B(men_men_n531_), .Y(men_men_n1190_));
  OAI210     u1162(.A0(men_men_n1190_), .A1(men_men_n1189_), .B0(men_men_n337_), .Y(men_men_n1191_));
  NA2        u1163(.A(men_men_n546_), .B(men_men_n544_), .Y(men_men_n1192_));
  NO3        u1164(.A(men_men_n77_), .B(men_men_n295_), .C(men_men_n45_), .Y(men_men_n1193_));
  NA2        u1165(.A(men_men_n1193_), .B(men_men_n528_), .Y(men_men_n1194_));
  NA3        u1166(.A(men_men_n1194_), .B(men_men_n1192_), .C(men_men_n640_), .Y(men_men_n1195_));
  NA2        u1167(.A(men_men_n1193_), .B(men_men_n780_), .Y(men_men_n1196_));
  NA2        u1168(.A(men_men_n1196_), .B(men_men_n376_), .Y(men_men_n1197_));
  NOi41      u1169(.An(men_men_n1191_), .B(men_men_n1197_), .C(men_men_n1195_), .D(men_men_n1188_), .Y(men_men_n1198_));
  NO2        u1170(.A(men_men_n130_), .B(men_men_n45_), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1200_));
  AO220      u1172(.A0(men_men_n1200_), .A1(men_men_n595_), .B0(men_men_n1199_), .B1(men_men_n671_), .Y(men_men_n1201_));
  NA2        u1173(.A(men_men_n1201_), .B(men_men_n337_), .Y(men_men_n1202_));
  INV        u1174(.A(men_men_n134_), .Y(men_men_n1203_));
  NO3        u1175(.A(men_men_n1027_), .B(men_men_n177_), .C(men_men_n85_), .Y(men_men_n1204_));
  AOI220     u1176(.A0(men_men_n1204_), .A1(men_men_n1203_), .B0(men_men_n1193_), .B1(men_men_n920_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n1205_), .B(men_men_n1202_), .Y(men_men_n1206_));
  NO2        u1178(.A(men_men_n586_), .B(men_men_n585_), .Y(men_men_n1207_));
  NO4        u1179(.A(men_men_n1027_), .B(men_men_n1207_), .C(men_men_n175_), .D(men_men_n85_), .Y(men_men_n1208_));
  NO3        u1180(.A(men_men_n1208_), .B(men_men_n1206_), .C(men_men_n611_), .Y(men_men_n1209_));
  NA4        u1181(.A(men_men_n1209_), .B(men_men_n1198_), .C(men_men_n1182_), .D(men_men_n1167_), .Y(men06));
  NO2        u1182(.A(men_men_n391_), .B(men_men_n535_), .Y(men_men_n1211_));
  NA2        u1183(.A(men_men_n266_), .B(men_men_n1211_), .Y(men_men_n1212_));
  NA2        u1184(.A(men_men_n1212_), .B(men_men_n1191_), .Y(men_men_n1213_));
  NO3        u1185(.A(men_men_n1213_), .B(men_men_n1195_), .C(men_men_n257_), .Y(men_men_n1214_));
  NO2        u1186(.A(men_men_n295_), .B(men_men_n45_), .Y(men_men_n1215_));
  AOI210     u1187(.A0(men_men_n1215_), .A1(men_men_n532_), .B0(men_men_n1201_), .Y(men_men_n1216_));
  NO2        u1188(.A(men_men_n1216_), .B(men_men_n334_), .Y(men_men_n1217_));
  NOi21      u1189(.An(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1218_));
  OAI210     u1190(.A0(men_men_n438_), .A1(men_men_n248_), .B0(men_men_n865_), .Y(men_men_n1219_));
  NO2        u1191(.A(men_men_n1219_), .B(men_men_n1218_), .Y(men_men_n1220_));
  OR2        u1192(.A(men_men_n571_), .B(men_men_n570_), .Y(men_men_n1221_));
  INV        u1193(.A(men_men_n1221_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n1222_), .B(men_men_n1220_), .Y(men_men_n1223_));
  NO2        u1195(.A(men_men_n714_), .B(men_men_n358_), .Y(men_men_n1224_));
  NOi21      u1196(.An(men_men_n1224_), .B(men_men_n150_), .Y(men_men_n1225_));
  AN2        u1197(.A(men_men_n902_), .B(men_men_n618_), .Y(men_men_n1226_));
  NO4        u1198(.A(men_men_n1226_), .B(men_men_n1225_), .C(men_men_n1223_), .D(men_men_n1217_), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n769_), .B(men_men_n275_), .Y(men_men_n1228_));
  OAI220     u1200(.A0(men_men_n700_), .A1(men_men_n47_), .B0(men_men_n223_), .B1(men_men_n588_), .Y(men_men_n1229_));
  OAI210     u1201(.A0(men_men_n275_), .A1(c), .B0(men_men_n614_), .Y(men_men_n1230_));
  AOI220     u1202(.A0(men_men_n1230_), .A1(men_men_n1229_), .B0(men_men_n1228_), .B1(men_men_n266_), .Y(men_men_n1231_));
  NO3        u1203(.A(men_men_n243_), .B(men_men_n102_), .C(men_men_n281_), .Y(men_men_n1232_));
  OAI220     u1204(.A0(men_men_n664_), .A1(men_men_n248_), .B0(men_men_n486_), .B1(men_men_n490_), .Y(men_men_n1233_));
  OAI210     u1205(.A0(l), .A1(i), .B0(k), .Y(men_men_n1234_));
  NO3        u1206(.A(men_men_n1234_), .B(men_men_n569_), .C(j), .Y(men_men_n1235_));
  NOi21      u1207(.An(men_men_n1235_), .B(men_men_n69_), .Y(men_men_n1236_));
  NO4        u1208(.A(men_men_n1236_), .B(men_men_n1233_), .C(men_men_n1232_), .D(men_men_n1053_), .Y(men_men_n1237_));
  NA3        u1209(.A(men_men_n1237_), .B(men_men_n1231_), .C(men_men_n1142_), .Y(men_men_n1238_));
  OR2        u1210(.A(men_men_n748_), .B(men_men_n518_), .Y(men_men_n1239_));
  OR3        u1211(.A(men_men_n361_), .B(men_men_n223_), .C(men_men_n588_), .Y(men_men_n1240_));
  NA2        u1212(.A(men_men_n1235_), .B(men_men_n756_), .Y(men_men_n1241_));
  NA3        u1213(.A(men_men_n1241_), .B(men_men_n1240_), .C(men_men_n1239_), .Y(men_men_n1242_));
  NA2        u1214(.A(men_men_n1224_), .B(men_men_n724_), .Y(men_men_n1243_));
  NO3        u1215(.A(men_men_n834_), .B(men_men_n475_), .C(men_men_n456_), .Y(men_men_n1244_));
  NA3        u1216(.A(men_men_n1244_), .B(men_men_n1243_), .C(men_men_n1196_), .Y(men_men_n1245_));
  NAi21      u1217(.An(j), .B(i), .Y(men_men_n1246_));
  NO4        u1218(.A(men_men_n1207_), .B(men_men_n1246_), .C(men_men_n423_), .D(men_men_n234_), .Y(men_men_n1247_));
  NO4        u1219(.A(men_men_n1247_), .B(men_men_n1245_), .C(men_men_n1242_), .D(men_men_n1238_), .Y(men_men_n1248_));
  NA4        u1220(.A(men_men_n1248_), .B(men_men_n1227_), .C(men_men_n1214_), .D(men_men_n1209_), .Y(men07));
  NAi32      u1221(.An(m), .Bn(b), .C(n), .Y(men_men_n1250_));
  NO3        u1222(.A(men_men_n1250_), .B(g), .C(f), .Y(men_men_n1251_));
  OAI210     u1223(.A0(men_men_n318_), .A1(men_men_n458_), .B0(men_men_n1251_), .Y(men_men_n1252_));
  NAi21      u1224(.An(f), .B(c), .Y(men_men_n1253_));
  NOi31      u1225(.An(n), .B(m), .C(b), .Y(men_men_n1254_));
  NO3        u1226(.A(men_men_n131_), .B(men_men_n430_), .C(h), .Y(men_men_n1255_));
  INV        u1227(.A(men_men_n1252_), .Y(men_men_n1256_));
  NOi41      u1228(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1257_));
  NA3        u1229(.A(men_men_n1257_), .B(men_men_n827_), .C(men_men_n393_), .Y(men_men_n1258_));
  NO2        u1230(.A(men_men_n1258_), .B(men_men_n53_), .Y(men_men_n1259_));
  NA2        u1231(.A(men_men_n1029_), .B(men_men_n219_), .Y(men_men_n1260_));
  NO2        u1232(.A(men_men_n1260_), .B(men_men_n57_), .Y(men_men_n1261_));
  NA2        u1233(.A(men_men_n85_), .B(men_men_n45_), .Y(men_men_n1262_));
  NO2        u1234(.A(men_men_n990_), .B(men_men_n423_), .Y(men_men_n1263_));
  NA3        u1235(.A(men_men_n1263_), .B(men_men_n1262_), .C(men_men_n213_), .Y(men_men_n1264_));
  NA2        u1236(.A(men_men_n1143_), .B(men_men_n289_), .Y(men_men_n1265_));
  NA2        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .Y(men_men_n1266_));
  NO4        u1238(.A(men_men_n1266_), .B(men_men_n1261_), .C(men_men_n1259_), .D(men_men_n1256_), .Y(men_men_n1267_));
  NO3        u1239(.A(e), .B(d), .C(c), .Y(men_men_n1268_));
  OAI210     u1240(.A0(men_men_n131_), .A1(men_men_n213_), .B0(men_men_n577_), .Y(men_men_n1269_));
  NA2        u1241(.A(men_men_n1269_), .B(men_men_n1268_), .Y(men_men_n1270_));
  INV        u1242(.A(men_men_n1270_), .Y(men_men_n1271_));
  OR2        u1243(.A(h), .B(f), .Y(men_men_n1272_));
  NO3        u1244(.A(n), .B(m), .C(i), .Y(men_men_n1273_));
  OAI210     u1245(.A0(men_men_n1051_), .A1(men_men_n158_), .B0(men_men_n1273_), .Y(men_men_n1274_));
  NO2        u1246(.A(i), .B(g), .Y(men_men_n1275_));
  OR3        u1247(.A(men_men_n1275_), .B(men_men_n1250_), .C(men_men_n68_), .Y(men_men_n1276_));
  OAI220     u1248(.A0(men_men_n1276_), .A1(men_men_n458_), .B0(men_men_n1274_), .B1(men_men_n1272_), .Y(men_men_n1277_));
  NA3        u1249(.A(men_men_n661_), .B(men_men_n649_), .C(men_men_n111_), .Y(men_men_n1278_));
  NA3        u1250(.A(men_men_n1254_), .B(l), .C(men_men_n642_), .Y(men_men_n1279_));
  AOI210     u1251(.A0(men_men_n1279_), .A1(men_men_n1278_), .B0(men_men_n45_), .Y(men_men_n1280_));
  NA2        u1252(.A(men_men_n1273_), .B(men_men_n613_), .Y(men_men_n1281_));
  NO2        u1253(.A(l), .B(k), .Y(men_men_n1282_));
  NO3        u1254(.A(men_men_n423_), .B(d), .C(c), .Y(men_men_n1283_));
  NO3        u1255(.A(men_men_n1280_), .B(men_men_n1277_), .C(men_men_n1271_), .Y(men_men_n1284_));
  NO2        u1256(.A(men_men_n148_), .B(h), .Y(men_men_n1285_));
  NO2        u1257(.A(g), .B(c), .Y(men_men_n1286_));
  NO2        u1258(.A(men_men_n431_), .B(a), .Y(men_men_n1287_));
  NA3        u1259(.A(men_men_n1287_), .B(k), .C(men_men_n112_), .Y(men_men_n1288_));
  NO2        u1260(.A(i), .B(h), .Y(men_men_n1289_));
  NA2        u1261(.A(men_men_n1289_), .B(men_men_n219_), .Y(men_men_n1290_));
  AOI210     u1262(.A0(men_men_n258_), .A1(men_men_n115_), .B0(men_men_n507_), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n1291_), .B(men_men_n1290_), .Y(men_men_n1292_));
  NO2        u1264(.A(men_men_n721_), .B(men_men_n187_), .Y(men_men_n1293_));
  NOi31      u1265(.An(m), .B(n), .C(b), .Y(men_men_n1294_));
  NOi31      u1266(.An(f), .B(d), .C(c), .Y(men_men_n1295_));
  NA2        u1267(.A(men_men_n1295_), .B(men_men_n1294_), .Y(men_men_n1296_));
  INV        u1268(.A(men_men_n1296_), .Y(men_men_n1297_));
  NO3        u1269(.A(men_men_n1297_), .B(men_men_n1293_), .C(men_men_n1292_), .Y(men_men_n1298_));
  OAI210     u1270(.A0(men_men_n182_), .A1(men_men_n502_), .B0(men_men_n999_), .Y(men_men_n1299_));
  AN3        u1271(.A(men_men_n1299_), .B(men_men_n1298_), .C(men_men_n1288_), .Y(men_men_n1300_));
  NA2        u1272(.A(men_men_n1254_), .B(men_men_n369_), .Y(men_men_n1301_));
  NO2        u1273(.A(i), .B(men_men_n212_), .Y(men_men_n1302_));
  NA4        u1274(.A(men_men_n1078_), .B(men_men_n1302_), .C(men_men_n103_), .D(m), .Y(men_men_n1303_));
  INV        u1275(.A(men_men_n1303_), .Y(men_men_n1304_));
  NO4        u1276(.A(men_men_n131_), .B(g), .C(f), .D(e), .Y(men_men_n1305_));
  NA2        u1277(.A(men_men_n290_), .B(h), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n194_), .B(men_men_n97_), .Y(men_men_n1307_));
  OR2        u1279(.A(e), .B(a), .Y(men_men_n1308_));
  NA2        u1280(.A(men_men_n30_), .B(h), .Y(men_men_n1309_));
  NO2        u1281(.A(men_men_n1309_), .B(men_men_n1018_), .Y(men_men_n1310_));
  NA2        u1282(.A(men_men_n1257_), .B(men_men_n1282_), .Y(men_men_n1311_));
  INV        u1283(.A(men_men_n1311_), .Y(men_men_n1312_));
  OR3        u1284(.A(men_men_n518_), .B(men_men_n517_), .C(men_men_n111_), .Y(men_men_n1313_));
  NA2        u1285(.A(men_men_n1049_), .B(men_men_n390_), .Y(men_men_n1314_));
  OAI220     u1286(.A0(men_men_n1314_), .A1(men_men_n416_), .B0(men_men_n1313_), .B1(men_men_n295_), .Y(men_men_n1315_));
  AO210      u1287(.A0(men_men_n1315_), .A1(men_men_n115_), .B0(men_men_n1312_), .Y(men_men_n1316_));
  NO3        u1288(.A(men_men_n1316_), .B(men_men_n1310_), .C(men_men_n1304_), .Y(men_men_n1317_));
  NA4        u1289(.A(men_men_n1317_), .B(men_men_n1300_), .C(men_men_n1284_), .D(men_men_n1267_), .Y(men_men_n1318_));
  NA2        u1290(.A(men_men_n369_), .B(men_men_n53_), .Y(men_men_n1319_));
  AOI210     u1291(.A0(men_men_n1319_), .A1(men_men_n990_), .B0(men_men_n1281_), .Y(men_men_n1320_));
  NA2        u1292(.A(men_men_n214_), .B(men_men_n179_), .Y(men_men_n1321_));
  AOI210     u1293(.A0(men_men_n1321_), .A1(men_men_n1117_), .B0(men_men_n1319_), .Y(men_men_n1322_));
  NO2        u1294(.A(men_men_n1022_), .B(men_men_n1018_), .Y(men_men_n1323_));
  NO3        u1295(.A(men_men_n1323_), .B(men_men_n1322_), .C(men_men_n1320_), .Y(men_men_n1324_));
  NO2        u1296(.A(men_men_n378_), .B(j), .Y(men_men_n1325_));
  NA3        u1297(.A(g), .B(men_men_n1325_), .C(men_men_n160_), .Y(men_men_n1326_));
  NO3        u1298(.A(men_men_n1018_), .B(men_men_n555_), .C(g), .Y(men_men_n1327_));
  NOi21      u1299(.An(men_men_n1321_), .B(men_men_n1327_), .Y(men_men_n1328_));
  AOI210     u1300(.A0(men_men_n1328_), .A1(men_men_n1307_), .B0(men_men_n990_), .Y(men_men_n1329_));
  OR2        u1301(.A(n), .B(i), .Y(men_men_n1330_));
  OAI210     u1302(.A0(men_men_n1330_), .A1(men_men_n1010_), .B0(men_men_n49_), .Y(men_men_n1331_));
  AOI220     u1303(.A0(men_men_n1331_), .A1(men_men_n1105_), .B0(men_men_n794_), .B1(men_men_n194_), .Y(men_men_n1332_));
  INV        u1304(.A(men_men_n1332_), .Y(men_men_n1333_));
  NO2        u1305(.A(men_men_n223_), .B(k), .Y(men_men_n1334_));
  NO2        u1306(.A(men_men_n1333_), .B(men_men_n1329_), .Y(men_men_n1335_));
  INV        u1307(.A(men_men_n49_), .Y(men_men_n1336_));
  NA2        u1308(.A(men_men_n1032_), .B(men_men_n1336_), .Y(men_men_n1337_));
  NO2        u1309(.A(men_men_n1337_), .B(j), .Y(men_men_n1338_));
  AOI210     u1310(.A0(men_men_n502_), .A1(h), .B0(men_men_n65_), .Y(men_men_n1339_));
  NA2        u1311(.A(men_men_n1339_), .B(men_men_n1287_), .Y(men_men_n1340_));
  NO2        u1312(.A(men_men_n1246_), .B(men_men_n175_), .Y(men_men_n1341_));
  NOi21      u1313(.An(d), .B(f), .Y(men_men_n1342_));
  NO3        u1314(.A(men_men_n1295_), .B(men_men_n1342_), .C(men_men_n40_), .Y(men_men_n1343_));
  NA2        u1315(.A(men_men_n1343_), .B(men_men_n1341_), .Y(men_men_n1344_));
  NO2        u1316(.A(men_men_n295_), .B(c), .Y(men_men_n1345_));
  NA2        u1317(.A(men_men_n1345_), .B(men_men_n519_), .Y(men_men_n1346_));
  NA3        u1318(.A(men_men_n1346_), .B(men_men_n1344_), .C(men_men_n1340_), .Y(men_men_n1347_));
  NO2        u1319(.A(men_men_n1347_), .B(men_men_n1338_), .Y(men_men_n1348_));
  NA4        u1320(.A(men_men_n1348_), .B(men_men_n1335_), .C(men_men_n1326_), .D(men_men_n1324_), .Y(men_men_n1349_));
  OAI210     u1321(.A0(men_men_n1305_), .A1(men_men_n1254_), .B0(men_men_n841_), .Y(men_men_n1350_));
  OAI220     u1322(.A0(men_men_n979_), .A1(men_men_n131_), .B0(h), .B1(men_men_n175_), .Y(men_men_n1351_));
  NA2        u1323(.A(men_men_n1351_), .B(men_men_n594_), .Y(men_men_n1352_));
  NA2        u1324(.A(men_men_n1352_), .B(men_men_n1350_), .Y(men_men_n1353_));
  NA2        u1325(.A(men_men_n1286_), .B(men_men_n1342_), .Y(men_men_n1354_));
  NO2        u1326(.A(men_men_n1354_), .B(m), .Y(men_men_n1355_));
  NA3        u1327(.A(men_men_n1029_), .B(men_men_n107_), .C(men_men_n219_), .Y(men_men_n1356_));
  NO2        u1328(.A(men_men_n152_), .B(men_men_n181_), .Y(men_men_n1357_));
  OAI210     u1329(.A0(men_men_n1357_), .A1(men_men_n109_), .B0(men_men_n1294_), .Y(men_men_n1358_));
  NA2        u1330(.A(men_men_n1358_), .B(men_men_n1356_), .Y(men_men_n1359_));
  NO3        u1331(.A(men_men_n1359_), .B(men_men_n1355_), .C(men_men_n1353_), .Y(men_men_n1360_));
  NO2        u1332(.A(men_men_n1253_), .B(e), .Y(men_men_n1361_));
  NA2        u1333(.A(men_men_n1361_), .B(men_men_n388_), .Y(men_men_n1362_));
  NA2        u1334(.A(men_men_n1060_), .B(men_men_n605_), .Y(men_men_n1363_));
  OR3        u1335(.A(men_men_n1334_), .B(men_men_n1143_), .C(men_men_n131_), .Y(men_men_n1364_));
  OAI220     u1336(.A0(men_men_n1364_), .A1(men_men_n1362_), .B0(men_men_n1363_), .B1(men_men_n425_), .Y(men_men_n1365_));
  NO2        u1337(.A(men_men_n1313_), .B(a), .Y(men_men_n1366_));
  NO2        u1338(.A(men_men_n1366_), .B(men_men_n1365_), .Y(men_men_n1367_));
  NO2        u1339(.A(men_men_n181_), .B(c), .Y(men_men_n1368_));
  OAI210     u1340(.A0(men_men_n1368_), .A1(men_men_n1361_), .B0(men_men_n179_), .Y(men_men_n1369_));
  AOI220     u1341(.A0(men_men_n1369_), .A1(men_men_n1012_), .B0(men_men_n509_), .B1(men_men_n358_), .Y(men_men_n1370_));
  NA2        u1342(.A(men_men_n517_), .B(g), .Y(men_men_n1371_));
  NA2        u1343(.A(men_men_n1371_), .B(men_men_n1283_), .Y(men_men_n1372_));
  NO2        u1344(.A(men_men_n1308_), .B(f), .Y(men_men_n1373_));
  AOI210     u1345(.A0(men_men_n1060_), .A1(a), .B0(men_men_n1373_), .Y(men_men_n1374_));
  OAI220     u1346(.A0(men_men_n1374_), .A1(men_men_n65_), .B0(men_men_n1372_), .B1(men_men_n212_), .Y(men_men_n1375_));
  AOI210     u1347(.A0(men_men_n858_), .A1(men_men_n400_), .B0(men_men_n104_), .Y(men_men_n1376_));
  OR2        u1348(.A(men_men_n1376_), .B(men_men_n517_), .Y(men_men_n1377_));
  NO2        u1349(.A(men_men_n1377_), .B(men_men_n175_), .Y(men_men_n1378_));
  NA2        u1350(.A(men_men_n1255_), .B(men_men_n182_), .Y(men_men_n1379_));
  NO2        u1351(.A(men_men_n49_), .B(l), .Y(men_men_n1380_));
  OAI210     u1352(.A0(men_men_n1308_), .A1(men_men_n822_), .B0(men_men_n458_), .Y(men_men_n1381_));
  OAI210     u1353(.A0(men_men_n1381_), .A1(men_men_n1032_), .B0(men_men_n1380_), .Y(men_men_n1382_));
  NO2        u1354(.A(men_men_n253_), .B(g), .Y(men_men_n1383_));
  NO2        u1355(.A(m), .B(i), .Y(men_men_n1384_));
  BUFFER     u1356(.A(men_men_n1384_), .Y(men_men_n1385_));
  AOI220     u1357(.A0(men_men_n1385_), .A1(men_men_n1285_), .B0(men_men_n1011_), .B1(men_men_n1383_), .Y(men_men_n1386_));
  NA3        u1358(.A(men_men_n1386_), .B(men_men_n1382_), .C(men_men_n1379_), .Y(men_men_n1387_));
  NO4        u1359(.A(men_men_n1387_), .B(men_men_n1378_), .C(men_men_n1375_), .D(men_men_n1370_), .Y(men_men_n1388_));
  NA3        u1360(.A(men_men_n1388_), .B(men_men_n1367_), .C(men_men_n1360_), .Y(men_men_n1389_));
  NA3        u1361(.A(men_men_n908_), .B(men_men_n138_), .C(men_men_n46_), .Y(men_men_n1390_));
  NO2        u1362(.A(men_men_n149_), .B(men_men_n1390_), .Y(men_men_n1391_));
  AO210      u1363(.A0(men_men_n132_), .A1(l), .B0(men_men_n1301_), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n68_), .B(c), .Y(men_men_n1393_));
  NO4        u1365(.A(men_men_n1272_), .B(men_men_n185_), .C(men_men_n430_), .D(men_men_n45_), .Y(men_men_n1394_));
  AOI210     u1366(.A0(men_men_n1341_), .A1(men_men_n1393_), .B0(men_men_n1394_), .Y(men_men_n1395_));
  NA2        u1367(.A(men_men_n1395_), .B(men_men_n1392_), .Y(men_men_n1396_));
  NO2        u1368(.A(men_men_n1396_), .B(men_men_n1391_), .Y(men_men_n1397_));
  NO4        u1369(.A(men_men_n223_), .B(men_men_n185_), .C(men_men_n258_), .D(k), .Y(men_men_n1398_));
  NO2        u1370(.A(men_men_n1390_), .B(men_men_n109_), .Y(men_men_n1399_));
  NOi21      u1371(.An(men_men_n1255_), .B(e), .Y(men_men_n1400_));
  NO3        u1372(.A(men_men_n1400_), .B(men_men_n1399_), .C(men_men_n1398_), .Y(men_men_n1401_));
  AOI220     u1373(.A0(men_men_n1384_), .A1(men_men_n613_), .B0(men_men_n996_), .B1(men_men_n161_), .Y(men_men_n1402_));
  NOi31      u1374(.An(men_men_n30_), .B(men_men_n1402_), .C(n), .Y(men_men_n1403_));
  INV        u1375(.A(men_men_n1403_), .Y(men_men_n1404_));
  NA3        u1376(.A(men_men_n1404_), .B(men_men_n1401_), .C(men_men_n1397_), .Y(men_men_n1405_));
  OR4        u1377(.A(men_men_n1405_), .B(men_men_n1389_), .C(men_men_n1349_), .D(men_men_n1318_), .Y(men04));
  NOi31      u1378(.An(men_men_n1305_), .B(men_men_n1306_), .C(men_men_n984_), .Y(men_men_n1407_));
  NO4        u1379(.A(d), .B(men_men_n974_), .C(men_men_n459_), .D(j), .Y(men_men_n1408_));
  OR3        u1380(.A(men_men_n1408_), .B(men_men_n1407_), .C(men_men_n1001_), .Y(men_men_n1409_));
  NO3        u1381(.A(men_men_n1262_), .B(men_men_n89_), .C(k), .Y(men_men_n1410_));
  AOI210     u1382(.A0(men_men_n1410_), .A1(men_men_n995_), .B0(men_men_n1119_), .Y(men_men_n1411_));
  NA2        u1383(.A(men_men_n1411_), .B(men_men_n1145_), .Y(men_men_n1412_));
  NO4        u1384(.A(men_men_n1412_), .B(men_men_n1409_), .C(men_men_n1009_), .D(men_men_n989_), .Y(men_men_n1413_));
  NA4        u1385(.A(men_men_n1413_), .B(men_men_n1062_), .C(men_men_n1047_), .D(men_men_n1035_), .Y(men05));
  INV        u1386(.A(men_men_n577_), .Y(men_men_n1417_));
  INV        u1387(.A(men_men_n135_), .Y(men_men_n1418_));
  INV        u1388(.A(men_men_n219_), .Y(men_men_n1419_));
  INV        u1389(.A(men_men_n166_), .Y(men_men_n1420_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule