//Benchmark atmr_alu4_1266_0.5

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n88_, ori_ori_n89_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n339_, ori_ori_n340_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n121_, mai_mai_n122_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n132_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  AO210      o008(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n31_));
  OR2        o009(.A(ori_ori_n31_), .B(i_11_), .Y(ori_ori_n32_));
  NA2        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .Y(ori_ori_n33_));
  XO2        o011(.A(ori_ori_n33_), .B(ori_ori_n23_), .Y(ori_ori_n34_));
  INV        o012(.A(i_4_), .Y(ori_ori_n35_));
  INV        o013(.A(i_10_), .Y(ori_ori_n36_));
  NAi21      o014(.An(i_11_), .B(i_9_), .Y(ori_ori_n37_));
  NO3        o015(.A(ori_ori_n37_), .B(i_12_), .C(ori_ori_n36_), .Y(ori_ori_n38_));
  INV        o016(.A(ori_ori_n34_), .Y(ori1));
  INV        o017(.A(i_11_), .Y(ori_ori_n40_));
  NO2        o018(.A(ori_ori_n40_), .B(i_6_), .Y(ori_ori_n41_));
  INV        o019(.A(i_2_), .Y(ori_ori_n42_));
  INV        o020(.A(i_5_), .Y(ori_ori_n43_));
  NA2        o021(.A(i_7_), .B(i_9_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n41_), .Y(ori_ori_n45_));
  NAi21      o023(.An(i_2_), .B(i_7_), .Y(ori_ori_n46_));
  INV        o024(.A(i_1_), .Y(ori_ori_n47_));
  NA2        o025(.A(ori_ori_n47_), .B(i_6_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n49_));
  INV        o027(.A(i_0_), .Y(ori_ori_n50_));
  NAi21      o028(.An(i_5_), .B(i_10_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_5_), .B(i_9_), .Y(ori_ori_n52_));
  AOI210     o030(.A0(ori_ori_n52_), .A1(ori_ori_n51_), .B0(ori_ori_n50_), .Y(ori_ori_n53_));
  INV        o031(.A(ori_ori_n53_), .Y(ori_ori_n54_));
  NA2        o032(.A(ori_ori_n49_), .B(ori_ori_n54_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n55_), .B(i_0_), .Y(ori_ori_n56_));
  NA2        o034(.A(i_12_), .B(i_5_), .Y(ori_ori_n57_));
  INV        o035(.A(i_6_), .Y(ori_ori_n58_));
  NO2        o036(.A(i_2_), .B(i_7_), .Y(ori_ori_n59_));
  INV        o037(.A(ori_ori_n59_), .Y(ori_ori_n60_));
  OAI210     o038(.A0(i_3_), .A1(i_8_), .B0(ori_ori_n60_), .Y(ori_ori_n61_));
  NAi21      o039(.An(i_6_), .B(i_10_), .Y(ori_ori_n62_));
  NA2        o040(.A(i_6_), .B(i_9_), .Y(ori_ori_n63_));
  AOI210     o041(.A0(ori_ori_n63_), .A1(ori_ori_n62_), .B0(ori_ori_n47_), .Y(ori_ori_n64_));
  NA2        o042(.A(i_2_), .B(i_6_), .Y(ori_ori_n65_));
  AOI210     o043(.A0(ori_ori_n62_), .A1(ori_ori_n61_), .B0(ori_ori_n57_), .Y(ori_ori_n66_));
  NAi21      o044(.An(i_6_), .B(i_11_), .Y(ori_ori_n67_));
  INV        o045(.A(i_7_), .Y(ori_ori_n68_));
  NA2        o046(.A(ori_ori_n42_), .B(ori_ori_n68_), .Y(ori_ori_n69_));
  NO2        o047(.A(i_0_), .B(i_5_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_12_), .B(i_3_), .Y(ori_ori_n71_));
  INV        o049(.A(i_7_), .Y(ori_ori_n72_));
  BUFFER     o050(.A(ori_ori_n57_), .Y(ori_ori_n73_));
  NA2        o051(.A(i_12_), .B(i_7_), .Y(ori_ori_n74_));
  NA2        o052(.A(i_11_), .B(i_12_), .Y(ori_ori_n75_));
  NOi21      o053(.An(i_1_), .B(i_5_), .Y(ori_ori_n76_));
  NA2        o054(.A(ori_ori_n76_), .B(i_11_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n78_));
  NA2        o056(.A(ori_ori_n78_), .B(i_10_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n42_), .Y(ori_ori_n80_));
  NA2        o058(.A(ori_ori_n63_), .B(ori_ori_n62_), .Y(ori_ori_n81_));
  NAi21      o059(.An(i_3_), .B(i_8_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_1_), .B(ori_ori_n58_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_6_), .B(i_5_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n77_), .Y(ori_ori_n85_));
  NO3        o063(.A(ori_ori_n85_), .B(ori_ori_n340_), .C(ori_ori_n66_), .Y(ori_ori_n86_));
  NA3        o064(.A(ori_ori_n86_), .B(ori_ori_n56_), .C(ori_ori_n45_), .Y(ori2));
  NO2        o065(.A(ori_ori_n47_), .B(ori_ori_n36_), .Y(ori_ori_n88_));
  INV        o066(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  NA3        o067(.A(ori_ori_n89_), .B(ori_ori_n54_), .C(ori_ori_n30_), .Y(ori0));
  NA2        o068(.A(i_7_), .B(i_6_), .Y(ori_ori_n91_));
  NO2        o069(.A(i_0_), .B(i_1_), .Y(ori_ori_n92_));
  NA2        o070(.A(i_2_), .B(i_3_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(i_4_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_1_), .B(i_5_), .Y(ori_ori_n95_));
  OR2        o073(.A(i_0_), .B(i_1_), .Y(ori_ori_n96_));
  NOi21      o074(.An(i_4_), .B(i_9_), .Y(ori_ori_n97_));
  NOi21      o075(.An(i_11_), .B(i_13_), .Y(ori_ori_n98_));
  NA2        o076(.A(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n100_));
  NAi21      o078(.An(i_4_), .B(i_12_), .Y(ori_ori_n101_));
  INV        o079(.A(i_8_), .Y(ori_ori_n102_));
  NO2        o080(.A(i_3_), .B(i_8_), .Y(ori_ori_n103_));
  NO3        o081(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n104_));
  NO2        o082(.A(i_13_), .B(i_9_), .Y(ori_ori_n105_));
  NAi21      o083(.An(i_12_), .B(i_3_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n40_), .B(i_5_), .Y(ori_ori_n107_));
  INV        o085(.A(i_13_), .Y(ori_ori_n108_));
  NO2        o086(.A(i_12_), .B(ori_ori_n108_), .Y(ori_ori_n109_));
  INV        o087(.A(i_12_), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n40_), .B(ori_ori_n110_), .Y(ori_ori_n111_));
  NO3        o089(.A(i_11_), .B(i_7_), .C(ori_ori_n36_), .Y(ori_ori_n112_));
  INV        o090(.A(i_0_), .Y(ori_ori_n113_));
  NOi41      o091(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n114_));
  NO2        o092(.A(i_11_), .B(ori_ori_n108_), .Y(ori_ori_n115_));
  INV        o093(.A(i_5_), .Y(ori_ori_n116_));
  NA2        o094(.A(i_3_), .B(i_9_), .Y(ori_ori_n117_));
  NAi21      o095(.An(i_7_), .B(i_10_), .Y(ori_ori_n118_));
  NO2        o096(.A(ori_ori_n118_), .B(ori_ori_n117_), .Y(ori_ori_n119_));
  NA3        o097(.A(ori_ori_n119_), .B(ori_ori_n116_), .C(ori_ori_n48_), .Y(ori_ori_n120_));
  INV        o098(.A(ori_ori_n120_), .Y(ori_ori_n121_));
  INV        o099(.A(ori_ori_n91_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n110_), .B(i_13_), .Y(ori_ori_n123_));
  NO2        o101(.A(ori_ori_n123_), .B(ori_ori_n52_), .Y(ori_ori_n124_));
  AOI220     o102(.A0(ori_ori_n124_), .A1(ori_ori_n122_), .B0(ori_ori_n121_), .B1(ori_ori_n115_), .Y(ori_ori_n125_));
  NA2        o103(.A(i_12_), .B(i_6_), .Y(ori_ori_n126_));
  AN2        o104(.A(i_3_), .B(i_10_), .Y(ori_ori_n127_));
  NO2        o105(.A(i_5_), .B(ori_ori_n36_), .Y(ori_ori_n128_));
  NO2        o106(.A(ori_ori_n42_), .B(ori_ori_n26_), .Y(ori_ori_n129_));
  NO2        o107(.A(i_2_), .B(i_3_), .Y(ori_ori_n130_));
  NO2        o108(.A(i_12_), .B(i_10_), .Y(ori_ori_n131_));
  INV        o109(.A(i_1_), .Y(ori_ori_n132_));
  NAi21      o110(.An(i_3_), .B(i_4_), .Y(ori_ori_n133_));
  AN2        o111(.A(i_12_), .B(i_5_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_5_), .B(i_10_), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n136_));
  NO3        o114(.A(ori_ori_n58_), .B(ori_ori_n43_), .C(i_9_), .Y(ori_ori_n137_));
  NO2        o115(.A(i_0_), .B(i_11_), .Y(ori_ori_n138_));
  NAi21      o116(.An(i_9_), .B(i_4_), .Y(ori_ori_n139_));
  OR2        o117(.A(i_13_), .B(i_10_), .Y(ori_ori_n140_));
  NO3        o118(.A(ori_ori_n140_), .B(ori_ori_n75_), .C(ori_ori_n139_), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n68_), .B(ori_ori_n25_), .Y(ori_ori_n142_));
  NO2        o120(.A(i_10_), .B(i_9_), .Y(ori_ori_n143_));
  NAi21      o121(.An(i_12_), .B(i_8_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n144_), .B(i_3_), .Y(ori_ori_n145_));
  NO3        o123(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n146_));
  NA2        o124(.A(ori_ori_n126_), .B(ori_ori_n67_), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n147_), .B(ori_ori_n146_), .Y(ori_ori_n148_));
  NA2        o126(.A(ori_ori_n115_), .B(ori_ori_n128_), .Y(ori_ori_n149_));
  NO3        o127(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n150_));
  INV        o128(.A(ori_ori_n150_), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n151_), .B(ori_ori_n149_), .Y(ori_ori_n152_));
  INV        o130(.A(ori_ori_n152_), .Y(ori_ori_n153_));
  NO2        o131(.A(i_11_), .B(i_1_), .Y(ori_ori_n154_));
  NA3        o132(.A(ori_ori_n114_), .B(ori_ori_n98_), .C(ori_ori_n84_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n42_), .B(ori_ori_n40_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n96_), .B(i_3_), .Y(ori_ori_n157_));
  NAi31      o135(.An(ori_ori_n156_), .B(ori_ori_n157_), .C(ori_ori_n109_), .Y(ori_ori_n158_));
  NA3        o136(.A(ori_ori_n136_), .B(ori_ori_n100_), .C(ori_ori_n94_), .Y(ori_ori_n159_));
  NA3        o137(.A(ori_ori_n159_), .B(ori_ori_n158_), .C(ori_ori_n155_), .Y(ori_ori_n160_));
  INV        o138(.A(ori_ori_n160_), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n146_), .B(ori_ori_n134_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n150_), .B(ori_ori_n135_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n161_), .B(ori_ori_n153_), .Y(ori_ori_n164_));
  NO2        o142(.A(ori_ori_n35_), .B(i_8_), .Y(ori_ori_n165_));
  AOI210     o143(.A0(ori_ori_n38_), .A1(i_13_), .B0(ori_ori_n141_), .Y(ori_ori_n166_));
  INV        o144(.A(ori_ori_n166_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n140_), .B(i_1_), .Y(ori_ori_n168_));
  NOi31      o146(.An(ori_ori_n168_), .B(ori_ori_n147_), .C(ori_ori_n50_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n74_), .B(ori_ori_n23_), .Y(ori_ori_n170_));
  NO2        o148(.A(i_12_), .B(ori_ori_n58_), .Y(ori_ori_n171_));
  NO2        o149(.A(ori_ori_n167_), .B(ori_ori_n164_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(ori_ori_n125_), .Y(ori7));
  NO2        o151(.A(ori_ori_n65_), .B(ori_ori_n44_), .Y(ori_ori_n174_));
  NA3        o152(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n175_));
  NO2        o153(.A(ori_ori_n110_), .B(i_4_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n176_), .B(i_8_), .Y(ori_ori_n177_));
  NO2        o155(.A(ori_ori_n71_), .B(ori_ori_n175_), .Y(ori_ori_n178_));
  NA2        o156(.A(i_2_), .B(ori_ori_n58_), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n103_), .B(ori_ori_n104_), .Y(ori_ori_n180_));
  NA2        o158(.A(i_4_), .B(i_8_), .Y(ori_ori_n181_));
  NA2        o159(.A(ori_ori_n181_), .B(ori_ori_n127_), .Y(ori_ori_n182_));
  OAI220     o160(.A0(ori_ori_n182_), .A1(ori_ori_n179_), .B0(ori_ori_n180_), .B1(i_13_), .Y(ori_ori_n183_));
  NO3        o161(.A(ori_ori_n183_), .B(ori_ori_n178_), .C(ori_ori_n174_), .Y(ori_ori_n184_));
  AOI210     o162(.A0(ori_ori_n82_), .A1(ori_ori_n46_), .B0(i_10_), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n185_), .B(ori_ori_n110_), .Y(ori_ori_n186_));
  OR2        o164(.A(i_6_), .B(i_10_), .Y(ori_ori_n187_));
  OR2        o165(.A(ori_ori_n186_), .B(i_9_), .Y(ori_ori_n188_));
  AOI210     o166(.A0(ori_ori_n188_), .A1(ori_ori_n184_), .B0(ori_ori_n47_), .Y(ori_ori_n189_));
  NOi21      o167(.An(i_11_), .B(i_7_), .Y(ori_ori_n190_));
  AO210      o168(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n191_), .B(ori_ori_n190_), .Y(ori_ori_n192_));
  NA2        o170(.A(ori_ori_n192_), .B(ori_ori_n105_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n193_), .B(ori_ori_n47_), .Y(ori_ori_n194_));
  NO2        o172(.A(i_1_), .B(i_12_), .Y(ori_ori_n195_));
  NA2        o173(.A(ori_ori_n194_), .B(i_6_), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n148_), .Y(ori_ori_n197_));
  NO3        o175(.A(ori_ori_n187_), .B(i_7_), .C(ori_ori_n23_), .Y(ori_ori_n198_));
  AOI210     o176(.A0(i_1_), .A1(ori_ori_n119_), .B0(ori_ori_n198_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(ori_ori_n40_), .Y(ori_ori_n200_));
  INV        o178(.A(i_2_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n88_), .B(i_9_), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n202_), .B(ori_ori_n201_), .Y(ori_ori_n203_));
  AOI210     o181(.A0(ori_ori_n154_), .A1(ori_ori_n142_), .B0(ori_ori_n112_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n204_), .B(ori_ori_n179_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_11_), .B(ori_ori_n36_), .Y(ori_ori_n206_));
  OR2        o184(.A(ori_ori_n205_), .B(ori_ori_n203_), .Y(ori_ori_n207_));
  NO3        o185(.A(ori_ori_n207_), .B(ori_ori_n200_), .C(ori_ori_n197_), .Y(ori_ori_n208_));
  NO2        o186(.A(i_7_), .B(ori_ori_n40_), .Y(ori_ori_n209_));
  NO3        o187(.A(ori_ori_n209_), .B(ori_ori_n129_), .C(ori_ori_n111_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n75_), .B(ori_ori_n36_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(i_6_), .Y(ori_ori_n212_));
  NO2        o190(.A(ori_ori_n58_), .B(i_9_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n213_), .B(ori_ori_n47_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n214_), .B(ori_ori_n195_), .Y(ori_ori_n215_));
  NO4        o193(.A(ori_ori_n215_), .B(ori_ori_n212_), .C(ori_ori_n210_), .D(i_4_), .Y(ori_ori_n216_));
  INV        o194(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  NA3        o195(.A(ori_ori_n217_), .B(ori_ori_n208_), .C(ori_ori_n196_), .Y(ori_ori_n218_));
  AOI210     o196(.A0(ori_ori_n126_), .A1(ori_ori_n67_), .B0(i_1_), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n133_), .B(i_2_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n221_));
  INV        o199(.A(ori_ori_n221_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n44_), .B(i_12_), .Y(ori_ori_n223_));
  INV        o201(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n224_), .B(ori_ori_n65_), .Y(ori_ori_n225_));
  INV        o203(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NA2        o204(.A(ori_ori_n81_), .B(i_13_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n219_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n64_), .B(ori_ori_n69_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n229_), .B(ori_ori_n177_), .Y(ori_ori_n230_));
  NO2        o208(.A(ori_ori_n230_), .B(ori_ori_n228_), .Y(ori_ori_n231_));
  OR2        o209(.A(i_11_), .B(i_6_), .Y(ori_ori_n232_));
  NO2        o210(.A(i_4_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NA2        o211(.A(ori_ori_n233_), .B(ori_ori_n47_), .Y(ori_ori_n234_));
  NO2        o212(.A(i_2_), .B(i_12_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n132_), .B(ori_ori_n235_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n236_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n237_), .B(ori_ori_n41_), .Y(ori_ori_n238_));
  NA4        o216(.A(ori_ori_n238_), .B(ori_ori_n234_), .C(ori_ori_n231_), .D(ori_ori_n226_), .Y(ori_ori_n239_));
  OR4        o217(.A(ori_ori_n239_), .B(ori_ori_n222_), .C(ori_ori_n218_), .D(ori_ori_n189_), .Y(ori5));
  AN2        o218(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n241_));
  NA3        o219(.A(ori_ori_n241_), .B(ori_ori_n235_), .C(i_7_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n177_), .B(i_11_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n59_), .B(ori_ori_n243_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n244_), .B(ori_ori_n242_), .Y(ori_ori_n245_));
  NO2        o223(.A(ori_ori_n78_), .B(ori_ori_n23_), .Y(ori_ori_n246_));
  NA2        o224(.A(i_12_), .B(i_8_), .Y(ori_ori_n247_));
  OAI210     o225(.A0(ori_ori_n42_), .A1(i_3_), .B0(ori_ori_n247_), .Y(ori_ori_n248_));
  INV        o226(.A(ori_ori_n143_), .Y(ori_ori_n249_));
  AOI220     o227(.A0(ori_ori_n130_), .A1(ori_ori_n170_), .B0(ori_ori_n248_), .B1(ori_ori_n246_), .Y(ori_ori_n250_));
  INV        o228(.A(ori_ori_n250_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n251_), .B(ori_ori_n245_), .Y(ori_ori_n252_));
  INV        o230(.A(ori_ori_n98_), .Y(ori_ori_n253_));
  INV        o231(.A(ori_ori_n114_), .Y(ori_ori_n254_));
  OAI210     o232(.A0(ori_ori_n220_), .A1(ori_ori_n145_), .B0(ori_ori_n72_), .Y(ori_ori_n255_));
  AOI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n254_), .B0(ori_ori_n253_), .Y(ori_ori_n256_));
  INV        o234(.A(ori_ori_n256_), .Y(ori_ori_n257_));
  INV        o235(.A(ori_ori_n99_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n191_), .B(ori_ori_n37_), .C(ori_ori_n26_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n258_), .B(ori_ori_n259_), .Y(ori_ori_n260_));
  NO2        o238(.A(ori_ori_n260_), .B(ori_ori_n102_), .Y(ori_ori_n261_));
  OA210      o239(.A0(ori_ori_n192_), .A1(ori_ori_n80_), .B0(i_13_), .Y(ori_ori_n262_));
  AOI210     o240(.A0(ori_ori_n106_), .A1(ori_ori_n93_), .B0(ori_ori_n165_), .Y(ori_ori_n263_));
  NA2        o241(.A(ori_ori_n263_), .B(ori_ori_n142_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n68_), .B(ori_ori_n127_), .Y(ori_ori_n265_));
  OAI210     o243(.A0(ori_ori_n265_), .A1(i_11_), .B0(ori_ori_n264_), .Y(ori_ori_n266_));
  NO3        o244(.A(ori_ori_n266_), .B(ori_ori_n262_), .C(ori_ori_n261_), .Y(ori_ori_n267_));
  NA2        o245(.A(ori_ori_n170_), .B(ori_ori_n28_), .Y(ori_ori_n268_));
  NA4        o246(.A(ori_ori_n268_), .B(ori_ori_n267_), .C(ori_ori_n257_), .D(ori_ori_n252_), .Y(ori6));
  NA2        o247(.A(ori_ori_n171_), .B(ori_ori_n47_), .Y(ori_ori_n270_));
  INV        o248(.A(ori_ori_n270_), .Y(ori_ori_n271_));
  NA2        o249(.A(ori_ori_n271_), .B(ori_ori_n50_), .Y(ori_ori_n272_));
  INV        o250(.A(ori_ori_n131_), .Y(ori_ori_n273_));
  NA2        o251(.A(ori_ori_n52_), .B(ori_ori_n83_), .Y(ori_ori_n274_));
  INV        o252(.A(ori_ori_n78_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n275_), .B(ori_ori_n42_), .Y(ori_ori_n276_));
  AOI210     o254(.A0(ori_ori_n276_), .A1(ori_ori_n274_), .B0(ori_ori_n273_), .Y(ori_ori_n277_));
  NAi32      o255(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n278_));
  NO2        o256(.A(ori_ori_n232_), .B(ori_ori_n278_), .Y(ori_ori_n279_));
  OR2        o257(.A(ori_ori_n279_), .B(ori_ori_n277_), .Y(ori_ori_n280_));
  BUFFER     o258(.A(ori_ori_n192_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n281_), .B(ori_ori_n92_), .Y(ori_ori_n282_));
  AO210      o260(.A0(ori_ori_n163_), .A1(ori_ori_n249_), .B0(ori_ori_n35_), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n283_), .B(ori_ori_n282_), .Y(ori_ori_n284_));
  NA2        o262(.A(ori_ori_n137_), .B(ori_ori_n49_), .Y(ori_ori_n285_));
  INV        o263(.A(ori_ori_n285_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n145_), .B(ori_ori_n143_), .Y(ori_ori_n287_));
  NA2        o265(.A(ori_ori_n73_), .B(ori_ori_n138_), .Y(ori_ori_n288_));
  NA2        o266(.A(ori_ori_n288_), .B(ori_ori_n287_), .Y(ori_ori_n289_));
  NO4        o267(.A(ori_ori_n289_), .B(ori_ori_n286_), .C(ori_ori_n284_), .D(ori_ori_n280_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n290_), .B(ori_ori_n272_), .Y(ori3));
  NO3        o269(.A(ori_ori_n134_), .B(ori_ori_n37_), .C(i_0_), .Y(ori_ori_n292_));
  INV        o270(.A(ori_ori_n292_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n293_), .B(ori_ori_n47_), .Y(ori_ori_n294_));
  NOi21      o272(.An(i_5_), .B(i_9_), .Y(ori_ori_n295_));
  NA2        o273(.A(ori_ori_n295_), .B(i_0_), .Y(ori_ori_n296_));
  BUFFER     o274(.A(ori_ori_n126_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n297_), .B(ori_ori_n154_), .Y(ori_ori_n298_));
  NO2        o276(.A(ori_ori_n298_), .B(ori_ori_n296_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n299_), .B(ori_ori_n294_), .Y(ori_ori_n300_));
  NA2        o278(.A(i_9_), .B(i_0_), .Y(ori_ori_n301_));
  NA2        o279(.A(i_0_), .B(i_10_), .Y(ori_ori_n302_));
  NA2        o280(.A(i_11_), .B(i_9_), .Y(ori_ori_n303_));
  NO3        o281(.A(i_12_), .B(ori_ori_n303_), .C(ori_ori_n179_), .Y(ori_ori_n304_));
  AN2        o282(.A(ori_ori_n304_), .B(i_5_), .Y(ori_ori_n305_));
  INV        o283(.A(ori_ori_n305_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n206_), .B(ori_ori_n76_), .Y(ori_ori_n307_));
  NO2        o285(.A(i_6_), .B(ori_ori_n307_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n98_), .B(ori_ori_n70_), .Y(ori_ori_n309_));
  INV        o287(.A(ori_ori_n308_), .Y(ori_ori_n310_));
  NA2        o288(.A(ori_ori_n310_), .B(ori_ori_n306_), .Y(ori_ori_n311_));
  INV        o289(.A(ori_ori_n311_), .Y(ori_ori_n312_));
  NO2        o290(.A(ori_ori_n270_), .B(ori_ori_n309_), .Y(ori_ori_n313_));
  INV        o291(.A(ori_ori_n313_), .Y(ori_ori_n314_));
  NA2        o292(.A(ori_ori_n113_), .B(ori_ori_n339_), .Y(ori_ori_n315_));
  AOI210     o293(.A0(ori_ori_n315_), .A1(ori_ori_n301_), .B0(ori_ori_n95_), .Y(ori_ori_n316_));
  INV        o294(.A(ori_ori_n316_), .Y(ori_ori_n317_));
  NA2        o295(.A(ori_ori_n317_), .B(ori_ori_n314_), .Y(ori_ori_n318_));
  NO3        o296(.A(ori_ori_n302_), .B(ori_ori_n295_), .C(ori_ori_n101_), .Y(ori_ori_n319_));
  AOI220     o297(.A0(ori_ori_n319_), .A1(i_11_), .B0(ori_ori_n169_), .B1(ori_ori_n52_), .Y(ori_ori_n320_));
  NO3        o298(.A(ori_ori_n107_), .B(ori_ori_n134_), .C(i_0_), .Y(ori_ori_n321_));
  OAI210     o299(.A0(ori_ori_n321_), .A1(ori_ori_n53_), .B0(i_13_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n322_), .B(ori_ori_n320_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n162_), .B(ori_ori_n155_), .Y(ori_ori_n324_));
  INV        o302(.A(ori_ori_n324_), .Y(ori_ori_n325_));
  NA3        o303(.A(ori_ori_n135_), .B(ori_ori_n98_), .C(ori_ori_n97_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n326_), .B(ori_ori_n325_), .Y(ori_ori_n327_));
  NO3        o305(.A(ori_ori_n327_), .B(ori_ori_n323_), .C(ori_ori_n318_), .Y(ori_ori_n328_));
  INV        o306(.A(ori_ori_n186_), .Y(ori_ori_n329_));
  NA2        o307(.A(ori_ori_n329_), .B(ori_ori_n105_), .Y(ori_ori_n330_));
  NA2        o308(.A(i_2_), .B(i_10_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n49_), .B(ori_ori_n331_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n332_), .B(ori_ori_n43_), .Y(ori_ori_n333_));
  AOI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n330_), .B0(ori_ori_n50_), .Y(ori_ori_n334_));
  INV        o312(.A(ori_ori_n334_), .Y(ori_ori_n335_));
  NA4        o313(.A(ori_ori_n335_), .B(ori_ori_n328_), .C(ori_ori_n312_), .D(ori_ori_n300_), .Y(ori4));
  INV        o314(.A(i_12_), .Y(ori_ori_n339_));
  INV        o315(.A(ori_ori_n75_), .Y(ori_ori_n340_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NOi21      m016(.An(i_12_), .B(i_13_), .Y(mai_mai_n39_));
  INV        m017(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NAi31      m018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n41_));
  INV        m019(.A(mai_mai_n35_), .Y(mai1));
  INV        m020(.A(i_11_), .Y(mai_mai_n43_));
  NO2        m021(.A(mai_mai_n43_), .B(i_6_), .Y(mai_mai_n44_));
  INV        m022(.A(i_2_), .Y(mai_mai_n45_));
  NA2        m023(.A(i_0_), .B(i_3_), .Y(mai_mai_n46_));
  INV        m024(.A(i_5_), .Y(mai_mai_n47_));
  NO2        m025(.A(i_7_), .B(i_10_), .Y(mai_mai_n48_));
  AOI210     m026(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n48_), .Y(mai_mai_n49_));
  OAI210     m027(.A0(mai_mai_n49_), .A1(i_3_), .B0(mai_mai_n47_), .Y(mai_mai_n50_));
  AOI210     m028(.A0(mai_mai_n50_), .A1(mai_mai_n46_), .B0(mai_mai_n45_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_0_), .B(i_2_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_7_), .B(i_9_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(mai_mai_n52_), .Y(mai_mai_n54_));
  NA2        m032(.A(mai_mai_n51_), .B(mai_mai_n44_), .Y(mai_mai_n55_));
  NA3        m033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n56_));
  NO2        m034(.A(i_1_), .B(i_6_), .Y(mai_mai_n57_));
  NA2        m035(.A(i_8_), .B(i_7_), .Y(mai_mai_n58_));
  OAI210     m036(.A0(mai_mai_n58_), .A1(mai_mai_n57_), .B0(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n60_));
  NAi21      m038(.An(i_2_), .B(i_7_), .Y(mai_mai_n61_));
  INV        m039(.A(i_1_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n62_), .B(i_6_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n61_), .B(mai_mai_n31_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n60_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n49_), .B(i_2_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n67_));
  NA2        m045(.A(i_1_), .B(i_6_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n25_), .Y(mai_mai_n69_));
  INV        m047(.A(i_0_), .Y(mai_mai_n70_));
  NAi21      m048(.An(i_5_), .B(i_10_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_5_), .B(i_9_), .Y(mai_mai_n72_));
  AOI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n71_), .B0(mai_mai_n70_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n69_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n74_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n65_), .B0(i_0_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_12_), .B(i_5_), .Y(mai_mai_n77_));
  NO2        m055(.A(i_3_), .B(i_9_), .Y(mai_mai_n78_));
  NO2        m056(.A(i_3_), .B(i_7_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n78_), .B(mai_mai_n62_), .Y(mai_mai_n80_));
  INV        m058(.A(i_6_), .Y(mai_mai_n81_));
  NA2        m059(.A(mai_mai_n80_), .B(i_2_), .Y(mai_mai_n82_));
  NAi21      m060(.An(i_6_), .B(i_10_), .Y(mai_mai_n83_));
  NA2        m061(.A(i_6_), .B(i_9_), .Y(mai_mai_n84_));
  AOI210     m062(.A0(mai_mai_n84_), .A1(mai_mai_n83_), .B0(mai_mai_n62_), .Y(mai_mai_n85_));
  NA2        m063(.A(i_2_), .B(i_6_), .Y(mai_mai_n86_));
  NO3        m064(.A(mai_mai_n86_), .B(mai_mai_n48_), .C(mai_mai_n25_), .Y(mai_mai_n87_));
  NO2        m065(.A(mai_mai_n87_), .B(mai_mai_n85_), .Y(mai_mai_n88_));
  AOI210     m066(.A0(mai_mai_n88_), .A1(mai_mai_n82_), .B0(mai_mai_n77_), .Y(mai_mai_n89_));
  NAi21      m067(.An(i_6_), .B(i_11_), .Y(mai_mai_n90_));
  INV        m068(.A(i_7_), .Y(mai_mai_n91_));
  NO2        m069(.A(i_0_), .B(i_5_), .Y(mai_mai_n92_));
  NAi21      m070(.An(i_7_), .B(i_11_), .Y(mai_mai_n93_));
  NO3        m071(.A(mai_mai_n93_), .B(mai_mai_n83_), .C(mai_mai_n52_), .Y(mai_mai_n94_));
  AN2        m072(.A(i_2_), .B(i_10_), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n95_), .B(i_7_), .Y(mai_mai_n96_));
  OR2        m074(.A(mai_mai_n77_), .B(mai_mai_n57_), .Y(mai_mai_n97_));
  NO3        m075(.A(i_7_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n98_));
  NA2        m076(.A(i_12_), .B(i_7_), .Y(mai_mai_n99_));
  NO2        m077(.A(mai_mai_n62_), .B(mai_mai_n26_), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n100_), .B(i_0_), .Y(mai_mai_n101_));
  NA2        m079(.A(i_11_), .B(i_12_), .Y(mai_mai_n102_));
  OAI210     m080(.A0(mai_mai_n101_), .A1(mai_mai_n99_), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n98_), .Y(mai_mai_n104_));
  NAi21      m082(.An(mai_mai_n94_), .B(mai_mai_n104_), .Y(mai_mai_n105_));
  NOi21      m083(.An(i_1_), .B(i_5_), .Y(mai_mai_n106_));
  NA2        m084(.A(mai_mai_n106_), .B(i_11_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n91_), .B(mai_mai_n37_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n109_));
  NA2        m087(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n110_), .B(mai_mai_n45_), .Y(mai_mai_n111_));
  NA2        m089(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n112_));
  NAi21      m090(.An(i_3_), .B(i_8_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n113_), .B(mai_mai_n61_), .Y(mai_mai_n114_));
  NOi31      m092(.An(mai_mai_n114_), .B(mai_mai_n112_), .C(mai_mai_n111_), .Y(mai_mai_n115_));
  NO2        m093(.A(i_1_), .B(mai_mai_n81_), .Y(mai_mai_n116_));
  NO2        m094(.A(i_6_), .B(i_5_), .Y(mai_mai_n117_));
  OAI220     m095(.A0(mai_mai_n46_), .A1(mai_mai_n93_), .B0(mai_mai_n115_), .B1(mai_mai_n107_), .Y(mai_mai_n118_));
  NO3        m096(.A(mai_mai_n118_), .B(mai_mai_n105_), .C(mai_mai_n89_), .Y(mai_mai_n119_));
  NA3        m097(.A(mai_mai_n119_), .B(mai_mai_n76_), .C(mai_mai_n55_), .Y(mai2));
  NO2        m098(.A(mai_mai_n62_), .B(mai_mai_n37_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n773_), .B(mai_mai_n121_), .Y(mai_mai_n122_));
  NA4        m100(.A(mai_mai_n122_), .B(mai_mai_n74_), .C(mai_mai_n66_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m101(.A(i_8_), .B(i_7_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(i_6_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_12_), .B(i_13_), .Y(mai_mai_n126_));
  NAi21      m104(.An(i_5_), .B(i_11_), .Y(mai_mai_n127_));
  NOi21      m105(.An(mai_mai_n126_), .B(mai_mai_n127_), .Y(mai_mai_n128_));
  NO2        m106(.A(i_0_), .B(i_1_), .Y(mai_mai_n129_));
  NA2        m107(.A(i_2_), .B(i_3_), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n130_), .B(i_4_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n131_), .B(mai_mai_n128_), .Y(mai_mai_n132_));
  AN2        m110(.A(mai_mai_n126_), .B(mai_mai_n78_), .Y(mai_mai_n133_));
  NA2        m111(.A(i_1_), .B(i_5_), .Y(mai_mai_n134_));
  NO3        m112(.A(mai_mai_n778_), .B(mai_mai_n134_), .C(mai_mai_n26_), .Y(mai_mai_n135_));
  OR2        m113(.A(i_0_), .B(i_1_), .Y(mai_mai_n136_));
  NO3        m114(.A(mai_mai_n136_), .B(mai_mai_n77_), .C(i_13_), .Y(mai_mai_n137_));
  NAi32      m115(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n138_));
  NAi21      m116(.An(mai_mai_n138_), .B(mai_mai_n137_), .Y(mai_mai_n139_));
  NOi21      m117(.An(i_4_), .B(i_10_), .Y(mai_mai_n140_));
  NA2        m118(.A(mai_mai_n140_), .B(mai_mai_n39_), .Y(mai_mai_n141_));
  NO2        m119(.A(i_3_), .B(i_5_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n137_), .B(mai_mai_n135_), .Y(mai_mai_n143_));
  AOI210     m121(.A0(mai_mai_n143_), .A1(mai_mai_n132_), .B0(mai_mai_n125_), .Y(mai_mai_n144_));
  NOi21      m122(.An(i_4_), .B(i_9_), .Y(mai_mai_n145_));
  NOi21      m123(.An(i_11_), .B(i_13_), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NO2        m125(.A(i_4_), .B(i_5_), .Y(mai_mai_n148_));
  NAi21      m126(.An(i_12_), .B(i_11_), .Y(mai_mai_n149_));
  NO2        m127(.A(mai_mai_n149_), .B(i_13_), .Y(mai_mai_n150_));
  NO2        m128(.A(mai_mai_n70_), .B(mai_mai_n62_), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n152_));
  NAi31      m130(.An(mai_mai_n152_), .B(mai_mai_n133_), .C(i_11_), .Y(mai_mai_n153_));
  NA2        m131(.A(i_3_), .B(i_5_), .Y(mai_mai_n154_));
  AOI210     m132(.A0(mai_mai_n147_), .A1(mai_mai_n153_), .B0(mai_mai_n62_), .Y(mai_mai_n155_));
  NO2        m133(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n156_));
  NO2        m134(.A(i_13_), .B(i_10_), .Y(mai_mai_n157_));
  NA3        m135(.A(mai_mai_n157_), .B(mai_mai_n156_), .C(mai_mai_n43_), .Y(mai_mai_n158_));
  NO2        m136(.A(i_2_), .B(i_1_), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n159_), .B(i_3_), .Y(mai_mai_n160_));
  NAi21      m138(.An(i_4_), .B(i_12_), .Y(mai_mai_n161_));
  NO3        m139(.A(mai_mai_n161_), .B(mai_mai_n158_), .C(mai_mai_n25_), .Y(mai_mai_n162_));
  NO2        m140(.A(mai_mai_n162_), .B(mai_mai_n155_), .Y(mai_mai_n163_));
  INV        m141(.A(i_8_), .Y(mai_mai_n164_));
  NA2        m142(.A(i_8_), .B(i_6_), .Y(mai_mai_n165_));
  NO3        m143(.A(i_3_), .B(mai_mai_n81_), .C(mai_mai_n47_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n166_), .B(i_7_), .Y(mai_mai_n167_));
  NO3        m145(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n168_));
  NA3        m146(.A(mai_mai_n168_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n169_));
  NO3        m147(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n169_), .B(mai_mai_n167_), .Y(mai_mai_n171_));
  NO3        m149(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n172_));
  NA2        m150(.A(mai_mai_n172_), .B(mai_mai_n39_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n92_), .B(mai_mai_n57_), .Y(mai_mai_n174_));
  NO2        m152(.A(i_13_), .B(i_9_), .Y(mai_mai_n175_));
  NA3        m153(.A(mai_mai_n175_), .B(i_6_), .C(mai_mai_n164_), .Y(mai_mai_n176_));
  NAi21      m154(.An(i_12_), .B(i_3_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n43_), .B(i_5_), .Y(mai_mai_n178_));
  OAI210     m156(.A0(mai_mai_n57_), .A1(mai_mai_n173_), .B0(mai_mai_n176_), .Y(mai_mai_n179_));
  AOI210     m157(.A0(mai_mai_n179_), .A1(i_7_), .B0(mai_mai_n171_), .Y(mai_mai_n180_));
  OAI220     m158(.A0(mai_mai_n180_), .A1(i_4_), .B0(mai_mai_n165_), .B1(mai_mai_n163_), .Y(mai_mai_n181_));
  NAi21      m159(.An(i_12_), .B(i_7_), .Y(mai_mai_n182_));
  NA3        m160(.A(i_13_), .B(mai_mai_n164_), .C(i_10_), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n183_), .B(mai_mai_n182_), .Y(mai_mai_n184_));
  NA2        m162(.A(i_0_), .B(i_5_), .Y(mai_mai_n185_));
  INV        m163(.A(mai_mai_n160_), .Y(mai_mai_n186_));
  NAi31      m164(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n187_));
  NO2        m165(.A(mai_mai_n45_), .B(mai_mai_n62_), .Y(mai_mai_n188_));
  INV        m166(.A(i_13_), .Y(mai_mai_n189_));
  NO2        m167(.A(i_12_), .B(mai_mai_n189_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n190_), .B(mai_mai_n166_), .Y(mai_mai_n191_));
  INV        m169(.A(mai_mai_n191_), .Y(mai_mai_n192_));
  AOI220     m170(.A0(mai_mai_n192_), .A1(mai_mai_n124_), .B0(mai_mai_n186_), .B1(mai_mai_n184_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n154_), .B(i_4_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(i_10_), .Y(mai_mai_n195_));
  OR2        m173(.A(i_8_), .B(i_7_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n52_), .B(i_1_), .Y(mai_mai_n197_));
  INV        m175(.A(i_12_), .Y(mai_mai_n198_));
  NO3        m176(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n199_));
  NA2        m177(.A(i_2_), .B(i_1_), .Y(mai_mai_n200_));
  NO3        m178(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n201_));
  NAi21      m179(.An(i_4_), .B(i_3_), .Y(mai_mai_n202_));
  NO2        m180(.A(i_0_), .B(i_6_), .Y(mai_mai_n203_));
  NOi41      m181(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n204_));
  NO2        m182(.A(i_11_), .B(mai_mai_n189_), .Y(mai_mai_n205_));
  NAi21      m183(.An(i_3_), .B(i_7_), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n198_), .B(i_9_), .Y(mai_mai_n207_));
  OR3        m185(.A(mai_mai_n207_), .B(mai_mai_n206_), .C(i_1_), .Y(mai_mai_n208_));
  NO2        m186(.A(i_12_), .B(i_3_), .Y(mai_mai_n209_));
  INV        m187(.A(mai_mai_n208_), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n210_), .B(mai_mai_n205_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n196_), .B(mai_mai_n37_), .Y(mai_mai_n212_));
  NA2        m190(.A(i_12_), .B(i_6_), .Y(mai_mai_n213_));
  OR2        m191(.A(i_13_), .B(i_9_), .Y(mai_mai_n214_));
  NO3        m192(.A(mai_mai_n214_), .B(mai_mai_n213_), .C(mai_mai_n47_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n202_), .B(i_2_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n205_), .B(i_9_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n62_), .B(mai_mai_n217_), .Y(mai_mai_n218_));
  NA2        m196(.A(i_2_), .B(mai_mai_n62_), .Y(mai_mai_n219_));
  NO3        m197(.A(i_11_), .B(mai_mai_n189_), .C(mai_mai_n25_), .Y(mai_mai_n220_));
  NO2        m198(.A(mai_mai_n206_), .B(i_8_), .Y(mai_mai_n221_));
  NA2        m199(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  NA3        m200(.A(i_3_), .B(mai_mai_n212_), .C(mai_mai_n190_), .Y(mai_mai_n223_));
  AOI210     m201(.A0(mai_mai_n223_), .A1(mai_mai_n222_), .B0(mai_mai_n219_), .Y(mai_mai_n224_));
  AOI210     m202(.A0(mai_mai_n218_), .A1(mai_mai_n212_), .B0(mai_mai_n224_), .Y(mai_mai_n225_));
  NA3        m203(.A(mai_mai_n225_), .B(mai_mai_n211_), .C(mai_mai_n193_), .Y(mai_mai_n226_));
  NO3        m204(.A(i_12_), .B(mai_mai_n189_), .C(mai_mai_n37_), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n227_), .Y(mai_mai_n228_));
  INV        m206(.A(i_8_), .Y(mai_mai_n229_));
  NO3        m207(.A(i_0_), .B(mai_mai_n45_), .C(i_1_), .Y(mai_mai_n230_));
  AOI220     m208(.A0(mai_mai_n230_), .A1(mai_mai_n166_), .B0(mai_mai_n142_), .B1(mai_mai_n197_), .Y(mai_mai_n231_));
  NO2        m209(.A(mai_mai_n231_), .B(mai_mai_n229_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n200_), .B(i_0_), .Y(mai_mai_n233_));
  NO2        m211(.A(i_6_), .B(i_0_), .Y(mai_mai_n234_));
  NA2        m212(.A(i_0_), .B(i_1_), .Y(mai_mai_n235_));
  NO2        m213(.A(mai_mai_n235_), .B(i_2_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n58_), .B(i_6_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  OAI210     m216(.A0(i_3_), .A1(mai_mai_n125_), .B0(mai_mai_n238_), .Y(mai_mai_n239_));
  NO3        m217(.A(mai_mai_n239_), .B(mai_mai_n234_), .C(mai_mai_n232_), .Y(mai_mai_n240_));
  NO2        m218(.A(i_3_), .B(i_10_), .Y(mai_mai_n241_));
  NA3        m219(.A(mai_mai_n241_), .B(mai_mai_n39_), .C(mai_mai_n43_), .Y(mai_mai_n242_));
  NA2        m220(.A(i_1_), .B(i_7_), .Y(mai_mai_n243_));
  AN2        m221(.A(i_3_), .B(i_10_), .Y(mai_mai_n244_));
  NA2        m222(.A(mai_mai_n150_), .B(mai_mai_n148_), .Y(mai_mai_n245_));
  OR2        m223(.A(mai_mai_n243_), .B(mai_mai_n242_), .Y(mai_mai_n246_));
  OAI220     m224(.A0(mai_mai_n246_), .A1(i_6_), .B0(mai_mai_n240_), .B1(mai_mai_n228_), .Y(mai_mai_n247_));
  NO4        m225(.A(mai_mai_n247_), .B(mai_mai_n226_), .C(mai_mai_n181_), .D(mai_mai_n144_), .Y(mai_mai_n248_));
  NO3        m226(.A(mai_mai_n43_), .B(i_13_), .C(i_9_), .Y(mai_mai_n249_));
  NO3        m227(.A(i_6_), .B(mai_mai_n164_), .C(i_7_), .Y(mai_mai_n250_));
  NO2        m228(.A(i_2_), .B(i_3_), .Y(mai_mai_n251_));
  OR2        m229(.A(i_0_), .B(i_5_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n185_), .B(mai_mai_n252_), .Y(mai_mai_n253_));
  NA3        m231(.A(mai_mai_n771_), .B(mai_mai_n251_), .C(i_1_), .Y(mai_mai_n254_));
  INV        m232(.A(i_6_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n136_), .B(mai_mai_n45_), .Y(mai_mai_n256_));
  INV        m234(.A(mai_mai_n256_), .Y(mai_mai_n257_));
  NA3        m235(.A(mai_mai_n257_), .B(mai_mai_n200_), .C(mai_mai_n254_), .Y(mai_mai_n258_));
  OAI210     m236(.A0(mai_mai_n258_), .A1(mai_mai_n250_), .B0(i_4_), .Y(mai_mai_n259_));
  NO2        m237(.A(i_12_), .B(i_10_), .Y(mai_mai_n260_));
  NOi21      m238(.An(i_5_), .B(i_0_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n769_), .B(mai_mai_n113_), .Y(mai_mai_n262_));
  INV        m240(.A(mai_mai_n262_), .Y(mai_mai_n263_));
  NO2        m241(.A(i_6_), .B(i_8_), .Y(mai_mai_n264_));
  NO2        m242(.A(i_1_), .B(i_7_), .Y(mai_mai_n265_));
  NA3        m243(.A(mai_mai_n264_), .B(i_4_), .C(i_5_), .Y(mai_mai_n266_));
  NA3        m244(.A(mai_mai_n266_), .B(mai_mai_n263_), .C(mai_mai_n259_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(i_7_), .A1(i_2_), .B0(i_6_), .Y(mai_mai_n268_));
  NA2        m246(.A(i_0_), .B(mai_mai_n117_), .Y(mai_mai_n269_));
  AOI210     m247(.A0(mai_mai_n164_), .A1(mai_mai_n253_), .B0(mai_mai_n141_), .Y(mai_mai_n270_));
  AOI210     m248(.A0(mai_mai_n267_), .A1(mai_mai_n249_), .B0(mai_mai_n270_), .Y(mai_mai_n271_));
  NOi32      m249(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n272_));
  INV        m250(.A(mai_mai_n272_), .Y(mai_mai_n273_));
  NAi21      m251(.An(i_1_), .B(i_5_), .Y(mai_mai_n274_));
  NA2        m252(.A(mai_mai_n274_), .B(i_0_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n275_), .B(mai_mai_n25_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(mai_mai_n138_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n138_), .B(mai_mai_n136_), .Y(mai_mai_n278_));
  NOi32      m256(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n279_), .B(mai_mai_n45_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n280_), .B(i_0_), .Y(mai_mai_n281_));
  OR2        m259(.A(mai_mai_n281_), .B(mai_mai_n278_), .Y(mai_mai_n282_));
  NO2        m260(.A(i_1_), .B(mai_mai_n91_), .Y(mai_mai_n283_));
  NAi21      m261(.An(i_3_), .B(i_4_), .Y(mai_mai_n284_));
  NO2        m262(.A(mai_mai_n284_), .B(i_9_), .Y(mai_mai_n285_));
  NA2        m263(.A(i_7_), .B(mai_mai_n285_), .Y(mai_mai_n286_));
  NA2        m264(.A(i_2_), .B(i_7_), .Y(mai_mai_n287_));
  NO2        m265(.A(mai_mai_n284_), .B(i_10_), .Y(mai_mai_n288_));
  NA3        m266(.A(mai_mai_n288_), .B(mai_mai_n287_), .C(mai_mai_n203_), .Y(mai_mai_n289_));
  AOI210     m267(.A0(mai_mai_n289_), .A1(mai_mai_n286_), .B0(mai_mai_n156_), .Y(mai_mai_n290_));
  AOI210     m268(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n291_));
  OAI210     m269(.A0(mai_mai_n291_), .A1(mai_mai_n159_), .B0(mai_mai_n288_), .Y(mai_mai_n292_));
  AOI220     m270(.A0(mai_mai_n288_), .A1(mai_mai_n265_), .B0(mai_mai_n199_), .B1(mai_mai_n159_), .Y(mai_mai_n293_));
  AOI210     m271(.A0(mai_mai_n293_), .A1(mai_mai_n292_), .B0(i_5_), .Y(mai_mai_n294_));
  NO4        m272(.A(mai_mai_n294_), .B(mai_mai_n290_), .C(mai_mai_n282_), .D(mai_mai_n277_), .Y(mai_mai_n295_));
  NO2        m273(.A(mai_mai_n295_), .B(mai_mai_n273_), .Y(mai_mai_n296_));
  AN2        m274(.A(i_12_), .B(i_5_), .Y(mai_mai_n297_));
  NA2        m275(.A(i_3_), .B(mai_mai_n297_), .Y(mai_mai_n298_));
  NO2        m276(.A(i_11_), .B(i_6_), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n136_), .B(mai_mai_n298_), .Y(mai_mai_n300_));
  NO2        m278(.A(mai_mai_n202_), .B(i_5_), .Y(mai_mai_n301_));
  NO2        m279(.A(i_5_), .B(i_10_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n300_), .B(i_9_), .Y(mai_mai_n303_));
  NO2        m281(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n304_));
  NO3        m282(.A(mai_mai_n81_), .B(mai_mai_n47_), .C(i_9_), .Y(mai_mai_n305_));
  NO2        m283(.A(i_11_), .B(i_12_), .Y(mai_mai_n306_));
  NA2        m284(.A(mai_mai_n302_), .B(mai_mai_n198_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n91_), .B(mai_mai_n187_), .Y(mai_mai_n308_));
  NO2        m286(.A(i_13_), .B(mai_mai_n200_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n308_), .B(mai_mai_n309_), .Y(mai_mai_n310_));
  NA3        m288(.A(mai_mai_n310_), .B(mai_mai_n132_), .C(mai_mai_n303_), .Y(mai_mai_n311_));
  NO2        m289(.A(i_0_), .B(i_11_), .Y(mai_mai_n312_));
  AN2        m290(.A(i_1_), .B(i_6_), .Y(mai_mai_n313_));
  OR2        m291(.A(i_13_), .B(i_10_), .Y(mai_mai_n314_));
  NO2        m292(.A(mai_mai_n147_), .B(mai_mai_n108_), .Y(mai_mai_n315_));
  BUFFER     m293(.A(mai_mai_n183_), .Y(mai_mai_n316_));
  NO2        m294(.A(mai_mai_n91_), .B(mai_mai_n25_), .Y(mai_mai_n317_));
  NA2        m295(.A(mai_mai_n227_), .B(mai_mai_n317_), .Y(mai_mai_n318_));
  OAI220     m296(.A0(i_6_), .A1(mai_mai_n316_), .B0(mai_mai_n318_), .B1(mai_mai_n92_), .Y(mai_mai_n319_));
  INV        m297(.A(mai_mai_n319_), .Y(mai_mai_n320_));
  NO2        m298(.A(mai_mai_n320_), .B(mai_mai_n26_), .Y(mai_mai_n321_));
  INV        m299(.A(mai_mai_n254_), .Y(mai_mai_n322_));
  AOI220     m300(.A0(mai_mai_n237_), .A1(mai_mai_n230_), .B0(mai_mai_n233_), .B1(i_7_), .Y(mai_mai_n323_));
  NO2        m301(.A(mai_mai_n323_), .B(i_5_), .Y(mai_mai_n324_));
  NO2        m302(.A(i_2_), .B(mai_mai_n229_), .Y(mai_mai_n325_));
  NO3        m303(.A(mai_mai_n325_), .B(mai_mai_n324_), .C(mai_mai_n322_), .Y(mai_mai_n326_));
  NA2        m304(.A(mai_mai_n166_), .B(i_1_), .Y(mai_mai_n327_));
  NO2        m305(.A(mai_mai_n327_), .B(i_8_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n63_), .B(i_2_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n237_), .B(mai_mai_n197_), .Y(mai_mai_n330_));
  OAI220     m308(.A0(mai_mai_n330_), .A1(mai_mai_n154_), .B0(mai_mai_n329_), .B1(mai_mai_n774_), .Y(mai_mai_n331_));
  NA3        m309(.A(mai_mai_n265_), .B(mai_mai_n264_), .C(i_5_), .Y(mai_mai_n332_));
  INV        m310(.A(mai_mai_n332_), .Y(mai_mai_n333_));
  NO3        m311(.A(mai_mai_n333_), .B(mai_mai_n331_), .C(mai_mai_n328_), .Y(mai_mai_n334_));
  AOI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n326_), .B0(mai_mai_n217_), .Y(mai_mai_n335_));
  NO4        m313(.A(mai_mai_n335_), .B(mai_mai_n321_), .C(mai_mai_n311_), .D(mai_mai_n296_), .Y(mai_mai_n336_));
  NO2        m314(.A(mai_mai_n70_), .B(i_13_), .Y(mai_mai_n337_));
  NO2        m315(.A(i_10_), .B(i_9_), .Y(mai_mai_n338_));
  NAi21      m316(.An(i_12_), .B(i_8_), .Y(mai_mai_n339_));
  NO2        m317(.A(mai_mai_n339_), .B(i_3_), .Y(mai_mai_n340_));
  NO3        m318(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n213_), .B(mai_mai_n90_), .Y(mai_mai_n342_));
  NA2        m320(.A(i_8_), .B(i_9_), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n227_), .B(mai_mai_n174_), .Y(mai_mai_n344_));
  NO2        m322(.A(mai_mai_n344_), .B(mai_mai_n343_), .Y(mai_mai_n345_));
  NO3        m323(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n346_));
  NA3        m324(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n100_), .B(mai_mai_n23_), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n349_), .B(mai_mai_n345_), .Y(mai_mai_n350_));
  OR2        m328(.A(mai_mai_n176_), .B(mai_mai_n195_), .Y(mai_mai_n351_));
  NO2        m329(.A(i_2_), .B(i_13_), .Y(mai_mai_n352_));
  NO3        m330(.A(i_4_), .B(mai_mai_n47_), .C(i_8_), .Y(mai_mai_n353_));
  NO2        m331(.A(i_6_), .B(i_7_), .Y(mai_mai_n354_));
  NO2        m332(.A(i_11_), .B(i_1_), .Y(mai_mai_n355_));
  NAi31      m333(.An(i_11_), .B(i_2_), .C(i_0_), .Y(mai_mai_n356_));
  NO2        m334(.A(mai_mai_n314_), .B(i_6_), .Y(mai_mai_n357_));
  NA2        m335(.A(mai_mai_n357_), .B(i_1_), .Y(mai_mai_n358_));
  NO2        m336(.A(mai_mai_n358_), .B(mai_mai_n356_), .Y(mai_mai_n359_));
  NO2        m337(.A(i_6_), .B(i_10_), .Y(mai_mai_n360_));
  INV        m338(.A(mai_mai_n359_), .Y(mai_mai_n361_));
  NAi21      m339(.An(mai_mai_n183_), .B(mai_mai_n306_), .Y(mai_mai_n362_));
  NA2        m340(.A(mai_mai_n265_), .B(mai_mai_n185_), .Y(mai_mai_n363_));
  NO2        m341(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n364_));
  NA3        m342(.A(i_6_), .B(mai_mai_n364_), .C(mai_mai_n124_), .Y(mai_mai_n365_));
  OR3        m343(.A(mai_mai_n769_), .B(mai_mai_n38_), .C(mai_mai_n45_), .Y(mai_mai_n366_));
  OAI220     m344(.A0(mai_mai_n366_), .A1(mai_mai_n365_), .B0(mai_mai_n363_), .B1(mai_mai_n362_), .Y(mai_mai_n367_));
  NA2        m345(.A(mai_mai_n249_), .B(mai_mai_n199_), .Y(mai_mai_n368_));
  NO2        m346(.A(mai_mai_n368_), .B(mai_mai_n329_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n369_), .B(mai_mai_n367_), .Y(mai_mai_n370_));
  NA4        m348(.A(mai_mai_n370_), .B(mai_mai_n361_), .C(mai_mai_n351_), .D(mai_mai_n350_), .Y(mai_mai_n371_));
  AN2        m349(.A(i_5_), .B(mai_mai_n341_), .Y(mai_mai_n372_));
  OAI210     m350(.A0(mai_mai_n70_), .A1(mai_mai_n195_), .B0(mai_mai_n245_), .Y(mai_mai_n373_));
  AOI220     m351(.A0(mai_mai_n373_), .A1(mai_mai_n255_), .B0(mai_mai_n372_), .B1(i_3_), .Y(mai_mai_n374_));
  NA3        m352(.A(mai_mai_n337_), .B(i_1_), .C(i_2_), .Y(mai_mai_n375_));
  INV        m353(.A(mai_mai_n375_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n297_), .B(mai_mai_n189_), .Y(mai_mai_n377_));
  NA2        m355(.A(mai_mai_n272_), .B(mai_mai_n70_), .Y(mai_mai_n378_));
  NA2        m356(.A(i_7_), .B(mai_mai_n279_), .Y(mai_mai_n379_));
  AO210      m357(.A0(mai_mai_n378_), .A1(mai_mai_n377_), .B0(mai_mai_n379_), .Y(mai_mai_n380_));
  NO2        m358(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n381_));
  NAi41      m359(.An(mai_mai_n378_), .B(mai_mai_n360_), .C(mai_mai_n381_), .D(mai_mai_n45_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n382_), .B(mai_mai_n380_), .Y(mai_mai_n383_));
  AOI210     m361(.A0(mai_mai_n376_), .A1(mai_mai_n172_), .B0(mai_mai_n383_), .Y(mai_mai_n384_));
  NO2        m362(.A(i_7_), .B(mai_mai_n169_), .Y(mai_mai_n385_));
  AOI220     m363(.A0(i_3_), .A1(mai_mai_n385_), .B0(mai_mai_n766_), .B1(mai_mai_n315_), .Y(mai_mai_n386_));
  NA3        m364(.A(mai_mai_n386_), .B(mai_mai_n384_), .C(mai_mai_n374_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n301_), .B(mai_mai_n236_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n298_), .B(mai_mai_n388_), .Y(mai_mai_n389_));
  NO2        m367(.A(i_12_), .B(mai_mai_n164_), .Y(mai_mai_n390_));
  OAI210     m368(.A0(mai_mai_n250_), .A1(mai_mai_n390_), .B0(mai_mai_n389_), .Y(mai_mai_n391_));
  NO2        m369(.A(i_8_), .B(i_7_), .Y(mai_mai_n392_));
  INV        m370(.A(mai_mai_n188_), .Y(mai_mai_n393_));
  NA2        m371(.A(mai_mai_n43_), .B(i_10_), .Y(mai_mai_n394_));
  NO2        m372(.A(mai_mai_n394_), .B(i_6_), .Y(mai_mai_n395_));
  NA3        m373(.A(mai_mai_n395_), .B(i_3_), .C(mai_mai_n392_), .Y(mai_mai_n396_));
  NA2        m374(.A(i_5_), .B(mai_mai_n203_), .Y(mai_mai_n397_));
  INV        m375(.A(mai_mai_n397_), .Y(mai_mai_n398_));
  NA2        m376(.A(mai_mai_n398_), .B(mai_mai_n212_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n242_), .B(mai_mai_n152_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n244_), .B(mai_mai_n148_), .Y(mai_mai_n401_));
  NA2        m379(.A(mai_mai_n780_), .B(mai_mai_n251_), .Y(mai_mai_n402_));
  NA2        m380(.A(mai_mai_n402_), .B(mai_mai_n401_), .Y(mai_mai_n403_));
  OAI210     m381(.A0(mai_mai_n403_), .A1(mai_mai_n400_), .B0(mai_mai_n346_), .Y(mai_mai_n404_));
  NA4        m382(.A(mai_mai_n404_), .B(mai_mai_n399_), .C(mai_mai_n396_), .D(mai_mai_n391_), .Y(mai_mai_n405_));
  NA3        m383(.A(mai_mai_n185_), .B(mai_mai_n68_), .C(mai_mai_n43_), .Y(mai_mai_n406_));
  NA2        m384(.A(mai_mai_n227_), .B(mai_mai_n79_), .Y(mai_mai_n407_));
  AOI210     m385(.A0(mai_mai_n406_), .A1(mai_mai_n269_), .B0(mai_mai_n407_), .Y(mai_mai_n408_));
  NA2        m386(.A(mai_mai_n390_), .B(mai_mai_n220_), .Y(mai_mai_n409_));
  NO2        m387(.A(mai_mai_n91_), .B(mai_mai_n409_), .Y(mai_mai_n410_));
  NO2        m388(.A(mai_mai_n410_), .B(mai_mai_n408_), .Y(mai_mai_n411_));
  NO4        m389(.A(i_1_), .B(mai_mai_n41_), .C(i_2_), .D(mai_mai_n47_), .Y(mai_mai_n412_));
  NO3        m390(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n413_));
  NO2        m391(.A(mai_mai_n196_), .B(mai_mai_n36_), .Y(mai_mai_n414_));
  AN2        m392(.A(mai_mai_n414_), .B(mai_mai_n413_), .Y(mai_mai_n415_));
  OA210      m393(.A0(mai_mai_n415_), .A1(mai_mai_n412_), .B0(mai_mai_n272_), .Y(mai_mai_n416_));
  NO2        m394(.A(mai_mai_n314_), .B(i_1_), .Y(mai_mai_n417_));
  NOi31      m395(.An(mai_mai_n417_), .B(mai_mai_n342_), .C(mai_mai_n70_), .Y(mai_mai_n418_));
  AN4        m396(.A(mai_mai_n418_), .B(mai_mai_n124_), .C(mai_mai_n364_), .D(i_2_), .Y(mai_mai_n419_));
  NO2        m397(.A(mai_mai_n419_), .B(mai_mai_n416_), .Y(mai_mai_n420_));
  NOi21      m398(.An(i_10_), .B(i_6_), .Y(mai_mai_n421_));
  NO2        m399(.A(mai_mai_n99_), .B(mai_mai_n23_), .Y(mai_mai_n422_));
  INV        m400(.A(mai_mai_n250_), .Y(mai_mai_n423_));
  AOI220     m401(.A0(mai_mai_n423_), .A1(mai_mai_n330_), .B0(mai_mai_n147_), .B1(mai_mai_n153_), .Y(mai_mai_n424_));
  INV        m402(.A(mai_mai_n424_), .Y(mai_mai_n425_));
  INV        m403(.A(mai_mai_n251_), .Y(mai_mai_n426_));
  NO2        m404(.A(i_12_), .B(mai_mai_n81_), .Y(mai_mai_n427_));
  NA2        m405(.A(mai_mai_n427_), .B(mai_mai_n220_), .Y(mai_mai_n428_));
  NA3        m406(.A(mai_mai_n299_), .B(mai_mai_n227_), .C(mai_mai_n185_), .Y(mai_mai_n429_));
  AOI210     m407(.A0(mai_mai_n429_), .A1(mai_mai_n428_), .B0(mai_mai_n426_), .Y(mai_mai_n430_));
  NO3        m408(.A(i_4_), .B(mai_mai_n268_), .C(mai_mai_n242_), .Y(mai_mai_n431_));
  OR2        m409(.A(i_5_), .B(mai_mai_n313_), .Y(mai_mai_n432_));
  NO2        m410(.A(mai_mai_n432_), .B(mai_mai_n362_), .Y(mai_mai_n433_));
  NO3        m411(.A(mai_mai_n433_), .B(mai_mai_n431_), .C(mai_mai_n430_), .Y(mai_mai_n434_));
  NA4        m412(.A(mai_mai_n434_), .B(mai_mai_n425_), .C(mai_mai_n420_), .D(mai_mai_n411_), .Y(mai_mai_n435_));
  NO4        m413(.A(mai_mai_n435_), .B(mai_mai_n405_), .C(mai_mai_n387_), .D(mai_mai_n371_), .Y(mai_mai_n436_));
  NA4        m414(.A(mai_mai_n436_), .B(mai_mai_n336_), .C(mai_mai_n271_), .D(mai_mai_n248_), .Y(mai7));
  NO2        m415(.A(mai_mai_n93_), .B(mai_mai_n83_), .Y(mai_mai_n438_));
  NA2        m416(.A(mai_mai_n360_), .B(mai_mai_n79_), .Y(mai_mai_n439_));
  NA2        m417(.A(i_11_), .B(mai_mai_n164_), .Y(mai_mai_n440_));
  NO2        m418(.A(mai_mai_n198_), .B(i_4_), .Y(mai_mai_n441_));
  NA2        m419(.A(mai_mai_n441_), .B(i_8_), .Y(mai_mai_n442_));
  INV        m420(.A(i_2_), .Y(mai_mai_n443_));
  INV        m421(.A(mai_mai_n172_), .Y(mai_mai_n444_));
  NO2        m422(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n445_));
  NA2        m423(.A(i_4_), .B(i_8_), .Y(mai_mai_n446_));
  INV        m424(.A(mai_mai_n438_), .Y(mai_mai_n447_));
  OR2        m425(.A(i_6_), .B(i_10_), .Y(mai_mai_n448_));
  NO2        m426(.A(mai_mai_n448_), .B(mai_mai_n23_), .Y(mai_mai_n449_));
  OR3        m427(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n450_));
  NO3        m428(.A(mai_mai_n450_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n451_));
  INV        m429(.A(mai_mai_n170_), .Y(mai_mai_n452_));
  NO2        m430(.A(mai_mai_n451_), .B(mai_mai_n449_), .Y(mai_mai_n453_));
  OA220      m431(.A0(mai_mai_n453_), .A1(mai_mai_n426_), .B0(mai_mai_n764_), .B1(mai_mai_n214_), .Y(mai_mai_n454_));
  AOI210     m432(.A0(mai_mai_n454_), .A1(mai_mai_n447_), .B0(mai_mai_n62_), .Y(mai_mai_n455_));
  NOi21      m433(.An(i_11_), .B(i_7_), .Y(mai_mai_n456_));
  AO210      m434(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n457_), .B(mai_mai_n456_), .Y(mai_mai_n458_));
  NA3        m436(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n459_));
  NAi31      m437(.An(mai_mai_n459_), .B(mai_mai_n182_), .C(i_11_), .Y(mai_mai_n460_));
  NO2        m438(.A(mai_mai_n460_), .B(mai_mai_n62_), .Y(mai_mai_n461_));
  AO210      m439(.A0(i_8_), .A1(mai_mai_n293_), .B0(mai_mai_n40_), .Y(mai_mai_n462_));
  NO3        m440(.A(i_7_), .B(mai_mai_n177_), .C(mai_mai_n440_), .Y(mai_mai_n463_));
  OAI210     m441(.A0(mai_mai_n463_), .A1(mai_mai_n190_), .B0(mai_mai_n62_), .Y(mai_mai_n464_));
  NA2        m442(.A(i_2_), .B(mai_mai_n31_), .Y(mai_mai_n465_));
  OR2        m443(.A(mai_mai_n177_), .B(mai_mai_n93_), .Y(mai_mai_n466_));
  NA2        m444(.A(mai_mai_n466_), .B(mai_mai_n465_), .Y(mai_mai_n467_));
  INV        m445(.A(i_4_), .Y(mai_mai_n468_));
  NA2        m446(.A(mai_mai_n468_), .B(mai_mai_n467_), .Y(mai_mai_n469_));
  NO2        m447(.A(i_1_), .B(i_12_), .Y(mai_mai_n470_));
  NA3        m448(.A(mai_mai_n470_), .B(mai_mai_n95_), .C(mai_mai_n24_), .Y(mai_mai_n471_));
  NA4        m449(.A(mai_mai_n471_), .B(mai_mai_n469_), .C(mai_mai_n464_), .D(mai_mai_n462_), .Y(mai_mai_n472_));
  OAI210     m450(.A0(mai_mai_n472_), .A1(mai_mai_n461_), .B0(i_6_), .Y(mai_mai_n473_));
  NO2        m451(.A(mai_mai_n459_), .B(mai_mai_n93_), .Y(mai_mai_n474_));
  NA2        m452(.A(mai_mai_n474_), .B(mai_mai_n427_), .Y(mai_mai_n475_));
  NO2        m453(.A(i_6_), .B(i_11_), .Y(mai_mai_n476_));
  INV        m454(.A(mai_mai_n475_), .Y(mai_mai_n477_));
  NA3        m455(.A(mai_mai_n392_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n478_));
  NA2        m456(.A(mai_mai_n121_), .B(i_9_), .Y(mai_mai_n479_));
  NA3        m457(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n480_));
  NA3        m458(.A(i_2_), .B(mai_mai_n213_), .C(mai_mai_n43_), .Y(mai_mai_n481_));
  OAI220     m459(.A0(mai_mai_n481_), .A1(mai_mai_n480_), .B0(mai_mai_n479_), .B1(mai_mai_n763_), .Y(mai_mai_n482_));
  AOI210     m460(.A0(mai_mai_n355_), .A1(mai_mai_n317_), .B0(mai_mai_n201_), .Y(mai_mai_n483_));
  NO2        m461(.A(mai_mai_n483_), .B(mai_mai_n443_), .Y(mai_mai_n484_));
  NO2        m462(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n485_));
  NA2        m463(.A(mai_mai_n485_), .B(mai_mai_n24_), .Y(mai_mai_n486_));
  NO2        m464(.A(mai_mai_n486_), .B(mai_mai_n45_), .Y(mai_mai_n487_));
  OR3        m465(.A(mai_mai_n487_), .B(mai_mai_n484_), .C(mai_mai_n482_), .Y(mai_mai_n488_));
  NO2        m466(.A(mai_mai_n488_), .B(mai_mai_n477_), .Y(mai_mai_n489_));
  NO2        m467(.A(mai_mai_n198_), .B(mai_mai_n91_), .Y(mai_mai_n490_));
  NO2        m468(.A(mai_mai_n490_), .B(mai_mai_n456_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n491_), .B(i_1_), .Y(mai_mai_n492_));
  NO2        m470(.A(mai_mai_n492_), .B(mai_mai_n450_), .Y(mai_mai_n493_));
  NA2        m471(.A(mai_mai_n493_), .B(mai_mai_n45_), .Y(mai_mai_n494_));
  NA2        m472(.A(i_3_), .B(mai_mai_n164_), .Y(mai_mai_n495_));
  NO2        m473(.A(mai_mai_n495_), .B(mai_mai_n99_), .Y(mai_mai_n496_));
  AN2        m474(.A(mai_mai_n496_), .B(mai_mai_n395_), .Y(mai_mai_n497_));
  NO2        m475(.A(mai_mai_n81_), .B(i_9_), .Y(mai_mai_n498_));
  NA2        m476(.A(i_1_), .B(i_3_), .Y(mai_mai_n499_));
  NO2        m477(.A(mai_mai_n86_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NO2        m478(.A(mai_mai_n500_), .B(mai_mai_n497_), .Y(mai_mai_n501_));
  NA4        m479(.A(mai_mai_n501_), .B(mai_mai_n494_), .C(mai_mai_n489_), .D(mai_mai_n473_), .Y(mai_mai_n502_));
  NO3        m480(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n503_));
  OR2        m481(.A(mai_mai_n503_), .B(mai_mai_n204_), .Y(mai_mai_n504_));
  NA3        m482(.A(mai_mai_n360_), .B(mai_mai_n381_), .C(mai_mai_n45_), .Y(mai_mai_n505_));
  NA2        m483(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n506_));
  NA2        m484(.A(mai_mai_n506_), .B(mai_mai_n505_), .Y(mai_mai_n507_));
  OAI210     m485(.A0(mai_mai_n507_), .A1(mai_mai_n504_), .B0(i_1_), .Y(mai_mai_n508_));
  AOI210     m486(.A0(mai_mai_n213_), .A1(mai_mai_n90_), .B0(i_1_), .Y(mai_mai_n509_));
  NO2        m487(.A(mai_mai_n284_), .B(i_2_), .Y(mai_mai_n510_));
  NA2        m488(.A(mai_mai_n510_), .B(mai_mai_n509_), .Y(mai_mai_n511_));
  AOI210     m489(.A0(mai_mai_n511_), .A1(mai_mai_n508_), .B0(i_13_), .Y(mai_mai_n512_));
  NA2        m490(.A(i_12_), .B(mai_mai_n121_), .Y(mai_mai_n513_));
  AOI220     m491(.A0(mai_mai_n352_), .A1(mai_mai_n140_), .B0(i_2_), .B1(mai_mai_n121_), .Y(mai_mai_n514_));
  OAI210     m492(.A0(mai_mai_n514_), .A1(mai_mai_n43_), .B0(mai_mai_n513_), .Y(mai_mai_n515_));
  NO2        m493(.A(mai_mai_n53_), .B(mai_mai_n86_), .Y(mai_mai_n516_));
  AOI210     m494(.A0(mai_mai_n515_), .A1(mai_mai_n264_), .B0(mai_mai_n516_), .Y(mai_mai_n517_));
  AOI220     m495(.A0(i_12_), .A1(mai_mai_n69_), .B0(mai_mai_n299_), .B1(i_2_), .Y(mai_mai_n518_));
  NO2        m496(.A(mai_mai_n518_), .B(mai_mai_n202_), .Y(mai_mai_n519_));
  AOI210     m497(.A0(mai_mai_n339_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n520_));
  NOi31      m498(.An(mai_mai_n520_), .B(mai_mai_n439_), .C(mai_mai_n43_), .Y(mai_mai_n521_));
  NA2        m499(.A(mai_mai_n112_), .B(i_13_), .Y(mai_mai_n522_));
  NO2        m500(.A(mai_mai_n480_), .B(mai_mai_n99_), .Y(mai_mai_n523_));
  INV        m501(.A(mai_mai_n523_), .Y(mai_mai_n524_));
  OAI220     m502(.A0(mai_mai_n524_), .A1(mai_mai_n68_), .B0(mai_mai_n522_), .B1(mai_mai_n509_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n198_), .B(mai_mai_n81_), .Y(mai_mai_n526_));
  INV        m504(.A(mai_mai_n526_), .Y(mai_mai_n527_));
  AOI210     m505(.A0(mai_mai_n299_), .A1(i_2_), .B0(mai_mai_n85_), .Y(mai_mai_n528_));
  OAI220     m506(.A0(mai_mai_n528_), .A1(mai_mai_n442_), .B0(mai_mai_n527_), .B1(mai_mai_n452_), .Y(mai_mai_n529_));
  NO4        m507(.A(mai_mai_n529_), .B(mai_mai_n525_), .C(mai_mai_n521_), .D(mai_mai_n519_), .Y(mai_mai_n530_));
  NO2        m508(.A(mai_mai_n524_), .B(i_11_), .Y(mai_mai_n531_));
  NA2        m509(.A(i_2_), .B(mai_mai_n445_), .Y(mai_mai_n532_));
  NA2        m510(.A(mai_mai_n476_), .B(i_13_), .Y(mai_mai_n533_));
  NAi21      m511(.An(i_11_), .B(i_12_), .Y(mai_mai_n534_));
  NOi41      m512(.An(mai_mai_n96_), .B(mai_mai_n534_), .C(i_13_), .D(mai_mai_n81_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n427_), .B(mai_mai_n446_), .Y(mai_mai_n536_));
  AOI210     m514(.A0(mai_mai_n536_), .A1(mai_mai_n249_), .B0(mai_mai_n535_), .Y(mai_mai_n537_));
  NA3        m515(.A(mai_mai_n537_), .B(mai_mai_n533_), .C(mai_mai_n532_), .Y(mai_mai_n538_));
  OAI210     m516(.A0(mai_mai_n538_), .A1(mai_mai_n531_), .B0(mai_mai_n62_), .Y(mai_mai_n539_));
  NO3        m517(.A(i_9_), .B(i_3_), .C(mai_mai_n441_), .Y(mai_mai_n540_));
  NA2        m518(.A(mai_mai_n540_), .B(mai_mai_n283_), .Y(mai_mai_n541_));
  NO2        m519(.A(mai_mai_n113_), .B(i_2_), .Y(mai_mai_n542_));
  NA2        m520(.A(mai_mai_n542_), .B(mai_mai_n470_), .Y(mai_mai_n543_));
  NA2        m521(.A(mai_mai_n543_), .B(mai_mai_n541_), .Y(mai_mai_n544_));
  NA3        m522(.A(mai_mai_n544_), .B(mai_mai_n44_), .C(mai_mai_n189_), .Y(mai_mai_n545_));
  NA4        m523(.A(mai_mai_n545_), .B(mai_mai_n539_), .C(mai_mai_n530_), .D(mai_mai_n517_), .Y(mai_mai_n546_));
  OR4        m524(.A(mai_mai_n546_), .B(mai_mai_n512_), .C(mai_mai_n502_), .D(mai_mai_n455_), .Y(mai5));
  NA2        m525(.A(mai_mai_n491_), .B(mai_mai_n216_), .Y(mai_mai_n548_));
  NO2        m526(.A(mai_mai_n442_), .B(i_11_), .Y(mai_mai_n549_));
  INV        m527(.A(mai_mai_n549_), .Y(mai_mai_n550_));
  NA2        m528(.A(mai_mai_n550_), .B(mai_mai_n548_), .Y(mai_mai_n551_));
  NO3        m529(.A(i_11_), .B(mai_mai_n198_), .C(i_13_), .Y(mai_mai_n552_));
  NO2        m530(.A(mai_mai_n109_), .B(mai_mai_n23_), .Y(mai_mai_n553_));
  NA2        m531(.A(i_12_), .B(i_8_), .Y(mai_mai_n554_));
  NA2        m532(.A(i_12_), .B(mai_mai_n553_), .Y(mai_mai_n555_));
  INV        m533(.A(mai_mai_n555_), .Y(mai_mai_n556_));
  NO2        m534(.A(mai_mai_n556_), .B(mai_mai_n551_), .Y(mai_mai_n557_));
  INV        m535(.A(mai_mai_n146_), .Y(mai_mai_n558_));
  INV        m536(.A(mai_mai_n204_), .Y(mai_mai_n559_));
  OAI210     m537(.A0(mai_mai_n510_), .A1(mai_mai_n340_), .B0(mai_mai_n96_), .Y(mai_mai_n560_));
  AOI210     m538(.A0(mai_mai_n560_), .A1(mai_mai_n559_), .B0(mai_mai_n558_), .Y(mai_mai_n561_));
  INV        m539(.A(mai_mai_n317_), .Y(mai_mai_n562_));
  NA2        m540(.A(mai_mai_n562_), .B(i_2_), .Y(mai_mai_n563_));
  INV        m541(.A(mai_mai_n563_), .Y(mai_mai_n564_));
  AOI210     m542(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n314_), .Y(mai_mai_n565_));
  AOI210     m543(.A0(mai_mai_n565_), .A1(mai_mai_n564_), .B0(mai_mai_n561_), .Y(mai_mai_n566_));
  NO2        m544(.A(mai_mai_n161_), .B(mai_mai_n110_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n567_), .B(i_2_), .Y(mai_mai_n568_));
  NO2        m546(.A(mai_mai_n568_), .B(mai_mai_n164_), .Y(mai_mai_n569_));
  OA210      m547(.A0(mai_mai_n458_), .A1(mai_mai_n111_), .B0(i_13_), .Y(mai_mai_n570_));
  INV        m548(.A(mai_mai_n170_), .Y(mai_mai_n571_));
  INV        m549(.A(mai_mai_n133_), .Y(mai_mai_n572_));
  AOI210     m550(.A0(mai_mai_n572_), .A1(mai_mai_n571_), .B0(mai_mai_n287_), .Y(mai_mai_n573_));
  AOI210     m551(.A0(mai_mai_n177_), .A1(mai_mai_n130_), .B0(mai_mai_n381_), .Y(mai_mai_n574_));
  NA2        m552(.A(mai_mai_n574_), .B(mai_mai_n317_), .Y(mai_mai_n575_));
  NO2        m553(.A(i_2_), .B(mai_mai_n43_), .Y(mai_mai_n576_));
  NA2        m554(.A(mai_mai_n244_), .B(mai_mai_n41_), .Y(mai_mai_n577_));
  OAI210     m555(.A0(mai_mai_n577_), .A1(mai_mai_n576_), .B0(mai_mai_n575_), .Y(mai_mai_n578_));
  NO4        m556(.A(mai_mai_n578_), .B(mai_mai_n573_), .C(mai_mai_n570_), .D(mai_mai_n569_), .Y(mai_mai_n579_));
  INV        m557(.A(mai_mai_n422_), .Y(mai_mai_n580_));
  NA2        m558(.A(mai_mai_n552_), .B(mai_mai_n221_), .Y(mai_mai_n581_));
  NA2        m559(.A(mai_mai_n581_), .B(mai_mai_n580_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n583_));
  NO2        m561(.A(mai_mai_n583_), .B(mai_mai_n111_), .Y(mai_mai_n584_));
  NO2        m562(.A(mai_mai_n584_), .B(mai_mai_n440_), .Y(mai_mai_n585_));
  AOI220     m563(.A0(mai_mai_n585_), .A1(mai_mai_n36_), .B0(mai_mai_n582_), .B1(mai_mai_n45_), .Y(mai_mai_n586_));
  NA4        m564(.A(mai_mai_n586_), .B(mai_mai_n579_), .C(mai_mai_n566_), .D(mai_mai_n557_), .Y(mai6));
  NA2        m565(.A(mai_mai_n25_), .B(mai_mai_n542_), .Y(mai_mai_n588_));
  NA3        m566(.A(mai_mai_n302_), .B(i_8_), .C(mai_mai_n68_), .Y(mai_mai_n589_));
  INV        m567(.A(mai_mai_n589_), .Y(mai_mai_n590_));
  NO2        m568(.A(mai_mai_n187_), .B(i_2_), .Y(mai_mai_n591_));
  INV        m569(.A(i_9_), .Y(mai_mai_n592_));
  NO2        m570(.A(mai_mai_n590_), .B(mai_mai_n261_), .Y(mai_mai_n593_));
  AO210      m571(.A0(mai_mai_n593_), .A1(mai_mai_n588_), .B0(i_12_), .Y(mai_mai_n594_));
  NA2        m572(.A(mai_mai_n288_), .B(mai_mai_n265_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n427_), .B(mai_mai_n62_), .Y(mai_mai_n596_));
  NA2        m574(.A(mai_mai_n596_), .B(mai_mai_n595_), .Y(mai_mai_n597_));
  INV        m575(.A(mai_mai_n167_), .Y(mai_mai_n598_));
  AOI220     m576(.A0(mai_mai_n598_), .A1(mai_mai_n592_), .B0(mai_mai_n597_), .B1(mai_mai_n70_), .Y(mai_mai_n599_));
  NA2        m577(.A(mai_mai_n767_), .B(mai_mai_n583_), .Y(mai_mai_n600_));
  AOI210     m578(.A0(mai_mai_n600_), .A1(mai_mai_n379_), .B0(mai_mai_n156_), .Y(mai_mai_n601_));
  NA3        m579(.A(mai_mai_n770_), .B(mai_mai_n354_), .C(mai_mai_n302_), .Y(mai_mai_n602_));
  NA2        m580(.A(mai_mai_n414_), .B(mai_mai_n413_), .Y(mai_mai_n603_));
  NA2        m581(.A(mai_mai_n603_), .B(mai_mai_n602_), .Y(mai_mai_n604_));
  OR2        m582(.A(mai_mai_n604_), .B(mai_mai_n601_), .Y(mai_mai_n605_));
  NO2        m583(.A(i_11_), .B(i_2_), .Y(mai_mai_n606_));
  NA2        m584(.A(mai_mai_n47_), .B(mai_mai_n37_), .Y(mai_mai_n607_));
  NO2        m585(.A(mai_mai_n607_), .B(mai_mai_n313_), .Y(mai_mai_n608_));
  NA2        m586(.A(mai_mai_n608_), .B(mai_mai_n606_), .Y(mai_mai_n609_));
  NA3        m587(.A(mai_mai_n772_), .B(mai_mai_n209_), .C(i_7_), .Y(mai_mai_n610_));
  BUFFER     m588(.A(mai_mai_n340_), .Y(mai_mai_n611_));
  NA2        m589(.A(mai_mai_n611_), .B(mai_mai_n129_), .Y(mai_mai_n612_));
  NA3        m590(.A(mai_mai_n612_), .B(mai_mai_n610_), .C(mai_mai_n609_), .Y(mai_mai_n613_));
  AOI210     m591(.A0(mai_mai_n765_), .A1(mai_mai_n413_), .B0(mai_mai_n591_), .Y(mai_mai_n614_));
  NA2        m592(.A(mai_mai_n199_), .B(mai_mai_n129_), .Y(mai_mai_n615_));
  OAI210     m593(.A0(mai_mai_n305_), .A1(mai_mai_n172_), .B0(mai_mai_n67_), .Y(mai_mai_n616_));
  NA4        m594(.A(mai_mai_n616_), .B(mai_mai_n615_), .C(mai_mai_n614_), .D(mai_mai_n444_), .Y(mai_mai_n617_));
  NA3        m595(.A(mai_mai_n381_), .B(mai_mai_n360_), .C(mai_mai_n185_), .Y(mai_mai_n618_));
  AOI210     m596(.A0(mai_mai_n340_), .A1(mai_mai_n338_), .B0(mai_mai_n412_), .Y(mai_mai_n619_));
  INV        m597(.A(mai_mai_n312_), .Y(mai_mai_n620_));
  INV        m598(.A(mai_mai_n432_), .Y(mai_mai_n621_));
  NA3        m599(.A(mai_mai_n621_), .B(mai_mai_n260_), .C(i_7_), .Y(mai_mai_n622_));
  NA4        m600(.A(mai_mai_n622_), .B(mai_mai_n620_), .C(mai_mai_n619_), .D(mai_mai_n618_), .Y(mai_mai_n623_));
  NO4        m601(.A(mai_mai_n623_), .B(mai_mai_n617_), .C(mai_mai_n613_), .D(mai_mai_n605_), .Y(mai_mai_n624_));
  NA4        m602(.A(mai_mai_n624_), .B(mai_mai_n599_), .C(mai_mai_n594_), .D(mai_mai_n295_), .Y(mai3));
  NA2        m603(.A(i_12_), .B(i_10_), .Y(mai_mai_n626_));
  NO2        m604(.A(i_11_), .B(mai_mai_n198_), .Y(mai_mai_n627_));
  NA2        m605(.A(mai_mai_n233_), .B(mai_mai_n627_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n628_), .B(mai_mai_n164_), .Y(mai_mai_n629_));
  NO2        m607(.A(mai_mai_n83_), .B(mai_mai_n43_), .Y(mai_mai_n630_));
  OA210      m608(.A0(mai_mai_n630_), .A1(mai_mai_n629_), .B0(mai_mai_n148_), .Y(mai_mai_n631_));
  NO3        m609(.A(mai_mai_n466_), .B(mai_mai_n343_), .C(mai_mai_n116_), .Y(mai_mai_n632_));
  NA2        m610(.A(i_2_), .B(mai_mai_n44_), .Y(mai_mai_n633_));
  AN2        m611(.A(mai_mai_n342_), .B(mai_mai_n54_), .Y(mai_mai_n634_));
  NO2        m612(.A(mai_mai_n634_), .B(mai_mai_n632_), .Y(mai_mai_n635_));
  INV        m613(.A(mai_mai_n635_), .Y(mai_mai_n636_));
  NO3        m614(.A(mai_mai_n291_), .B(mai_mai_n38_), .C(i_0_), .Y(mai_mai_n637_));
  NO2        m615(.A(mai_mai_n779_), .B(mai_mai_n62_), .Y(mai_mai_n638_));
  NOi21      m616(.An(i_5_), .B(i_9_), .Y(mai_mai_n639_));
  NA2        m617(.A(mai_mai_n639_), .B(mai_mai_n337_), .Y(mai_mai_n640_));
  NO2        m618(.A(mai_mai_n149_), .B(mai_mai_n130_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n641_), .B(mai_mai_n203_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n642_), .B(mai_mai_n152_), .Y(mai_mai_n643_));
  NO4        m621(.A(mai_mai_n643_), .B(mai_mai_n638_), .C(mai_mai_n636_), .D(mai_mai_n631_), .Y(mai_mai_n644_));
  NA2        m622(.A(mai_mai_n156_), .B(mai_mai_n24_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n102_), .B(mai_mai_n645_), .Y(mai_mai_n646_));
  NA2        m624(.A(mai_mai_n249_), .B(mai_mai_n114_), .Y(mai_mai_n647_));
  NO2        m625(.A(mai_mai_n647_), .B(mai_mai_n307_), .Y(mai_mai_n648_));
  NO2        m626(.A(mai_mai_n648_), .B(mai_mai_n646_), .Y(mai_mai_n649_));
  NA2        m627(.A(i_6_), .B(i_0_), .Y(mai_mai_n650_));
  NO4        m628(.A(i_5_), .B(mai_mai_n182_), .C(mai_mai_n314_), .D(mai_mai_n313_), .Y(mai_mai_n651_));
  NA2        m629(.A(mai_mai_n651_), .B(i_11_), .Y(mai_mai_n652_));
  NA2        m630(.A(mai_mai_n552_), .B(mai_mai_n261_), .Y(mai_mai_n653_));
  OAI220     m631(.A0(i_6_), .A1(mai_mai_n653_), .B0(mai_mai_n486_), .B1(mai_mai_n393_), .Y(mai_mai_n654_));
  NO2        m632(.A(mai_mai_n207_), .B(mai_mai_n134_), .Y(mai_mai_n655_));
  NA2        m633(.A(i_0_), .B(i_10_), .Y(mai_mai_n656_));
  NO4        m634(.A(mai_mai_n99_), .B(mai_mai_n57_), .C(mai_mai_n495_), .D(i_5_), .Y(mai_mai_n657_));
  AO220      m635(.A0(mai_mai_n657_), .A1(i_0_), .B0(mai_mai_n655_), .B1(i_6_), .Y(mai_mai_n658_));
  NO2        m636(.A(mai_mai_n658_), .B(mai_mai_n654_), .Y(mai_mai_n659_));
  NA3        m637(.A(mai_mai_n659_), .B(mai_mai_n652_), .C(mai_mai_n649_), .Y(mai_mai_n660_));
  NA2        m638(.A(i_11_), .B(i_9_), .Y(mai_mai_n661_));
  NA2        m639(.A(mai_mai_n304_), .B(mai_mai_n151_), .Y(mai_mai_n662_));
  NA2        m640(.A(mai_mai_n662_), .B(mai_mai_n139_), .Y(mai_mai_n663_));
  NO2        m641(.A(mai_mai_n661_), .B(mai_mai_n70_), .Y(mai_mai_n664_));
  NO2        m642(.A(mai_mai_n149_), .B(i_0_), .Y(mai_mai_n665_));
  NA2        m643(.A(mai_mai_n354_), .B(mai_mai_n194_), .Y(mai_mai_n666_));
  OAI220     m644(.A0(i_12_), .A1(mai_mai_n640_), .B0(mai_mai_n666_), .B1(mai_mai_n149_), .Y(mai_mai_n667_));
  NO2        m645(.A(mai_mai_n667_), .B(mai_mai_n663_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n485_), .B(mai_mai_n106_), .Y(mai_mai_n669_));
  NO2        m647(.A(i_6_), .B(mai_mai_n669_), .Y(mai_mai_n670_));
  AOI210     m648(.A0(mai_mai_n339_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n146_), .B(mai_mai_n92_), .Y(mai_mai_n672_));
  NOi32      m650(.An(mai_mai_n671_), .Bn(mai_mai_n159_), .C(mai_mai_n672_), .Y(mai_mai_n673_));
  NO2        m651(.A(mai_mai_n37_), .B(mai_mai_n633_), .Y(mai_mai_n674_));
  NO3        m652(.A(mai_mai_n674_), .B(mai_mai_n673_), .C(mai_mai_n670_), .Y(mai_mai_n675_));
  NOi31      m653(.An(i_7_), .B(i_0_), .C(mai_mai_n534_), .Y(mai_mai_n676_));
  NA2        m654(.A(mai_mai_n675_), .B(mai_mai_n668_), .Y(mai_mai_n677_));
  INV        m655(.A(mai_mai_n626_), .Y(mai_mai_n678_));
  OA210      m656(.A0(mai_mai_n354_), .A1(mai_mai_n188_), .B0(mai_mai_n353_), .Y(mai_mai_n679_));
  NA2        m657(.A(mai_mai_n678_), .B(mai_mai_n664_), .Y(mai_mai_n680_));
  NA3        m658(.A(mai_mai_n353_), .B(i_2_), .C(mai_mai_n44_), .Y(mai_mai_n681_));
  INV        m659(.A(mai_mai_n681_), .Y(mai_mai_n682_));
  INV        m660(.A(mai_mai_n158_), .Y(mai_mai_n683_));
  AOI220     m661(.A0(mai_mai_n683_), .A1(mai_mai_n354_), .B0(mai_mai_n682_), .B1(mai_mai_n70_), .Y(mai_mai_n684_));
  NA2        m662(.A(mai_mai_n86_), .B(mai_mai_n43_), .Y(mai_mai_n685_));
  NO2        m663(.A(mai_mai_n72_), .B(mai_mai_n554_), .Y(mai_mai_n686_));
  NA2        m664(.A(mai_mai_n686_), .B(mai_mai_n685_), .Y(mai_mai_n687_));
  NO2        m665(.A(mai_mai_n687_), .B(mai_mai_n46_), .Y(mai_mai_n688_));
  NO3        m666(.A(i_5_), .B(i_0_), .C(mai_mai_n24_), .Y(mai_mai_n689_));
  INV        m667(.A(mai_mai_n689_), .Y(mai_mai_n690_));
  NO2        m668(.A(mai_mai_n690_), .B(mai_mai_n147_), .Y(mai_mai_n691_));
  NO3        m669(.A(mai_mai_n691_), .B(mai_mai_n688_), .C(mai_mai_n383_), .Y(mai_mai_n692_));
  NA3        m670(.A(mai_mai_n692_), .B(mai_mai_n684_), .C(mai_mai_n680_), .Y(mai_mai_n693_));
  NO3        m671(.A(mai_mai_n693_), .B(mai_mai_n677_), .C(mai_mai_n660_), .Y(mai_mai_n694_));
  NO2        m672(.A(i_0_), .B(mai_mai_n534_), .Y(mai_mai_n695_));
  NO2        m673(.A(mai_mai_n596_), .B(mai_mai_n672_), .Y(mai_mai_n696_));
  INV        m674(.A(mai_mai_n696_), .Y(mai_mai_n697_));
  NA3        m675(.A(mai_mai_n128_), .B(mai_mai_n498_), .C(mai_mai_n70_), .Y(mai_mai_n698_));
  NA2        m676(.A(mai_mai_n627_), .B(i_9_), .Y(mai_mai_n699_));
  AOI210     m677(.A0(mai_mai_n775_), .A1(mai_mai_n365_), .B0(mai_mai_n699_), .Y(mai_mai_n700_));
  NA2        m678(.A(mai_mai_n203_), .B(i_10_), .Y(mai_mai_n701_));
  AOI210     m679(.A0(mai_mai_n701_), .A1(mai_mai_n650_), .B0(mai_mai_n134_), .Y(mai_mai_n702_));
  NO2        m680(.A(mai_mai_n702_), .B(mai_mai_n700_), .Y(mai_mai_n703_));
  NA3        m681(.A(mai_mai_n703_), .B(mai_mai_n698_), .C(mai_mai_n697_), .Y(mai_mai_n704_));
  NO2        m682(.A(mai_mai_n141_), .B(mai_mai_n768_), .Y(mai_mai_n705_));
  INV        m683(.A(mai_mai_n705_), .Y(mai_mai_n706_));
  NA2        m684(.A(mai_mai_n418_), .B(mai_mai_n72_), .Y(mai_mai_n707_));
  NO3        m685(.A(mai_mai_n178_), .B(mai_mai_n297_), .C(i_0_), .Y(mai_mai_n708_));
  OAI210     m686(.A0(mai_mai_n708_), .A1(mai_mai_n73_), .B0(i_13_), .Y(mai_mai_n709_));
  NA3        m687(.A(mai_mai_n709_), .B(mai_mai_n707_), .C(mai_mai_n706_), .Y(mai_mai_n710_));
  AOI210     m688(.A0(i_6_), .A1(mai_mai_n695_), .B0(mai_mai_n94_), .Y(mai_mai_n711_));
  BUFFER     m689(.A(mai_mai_n711_), .Y(mai_mai_n712_));
  AOI210     m690(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n149_), .Y(mai_mai_n713_));
  NA2        m691(.A(mai_mai_n713_), .B(mai_mai_n679_), .Y(mai_mai_n714_));
  NOi31      m692(.An(mai_mai_n301_), .B(i_11_), .C(mai_mai_n200_), .Y(mai_mai_n715_));
  NO3        m693(.A(mai_mai_n661_), .B(mai_mai_n185_), .C(mai_mai_n161_), .Y(mai_mai_n716_));
  NO2        m694(.A(mai_mai_n716_), .B(mai_mai_n715_), .Y(mai_mai_n717_));
  NA3        m695(.A(mai_mai_n717_), .B(mai_mai_n714_), .C(mai_mai_n712_), .Y(mai_mai_n718_));
  NAi21      m696(.An(mai_mai_n201_), .B(mai_mai_n202_), .Y(mai_mai_n719_));
  NO4        m697(.A(mai_mai_n200_), .B(mai_mai_n178_), .C(i_0_), .D(i_12_), .Y(mai_mai_n720_));
  AOI220     m698(.A0(mai_mai_n720_), .A1(mai_mai_n719_), .B0(mai_mai_n590_), .B1(mai_mai_n150_), .Y(mai_mai_n721_));
  AN2        m699(.A(mai_mai_n656_), .B(mai_mai_n134_), .Y(mai_mai_n722_));
  NO4        m700(.A(mai_mai_n722_), .B(i_12_), .C(mai_mai_n478_), .D(mai_mai_n116_), .Y(mai_mai_n723_));
  INV        m701(.A(mai_mai_n723_), .Y(mai_mai_n724_));
  NA2        m702(.A(mai_mai_n421_), .B(i_11_), .Y(mai_mai_n725_));
  NO2        m703(.A(mai_mai_n725_), .B(mai_mai_n778_), .Y(mai_mai_n726_));
  NA2        m704(.A(i_7_), .B(mai_mai_n352_), .Y(mai_mai_n727_));
  OAI220     m705(.A0(i_6_), .A1(mai_mai_n776_), .B0(mai_mai_n727_), .B1(i_1_), .Y(mai_mai_n728_));
  AOI210     m706(.A0(mai_mai_n728_), .A1(mai_mai_n665_), .B0(mai_mai_n726_), .Y(mai_mai_n729_));
  NA3        m707(.A(mai_mai_n729_), .B(mai_mai_n724_), .C(mai_mai_n721_), .Y(mai_mai_n730_));
  NO4        m708(.A(mai_mai_n730_), .B(mai_mai_n718_), .C(mai_mai_n710_), .D(mai_mai_n704_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n770_), .B(mai_mai_n37_), .Y(mai_mai_n732_));
  NA2        m710(.A(mai_mai_n732_), .B(mai_mai_n764_), .Y(mai_mai_n733_));
  NA2        m711(.A(mai_mai_n733_), .B(mai_mai_n175_), .Y(mai_mai_n734_));
  OAI210     m712(.A0(mai_mai_n451_), .A1(mai_mai_n449_), .B0(mai_mai_n251_), .Y(mai_mai_n735_));
  INV        m713(.A(mai_mai_n735_), .Y(mai_mai_n736_));
  NO4        m714(.A(mai_mai_n196_), .B(mai_mai_n127_), .C(mai_mai_n499_), .D(mai_mai_n37_), .Y(mai_mai_n737_));
  NO2        m715(.A(mai_mai_n737_), .B(mai_mai_n651_), .Y(mai_mai_n738_));
  NA2        m716(.A(mai_mai_n725_), .B(mai_mai_n738_), .Y(mai_mai_n739_));
  AOI210     m717(.A0(mai_mai_n736_), .A1(mai_mai_n47_), .B0(mai_mai_n739_), .Y(mai_mai_n740_));
  AOI210     m718(.A0(mai_mai_n740_), .A1(mai_mai_n734_), .B0(mai_mai_n70_), .Y(mai_mai_n741_));
  NO2        m719(.A(mai_mai_n415_), .B(mai_mai_n294_), .Y(mai_mai_n742_));
  NO2        m720(.A(mai_mai_n742_), .B(mai_mai_n558_), .Y(mai_mai_n743_));
  INV        m721(.A(mai_mai_n93_), .Y(mai_mai_n744_));
  NA2        m722(.A(mai_mai_n744_), .B(mai_mai_n73_), .Y(mai_mai_n745_));
  AOI210     m723(.A0(mai_mai_n713_), .A1(mai_mai_n777_), .B0(mai_mai_n676_), .Y(mai_mai_n746_));
  AOI210     m724(.A0(mai_mai_n746_), .A1(mai_mai_n745_), .B0(mai_mai_n499_), .Y(mai_mai_n747_));
  INV        m725(.A(mai_mai_n56_), .Y(mai_mai_n748_));
  NA2        m726(.A(mai_mai_n748_), .B(mai_mai_n73_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n749_), .B(mai_mai_n198_), .Y(mai_mai_n750_));
  NO2        m728(.A(mai_mai_n750_), .B(mai_mai_n747_), .Y(mai_mai_n751_));
  NO3        m729(.A(mai_mai_n58_), .B(mai_mai_n57_), .C(i_4_), .Y(mai_mai_n752_));
  INV        m730(.A(mai_mai_n752_), .Y(mai_mai_n753_));
  NO2        m731(.A(mai_mai_n753_), .B(mai_mai_n534_), .Y(mai_mai_n754_));
  INV        m732(.A(mai_mai_n412_), .Y(mai_mai_n755_));
  NO2        m733(.A(mai_mai_n755_), .B(mai_mai_n40_), .Y(mai_mai_n756_));
  NO3        m734(.A(mai_mai_n756_), .B(mai_mai_n754_), .C(mai_mai_n215_), .Y(mai_mai_n757_));
  OAI210     m735(.A0(mai_mai_n751_), .A1(i_4_), .B0(mai_mai_n757_), .Y(mai_mai_n758_));
  NO3        m736(.A(mai_mai_n758_), .B(mai_mai_n743_), .C(mai_mai_n741_), .Y(mai_mai_n759_));
  NA4        m737(.A(mai_mai_n759_), .B(mai_mai_n731_), .C(mai_mai_n694_), .D(mai_mai_n644_), .Y(mai4));
  INV        m738(.A(i_2_), .Y(mai_mai_n763_));
  INV        m739(.A(mai_mai_n140_), .Y(mai_mai_n764_));
  INV        m740(.A(i_11_), .Y(mai_mai_n765_));
  INV        m741(.A(mai_mai_n116_), .Y(mai_mai_n766_));
  INV        m742(.A(i_9_), .Y(mai_mai_n767_));
  INV        m743(.A(mai_mai_n261_), .Y(mai_mai_n768_));
  INV        m744(.A(i_1_), .Y(mai_mai_n769_));
  INV        m745(.A(i_11_), .Y(mai_mai_n770_));
  INV        m746(.A(i_7_), .Y(mai_mai_n771_));
  INV        m747(.A(i_9_), .Y(mai_mai_n772_));
  INV        m748(.A(i_6_), .Y(mai_mai_n773_));
  INV        m749(.A(i_10_), .Y(mai_mai_n774_));
  INV        m750(.A(i_6_), .Y(mai_mai_n775_));
  INV        m751(.A(i_10_), .Y(mai_mai_n776_));
  INV        m752(.A(i_7_), .Y(mai_mai_n777_));
  INV        m753(.A(i_2_), .Y(mai_mai_n778_));
  INV        m754(.A(mai_mai_n637_), .Y(mai_mai_n779_));
  INV        m755(.A(i_0_), .Y(mai_mai_n780_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  OAI210     u0006(.A0(men_men_n27_), .A1(men_men_n24_), .B0(i_10_), .Y(men_men_n29_));
  NOi21      u0007(.An(i_11_), .B(i_8_), .Y(men_men_n30_));
  AO210      u0008(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n31_));
  OR2        u0009(.A(men_men_n31_), .B(men_men_n30_), .Y(men_men_n32_));
  NA2        u0010(.A(men_men_n32_), .B(men_men_n29_), .Y(men_men_n33_));
  XO2        u0011(.A(men_men_n33_), .B(men_men_n23_), .Y(men_men_n34_));
  INV        u0012(.A(i_4_), .Y(men_men_n35_));
  INV        u0013(.A(i_10_), .Y(men_men_n36_));
  NAi21      u0014(.An(i_11_), .B(i_9_), .Y(men_men_n37_));
  NO3        u0015(.A(men_men_n37_), .B(i_12_), .C(men_men_n36_), .Y(men_men_n38_));
  NOi21      u0016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u0017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u0018(.A(men_men_n35_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n34_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NA2        u0026(.A(i_7_), .B(men_men_n25_), .Y(men_men_n49_));
  NO2        u0027(.A(men_men_n47_), .B(men_men_n46_), .Y(men_men_n50_));
  NA2        u0028(.A(i_0_), .B(i_2_), .Y(men_men_n51_));
  NA2        u0029(.A(i_7_), .B(i_9_), .Y(men_men_n52_));
  NO2        u0030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NA2        u0031(.A(men_men_n50_), .B(men_men_n45_), .Y(men_men_n54_));
  NA3        u0032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n55_));
  NO2        u0033(.A(i_1_), .B(i_6_), .Y(men_men_n56_));
  NA2        u0034(.A(i_8_), .B(i_7_), .Y(men_men_n57_));
  OAI210     u0035(.A0(men_men_n57_), .A1(men_men_n56_), .B0(men_men_n55_), .Y(men_men_n58_));
  NA2        u0036(.A(men_men_n58_), .B(i_12_), .Y(men_men_n59_));
  NAi21      u0037(.An(i_2_), .B(i_7_), .Y(men_men_n60_));
  INV        u0038(.A(i_1_), .Y(men_men_n61_));
  NA2        u0039(.A(men_men_n61_), .B(i_6_), .Y(men_men_n62_));
  NA2        u0040(.A(i_1_), .B(i_10_), .Y(men_men_n63_));
  NO2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NAi21      u0042(.An(men_men_n64_), .B(men_men_n59_), .Y(men_men_n65_));
  NA2        u0043(.A(men_men_n49_), .B(i_2_), .Y(men_men_n66_));
  NA2        u0044(.A(i_1_), .B(i_6_), .Y(men_men_n67_));
  NO2        u0045(.A(men_men_n67_), .B(men_men_n25_), .Y(men_men_n68_));
  INV        u0046(.A(i_0_), .Y(men_men_n69_));
  NAi21      u0047(.An(i_5_), .B(i_10_), .Y(men_men_n70_));
  NA2        u0048(.A(i_5_), .B(i_9_), .Y(men_men_n71_));
  AOI210     u0049(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n69_), .Y(men_men_n72_));
  NO2        u0050(.A(men_men_n72_), .B(men_men_n68_), .Y(men_men_n73_));
  OAI210     u0051(.A0(men_men_n72_), .A1(men_men_n65_), .B0(i_0_), .Y(men_men_n74_));
  NA2        u0052(.A(i_12_), .B(i_5_), .Y(men_men_n75_));
  NA2        u0053(.A(i_2_), .B(i_8_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n56_), .Y(men_men_n77_));
  NO2        u0055(.A(i_3_), .B(i_9_), .Y(men_men_n78_));
  NO2        u0056(.A(i_3_), .B(i_7_), .Y(men_men_n79_));
  NO3        u0057(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n61_), .Y(men_men_n80_));
  INV        u0058(.A(i_6_), .Y(men_men_n81_));
  OR4        u0059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n82_));
  INV        u0060(.A(men_men_n82_), .Y(men_men_n83_));
  NO2        u0061(.A(i_2_), .B(i_7_), .Y(men_men_n84_));
  OAI210     u0062(.A0(men_men_n80_), .A1(men_men_n77_), .B0(i_2_), .Y(men_men_n85_));
  NAi21      u0063(.An(i_6_), .B(i_10_), .Y(men_men_n86_));
  NA2        u0064(.A(i_6_), .B(i_9_), .Y(men_men_n87_));
  NA2        u0065(.A(i_2_), .B(i_6_), .Y(men_men_n88_));
  AOI210     u0066(.A0(men_men_n87_), .A1(men_men_n85_), .B0(men_men_n75_), .Y(men_men_n89_));
  AN3        u0067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n90_));
  NAi21      u0068(.An(i_6_), .B(i_11_), .Y(men_men_n91_));
  NO2        u0069(.A(i_5_), .B(i_8_), .Y(men_men_n92_));
  NOi21      u0070(.An(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  AOI220     u0071(.A0(men_men_n93_), .A1(men_men_n60_), .B0(men_men_n90_), .B1(men_men_n31_), .Y(men_men_n94_));
  INV        u0072(.A(i_7_), .Y(men_men_n95_));
  NA2        u0073(.A(men_men_n46_), .B(men_men_n95_), .Y(men_men_n96_));
  NO2        u0074(.A(i_0_), .B(i_5_), .Y(men_men_n97_));
  NO2        u0075(.A(men_men_n97_), .B(men_men_n81_), .Y(men_men_n98_));
  NA2        u0076(.A(i_12_), .B(i_3_), .Y(men_men_n99_));
  INV        u0077(.A(men_men_n99_), .Y(men_men_n100_));
  NA3        u0078(.A(men_men_n100_), .B(men_men_n98_), .C(men_men_n96_), .Y(men_men_n101_));
  NAi21      u0079(.An(i_7_), .B(i_11_), .Y(men_men_n102_));
  NO3        u0080(.A(men_men_n102_), .B(men_men_n86_), .C(men_men_n51_), .Y(men_men_n103_));
  AN2        u0081(.A(i_2_), .B(i_10_), .Y(men_men_n104_));
  NO2        u0082(.A(men_men_n104_), .B(i_7_), .Y(men_men_n105_));
  OR2        u0083(.A(men_men_n75_), .B(men_men_n56_), .Y(men_men_n106_));
  NO2        u0084(.A(i_8_), .B(men_men_n95_), .Y(men_men_n107_));
  NO3        u0085(.A(men_men_n107_), .B(men_men_n106_), .C(men_men_n105_), .Y(men_men_n108_));
  NA2        u0086(.A(i_12_), .B(i_7_), .Y(men_men_n109_));
  NO2        u0087(.A(men_men_n61_), .B(men_men_n26_), .Y(men_men_n110_));
  INV        u0088(.A(men_men_n110_), .Y(men_men_n111_));
  NA2        u0089(.A(i_11_), .B(i_12_), .Y(men_men_n112_));
  OAI210     u0090(.A0(men_men_n111_), .A1(men_men_n109_), .B0(men_men_n112_), .Y(men_men_n113_));
  NO2        u0091(.A(men_men_n113_), .B(men_men_n108_), .Y(men_men_n114_));
  NAi41      u0092(.An(men_men_n103_), .B(men_men_n114_), .C(men_men_n101_), .D(men_men_n94_), .Y(men_men_n115_));
  NOi21      u0093(.An(i_1_), .B(i_5_), .Y(men_men_n116_));
  NA2        u0094(.A(men_men_n116_), .B(i_11_), .Y(men_men_n117_));
  NA2        u0095(.A(men_men_n95_), .B(men_men_n36_), .Y(men_men_n118_));
  NA2        u0096(.A(i_7_), .B(men_men_n25_), .Y(men_men_n119_));
  NA2        u0097(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NO2        u0098(.A(men_men_n120_), .B(men_men_n46_), .Y(men_men_n121_));
  NAi21      u0099(.An(i_3_), .B(i_8_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n122_), .B(men_men_n60_), .Y(men_men_n123_));
  INV        u0101(.A(men_men_n121_), .Y(men_men_n124_));
  NO2        u0102(.A(i_1_), .B(men_men_n81_), .Y(men_men_n125_));
  NO2        u0103(.A(i_6_), .B(i_5_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n126_), .B(i_3_), .Y(men_men_n127_));
  AO210      u0105(.A0(men_men_n127_), .A1(men_men_n47_), .B0(men_men_n125_), .Y(men_men_n128_));
  OAI220     u0106(.A0(men_men_n128_), .A1(men_men_n102_), .B0(men_men_n124_), .B1(men_men_n117_), .Y(men_men_n129_));
  NO3        u0107(.A(men_men_n129_), .B(men_men_n115_), .C(men_men_n89_), .Y(men_men_n130_));
  NA3        u0108(.A(men_men_n130_), .B(men_men_n74_), .C(men_men_n54_), .Y(men2));
  NO2        u0109(.A(men_men_n61_), .B(men_men_n36_), .Y(men_men_n132_));
  NA3        u0110(.A(men_men_n73_), .B(men_men_n66_), .C(men_men_n29_), .Y(men0));
  AN2        u0111(.A(i_8_), .B(i_7_), .Y(men_men_n134_));
  NA2        u0112(.A(men_men_n134_), .B(i_6_), .Y(men_men_n135_));
  NO2        u0113(.A(i_12_), .B(i_13_), .Y(men_men_n136_));
  NAi21      u0114(.An(i_5_), .B(i_11_), .Y(men_men_n137_));
  NOi21      u0115(.An(men_men_n136_), .B(men_men_n137_), .Y(men_men_n138_));
  NO2        u0116(.A(i_0_), .B(i_1_), .Y(men_men_n139_));
  NA2        u0117(.A(i_2_), .B(i_3_), .Y(men_men_n140_));
  NO2        u0118(.A(men_men_n140_), .B(i_4_), .Y(men_men_n141_));
  NA3        u0119(.A(men_men_n141_), .B(men_men_n139_), .C(men_men_n138_), .Y(men_men_n142_));
  OR2        u0120(.A(men_men_n142_), .B(men_men_n25_), .Y(men_men_n143_));
  AN2        u0121(.A(men_men_n136_), .B(men_men_n78_), .Y(men_men_n144_));
  NO2        u0122(.A(men_men_n144_), .B(men_men_n27_), .Y(men_men_n145_));
  NA2        u0123(.A(i_1_), .B(i_5_), .Y(men_men_n146_));
  NO2        u0124(.A(men_men_n69_), .B(men_men_n46_), .Y(men_men_n147_));
  NA2        u0125(.A(men_men_n147_), .B(men_men_n35_), .Y(men_men_n148_));
  NO3        u0126(.A(men_men_n148_), .B(men_men_n146_), .C(men_men_n145_), .Y(men_men_n149_));
  OR2        u0127(.A(i_0_), .B(i_1_), .Y(men_men_n150_));
  NO3        u0128(.A(men_men_n150_), .B(men_men_n75_), .C(i_13_), .Y(men_men_n151_));
  NAi32      u0129(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n152_));
  NAi21      u0130(.An(men_men_n152_), .B(men_men_n151_), .Y(men_men_n153_));
  NOi21      u0131(.An(i_4_), .B(i_10_), .Y(men_men_n154_));
  NA2        u0132(.A(men_men_n154_), .B(men_men_n39_), .Y(men_men_n155_));
  NO2        u0133(.A(i_3_), .B(i_5_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n69_), .B(i_2_), .C(i_1_), .Y(men_men_n157_));
  NA2        u0135(.A(men_men_n157_), .B(men_men_n156_), .Y(men_men_n158_));
  OAI210     u0136(.A0(men_men_n158_), .A1(men_men_n155_), .B0(men_men_n153_), .Y(men_men_n159_));
  NO2        u0137(.A(men_men_n159_), .B(men_men_n149_), .Y(men_men_n160_));
  AOI210     u0138(.A0(men_men_n160_), .A1(men_men_n143_), .B0(men_men_n135_), .Y(men_men_n161_));
  NA3        u0139(.A(men_men_n69_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n162_));
  NA2        u0140(.A(i_3_), .B(men_men_n48_), .Y(men_men_n163_));
  NOi21      u0141(.An(i_4_), .B(i_9_), .Y(men_men_n164_));
  NOi21      u0142(.An(i_11_), .B(i_13_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  OR2        u0144(.A(men_men_n166_), .B(men_men_n163_), .Y(men_men_n167_));
  NO2        u0145(.A(i_4_), .B(i_5_), .Y(men_men_n168_));
  NAi21      u0146(.An(i_12_), .B(i_11_), .Y(men_men_n169_));
  NO2        u0147(.A(men_men_n169_), .B(i_13_), .Y(men_men_n170_));
  NA3        u0148(.A(men_men_n170_), .B(men_men_n168_), .C(men_men_n78_), .Y(men_men_n171_));
  AOI210     u0149(.A0(men_men_n171_), .A1(men_men_n167_), .B0(men_men_n162_), .Y(men_men_n172_));
  NO2        u0150(.A(men_men_n69_), .B(men_men_n61_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n46_), .Y(men_men_n174_));
  NA2        u0152(.A(men_men_n35_), .B(i_5_), .Y(men_men_n175_));
  NAi31      u0153(.An(men_men_n175_), .B(men_men_n144_), .C(i_11_), .Y(men_men_n176_));
  NA2        u0154(.A(i_3_), .B(i_5_), .Y(men_men_n177_));
  OR2        u0155(.A(men_men_n177_), .B(men_men_n166_), .Y(men_men_n178_));
  AOI210     u0156(.A0(men_men_n178_), .A1(men_men_n176_), .B0(men_men_n174_), .Y(men_men_n179_));
  NO2        u0157(.A(men_men_n69_), .B(i_5_), .Y(men_men_n180_));
  NO2        u0158(.A(i_13_), .B(i_10_), .Y(men_men_n181_));
  NA3        u0159(.A(men_men_n181_), .B(men_men_n180_), .C(men_men_n44_), .Y(men_men_n182_));
  NO2        u0160(.A(i_2_), .B(i_1_), .Y(men_men_n183_));
  NA2        u0161(.A(men_men_n183_), .B(i_3_), .Y(men_men_n184_));
  NAi21      u0162(.An(i_4_), .B(i_12_), .Y(men_men_n185_));
  NO3        u0163(.A(men_men_n185_), .B(men_men_n184_), .C(men_men_n182_), .Y(men_men_n186_));
  NO3        u0164(.A(men_men_n186_), .B(men_men_n179_), .C(men_men_n172_), .Y(men_men_n187_));
  INV        u0165(.A(i_8_), .Y(men_men_n188_));
  NO2        u0166(.A(men_men_n188_), .B(i_7_), .Y(men_men_n189_));
  NA2        u0167(.A(men_men_n189_), .B(i_6_), .Y(men_men_n190_));
  NO3        u0168(.A(i_3_), .B(men_men_n81_), .C(men_men_n48_), .Y(men_men_n191_));
  NA2        u0169(.A(men_men_n191_), .B(men_men_n107_), .Y(men_men_n192_));
  NO3        u0170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n193_));
  NA3        u0171(.A(men_men_n193_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n194_));
  NO3        u0172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n195_));
  OAI210     u0173(.A0(men_men_n90_), .A1(i_12_), .B0(men_men_n195_), .Y(men_men_n196_));
  AOI210     u0174(.A0(men_men_n196_), .A1(men_men_n194_), .B0(men_men_n192_), .Y(men_men_n197_));
  NO2        u0175(.A(i_3_), .B(i_8_), .Y(men_men_n198_));
  NO3        u0176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n199_));
  NA3        u0177(.A(men_men_n199_), .B(men_men_n198_), .C(men_men_n39_), .Y(men_men_n200_));
  NO2        u0178(.A(men_men_n97_), .B(men_men_n56_), .Y(men_men_n201_));
  NO2        u0179(.A(i_13_), .B(i_9_), .Y(men_men_n202_));
  NAi21      u0180(.An(i_12_), .B(i_3_), .Y(men_men_n203_));
  OR2        u0181(.A(men_men_n203_), .B(men_men_n1081_), .Y(men_men_n204_));
  NO2        u0182(.A(men_men_n44_), .B(i_5_), .Y(men_men_n205_));
  NO3        u0183(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n206_));
  NA3        u0184(.A(men_men_n206_), .B(men_men_n205_), .C(i_10_), .Y(men_men_n207_));
  OAI220     u0185(.A0(men_men_n207_), .A1(men_men_n204_), .B0(men_men_n97_), .B1(men_men_n200_), .Y(men_men_n208_));
  AOI210     u0186(.A0(men_men_n208_), .A1(i_7_), .B0(men_men_n197_), .Y(men_men_n209_));
  OAI220     u0187(.A0(men_men_n209_), .A1(i_4_), .B0(men_men_n190_), .B1(men_men_n187_), .Y(men_men_n210_));
  NAi21      u0188(.An(i_12_), .B(i_7_), .Y(men_men_n211_));
  NA3        u0189(.A(i_13_), .B(men_men_n188_), .C(i_10_), .Y(men_men_n212_));
  NO2        u0190(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n213_));
  NA2        u0191(.A(i_0_), .B(i_5_), .Y(men_men_n214_));
  NA2        u0192(.A(men_men_n214_), .B(men_men_n98_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(men_men_n184_), .B0(men_men_n174_), .B1(men_men_n127_), .Y(men_men_n216_));
  NAi31      u0194(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n217_));
  NO2        u0195(.A(men_men_n35_), .B(i_13_), .Y(men_men_n218_));
  NO2        u0196(.A(men_men_n69_), .B(men_men_n26_), .Y(men_men_n219_));
  NO2        u0197(.A(men_men_n46_), .B(men_men_n61_), .Y(men_men_n220_));
  NA3        u0198(.A(men_men_n220_), .B(men_men_n219_), .C(men_men_n218_), .Y(men_men_n221_));
  INV        u0199(.A(i_13_), .Y(men_men_n222_));
  NO2        u0200(.A(i_12_), .B(men_men_n222_), .Y(men_men_n223_));
  NA3        u0201(.A(men_men_n223_), .B(men_men_n193_), .C(men_men_n191_), .Y(men_men_n224_));
  OAI210     u0202(.A0(men_men_n221_), .A1(men_men_n217_), .B0(men_men_n224_), .Y(men_men_n225_));
  AOI220     u0203(.A0(men_men_n225_), .A1(men_men_n134_), .B0(men_men_n216_), .B1(men_men_n213_), .Y(men_men_n226_));
  NO2        u0204(.A(i_12_), .B(men_men_n36_), .Y(men_men_n227_));
  NO2        u0205(.A(men_men_n177_), .B(i_4_), .Y(men_men_n228_));
  NA2        u0206(.A(men_men_n228_), .B(men_men_n227_), .Y(men_men_n229_));
  OR2        u0207(.A(i_8_), .B(i_7_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n230_), .B(men_men_n81_), .Y(men_men_n231_));
  NO2        u0209(.A(men_men_n51_), .B(i_1_), .Y(men_men_n232_));
  NA2        u0210(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  INV        u0211(.A(i_12_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n44_), .B(men_men_n234_), .Y(men_men_n235_));
  NO3        u0213(.A(men_men_n35_), .B(i_8_), .C(i_10_), .Y(men_men_n236_));
  NA2        u0214(.A(i_2_), .B(i_1_), .Y(men_men_n237_));
  NO2        u0215(.A(men_men_n233_), .B(men_men_n229_), .Y(men_men_n238_));
  NO3        u0216(.A(i_11_), .B(i_7_), .C(men_men_n36_), .Y(men_men_n239_));
  NAi21      u0217(.An(i_4_), .B(i_3_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n240_), .B(men_men_n71_), .Y(men_men_n241_));
  NO2        u0219(.A(i_0_), .B(i_6_), .Y(men_men_n242_));
  NOi41      u0220(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n243_));
  NA2        u0221(.A(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  NO2        u0222(.A(men_men_n237_), .B(men_men_n177_), .Y(men_men_n245_));
  NAi21      u0223(.An(men_men_n244_), .B(men_men_n245_), .Y(men_men_n246_));
  INV        u0224(.A(men_men_n246_), .Y(men_men_n247_));
  AOI220     u0225(.A0(men_men_n247_), .A1(men_men_n39_), .B0(men_men_n238_), .B1(men_men_n202_), .Y(men_men_n248_));
  NO2        u0226(.A(i_11_), .B(men_men_n222_), .Y(men_men_n249_));
  NOi21      u0227(.An(i_1_), .B(i_6_), .Y(men_men_n250_));
  NAi21      u0228(.An(i_3_), .B(i_7_), .Y(men_men_n251_));
  NA2        u0229(.A(men_men_n234_), .B(i_9_), .Y(men_men_n252_));
  OR4        u0230(.A(men_men_n252_), .B(men_men_n251_), .C(men_men_n250_), .D(men_men_n180_), .Y(men_men_n253_));
  NO2        u0231(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n254_));
  NO2        u0232(.A(i_12_), .B(i_3_), .Y(men_men_n255_));
  NA2        u0233(.A(men_men_n69_), .B(i_5_), .Y(men_men_n256_));
  NA2        u0234(.A(i_3_), .B(i_9_), .Y(men_men_n257_));
  NAi21      u0235(.An(i_7_), .B(i_10_), .Y(men_men_n258_));
  NO2        u0236(.A(men_men_n258_), .B(men_men_n257_), .Y(men_men_n259_));
  NA3        u0237(.A(men_men_n259_), .B(men_men_n256_), .C(men_men_n62_), .Y(men_men_n260_));
  NA2        u0238(.A(men_men_n260_), .B(men_men_n253_), .Y(men_men_n261_));
  NA3        u0239(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n262_));
  INV        u0240(.A(men_men_n135_), .Y(men_men_n263_));
  NA2        u0241(.A(men_men_n234_), .B(i_13_), .Y(men_men_n264_));
  NO2        u0242(.A(men_men_n264_), .B(men_men_n71_), .Y(men_men_n265_));
  AOI220     u0243(.A0(men_men_n265_), .A1(men_men_n263_), .B0(men_men_n261_), .B1(men_men_n249_), .Y(men_men_n266_));
  NO2        u0244(.A(men_men_n230_), .B(men_men_n36_), .Y(men_men_n267_));
  NA2        u0245(.A(i_12_), .B(i_6_), .Y(men_men_n268_));
  OR2        u0246(.A(i_13_), .B(i_9_), .Y(men_men_n269_));
  NO3        u0247(.A(men_men_n269_), .B(men_men_n268_), .C(men_men_n48_), .Y(men_men_n270_));
  NO2        u0248(.A(men_men_n240_), .B(i_2_), .Y(men_men_n271_));
  NA3        u0249(.A(men_men_n271_), .B(men_men_n270_), .C(men_men_n44_), .Y(men_men_n272_));
  NA2        u0250(.A(men_men_n249_), .B(i_9_), .Y(men_men_n273_));
  OAI210     u0251(.A0(men_men_n69_), .A1(men_men_n273_), .B0(men_men_n272_), .Y(men_men_n274_));
  NO3        u0252(.A(i_11_), .B(men_men_n222_), .C(men_men_n25_), .Y(men_men_n275_));
  NO2        u0253(.A(men_men_n251_), .B(i_8_), .Y(men_men_n276_));
  NO2        u0254(.A(i_6_), .B(men_men_n48_), .Y(men_men_n277_));
  NA3        u0255(.A(men_men_n277_), .B(men_men_n276_), .C(men_men_n275_), .Y(men_men_n278_));
  NO3        u0256(.A(men_men_n26_), .B(men_men_n81_), .C(i_5_), .Y(men_men_n279_));
  NA3        u0257(.A(men_men_n279_), .B(men_men_n267_), .C(men_men_n223_), .Y(men_men_n280_));
  AOI210     u0258(.A0(men_men_n280_), .A1(men_men_n278_), .B0(men_men_n69_), .Y(men_men_n281_));
  AOI210     u0259(.A0(men_men_n274_), .A1(men_men_n267_), .B0(men_men_n281_), .Y(men_men_n282_));
  NA4        u0260(.A(men_men_n282_), .B(men_men_n266_), .C(men_men_n248_), .D(men_men_n226_), .Y(men_men_n283_));
  NO3        u0261(.A(i_12_), .B(men_men_n222_), .C(men_men_n36_), .Y(men_men_n284_));
  INV        u0262(.A(men_men_n284_), .Y(men_men_n285_));
  NOi21      u0263(.An(men_men_n156_), .B(men_men_n81_), .Y(men_men_n286_));
  NO3        u0264(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n287_));
  AOI220     u0265(.A0(men_men_n287_), .A1(men_men_n191_), .B0(men_men_n286_), .B1(men_men_n232_), .Y(men_men_n288_));
  NO2        u0266(.A(men_men_n288_), .B(i_7_), .Y(men_men_n289_));
  NO3        u0267(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n237_), .B(i_0_), .Y(men_men_n291_));
  AOI220     u0269(.A0(men_men_n291_), .A1(men_men_n189_), .B0(men_men_n290_), .B1(men_men_n134_), .Y(men_men_n292_));
  NA2        u0270(.A(men_men_n277_), .B(men_men_n26_), .Y(men_men_n293_));
  NO2        u0271(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n294_));
  NA2        u0272(.A(i_0_), .B(i_1_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n295_), .B(i_2_), .Y(men_men_n296_));
  NO2        u0274(.A(men_men_n57_), .B(i_6_), .Y(men_men_n297_));
  NA3        u0275(.A(men_men_n297_), .B(men_men_n296_), .C(men_men_n156_), .Y(men_men_n298_));
  OAI210     u0276(.A0(men_men_n158_), .A1(men_men_n135_), .B0(men_men_n298_), .Y(men_men_n299_));
  NO3        u0277(.A(men_men_n299_), .B(men_men_n294_), .C(men_men_n289_), .Y(men_men_n300_));
  NO2        u0278(.A(i_3_), .B(i_10_), .Y(men_men_n301_));
  NA3        u0279(.A(men_men_n301_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n302_));
  NO2        u0280(.A(i_2_), .B(men_men_n95_), .Y(men_men_n303_));
  NO2        u0281(.A(i_4_), .B(i_8_), .Y(men_men_n304_));
  NOi21      u0282(.An(men_men_n214_), .B(men_men_n97_), .Y(men_men_n305_));
  NA3        u0283(.A(men_men_n305_), .B(men_men_n304_), .C(men_men_n303_), .Y(men_men_n306_));
  AN2        u0284(.A(i_3_), .B(i_10_), .Y(men_men_n307_));
  NA4        u0285(.A(men_men_n307_), .B(men_men_n193_), .C(men_men_n170_), .D(men_men_n168_), .Y(men_men_n308_));
  NO2        u0286(.A(i_5_), .B(men_men_n36_), .Y(men_men_n309_));
  NO2        u0287(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n310_));
  OR2        u0288(.A(men_men_n306_), .B(men_men_n302_), .Y(men_men_n311_));
  OAI220     u0289(.A0(men_men_n311_), .A1(i_6_), .B0(men_men_n300_), .B1(men_men_n285_), .Y(men_men_n312_));
  NO4        u0290(.A(men_men_n312_), .B(men_men_n283_), .C(men_men_n210_), .D(men_men_n161_), .Y(men_men_n313_));
  NO3        u0291(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n314_));
  NO2        u0292(.A(men_men_n57_), .B(men_men_n81_), .Y(men_men_n315_));
  NA2        u0293(.A(men_men_n291_), .B(men_men_n315_), .Y(men_men_n316_));
  NO3        u0294(.A(i_6_), .B(men_men_n188_), .C(i_7_), .Y(men_men_n317_));
  AOI210     u0295(.A0(men_men_n1084_), .A1(men_men_n316_), .B0(men_men_n163_), .Y(men_men_n318_));
  NO2        u0296(.A(i_2_), .B(i_3_), .Y(men_men_n319_));
  OR2        u0297(.A(i_0_), .B(i_5_), .Y(men_men_n320_));
  NA2        u0298(.A(men_men_n214_), .B(men_men_n320_), .Y(men_men_n321_));
  NA4        u0299(.A(men_men_n321_), .B(men_men_n231_), .C(men_men_n319_), .D(i_1_), .Y(men_men_n322_));
  NA3        u0300(.A(men_men_n291_), .B(men_men_n286_), .C(men_men_n107_), .Y(men_men_n323_));
  NAi21      u0301(.An(i_8_), .B(i_7_), .Y(men_men_n324_));
  NO2        u0302(.A(men_men_n324_), .B(i_6_), .Y(men_men_n325_));
  NO2        u0303(.A(men_men_n150_), .B(men_men_n46_), .Y(men_men_n326_));
  NA3        u0304(.A(men_men_n326_), .B(men_men_n325_), .C(men_men_n156_), .Y(men_men_n327_));
  NA3        u0305(.A(men_men_n327_), .B(men_men_n323_), .C(men_men_n322_), .Y(men_men_n328_));
  OAI210     u0306(.A0(men_men_n328_), .A1(men_men_n318_), .B0(i_4_), .Y(men_men_n329_));
  NO2        u0307(.A(i_12_), .B(i_10_), .Y(men_men_n330_));
  NOi21      u0308(.An(i_5_), .B(i_0_), .Y(men_men_n331_));
  AOI210     u0309(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n95_), .Y(men_men_n332_));
  NO4        u0310(.A(men_men_n332_), .B(i_4_), .C(men_men_n331_), .D(men_men_n122_), .Y(men_men_n333_));
  NA4        u0311(.A(men_men_n79_), .B(men_men_n35_), .C(men_men_n81_), .D(i_8_), .Y(men_men_n334_));
  NA2        u0312(.A(men_men_n333_), .B(men_men_n330_), .Y(men_men_n335_));
  NO2        u0313(.A(i_6_), .B(i_8_), .Y(men_men_n336_));
  NOi21      u0314(.An(i_0_), .B(i_2_), .Y(men_men_n337_));
  AN2        u0315(.A(men_men_n337_), .B(men_men_n336_), .Y(men_men_n338_));
  NO2        u0316(.A(i_1_), .B(i_7_), .Y(men_men_n339_));
  AO220      u0317(.A0(men_men_n339_), .A1(men_men_n338_), .B0(men_men_n325_), .B1(men_men_n232_), .Y(men_men_n340_));
  NA2        u0318(.A(men_men_n340_), .B(men_men_n41_), .Y(men_men_n341_));
  NA3        u0319(.A(men_men_n341_), .B(men_men_n335_), .C(men_men_n329_), .Y(men_men_n342_));
  NO3        u0320(.A(men_men_n230_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n343_));
  NO3        u0321(.A(men_men_n324_), .B(i_2_), .C(i_1_), .Y(men_men_n344_));
  OAI210     u0322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(i_6_), .Y(men_men_n345_));
  NA3        u0323(.A(men_men_n250_), .B(men_men_n303_), .C(men_men_n188_), .Y(men_men_n346_));
  NA2        u0324(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  NOi21      u0325(.An(men_men_n146_), .B(men_men_n98_), .Y(men_men_n348_));
  NO2        u0326(.A(men_men_n348_), .B(men_men_n119_), .Y(men_men_n349_));
  OAI210     u0327(.A0(men_men_n349_), .A1(men_men_n347_), .B0(i_3_), .Y(men_men_n350_));
  INV        u0328(.A(men_men_n79_), .Y(men_men_n351_));
  NO2        u0329(.A(men_men_n295_), .B(men_men_n76_), .Y(men_men_n352_));
  NA2        u0330(.A(men_men_n352_), .B(men_men_n126_), .Y(men_men_n353_));
  NO2        u0331(.A(men_men_n88_), .B(men_men_n188_), .Y(men_men_n354_));
  NA3        u0332(.A(men_men_n305_), .B(men_men_n354_), .C(men_men_n61_), .Y(men_men_n355_));
  AOI210     u0333(.A0(men_men_n355_), .A1(men_men_n353_), .B0(men_men_n351_), .Y(men_men_n356_));
  NO2        u0334(.A(men_men_n188_), .B(i_9_), .Y(men_men_n357_));
  NA2        u0335(.A(men_men_n357_), .B(men_men_n201_), .Y(men_men_n358_));
  NO2        u0336(.A(men_men_n358_), .B(men_men_n46_), .Y(men_men_n359_));
  NO3        u0337(.A(men_men_n359_), .B(men_men_n356_), .C(men_men_n294_), .Y(men_men_n360_));
  AOI210     u0338(.A0(men_men_n360_), .A1(men_men_n350_), .B0(men_men_n155_), .Y(men_men_n361_));
  AOI210     u0339(.A0(men_men_n342_), .A1(men_men_n314_), .B0(men_men_n361_), .Y(men_men_n362_));
  NOi32      u0340(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n363_));
  INV        u0341(.A(men_men_n363_), .Y(men_men_n364_));
  NAi21      u0342(.An(i_0_), .B(i_6_), .Y(men_men_n365_));
  NAi21      u0343(.An(i_1_), .B(i_5_), .Y(men_men_n366_));
  NA2        u0344(.A(men_men_n366_), .B(men_men_n365_), .Y(men_men_n367_));
  NA2        u0345(.A(men_men_n367_), .B(men_men_n25_), .Y(men_men_n368_));
  OAI210     u0346(.A0(men_men_n368_), .A1(men_men_n152_), .B0(men_men_n244_), .Y(men_men_n369_));
  NAi41      u0347(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n370_));
  OAI220     u0348(.A0(men_men_n370_), .A1(men_men_n366_), .B0(men_men_n217_), .B1(men_men_n152_), .Y(men_men_n371_));
  AOI210     u0349(.A0(men_men_n370_), .A1(men_men_n152_), .B0(men_men_n150_), .Y(men_men_n372_));
  NOi32      u0350(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n373_));
  NAi21      u0351(.An(i_6_), .B(i_1_), .Y(men_men_n374_));
  NA3        u0352(.A(men_men_n374_), .B(men_men_n373_), .C(men_men_n46_), .Y(men_men_n375_));
  NO2        u0353(.A(men_men_n375_), .B(i_0_), .Y(men_men_n376_));
  OR3        u0354(.A(men_men_n376_), .B(men_men_n372_), .C(men_men_n371_), .Y(men_men_n377_));
  NO2        u0355(.A(i_1_), .B(men_men_n95_), .Y(men_men_n378_));
  NAi21      u0356(.An(i_3_), .B(i_4_), .Y(men_men_n379_));
  NO2        u0357(.A(men_men_n379_), .B(i_9_), .Y(men_men_n380_));
  AN2        u0358(.A(i_6_), .B(i_7_), .Y(men_men_n381_));
  OAI210     u0359(.A0(men_men_n381_), .A1(men_men_n378_), .B0(men_men_n380_), .Y(men_men_n382_));
  NA2        u0360(.A(i_2_), .B(i_7_), .Y(men_men_n383_));
  NO2        u0361(.A(men_men_n379_), .B(i_10_), .Y(men_men_n384_));
  NA3        u0362(.A(men_men_n384_), .B(men_men_n383_), .C(men_men_n242_), .Y(men_men_n385_));
  AOI210     u0363(.A0(men_men_n385_), .A1(men_men_n382_), .B0(men_men_n180_), .Y(men_men_n386_));
  AOI210     u0364(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n387_));
  OAI210     u0365(.A0(men_men_n387_), .A1(men_men_n183_), .B0(men_men_n384_), .Y(men_men_n388_));
  AOI220     u0366(.A0(men_men_n384_), .A1(men_men_n339_), .B0(men_men_n236_), .B1(men_men_n183_), .Y(men_men_n389_));
  AOI210     u0367(.A0(men_men_n389_), .A1(men_men_n388_), .B0(i_5_), .Y(men_men_n390_));
  NO4        u0368(.A(men_men_n390_), .B(men_men_n386_), .C(men_men_n377_), .D(men_men_n369_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n391_), .B(men_men_n364_), .Y(men_men_n392_));
  NO2        u0370(.A(men_men_n57_), .B(men_men_n25_), .Y(men_men_n393_));
  AN2        u0371(.A(i_12_), .B(i_5_), .Y(men_men_n394_));
  NO2        u0372(.A(i_4_), .B(men_men_n26_), .Y(men_men_n395_));
  NA2        u0373(.A(men_men_n395_), .B(men_men_n394_), .Y(men_men_n396_));
  NO2        u0374(.A(i_11_), .B(i_6_), .Y(men_men_n397_));
  NA3        u0375(.A(men_men_n397_), .B(men_men_n326_), .C(men_men_n222_), .Y(men_men_n398_));
  NO2        u0376(.A(men_men_n398_), .B(men_men_n396_), .Y(men_men_n399_));
  NO2        u0377(.A(men_men_n240_), .B(i_5_), .Y(men_men_n400_));
  NO2        u0378(.A(i_5_), .B(i_10_), .Y(men_men_n401_));
  AOI220     u0379(.A0(men_men_n401_), .A1(men_men_n271_), .B0(men_men_n400_), .B1(men_men_n193_), .Y(men_men_n402_));
  NA2        u0380(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n403_));
  NO2        u0381(.A(men_men_n403_), .B(men_men_n402_), .Y(men_men_n404_));
  OAI210     u0382(.A0(men_men_n404_), .A1(men_men_n399_), .B0(men_men_n393_), .Y(men_men_n405_));
  NO2        u0383(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n406_));
  NO2        u0384(.A(men_men_n142_), .B(men_men_n81_), .Y(men_men_n407_));
  OAI210     u0385(.A0(men_men_n407_), .A1(men_men_n399_), .B0(men_men_n406_), .Y(men_men_n408_));
  NO3        u0386(.A(men_men_n81_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n409_));
  NO2        u0387(.A(i_3_), .B(men_men_n95_), .Y(men_men_n410_));
  NO2        u0388(.A(i_11_), .B(i_12_), .Y(men_men_n411_));
  NA2        u0389(.A(men_men_n401_), .B(men_men_n234_), .Y(men_men_n412_));
  NA3        u0390(.A(men_men_n107_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n413_));
  OAI220     u0391(.A0(men_men_n413_), .A1(men_men_n217_), .B0(men_men_n412_), .B1(men_men_n334_), .Y(men_men_n414_));
  NAi21      u0392(.An(i_13_), .B(i_0_), .Y(men_men_n415_));
  INV        u0393(.A(men_men_n415_), .Y(men_men_n416_));
  NA2        u0394(.A(men_men_n414_), .B(men_men_n416_), .Y(men_men_n417_));
  NA3        u0395(.A(men_men_n417_), .B(men_men_n408_), .C(men_men_n405_), .Y(men_men_n418_));
  NA2        u0396(.A(men_men_n44_), .B(men_men_n222_), .Y(men_men_n419_));
  NO3        u0397(.A(i_1_), .B(i_12_), .C(men_men_n81_), .Y(men_men_n420_));
  NO2        u0398(.A(i_0_), .B(i_11_), .Y(men_men_n421_));
  NOi21      u0399(.An(i_2_), .B(i_12_), .Y(men_men_n422_));
  NA2        u0400(.A(men_men_n422_), .B(i_6_), .Y(men_men_n423_));
  NO2        u0401(.A(men_men_n423_), .B(men_men_n1078_), .Y(men_men_n424_));
  NA2        u0402(.A(men_men_n134_), .B(i_9_), .Y(men_men_n425_));
  NO2        u0403(.A(men_men_n425_), .B(i_4_), .Y(men_men_n426_));
  NA2        u0404(.A(men_men_n424_), .B(men_men_n426_), .Y(men_men_n427_));
  NAi21      u0405(.An(i_9_), .B(i_4_), .Y(men_men_n428_));
  OR2        u0406(.A(i_13_), .B(i_10_), .Y(men_men_n429_));
  NO3        u0407(.A(men_men_n429_), .B(men_men_n112_), .C(men_men_n428_), .Y(men_men_n430_));
  NO2        u0408(.A(men_men_n166_), .B(men_men_n118_), .Y(men_men_n431_));
  OR2        u0409(.A(men_men_n212_), .B(men_men_n211_), .Y(men_men_n432_));
  NO2        u0410(.A(men_men_n95_), .B(men_men_n25_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n284_), .B(men_men_n433_), .Y(men_men_n434_));
  NA2        u0412(.A(men_men_n277_), .B(men_men_n206_), .Y(men_men_n435_));
  OAI220     u0413(.A0(men_men_n435_), .A1(men_men_n432_), .B0(men_men_n434_), .B1(men_men_n348_), .Y(men_men_n436_));
  INV        u0414(.A(men_men_n436_), .Y(men_men_n437_));
  AOI210     u0415(.A0(men_men_n437_), .A1(men_men_n427_), .B0(men_men_n26_), .Y(men_men_n438_));
  NA2        u0416(.A(men_men_n323_), .B(men_men_n322_), .Y(men_men_n439_));
  AOI220     u0417(.A0(men_men_n297_), .A1(men_men_n287_), .B0(men_men_n291_), .B1(men_men_n315_), .Y(men_men_n440_));
  NO2        u0418(.A(men_men_n440_), .B(men_men_n163_), .Y(men_men_n441_));
  NO2        u0419(.A(men_men_n177_), .B(men_men_n81_), .Y(men_men_n442_));
  AOI220     u0420(.A0(men_men_n442_), .A1(men_men_n296_), .B0(men_men_n279_), .B1(men_men_n206_), .Y(men_men_n443_));
  NO2        u0421(.A(men_men_n443_), .B(i_7_), .Y(men_men_n444_));
  NO3        u0422(.A(men_men_n444_), .B(men_men_n441_), .C(men_men_n439_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n191_), .B(men_men_n90_), .Y(men_men_n446_));
  NA3        u0424(.A(men_men_n326_), .B(men_men_n156_), .C(men_men_n81_), .Y(men_men_n447_));
  AOI210     u0425(.A0(men_men_n447_), .A1(men_men_n446_), .B0(men_men_n324_), .Y(men_men_n448_));
  NA2        u0426(.A(men_men_n188_), .B(i_10_), .Y(men_men_n449_));
  NA3        u0427(.A(men_men_n256_), .B(men_men_n62_), .C(i_2_), .Y(men_men_n450_));
  NA2        u0428(.A(men_men_n297_), .B(men_men_n232_), .Y(men_men_n451_));
  OAI220     u0429(.A0(men_men_n451_), .A1(men_men_n177_), .B0(men_men_n450_), .B1(men_men_n449_), .Y(men_men_n452_));
  NO2        u0430(.A(i_3_), .B(men_men_n48_), .Y(men_men_n453_));
  NA3        u0431(.A(men_men_n339_), .B(men_men_n338_), .C(men_men_n453_), .Y(men_men_n454_));
  NA2        u0432(.A(men_men_n317_), .B(men_men_n321_), .Y(men_men_n455_));
  OAI210     u0433(.A0(men_men_n455_), .A1(men_men_n184_), .B0(men_men_n454_), .Y(men_men_n456_));
  NO3        u0434(.A(men_men_n456_), .B(men_men_n452_), .C(men_men_n448_), .Y(men_men_n457_));
  AOI210     u0435(.A0(men_men_n457_), .A1(men_men_n445_), .B0(men_men_n273_), .Y(men_men_n458_));
  NO4        u0436(.A(men_men_n458_), .B(men_men_n438_), .C(men_men_n418_), .D(men_men_n392_), .Y(men_men_n459_));
  NO2        u0437(.A(men_men_n61_), .B(i_4_), .Y(men_men_n460_));
  NO2        u0438(.A(men_men_n69_), .B(i_13_), .Y(men_men_n461_));
  NA3        u0439(.A(men_men_n461_), .B(men_men_n460_), .C(i_2_), .Y(men_men_n462_));
  NO2        u0440(.A(i_10_), .B(i_9_), .Y(men_men_n463_));
  NAi21      u0441(.An(i_12_), .B(i_8_), .Y(men_men_n464_));
  NO2        u0442(.A(men_men_n464_), .B(i_3_), .Y(men_men_n465_));
  NA2        u0443(.A(men_men_n465_), .B(men_men_n463_), .Y(men_men_n466_));
  NA2        u0444(.A(men_men_n1086_), .B(men_men_n98_), .Y(men_men_n467_));
  OAI220     u0445(.A0(men_men_n467_), .A1(men_men_n200_), .B0(men_men_n466_), .B1(men_men_n462_), .Y(men_men_n468_));
  NA2        u0446(.A(men_men_n310_), .B(i_0_), .Y(men_men_n469_));
  NO3        u0447(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n470_));
  NA2        u0448(.A(men_men_n268_), .B(men_men_n91_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n471_), .B(men_men_n470_), .Y(men_men_n472_));
  NA2        u0450(.A(i_8_), .B(i_9_), .Y(men_men_n473_));
  AOI210     u0451(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n474_));
  OR2        u0452(.A(men_men_n474_), .B(men_men_n473_), .Y(men_men_n475_));
  NA2        u0453(.A(men_men_n284_), .B(men_men_n201_), .Y(men_men_n476_));
  OAI220     u0454(.A0(men_men_n476_), .A1(men_men_n475_), .B0(men_men_n472_), .B1(men_men_n469_), .Y(men_men_n477_));
  NA2        u0455(.A(men_men_n249_), .B(men_men_n309_), .Y(men_men_n478_));
  NO3        u0456(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n479_));
  INV        u0457(.A(men_men_n479_), .Y(men_men_n480_));
  NA3        u0458(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n481_));
  NA4        u0459(.A(men_men_n137_), .B(men_men_n110_), .C(men_men_n75_), .D(men_men_n23_), .Y(men_men_n482_));
  OAI220     u0460(.A0(men_men_n482_), .A1(men_men_n481_), .B0(men_men_n480_), .B1(men_men_n478_), .Y(men_men_n483_));
  NO3        u0461(.A(men_men_n483_), .B(men_men_n477_), .C(men_men_n468_), .Y(men_men_n484_));
  NA2        u0462(.A(men_men_n296_), .B(men_men_n102_), .Y(men_men_n485_));
  OR2        u0463(.A(men_men_n485_), .B(men_men_n1081_), .Y(men_men_n486_));
  OA210      u0464(.A0(men_men_n358_), .A1(men_men_n95_), .B0(men_men_n298_), .Y(men_men_n487_));
  OA220      u0465(.A0(men_men_n487_), .A1(men_men_n155_), .B0(men_men_n486_), .B1(men_men_n229_), .Y(men_men_n488_));
  NA2        u0466(.A(men_men_n90_), .B(i_13_), .Y(men_men_n489_));
  NA2        u0467(.A(men_men_n442_), .B(men_men_n393_), .Y(men_men_n490_));
  NO2        u0468(.A(i_2_), .B(i_13_), .Y(men_men_n491_));
  NO2        u0469(.A(men_men_n490_), .B(men_men_n489_), .Y(men_men_n492_));
  NO3        u0470(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n493_));
  NO2        u0471(.A(i_6_), .B(i_7_), .Y(men_men_n494_));
  NA2        u0472(.A(men_men_n494_), .B(men_men_n493_), .Y(men_men_n495_));
  OR2        u0473(.A(i_11_), .B(i_8_), .Y(men_men_n496_));
  NOi21      u0474(.An(i_2_), .B(i_7_), .Y(men_men_n497_));
  NAi31      u0475(.An(men_men_n496_), .B(men_men_n497_), .C(men_men_n1080_), .Y(men_men_n498_));
  NO2        u0476(.A(men_men_n429_), .B(i_6_), .Y(men_men_n499_));
  NA3        u0477(.A(men_men_n499_), .B(men_men_n460_), .C(men_men_n71_), .Y(men_men_n500_));
  NO2        u0478(.A(men_men_n500_), .B(men_men_n498_), .Y(men_men_n501_));
  NO2        u0479(.A(i_6_), .B(i_10_), .Y(men_men_n502_));
  NA3        u0480(.A(men_men_n243_), .B(men_men_n165_), .C(men_men_n126_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n504_));
  NO2        u0482(.A(men_men_n150_), .B(i_3_), .Y(men_men_n505_));
  NAi31      u0483(.An(men_men_n504_), .B(men_men_n505_), .C(men_men_n223_), .Y(men_men_n506_));
  NA3        u0484(.A(men_men_n406_), .B(men_men_n173_), .C(men_men_n141_), .Y(men_men_n507_));
  NA3        u0485(.A(men_men_n507_), .B(men_men_n506_), .C(men_men_n503_), .Y(men_men_n508_));
  NO3        u0486(.A(men_men_n508_), .B(men_men_n501_), .C(men_men_n492_), .Y(men_men_n509_));
  NA2        u0487(.A(men_men_n479_), .B(men_men_n401_), .Y(men_men_n510_));
  NO2        u0488(.A(men_men_n510_), .B(men_men_n221_), .Y(men_men_n511_));
  NAi21      u0489(.An(men_men_n212_), .B(men_men_n411_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n339_), .B(men_men_n214_), .Y(men_men_n513_));
  NO2        u0491(.A(men_men_n26_), .B(i_5_), .Y(men_men_n514_));
  NO2        u0492(.A(i_0_), .B(men_men_n81_), .Y(men_men_n515_));
  NA3        u0493(.A(men_men_n515_), .B(men_men_n514_), .C(men_men_n134_), .Y(men_men_n516_));
  OR3        u0494(.A(i_4_), .B(men_men_n37_), .C(men_men_n46_), .Y(men_men_n517_));
  OAI220     u0495(.A0(men_men_n517_), .A1(men_men_n516_), .B0(men_men_n513_), .B1(men_men_n512_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n27_), .B(i_10_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n314_), .B(men_men_n236_), .Y(men_men_n520_));
  OAI220     u0498(.A0(men_men_n520_), .A1(men_men_n450_), .B0(men_men_n519_), .B1(men_men_n489_), .Y(men_men_n521_));
  NA4        u0499(.A(men_men_n307_), .B(men_men_n220_), .C(men_men_n69_), .D(men_men_n234_), .Y(men_men_n522_));
  NO2        u0500(.A(men_men_n522_), .B(men_men_n495_), .Y(men_men_n523_));
  NO4        u0501(.A(men_men_n523_), .B(men_men_n521_), .C(men_men_n518_), .D(men_men_n511_), .Y(men_men_n524_));
  NA4        u0502(.A(men_men_n524_), .B(men_men_n509_), .C(men_men_n488_), .D(men_men_n484_), .Y(men_men_n525_));
  NA3        u0503(.A(men_men_n307_), .B(men_men_n170_), .C(men_men_n168_), .Y(men_men_n526_));
  OAI210     u0504(.A0(men_men_n302_), .A1(men_men_n175_), .B0(men_men_n526_), .Y(men_men_n527_));
  AN2        u0505(.A(men_men_n287_), .B(men_men_n231_), .Y(men_men_n528_));
  NA2        u0506(.A(men_men_n528_), .B(men_men_n527_), .Y(men_men_n529_));
  NA2        u0507(.A(men_men_n117_), .B(men_men_n106_), .Y(men_men_n530_));
  AO220      u0508(.A0(men_men_n530_), .A1(men_men_n470_), .B0(men_men_n430_), .B1(i_6_), .Y(men_men_n531_));
  NA2        u0509(.A(men_men_n314_), .B(men_men_n157_), .Y(men_men_n532_));
  OAI210     u0510(.A0(men_men_n532_), .A1(men_men_n229_), .B0(men_men_n308_), .Y(men_men_n533_));
  AOI220     u0511(.A0(men_men_n533_), .A1(men_men_n325_), .B0(men_men_n531_), .B1(men_men_n310_), .Y(men_men_n534_));
  NA4        u0512(.A(men_men_n461_), .B(men_men_n460_), .C(men_men_n198_), .D(i_2_), .Y(men_men_n535_));
  INV        u0513(.A(men_men_n535_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n394_), .B(men_men_n222_), .Y(men_men_n537_));
  NA2        u0515(.A(men_men_n363_), .B(men_men_n69_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n381_), .B(men_men_n373_), .Y(men_men_n539_));
  AO210      u0517(.A0(men_men_n538_), .A1(men_men_n537_), .B0(men_men_n539_), .Y(men_men_n540_));
  NO2        u0518(.A(men_men_n35_), .B(i_8_), .Y(men_men_n541_));
  NAi41      u0519(.An(men_men_n538_), .B(men_men_n502_), .C(men_men_n541_), .D(men_men_n46_), .Y(men_men_n542_));
  AOI210     u0520(.A0(men_men_n38_), .A1(i_13_), .B0(men_men_n430_), .Y(men_men_n543_));
  NA3        u0521(.A(men_men_n543_), .B(men_men_n542_), .C(men_men_n540_), .Y(men_men_n544_));
  AOI210     u0522(.A0(men_men_n536_), .A1(men_men_n199_), .B0(men_men_n544_), .Y(men_men_n545_));
  NA2        u0523(.A(men_men_n256_), .B(men_men_n62_), .Y(men_men_n546_));
  OAI210     u0524(.A0(i_8_), .A1(men_men_n546_), .B0(men_men_n128_), .Y(men_men_n547_));
  AOI210     u0525(.A0(men_men_n189_), .A1(i_9_), .B0(men_men_n267_), .Y(men_men_n548_));
  NO2        u0526(.A(men_men_n548_), .B(men_men_n194_), .Y(men_men_n549_));
  OR2        u0527(.A(men_men_n177_), .B(i_4_), .Y(men_men_n550_));
  NO2        u0528(.A(men_men_n550_), .B(men_men_n81_), .Y(men_men_n551_));
  AOI220     u0529(.A0(men_men_n551_), .A1(men_men_n549_), .B0(men_men_n547_), .B1(men_men_n431_), .Y(men_men_n552_));
  NA4        u0530(.A(men_men_n552_), .B(men_men_n545_), .C(men_men_n534_), .D(men_men_n529_), .Y(men_men_n553_));
  NA2        u0531(.A(men_men_n400_), .B(men_men_n296_), .Y(men_men_n554_));
  OAI210     u0532(.A0(men_men_n396_), .A1(men_men_n162_), .B0(men_men_n554_), .Y(men_men_n555_));
  NO2        u0533(.A(i_12_), .B(men_men_n188_), .Y(men_men_n556_));
  NA2        u0534(.A(men_men_n556_), .B(men_men_n222_), .Y(men_men_n557_));
  NA3        u0535(.A(men_men_n502_), .B(men_men_n168_), .C(men_men_n27_), .Y(men_men_n558_));
  NO3        u0536(.A(men_men_n558_), .B(men_men_n557_), .C(men_men_n485_), .Y(men_men_n559_));
  NOi31      u0537(.An(men_men_n317_), .B(men_men_n429_), .C(men_men_n37_), .Y(men_men_n560_));
  OAI210     u0538(.A0(men_men_n560_), .A1(men_men_n559_), .B0(men_men_n555_), .Y(men_men_n561_));
  NO2        u0539(.A(i_8_), .B(i_7_), .Y(men_men_n562_));
  OAI210     u0540(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n563_), .B(men_men_n220_), .Y(men_men_n564_));
  AOI220     u0542(.A0(men_men_n326_), .A1(men_men_n39_), .B0(men_men_n232_), .B1(men_men_n202_), .Y(men_men_n565_));
  OAI220     u0543(.A0(men_men_n565_), .A1(men_men_n550_), .B0(men_men_n564_), .B1(men_men_n240_), .Y(men_men_n566_));
  NA2        u0544(.A(men_men_n44_), .B(i_10_), .Y(men_men_n567_));
  NO2        u0545(.A(men_men_n567_), .B(i_6_), .Y(men_men_n568_));
  NA3        u0546(.A(men_men_n568_), .B(men_men_n566_), .C(men_men_n562_), .Y(men_men_n569_));
  AOI220     u0547(.A0(men_men_n442_), .A1(men_men_n326_), .B0(men_men_n245_), .B1(men_men_n242_), .Y(men_men_n570_));
  OAI220     u0548(.A0(men_men_n570_), .A1(men_men_n264_), .B0(men_men_n489_), .B1(men_men_n127_), .Y(men_men_n571_));
  NA2        u0549(.A(men_men_n571_), .B(men_men_n267_), .Y(men_men_n572_));
  NOi31      u0550(.An(men_men_n291_), .B(men_men_n302_), .C(men_men_n175_), .Y(men_men_n573_));
  NA3        u0551(.A(men_men_n307_), .B(men_men_n168_), .C(men_men_n90_), .Y(men_men_n574_));
  NO2        u0552(.A(men_men_n218_), .B(men_men_n44_), .Y(men_men_n575_));
  NO2        u0553(.A(men_men_n150_), .B(i_5_), .Y(men_men_n576_));
  NA3        u0554(.A(men_men_n576_), .B(men_men_n419_), .C(men_men_n319_), .Y(men_men_n577_));
  OAI210     u0555(.A0(men_men_n577_), .A1(men_men_n575_), .B0(men_men_n574_), .Y(men_men_n578_));
  OAI210     u0556(.A0(men_men_n578_), .A1(men_men_n573_), .B0(men_men_n479_), .Y(men_men_n579_));
  NA4        u0557(.A(men_men_n579_), .B(men_men_n572_), .C(men_men_n569_), .D(men_men_n561_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n284_), .B(men_men_n79_), .Y(men_men_n581_));
  AOI210     u0559(.A0(i_11_), .A1(men_men_n353_), .B0(men_men_n581_), .Y(men_men_n582_));
  NA2        u0560(.A(men_men_n297_), .B(men_men_n287_), .Y(men_men_n583_));
  NO2        u0561(.A(men_men_n583_), .B(men_men_n167_), .Y(men_men_n584_));
  NA2        u0562(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n585_));
  NA2        u0563(.A(men_men_n463_), .B(men_men_n218_), .Y(men_men_n586_));
  NO2        u0564(.A(men_men_n585_), .B(men_men_n586_), .Y(men_men_n587_));
  NA2        u0565(.A(i_0_), .B(men_men_n48_), .Y(men_men_n588_));
  NA3        u0566(.A(men_men_n556_), .B(men_men_n275_), .C(men_men_n588_), .Y(men_men_n589_));
  NO2        u0567(.A(men_men_n1085_), .B(men_men_n589_), .Y(men_men_n590_));
  NO4        u0568(.A(men_men_n590_), .B(men_men_n587_), .C(men_men_n584_), .D(men_men_n582_), .Y(men_men_n591_));
  NO4        u0569(.A(men_men_n250_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n592_));
  NO3        u0570(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n593_));
  NO2        u0571(.A(men_men_n230_), .B(men_men_n35_), .Y(men_men_n594_));
  AN2        u0572(.A(men_men_n594_), .B(men_men_n593_), .Y(men_men_n595_));
  AN2        u0573(.A(men_men_n592_), .B(men_men_n363_), .Y(men_men_n596_));
  NO2        u0574(.A(men_men_n429_), .B(i_1_), .Y(men_men_n597_));
  NOi31      u0575(.An(men_men_n597_), .B(men_men_n471_), .C(men_men_n69_), .Y(men_men_n598_));
  AN3        u0576(.A(men_men_n598_), .B(men_men_n426_), .C(i_2_), .Y(men_men_n599_));
  NO2        u0577(.A(men_men_n440_), .B(men_men_n171_), .Y(men_men_n600_));
  NO3        u0578(.A(men_men_n600_), .B(men_men_n599_), .C(men_men_n596_), .Y(men_men_n601_));
  NOi21      u0579(.An(i_10_), .B(i_6_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n81_), .B(men_men_n25_), .Y(men_men_n603_));
  AOI220     u0581(.A0(men_men_n284_), .A1(men_men_n603_), .B0(men_men_n275_), .B1(men_men_n602_), .Y(men_men_n604_));
  NO2        u0582(.A(men_men_n604_), .B(men_men_n469_), .Y(men_men_n605_));
  NA2        u0583(.A(men_men_n317_), .B(men_men_n157_), .Y(men_men_n606_));
  AOI220     u0584(.A0(men_men_n606_), .A1(men_men_n451_), .B0(men_men_n178_), .B1(men_men_n176_), .Y(men_men_n607_));
  NO2        u0585(.A(men_men_n193_), .B(men_men_n36_), .Y(men_men_n608_));
  NOi31      u0586(.An(men_men_n138_), .B(men_men_n608_), .C(men_men_n334_), .Y(men_men_n609_));
  NO3        u0587(.A(men_men_n609_), .B(men_men_n607_), .C(men_men_n605_), .Y(men_men_n610_));
  NO2        u0588(.A(men_men_n538_), .B(men_men_n389_), .Y(men_men_n611_));
  INV        u0589(.A(men_men_n319_), .Y(men_men_n612_));
  NO2        u0590(.A(i_12_), .B(men_men_n81_), .Y(men_men_n613_));
  NA3        u0591(.A(men_men_n613_), .B(men_men_n275_), .C(men_men_n588_), .Y(men_men_n614_));
  NA3        u0592(.A(men_men_n397_), .B(men_men_n284_), .C(men_men_n214_), .Y(men_men_n615_));
  AOI210     u0593(.A0(men_men_n615_), .A1(men_men_n614_), .B0(men_men_n612_), .Y(men_men_n616_));
  NA2        u0594(.A(men_men_n168_), .B(i_0_), .Y(men_men_n617_));
  NO3        u0595(.A(men_men_n617_), .B(men_men_n345_), .C(men_men_n302_), .Y(men_men_n618_));
  OR2        u0596(.A(i_2_), .B(i_5_), .Y(men_men_n619_));
  BUFFER     u0597(.A(men_men_n619_), .Y(men_men_n620_));
  AOI210     u0598(.A0(men_men_n383_), .A1(men_men_n242_), .B0(men_men_n193_), .Y(men_men_n621_));
  AOI210     u0599(.A0(men_men_n621_), .A1(men_men_n620_), .B0(men_men_n512_), .Y(men_men_n622_));
  NO4        u0600(.A(men_men_n622_), .B(men_men_n618_), .C(men_men_n616_), .D(men_men_n611_), .Y(men_men_n623_));
  NA4        u0601(.A(men_men_n623_), .B(men_men_n610_), .C(men_men_n601_), .D(men_men_n591_), .Y(men_men_n624_));
  NO4        u0602(.A(men_men_n624_), .B(men_men_n580_), .C(men_men_n553_), .D(men_men_n525_), .Y(men_men_n625_));
  NA4        u0603(.A(men_men_n625_), .B(men_men_n459_), .C(men_men_n362_), .D(men_men_n313_), .Y(men7));
  NO2        u0604(.A(men_men_n88_), .B(men_men_n52_), .Y(men_men_n627_));
  NO2        u0605(.A(men_men_n102_), .B(men_men_n86_), .Y(men_men_n628_));
  NA2        u0606(.A(men_men_n395_), .B(men_men_n628_), .Y(men_men_n629_));
  NA2        u0607(.A(men_men_n502_), .B(men_men_n79_), .Y(men_men_n630_));
  OAI210     u0608(.A0(men_men_n1082_), .A1(men_men_n630_), .B0(men_men_n629_), .Y(men_men_n631_));
  NA3        u0609(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n632_));
  NA2        u0610(.A(i_12_), .B(i_8_), .Y(men_men_n633_));
  AOI210     u0611(.A0(men_men_n633_), .A1(men_men_n99_), .B0(men_men_n632_), .Y(men_men_n634_));
  NA2        u0612(.A(i_2_), .B(men_men_n81_), .Y(men_men_n635_));
  OAI210     u0613(.A0(men_men_n84_), .A1(men_men_n198_), .B0(men_men_n199_), .Y(men_men_n636_));
  NO2        u0614(.A(i_7_), .B(men_men_n36_), .Y(men_men_n637_));
  NA2        u0615(.A(i_4_), .B(i_8_), .Y(men_men_n638_));
  NO2        u0616(.A(men_men_n307_), .B(men_men_n637_), .Y(men_men_n639_));
  OAI220     u0617(.A0(men_men_n639_), .A1(men_men_n635_), .B0(men_men_n636_), .B1(i_13_), .Y(men_men_n640_));
  NO4        u0618(.A(men_men_n640_), .B(men_men_n634_), .C(men_men_n631_), .D(men_men_n627_), .Y(men_men_n641_));
  AOI210     u0619(.A0(men_men_n122_), .A1(men_men_n60_), .B0(i_10_), .Y(men_men_n642_));
  AOI210     u0620(.A0(men_men_n642_), .A1(men_men_n234_), .B0(men_men_n154_), .Y(men_men_n643_));
  OR2        u0621(.A(i_6_), .B(i_10_), .Y(men_men_n644_));
  NO2        u0622(.A(men_men_n644_), .B(men_men_n23_), .Y(men_men_n645_));
  OR3        u0623(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n646_));
  NO2        u0624(.A(men_men_n646_), .B(i_8_), .Y(men_men_n647_));
  INV        u0625(.A(men_men_n195_), .Y(men_men_n648_));
  OA220      u0626(.A0(men_men_n646_), .A1(men_men_n612_), .B0(men_men_n643_), .B1(men_men_n269_), .Y(men_men_n649_));
  AOI210     u0627(.A0(men_men_n649_), .A1(men_men_n641_), .B0(men_men_n61_), .Y(men_men_n650_));
  NOi21      u0628(.An(i_11_), .B(i_7_), .Y(men_men_n651_));
  AO210      u0629(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n652_), .B(men_men_n651_), .Y(men_men_n653_));
  NA3        u0631(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n654_));
  NAi21      u0632(.An(men_men_n654_), .B(i_11_), .Y(men_men_n655_));
  NO2        u0633(.A(men_men_n655_), .B(men_men_n61_), .Y(men_men_n656_));
  NA2        u0634(.A(men_men_n83_), .B(men_men_n61_), .Y(men_men_n657_));
  AO210      u0635(.A0(men_men_n657_), .A1(men_men_n389_), .B0(men_men_n40_), .Y(men_men_n658_));
  NO3        u0636(.A(men_men_n258_), .B(men_men_n203_), .C(i_8_), .Y(men_men_n659_));
  OAI210     u0637(.A0(men_men_n659_), .A1(men_men_n223_), .B0(men_men_n61_), .Y(men_men_n660_));
  NA2        u0638(.A(men_men_n422_), .B(men_men_n30_), .Y(men_men_n661_));
  OR2        u0639(.A(men_men_n203_), .B(men_men_n102_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(men_men_n661_), .Y(men_men_n663_));
  NO2        u0641(.A(men_men_n61_), .B(i_9_), .Y(men_men_n664_));
  NO2        u0642(.A(men_men_n664_), .B(i_4_), .Y(men_men_n665_));
  NA2        u0643(.A(men_men_n665_), .B(men_men_n663_), .Y(men_men_n666_));
  NO2        u0644(.A(i_1_), .B(i_12_), .Y(men_men_n667_));
  NA2        u0645(.A(men_men_n667_), .B(men_men_n104_), .Y(men_men_n668_));
  NA4        u0646(.A(men_men_n668_), .B(men_men_n666_), .C(men_men_n660_), .D(men_men_n658_), .Y(men_men_n669_));
  OAI210     u0647(.A0(men_men_n669_), .A1(men_men_n656_), .B0(i_6_), .Y(men_men_n670_));
  OAI210     u0648(.A0(men_men_n654_), .A1(men_men_n102_), .B0(men_men_n481_), .Y(men_men_n671_));
  NA2        u0649(.A(men_men_n671_), .B(men_men_n613_), .Y(men_men_n672_));
  NO2        u0650(.A(i_6_), .B(i_11_), .Y(men_men_n673_));
  NA2        u0651(.A(men_men_n672_), .B(men_men_n472_), .Y(men_men_n674_));
  NO4        u0652(.A(men_men_n211_), .B(men_men_n122_), .C(i_13_), .D(men_men_n81_), .Y(men_men_n675_));
  INV        u0653(.A(men_men_n675_), .Y(men_men_n676_));
  NA2        u0654(.A(men_men_n234_), .B(i_6_), .Y(men_men_n677_));
  NO3        u0655(.A(men_men_n644_), .B(men_men_n230_), .C(men_men_n23_), .Y(men_men_n678_));
  AOI210     u0656(.A0(i_1_), .A1(men_men_n259_), .B0(men_men_n678_), .Y(men_men_n679_));
  OAI210     u0657(.A0(men_men_n679_), .A1(men_men_n44_), .B0(men_men_n676_), .Y(men_men_n680_));
  NA3        u0658(.A(men_men_n562_), .B(i_11_), .C(men_men_n35_), .Y(men_men_n681_));
  NA3        u0659(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n682_));
  NO2        u0660(.A(men_men_n46_), .B(i_1_), .Y(men_men_n683_));
  NA3        u0661(.A(men_men_n683_), .B(men_men_n268_), .C(men_men_n44_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n684_), .B(men_men_n682_), .Y(men_men_n685_));
  NA3        u0663(.A(men_men_n664_), .B(men_men_n319_), .C(i_6_), .Y(men_men_n686_));
  NO2        u0664(.A(men_men_n686_), .B(men_men_n23_), .Y(men_men_n687_));
  NA2        u0665(.A(men_men_n683_), .B(men_men_n268_), .Y(men_men_n688_));
  NO2        u0666(.A(i_11_), .B(men_men_n36_), .Y(men_men_n689_));
  NA2        u0667(.A(men_men_n689_), .B(men_men_n24_), .Y(men_men_n690_));
  NO2        u0668(.A(men_men_n690_), .B(men_men_n688_), .Y(men_men_n691_));
  OR3        u0669(.A(men_men_n691_), .B(men_men_n687_), .C(men_men_n685_), .Y(men_men_n692_));
  NO3        u0670(.A(men_men_n692_), .B(men_men_n680_), .C(men_men_n674_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n234_), .B(men_men_n95_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n694_), .B(men_men_n651_), .Y(men_men_n695_));
  NA2        u0673(.A(men_men_n695_), .B(i_1_), .Y(men_men_n696_));
  NO2        u0674(.A(men_men_n696_), .B(men_men_n646_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n428_), .B(men_men_n81_), .Y(men_men_n698_));
  NA2        u0676(.A(men_men_n697_), .B(men_men_n46_), .Y(men_men_n699_));
  NA2        u0677(.A(i_3_), .B(men_men_n188_), .Y(men_men_n700_));
  NO2        u0678(.A(men_men_n230_), .B(men_men_n44_), .Y(men_men_n701_));
  NO3        u0679(.A(men_men_n701_), .B(men_men_n310_), .C(men_men_n235_), .Y(men_men_n702_));
  NO2        u0680(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n703_));
  NO2        u0681(.A(men_men_n81_), .B(i_9_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n704_), .B(men_men_n61_), .Y(men_men_n705_));
  NO2        u0683(.A(men_men_n705_), .B(men_men_n667_), .Y(men_men_n706_));
  NO4        u0684(.A(men_men_n706_), .B(men_men_n1088_), .C(men_men_n702_), .D(i_4_), .Y(men_men_n707_));
  NA2        u0685(.A(i_1_), .B(i_3_), .Y(men_men_n708_));
  NO2        u0686(.A(men_men_n473_), .B(men_men_n88_), .Y(men_men_n709_));
  AOI210     u0687(.A0(men_men_n701_), .A1(men_men_n602_), .B0(men_men_n709_), .Y(men_men_n710_));
  NO2        u0688(.A(men_men_n710_), .B(men_men_n708_), .Y(men_men_n711_));
  NO2        u0689(.A(men_men_n711_), .B(men_men_n707_), .Y(men_men_n712_));
  NA4        u0690(.A(men_men_n712_), .B(men_men_n699_), .C(men_men_n693_), .D(men_men_n670_), .Y(men_men_n713_));
  NO3        u0691(.A(men_men_n496_), .B(i_3_), .C(i_7_), .Y(men_men_n714_));
  NOi21      u0692(.An(men_men_n714_), .B(i_10_), .Y(men_men_n715_));
  OA210      u0693(.A0(men_men_n715_), .A1(men_men_n243_), .B0(men_men_n81_), .Y(men_men_n716_));
  NA2        u0694(.A(men_men_n381_), .B(men_men_n380_), .Y(men_men_n717_));
  NA3        u0695(.A(men_men_n502_), .B(men_men_n541_), .C(men_men_n46_), .Y(men_men_n718_));
  NO3        u0696(.A(men_men_n497_), .B(men_men_n638_), .C(men_men_n81_), .Y(men_men_n719_));
  NA2        u0697(.A(men_men_n719_), .B(men_men_n25_), .Y(men_men_n720_));
  NA3        u0698(.A(men_men_n154_), .B(men_men_n79_), .C(men_men_n81_), .Y(men_men_n721_));
  NA4        u0699(.A(men_men_n721_), .B(men_men_n720_), .C(men_men_n718_), .D(men_men_n717_), .Y(men_men_n722_));
  OAI210     u0700(.A0(men_men_n722_), .A1(men_men_n716_), .B0(i_1_), .Y(men_men_n723_));
  NO2        u0701(.A(men_men_n686_), .B(men_men_n464_), .Y(men_men_n724_));
  INV        u0702(.A(men_men_n724_), .Y(men_men_n725_));
  AOI210     u0703(.A0(men_men_n725_), .A1(men_men_n723_), .B0(i_13_), .Y(men_men_n726_));
  OR2        u0704(.A(i_11_), .B(i_7_), .Y(men_men_n727_));
  NA3        u0705(.A(men_men_n727_), .B(men_men_n100_), .C(men_men_n132_), .Y(men_men_n728_));
  AOI220     u0706(.A0(men_men_n491_), .A1(men_men_n154_), .B0(men_men_n1086_), .B1(men_men_n132_), .Y(men_men_n729_));
  OAI210     u0707(.A0(men_men_n729_), .A1(men_men_n44_), .B0(men_men_n728_), .Y(men_men_n730_));
  NO2        u0708(.A(men_men_n497_), .B(men_men_n24_), .Y(men_men_n731_));
  AOI220     u0709(.A0(men_men_n731_), .A1(men_men_n698_), .B0(men_men_n243_), .B1(men_men_n125_), .Y(men_men_n732_));
  NO2        u0710(.A(men_men_n732_), .B(men_men_n40_), .Y(men_men_n733_));
  AOI210     u0711(.A0(men_men_n730_), .A1(men_men_n336_), .B0(men_men_n733_), .Y(men_men_n734_));
  NA2        u0712(.A(i_7_), .B(men_men_n68_), .Y(men_men_n735_));
  NO2        u0713(.A(men_men_n735_), .B(men_men_n240_), .Y(men_men_n736_));
  AOI210     u0714(.A0(men_men_n464_), .A1(men_men_n35_), .B0(i_13_), .Y(men_men_n737_));
  NOi31      u0715(.An(men_men_n737_), .B(men_men_n630_), .C(men_men_n44_), .Y(men_men_n738_));
  NO2        u0716(.A(men_men_n682_), .B(men_men_n109_), .Y(men_men_n739_));
  INV        u0717(.A(men_men_n739_), .Y(men_men_n740_));
  NO2        u0718(.A(men_men_n740_), .B(men_men_n67_), .Y(men_men_n741_));
  NO3        u0719(.A(men_men_n67_), .B(men_men_n31_), .C(men_men_n95_), .Y(men_men_n742_));
  NA2        u0720(.A(men_men_n26_), .B(men_men_n188_), .Y(men_men_n743_));
  NA2        u0721(.A(men_men_n743_), .B(i_7_), .Y(men_men_n744_));
  NO3        u0722(.A(men_men_n497_), .B(men_men_n234_), .C(men_men_n81_), .Y(men_men_n745_));
  AOI210     u0723(.A0(men_men_n745_), .A1(men_men_n744_), .B0(men_men_n742_), .Y(men_men_n746_));
  NA2        u0724(.A(men_men_n397_), .B(men_men_n683_), .Y(men_men_n747_));
  OAI220     u0725(.A0(men_men_n747_), .A1(men_men_n633_), .B0(men_men_n746_), .B1(men_men_n648_), .Y(men_men_n748_));
  NO4        u0726(.A(men_men_n748_), .B(men_men_n741_), .C(men_men_n738_), .D(men_men_n736_), .Y(men_men_n749_));
  OR2        u0727(.A(i_11_), .B(i_6_), .Y(men_men_n750_));
  NA3        u0728(.A(i_12_), .B(men_men_n743_), .C(i_7_), .Y(men_men_n751_));
  NO2        u0729(.A(men_men_n751_), .B(men_men_n750_), .Y(men_men_n752_));
  NA2        u0730(.A(men_men_n673_), .B(i_13_), .Y(men_men_n753_));
  NA2        u0731(.A(men_men_n96_), .B(men_men_n743_), .Y(men_men_n754_));
  NAi21      u0732(.An(i_11_), .B(i_12_), .Y(men_men_n755_));
  NOi41      u0733(.An(men_men_n105_), .B(men_men_n755_), .C(i_13_), .D(men_men_n81_), .Y(men_men_n756_));
  NO3        u0734(.A(men_men_n497_), .B(men_men_n613_), .C(men_men_n638_), .Y(men_men_n757_));
  AOI220     u0735(.A0(men_men_n757_), .A1(men_men_n314_), .B0(men_men_n756_), .B1(men_men_n754_), .Y(men_men_n758_));
  NA2        u0736(.A(men_men_n758_), .B(men_men_n753_), .Y(men_men_n759_));
  OAI210     u0737(.A0(men_men_n759_), .A1(men_men_n752_), .B0(men_men_n61_), .Y(men_men_n760_));
  NO2        u0738(.A(i_2_), .B(i_12_), .Y(men_men_n761_));
  NA2        u0739(.A(men_men_n378_), .B(men_men_n761_), .Y(men_men_n762_));
  OAI210     u0740(.A0(i_8_), .A1(men_men_n380_), .B0(men_men_n378_), .Y(men_men_n763_));
  NO2        u0741(.A(men_men_n122_), .B(i_2_), .Y(men_men_n764_));
  NA2        u0742(.A(men_men_n764_), .B(men_men_n667_), .Y(men_men_n765_));
  NA3        u0743(.A(men_men_n765_), .B(men_men_n763_), .C(men_men_n762_), .Y(men_men_n766_));
  NA3        u0744(.A(men_men_n766_), .B(men_men_n45_), .C(men_men_n222_), .Y(men_men_n767_));
  NA4        u0745(.A(men_men_n767_), .B(men_men_n760_), .C(men_men_n749_), .D(men_men_n734_), .Y(men_men_n768_));
  OR4        u0746(.A(men_men_n768_), .B(men_men_n726_), .C(men_men_n713_), .D(men_men_n650_), .Y(men5));
  AOI210     u0747(.A0(men_men_n695_), .A1(men_men_n271_), .B0(men_men_n431_), .Y(men_men_n770_));
  NA3        u0748(.A(men_men_n24_), .B(men_men_n761_), .C(men_men_n102_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n771_), .B(men_men_n770_), .Y(men_men_n772_));
  NO3        u0750(.A(i_11_), .B(men_men_n234_), .C(i_13_), .Y(men_men_n773_));
  NO2        u0751(.A(men_men_n119_), .B(men_men_n23_), .Y(men_men_n774_));
  NA2        u0752(.A(i_12_), .B(i_8_), .Y(men_men_n775_));
  INV        u0753(.A(men_men_n463_), .Y(men_men_n776_));
  INV        u0754(.A(men_men_n772_), .Y(men_men_n777_));
  INV        u0755(.A(men_men_n165_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n473_), .B(men_men_n26_), .Y(men_men_n779_));
  NO2        u0757(.A(men_men_n779_), .B(men_men_n433_), .Y(men_men_n780_));
  NA2        u0758(.A(men_men_n780_), .B(i_2_), .Y(men_men_n781_));
  INV        u0759(.A(men_men_n781_), .Y(men_men_n782_));
  AOI210     u0760(.A0(men_men_n32_), .A1(men_men_n35_), .B0(men_men_n429_), .Y(men_men_n783_));
  NA2        u0761(.A(men_men_n783_), .B(men_men_n782_), .Y(men_men_n784_));
  NO2        u0762(.A(men_men_n185_), .B(men_men_n120_), .Y(men_men_n785_));
  OAI210     u0763(.A0(men_men_n785_), .A1(men_men_n774_), .B0(i_2_), .Y(men_men_n786_));
  NO3        u0764(.A(men_men_n652_), .B(men_men_n37_), .C(men_men_n26_), .Y(men_men_n787_));
  AOI210     u0765(.A0(men_men_n165_), .A1(men_men_n84_), .B0(men_men_n787_), .Y(men_men_n788_));
  AOI210     u0766(.A0(men_men_n788_), .A1(men_men_n786_), .B0(men_men_n188_), .Y(men_men_n789_));
  AN2        u0767(.A(men_men_n121_), .B(i_13_), .Y(men_men_n790_));
  NA2        u0768(.A(men_men_n195_), .B(men_men_n198_), .Y(men_men_n791_));
  NA2        u0769(.A(men_men_n144_), .B(i_8_), .Y(men_men_n792_));
  AOI210     u0770(.A0(men_men_n792_), .A1(men_men_n791_), .B0(men_men_n383_), .Y(men_men_n793_));
  NA3        u0771(.A(men_men_n307_), .B(men_men_n119_), .C(men_men_n42_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n794_), .B(men_men_n46_), .Y(men_men_n795_));
  NO4        u0773(.A(men_men_n795_), .B(men_men_n793_), .C(men_men_n790_), .D(men_men_n789_), .Y(men_men_n796_));
  NO2        u0774(.A(men_men_n60_), .B(i_12_), .Y(men_men_n797_));
  INV        u0775(.A(men_men_n121_), .Y(men_men_n798_));
  NO2        u0776(.A(men_men_n798_), .B(i_8_), .Y(men_men_n799_));
  AOI220     u0777(.A0(men_men_n799_), .A1(men_men_n35_), .B0(men_men_n276_), .B1(men_men_n46_), .Y(men_men_n800_));
  NA4        u0778(.A(men_men_n800_), .B(men_men_n796_), .C(men_men_n784_), .D(men_men_n777_), .Y(men6));
  NA4        u0779(.A(men_men_n401_), .B(men_men_n1089_), .C(men_men_n67_), .D(men_men_n95_), .Y(men_men_n802_));
  INV        u0780(.A(men_men_n802_), .Y(men_men_n803_));
  NO2        u0781(.A(men_men_n217_), .B(men_men_n504_), .Y(men_men_n804_));
  NO2        u0782(.A(i_11_), .B(i_9_), .Y(men_men_n805_));
  NO2        u0783(.A(men_men_n803_), .B(men_men_n331_), .Y(men_men_n806_));
  OR2        u0784(.A(men_men_n806_), .B(i_12_), .Y(men_men_n807_));
  NA2        u0785(.A(men_men_n384_), .B(men_men_n339_), .Y(men_men_n808_));
  NA2        u0786(.A(men_men_n715_), .B(men_men_n67_), .Y(men_men_n809_));
  NA3        u0787(.A(men_men_n657_), .B(men_men_n809_), .C(men_men_n808_), .Y(men_men_n810_));
  INV        u0788(.A(men_men_n192_), .Y(men_men_n811_));
  AOI220     u0789(.A0(men_men_n811_), .A1(men_men_n805_), .B0(men_men_n810_), .B1(men_men_n69_), .Y(men_men_n812_));
  INV        u0790(.A(men_men_n330_), .Y(men_men_n813_));
  INV        u0791(.A(men_men_n125_), .Y(men_men_n814_));
  NO2        u0792(.A(men_men_n814_), .B(men_men_n813_), .Y(men_men_n815_));
  NO3        u0793(.A(men_men_n250_), .B(men_men_n126_), .C(i_9_), .Y(men_men_n816_));
  NA2        u0794(.A(men_men_n816_), .B(men_men_n797_), .Y(men_men_n817_));
  AOI210     u0795(.A0(men_men_n817_), .A1(men_men_n539_), .B0(men_men_n180_), .Y(men_men_n818_));
  NO2        u0796(.A(men_men_n31_), .B(i_11_), .Y(men_men_n819_));
  NA3        u0797(.A(men_men_n819_), .B(men_men_n494_), .C(men_men_n401_), .Y(men_men_n820_));
  NAi32      u0798(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n821_));
  AOI210     u0799(.A0(men_men_n750_), .A1(men_men_n82_), .B0(men_men_n821_), .Y(men_men_n822_));
  OAI210     u0800(.A0(men_men_n714_), .A1(men_men_n594_), .B0(men_men_n593_), .Y(men_men_n823_));
  NAi31      u0801(.An(men_men_n822_), .B(men_men_n823_), .C(men_men_n820_), .Y(men_men_n824_));
  OR3        u0802(.A(men_men_n824_), .B(men_men_n818_), .C(men_men_n815_), .Y(men_men_n825_));
  NO2        u0803(.A(men_men_n727_), .B(i_2_), .Y(men_men_n826_));
  NA2        u0804(.A(men_men_n48_), .B(men_men_n36_), .Y(men_men_n827_));
  NA2        u0805(.A(men_men_n1083_), .B(men_men_n826_), .Y(men_men_n828_));
  AO220      u0806(.A0(men_men_n367_), .A1(men_men_n357_), .B0(men_men_n409_), .B1(i_8_), .Y(men_men_n829_));
  NA2        u0807(.A(men_men_n829_), .B(men_men_n255_), .Y(men_men_n830_));
  OR2        u0808(.A(men_men_n653_), .B(men_men_n465_), .Y(men_men_n831_));
  NA3        u0809(.A(men_men_n831_), .B(men_men_n139_), .C(men_men_n66_), .Y(men_men_n832_));
  AO210      u0810(.A0(men_men_n510_), .A1(men_men_n776_), .B0(men_men_n35_), .Y(men_men_n833_));
  NA4        u0811(.A(men_men_n833_), .B(men_men_n832_), .C(men_men_n830_), .D(men_men_n828_), .Y(men_men_n834_));
  OAI210     u0812(.A0(i_6_), .A1(i_11_), .B0(men_men_n82_), .Y(men_men_n835_));
  AOI220     u0813(.A0(men_men_n835_), .A1(men_men_n593_), .B0(men_men_n804_), .B1(men_men_n744_), .Y(men_men_n836_));
  NA3        u0814(.A(men_men_n383_), .B(men_men_n236_), .C(men_men_n139_), .Y(men_men_n837_));
  NA3        u0815(.A(men_men_n837_), .B(men_men_n836_), .C(men_men_n636_), .Y(men_men_n838_));
  AO210      u0816(.A0(men_men_n541_), .A1(men_men_n46_), .B0(men_men_n83_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n839_), .B(men_men_n502_), .Y(men_men_n840_));
  INV        u0818(.A(men_men_n592_), .Y(men_men_n841_));
  NO2        u0819(.A(men_men_n644_), .B(men_men_n96_), .Y(men_men_n842_));
  OAI210     u0820(.A0(men_men_n842_), .A1(men_men_n106_), .B0(men_men_n421_), .Y(men_men_n843_));
  NA2        u0821(.A(men_men_n242_), .B(men_men_n46_), .Y(men_men_n844_));
  INV        u0822(.A(men_men_n620_), .Y(men_men_n845_));
  NA3        u0823(.A(men_men_n845_), .B(men_men_n330_), .C(i_7_), .Y(men_men_n846_));
  NA4        u0824(.A(men_men_n846_), .B(men_men_n843_), .C(men_men_n841_), .D(men_men_n840_), .Y(men_men_n847_));
  NO4        u0825(.A(men_men_n847_), .B(men_men_n838_), .C(men_men_n834_), .D(men_men_n825_), .Y(men_men_n848_));
  NA4        u0826(.A(men_men_n848_), .B(men_men_n812_), .C(men_men_n807_), .D(men_men_n391_), .Y(men3));
  NA2        u0827(.A(i_12_), .B(i_10_), .Y(men_men_n850_));
  NA2        u0828(.A(i_6_), .B(i_7_), .Y(men_men_n851_));
  NO2        u0829(.A(men_men_n851_), .B(i_0_), .Y(men_men_n852_));
  NO2        u0830(.A(i_11_), .B(men_men_n234_), .Y(men_men_n853_));
  OAI210     u0831(.A0(men_men_n852_), .A1(men_men_n291_), .B0(men_men_n853_), .Y(men_men_n854_));
  NO2        u0832(.A(men_men_n854_), .B(men_men_n188_), .Y(men_men_n855_));
  NO3        u0833(.A(men_men_n469_), .B(men_men_n86_), .C(men_men_n44_), .Y(men_men_n856_));
  OA210      u0834(.A0(men_men_n856_), .A1(men_men_n855_), .B0(men_men_n168_), .Y(men_men_n857_));
  NA3        u0835(.A(men_men_n837_), .B(men_men_n636_), .C(men_men_n382_), .Y(men_men_n858_));
  NA2        u0836(.A(men_men_n858_), .B(men_men_n39_), .Y(men_men_n859_));
  NOi21      u0837(.An(men_men_n90_), .B(men_men_n780_), .Y(men_men_n860_));
  NO3        u0838(.A(men_men_n662_), .B(men_men_n473_), .C(men_men_n125_), .Y(men_men_n861_));
  NA2        u0839(.A(men_men_n422_), .B(men_men_n45_), .Y(men_men_n862_));
  NO3        u0840(.A(men_men_n53_), .B(men_men_n861_), .C(men_men_n860_), .Y(men_men_n863_));
  AOI210     u0841(.A0(men_men_n863_), .A1(men_men_n859_), .B0(men_men_n48_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n180_), .B(men_men_n602_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n737_), .B(men_men_n704_), .Y(men_men_n866_));
  NA2        u0844(.A(men_men_n337_), .B(men_men_n453_), .Y(men_men_n867_));
  OAI220     u0845(.A0(men_men_n867_), .A1(men_men_n866_), .B0(men_men_n865_), .B1(men_men_n61_), .Y(men_men_n868_));
  NOi21      u0846(.An(i_5_), .B(i_9_), .Y(men_men_n869_));
  NA2        u0847(.A(men_men_n869_), .B(men_men_n461_), .Y(men_men_n870_));
  INV        u0848(.A(men_men_n719_), .Y(men_men_n871_));
  NO3        u0849(.A(men_men_n425_), .B(men_men_n268_), .C(men_men_n69_), .Y(men_men_n872_));
  NO2        u0850(.A(men_men_n169_), .B(men_men_n140_), .Y(men_men_n873_));
  AOI210     u0851(.A0(men_men_n873_), .A1(men_men_n242_), .B0(men_men_n872_), .Y(men_men_n874_));
  OAI220     u0852(.A0(men_men_n874_), .A1(men_men_n175_), .B0(men_men_n871_), .B1(men_men_n870_), .Y(men_men_n875_));
  NO4        u0853(.A(men_men_n875_), .B(men_men_n868_), .C(men_men_n864_), .D(men_men_n857_), .Y(men_men_n876_));
  NA2        u0854(.A(men_men_n180_), .B(men_men_n24_), .Y(men_men_n877_));
  NO2        u0855(.A(men_men_n703_), .B(men_men_n628_), .Y(men_men_n878_));
  NO2        u0856(.A(men_men_n878_), .B(men_men_n877_), .Y(men_men_n879_));
  NA2        u0857(.A(men_men_n314_), .B(men_men_n123_), .Y(men_men_n880_));
  NAi21      u0858(.An(men_men_n155_), .B(men_men_n453_), .Y(men_men_n881_));
  OAI220     u0859(.A0(men_men_n881_), .A1(men_men_n844_), .B0(men_men_n880_), .B1(men_men_n412_), .Y(men_men_n882_));
  NO2        u0860(.A(men_men_n882_), .B(men_men_n879_), .Y(men_men_n883_));
  NO2        u0861(.A(men_men_n401_), .B(men_men_n295_), .Y(men_men_n884_));
  NA2        u0862(.A(men_men_n884_), .B(men_men_n739_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n603_), .B(i_0_), .Y(men_men_n886_));
  NO3        u0864(.A(men_men_n886_), .B(men_men_n396_), .C(men_men_n84_), .Y(men_men_n887_));
  NO3        u0865(.A(men_men_n619_), .B(men_men_n211_), .C(men_men_n429_), .Y(men_men_n888_));
  AOI210     u0866(.A0(men_men_n888_), .A1(i_11_), .B0(men_men_n887_), .Y(men_men_n889_));
  INV        u0867(.A(men_men_n494_), .Y(men_men_n890_));
  AN2        u0868(.A(men_men_n90_), .B(men_men_n241_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n773_), .B(men_men_n331_), .Y(men_men_n892_));
  AOI210     u0870(.A0(men_men_n502_), .A1(men_men_n84_), .B0(men_men_n56_), .Y(men_men_n893_));
  OAI220     u0871(.A0(men_men_n893_), .A1(men_men_n892_), .B0(men_men_n690_), .B1(men_men_n564_), .Y(men_men_n894_));
  NO2        u0872(.A(men_men_n252_), .B(men_men_n146_), .Y(men_men_n895_));
  NA2        u0873(.A(i_0_), .B(i_10_), .Y(men_men_n896_));
  OAI210     u0874(.A0(men_men_n896_), .A1(men_men_n81_), .B0(men_men_n567_), .Y(men_men_n897_));
  NO4        u0875(.A(men_men_n109_), .B(men_men_n56_), .C(men_men_n700_), .D(i_5_), .Y(men_men_n898_));
  AO220      u0876(.A0(men_men_n898_), .A1(men_men_n897_), .B0(men_men_n895_), .B1(i_6_), .Y(men_men_n899_));
  AOI220     u0877(.A0(men_men_n337_), .A1(men_men_n92_), .B0(men_men_n180_), .B1(men_men_n79_), .Y(men_men_n900_));
  NA2        u0878(.A(men_men_n597_), .B(i_4_), .Y(men_men_n901_));
  NA2        u0879(.A(men_men_n183_), .B(men_men_n198_), .Y(men_men_n902_));
  OAI220     u0880(.A0(men_men_n902_), .A1(men_men_n892_), .B0(men_men_n901_), .B1(men_men_n900_), .Y(men_men_n903_));
  NO4        u0881(.A(men_men_n903_), .B(men_men_n899_), .C(men_men_n894_), .D(men_men_n891_), .Y(men_men_n904_));
  NA4        u0882(.A(men_men_n904_), .B(men_men_n889_), .C(men_men_n885_), .D(men_men_n883_), .Y(men_men_n905_));
  NO2        u0883(.A(men_men_n97_), .B(men_men_n36_), .Y(men_men_n906_));
  NA2        u0884(.A(i_11_), .B(i_9_), .Y(men_men_n907_));
  NO3        u0885(.A(i_12_), .B(men_men_n907_), .C(men_men_n635_), .Y(men_men_n908_));
  AN2        u0886(.A(men_men_n908_), .B(men_men_n906_), .Y(men_men_n909_));
  NO2        u0887(.A(men_men_n48_), .B(i_7_), .Y(men_men_n910_));
  NA2        u0888(.A(men_men_n406_), .B(men_men_n173_), .Y(men_men_n911_));
  NAi41      u0889(.An(men_men_n265_), .B(men_men_n911_), .C(men_men_n478_), .D(men_men_n153_), .Y(men_men_n912_));
  NO2        u0890(.A(men_men_n907_), .B(men_men_n69_), .Y(men_men_n913_));
  NO2        u0891(.A(men_men_n169_), .B(i_0_), .Y(men_men_n914_));
  INV        u0892(.A(men_men_n914_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n494_), .B(men_men_n228_), .Y(men_men_n916_));
  AOI210     u0894(.A0(men_men_n381_), .A1(men_men_n41_), .B0(men_men_n420_), .Y(men_men_n917_));
  OAI220     u0895(.A0(men_men_n917_), .A1(men_men_n870_), .B0(men_men_n916_), .B1(men_men_n915_), .Y(men_men_n918_));
  NO3        u0896(.A(men_men_n918_), .B(men_men_n912_), .C(men_men_n909_), .Y(men_men_n919_));
  AOI210     u0897(.A0(men_men_n464_), .A1(men_men_n35_), .B0(i_3_), .Y(men_men_n920_));
  NA2        u0898(.A(men_men_n165_), .B(men_men_n97_), .Y(men_men_n921_));
  NOi32      u0899(.An(men_men_n920_), .Bn(men_men_n183_), .C(men_men_n921_), .Y(men_men_n922_));
  AOI210     u0900(.A0(men_men_n637_), .A1(men_men_n331_), .B0(men_men_n241_), .Y(men_men_n923_));
  NO2        u0901(.A(men_men_n923_), .B(men_men_n862_), .Y(men_men_n924_));
  NO2        u0902(.A(men_men_n924_), .B(men_men_n922_), .Y(men_men_n925_));
  NOi21      u0903(.An(i_7_), .B(i_5_), .Y(men_men_n926_));
  NOi31      u0904(.An(men_men_n926_), .B(i_0_), .C(men_men_n755_), .Y(men_men_n927_));
  NA3        u0905(.A(men_men_n927_), .B(men_men_n395_), .C(i_6_), .Y(men_men_n928_));
  OA210      u0906(.A0(men_men_n921_), .A1(men_men_n539_), .B0(men_men_n928_), .Y(men_men_n929_));
  NO3        u0907(.A(men_men_n415_), .B(men_men_n370_), .C(men_men_n366_), .Y(men_men_n930_));
  NO2        u0908(.A(men_men_n262_), .B(men_men_n320_), .Y(men_men_n931_));
  NO2        u0909(.A(men_men_n755_), .B(men_men_n257_), .Y(men_men_n932_));
  AOI210     u0910(.A0(men_men_n932_), .A1(men_men_n931_), .B0(men_men_n930_), .Y(men_men_n933_));
  NA4        u0911(.A(men_men_n933_), .B(men_men_n929_), .C(men_men_n925_), .D(men_men_n919_), .Y(men_men_n934_));
  NO2        u0912(.A(men_men_n877_), .B(men_men_n237_), .Y(men_men_n935_));
  AN2        u0913(.A(men_men_n336_), .B(men_men_n331_), .Y(men_men_n936_));
  AN2        u0914(.A(men_men_n936_), .B(men_men_n873_), .Y(men_men_n937_));
  OAI210     u0915(.A0(men_men_n937_), .A1(men_men_n935_), .B0(i_10_), .Y(men_men_n938_));
  NO2        u0916(.A(men_men_n850_), .B(men_men_n319_), .Y(men_men_n939_));
  OA210      u0917(.A0(men_men_n494_), .A1(men_men_n220_), .B0(men_men_n493_), .Y(men_men_n940_));
  NA2        u0918(.A(men_men_n939_), .B(men_men_n913_), .Y(men_men_n941_));
  NA3        u0919(.A(men_men_n493_), .B(men_men_n422_), .C(men_men_n45_), .Y(men_men_n942_));
  OAI210     u0920(.A0(men_men_n881_), .A1(men_men_n890_), .B0(men_men_n942_), .Y(men_men_n943_));
  NO2        u0921(.A(men_men_n255_), .B(men_men_n46_), .Y(men_men_n944_));
  NA2        u0922(.A(men_men_n913_), .B(men_men_n307_), .Y(men_men_n945_));
  OAI210     u0923(.A0(men_men_n944_), .A1(men_men_n182_), .B0(men_men_n945_), .Y(men_men_n946_));
  AOI220     u0924(.A0(men_men_n946_), .A1(men_men_n494_), .B0(men_men_n943_), .B1(men_men_n69_), .Y(men_men_n947_));
  NA3        u0925(.A(men_men_n827_), .B(men_men_n393_), .C(i_6_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n88_), .B(men_men_n44_), .Y(men_men_n949_));
  NO2        u0927(.A(men_men_n71_), .B(men_men_n775_), .Y(men_men_n950_));
  AOI220     u0928(.A0(men_men_n950_), .A1(men_men_n949_), .B0(men_men_n168_), .B1(men_men_n628_), .Y(men_men_n951_));
  AOI210     u0929(.A0(men_men_n951_), .A1(men_men_n948_), .B0(men_men_n47_), .Y(men_men_n952_));
  NO3        u0930(.A(men_men_n619_), .B(men_men_n365_), .C(men_men_n24_), .Y(men_men_n953_));
  AOI210     u0931(.A0(men_men_n731_), .A1(men_men_n576_), .B0(men_men_n953_), .Y(men_men_n954_));
  NAi21      u0932(.An(i_9_), .B(i_5_), .Y(men_men_n955_));
  NO2        u0933(.A(men_men_n955_), .B(men_men_n415_), .Y(men_men_n956_));
  NO2        u0934(.A(men_men_n632_), .B(men_men_n99_), .Y(men_men_n957_));
  AOI220     u0935(.A0(men_men_n957_), .A1(i_0_), .B0(men_men_n956_), .B1(men_men_n653_), .Y(men_men_n958_));
  OAI220     u0936(.A0(men_men_n958_), .A1(men_men_n81_), .B0(men_men_n954_), .B1(men_men_n166_), .Y(men_men_n959_));
  NO3        u0937(.A(men_men_n959_), .B(men_men_n952_), .C(men_men_n544_), .Y(men_men_n960_));
  NA4        u0938(.A(men_men_n960_), .B(men_men_n947_), .C(men_men_n941_), .D(men_men_n938_), .Y(men_men_n961_));
  NO3        u0939(.A(men_men_n961_), .B(men_men_n934_), .C(men_men_n905_), .Y(men_men_n962_));
  NO2        u0940(.A(i_0_), .B(men_men_n755_), .Y(men_men_n963_));
  NA2        u0941(.A(men_men_n69_), .B(men_men_n44_), .Y(men_men_n964_));
  NO3        u0942(.A(men_men_n99_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n965_));
  AO220      u0943(.A0(men_men_n965_), .A1(men_men_n69_), .B0(men_men_n963_), .B1(men_men_n168_), .Y(men_men_n966_));
  NO2        u0944(.A(men_men_n717_), .B(men_men_n921_), .Y(men_men_n967_));
  AOI210     u0945(.A0(men_men_n966_), .A1(men_men_n354_), .B0(men_men_n967_), .Y(men_men_n968_));
  NA2        u0946(.A(men_men_n764_), .B(men_men_n138_), .Y(men_men_n969_));
  INV        u0947(.A(men_men_n969_), .Y(men_men_n970_));
  NA2        u0948(.A(men_men_n970_), .B(men_men_n704_), .Y(men_men_n971_));
  NO2        u0949(.A(men_men_n823_), .B(men_men_n415_), .Y(men_men_n972_));
  NA3        u0950(.A(men_men_n852_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n973_));
  AOI210     u0951(.A0(men_men_n973_), .A1(men_men_n516_), .B0(men_men_n1091_), .Y(men_men_n974_));
  NO2        u0952(.A(men_men_n974_), .B(men_men_n972_), .Y(men_men_n975_));
  NA3        u0953(.A(men_men_n975_), .B(men_men_n971_), .C(men_men_n968_), .Y(men_men_n976_));
  NA2        u0954(.A(men_men_n936_), .B(men_men_n383_), .Y(men_men_n977_));
  AOI210     u0955(.A0(men_men_n302_), .A1(men_men_n155_), .B0(men_men_n977_), .Y(men_men_n978_));
  NA3        u0956(.A(men_men_n39_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n979_));
  NA2        u0957(.A(men_men_n910_), .B(men_men_n505_), .Y(men_men_n980_));
  AOI210     u0958(.A0(men_men_n979_), .A1(men_men_n155_), .B0(men_men_n980_), .Y(men_men_n981_));
  NO2        u0959(.A(men_men_n981_), .B(men_men_n978_), .Y(men_men_n982_));
  NO3        u0960(.A(men_men_n896_), .B(men_men_n869_), .C(men_men_n185_), .Y(men_men_n983_));
  NA2        u0961(.A(men_men_n983_), .B(i_11_), .Y(men_men_n984_));
  INV        u0962(.A(men_men_n214_), .Y(men_men_n985_));
  OAI220     u0963(.A0(men_men_n557_), .A1(men_men_n1090_), .B0(men_men_n677_), .B1(men_men_n648_), .Y(men_men_n986_));
  NA3        u0964(.A(men_men_n986_), .B(men_men_n410_), .C(men_men_n985_), .Y(men_men_n987_));
  NA3        u0965(.A(men_men_n987_), .B(men_men_n984_), .C(men_men_n982_), .Y(men_men_n988_));
  NO2        u0966(.A(men_men_n240_), .B(men_men_n88_), .Y(men_men_n989_));
  NA2        u0967(.A(men_men_n989_), .B(men_men_n963_), .Y(men_men_n990_));
  AOI220     u0968(.A0(men_men_n926_), .A1(men_men_n505_), .B0(men_men_n852_), .B1(men_men_n156_), .Y(men_men_n991_));
  NA2        u0969(.A(men_men_n357_), .B(men_men_n170_), .Y(men_men_n992_));
  OA220      u0970(.A0(men_men_n992_), .A1(men_men_n991_), .B0(men_men_n990_), .B1(i_5_), .Y(men_men_n993_));
  AOI210     u0971(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n169_), .Y(men_men_n994_));
  NA2        u0972(.A(men_men_n994_), .B(men_men_n940_), .Y(men_men_n995_));
  NA3        u0973(.A(men_men_n645_), .B(men_men_n180_), .C(men_men_n79_), .Y(men_men_n996_));
  NA2        u0974(.A(men_men_n996_), .B(men_men_n574_), .Y(men_men_n997_));
  NO3        u0975(.A(men_men_n862_), .B(men_men_n52_), .C(men_men_n48_), .Y(men_men_n998_));
  NO3        u0976(.A(men_men_n1079_), .B(men_men_n998_), .C(men_men_n997_), .Y(men_men_n999_));
  NA3        u0977(.A(men_men_n401_), .B(men_men_n165_), .C(men_men_n164_), .Y(men_men_n1000_));
  NA3        u0978(.A(men_men_n910_), .B(men_men_n291_), .C(men_men_n227_), .Y(men_men_n1001_));
  NA2        u0979(.A(men_men_n1001_), .B(men_men_n1000_), .Y(men_men_n1002_));
  NA3        u0980(.A(men_men_n401_), .B(men_men_n338_), .C(men_men_n218_), .Y(men_men_n1003_));
  INV        u0981(.A(men_men_n1003_), .Y(men_men_n1004_));
  NOi31      u0982(.An(men_men_n400_), .B(men_men_n964_), .C(men_men_n237_), .Y(men_men_n1005_));
  NO3        u0983(.A(men_men_n907_), .B(men_men_n214_), .C(men_men_n185_), .Y(men_men_n1006_));
  NO4        u0984(.A(men_men_n1006_), .B(men_men_n1005_), .C(men_men_n1004_), .D(men_men_n1002_), .Y(men_men_n1007_));
  NA4        u0985(.A(men_men_n1007_), .B(men_men_n999_), .C(men_men_n995_), .D(men_men_n993_), .Y(men_men_n1008_));
  INV        u0986(.A(men_men_n647_), .Y(men_men_n1009_));
  NO3        u0987(.A(men_men_n1009_), .B(men_men_n588_), .C(men_men_n351_), .Y(men_men_n1010_));
  NA3        u0988(.A(men_men_n853_), .B(men_men_n104_), .C(men_men_n119_), .Y(men_men_n1011_));
  INV        u0989(.A(men_men_n1011_), .Y(men_men_n1012_));
  AOI210     u0990(.A0(men_men_n1012_), .A1(men_men_n1087_), .B0(men_men_n1010_), .Y(men_men_n1013_));
  NA3        u0991(.A(men_men_n307_), .B(i_5_), .C(men_men_n188_), .Y(men_men_n1014_));
  NAi31      u0992(.An(men_men_n239_), .B(men_men_n1014_), .C(men_men_n240_), .Y(men_men_n1015_));
  NO4        u0993(.A(men_men_n237_), .B(men_men_n205_), .C(i_0_), .D(i_12_), .Y(men_men_n1016_));
  AOI220     u0994(.A0(men_men_n1016_), .A1(men_men_n1015_), .B0(men_men_n803_), .B1(men_men_n170_), .Y(men_men_n1017_));
  AN2        u0995(.A(men_men_n896_), .B(men_men_n146_), .Y(men_men_n1018_));
  NO4        u0996(.A(men_men_n1018_), .B(i_12_), .C(men_men_n681_), .D(men_men_n125_), .Y(men_men_n1019_));
  NA2        u0997(.A(men_men_n1019_), .B(men_men_n214_), .Y(men_men_n1020_));
  NA3        u0998(.A(men_men_n92_), .B(men_men_n602_), .C(i_11_), .Y(men_men_n1021_));
  NO2        u0999(.A(men_men_n1021_), .B(men_men_n148_), .Y(men_men_n1022_));
  NA2        u1000(.A(men_men_n926_), .B(men_men_n491_), .Y(men_men_n1023_));
  OAI220     u1001(.A0(i_7_), .A1(men_men_n1014_), .B0(men_men_n1023_), .B1(men_men_n705_), .Y(men_men_n1024_));
  AOI210     u1002(.A0(men_men_n1024_), .A1(men_men_n914_), .B0(men_men_n1022_), .Y(men_men_n1025_));
  NA4        u1003(.A(men_men_n1025_), .B(men_men_n1020_), .C(men_men_n1017_), .D(men_men_n1013_), .Y(men_men_n1026_));
  NO4        u1004(.A(men_men_n1026_), .B(men_men_n1008_), .C(men_men_n988_), .D(men_men_n976_), .Y(men_men_n1027_));
  OAI210     u1005(.A0(men_men_n826_), .A1(men_men_n819_), .B0(men_men_n36_), .Y(men_men_n1028_));
  NA3        u1006(.A(men_men_n920_), .B(men_men_n378_), .C(i_5_), .Y(men_men_n1029_));
  NA3        u1007(.A(men_men_n1029_), .B(men_men_n1028_), .C(men_men_n643_), .Y(men_men_n1030_));
  NA2        u1008(.A(men_men_n1030_), .B(men_men_n202_), .Y(men_men_n1031_));
  AN2        u1009(.A(men_men_n727_), .B(men_men_n379_), .Y(men_men_n1032_));
  NA2        u1010(.A(men_men_n181_), .B(men_men_n183_), .Y(men_men_n1033_));
  AO210      u1011(.A0(men_men_n1032_), .A1(men_men_n32_), .B0(men_men_n1033_), .Y(men_men_n1034_));
  OAI210     u1012(.A0(men_men_n647_), .A1(men_men_n645_), .B0(men_men_n319_), .Y(men_men_n1035_));
  NAi31      u1013(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1036_));
  INV        u1014(.A(men_men_n1036_), .Y(men_men_n1037_));
  NO2        u1015(.A(men_men_n1037_), .B(men_men_n678_), .Y(men_men_n1038_));
  NA3        u1016(.A(men_men_n1038_), .B(men_men_n1035_), .C(men_men_n1034_), .Y(men_men_n1039_));
  NO2        u1017(.A(men_men_n481_), .B(men_men_n268_), .Y(men_men_n1040_));
  NO4        u1018(.A(men_men_n230_), .B(men_men_n137_), .C(men_men_n708_), .D(men_men_n36_), .Y(men_men_n1041_));
  NO3        u1019(.A(men_men_n1041_), .B(men_men_n1040_), .C(men_men_n888_), .Y(men_men_n1042_));
  OAI210     u1020(.A0(men_men_n1021_), .A1(men_men_n140_), .B0(men_men_n1042_), .Y(men_men_n1043_));
  AOI210     u1021(.A0(men_men_n1039_), .A1(men_men_n48_), .B0(men_men_n1043_), .Y(men_men_n1044_));
  AOI210     u1022(.A0(men_men_n1044_), .A1(men_men_n1031_), .B0(men_men_n69_), .Y(men_men_n1045_));
  NO2        u1023(.A(men_men_n595_), .B(men_men_n390_), .Y(men_men_n1046_));
  NO2        u1024(.A(men_men_n1046_), .B(men_men_n778_), .Y(men_men_n1047_));
  OAI210     u1025(.A0(men_men_n75_), .A1(men_men_n52_), .B0(men_men_n102_), .Y(men_men_n1048_));
  NA2        u1026(.A(men_men_n1048_), .B(men_men_n72_), .Y(men_men_n1049_));
  AOI210     u1027(.A0(men_men_n994_), .A1(men_men_n910_), .B0(men_men_n927_), .Y(men_men_n1050_));
  AOI210     u1028(.A0(men_men_n1050_), .A1(men_men_n1049_), .B0(men_men_n708_), .Y(men_men_n1051_));
  NA2        u1029(.A(men_men_n262_), .B(men_men_n55_), .Y(men_men_n1052_));
  AOI220     u1030(.A0(men_men_n1052_), .A1(men_men_n72_), .B0(men_men_n352_), .B1(men_men_n254_), .Y(men_men_n1053_));
  NO2        u1031(.A(men_men_n1053_), .B(men_men_n234_), .Y(men_men_n1054_));
  NA3        u1032(.A(men_men_n90_), .B(men_men_n309_), .C(men_men_n30_), .Y(men_men_n1055_));
  INV        u1033(.A(men_men_n1055_), .Y(men_men_n1056_));
  NO3        u1034(.A(men_men_n1056_), .B(men_men_n1054_), .C(men_men_n1051_), .Y(men_men_n1057_));
  OAI210     u1035(.A0(men_men_n270_), .A1(men_men_n151_), .B0(men_men_n84_), .Y(men_men_n1058_));
  NA3        u1036(.A(men_men_n779_), .B(men_men_n291_), .C(men_men_n75_), .Y(men_men_n1059_));
  AOI210     u1037(.A0(men_men_n1059_), .A1(men_men_n1058_), .B0(i_11_), .Y(men_men_n1060_));
  NA2        u1038(.A(men_men_n638_), .B(men_men_n211_), .Y(men_men_n1061_));
  OAI210     u1039(.A0(men_men_n1061_), .A1(men_men_n920_), .B0(men_men_n202_), .Y(men_men_n1062_));
  NA2        u1040(.A(men_men_n157_), .B(i_5_), .Y(men_men_n1063_));
  AOI210     u1041(.A0(men_men_n1062_), .A1(men_men_n791_), .B0(men_men_n1063_), .Y(men_men_n1064_));
  NO3        u1042(.A(men_men_n57_), .B(men_men_n56_), .C(i_4_), .Y(men_men_n1065_));
  OAI210     u1043(.A0(men_men_n931_), .A1(men_men_n309_), .B0(men_men_n1065_), .Y(men_men_n1066_));
  NO2        u1044(.A(men_men_n1066_), .B(men_men_n755_), .Y(men_men_n1067_));
  NO4        u1045(.A(men_men_n955_), .B(men_men_n496_), .C(men_men_n251_), .D(men_men_n250_), .Y(men_men_n1068_));
  NO2        u1046(.A(men_men_n1068_), .B(men_men_n592_), .Y(men_men_n1069_));
  NO2        u1047(.A(men_men_n822_), .B(men_men_n371_), .Y(men_men_n1070_));
  AOI210     u1048(.A0(men_men_n1070_), .A1(men_men_n1069_), .B0(men_men_n40_), .Y(men_men_n1071_));
  NO4        u1049(.A(men_men_n1071_), .B(men_men_n1067_), .C(men_men_n1064_), .D(men_men_n1060_), .Y(men_men_n1072_));
  OAI210     u1050(.A0(men_men_n1057_), .A1(i_4_), .B0(men_men_n1072_), .Y(men_men_n1073_));
  NO3        u1051(.A(men_men_n1073_), .B(men_men_n1047_), .C(men_men_n1045_), .Y(men_men_n1074_));
  NA4        u1052(.A(men_men_n1074_), .B(men_men_n1027_), .C(men_men_n962_), .D(men_men_n876_), .Y(men4));
  INV        u1053(.A(i_5_), .Y(men_men_n1078_));
  INV        u1054(.A(men_men_n503_), .Y(men_men_n1079_));
  INV        u1055(.A(i_3_), .Y(men_men_n1080_));
  INV        u1056(.A(i_6_), .Y(men_men_n1081_));
  INV        u1057(.A(men_men_n136_), .Y(men_men_n1082_));
  INV        u1058(.A(men_men_n827_), .Y(men_men_n1083_));
  INV        u1059(.A(men_men_n193_), .Y(men_men_n1084_));
  INV        u1060(.A(men_men_n374_), .Y(men_men_n1085_));
  INV        u1061(.A(i_4_), .Y(men_men_n1086_));
  INV        u1062(.A(i_5_), .Y(men_men_n1087_));
  INV        u1063(.A(i_6_), .Y(men_men_n1088_));
  INV        u1064(.A(i_3_), .Y(men_men_n1089_));
  INV        u1065(.A(i_6_), .Y(men_men_n1090_));
  INV        u1066(.A(i_9_), .Y(men_men_n1091_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule