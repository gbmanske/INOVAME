// Benchmark "top" written by ABC on Thu Jun 20 14:59:14 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n141_, new_new_n142_, new_new_n143_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n700_, new_new_n701_, new_new_n702_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n973_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g040(.A(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g063(.A(i_6_), .Y(new_new_n86_));
  OR4        g064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n88_), .B(new_new_n89_), .Y(new_new_n90_));
  OAI210     g068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g073(.A(new_new_n95_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n98_));
  AN3        g076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g080(.A0(new_new_n102_), .A1(new_new_n62_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g081(.A(i_7_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n46_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(new_new_n86_), .Y(new_new_n107_));
  NA2        g085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  AN2        g089(.A(i_2_), .B(i_10_), .Y(new_new_n112_));
  NO2        g090(.A(new_new_n112_), .B(i_7_), .Y(new_new_n113_));
  OR2        g091(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n114_));
  NO2        g092(.A(i_8_), .B(new_new_n104_), .Y(new_new_n115_));
  NO3        g093(.A(new_new_n115_), .B(new_new_n114_), .C(new_new_n113_), .Y(new_new_n116_));
  NA2        g094(.A(i_12_), .B(i_7_), .Y(new_new_n117_));
  NO2        g095(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(i_0_), .Y(new_new_n119_));
  NA2        g097(.A(i_11_), .B(i_12_), .Y(new_new_n120_));
  OAI210     g098(.A0(new_new_n119_), .A1(new_new_n117_), .B0(new_new_n120_), .Y(new_new_n121_));
  NO2        g099(.A(new_new_n121_), .B(new_new_n116_), .Y(new_new_n122_));
  NA3        g100(.A(new_new_n122_), .B(new_new_n110_), .C(new_new_n103_), .Y(new_new_n123_));
  NOi21      g101(.An(i_1_), .B(i_5_), .Y(new_new_n124_));
  NA2        g102(.A(new_new_n124_), .B(i_11_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n126_));
  NA2        g104(.A(i_7_), .B(new_new_n25_), .Y(new_new_n127_));
  NA2        g105(.A(new_new_n127_), .B(new_new_n126_), .Y(new_new_n128_));
  NO2        g106(.A(new_new_n128_), .B(new_new_n46_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n130_));
  NAi21      g108(.An(i_3_), .B(i_8_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(new_new_n62_), .Y(new_new_n132_));
  NOi31      g110(.An(new_new_n132_), .B(new_new_n130_), .C(new_new_n129_), .Y(new_new_n133_));
  NO2        g111(.A(i_1_), .B(new_new_n86_), .Y(new_new_n134_));
  NO2        g112(.A(i_6_), .B(i_5_), .Y(new_new_n135_));
  NA2        g113(.A(new_new_n135_), .B(i_3_), .Y(new_new_n136_));
  AO210      g114(.A0(new_new_n136_), .A1(new_new_n47_), .B0(new_new_n134_), .Y(new_new_n137_));
  OAI220     g115(.A0(new_new_n137_), .A1(new_new_n111_), .B0(new_new_n133_), .B1(new_new_n125_), .Y(new_new_n138_));
  NO3        g116(.A(new_new_n138_), .B(new_new_n123_), .C(new_new_n98_), .Y(new_new_n139_));
  NA3        g117(.A(new_new_n139_), .B(new_new_n79_), .C(new_new_n56_), .Y(ori2));
  NO2        g118(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n141_));
  INV        g119(.A(i_6_), .Y(new_new_n142_));
  NA2        g120(.A(new_new_n142_), .B(new_new_n141_), .Y(new_new_n143_));
  NA4        g121(.A(new_new_n143_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(ori0));
  AN2        g122(.A(i_8_), .B(i_7_), .Y(new_new_n145_));
  NA2        g123(.A(new_new_n145_), .B(i_6_), .Y(new_new_n146_));
  NO2        g124(.A(i_12_), .B(i_13_), .Y(new_new_n147_));
  NAi21      g125(.An(i_5_), .B(i_11_), .Y(new_new_n148_));
  NOi21      g126(.An(new_new_n147_), .B(new_new_n148_), .Y(new_new_n149_));
  NO2        g127(.A(i_0_), .B(i_1_), .Y(new_new_n150_));
  NA2        g128(.A(i_2_), .B(i_3_), .Y(new_new_n151_));
  NO2        g129(.A(new_new_n151_), .B(i_4_), .Y(new_new_n152_));
  NA3        g130(.A(new_new_n152_), .B(new_new_n150_), .C(new_new_n149_), .Y(new_new_n153_));
  AN2        g131(.A(new_new_n147_), .B(new_new_n83_), .Y(new_new_n154_));
  NA2        g132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g133(.A(new_new_n73_), .B(new_new_n46_), .Y(new_new_n156_));
  NA2        g134(.A(new_new_n156_), .B(new_new_n36_), .Y(new_new_n157_));
  OR2        g135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NO3        g136(.A(new_new_n158_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n159_));
  NAi32      g137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n160_));
  NAi21      g138(.An(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  NOi21      g139(.An(i_4_), .B(i_10_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n40_), .Y(new_new_n163_));
  NO2        g141(.A(i_3_), .B(i_5_), .Y(new_new_n164_));
  NO3        g142(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  OAI210     g144(.A0(new_new_n166_), .A1(new_new_n163_), .B0(new_new_n161_), .Y(new_new_n167_));
  INV        g145(.A(new_new_n167_), .Y(new_new_n168_));
  NO2        g146(.A(new_new_n168_), .B(new_new_n146_), .Y(new_new_n169_));
  NA2        g147(.A(i_3_), .B(new_new_n48_), .Y(new_new_n170_));
  NOi21      g148(.An(i_4_), .B(i_9_), .Y(new_new_n171_));
  NOi21      g149(.An(i_11_), .B(i_13_), .Y(new_new_n172_));
  NA2        g150(.A(new_new_n172_), .B(new_new_n171_), .Y(new_new_n173_));
  NO2        g151(.A(i_4_), .B(i_5_), .Y(new_new_n174_));
  NAi21      g152(.An(i_12_), .B(i_11_), .Y(new_new_n175_));
  NO2        g153(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n176_));
  NA2        g154(.A(new_new_n176_), .B(new_new_n46_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n36_), .B(i_5_), .Y(new_new_n178_));
  NAi31      g156(.An(new_new_n178_), .B(new_new_n154_), .C(i_11_), .Y(new_new_n179_));
  NA2        g157(.A(i_3_), .B(i_5_), .Y(new_new_n180_));
  OR2        g158(.A(new_new_n180_), .B(new_new_n173_), .Y(new_new_n181_));
  AOI210     g159(.A0(new_new_n181_), .A1(new_new_n179_), .B0(new_new_n177_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n73_), .B(i_5_), .Y(new_new_n183_));
  NO2        g161(.A(i_13_), .B(i_10_), .Y(new_new_n184_));
  NA3        g162(.A(new_new_n184_), .B(new_new_n183_), .C(new_new_n44_), .Y(new_new_n185_));
  NO2        g163(.A(i_2_), .B(i_1_), .Y(new_new_n186_));
  NAi21      g164(.An(i_4_), .B(i_12_), .Y(new_new_n187_));
  INV        g165(.A(new_new_n182_), .Y(new_new_n188_));
  INV        g166(.A(i_8_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n189_), .B(i_7_), .Y(new_new_n190_));
  NA2        g168(.A(new_new_n190_), .B(i_6_), .Y(new_new_n191_));
  NO3        g169(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n192_));
  NO3        g170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n193_));
  NO3        g171(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n194_));
  NO2        g172(.A(i_3_), .B(i_8_), .Y(new_new_n195_));
  NO3        g173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n40_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n106_), .B(new_new_n58_), .Y(new_new_n198_));
  INV        g176(.A(new_new_n198_), .Y(new_new_n199_));
  NO2        g177(.A(i_13_), .B(i_9_), .Y(new_new_n200_));
  NAi21      g178(.An(i_12_), .B(i_3_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n44_), .B(i_5_), .Y(new_new_n202_));
  NO3        g180(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n199_), .B(new_new_n197_), .Y(new_new_n204_));
  NA2        g182(.A(new_new_n204_), .B(i_7_), .Y(new_new_n205_));
  OAI220     g183(.A0(new_new_n205_), .A1(i_4_), .B0(new_new_n191_), .B1(new_new_n188_), .Y(new_new_n206_));
  NAi21      g184(.An(i_12_), .B(i_7_), .Y(new_new_n207_));
  NA3        g185(.A(i_13_), .B(new_new_n189_), .C(i_10_), .Y(new_new_n208_));
  NA2        g186(.A(i_0_), .B(i_5_), .Y(new_new_n209_));
  NAi31      g187(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n36_), .B(i_13_), .Y(new_new_n211_));
  NO2        g189(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n212_));
  NO2        g190(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n213_));
  NA3        g191(.A(new_new_n213_), .B(new_new_n212_), .C(new_new_n211_), .Y(new_new_n214_));
  INV        g192(.A(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(i_12_), .B(new_new_n215_), .Y(new_new_n216_));
  NA3        g194(.A(new_new_n216_), .B(new_new_n193_), .C(new_new_n192_), .Y(new_new_n217_));
  OAI210     g195(.A0(new_new_n214_), .A1(new_new_n210_), .B0(new_new_n217_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n218_), .B(new_new_n145_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n37_), .Y(new_new_n220_));
  OR2        g198(.A(i_8_), .B(i_7_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n53_), .B(i_1_), .Y(new_new_n222_));
  INV        g200(.A(i_12_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n44_), .B(new_new_n223_), .Y(new_new_n224_));
  NO3        g202(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n225_));
  NA2        g203(.A(i_2_), .B(i_1_), .Y(new_new_n226_));
  NO3        g204(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n227_));
  NAi21      g205(.An(i_4_), .B(i_3_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n228_), .B(new_new_n75_), .Y(new_new_n229_));
  NO2        g207(.A(i_0_), .B(i_6_), .Y(new_new_n230_));
  NOi41      g208(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n226_), .B(new_new_n180_), .Y(new_new_n232_));
  NO2        g210(.A(i_11_), .B(new_new_n215_), .Y(new_new_n233_));
  NOi21      g211(.An(i_1_), .B(i_6_), .Y(new_new_n234_));
  NAi21      g212(.An(i_3_), .B(i_7_), .Y(new_new_n235_));
  NA2        g213(.A(new_new_n223_), .B(i_9_), .Y(new_new_n236_));
  OR4        g214(.A(new_new_n236_), .B(new_new_n235_), .C(new_new_n234_), .D(new_new_n183_), .Y(new_new_n237_));
  NA2        g215(.A(new_new_n73_), .B(i_5_), .Y(new_new_n238_));
  NA2        g216(.A(i_3_), .B(i_9_), .Y(new_new_n239_));
  NAi21      g217(.An(i_7_), .B(i_10_), .Y(new_new_n240_));
  NO2        g218(.A(new_new_n240_), .B(new_new_n239_), .Y(new_new_n241_));
  NA3        g219(.A(new_new_n241_), .B(new_new_n238_), .C(new_new_n64_), .Y(new_new_n242_));
  NA2        g220(.A(new_new_n242_), .B(new_new_n237_), .Y(new_new_n243_));
  INV        g221(.A(new_new_n146_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n223_), .B(i_13_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n245_), .B(new_new_n75_), .Y(new_new_n246_));
  AOI220     g224(.A0(new_new_n246_), .A1(new_new_n244_), .B0(new_new_n243_), .B1(new_new_n233_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n221_), .B(new_new_n37_), .Y(new_new_n248_));
  NA2        g226(.A(i_12_), .B(i_6_), .Y(new_new_n249_));
  OR2        g227(.A(i_13_), .B(i_9_), .Y(new_new_n250_));
  NO3        g228(.A(new_new_n250_), .B(new_new_n249_), .C(new_new_n48_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n228_), .B(i_2_), .Y(new_new_n252_));
  NA3        g230(.A(new_new_n252_), .B(new_new_n251_), .C(new_new_n44_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n233_), .B(i_9_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n238_), .B(new_new_n64_), .Y(new_new_n255_));
  OAI210     g233(.A0(new_new_n255_), .A1(new_new_n254_), .B0(new_new_n253_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n156_), .B(new_new_n63_), .Y(new_new_n257_));
  NO3        g235(.A(i_11_), .B(new_new_n215_), .C(new_new_n25_), .Y(new_new_n258_));
  NO2        g236(.A(new_new_n235_), .B(i_8_), .Y(new_new_n259_));
  NO2        g237(.A(i_6_), .B(new_new_n48_), .Y(new_new_n260_));
  NA3        g238(.A(new_new_n260_), .B(new_new_n259_), .C(new_new_n258_), .Y(new_new_n261_));
  NO3        g239(.A(new_new_n26_), .B(new_new_n86_), .C(i_5_), .Y(new_new_n262_));
  NA3        g240(.A(new_new_n262_), .B(new_new_n248_), .C(new_new_n216_), .Y(new_new_n263_));
  AOI210     g241(.A0(new_new_n263_), .A1(new_new_n261_), .B0(new_new_n257_), .Y(new_new_n264_));
  AOI210     g242(.A0(new_new_n256_), .A1(new_new_n248_), .B0(new_new_n264_), .Y(new_new_n265_));
  NA3        g243(.A(new_new_n265_), .B(new_new_n247_), .C(new_new_n219_), .Y(new_new_n266_));
  NO3        g244(.A(i_12_), .B(new_new_n215_), .C(new_new_n37_), .Y(new_new_n267_));
  INV        g245(.A(new_new_n267_), .Y(new_new_n268_));
  NA2        g246(.A(i_8_), .B(new_new_n104_), .Y(new_new_n269_));
  NOi21      g247(.An(new_new_n164_), .B(new_new_n86_), .Y(new_new_n270_));
  NO3        g248(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n271_));
  AOI220     g249(.A0(new_new_n271_), .A1(new_new_n192_), .B0(new_new_n270_), .B1(new_new_n222_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n272_), .B(new_new_n269_), .Y(new_new_n273_));
  NO3        g251(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n226_), .B(i_0_), .Y(new_new_n275_));
  AOI220     g253(.A0(new_new_n275_), .A1(new_new_n190_), .B0(new_new_n274_), .B1(new_new_n145_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n260_), .B(new_new_n26_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n277_), .B(new_new_n276_), .Y(new_new_n278_));
  NA2        g256(.A(i_0_), .B(i_1_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(i_2_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n59_), .B(i_6_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n166_), .B(new_new_n146_), .Y(new_new_n282_));
  NO3        g260(.A(new_new_n282_), .B(new_new_n278_), .C(new_new_n273_), .Y(new_new_n283_));
  NO2        g261(.A(i_2_), .B(new_new_n104_), .Y(new_new_n284_));
  NA2        g262(.A(i_1_), .B(new_new_n36_), .Y(new_new_n285_));
  AN2        g263(.A(i_3_), .B(i_10_), .Y(new_new_n286_));
  NO2        g264(.A(i_5_), .B(new_new_n37_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n283_), .B(new_new_n268_), .Y(new_new_n289_));
  NO4        g267(.A(new_new_n289_), .B(new_new_n266_), .C(new_new_n206_), .D(new_new_n169_), .Y(new_new_n290_));
  NO3        g268(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n59_), .B(new_new_n86_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n275_), .B(new_new_n292_), .Y(new_new_n293_));
  NO3        g271(.A(i_6_), .B(new_new_n189_), .C(i_7_), .Y(new_new_n294_));
  NA2        g272(.A(new_new_n294_), .B(new_new_n193_), .Y(new_new_n295_));
  AOI210     g273(.A0(new_new_n295_), .A1(new_new_n293_), .B0(new_new_n170_), .Y(new_new_n296_));
  NO2        g274(.A(i_2_), .B(i_3_), .Y(new_new_n297_));
  OR2        g275(.A(i_0_), .B(i_5_), .Y(new_new_n298_));
  NA3        g276(.A(new_new_n275_), .B(new_new_n270_), .C(new_new_n115_), .Y(new_new_n299_));
  NAi21      g277(.An(i_8_), .B(i_7_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n158_), .B(new_new_n46_), .Y(new_new_n301_));
  INV        g279(.A(new_new_n299_), .Y(new_new_n302_));
  OAI210     g280(.A0(new_new_n302_), .A1(new_new_n296_), .B0(i_4_), .Y(new_new_n303_));
  NO2        g281(.A(i_12_), .B(i_10_), .Y(new_new_n304_));
  NOi21      g282(.An(i_5_), .B(i_0_), .Y(new_new_n305_));
  AOI210     g283(.A0(i_2_), .A1(new_new_n48_), .B0(new_new_n104_), .Y(new_new_n306_));
  NO4        g284(.A(new_new_n306_), .B(new_new_n285_), .C(new_new_n305_), .D(new_new_n131_), .Y(new_new_n307_));
  NA4        g285(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n308_));
  NA2        g286(.A(new_new_n307_), .B(new_new_n304_), .Y(new_new_n309_));
  NO2        g287(.A(i_6_), .B(i_8_), .Y(new_new_n310_));
  NOi21      g288(.An(i_0_), .B(i_2_), .Y(new_new_n311_));
  AN2        g289(.A(new_new_n311_), .B(new_new_n310_), .Y(new_new_n312_));
  NO2        g290(.A(i_1_), .B(i_7_), .Y(new_new_n313_));
  NA2        g291(.A(new_new_n309_), .B(new_new_n303_), .Y(new_new_n314_));
  NOi21      g292(.An(new_new_n155_), .B(new_new_n107_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n315_), .B(new_new_n127_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(i_3_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n189_), .B(i_9_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n318_), .B(new_new_n198_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n319_), .B(new_new_n46_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n320_), .B(new_new_n278_), .Y(new_new_n321_));
  AOI210     g299(.A0(new_new_n321_), .A1(new_new_n317_), .B0(new_new_n163_), .Y(new_new_n322_));
  AOI210     g300(.A0(new_new_n314_), .A1(new_new_n291_), .B0(new_new_n322_), .Y(new_new_n323_));
  NOi32      g301(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n324_));
  INV        g302(.A(new_new_n324_), .Y(new_new_n325_));
  NAi21      g303(.An(i_1_), .B(i_5_), .Y(new_new_n326_));
  NAi41      g304(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n327_));
  OAI220     g305(.A0(new_new_n327_), .A1(new_new_n326_), .B0(new_new_n210_), .B1(new_new_n160_), .Y(new_new_n328_));
  AOI210     g306(.A0(new_new_n327_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n329_));
  NOi32      g307(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n330_));
  NAi21      g308(.An(i_6_), .B(i_1_), .Y(new_new_n331_));
  NA3        g309(.A(new_new_n331_), .B(new_new_n330_), .C(new_new_n46_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n332_), .B(i_0_), .Y(new_new_n333_));
  OR3        g311(.A(new_new_n333_), .B(new_new_n329_), .C(new_new_n328_), .Y(new_new_n334_));
  NO2        g312(.A(i_1_), .B(new_new_n104_), .Y(new_new_n335_));
  NAi21      g313(.An(i_3_), .B(i_4_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n336_), .B(i_9_), .Y(new_new_n337_));
  AN2        g315(.A(i_6_), .B(i_7_), .Y(new_new_n338_));
  OAI210     g316(.A0(new_new_n338_), .A1(new_new_n335_), .B0(new_new_n337_), .Y(new_new_n339_));
  NA2        g317(.A(i_2_), .B(i_7_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n336_), .B(i_10_), .Y(new_new_n341_));
  NA3        g319(.A(new_new_n341_), .B(new_new_n340_), .C(new_new_n230_), .Y(new_new_n342_));
  AOI210     g320(.A0(new_new_n342_), .A1(new_new_n339_), .B0(new_new_n183_), .Y(new_new_n343_));
  AOI210     g321(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n344_));
  OAI210     g322(.A0(new_new_n344_), .A1(new_new_n186_), .B0(new_new_n341_), .Y(new_new_n345_));
  AOI220     g323(.A0(new_new_n341_), .A1(new_new_n313_), .B0(new_new_n225_), .B1(new_new_n186_), .Y(new_new_n346_));
  AOI210     g324(.A0(new_new_n346_), .A1(new_new_n345_), .B0(i_5_), .Y(new_new_n347_));
  NO3        g325(.A(new_new_n347_), .B(new_new_n343_), .C(new_new_n334_), .Y(new_new_n348_));
  NO2        g326(.A(new_new_n348_), .B(new_new_n325_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n350_));
  AN2        g328(.A(i_12_), .B(i_5_), .Y(new_new_n351_));
  NO2        g329(.A(i_4_), .B(new_new_n26_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n352_), .B(new_new_n351_), .Y(new_new_n353_));
  NO2        g331(.A(i_11_), .B(i_6_), .Y(new_new_n354_));
  NA3        g332(.A(new_new_n354_), .B(new_new_n301_), .C(new_new_n215_), .Y(new_new_n355_));
  NO2        g333(.A(new_new_n355_), .B(new_new_n353_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n228_), .B(i_5_), .Y(new_new_n357_));
  NO2        g335(.A(i_5_), .B(i_10_), .Y(new_new_n358_));
  AOI220     g336(.A0(new_new_n358_), .A1(new_new_n252_), .B0(new_new_n357_), .B1(new_new_n193_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n147_), .B(new_new_n45_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n361_));
  OAI210     g339(.A0(new_new_n361_), .A1(new_new_n356_), .B0(new_new_n350_), .Y(new_new_n362_));
  NO2        g340(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n153_), .B(new_new_n86_), .Y(new_new_n364_));
  OAI210     g342(.A0(new_new_n364_), .A1(new_new_n356_), .B0(new_new_n363_), .Y(new_new_n365_));
  NO3        g343(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n366_));
  NO2        g344(.A(i_11_), .B(i_12_), .Y(new_new_n367_));
  NA2        g345(.A(new_new_n358_), .B(new_new_n223_), .Y(new_new_n368_));
  NAi21      g346(.An(i_13_), .B(i_0_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n365_), .B(new_new_n362_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n44_), .B(new_new_n215_), .Y(new_new_n371_));
  NO3        g349(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n372_));
  NO2        g350(.A(i_0_), .B(i_11_), .Y(new_new_n373_));
  AN2        g351(.A(i_1_), .B(i_6_), .Y(new_new_n374_));
  NOi21      g352(.An(i_2_), .B(i_12_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n145_), .B(i_9_), .Y(new_new_n376_));
  NO2        g354(.A(new_new_n376_), .B(i_4_), .Y(new_new_n377_));
  NAi21      g355(.An(i_9_), .B(i_4_), .Y(new_new_n378_));
  OR2        g356(.A(i_13_), .B(i_10_), .Y(new_new_n379_));
  NO3        g357(.A(new_new_n379_), .B(new_new_n120_), .C(new_new_n378_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n173_), .B(new_new_n126_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n267_), .B(new_new_n382_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n315_), .Y(new_new_n384_));
  INV        g362(.A(new_new_n384_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n385_), .B(new_new_n26_), .Y(new_new_n386_));
  INV        g364(.A(new_new_n299_), .Y(new_new_n387_));
  NO2        g365(.A(new_new_n180_), .B(new_new_n86_), .Y(new_new_n388_));
  AOI220     g366(.A0(new_new_n388_), .A1(new_new_n280_), .B0(new_new_n262_), .B1(new_new_n203_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(new_new_n269_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n387_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n192_), .B(new_new_n99_), .Y(new_new_n392_));
  NA3        g370(.A(new_new_n301_), .B(new_new_n164_), .C(new_new_n86_), .Y(new_new_n393_));
  AOI210     g371(.A0(new_new_n393_), .A1(new_new_n392_), .B0(new_new_n300_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n189_), .B(i_10_), .Y(new_new_n395_));
  NA3        g373(.A(new_new_n238_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n281_), .B(new_new_n222_), .Y(new_new_n397_));
  OAI220     g375(.A0(new_new_n397_), .A1(new_new_n180_), .B0(new_new_n396_), .B1(new_new_n395_), .Y(new_new_n398_));
  NO2        g376(.A(i_3_), .B(new_new_n48_), .Y(new_new_n399_));
  NA3        g377(.A(new_new_n313_), .B(new_new_n312_), .C(new_new_n399_), .Y(new_new_n400_));
  INV        g378(.A(new_new_n400_), .Y(new_new_n401_));
  NO3        g379(.A(new_new_n401_), .B(new_new_n398_), .C(new_new_n394_), .Y(new_new_n402_));
  AOI210     g380(.A0(new_new_n402_), .A1(new_new_n391_), .B0(new_new_n254_), .Y(new_new_n403_));
  NO4        g381(.A(new_new_n403_), .B(new_new_n386_), .C(new_new_n370_), .D(new_new_n349_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n63_), .B(i_4_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n73_), .B(i_13_), .Y(new_new_n406_));
  NA3        g384(.A(new_new_n406_), .B(new_new_n405_), .C(i_2_), .Y(new_new_n407_));
  NO2        g385(.A(i_10_), .B(i_9_), .Y(new_new_n408_));
  NAi21      g386(.An(i_12_), .B(i_8_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n409_), .B(i_3_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n410_), .B(new_new_n408_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n46_), .B(i_4_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n412_), .B(new_new_n107_), .Y(new_new_n413_));
  OAI220     g391(.A0(new_new_n413_), .A1(new_new_n197_), .B0(new_new_n411_), .B1(new_new_n407_), .Y(new_new_n414_));
  NA2        g392(.A(new_new_n288_), .B(i_0_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n249_), .B(new_new_n100_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n417_), .B(new_new_n416_), .Y(new_new_n418_));
  NA2        g396(.A(i_8_), .B(i_9_), .Y(new_new_n419_));
  AOI210     g397(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n420_));
  OR2        g398(.A(new_new_n420_), .B(new_new_n419_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n267_), .B(new_new_n198_), .Y(new_new_n422_));
  OAI220     g400(.A0(new_new_n422_), .A1(new_new_n421_), .B0(new_new_n418_), .B1(new_new_n415_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n233_), .B(new_new_n287_), .Y(new_new_n424_));
  NO3        g402(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n425_));
  INV        g403(.A(new_new_n425_), .Y(new_new_n426_));
  NA3        g404(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n427_));
  NA4        g405(.A(new_new_n148_), .B(new_new_n118_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n428_));
  OAI220     g406(.A0(new_new_n428_), .A1(new_new_n427_), .B0(new_new_n426_), .B1(new_new_n424_), .Y(new_new_n429_));
  NO3        g407(.A(new_new_n429_), .B(new_new_n423_), .C(new_new_n414_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n99_), .B(i_13_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n388_), .B(new_new_n350_), .Y(new_new_n432_));
  NO2        g410(.A(i_2_), .B(i_13_), .Y(new_new_n433_));
  NO2        g411(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n434_));
  NO3        g412(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n435_));
  NO2        g413(.A(i_6_), .B(i_7_), .Y(new_new_n436_));
  NO2        g414(.A(i_11_), .B(i_1_), .Y(new_new_n437_));
  OR2        g415(.A(i_11_), .B(i_8_), .Y(new_new_n438_));
  NOi21      g416(.An(i_2_), .B(i_7_), .Y(new_new_n439_));
  NO2        g417(.A(i_6_), .B(i_10_), .Y(new_new_n440_));
  NA3        g418(.A(new_new_n231_), .B(new_new_n172_), .C(new_new_n135_), .Y(new_new_n441_));
  NA2        g419(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n442_));
  NO2        g420(.A(new_new_n158_), .B(i_3_), .Y(new_new_n443_));
  NAi31      g421(.An(new_new_n442_), .B(new_new_n443_), .C(new_new_n216_), .Y(new_new_n444_));
  NA3        g422(.A(new_new_n363_), .B(new_new_n176_), .C(new_new_n152_), .Y(new_new_n445_));
  NA3        g423(.A(new_new_n445_), .B(new_new_n444_), .C(new_new_n441_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n446_), .B(new_new_n434_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n416_), .B(new_new_n351_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n425_), .B(new_new_n358_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n449_), .B(new_new_n214_), .Y(new_new_n450_));
  NAi21      g428(.An(new_new_n208_), .B(new_new_n367_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n313_), .B(new_new_n209_), .Y(new_new_n452_));
  NO2        g430(.A(new_new_n26_), .B(i_5_), .Y(new_new_n453_));
  NO2        g431(.A(i_0_), .B(new_new_n86_), .Y(new_new_n454_));
  NA3        g432(.A(new_new_n454_), .B(new_new_n453_), .C(new_new_n145_), .Y(new_new_n455_));
  OR3        g433(.A(new_new_n285_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n456_));
  OAI220     g434(.A0(new_new_n456_), .A1(new_new_n455_), .B0(new_new_n452_), .B1(new_new_n451_), .Y(new_new_n457_));
  NA2        g435(.A(new_new_n27_), .B(i_10_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n291_), .B(new_new_n225_), .Y(new_new_n459_));
  OAI220     g437(.A0(new_new_n459_), .A1(new_new_n396_), .B0(new_new_n458_), .B1(new_new_n431_), .Y(new_new_n460_));
  NO3        g438(.A(new_new_n460_), .B(new_new_n457_), .C(new_new_n450_), .Y(new_new_n461_));
  NA3        g439(.A(new_new_n461_), .B(new_new_n447_), .C(new_new_n430_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n125_), .B(new_new_n114_), .Y(new_new_n463_));
  AN2        g441(.A(new_new_n463_), .B(new_new_n416_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n464_), .B(new_new_n288_), .Y(new_new_n465_));
  NA4        g443(.A(new_new_n406_), .B(new_new_n405_), .C(new_new_n195_), .D(i_2_), .Y(new_new_n466_));
  INV        g444(.A(new_new_n466_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n351_), .B(new_new_n215_), .Y(new_new_n468_));
  NA2        g446(.A(new_new_n324_), .B(new_new_n73_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n338_), .B(new_new_n330_), .Y(new_new_n470_));
  OR2        g448(.A(new_new_n468_), .B(new_new_n470_), .Y(new_new_n471_));
  NO2        g449(.A(new_new_n36_), .B(i_8_), .Y(new_new_n472_));
  AOI210     g450(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n380_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n473_), .B(new_new_n471_), .Y(new_new_n474_));
  AOI210     g452(.A0(new_new_n467_), .A1(new_new_n196_), .B0(new_new_n474_), .Y(new_new_n475_));
  NA2        g453(.A(new_new_n238_), .B(new_new_n64_), .Y(new_new_n476_));
  OAI210     g454(.A0(i_8_), .A1(new_new_n476_), .B0(new_new_n137_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n477_), .B(new_new_n381_), .Y(new_new_n478_));
  NA3        g456(.A(new_new_n478_), .B(new_new_n475_), .C(new_new_n465_), .Y(new_new_n479_));
  NO2        g457(.A(i_12_), .B(new_new_n189_), .Y(new_new_n480_));
  NO2        g458(.A(i_8_), .B(i_7_), .Y(new_new_n481_));
  OAI210     g459(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n482_), .B(new_new_n213_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n228_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n44_), .B(i_10_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n485_), .B(i_6_), .Y(new_new_n486_));
  NA3        g464(.A(new_new_n486_), .B(new_new_n484_), .C(new_new_n481_), .Y(new_new_n487_));
  AOI220     g465(.A0(new_new_n388_), .A1(new_new_n301_), .B0(new_new_n232_), .B1(new_new_n230_), .Y(new_new_n488_));
  OAI220     g466(.A0(new_new_n488_), .A1(new_new_n245_), .B0(new_new_n431_), .B1(new_new_n136_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n489_), .B(new_new_n248_), .Y(new_new_n490_));
  NA3        g468(.A(new_new_n286_), .B(new_new_n174_), .C(new_new_n99_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n211_), .B(new_new_n44_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n158_), .B(i_5_), .Y(new_new_n493_));
  NA3        g471(.A(new_new_n493_), .B(new_new_n371_), .C(new_new_n297_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n494_), .A1(new_new_n492_), .B0(new_new_n491_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n425_), .Y(new_new_n496_));
  NA3        g474(.A(new_new_n496_), .B(new_new_n490_), .C(new_new_n487_), .Y(new_new_n497_));
  NA3        g475(.A(new_new_n209_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n267_), .B(new_new_n84_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n498_), .B(new_new_n499_), .Y(new_new_n500_));
  NA2        g478(.A(new_new_n213_), .B(new_new_n212_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n408_), .B(new_new_n211_), .Y(new_new_n502_));
  NO2        g480(.A(new_new_n501_), .B(new_new_n502_), .Y(new_new_n503_));
  AOI210     g481(.A0(new_new_n331_), .A1(new_new_n46_), .B0(new_new_n335_), .Y(new_new_n504_));
  NA2        g482(.A(i_0_), .B(new_new_n48_), .Y(new_new_n505_));
  NA3        g483(.A(new_new_n480_), .B(new_new_n258_), .C(new_new_n505_), .Y(new_new_n506_));
  NO2        g484(.A(new_new_n504_), .B(new_new_n506_), .Y(new_new_n507_));
  NO3        g485(.A(new_new_n507_), .B(new_new_n503_), .C(new_new_n500_), .Y(new_new_n508_));
  NO4        g486(.A(new_new_n234_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n509_));
  NO3        g487(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n221_), .B(new_new_n36_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n379_), .B(i_1_), .Y(new_new_n512_));
  NOi31      g490(.An(new_new_n512_), .B(new_new_n417_), .C(new_new_n73_), .Y(new_new_n513_));
  AN4        g491(.A(new_new_n513_), .B(new_new_n377_), .C(new_new_n453_), .D(i_2_), .Y(new_new_n514_));
  INV        g492(.A(new_new_n514_), .Y(new_new_n515_));
  NOi21      g493(.An(i_10_), .B(i_6_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n517_));
  AOI220     g495(.A0(new_new_n267_), .A1(new_new_n517_), .B0(new_new_n258_), .B1(new_new_n516_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(new_new_n415_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n294_), .B(new_new_n165_), .Y(new_new_n521_));
  AOI220     g499(.A0(new_new_n521_), .A1(new_new_n397_), .B0(new_new_n181_), .B1(new_new_n179_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n193_), .B(new_new_n37_), .Y(new_new_n523_));
  NOi31      g501(.An(new_new_n149_), .B(new_new_n523_), .C(new_new_n308_), .Y(new_new_n524_));
  NO3        g502(.A(new_new_n524_), .B(new_new_n522_), .C(new_new_n519_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n469_), .B(new_new_n346_), .Y(new_new_n526_));
  INV        g504(.A(new_new_n297_), .Y(new_new_n527_));
  NO2        g505(.A(i_12_), .B(new_new_n86_), .Y(new_new_n528_));
  NA3        g506(.A(new_new_n528_), .B(new_new_n258_), .C(new_new_n505_), .Y(new_new_n529_));
  NA3        g507(.A(new_new_n354_), .B(new_new_n267_), .C(new_new_n209_), .Y(new_new_n530_));
  AOI210     g508(.A0(new_new_n530_), .A1(new_new_n529_), .B0(new_new_n527_), .Y(new_new_n531_));
  OR2        g509(.A(i_2_), .B(i_5_), .Y(new_new_n532_));
  OR2        g510(.A(new_new_n532_), .B(new_new_n374_), .Y(new_new_n533_));
  AOI210     g511(.A0(new_new_n340_), .A1(new_new_n230_), .B0(new_new_n193_), .Y(new_new_n534_));
  AOI210     g512(.A0(new_new_n534_), .A1(new_new_n533_), .B0(new_new_n451_), .Y(new_new_n535_));
  NO3        g513(.A(new_new_n535_), .B(new_new_n531_), .C(new_new_n526_), .Y(new_new_n536_));
  NA4        g514(.A(new_new_n536_), .B(new_new_n525_), .C(new_new_n515_), .D(new_new_n508_), .Y(new_new_n537_));
  NO4        g515(.A(new_new_n537_), .B(new_new_n497_), .C(new_new_n479_), .D(new_new_n462_), .Y(new_new_n538_));
  NA4        g516(.A(new_new_n538_), .B(new_new_n404_), .C(new_new_n323_), .D(new_new_n290_), .Y(ori7));
  NO2        g517(.A(new_new_n95_), .B(new_new_n54_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n111_), .B(new_new_n92_), .Y(new_new_n541_));
  NA2        g519(.A(new_new_n352_), .B(new_new_n541_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n440_), .B(new_new_n84_), .Y(new_new_n543_));
  NA2        g521(.A(i_11_), .B(new_new_n189_), .Y(new_new_n544_));
  NA2        g522(.A(new_new_n147_), .B(new_new_n544_), .Y(new_new_n545_));
  OAI210     g523(.A0(new_new_n545_), .A1(new_new_n543_), .B0(new_new_n542_), .Y(new_new_n546_));
  NA3        g524(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n223_), .B(i_4_), .Y(new_new_n548_));
  NA2        g526(.A(new_new_n548_), .B(i_8_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n108_), .B(new_new_n547_), .Y(new_new_n550_));
  NA2        g528(.A(i_2_), .B(new_new_n86_), .Y(new_new_n551_));
  OAI210     g529(.A0(new_new_n89_), .A1(new_new_n195_), .B0(new_new_n196_), .Y(new_new_n552_));
  NO2        g530(.A(i_7_), .B(new_new_n37_), .Y(new_new_n553_));
  NA2        g531(.A(i_4_), .B(i_8_), .Y(new_new_n554_));
  AOI210     g532(.A0(new_new_n554_), .A1(new_new_n286_), .B0(new_new_n553_), .Y(new_new_n555_));
  OAI220     g533(.A0(new_new_n555_), .A1(new_new_n551_), .B0(new_new_n552_), .B1(i_13_), .Y(new_new_n556_));
  NO4        g534(.A(new_new_n556_), .B(new_new_n550_), .C(new_new_n546_), .D(new_new_n540_), .Y(new_new_n557_));
  AOI210     g535(.A0(new_new_n131_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n558_));
  AOI210     g536(.A0(new_new_n558_), .A1(new_new_n223_), .B0(new_new_n162_), .Y(new_new_n559_));
  OR2        g537(.A(i_6_), .B(i_10_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n560_), .B(new_new_n23_), .Y(new_new_n561_));
  OR3        g539(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n562_));
  INV        g540(.A(new_new_n194_), .Y(new_new_n563_));
  INV        g541(.A(new_new_n561_), .Y(new_new_n564_));
  OA220      g542(.A0(new_new_n564_), .A1(new_new_n527_), .B0(new_new_n559_), .B1(new_new_n250_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n565_), .A1(new_new_n557_), .B0(new_new_n63_), .Y(new_new_n566_));
  NOi21      g544(.An(i_11_), .B(i_7_), .Y(new_new_n567_));
  AO210      g545(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n568_));
  NO2        g546(.A(new_new_n568_), .B(new_new_n567_), .Y(new_new_n569_));
  NA2        g547(.A(new_new_n569_), .B(new_new_n200_), .Y(new_new_n570_));
  NA3        g548(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n571_));
  NAi31      g549(.An(new_new_n571_), .B(new_new_n207_), .C(i_11_), .Y(new_new_n572_));
  AOI210     g550(.A0(new_new_n572_), .A1(new_new_n570_), .B0(new_new_n63_), .Y(new_new_n573_));
  NA2        g551(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n574_));
  AO210      g552(.A0(new_new_n574_), .A1(new_new_n346_), .B0(new_new_n41_), .Y(new_new_n575_));
  NO3        g553(.A(new_new_n240_), .B(new_new_n201_), .C(new_new_n544_), .Y(new_new_n576_));
  OAI210     g554(.A0(new_new_n576_), .A1(new_new_n216_), .B0(new_new_n63_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n375_), .B(new_new_n31_), .Y(new_new_n578_));
  OR2        g556(.A(new_new_n201_), .B(new_new_n111_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n579_), .B(new_new_n578_), .Y(new_new_n580_));
  NO2        g558(.A(i_1_), .B(i_4_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n581_), .B(new_new_n580_), .Y(new_new_n582_));
  NO2        g560(.A(i_1_), .B(i_12_), .Y(new_new_n583_));
  NA3        g561(.A(new_new_n583_), .B(new_new_n112_), .C(new_new_n24_), .Y(new_new_n584_));
  BUFFER     g562(.A(new_new_n584_), .Y(new_new_n585_));
  NA4        g563(.A(new_new_n585_), .B(new_new_n582_), .C(new_new_n577_), .D(new_new_n575_), .Y(new_new_n586_));
  OAI210     g564(.A0(new_new_n586_), .A1(new_new_n573_), .B0(i_6_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n571_), .B(new_new_n111_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(new_new_n528_), .Y(new_new_n589_));
  NO2        g567(.A(new_new_n223_), .B(new_new_n86_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n590_), .B(i_11_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n589_), .B(new_new_n418_), .Y(new_new_n592_));
  NO3        g570(.A(new_new_n560_), .B(new_new_n221_), .C(new_new_n23_), .Y(new_new_n593_));
  AOI210     g571(.A0(i_1_), .A1(new_new_n241_), .B0(new_new_n593_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n594_), .B(new_new_n44_), .Y(new_new_n595_));
  NA3        g573(.A(new_new_n481_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n596_));
  INV        g574(.A(i_2_), .Y(new_new_n597_));
  NA2        g575(.A(new_new_n141_), .B(i_9_), .Y(new_new_n598_));
  NA3        g576(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n46_), .B(i_1_), .Y(new_new_n600_));
  NA3        g578(.A(new_new_n600_), .B(new_new_n249_), .C(new_new_n44_), .Y(new_new_n601_));
  OAI220     g579(.A0(new_new_n601_), .A1(new_new_n599_), .B0(new_new_n598_), .B1(new_new_n597_), .Y(new_new_n602_));
  AOI210     g580(.A0(new_new_n437_), .A1(new_new_n382_), .B0(new_new_n227_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n603_), .B(new_new_n551_), .Y(new_new_n604_));
  NAi21      g582(.An(new_new_n596_), .B(new_new_n94_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n600_), .B(new_new_n249_), .Y(new_new_n606_));
  NO2        g584(.A(i_11_), .B(new_new_n37_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n607_), .B(new_new_n24_), .Y(new_new_n608_));
  OAI210     g586(.A0(new_new_n608_), .A1(new_new_n606_), .B0(new_new_n605_), .Y(new_new_n609_));
  OR3        g587(.A(new_new_n609_), .B(new_new_n604_), .C(new_new_n602_), .Y(new_new_n610_));
  NO3        g588(.A(new_new_n610_), .B(new_new_n595_), .C(new_new_n592_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n223_), .B(new_new_n104_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n567_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n613_), .B(i_1_), .Y(new_new_n614_));
  NO2        g592(.A(new_new_n614_), .B(new_new_n562_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n378_), .B(new_new_n86_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n615_), .B(new_new_n46_), .Y(new_new_n617_));
  NA2        g595(.A(i_3_), .B(new_new_n189_), .Y(new_new_n618_));
  NO2        g596(.A(new_new_n618_), .B(new_new_n117_), .Y(new_new_n619_));
  AN2        g597(.A(new_new_n619_), .B(new_new_n486_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n221_), .B(new_new_n44_), .Y(new_new_n621_));
  NO3        g599(.A(new_new_n621_), .B(new_new_n288_), .C(new_new_n224_), .Y(new_new_n622_));
  NO2        g600(.A(new_new_n120_), .B(new_new_n37_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n623_), .B(i_6_), .Y(new_new_n624_));
  NO2        g602(.A(new_new_n86_), .B(i_9_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n63_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n626_), .B(new_new_n583_), .Y(new_new_n627_));
  NO4        g605(.A(new_new_n627_), .B(new_new_n624_), .C(new_new_n622_), .D(i_4_), .Y(new_new_n628_));
  NA2        g606(.A(i_1_), .B(i_3_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n419_), .B(new_new_n95_), .Y(new_new_n630_));
  AOI210     g608(.A0(new_new_n621_), .A1(new_new_n516_), .B0(new_new_n630_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n629_), .Y(new_new_n632_));
  NO3        g610(.A(new_new_n632_), .B(new_new_n628_), .C(new_new_n620_), .Y(new_new_n633_));
  NA4        g611(.A(new_new_n633_), .B(new_new_n617_), .C(new_new_n611_), .D(new_new_n587_), .Y(new_new_n634_));
  NO3        g612(.A(new_new_n438_), .B(i_3_), .C(i_7_), .Y(new_new_n635_));
  NOi21      g613(.An(new_new_n635_), .B(i_10_), .Y(new_new_n636_));
  OA210      g614(.A0(new_new_n636_), .A1(new_new_n231_), .B0(new_new_n86_), .Y(new_new_n637_));
  NO3        g615(.A(new_new_n439_), .B(new_new_n554_), .C(new_new_n86_), .Y(new_new_n638_));
  NA2        g616(.A(new_new_n638_), .B(new_new_n25_), .Y(new_new_n639_));
  INV        g617(.A(new_new_n639_), .Y(new_new_n640_));
  OAI210     g618(.A0(new_new_n640_), .A1(new_new_n637_), .B0(i_1_), .Y(new_new_n641_));
  AOI210     g619(.A0(new_new_n249_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n336_), .B(i_2_), .Y(new_new_n643_));
  NA2        g621(.A(new_new_n643_), .B(new_new_n642_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n644_), .A1(new_new_n641_), .B0(i_13_), .Y(new_new_n645_));
  OR2        g623(.A(i_11_), .B(i_7_), .Y(new_new_n646_));
  NA3        g624(.A(new_new_n646_), .B(new_new_n109_), .C(new_new_n141_), .Y(new_new_n647_));
  AOI220     g625(.A0(new_new_n433_), .A1(new_new_n162_), .B0(new_new_n412_), .B1(new_new_n141_), .Y(new_new_n648_));
  OAI210     g626(.A0(new_new_n648_), .A1(new_new_n44_), .B0(new_new_n647_), .Y(new_new_n649_));
  AOI210     g627(.A0(new_new_n599_), .A1(new_new_n54_), .B0(i_12_), .Y(new_new_n650_));
  NO2        g628(.A(new_new_n439_), .B(new_new_n24_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n651_), .B(new_new_n616_), .Y(new_new_n652_));
  OAI220     g630(.A0(new_new_n652_), .A1(new_new_n41_), .B0(new_new_n973_), .B1(new_new_n95_), .Y(new_new_n653_));
  AOI210     g631(.A0(new_new_n649_), .A1(new_new_n310_), .B0(new_new_n653_), .Y(new_new_n654_));
  NA2        g632(.A(new_new_n354_), .B(new_new_n600_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n655_), .B(new_new_n228_), .Y(new_new_n656_));
  AOI210     g634(.A0(new_new_n409_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n657_));
  NOi31      g635(.An(new_new_n657_), .B(new_new_n543_), .C(new_new_n44_), .Y(new_new_n658_));
  NA2        g636(.A(new_new_n130_), .B(i_13_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n599_), .B(new_new_n117_), .Y(new_new_n660_));
  INV        g638(.A(new_new_n660_), .Y(new_new_n661_));
  OAI220     g639(.A0(new_new_n661_), .A1(new_new_n71_), .B0(new_new_n659_), .B1(new_new_n642_), .Y(new_new_n662_));
  NO3        g640(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n26_), .B(new_new_n189_), .Y(new_new_n664_));
  NA2        g642(.A(new_new_n664_), .B(i_7_), .Y(new_new_n665_));
  INV        g643(.A(new_new_n663_), .Y(new_new_n666_));
  AOI220     g644(.A0(new_new_n354_), .A1(new_new_n600_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n667_));
  OAI220     g645(.A0(new_new_n667_), .A1(new_new_n549_), .B0(new_new_n666_), .B1(new_new_n563_), .Y(new_new_n668_));
  NO4        g646(.A(new_new_n668_), .B(new_new_n662_), .C(new_new_n658_), .D(new_new_n656_), .Y(new_new_n669_));
  OR2        g647(.A(i_11_), .B(i_6_), .Y(new_new_n670_));
  NA3        g648(.A(new_new_n548_), .B(new_new_n664_), .C(i_7_), .Y(new_new_n671_));
  AOI210     g649(.A0(new_new_n671_), .A1(new_new_n661_), .B0(new_new_n670_), .Y(new_new_n672_));
  NA3        g650(.A(new_new_n375_), .B(new_new_n553_), .C(new_new_n100_), .Y(new_new_n673_));
  NA2        g651(.A(new_new_n591_), .B(i_13_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n105_), .B(new_new_n664_), .Y(new_new_n675_));
  NAi21      g653(.An(i_11_), .B(i_12_), .Y(new_new_n676_));
  NOi41      g654(.An(new_new_n113_), .B(new_new_n676_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n677_));
  NO3        g655(.A(new_new_n439_), .B(new_new_n528_), .C(new_new_n554_), .Y(new_new_n678_));
  AOI220     g656(.A0(new_new_n678_), .A1(new_new_n291_), .B0(new_new_n677_), .B1(new_new_n675_), .Y(new_new_n679_));
  NA3        g657(.A(new_new_n679_), .B(new_new_n674_), .C(new_new_n673_), .Y(new_new_n680_));
  OAI210     g658(.A0(new_new_n680_), .A1(new_new_n672_), .B0(new_new_n63_), .Y(new_new_n681_));
  NO2        g659(.A(i_2_), .B(i_12_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n335_), .B(new_new_n682_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n337_), .B(new_new_n335_), .Y(new_new_n684_));
  NO2        g662(.A(new_new_n131_), .B(i_2_), .Y(new_new_n685_));
  NA2        g663(.A(new_new_n685_), .B(new_new_n583_), .Y(new_new_n686_));
  NA3        g664(.A(new_new_n686_), .B(new_new_n684_), .C(new_new_n683_), .Y(new_new_n687_));
  NA3        g665(.A(new_new_n687_), .B(new_new_n45_), .C(new_new_n215_), .Y(new_new_n688_));
  NA4        g666(.A(new_new_n688_), .B(new_new_n681_), .C(new_new_n669_), .D(new_new_n654_), .Y(new_new_n689_));
  OR4        g667(.A(new_new_n689_), .B(new_new_n645_), .C(new_new_n634_), .D(new_new_n566_), .Y(ori5));
  NA2        g668(.A(new_new_n613_), .B(new_new_n252_), .Y(new_new_n691_));
  AN2        g669(.A(new_new_n24_), .B(i_10_), .Y(new_new_n692_));
  NA3        g670(.A(new_new_n692_), .B(new_new_n682_), .C(new_new_n111_), .Y(new_new_n693_));
  NO2        g671(.A(new_new_n549_), .B(i_11_), .Y(new_new_n694_));
  NA2        g672(.A(new_new_n89_), .B(new_new_n694_), .Y(new_new_n695_));
  NA3        g673(.A(new_new_n695_), .B(new_new_n693_), .C(new_new_n691_), .Y(new_new_n696_));
  NO3        g674(.A(i_11_), .B(new_new_n223_), .C(i_13_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n127_), .B(new_new_n23_), .Y(new_new_n698_));
  NA2        g676(.A(i_12_), .B(i_8_), .Y(new_new_n699_));
  OAI210     g677(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n699_), .Y(new_new_n700_));
  INV        g678(.A(new_new_n408_), .Y(new_new_n701_));
  AOI220     g679(.A0(new_new_n297_), .A1(new_new_n520_), .B0(new_new_n700_), .B1(new_new_n698_), .Y(new_new_n702_));
  INV        g680(.A(new_new_n702_), .Y(new_new_n703_));
  NO2        g681(.A(new_new_n703_), .B(new_new_n696_), .Y(new_new_n704_));
  INV        g682(.A(new_new_n172_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n231_), .Y(new_new_n706_));
  OAI210     g684(.A0(new_new_n643_), .A1(new_new_n410_), .B0(new_new_n113_), .Y(new_new_n707_));
  AOI210     g685(.A0(new_new_n707_), .A1(new_new_n706_), .B0(new_new_n705_), .Y(new_new_n708_));
  NO2        g686(.A(new_new_n419_), .B(new_new_n26_), .Y(new_new_n709_));
  NO2        g687(.A(new_new_n709_), .B(new_new_n382_), .Y(new_new_n710_));
  NA2        g688(.A(new_new_n710_), .B(i_2_), .Y(new_new_n711_));
  INV        g689(.A(new_new_n711_), .Y(new_new_n712_));
  AOI210     g690(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n379_), .Y(new_new_n713_));
  AOI210     g691(.A0(new_new_n713_), .A1(new_new_n712_), .B0(new_new_n708_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n187_), .B(new_new_n128_), .Y(new_new_n715_));
  OAI210     g693(.A0(new_new_n715_), .A1(new_new_n698_), .B0(i_2_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n173_), .Y(new_new_n717_));
  NO3        g695(.A(new_new_n568_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n718_));
  AOI210     g696(.A0(new_new_n717_), .A1(new_new_n89_), .B0(new_new_n718_), .Y(new_new_n719_));
  AOI210     g697(.A0(new_new_n719_), .A1(new_new_n716_), .B0(new_new_n189_), .Y(new_new_n720_));
  OA210      g698(.A0(new_new_n569_), .A1(new_new_n129_), .B0(i_13_), .Y(new_new_n721_));
  NA2        g699(.A(new_new_n194_), .B(new_new_n195_), .Y(new_new_n722_));
  NA2        g700(.A(new_new_n154_), .B(new_new_n544_), .Y(new_new_n723_));
  AOI210     g701(.A0(new_new_n723_), .A1(new_new_n722_), .B0(new_new_n340_), .Y(new_new_n724_));
  AOI210     g702(.A0(new_new_n201_), .A1(new_new_n151_), .B0(new_new_n472_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(new_new_n382_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n105_), .B(new_new_n44_), .Y(new_new_n727_));
  INV        g705(.A(new_new_n284_), .Y(new_new_n728_));
  NA4        g706(.A(new_new_n728_), .B(new_new_n286_), .C(new_new_n127_), .D(new_new_n42_), .Y(new_new_n729_));
  OAI210     g707(.A0(new_new_n729_), .A1(new_new_n727_), .B0(new_new_n726_), .Y(new_new_n730_));
  NO4        g708(.A(new_new_n730_), .B(new_new_n724_), .C(new_new_n721_), .D(new_new_n720_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n520_), .B(new_new_n28_), .Y(new_new_n732_));
  NA2        g710(.A(new_new_n697_), .B(new_new_n259_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n733_), .B(new_new_n732_), .Y(new_new_n734_));
  NO2        g712(.A(new_new_n62_), .B(i_12_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n735_), .B(new_new_n129_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n736_), .B(new_new_n544_), .Y(new_new_n737_));
  AOI220     g715(.A0(new_new_n737_), .A1(new_new_n36_), .B0(new_new_n734_), .B1(new_new_n46_), .Y(new_new_n738_));
  NA4        g716(.A(new_new_n738_), .B(new_new_n731_), .C(new_new_n714_), .D(new_new_n704_), .Y(ori6));
  NO3        g717(.A(i_9_), .B(new_new_n287_), .C(i_1_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n740_), .B(new_new_n685_), .Y(new_new_n741_));
  NO2        g719(.A(new_new_n210_), .B(new_new_n442_), .Y(new_new_n742_));
  INV        g720(.A(new_new_n305_), .Y(new_new_n743_));
  AO210      g721(.A0(new_new_n743_), .A1(new_new_n741_), .B0(i_12_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n528_), .B(new_new_n63_), .Y(new_new_n745_));
  NA2        g723(.A(new_new_n636_), .B(new_new_n71_), .Y(new_new_n746_));
  BUFFER     g724(.A(new_new_n574_), .Y(new_new_n747_));
  NA3        g725(.A(new_new_n747_), .B(new_new_n746_), .C(new_new_n745_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n748_), .B(new_new_n73_), .Y(new_new_n749_));
  INV        g727(.A(new_new_n304_), .Y(new_new_n750_));
  NA2        g728(.A(new_new_n75_), .B(new_new_n134_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n127_), .Y(new_new_n752_));
  NA2        g730(.A(new_new_n752_), .B(new_new_n46_), .Y(new_new_n753_));
  AOI210     g731(.A0(new_new_n753_), .A1(new_new_n751_), .B0(new_new_n750_), .Y(new_new_n754_));
  NO3        g732(.A(new_new_n234_), .B(new_new_n135_), .C(i_9_), .Y(new_new_n755_));
  NA2        g733(.A(new_new_n755_), .B(new_new_n735_), .Y(new_new_n756_));
  AOI210     g734(.A0(new_new_n756_), .A1(new_new_n470_), .B0(new_new_n183_), .Y(new_new_n757_));
  NO2        g735(.A(new_new_n32_), .B(i_11_), .Y(new_new_n758_));
  NA3        g736(.A(new_new_n758_), .B(new_new_n436_), .C(new_new_n358_), .Y(new_new_n759_));
  NAi32      g737(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n670_), .B(new_new_n760_), .Y(new_new_n761_));
  OAI210     g739(.A0(new_new_n635_), .A1(new_new_n511_), .B0(new_new_n510_), .Y(new_new_n762_));
  NAi31      g740(.An(new_new_n761_), .B(new_new_n762_), .C(new_new_n759_), .Y(new_new_n763_));
  OR3        g741(.A(new_new_n763_), .B(new_new_n757_), .C(new_new_n754_), .Y(new_new_n764_));
  NO2        g742(.A(new_new_n646_), .B(i_2_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n766_), .B(new_new_n374_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n767_), .B(new_new_n765_), .Y(new_new_n768_));
  OR2        g746(.A(new_new_n569_), .B(new_new_n410_), .Y(new_new_n769_));
  NA3        g747(.A(new_new_n769_), .B(new_new_n150_), .C(new_new_n69_), .Y(new_new_n770_));
  AO210      g748(.A0(new_new_n449_), .A1(new_new_n701_), .B0(new_new_n36_), .Y(new_new_n771_));
  NA3        g749(.A(new_new_n771_), .B(new_new_n770_), .C(new_new_n768_), .Y(new_new_n772_));
  OAI210     g750(.A0(new_new_n590_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n773_));
  AOI220     g751(.A0(new_new_n773_), .A1(new_new_n510_), .B0(new_new_n742_), .B1(new_new_n665_), .Y(new_new_n774_));
  NA3        g752(.A(new_new_n340_), .B(new_new_n225_), .C(new_new_n150_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n366_), .B(new_new_n70_), .Y(new_new_n776_));
  NA4        g754(.A(new_new_n776_), .B(new_new_n775_), .C(new_new_n774_), .D(new_new_n552_), .Y(new_new_n777_));
  AO210      g755(.A0(new_new_n472_), .A1(new_new_n46_), .B0(new_new_n88_), .Y(new_new_n778_));
  NA3        g756(.A(new_new_n778_), .B(new_new_n440_), .C(new_new_n209_), .Y(new_new_n779_));
  AOI210     g757(.A0(new_new_n410_), .A1(new_new_n408_), .B0(new_new_n509_), .Y(new_new_n780_));
  NO2        g758(.A(new_new_n560_), .B(new_new_n105_), .Y(new_new_n781_));
  OAI210     g759(.A0(new_new_n781_), .A1(new_new_n114_), .B0(new_new_n373_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n230_), .B(new_new_n46_), .Y(new_new_n783_));
  INV        g761(.A(new_new_n533_), .Y(new_new_n784_));
  NA3        g762(.A(new_new_n784_), .B(new_new_n304_), .C(i_7_), .Y(new_new_n785_));
  NA4        g763(.A(new_new_n785_), .B(new_new_n782_), .C(new_new_n780_), .D(new_new_n779_), .Y(new_new_n786_));
  NO4        g764(.A(new_new_n786_), .B(new_new_n777_), .C(new_new_n772_), .D(new_new_n764_), .Y(new_new_n787_));
  NA4        g765(.A(new_new_n787_), .B(new_new_n749_), .C(new_new_n744_), .D(new_new_n348_), .Y(ori3));
  NA2        g766(.A(i_12_), .B(i_10_), .Y(new_new_n789_));
  NO2        g767(.A(i_11_), .B(new_new_n223_), .Y(new_new_n790_));
  NA3        g768(.A(new_new_n775_), .B(new_new_n552_), .C(new_new_n339_), .Y(new_new_n791_));
  NA2        g769(.A(new_new_n791_), .B(new_new_n40_), .Y(new_new_n792_));
  NOi21      g770(.An(new_new_n99_), .B(new_new_n710_), .Y(new_new_n793_));
  NO3        g771(.A(new_new_n579_), .B(new_new_n419_), .C(new_new_n134_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n375_), .B(new_new_n45_), .Y(new_new_n795_));
  AN2        g773(.A(new_new_n417_), .B(new_new_n55_), .Y(new_new_n796_));
  NO3        g774(.A(new_new_n796_), .B(new_new_n794_), .C(new_new_n793_), .Y(new_new_n797_));
  AOI210     g775(.A0(new_new_n797_), .A1(new_new_n792_), .B0(new_new_n48_), .Y(new_new_n798_));
  NO4        g776(.A(new_new_n344_), .B(new_new_n351_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n799_));
  NA2        g777(.A(new_new_n183_), .B(new_new_n516_), .Y(new_new_n800_));
  NOi21      g778(.An(new_new_n800_), .B(new_new_n799_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n657_), .B(new_new_n625_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n311_), .B(new_new_n399_), .Y(new_new_n803_));
  OAI220     g781(.A0(new_new_n803_), .A1(new_new_n802_), .B0(new_new_n801_), .B1(new_new_n63_), .Y(new_new_n804_));
  NOi21      g782(.An(i_5_), .B(i_9_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n805_), .B(new_new_n406_), .Y(new_new_n806_));
  BUFFER     g784(.A(new_new_n249_), .Y(new_new_n807_));
  AOI210     g785(.A0(new_new_n807_), .A1(new_new_n437_), .B0(new_new_n638_), .Y(new_new_n808_));
  NO3        g786(.A(new_new_n376_), .B(new_new_n249_), .C(new_new_n73_), .Y(new_new_n809_));
  NO2        g787(.A(new_new_n175_), .B(new_new_n151_), .Y(new_new_n810_));
  AOI210     g788(.A0(new_new_n810_), .A1(new_new_n230_), .B0(new_new_n809_), .Y(new_new_n811_));
  OAI220     g789(.A0(new_new_n811_), .A1(new_new_n178_), .B0(new_new_n808_), .B1(new_new_n806_), .Y(new_new_n812_));
  NO3        g790(.A(new_new_n812_), .B(new_new_n804_), .C(new_new_n798_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n183_), .B(new_new_n24_), .Y(new_new_n814_));
  NO2        g792(.A(new_new_n623_), .B(new_new_n541_), .Y(new_new_n815_));
  NO2        g793(.A(new_new_n815_), .B(new_new_n814_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n291_), .B(new_new_n132_), .Y(new_new_n817_));
  NAi21      g795(.An(new_new_n163_), .B(new_new_n399_), .Y(new_new_n818_));
  OAI220     g796(.A0(new_new_n818_), .A1(new_new_n783_), .B0(new_new_n817_), .B1(new_new_n368_), .Y(new_new_n819_));
  NO2        g797(.A(new_new_n819_), .B(new_new_n816_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n517_), .B(i_0_), .Y(new_new_n821_));
  NO3        g799(.A(new_new_n821_), .B(new_new_n353_), .C(new_new_n89_), .Y(new_new_n822_));
  NO4        g800(.A(new_new_n532_), .B(new_new_n207_), .C(new_new_n379_), .D(new_new_n374_), .Y(new_new_n823_));
  AOI210     g801(.A0(new_new_n823_), .A1(i_11_), .B0(new_new_n822_), .Y(new_new_n824_));
  INV        g802(.A(new_new_n436_), .Y(new_new_n825_));
  AN2        g803(.A(new_new_n99_), .B(new_new_n229_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n697_), .B(new_new_n305_), .Y(new_new_n827_));
  AOI210     g805(.A0(new_new_n440_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n828_));
  OAI220     g806(.A0(new_new_n828_), .A1(new_new_n827_), .B0(new_new_n608_), .B1(new_new_n483_), .Y(new_new_n829_));
  NO2        g807(.A(new_new_n236_), .B(new_new_n155_), .Y(new_new_n830_));
  NA2        g808(.A(i_0_), .B(i_10_), .Y(new_new_n831_));
  INV        g809(.A(new_new_n485_), .Y(new_new_n832_));
  NO4        g810(.A(new_new_n117_), .B(new_new_n58_), .C(new_new_n618_), .D(i_5_), .Y(new_new_n833_));
  AO220      g811(.A0(new_new_n833_), .A1(new_new_n832_), .B0(new_new_n830_), .B1(i_6_), .Y(new_new_n834_));
  NA2        g812(.A(new_new_n186_), .B(new_new_n195_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n835_), .B(new_new_n827_), .Y(new_new_n836_));
  NO4        g814(.A(new_new_n836_), .B(new_new_n834_), .C(new_new_n829_), .D(new_new_n826_), .Y(new_new_n837_));
  NA3        g815(.A(new_new_n837_), .B(new_new_n824_), .C(new_new_n820_), .Y(new_new_n838_));
  NO2        g816(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n839_));
  NA2        g817(.A(i_11_), .B(i_9_), .Y(new_new_n840_));
  NO3        g818(.A(i_12_), .B(new_new_n840_), .C(new_new_n551_), .Y(new_new_n841_));
  AN2        g819(.A(new_new_n841_), .B(new_new_n839_), .Y(new_new_n842_));
  NO2        g820(.A(new_new_n48_), .B(i_7_), .Y(new_new_n843_));
  NA2        g821(.A(new_new_n363_), .B(new_new_n176_), .Y(new_new_n844_));
  NA2        g822(.A(new_new_n844_), .B(new_new_n161_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n840_), .B(new_new_n73_), .Y(new_new_n846_));
  NO2        g824(.A(new_new_n175_), .B(i_0_), .Y(new_new_n847_));
  INV        g825(.A(new_new_n372_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n848_), .B(new_new_n806_), .Y(new_new_n849_));
  NO3        g827(.A(new_new_n849_), .B(new_new_n845_), .C(new_new_n842_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n607_), .B(new_new_n124_), .Y(new_new_n851_));
  NO2        g829(.A(i_6_), .B(new_new_n851_), .Y(new_new_n852_));
  AOI210     g830(.A0(new_new_n409_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n853_));
  NA2        g831(.A(new_new_n172_), .B(new_new_n106_), .Y(new_new_n854_));
  NOi32      g832(.An(new_new_n853_), .Bn(new_new_n186_), .C(new_new_n854_), .Y(new_new_n855_));
  NA2        g833(.A(new_new_n553_), .B(new_new_n305_), .Y(new_new_n856_));
  NO2        g834(.A(new_new_n856_), .B(new_new_n795_), .Y(new_new_n857_));
  NO3        g835(.A(new_new_n857_), .B(new_new_n855_), .C(new_new_n852_), .Y(new_new_n858_));
  NOi21      g836(.An(i_7_), .B(i_5_), .Y(new_new_n859_));
  OR2        g837(.A(new_new_n854_), .B(new_new_n470_), .Y(new_new_n860_));
  INV        g838(.A(new_new_n298_), .Y(new_new_n861_));
  NA3        g839(.A(new_new_n860_), .B(new_new_n858_), .C(new_new_n850_), .Y(new_new_n862_));
  NO2        g840(.A(new_new_n789_), .B(new_new_n297_), .Y(new_new_n863_));
  OA210      g841(.A0(new_new_n436_), .A1(new_new_n213_), .B0(new_new_n435_), .Y(new_new_n864_));
  NA2        g842(.A(new_new_n863_), .B(new_new_n846_), .Y(new_new_n865_));
  NA3        g843(.A(new_new_n435_), .B(new_new_n375_), .C(new_new_n45_), .Y(new_new_n866_));
  OAI210     g844(.A0(new_new_n818_), .A1(new_new_n825_), .B0(new_new_n866_), .Y(new_new_n867_));
  NO2        g845(.A(i_2_), .B(new_new_n185_), .Y(new_new_n868_));
  AOI220     g846(.A0(new_new_n868_), .A1(new_new_n436_), .B0(new_new_n867_), .B1(new_new_n73_), .Y(new_new_n869_));
  NA3        g847(.A(new_new_n766_), .B(new_new_n350_), .C(new_new_n590_), .Y(new_new_n870_));
  NA2        g848(.A(new_new_n95_), .B(new_new_n44_), .Y(new_new_n871_));
  NO2        g849(.A(new_new_n75_), .B(new_new_n699_), .Y(new_new_n872_));
  AOI220     g850(.A0(new_new_n872_), .A1(new_new_n871_), .B0(new_new_n174_), .B1(new_new_n541_), .Y(new_new_n873_));
  AOI210     g851(.A0(new_new_n873_), .A1(new_new_n870_), .B0(new_new_n47_), .Y(new_new_n874_));
  NA2        g852(.A(new_new_n651_), .B(new_new_n493_), .Y(new_new_n875_));
  NO2        g853(.A(new_new_n875_), .B(new_new_n173_), .Y(new_new_n876_));
  NO3        g854(.A(new_new_n876_), .B(new_new_n874_), .C(new_new_n474_), .Y(new_new_n877_));
  NA3        g855(.A(new_new_n877_), .B(new_new_n869_), .C(new_new_n865_), .Y(new_new_n878_));
  NO3        g856(.A(new_new_n878_), .B(new_new_n862_), .C(new_new_n838_), .Y(new_new_n879_));
  NO2        g857(.A(i_0_), .B(new_new_n676_), .Y(new_new_n880_));
  NA2        g858(.A(new_new_n73_), .B(new_new_n44_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n745_), .B(new_new_n854_), .Y(new_new_n882_));
  INV        g860(.A(new_new_n882_), .Y(new_new_n883_));
  NO2        g861(.A(new_new_n762_), .B(new_new_n369_), .Y(new_new_n884_));
  NA2        g862(.A(new_new_n790_), .B(i_9_), .Y(new_new_n885_));
  NO2        g863(.A(new_new_n455_), .B(new_new_n885_), .Y(new_new_n886_));
  OAI210     g864(.A0(new_new_n230_), .A1(i_9_), .B0(new_new_n220_), .Y(new_new_n887_));
  AOI210     g865(.A0(new_new_n887_), .A1(new_new_n821_), .B0(new_new_n155_), .Y(new_new_n888_));
  NO3        g866(.A(new_new_n888_), .B(new_new_n886_), .C(new_new_n884_), .Y(new_new_n889_));
  NA2        g867(.A(new_new_n889_), .B(new_new_n883_), .Y(new_new_n890_));
  NO3        g868(.A(new_new_n831_), .B(new_new_n805_), .C(new_new_n187_), .Y(new_new_n891_));
  AOI220     g869(.A0(new_new_n891_), .A1(i_11_), .B0(new_new_n513_), .B1(new_new_n75_), .Y(new_new_n892_));
  NO3        g870(.A(new_new_n202_), .B(new_new_n351_), .C(i_0_), .Y(new_new_n893_));
  OAI210     g871(.A0(new_new_n893_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n894_));
  NA2        g872(.A(new_new_n894_), .B(new_new_n892_), .Y(new_new_n895_));
  NO2        g873(.A(new_new_n228_), .B(new_new_n95_), .Y(new_new_n896_));
  NA2        g874(.A(new_new_n896_), .B(new_new_n880_), .Y(new_new_n897_));
  OR2        g875(.A(new_new_n897_), .B(i_5_), .Y(new_new_n898_));
  AOI210     g876(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n175_), .Y(new_new_n899_));
  NA2        g877(.A(new_new_n899_), .B(new_new_n864_), .Y(new_new_n900_));
  INV        g878(.A(new_new_n491_), .Y(new_new_n901_));
  NO3        g879(.A(new_new_n795_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n448_), .B(new_new_n441_), .Y(new_new_n903_));
  NO3        g881(.A(new_new_n903_), .B(new_new_n902_), .C(new_new_n901_), .Y(new_new_n904_));
  NA3        g882(.A(new_new_n358_), .B(new_new_n172_), .C(new_new_n171_), .Y(new_new_n905_));
  INV        g883(.A(new_new_n905_), .Y(new_new_n906_));
  NA3        g884(.A(new_new_n358_), .B(new_new_n312_), .C(new_new_n211_), .Y(new_new_n907_));
  INV        g885(.A(new_new_n907_), .Y(new_new_n908_));
  NOi31      g886(.An(new_new_n357_), .B(new_new_n881_), .C(new_new_n226_), .Y(new_new_n909_));
  NO3        g887(.A(new_new_n840_), .B(new_new_n209_), .C(new_new_n187_), .Y(new_new_n910_));
  NO4        g888(.A(new_new_n910_), .B(new_new_n909_), .C(new_new_n908_), .D(new_new_n906_), .Y(new_new_n911_));
  NA4        g889(.A(new_new_n911_), .B(new_new_n904_), .C(new_new_n900_), .D(new_new_n898_), .Y(new_new_n912_));
  NO2        g890(.A(new_new_n86_), .B(i_5_), .Y(new_new_n913_));
  NA3        g891(.A(new_new_n790_), .B(new_new_n112_), .C(new_new_n127_), .Y(new_new_n914_));
  INV        g892(.A(new_new_n914_), .Y(new_new_n915_));
  NA2        g893(.A(new_new_n915_), .B(new_new_n913_), .Y(new_new_n916_));
  NA3        g894(.A(new_new_n286_), .B(i_5_), .C(new_new_n189_), .Y(new_new_n917_));
  NAi31      g895(.An(new_new_n227_), .B(new_new_n917_), .C(new_new_n228_), .Y(new_new_n918_));
  NO4        g896(.A(new_new_n226_), .B(new_new_n202_), .C(i_0_), .D(i_12_), .Y(new_new_n919_));
  NA2        g897(.A(new_new_n919_), .B(new_new_n918_), .Y(new_new_n920_));
  AN2        g898(.A(new_new_n831_), .B(new_new_n155_), .Y(new_new_n921_));
  NO4        g899(.A(new_new_n921_), .B(i_12_), .C(new_new_n596_), .D(new_new_n134_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n922_), .B(new_new_n209_), .Y(new_new_n923_));
  NA3        g901(.A(new_new_n101_), .B(new_new_n516_), .C(i_11_), .Y(new_new_n924_));
  NO2        g902(.A(new_new_n924_), .B(new_new_n157_), .Y(new_new_n925_));
  NA2        g903(.A(new_new_n859_), .B(new_new_n433_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n64_), .B(new_new_n104_), .Y(new_new_n927_));
  OAI220     g905(.A0(new_new_n927_), .A1(new_new_n917_), .B0(new_new_n926_), .B1(new_new_n626_), .Y(new_new_n928_));
  AOI210     g906(.A0(new_new_n928_), .A1(new_new_n847_), .B0(new_new_n925_), .Y(new_new_n929_));
  NA4        g907(.A(new_new_n929_), .B(new_new_n923_), .C(new_new_n920_), .D(new_new_n916_), .Y(new_new_n930_));
  NO4        g908(.A(new_new_n930_), .B(new_new_n912_), .C(new_new_n895_), .D(new_new_n890_), .Y(new_new_n931_));
  OAI210     g909(.A0(new_new_n765_), .A1(new_new_n758_), .B0(new_new_n37_), .Y(new_new_n932_));
  NA3        g910(.A(new_new_n853_), .B(new_new_n335_), .C(i_5_), .Y(new_new_n933_));
  NA3        g911(.A(new_new_n933_), .B(new_new_n932_), .C(new_new_n559_), .Y(new_new_n934_));
  NA2        g912(.A(new_new_n934_), .B(new_new_n200_), .Y(new_new_n935_));
  AN2        g913(.A(new_new_n646_), .B(new_new_n336_), .Y(new_new_n936_));
  NA2        g914(.A(new_new_n184_), .B(new_new_n186_), .Y(new_new_n937_));
  AO210      g915(.A0(new_new_n936_), .A1(new_new_n33_), .B0(new_new_n937_), .Y(new_new_n938_));
  NAi31      g916(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n939_));
  AOI210     g917(.A0(new_new_n120_), .A1(new_new_n70_), .B0(new_new_n939_), .Y(new_new_n940_));
  NO2        g918(.A(new_new_n940_), .B(new_new_n593_), .Y(new_new_n941_));
  NA2        g919(.A(new_new_n941_), .B(new_new_n938_), .Y(new_new_n942_));
  NO2        g920(.A(new_new_n427_), .B(new_new_n249_), .Y(new_new_n943_));
  NO2        g921(.A(new_new_n943_), .B(new_new_n823_), .Y(new_new_n944_));
  OAI210     g922(.A0(new_new_n924_), .A1(new_new_n151_), .B0(new_new_n944_), .Y(new_new_n945_));
  AOI210     g923(.A0(new_new_n942_), .A1(new_new_n48_), .B0(new_new_n945_), .Y(new_new_n946_));
  AOI210     g924(.A0(new_new_n946_), .A1(new_new_n935_), .B0(new_new_n73_), .Y(new_new_n947_));
  INV        g925(.A(new_new_n347_), .Y(new_new_n948_));
  NO2        g926(.A(new_new_n948_), .B(new_new_n705_), .Y(new_new_n949_));
  OAI210     g927(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n111_), .Y(new_new_n950_));
  NA2        g928(.A(new_new_n950_), .B(new_new_n76_), .Y(new_new_n951_));
  NA2        g929(.A(new_new_n899_), .B(new_new_n843_), .Y(new_new_n952_));
  AOI210     g930(.A0(new_new_n952_), .A1(new_new_n951_), .B0(new_new_n629_), .Y(new_new_n953_));
  INV        g931(.A(new_new_n953_), .Y(new_new_n954_));
  OAI210     g932(.A0(new_new_n251_), .A1(new_new_n159_), .B0(new_new_n89_), .Y(new_new_n955_));
  NO2        g933(.A(new_new_n955_), .B(i_11_), .Y(new_new_n956_));
  NA2        g934(.A(new_new_n554_), .B(new_new_n207_), .Y(new_new_n957_));
  OAI210     g935(.A0(new_new_n957_), .A1(new_new_n853_), .B0(new_new_n200_), .Y(new_new_n958_));
  NA2        g936(.A(new_new_n165_), .B(i_5_), .Y(new_new_n959_));
  NO2        g937(.A(new_new_n958_), .B(new_new_n959_), .Y(new_new_n960_));
  NO3        g938(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n961_));
  OAI210     g939(.A0(new_new_n861_), .A1(new_new_n287_), .B0(new_new_n961_), .Y(new_new_n962_));
  NO2        g940(.A(new_new_n962_), .B(new_new_n676_), .Y(new_new_n963_));
  INV        g941(.A(new_new_n509_), .Y(new_new_n964_));
  INV        g942(.A(new_new_n328_), .Y(new_new_n965_));
  AOI210     g943(.A0(new_new_n965_), .A1(new_new_n964_), .B0(new_new_n41_), .Y(new_new_n966_));
  NO4        g944(.A(new_new_n966_), .B(new_new_n963_), .C(new_new_n960_), .D(new_new_n956_), .Y(new_new_n967_));
  OAI210     g945(.A0(new_new_n954_), .A1(i_4_), .B0(new_new_n967_), .Y(new_new_n968_));
  NO3        g946(.A(new_new_n968_), .B(new_new_n949_), .C(new_new_n947_), .Y(new_new_n969_));
  NA4        g947(.A(new_new_n969_), .B(new_new_n931_), .C(new_new_n879_), .D(new_new_n813_), .Y(ori4));
  INV        g948(.A(new_new_n650_), .Y(new_new_n973_));
endmodule


