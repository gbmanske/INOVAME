//Benchmark atmr_intb_466_0.0156

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n374_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n433_, ori_ori_n434_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n378_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n384_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n445_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  NO3        o027(.A(ori_ori_n49_), .B(x11), .C(x09), .Y(ori_ori_n50_));
  INV        o028(.A(x09), .Y(ori_ori_n51_));
  NO2        o029(.A(x10), .B(x02), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x07), .Y(ori_ori_n54_));
  OAI210     o032(.A0(ori_ori_n54_), .A1(ori_ori_n50_), .B0(ori_ori_n47_), .Y(ori_ori_n55_));
  NOi21      o033(.An(x01), .B(x09), .Y(ori_ori_n56_));
  INV        o034(.A(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(ori_ori_n51_), .B(ori_ori_n57_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n56_), .Y(ori_ori_n59_));
  NA2        o037(.A(x09), .B(ori_ori_n57_), .Y(ori_ori_n60_));
  INV        o038(.A(x07), .Y(ori_ori_n61_));
  INV        o039(.A(ori_ori_n59_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n63_));
  NA2        o041(.A(ori_ori_n63_), .B(ori_ori_n24_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(ori_ori_n62_), .Y(ori_ori_n65_));
  NA2        o043(.A(ori_ori_n61_), .B(ori_ori_n48_), .Y(ori_ori_n66_));
  OAI210     o044(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n66_), .Y(ori_ori_n67_));
  AOI220     o045(.A0(ori_ori_n67_), .A1(ori_ori_n59_), .B0(ori_ori_n65_), .B1(ori_ori_n31_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(ori_ori_n68_), .A1(ori_ori_n55_), .B0(x05), .Y(ori_ori_n69_));
  NA2        o047(.A(x10), .B(x09), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n61_), .B(ori_ori_n23_), .Y(ori_ori_n71_));
  NA2        o049(.A(x09), .B(x05), .Y(ori_ori_n72_));
  NA2        o050(.A(x10), .B(x06), .Y(ori_ori_n73_));
  NA3        o051(.A(ori_ori_n73_), .B(ori_ori_n72_), .C(ori_ori_n28_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n71_), .B0(x03), .Y(ori_ori_n75_));
  NOi31      o053(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n76_));
  INV        o054(.A(x07), .Y(ori_ori_n77_));
  NO2        o055(.A(ori_ori_n77_), .B(ori_ori_n24_), .Y(ori_ori_n78_));
  NO2        o056(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n36_), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n79_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n81_));
  AOI210     o059(.A0(ori_ori_n80_), .A1(ori_ori_n48_), .B0(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o060(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n83_));
  NO2        o061(.A(x08), .B(x01), .Y(ori_ori_n84_));
  OAI210     o062(.A0(ori_ori_n84_), .A1(ori_ori_n83_), .B0(ori_ori_n35_), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n86_));
  NO3        o064(.A(ori_ori_n85_), .B(ori_ori_n82_), .C(ori_ori_n78_), .Y(ori_ori_n87_));
  AN2        o065(.A(ori_ori_n87_), .B(ori_ori_n75_), .Y(ori_ori_n88_));
  INV        o066(.A(ori_ori_n85_), .Y(ori_ori_n89_));
  NO2        o067(.A(x06), .B(x05), .Y(ori_ori_n90_));
  NA2        o068(.A(x11), .B(x00), .Y(ori_ori_n91_));
  NO2        o069(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n92_));
  NOi21      o070(.An(ori_ori_n91_), .B(ori_ori_n92_), .Y(ori_ori_n93_));
  AOI210     o071(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NOi21      o072(.An(x01), .B(x10), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n29_), .B(ori_ori_n57_), .Y(ori_ori_n96_));
  NO3        o074(.A(ori_ori_n96_), .B(ori_ori_n95_), .C(x06), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n97_), .B(ori_ori_n27_), .Y(ori_ori_n98_));
  OAI210     o076(.A0(ori_ori_n94_), .A1(x07), .B0(ori_ori_n98_), .Y(ori_ori_n99_));
  NO3        o077(.A(ori_ori_n99_), .B(ori_ori_n88_), .C(ori_ori_n69_), .Y(ori01));
  INV        o078(.A(x12), .Y(ori_ori_n101_));
  INV        o079(.A(x13), .Y(ori_ori_n102_));
  NA2        o080(.A(x08), .B(x04), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n95_), .B(ori_ori_n28_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(ori_ori_n72_), .Y(ori_ori_n105_));
  NO2        o083(.A(x10), .B(x01), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n107_), .B(ori_ori_n106_), .Y(ori_ori_n108_));
  NA2        o086(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n109_));
  NO3        o087(.A(ori_ori_n109_), .B(ori_ori_n36_), .C(ori_ori_n41_), .Y(ori_ori_n110_));
  AOI210     o088(.A0(ori_ori_n110_), .A1(ori_ori_n108_), .B0(ori_ori_n105_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n111_), .B(ori_ori_n102_), .Y(ori_ori_n112_));
  NO2        o090(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n113_));
  NOi21      o091(.An(ori_ori_n113_), .B(ori_ori_n58_), .Y(ori_ori_n114_));
  NO2        o092(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n115_));
  NA3        o093(.A(x13), .B(ori_ori_n115_), .C(x06), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n114_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n84_), .B(x13), .Y(ori_ori_n118_));
  NA2        o096(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NA2        o098(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n121_), .B(x05), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n122_), .B(ori_ori_n120_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n35_), .B(ori_ori_n57_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n124_), .B(ori_ori_n102_), .Y(ori_ori_n125_));
  AOI210     o103(.A0(ori_ori_n125_), .A1(ori_ori_n80_), .B0(ori_ori_n114_), .Y(ori_ori_n126_));
  AOI210     o104(.A0(ori_ori_n126_), .A1(ori_ori_n123_), .B0(ori_ori_n73_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n128_));
  NA2        o106(.A(x10), .B(ori_ori_n57_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(ori_ori_n128_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n51_), .B(x05), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n132_));
  NA3        o110(.A(ori_ori_n132_), .B(ori_ori_n131_), .C(x13), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n60_), .B(x05), .Y(ori_ori_n134_));
  NOi31      o112(.An(ori_ori_n133_), .B(ori_ori_n134_), .C(ori_ori_n130_), .Y(ori_ori_n135_));
  NO3        o113(.A(ori_ori_n135_), .B(x06), .C(x03), .Y(ori_ori_n136_));
  NO4        o114(.A(ori_ori_n136_), .B(ori_ori_n127_), .C(ori_ori_n117_), .D(ori_ori_n112_), .Y(ori_ori_n137_));
  NA2        o115(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n138_));
  OAI210     o116(.A0(ori_ori_n84_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n139_), .B(ori_ori_n138_), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n142_));
  AOI210     o120(.A0(ori_ori_n142_), .A1(ori_ori_n49_), .B0(ori_ori_n141_), .Y(ori_ori_n143_));
  AN2        o121(.A(ori_ori_n143_), .B(ori_ori_n140_), .Y(ori_ori_n144_));
  NO2        o122(.A(x09), .B(x05), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n145_), .B(ori_ori_n47_), .Y(ori_ori_n146_));
  AOI210     o124(.A0(ori_ori_n146_), .A1(ori_ori_n108_), .B0(ori_ori_n49_), .Y(ori_ori_n147_));
  NA2        o125(.A(x09), .B(x00), .Y(ori_ori_n148_));
  NA2        o126(.A(ori_ori_n113_), .B(ori_ori_n148_), .Y(ori_ori_n149_));
  NA2        o127(.A(ori_ori_n76_), .B(ori_ori_n51_), .Y(ori_ori_n150_));
  AOI210     o128(.A0(ori_ori_n150_), .A1(ori_ori_n149_), .B0(ori_ori_n142_), .Y(ori_ori_n151_));
  NO3        o129(.A(ori_ori_n151_), .B(ori_ori_n147_), .C(ori_ori_n144_), .Y(ori_ori_n152_));
  NO2        o130(.A(x03), .B(x02), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n85_), .B(ori_ori_n102_), .Y(ori_ori_n154_));
  OAI210     o132(.A0(ori_ori_n154_), .A1(ori_ori_n114_), .B0(ori_ori_n153_), .Y(ori_ori_n155_));
  OA210      o133(.A0(ori_ori_n152_), .A1(x11), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  OAI210     o134(.A0(ori_ori_n137_), .A1(ori_ori_n23_), .B0(ori_ori_n156_), .Y(ori_ori_n157_));
  NA2        o135(.A(ori_ori_n108_), .B(ori_ori_n40_), .Y(ori_ori_n158_));
  NAi21      o136(.An(x06), .B(x10), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n158_), .B(ori_ori_n41_), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n102_), .B(x01), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n162_), .B(x08), .Y(ori_ori_n163_));
  OAI210     o141(.A0(x05), .A1(ori_ori_n163_), .B0(ori_ori_n51_), .Y(ori_ori_n164_));
  AOI210     o142(.A0(ori_ori_n164_), .A1(ori_ori_n161_), .B0(ori_ori_n48_), .Y(ori_ori_n165_));
  AOI210     o143(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n166_));
  OAI210     o144(.A0(ori_ori_n165_), .A1(ori_ori_n160_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  NA2        o145(.A(x04), .B(x02), .Y(ori_ori_n168_));
  NA2        o146(.A(x10), .B(x05), .Y(ori_ori_n169_));
  NO2        o147(.A(x09), .B(x01), .Y(ori_ori_n170_));
  NO3        o148(.A(ori_ori_n170_), .B(ori_ori_n106_), .C(ori_ori_n31_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(x00), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n113_), .B(x08), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n95_), .B(x05), .Y(ori_ori_n174_));
  INV        o152(.A(ori_ori_n174_), .Y(ori_ori_n175_));
  AOI210     o153(.A0(ori_ori_n173_), .A1(x06), .B0(ori_ori_n175_), .Y(ori_ori_n176_));
  OAI210     o154(.A0(ori_ori_n176_), .A1(x11), .B0(ori_ori_n172_), .Y(ori_ori_n177_));
  NAi21      o155(.An(ori_ori_n168_), .B(ori_ori_n177_), .Y(ori_ori_n178_));
  INV        o156(.A(ori_ori_n25_), .Y(ori_ori_n179_));
  NAi21      o157(.An(x13), .B(x00), .Y(ori_ori_n180_));
  AOI210     o158(.A0(ori_ori_n29_), .A1(ori_ori_n48_), .B0(ori_ori_n180_), .Y(ori_ori_n181_));
  AOI220     o159(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(ori_ori_n182_));
  OAI210     o160(.A0(ori_ori_n169_), .A1(ori_ori_n35_), .B0(ori_ori_n182_), .Y(ori_ori_n183_));
  AN2        o161(.A(ori_ori_n183_), .B(ori_ori_n181_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n96_), .B(x06), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n180_), .B(ori_ori_n36_), .Y(ori_ori_n186_));
  INV        o164(.A(ori_ori_n186_), .Y(ori_ori_n187_));
  OAI210     o165(.A0(ori_ori_n433_), .A1(ori_ori_n184_), .B0(ori_ori_n179_), .Y(ori_ori_n188_));
  NOi21      o166(.An(x09), .B(x00), .Y(ori_ori_n189_));
  NO3        o167(.A(ori_ori_n83_), .B(ori_ori_n189_), .C(ori_ori_n47_), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n190_), .B(ori_ori_n129_), .Y(ori_ori_n191_));
  NA2        o169(.A(x10), .B(x08), .Y(ori_ori_n192_));
  INV        o170(.A(ori_ori_n192_), .Y(ori_ori_n193_));
  NA2        o171(.A(x06), .B(x05), .Y(ori_ori_n194_));
  OAI210     o172(.A0(ori_ori_n194_), .A1(ori_ori_n35_), .B0(ori_ori_n101_), .Y(ori_ori_n195_));
  AOI210     o173(.A0(ori_ori_n193_), .A1(ori_ori_n58_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n196_), .B(ori_ori_n191_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n102_), .B(x12), .Y(ori_ori_n198_));
  AOI210     o176(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n198_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n95_), .B(ori_ori_n51_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n201_));
  NA2        o179(.A(ori_ori_n201_), .B(x02), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n202_), .B(ori_ori_n200_), .Y(ori_ori_n203_));
  AOI210     o181(.A0(ori_ori_n199_), .A1(ori_ori_n197_), .B0(ori_ori_n203_), .Y(ori_ori_n204_));
  NA4        o182(.A(ori_ori_n204_), .B(ori_ori_n188_), .C(ori_ori_n178_), .D(ori_ori_n167_), .Y(ori_ori_n205_));
  AOI210     o183(.A0(ori_ori_n157_), .A1(ori_ori_n101_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  INV        o184(.A(ori_ori_n74_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n207_), .B(ori_ori_n140_), .Y(ori_ori_n208_));
  NA2        o186(.A(ori_ori_n51_), .B(ori_ori_n47_), .Y(ori_ori_n209_));
  NA2        o187(.A(ori_ori_n209_), .B(ori_ori_n139_), .Y(ori_ori_n210_));
  AOI210     o188(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n128_), .B(x06), .Y(ori_ori_n212_));
  AOI210     o190(.A0(ori_ori_n211_), .A1(ori_ori_n210_), .B0(ori_ori_n212_), .Y(ori_ori_n213_));
  AOI210     o191(.A0(ori_ori_n213_), .A1(ori_ori_n208_), .B0(x12), .Y(ori_ori_n214_));
  INV        o192(.A(ori_ori_n76_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n95_), .B(x06), .Y(ori_ori_n216_));
  AOI210     o194(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n51_), .Y(ori_ori_n217_));
  NO3        o195(.A(ori_ori_n217_), .B(ori_ori_n216_), .C(ori_ori_n41_), .Y(ori_ori_n218_));
  NA4        o196(.A(ori_ori_n159_), .B(ori_ori_n56_), .C(ori_ori_n36_), .D(x04), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n219_), .B(ori_ori_n142_), .Y(ori_ori_n220_));
  OAI210     o198(.A0(ori_ori_n220_), .A1(ori_ori_n218_), .B0(x02), .Y(ori_ori_n221_));
  AOI210     o199(.A0(ori_ori_n221_), .A1(ori_ori_n57_), .B0(ori_ori_n23_), .Y(ori_ori_n222_));
  OAI210     o200(.A0(ori_ori_n214_), .A1(ori_ori_n57_), .B0(ori_ori_n222_), .Y(ori_ori_n223_));
  INV        o201(.A(ori_ori_n142_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n51_), .B(x03), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n79_), .A1(ori_ori_n36_), .B0(ori_ori_n119_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n102_), .B(x03), .Y(ori_ori_n227_));
  AOI220     o205(.A0(ori_ori_n227_), .A1(ori_ori_n226_), .B0(ori_ori_n76_), .B1(ori_ori_n225_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n229_));
  INV        o207(.A(ori_ori_n159_), .Y(ori_ori_n230_));
  NOi21      o208(.An(x13), .B(x04), .Y(ori_ori_n231_));
  NO3        o209(.A(ori_ori_n231_), .B(ori_ori_n76_), .C(ori_ori_n189_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n232_), .B(x05), .Y(ori_ori_n233_));
  AOI220     o211(.A0(ori_ori_n233_), .A1(ori_ori_n229_), .B0(ori_ori_n230_), .B1(ori_ori_n57_), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n228_), .A1(ori_ori_n224_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  INV        o213(.A(ori_ori_n92_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(x12), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n51_), .B(ori_ori_n36_), .Y(ori_ori_n239_));
  OAI210     o217(.A0(ori_ori_n239_), .A1(ori_ori_n183_), .B0(ori_ori_n181_), .Y(ori_ori_n240_));
  AOI210     o218(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n241_));
  NO2        o219(.A(x06), .B(x00), .Y(ori_ori_n242_));
  NO3        o220(.A(ori_ori_n242_), .B(ori_ori_n241_), .C(ori_ori_n41_), .Y(ori_ori_n243_));
  OAI210     o221(.A0(ori_ori_n103_), .A1(ori_ori_n148_), .B0(ori_ori_n73_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(ori_ori_n243_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(x03), .Y(ori_ori_n247_));
  OA210      o225(.A0(ori_ori_n247_), .A1(ori_ori_n245_), .B0(ori_ori_n240_), .Y(ori_ori_n248_));
  NA2        o226(.A(x13), .B(ori_ori_n101_), .Y(ori_ori_n249_));
  NA3        o227(.A(ori_ori_n249_), .B(ori_ori_n195_), .C(ori_ori_n93_), .Y(ori_ori_n250_));
  OAI210     o228(.A0(ori_ori_n248_), .A1(ori_ori_n238_), .B0(ori_ori_n250_), .Y(ori_ori_n251_));
  AOI210     o229(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(ori_ori_n251_), .Y(ori_ori_n252_));
  AOI210     o230(.A0(ori_ori_n252_), .A1(ori_ori_n223_), .B0(x07), .Y(ori_ori_n253_));
  NA2        o231(.A(ori_ori_n72_), .B(ori_ori_n29_), .Y(ori_ori_n254_));
  NOi31      o232(.An(ori_ori_n138_), .B(ori_ori_n231_), .C(ori_ori_n189_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n255_), .B(ori_ori_n254_), .Y(ori_ori_n256_));
  NO2        o234(.A(x08), .B(x05), .Y(ori_ori_n257_));
  INV        o235(.A(ori_ori_n241_), .Y(ori_ori_n258_));
  NA2        o236(.A(x13), .B(ori_ori_n31_), .Y(ori_ori_n259_));
  INV        o237(.A(ori_ori_n259_), .Y(ori_ori_n260_));
  NO2        o238(.A(x12), .B(x02), .Y(ori_ori_n261_));
  INV        o239(.A(ori_ori_n261_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n236_), .Y(ori_ori_n263_));
  OA210      o241(.A0(ori_ori_n260_), .A1(ori_ori_n256_), .B0(ori_ori_n263_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n51_), .B(ori_ori_n41_), .Y(ori_ori_n265_));
  NO2        o243(.A(ori_ori_n265_), .B(x01), .Y(ori_ori_n266_));
  INV        o244(.A(ori_ori_n266_), .Y(ori_ori_n267_));
  AOI210     o245(.A0(ori_ori_n267_), .A1(ori_ori_n133_), .B0(ori_ori_n29_), .Y(ori_ori_n268_));
  NA2        o246(.A(ori_ori_n102_), .B(x04), .Y(ori_ori_n269_));
  NA2        o247(.A(ori_ori_n269_), .B(ori_ori_n28_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n270_), .B(ori_ori_n118_), .Y(ori_ori_n271_));
  NO3        o249(.A(ori_ori_n91_), .B(x12), .C(x03), .Y(ori_ori_n272_));
  OAI210     o250(.A0(ori_ori_n271_), .A1(ori_ori_n268_), .B0(ori_ori_n272_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n200_), .A1(ori_ori_n194_), .B0(ori_ori_n103_), .Y(ori_ori_n274_));
  NOi21      o252(.An(ori_ori_n254_), .B(ori_ori_n216_), .Y(ori_ori_n275_));
  NO2        o253(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n276_));
  OAI210     o254(.A0(ori_ori_n275_), .A1(ori_ori_n274_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  NO2        o255(.A(ori_ori_n58_), .B(x05), .Y(ori_ori_n278_));
  NO3        o256(.A(ori_ori_n278_), .B(ori_ori_n217_), .C(ori_ori_n185_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n238_), .B(ori_ori_n28_), .Y(ori_ori_n280_));
  OAI210     o258(.A0(ori_ori_n279_), .A1(ori_ori_n224_), .B0(ori_ori_n280_), .Y(ori_ori_n281_));
  NA3        o259(.A(ori_ori_n281_), .B(ori_ori_n277_), .C(ori_ori_n273_), .Y(ori_ori_n282_));
  NO3        o260(.A(ori_ori_n282_), .B(ori_ori_n264_), .C(ori_ori_n253_), .Y(ori_ori_n283_));
  OAI210     o261(.A0(ori_ori_n206_), .A1(ori_ori_n61_), .B0(ori_ori_n283_), .Y(ori02));
  AOI210     o262(.A0(ori_ori_n138_), .A1(ori_ori_n85_), .B0(ori_ori_n131_), .Y(ori_ori_n285_));
  NOi21      o263(.An(ori_ori_n232_), .B(ori_ori_n170_), .Y(ori_ori_n286_));
  NO2        o264(.A(ori_ori_n102_), .B(ori_ori_n35_), .Y(ori_ori_n287_));
  NA3        o265(.A(ori_ori_n287_), .B(ori_ori_n193_), .C(ori_ori_n56_), .Y(ori_ori_n288_));
  OAI210     o266(.A0(ori_ori_n286_), .A1(ori_ori_n32_), .B0(ori_ori_n288_), .Y(ori_ori_n289_));
  OAI210     o267(.A0(ori_ori_n289_), .A1(ori_ori_n285_), .B0(ori_ori_n169_), .Y(ori_ori_n290_));
  INV        o268(.A(ori_ori_n169_), .Y(ori_ori_n291_));
  AOI210     o269(.A0(ori_ori_n115_), .A1(ori_ori_n86_), .B0(ori_ori_n217_), .Y(ori_ori_n292_));
  OAI220     o270(.A0(ori_ori_n292_), .A1(ori_ori_n102_), .B0(ori_ori_n85_), .B1(ori_ori_n51_), .Y(ori_ori_n293_));
  AOI220     o271(.A0(ori_ori_n293_), .A1(ori_ori_n291_), .B0(ori_ori_n154_), .B1(ori_ori_n153_), .Y(ori_ori_n294_));
  AOI210     o272(.A0(ori_ori_n294_), .A1(ori_ori_n290_), .B0(ori_ori_n48_), .Y(ori_ori_n295_));
  NO2        o273(.A(x05), .B(x02), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n210_), .A1(ori_ori_n189_), .B0(ori_ori_n296_), .Y(ori_ori_n297_));
  AOI220     o275(.A0(ori_ori_n257_), .A1(ori_ori_n58_), .B0(ori_ori_n56_), .B1(ori_ori_n36_), .Y(ori_ori_n298_));
  NOi21      o276(.An(ori_ori_n287_), .B(ori_ori_n298_), .Y(ori_ori_n299_));
  INV        o277(.A(ori_ori_n299_), .Y(ori_ori_n300_));
  AOI210     o278(.A0(ori_ori_n300_), .A1(ori_ori_n297_), .B0(ori_ori_n142_), .Y(ori_ori_n301_));
  NAi21      o279(.An(ori_ori_n233_), .B(ori_ori_n228_), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n246_), .B(ori_ori_n47_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n303_), .B(ori_ori_n302_), .Y(ori_ori_n304_));
  AN2        o282(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n305_));
  OAI210     o283(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n306_));
  NA2        o284(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n307_));
  OA210      o285(.A0(ori_ori_n307_), .A1(x08), .B0(ori_ori_n146_), .Y(ori_ori_n308_));
  AOI210     o286(.A0(ori_ori_n308_), .A1(ori_ori_n139_), .B0(ori_ori_n306_), .Y(ori_ori_n309_));
  OAI210     o287(.A0(ori_ori_n309_), .A1(ori_ori_n305_), .B0(ori_ori_n96_), .Y(ori_ori_n310_));
  INV        o288(.A(ori_ori_n153_), .Y(ori_ori_n311_));
  OAI220     o289(.A0(ori_ori_n258_), .A1(ori_ori_n104_), .B0(ori_ori_n311_), .B1(ori_ori_n130_), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n312_), .B(x13), .Y(ori_ori_n313_));
  NA3        o291(.A(ori_ori_n313_), .B(ori_ori_n310_), .C(ori_ori_n304_), .Y(ori_ori_n314_));
  NO3        o292(.A(ori_ori_n314_), .B(ori_ori_n301_), .C(ori_ori_n295_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n141_), .B(x03), .Y(ori_ori_n316_));
  INV        o294(.A(ori_ori_n180_), .Y(ori_ori_n317_));
  AOI220     o295(.A0(x08), .A1(ori_ori_n317_), .B0(ori_ori_n201_), .B1(x08), .Y(ori_ori_n318_));
  OAI210     o296(.A0(ori_ori_n318_), .A1(ori_ori_n278_), .B0(ori_ori_n316_), .Y(ori_ori_n319_));
  NA2        o297(.A(ori_ori_n319_), .B(ori_ori_n106_), .Y(ori_ori_n320_));
  NA2        o298(.A(ori_ori_n168_), .B(ori_ori_n162_), .Y(ori_ori_n321_));
  AN2        o299(.A(ori_ori_n321_), .B(ori_ori_n173_), .Y(ori_ori_n322_));
  INV        o300(.A(ori_ori_n56_), .Y(ori_ori_n323_));
  OAI220     o301(.A0(ori_ori_n269_), .A1(ori_ori_n323_), .B0(ori_ori_n131_), .B1(ori_ori_n28_), .Y(ori_ori_n324_));
  OAI210     o302(.A0(ori_ori_n324_), .A1(ori_ori_n322_), .B0(ori_ori_n107_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n269_), .B(ori_ori_n101_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n101_), .B(ori_ori_n41_), .Y(ori_ori_n327_));
  NA3        o305(.A(ori_ori_n327_), .B(ori_ori_n326_), .C(ori_ori_n130_), .Y(ori_ori_n328_));
  NA4        o306(.A(ori_ori_n328_), .B(ori_ori_n325_), .C(ori_ori_n320_), .D(ori_ori_n48_), .Y(ori_ori_n329_));
  INV        o307(.A(ori_ori_n201_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n331_));
  OAI220     o309(.A0(ori_ori_n331_), .A1(ori_ori_n434_), .B0(ori_ori_n330_), .B1(ori_ori_n59_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n332_), .B(x02), .Y(ori_ori_n333_));
  INV        o311(.A(ori_ori_n239_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n198_), .B(x04), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n335_), .B(ori_ori_n334_), .Y(ori_ori_n336_));
  NO3        o314(.A(ori_ori_n182_), .B(x13), .C(ori_ori_n31_), .Y(ori_ori_n337_));
  OAI210     o315(.A0(ori_ori_n337_), .A1(ori_ori_n336_), .B0(ori_ori_n96_), .Y(ori_ori_n338_));
  NO3        o316(.A(ori_ori_n198_), .B(ori_ori_n161_), .C(ori_ori_n52_), .Y(ori_ori_n339_));
  OAI210     o317(.A0(ori_ori_n148_), .A1(ori_ori_n36_), .B0(ori_ori_n101_), .Y(ori_ori_n340_));
  OAI210     o318(.A0(ori_ori_n340_), .A1(ori_ori_n190_), .B0(ori_ori_n339_), .Y(ori_ori_n341_));
  NA4        o319(.A(ori_ori_n341_), .B(ori_ori_n338_), .C(ori_ori_n333_), .D(x06), .Y(ori_ori_n342_));
  NA2        o320(.A(x09), .B(x03), .Y(ori_ori_n343_));
  OAI220     o321(.A0(ori_ori_n343_), .A1(ori_ori_n129_), .B0(ori_ori_n209_), .B1(ori_ori_n63_), .Y(ori_ori_n344_));
  NO3        o322(.A(ori_ori_n278_), .B(ori_ori_n128_), .C(x08), .Y(ori_ori_n345_));
  INV        o323(.A(ori_ori_n345_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n347_));
  NO3        o325(.A(ori_ori_n113_), .B(ori_ori_n129_), .C(ori_ori_n38_), .Y(ori_ori_n348_));
  AOI210     o326(.A0(ori_ori_n339_), .A1(ori_ori_n347_), .B0(ori_ori_n348_), .Y(ori_ori_n349_));
  OAI210     o327(.A0(ori_ori_n346_), .A1(ori_ori_n28_), .B0(ori_ori_n349_), .Y(ori_ori_n350_));
  AO220      o328(.A0(ori_ori_n350_), .A1(x04), .B0(ori_ori_n344_), .B1(x05), .Y(ori_ori_n351_));
  AOI210     o329(.A0(ori_ori_n342_), .A1(ori_ori_n329_), .B0(ori_ori_n351_), .Y(ori_ori_n352_));
  OAI210     o330(.A0(ori_ori_n315_), .A1(x12), .B0(ori_ori_n352_), .Y(ori03));
  OR2        o331(.A(ori_ori_n42_), .B(ori_ori_n225_), .Y(ori_ori_n354_));
  AOI210     o332(.A0(ori_ori_n154_), .A1(ori_ori_n101_), .B0(ori_ori_n354_), .Y(ori_ori_n355_));
  AO210      o333(.A0(ori_ori_n334_), .A1(ori_ori_n86_), .B0(ori_ori_n335_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n198_), .B(ori_ori_n153_), .Y(ori_ori_n357_));
  NA3        o335(.A(ori_ori_n357_), .B(ori_ori_n356_), .C(ori_ori_n202_), .Y(ori_ori_n358_));
  OAI210     o336(.A0(ori_ori_n358_), .A1(ori_ori_n355_), .B0(x05), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n354_), .B(x05), .Y(ori_ori_n360_));
  AOI210     o338(.A0(ori_ori_n139_), .A1(ori_ori_n215_), .B0(ori_ori_n360_), .Y(ori_ori_n361_));
  AOI210     o339(.A0(ori_ori_n227_), .A1(ori_ori_n80_), .B0(ori_ori_n122_), .Y(ori_ori_n362_));
  OAI220     o340(.A0(ori_ori_n362_), .A1(ori_ori_n59_), .B0(ori_ori_n307_), .B1(ori_ori_n298_), .Y(ori_ori_n363_));
  OAI210     o341(.A0(ori_ori_n363_), .A1(ori_ori_n361_), .B0(ori_ori_n101_), .Y(ori_ori_n364_));
  AOI210     o342(.A0(ori_ori_n146_), .A1(ori_ori_n60_), .B0(ori_ori_n38_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n170_), .B(ori_ori_n134_), .Y(ori_ori_n366_));
  OAI220     o344(.A0(ori_ori_n366_), .A1(ori_ori_n37_), .B0(ori_ori_n149_), .B1(x13), .Y(ori_ori_n367_));
  OAI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n365_), .B0(x04), .Y(ori_ori_n368_));
  NO3        o346(.A(ori_ori_n327_), .B(ori_ori_n85_), .C(ori_ori_n59_), .Y(ori_ori_n369_));
  AOI210     o347(.A0(ori_ori_n187_), .A1(ori_ori_n101_), .B0(ori_ori_n146_), .Y(ori_ori_n370_));
  OA210      o348(.A0(ori_ori_n163_), .A1(x12), .B0(ori_ori_n134_), .Y(ori_ori_n371_));
  NO3        o349(.A(ori_ori_n371_), .B(ori_ori_n370_), .C(ori_ori_n369_), .Y(ori_ori_n372_));
  NA4        o350(.A(ori_ori_n372_), .B(ori_ori_n368_), .C(ori_ori_n364_), .D(ori_ori_n359_), .Y(ori04));
  NO2        o351(.A(ori_ori_n89_), .B(ori_ori_n39_), .Y(ori_ori_n374_));
  XO2        o352(.A(ori_ori_n374_), .B(ori_ori_n249_), .Y(ori05));
  NO2        o353(.A(ori_ori_n306_), .B(ori_ori_n25_), .Y(ori_ori_n376_));
  NA3        o354(.A(ori_ori_n142_), .B(ori_ori_n131_), .C(ori_ori_n31_), .Y(ori_ori_n377_));
  AOI210     o355(.A0(ori_ori_n230_), .A1(ori_ori_n57_), .B0(ori_ori_n90_), .Y(ori_ori_n378_));
  AOI210     o356(.A0(ori_ori_n378_), .A1(ori_ori_n377_), .B0(ori_ori_n24_), .Y(ori_ori_n379_));
  OAI210     o357(.A0(ori_ori_n379_), .A1(ori_ori_n376_), .B0(ori_ori_n101_), .Y(ori_ori_n380_));
  NA2        o358(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n381_));
  NA2        o359(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n254_), .B(x03), .Y(ori_ori_n383_));
  OAI220     o361(.A0(ori_ori_n383_), .A1(ori_ori_n382_), .B0(ori_ori_n381_), .B1(ori_ori_n81_), .Y(ori_ori_n384_));
  OAI210     o362(.A0(ori_ori_n26_), .A1(ori_ori_n101_), .B0(x07), .Y(ori_ori_n385_));
  AOI210     o363(.A0(ori_ori_n384_), .A1(x06), .B0(ori_ori_n385_), .Y(ori_ori_n386_));
  AOI210     o364(.A0(ori_ori_n81_), .A1(ori_ori_n31_), .B0(ori_ori_n52_), .Y(ori_ori_n387_));
  NO3        o365(.A(ori_ori_n387_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n388_));
  NA2        o366(.A(ori_ori_n70_), .B(x02), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n389_), .B(ori_ori_n383_), .Y(ori_ori_n390_));
  OR2        o368(.A(ori_ori_n390_), .B(ori_ori_n238_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n242_), .B(ori_ori_n236_), .Y(ori_ori_n392_));
  OAI210     o370(.A0(x11), .A1(ori_ori_n29_), .B0(ori_ori_n48_), .Y(ori_ori_n393_));
  OR2        o371(.A(ori_ori_n393_), .B(ori_ori_n44_), .Y(ori_ori_n394_));
  NA3        o372(.A(ori_ori_n394_), .B(ori_ori_n392_), .C(ori_ori_n391_), .Y(ori_ori_n395_));
  OAI210     o373(.A0(ori_ori_n395_), .A1(ori_ori_n388_), .B0(ori_ori_n101_), .Y(ori_ori_n396_));
  NA2        o374(.A(ori_ori_n33_), .B(ori_ori_n101_), .Y(ori_ori_n397_));
  AOI210     o375(.A0(ori_ori_n397_), .A1(ori_ori_n92_), .B0(x07), .Y(ori_ori_n398_));
  AOI220     o376(.A0(ori_ori_n398_), .A1(ori_ori_n396_), .B0(ori_ori_n386_), .B1(ori_ori_n380_), .Y(ori_ori_n399_));
  OR2        o377(.A(ori_ori_n265_), .B(ori_ori_n262_), .Y(ori_ori_n400_));
  NO2        o378(.A(ori_ori_n145_), .B(ori_ori_n28_), .Y(ori_ori_n401_));
  AOI210     o379(.A0(ori_ori_n400_), .A1(ori_ori_n47_), .B0(ori_ori_n401_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n402_), .B(ori_ori_n102_), .Y(ori_ori_n403_));
  AOI210     o381(.A0(ori_ori_n335_), .A1(ori_ori_n109_), .B0(ori_ori_n261_), .Y(ori_ori_n404_));
  NOi21      o382(.An(ori_ori_n316_), .B(ori_ori_n134_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n405_), .B(ori_ori_n262_), .Y(ori_ori_n406_));
  OAI210     o384(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n407_));
  AOI210     o385(.A0(ori_ori_n249_), .A1(ori_ori_n47_), .B0(ori_ori_n407_), .Y(ori_ori_n408_));
  NO4        o386(.A(ori_ori_n408_), .B(ori_ori_n406_), .C(ori_ori_n404_), .D(x08), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n131_), .B(ori_ori_n28_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n410_), .B(ori_ori_n266_), .Y(ori_ori_n411_));
  OR3        o389(.A(ori_ori_n411_), .B(x12), .C(x03), .Y(ori_ori_n412_));
  NA3        o390(.A(ori_ori_n330_), .B(ori_ori_n124_), .C(x12), .Y(ori_ori_n413_));
  AO210      o391(.A0(ori_ori_n330_), .A1(ori_ori_n124_), .B0(ori_ori_n249_), .Y(ori_ori_n414_));
  NA4        o392(.A(ori_ori_n414_), .B(ori_ori_n413_), .C(ori_ori_n412_), .D(x08), .Y(ori_ori_n415_));
  INV        o393(.A(ori_ori_n415_), .Y(ori_ori_n416_));
  AOI210     o394(.A0(ori_ori_n409_), .A1(ori_ori_n403_), .B0(ori_ori_n416_), .Y(ori_ori_n417_));
  INV        o395(.A(x03), .Y(ori_ori_n418_));
  NO2        o396(.A(ori_ori_n145_), .B(ori_ori_n43_), .Y(ori_ori_n419_));
  OAI210     o397(.A0(ori_ori_n419_), .A1(ori_ori_n418_), .B0(ori_ori_n186_), .Y(ori_ori_n420_));
  NA3        o398(.A(ori_ori_n411_), .B(ori_ori_n405_), .C(ori_ori_n326_), .Y(ori_ori_n421_));
  NA3        o399(.A(x14), .B(ori_ori_n421_), .C(ori_ori_n420_), .Y(ori_ori_n422_));
  AOI220     o400(.A0(ori_ori_n397_), .A1(ori_ori_n61_), .B0(ori_ori_n410_), .B1(ori_ori_n161_), .Y(ori_ori_n423_));
  NOi21      o401(.An(ori_ori_n269_), .B(ori_ori_n149_), .Y(ori_ori_n424_));
  NO3        o402(.A(ori_ori_n128_), .B(ori_ori_n24_), .C(x06), .Y(ori_ori_n425_));
  AOI210     o403(.A0(ori_ori_n276_), .A1(ori_ori_n230_), .B0(ori_ori_n425_), .Y(ori_ori_n426_));
  OAI210     o404(.A0(ori_ori_n44_), .A1(x04), .B0(ori_ori_n426_), .Y(ori_ori_n427_));
  OAI210     o405(.A0(ori_ori_n427_), .A1(ori_ori_n424_), .B0(ori_ori_n101_), .Y(ori_ori_n428_));
  OAI210     o406(.A0(ori_ori_n423_), .A1(ori_ori_n91_), .B0(ori_ori_n428_), .Y(ori_ori_n429_));
  NO4        o407(.A(ori_ori_n429_), .B(ori_ori_n422_), .C(ori_ori_n417_), .D(ori_ori_n399_), .Y(ori06));
  INV        o408(.A(ori_ori_n73_), .Y(ori_ori_n433_));
  INV        o409(.A(ori_ori_n40_), .Y(ori_ori_n434_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x10), .B(x09), .Y(mai_mai_n71_));
  NO2        m049(.A(mai_mai_n61_), .B(mai_mai_n23_), .Y(mai_mai_n72_));
  NA2        m050(.A(x09), .B(x05), .Y(mai_mai_n73_));
  NA2        m051(.A(x10), .B(x06), .Y(mai_mai_n74_));
  NA3        m052(.A(mai_mai_n74_), .B(mai_mai_n73_), .C(mai_mai_n28_), .Y(mai_mai_n75_));
  NO2        m053(.A(mai_mai_n61_), .B(mai_mai_n41_), .Y(mai_mai_n76_));
  OAI210     m054(.A0(mai_mai_n75_), .A1(mai_mai_n72_), .B0(x03), .Y(mai_mai_n77_));
  NOi31      m055(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n78_));
  NO2        m056(.A(x10), .B(x09), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n447_), .B(mai_mai_n24_), .Y(mai_mai_n80_));
  NO2        m058(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n81_));
  NO2        m059(.A(mai_mai_n81_), .B(mai_mai_n36_), .Y(mai_mai_n82_));
  OAI210     m060(.A0(mai_mai_n81_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n83_));
  AOI210     m061(.A0(mai_mai_n82_), .A1(mai_mai_n48_), .B0(mai_mai_n83_), .Y(mai_mai_n84_));
  NO2        m062(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n85_));
  NO2        m063(.A(x08), .B(x01), .Y(mai_mai_n86_));
  OAI210     m064(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n35_), .Y(mai_mai_n87_));
  NA2        m065(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n88_));
  NO3        m066(.A(mai_mai_n87_), .B(mai_mai_n84_), .C(mai_mai_n80_), .Y(mai_mai_n89_));
  AN2        m067(.A(mai_mai_n89_), .B(mai_mai_n77_), .Y(mai_mai_n90_));
  INV        m068(.A(mai_mai_n87_), .Y(mai_mai_n91_));
  NA2        m069(.A(x11), .B(x00), .Y(mai_mai_n92_));
  NO2        m070(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n93_));
  NOi21      m071(.An(mai_mai_n92_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  INV        m072(.A(mai_mai_n94_), .Y(mai_mai_n95_));
  NOi21      m073(.An(x01), .B(x10), .Y(mai_mai_n96_));
  NO2        m074(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n97_));
  NO3        m075(.A(mai_mai_n97_), .B(mai_mai_n96_), .C(x06), .Y(mai_mai_n98_));
  NA2        m076(.A(mai_mai_n98_), .B(mai_mai_n27_), .Y(mai_mai_n99_));
  OAI210     m077(.A0(mai_mai_n95_), .A1(x07), .B0(mai_mai_n99_), .Y(mai_mai_n100_));
  NO3        m078(.A(mai_mai_n100_), .B(mai_mai_n90_), .C(mai_mai_n70_), .Y(mai01));
  INV        m079(.A(x12), .Y(mai_mai_n102_));
  INV        m080(.A(x13), .Y(mai_mai_n103_));
  NA2        m081(.A(mai_mai_n449_), .B(mai_mai_n71_), .Y(mai_mai_n104_));
  NA2        m082(.A(x08), .B(x04), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n105_), .B(mai_mai_n57_), .Y(mai_mai_n106_));
  NA2        m084(.A(mai_mai_n106_), .B(mai_mai_n104_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n96_), .B(mai_mai_n28_), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n108_), .B(mai_mai_n73_), .Y(mai_mai_n109_));
  NO2        m087(.A(x10), .B(x01), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n111_), .B(mai_mai_n110_), .Y(mai_mai_n112_));
  NA2        m090(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n113_));
  INV        m091(.A(mai_mai_n109_), .Y(mai_mai_n114_));
  AOI210     m092(.A0(mai_mai_n114_), .A1(mai_mai_n107_), .B0(mai_mai_n103_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n116_));
  NOi21      m094(.An(mai_mai_n116_), .B(mai_mai_n58_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n86_), .B(x13), .Y(mai_mai_n118_));
  NA2        m096(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NA2        m098(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n121_), .B(x05), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n122_), .B(mai_mai_n120_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n124_));
  INV        m102(.A(mai_mai_n117_), .Y(mai_mai_n125_));
  AOI210     m103(.A0(mai_mai_n125_), .A1(mai_mai_n123_), .B0(mai_mai_n74_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n127_));
  NA2        m105(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n130_));
  NO2        m108(.A(mai_mai_n124_), .B(mai_mai_n36_), .Y(mai_mai_n131_));
  NO2        m109(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n132_));
  NO3        m110(.A(mai_mai_n132_), .B(mai_mai_n131_), .C(mai_mai_n129_), .Y(mai_mai_n133_));
  NO3        m111(.A(mai_mai_n133_), .B(x06), .C(x03), .Y(mai_mai_n134_));
  NO3        m112(.A(mai_mai_n134_), .B(mai_mai_n126_), .C(mai_mai_n115_), .Y(mai_mai_n135_));
  NA2        m113(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n136_));
  OAI210     m114(.A0(mai_mai_n86_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n138_));
  NO2        m116(.A(mai_mai_n35_), .B(mai_mai_n47_), .Y(mai_mai_n139_));
  OA210      m117(.A0(x00), .A1(mai_mai_n79_), .B0(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m118(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n142_));
  AOI210     m120(.A0(mai_mai_n142_), .A1(mai_mai_n49_), .B0(mai_mai_n141_), .Y(mai_mai_n143_));
  OA210      m121(.A0(mai_mai_n143_), .A1(mai_mai_n140_), .B0(mai_mai_n138_), .Y(mai_mai_n144_));
  NO2        m122(.A(x09), .B(x05), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n145_), .B(mai_mai_n47_), .Y(mai_mai_n146_));
  AOI210     m124(.A0(mai_mai_n146_), .A1(mai_mai_n112_), .B0(mai_mai_n49_), .Y(mai_mai_n147_));
  NA2        m125(.A(x09), .B(x00), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n116_), .B(mai_mai_n148_), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n78_), .B(mai_mai_n51_), .Y(mai_mai_n150_));
  AOI210     m128(.A0(mai_mai_n150_), .A1(mai_mai_n149_), .B0(mai_mai_n142_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n147_), .C(mai_mai_n144_), .Y(mai_mai_n152_));
  NO2        m130(.A(x03), .B(x02), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n87_), .B(mai_mai_n103_), .Y(mai_mai_n154_));
  OAI210     m132(.A0(mai_mai_n154_), .A1(mai_mai_n117_), .B0(mai_mai_n153_), .Y(mai_mai_n155_));
  OA210      m133(.A0(mai_mai_n152_), .A1(x11), .B0(mai_mai_n155_), .Y(mai_mai_n156_));
  OAI210     m134(.A0(mai_mai_n135_), .A1(mai_mai_n23_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NA2        m135(.A(mai_mai_n112_), .B(mai_mai_n40_), .Y(mai_mai_n158_));
  NAi21      m136(.An(x06), .B(x10), .Y(mai_mai_n159_));
  NOi21      m137(.An(x01), .B(x13), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  BUFFER     m139(.A(mai_mai_n161_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n162_), .A1(mai_mai_n158_), .B0(mai_mai_n41_), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n164_));
  NA2        m142(.A(mai_mai_n103_), .B(x01), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n165_), .B(x08), .Y(mai_mai_n166_));
  OAI210     m144(.A0(x05), .A1(mai_mai_n166_), .B0(mai_mai_n51_), .Y(mai_mai_n167_));
  AOI210     m145(.A0(mai_mai_n167_), .A1(mai_mai_n164_), .B0(mai_mai_n48_), .Y(mai_mai_n168_));
  AOI210     m146(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n169_));
  OAI210     m147(.A0(mai_mai_n168_), .A1(mai_mai_n163_), .B0(mai_mai_n169_), .Y(mai_mai_n170_));
  NA2        m148(.A(x04), .B(x02), .Y(mai_mai_n171_));
  NA2        m149(.A(x10), .B(x05), .Y(mai_mai_n172_));
  INV        m150(.A(x06), .Y(mai_mai_n173_));
  NO2        m151(.A(x09), .B(x01), .Y(mai_mai_n174_));
  NO2        m152(.A(mai_mai_n116_), .B(x08), .Y(mai_mai_n175_));
  NA3        m153(.A(mai_mai_n160_), .B(mai_mai_n159_), .C(mai_mai_n51_), .Y(mai_mai_n176_));
  NO2        m154(.A(mai_mai_n176_), .B(x11), .Y(mai_mai_n177_));
  NAi21      m155(.An(mai_mai_n171_), .B(mai_mai_n177_), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n25_), .Y(mai_mai_n179_));
  NAi21      m157(.An(x13), .B(x00), .Y(mai_mai_n180_));
  AOI220     m158(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n181_));
  BUFFER     m159(.A(mai_mai_n73_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n97_), .B(x06), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n180_), .B(mai_mai_n36_), .Y(mai_mai_n184_));
  INV        m162(.A(mai_mai_n184_), .Y(mai_mai_n185_));
  OAI220     m163(.A0(mai_mai_n185_), .A1(mai_mai_n173_), .B0(mai_mai_n183_), .B1(mai_mai_n182_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n186_), .B(mai_mai_n179_), .Y(mai_mai_n187_));
  NOi21      m165(.An(x09), .B(x00), .Y(mai_mai_n188_));
  NO3        m166(.A(mai_mai_n85_), .B(mai_mai_n188_), .C(mai_mai_n47_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n128_), .Y(mai_mai_n190_));
  NA2        m168(.A(x06), .B(x05), .Y(mai_mai_n191_));
  OAI210     m169(.A0(mai_mai_n191_), .A1(mai_mai_n35_), .B0(mai_mai_n102_), .Y(mai_mai_n192_));
  AOI210     m170(.A0(x10), .A1(mai_mai_n58_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n193_), .B(mai_mai_n190_), .Y(mai_mai_n194_));
  NO2        m172(.A(mai_mai_n103_), .B(x12), .Y(mai_mai_n195_));
  AOI210     m173(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n195_), .Y(mai_mai_n196_));
  NA2        m174(.A(mai_mai_n96_), .B(mai_mai_n51_), .Y(mai_mai_n197_));
  NO2        m175(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n198_), .B(x02), .Y(mai_mai_n199_));
  NA2        m177(.A(mai_mai_n196_), .B(mai_mai_n194_), .Y(mai_mai_n200_));
  NA4        m178(.A(mai_mai_n200_), .B(mai_mai_n187_), .C(mai_mai_n178_), .D(mai_mai_n170_), .Y(mai_mai_n201_));
  AOI210     m179(.A0(mai_mai_n157_), .A1(mai_mai_n102_), .B0(mai_mai_n201_), .Y(mai_mai_n202_));
  INV        m180(.A(mai_mai_n75_), .Y(mai_mai_n203_));
  NA2        m181(.A(mai_mai_n203_), .B(mai_mai_n138_), .Y(mai_mai_n204_));
  NA2        m182(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n205_), .B(mai_mai_n137_), .Y(mai_mai_n206_));
  AOI210     m184(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n127_), .B(x06), .Y(mai_mai_n208_));
  AOI210     m186(.A0(mai_mai_n207_), .A1(mai_mai_n206_), .B0(mai_mai_n208_), .Y(mai_mai_n209_));
  AOI210     m187(.A0(mai_mai_n209_), .A1(mai_mai_n204_), .B0(x12), .Y(mai_mai_n210_));
  INV        m188(.A(mai_mai_n78_), .Y(mai_mai_n211_));
  NO2        m189(.A(x05), .B(mai_mai_n51_), .Y(mai_mai_n212_));
  OAI210     m190(.A0(mai_mai_n212_), .A1(mai_mai_n161_), .B0(mai_mai_n57_), .Y(mai_mai_n213_));
  NA2        m191(.A(mai_mai_n213_), .B(mai_mai_n211_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n96_), .B(x06), .Y(mai_mai_n215_));
  AOI210     m193(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n216_));
  NO3        m194(.A(mai_mai_n216_), .B(mai_mai_n215_), .C(mai_mai_n41_), .Y(mai_mai_n217_));
  INV        m195(.A(mai_mai_n142_), .Y(mai_mai_n218_));
  OAI210     m196(.A0(mai_mai_n218_), .A1(mai_mai_n217_), .B0(x02), .Y(mai_mai_n219_));
  AOI210     m197(.A0(mai_mai_n219_), .A1(mai_mai_n214_), .B0(mai_mai_n23_), .Y(mai_mai_n220_));
  OAI210     m198(.A0(mai_mai_n210_), .A1(mai_mai_n57_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  INV        m199(.A(mai_mai_n142_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n223_));
  OAI210     m201(.A0(mai_mai_n81_), .A1(mai_mai_n36_), .B0(mai_mai_n119_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n103_), .B(x03), .Y(mai_mai_n225_));
  AOI220     m203(.A0(mai_mai_n225_), .A1(mai_mai_n224_), .B0(mai_mai_n78_), .B1(mai_mai_n223_), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n159_), .Y(mai_mai_n228_));
  NOi21      m206(.An(x13), .B(x04), .Y(mai_mai_n229_));
  NO3        m207(.A(mai_mai_n229_), .B(mai_mai_n78_), .C(mai_mai_n188_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n230_), .B(x05), .Y(mai_mai_n231_));
  AOI220     m209(.A0(mai_mai_n231_), .A1(mai_mai_n227_), .B0(mai_mai_n228_), .B1(mai_mai_n57_), .Y(mai_mai_n232_));
  OAI210     m210(.A0(mai_mai_n226_), .A1(mai_mai_n222_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  INV        m211(.A(mai_mai_n93_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n234_), .B(x12), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n237_));
  AOI210     m215(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n238_));
  NO2        m216(.A(x06), .B(x00), .Y(mai_mai_n239_));
  NO3        m217(.A(mai_mai_n239_), .B(mai_mai_n238_), .C(mai_mai_n41_), .Y(mai_mai_n240_));
  INV        m218(.A(mai_mai_n74_), .Y(mai_mai_n241_));
  NO2        m219(.A(mai_mai_n241_), .B(mai_mai_n240_), .Y(mai_mai_n242_));
  NA2        m220(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n243_));
  NA2        m221(.A(mai_mai_n243_), .B(x03), .Y(mai_mai_n244_));
  OR2        m222(.A(mai_mai_n244_), .B(mai_mai_n242_), .Y(mai_mai_n245_));
  NA2        m223(.A(x13), .B(mai_mai_n102_), .Y(mai_mai_n246_));
  NA3        m224(.A(mai_mai_n246_), .B(mai_mai_n192_), .C(mai_mai_n94_), .Y(mai_mai_n247_));
  OAI210     m225(.A0(mai_mai_n245_), .A1(mai_mai_n236_), .B0(mai_mai_n247_), .Y(mai_mai_n248_));
  AOI210     m226(.A0(mai_mai_n235_), .A1(mai_mai_n233_), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  AOI210     m227(.A0(mai_mai_n249_), .A1(mai_mai_n221_), .B0(x07), .Y(mai_mai_n250_));
  NA2        m228(.A(mai_mai_n73_), .B(mai_mai_n29_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n229_), .B(mai_mai_n188_), .Y(mai_mai_n252_));
  AOI210     m230(.A0(mai_mai_n252_), .A1(mai_mai_n150_), .B0(mai_mai_n251_), .Y(mai_mai_n253_));
  NO2        m231(.A(mai_mai_n103_), .B(x06), .Y(mai_mai_n254_));
  INV        m232(.A(mai_mai_n254_), .Y(mai_mai_n255_));
  NO2        m233(.A(x08), .B(x05), .Y(mai_mai_n256_));
  NO2        m234(.A(mai_mai_n256_), .B(mai_mai_n238_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n78_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n258_));
  OAI210     m236(.A0(mai_mai_n257_), .A1(mai_mai_n255_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  NO2        m237(.A(x12), .B(x02), .Y(mai_mai_n260_));
  INV        m238(.A(mai_mai_n260_), .Y(mai_mai_n261_));
  NO2        m239(.A(mai_mai_n261_), .B(mai_mai_n234_), .Y(mai_mai_n262_));
  OA210      m240(.A0(mai_mai_n259_), .A1(mai_mai_n253_), .B0(mai_mai_n262_), .Y(mai_mai_n263_));
  NA2        m241(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n264_), .B(x01), .Y(mai_mai_n265_));
  NOi21      m243(.An(mai_mai_n86_), .B(mai_mai_n119_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n266_), .B(mai_mai_n265_), .Y(mai_mai_n267_));
  NO2        m245(.A(mai_mai_n267_), .B(mai_mai_n29_), .Y(mai_mai_n268_));
  NA2        m246(.A(mai_mai_n254_), .B(mai_mai_n224_), .Y(mai_mai_n269_));
  NA2        m247(.A(mai_mai_n103_), .B(x04), .Y(mai_mai_n270_));
  NA2        m248(.A(mai_mai_n270_), .B(mai_mai_n28_), .Y(mai_mai_n271_));
  OAI210     m249(.A0(mai_mai_n271_), .A1(mai_mai_n118_), .B0(mai_mai_n269_), .Y(mai_mai_n272_));
  NO3        m250(.A(mai_mai_n92_), .B(x12), .C(x03), .Y(mai_mai_n273_));
  OAI210     m251(.A0(mai_mai_n272_), .A1(mai_mai_n268_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  AOI210     m252(.A0(mai_mai_n197_), .A1(mai_mai_n191_), .B0(mai_mai_n105_), .Y(mai_mai_n275_));
  NOi21      m253(.An(mai_mai_n251_), .B(mai_mai_n215_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n277_));
  OAI210     m255(.A0(mai_mai_n276_), .A1(mai_mai_n275_), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n279_));
  NO3        m257(.A(mai_mai_n279_), .B(mai_mai_n216_), .C(mai_mai_n183_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n236_), .B(mai_mai_n28_), .Y(mai_mai_n281_));
  OAI210     m259(.A0(mai_mai_n280_), .A1(mai_mai_n222_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  NA3        m260(.A(mai_mai_n282_), .B(mai_mai_n278_), .C(mai_mai_n274_), .Y(mai_mai_n283_));
  NO3        m261(.A(mai_mai_n283_), .B(mai_mai_n263_), .C(mai_mai_n250_), .Y(mai_mai_n284_));
  OAI210     m262(.A0(mai_mai_n202_), .A1(mai_mai_n61_), .B0(mai_mai_n284_), .Y(mai02));
  AOI210     m263(.A0(mai_mai_n136_), .A1(mai_mai_n87_), .B0(mai_mai_n130_), .Y(mai_mai_n286_));
  NOi21      m264(.An(mai_mai_n230_), .B(mai_mai_n174_), .Y(mai_mai_n287_));
  NO2        m265(.A(mai_mai_n287_), .B(mai_mai_n32_), .Y(mai_mai_n288_));
  OAI210     m266(.A0(mai_mai_n288_), .A1(mai_mai_n286_), .B0(mai_mai_n172_), .Y(mai_mai_n289_));
  INV        m267(.A(mai_mai_n172_), .Y(mai_mai_n290_));
  INV        m268(.A(mai_mai_n216_), .Y(mai_mai_n291_));
  OAI220     m269(.A0(mai_mai_n291_), .A1(mai_mai_n103_), .B0(mai_mai_n87_), .B1(mai_mai_n51_), .Y(mai_mai_n292_));
  AOI220     m270(.A0(mai_mai_n292_), .A1(mai_mai_n290_), .B0(mai_mai_n154_), .B1(mai_mai_n153_), .Y(mai_mai_n293_));
  AOI210     m271(.A0(mai_mai_n293_), .A1(mai_mai_n289_), .B0(mai_mai_n48_), .Y(mai_mai_n294_));
  NO2        m272(.A(x05), .B(x02), .Y(mai_mai_n295_));
  OAI210     m273(.A0(mai_mai_n206_), .A1(mai_mai_n188_), .B0(mai_mai_n295_), .Y(mai_mai_n296_));
  AOI220     m274(.A0(mai_mai_n256_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n297_));
  NA2        m275(.A(mai_mai_n229_), .B(mai_mai_n81_), .Y(mai_mai_n298_));
  AOI210     m276(.A0(mai_mai_n298_), .A1(mai_mai_n296_), .B0(mai_mai_n142_), .Y(mai_mai_n299_));
  NAi21      m277(.An(mai_mai_n231_), .B(mai_mai_n226_), .Y(mai_mai_n300_));
  NO2        m278(.A(mai_mai_n243_), .B(mai_mai_n47_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n301_), .B(mai_mai_n300_), .Y(mai_mai_n302_));
  AN2        m280(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n303_));
  OAI210     m281(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n304_));
  NA2        m282(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n305_));
  OA210      m283(.A0(mai_mai_n305_), .A1(x08), .B0(mai_mai_n146_), .Y(mai_mai_n306_));
  AOI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n137_), .B0(mai_mai_n304_), .Y(mai_mai_n307_));
  OAI210     m285(.A0(mai_mai_n307_), .A1(mai_mai_n303_), .B0(mai_mai_n97_), .Y(mai_mai_n308_));
  NA3        m286(.A(mai_mai_n97_), .B(mai_mai_n86_), .C(mai_mai_n223_), .Y(mai_mai_n309_));
  NA3        m287(.A(mai_mai_n96_), .B(mai_mai_n85_), .C(mai_mai_n42_), .Y(mai_mai_n310_));
  AOI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n309_), .B0(x04), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n153_), .Y(mai_mai_n312_));
  OAI220     m290(.A0(mai_mai_n257_), .A1(mai_mai_n108_), .B0(mai_mai_n312_), .B1(mai_mai_n129_), .Y(mai_mai_n313_));
  AOI210     m291(.A0(mai_mai_n313_), .A1(x13), .B0(mai_mai_n311_), .Y(mai_mai_n314_));
  NA3        m292(.A(mai_mai_n314_), .B(mai_mai_n308_), .C(mai_mai_n302_), .Y(mai_mai_n315_));
  NO3        m293(.A(mai_mai_n315_), .B(mai_mai_n299_), .C(mai_mai_n294_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n141_), .B(x03), .Y(mai_mai_n317_));
  INV        m295(.A(mai_mai_n180_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n51_), .A1(mai_mai_n35_), .B0(mai_mai_n36_), .Y(mai_mai_n319_));
  AOI220     m297(.A0(mai_mai_n319_), .A1(mai_mai_n318_), .B0(mai_mai_n198_), .B1(x08), .Y(mai_mai_n320_));
  OAI210     m298(.A0(mai_mai_n320_), .A1(mai_mai_n279_), .B0(mai_mai_n317_), .Y(mai_mai_n321_));
  NA2        m299(.A(mai_mai_n321_), .B(mai_mai_n110_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n171_), .B(mai_mai_n165_), .Y(mai_mai_n323_));
  AN2        m301(.A(mai_mai_n323_), .B(mai_mai_n175_), .Y(mai_mai_n324_));
  INV        m302(.A(mai_mai_n56_), .Y(mai_mai_n325_));
  OAI220     m303(.A0(mai_mai_n270_), .A1(mai_mai_n325_), .B0(mai_mai_n130_), .B1(mai_mai_n28_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n326_), .A1(mai_mai_n324_), .B0(mai_mai_n111_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n270_), .B(mai_mai_n102_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n102_), .B(mai_mai_n41_), .Y(mai_mai_n329_));
  NA3        m307(.A(mai_mai_n329_), .B(mai_mai_n328_), .C(mai_mai_n129_), .Y(mai_mai_n330_));
  NA4        m308(.A(mai_mai_n330_), .B(mai_mai_n327_), .C(mai_mai_n322_), .D(mai_mai_n48_), .Y(mai_mai_n331_));
  INV        m309(.A(mai_mai_n198_), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n166_), .B(mai_mai_n40_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n334_));
  OAI220     m312(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n332_), .B1(mai_mai_n59_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n335_), .B(x02), .Y(mai_mai_n336_));
  INV        m314(.A(mai_mai_n237_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n195_), .B(x04), .Y(mai_mai_n338_));
  NO2        m316(.A(mai_mai_n338_), .B(mai_mai_n337_), .Y(mai_mai_n339_));
  NO3        m317(.A(mai_mai_n181_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n340_));
  OAI210     m318(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(mai_mai_n97_), .Y(mai_mai_n341_));
  NO3        m319(.A(mai_mai_n195_), .B(mai_mai_n164_), .C(mai_mai_n52_), .Y(mai_mai_n342_));
  OAI210     m320(.A0(mai_mai_n148_), .A1(mai_mai_n36_), .B0(mai_mai_n102_), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n189_), .B0(mai_mai_n342_), .Y(mai_mai_n344_));
  NA4        m322(.A(mai_mai_n344_), .B(mai_mai_n341_), .C(mai_mai_n336_), .D(x06), .Y(mai_mai_n345_));
  NA2        m323(.A(x09), .B(x03), .Y(mai_mai_n346_));
  OAI220     m324(.A0(mai_mai_n346_), .A1(mai_mai_n128_), .B0(mai_mai_n205_), .B1(mai_mai_n64_), .Y(mai_mai_n347_));
  OAI220     m325(.A0(mai_mai_n165_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n348_));
  NO3        m326(.A(mai_mai_n279_), .B(mai_mai_n127_), .C(x08), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n348_), .A1(mai_mai_n222_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n351_));
  NO3        m329(.A(mai_mai_n116_), .B(mai_mai_n128_), .C(mai_mai_n38_), .Y(mai_mai_n352_));
  AOI210     m330(.A0(mai_mai_n342_), .A1(mai_mai_n351_), .B0(mai_mai_n352_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n350_), .A1(mai_mai_n28_), .B0(mai_mai_n353_), .Y(mai_mai_n354_));
  AO220      m332(.A0(mai_mai_n354_), .A1(x04), .B0(mai_mai_n347_), .B1(x05), .Y(mai_mai_n355_));
  AOI210     m333(.A0(mai_mai_n345_), .A1(mai_mai_n331_), .B0(mai_mai_n355_), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n316_), .A1(x12), .B0(mai_mai_n356_), .Y(mai03));
  OR2        m335(.A(mai_mai_n42_), .B(mai_mai_n223_), .Y(mai_mai_n358_));
  AOI210     m336(.A0(mai_mai_n154_), .A1(mai_mai_n102_), .B0(mai_mai_n358_), .Y(mai_mai_n359_));
  AO210      m337(.A0(mai_mai_n337_), .A1(mai_mai_n88_), .B0(mai_mai_n338_), .Y(mai_mai_n360_));
  NA2        m338(.A(mai_mai_n195_), .B(mai_mai_n153_), .Y(mai_mai_n361_));
  NA3        m339(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n199_), .Y(mai_mai_n362_));
  OAI210     m340(.A0(mai_mai_n362_), .A1(mai_mai_n359_), .B0(x05), .Y(mai_mai_n363_));
  NA2        m341(.A(mai_mai_n358_), .B(x05), .Y(mai_mai_n364_));
  AOI210     m342(.A0(mai_mai_n137_), .A1(mai_mai_n211_), .B0(mai_mai_n364_), .Y(mai_mai_n365_));
  AOI210     m343(.A0(mai_mai_n225_), .A1(mai_mai_n82_), .B0(mai_mai_n122_), .Y(mai_mai_n366_));
  OAI220     m344(.A0(mai_mai_n366_), .A1(mai_mai_n59_), .B0(mai_mai_n305_), .B1(mai_mai_n297_), .Y(mai_mai_n367_));
  OAI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n365_), .B0(mai_mai_n102_), .Y(mai_mai_n368_));
  AOI210     m346(.A0(mai_mai_n146_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n174_), .B(mai_mai_n132_), .Y(mai_mai_n370_));
  OAI220     m348(.A0(mai_mai_n370_), .A1(mai_mai_n37_), .B0(mai_mai_n149_), .B1(x13), .Y(mai_mai_n371_));
  OAI210     m349(.A0(mai_mai_n371_), .A1(mai_mai_n369_), .B0(x04), .Y(mai_mai_n372_));
  NO3        m350(.A(mai_mai_n329_), .B(mai_mai_n87_), .C(mai_mai_n59_), .Y(mai_mai_n373_));
  AOI210     m351(.A0(mai_mai_n185_), .A1(mai_mai_n102_), .B0(mai_mai_n146_), .Y(mai_mai_n374_));
  OA210      m352(.A0(mai_mai_n166_), .A1(x12), .B0(mai_mai_n132_), .Y(mai_mai_n375_));
  NO3        m353(.A(mai_mai_n375_), .B(mai_mai_n374_), .C(mai_mai_n373_), .Y(mai_mai_n376_));
  NA4        m354(.A(mai_mai_n376_), .B(mai_mai_n372_), .C(mai_mai_n368_), .D(mai_mai_n363_), .Y(mai04));
  NO2        m355(.A(mai_mai_n91_), .B(mai_mai_n39_), .Y(mai_mai_n378_));
  XO2        m356(.A(mai_mai_n378_), .B(mai_mai_n246_), .Y(mai05));
  AOI210     m357(.A0(mai_mai_n73_), .A1(mai_mai_n52_), .B0(mai_mai_n208_), .Y(mai_mai_n380_));
  AOI210     m358(.A0(mai_mai_n380_), .A1(mai_mai_n304_), .B0(mai_mai_n25_), .Y(mai_mai_n381_));
  NA3        m359(.A(mai_mai_n142_), .B(mai_mai_n130_), .C(mai_mai_n31_), .Y(mai_mai_n382_));
  NO2        m360(.A(mai_mai_n382_), .B(mai_mai_n24_), .Y(mai_mai_n383_));
  OAI210     m361(.A0(mai_mai_n383_), .A1(mai_mai_n381_), .B0(mai_mai_n102_), .Y(mai_mai_n384_));
  NA2        m362(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n251_), .B(x03), .Y(mai_mai_n387_));
  OAI220     m365(.A0(mai_mai_n387_), .A1(mai_mai_n386_), .B0(mai_mai_n385_), .B1(mai_mai_n83_), .Y(mai_mai_n388_));
  OAI210     m366(.A0(mai_mai_n26_), .A1(mai_mai_n102_), .B0(x07), .Y(mai_mai_n389_));
  AOI210     m367(.A0(mai_mai_n388_), .A1(x06), .B0(mai_mai_n389_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n71_), .B(x02), .Y(mai_mai_n391_));
  AOI210     m369(.A0(mai_mai_n391_), .A1(mai_mai_n387_), .B0(mai_mai_n254_), .Y(mai_mai_n392_));
  OR2        m370(.A(mai_mai_n392_), .B(mai_mai_n236_), .Y(mai_mai_n393_));
  NA2        m371(.A(mai_mai_n160_), .B(x05), .Y(mai_mai_n394_));
  NA3        m372(.A(mai_mai_n394_), .B(mai_mai_n239_), .C(mai_mai_n234_), .Y(mai_mai_n395_));
  NA2        m373(.A(mai_mai_n395_), .B(mai_mai_n393_), .Y(mai_mai_n396_));
  NA2        m374(.A(mai_mai_n396_), .B(mai_mai_n102_), .Y(mai_mai_n397_));
  NA2        m375(.A(mai_mai_n33_), .B(mai_mai_n102_), .Y(mai_mai_n398_));
  AOI210     m376(.A0(mai_mai_n398_), .A1(mai_mai_n93_), .B0(x07), .Y(mai_mai_n399_));
  AOI220     m377(.A0(mai_mai_n399_), .A1(mai_mai_n397_), .B0(mai_mai_n390_), .B1(mai_mai_n384_), .Y(mai_mai_n400_));
  NA3        m378(.A(mai_mai_n23_), .B(mai_mai_n61_), .C(mai_mai_n48_), .Y(mai_mai_n401_));
  AO210      m379(.A0(mai_mai_n401_), .A1(mai_mai_n264_), .B0(mai_mai_n261_), .Y(mai_mai_n402_));
  AOI210     m380(.A0(x11), .A1(mai_mai_n76_), .B0(mai_mai_n141_), .Y(mai_mai_n403_));
  OR2        m381(.A(mai_mai_n403_), .B(x03), .Y(mai_mai_n404_));
  NA2        m382(.A(mai_mai_n351_), .B(mai_mai_n61_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n405_), .B(x11), .Y(mai_mai_n406_));
  NO3        m384(.A(mai_mai_n406_), .B(mai_mai_n145_), .C(mai_mai_n28_), .Y(mai_mai_n407_));
  AOI220     m385(.A0(mai_mai_n407_), .A1(mai_mai_n404_), .B0(mai_mai_n402_), .B1(mai_mai_n47_), .Y(mai_mai_n408_));
  NO3        m386(.A(mai_mai_n329_), .B(mai_mai_n32_), .C(x11), .Y(mai_mai_n409_));
  OAI210     m387(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(mai_mai_n103_), .Y(mai_mai_n410_));
  AOI210     m388(.A0(mai_mai_n338_), .A1(mai_mai_n113_), .B0(mai_mai_n260_), .Y(mai_mai_n411_));
  NOi21      m389(.An(mai_mai_n317_), .B(mai_mai_n132_), .Y(mai_mai_n412_));
  NO2        m390(.A(mai_mai_n412_), .B(mai_mai_n261_), .Y(mai_mai_n413_));
  OAI210     m391(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n414_));
  AOI210     m392(.A0(mai_mai_n246_), .A1(mai_mai_n47_), .B0(mai_mai_n414_), .Y(mai_mai_n415_));
  NO4        m393(.A(mai_mai_n415_), .B(mai_mai_n413_), .C(mai_mai_n411_), .D(x08), .Y(mai_mai_n416_));
  OAI210     m394(.A0(x05), .A1(x03), .B0(mai_mai_n385_), .Y(mai_mai_n417_));
  NO2        m395(.A(x13), .B(x12), .Y(mai_mai_n418_));
  NO2        m396(.A(mai_mai_n130_), .B(mai_mai_n28_), .Y(mai_mai_n419_));
  NO2        m397(.A(mai_mai_n419_), .B(mai_mai_n265_), .Y(mai_mai_n420_));
  OR3        m398(.A(mai_mai_n420_), .B(x12), .C(x03), .Y(mai_mai_n421_));
  NA3        m399(.A(mai_mai_n332_), .B(mai_mai_n124_), .C(x12), .Y(mai_mai_n422_));
  AO210      m400(.A0(mai_mai_n332_), .A1(mai_mai_n124_), .B0(mai_mai_n246_), .Y(mai_mai_n423_));
  NA4        m401(.A(mai_mai_n423_), .B(mai_mai_n422_), .C(mai_mai_n421_), .D(x08), .Y(mai_mai_n424_));
  AOI210     m402(.A0(mai_mai_n418_), .A1(mai_mai_n417_), .B0(mai_mai_n424_), .Y(mai_mai_n425_));
  AOI210     m403(.A0(mai_mai_n416_), .A1(mai_mai_n410_), .B0(mai_mai_n425_), .Y(mai_mai_n426_));
  OAI210     m404(.A0(mai_mai_n405_), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n427_));
  OAI220     m405(.A0(mai_mai_n448_), .A1(mai_mai_n386_), .B0(mai_mai_n145_), .B1(mai_mai_n43_), .Y(mai_mai_n428_));
  OAI210     m406(.A0(mai_mai_n428_), .A1(mai_mai_n427_), .B0(mai_mai_n184_), .Y(mai_mai_n429_));
  NA3        m407(.A(mai_mai_n420_), .B(mai_mai_n412_), .C(mai_mai_n328_), .Y(mai_mai_n430_));
  INV        m408(.A(x14), .Y(mai_mai_n431_));
  NO3        m409(.A(mai_mai_n317_), .B(mai_mai_n108_), .C(x11), .Y(mai_mai_n432_));
  NO3        m410(.A(mai_mai_n165_), .B(mai_mai_n76_), .C(mai_mai_n57_), .Y(mai_mai_n433_));
  NO3        m411(.A(mai_mai_n401_), .B(mai_mai_n329_), .C(mai_mai_n180_), .Y(mai_mai_n434_));
  NO4        m412(.A(mai_mai_n434_), .B(mai_mai_n433_), .C(mai_mai_n432_), .D(mai_mai_n431_), .Y(mai_mai_n435_));
  NA3        m413(.A(mai_mai_n435_), .B(mai_mai_n430_), .C(mai_mai_n429_), .Y(mai_mai_n436_));
  AOI220     m414(.A0(mai_mai_n398_), .A1(mai_mai_n61_), .B0(mai_mai_n419_), .B1(mai_mai_n164_), .Y(mai_mai_n437_));
  NOi21      m415(.An(mai_mai_n270_), .B(mai_mai_n149_), .Y(mai_mai_n438_));
  NO3        m416(.A(mai_mai_n127_), .B(mai_mai_n24_), .C(x06), .Y(mai_mai_n439_));
  AOI210     m417(.A0(mai_mai_n277_), .A1(mai_mai_n228_), .B0(mai_mai_n439_), .Y(mai_mai_n440_));
  OAI210     m418(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n440_), .Y(mai_mai_n441_));
  OAI210     m419(.A0(mai_mai_n441_), .A1(mai_mai_n438_), .B0(mai_mai_n102_), .Y(mai_mai_n442_));
  OAI210     m420(.A0(mai_mai_n437_), .A1(mai_mai_n92_), .B0(mai_mai_n442_), .Y(mai_mai_n443_));
  NO4        m421(.A(mai_mai_n443_), .B(mai_mai_n436_), .C(mai_mai_n426_), .D(mai_mai_n400_), .Y(mai06));
  INV        m422(.A(x07), .Y(mai_mai_n447_));
  INV        m423(.A(x07), .Y(mai_mai_n448_));
  INV        m424(.A(x01), .Y(mai_mai_n449_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  INV        u027(.A(x09), .Y(men_men_n50_));
  NO2        u028(.A(x10), .B(x02), .Y(men_men_n51_));
  NOi21      u029(.An(x01), .B(x09), .Y(men_men_n52_));
  INV        u030(.A(x00), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n50_), .B(men_men_n53_), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n54_), .B(men_men_n52_), .Y(men_men_n55_));
  NA2        u033(.A(x09), .B(men_men_n53_), .Y(men_men_n56_));
  INV        u034(.A(x07), .Y(men_men_n57_));
  AOI220     u035(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n57_), .Y(men_men_n58_));
  INV        u036(.A(men_men_n55_), .Y(men_men_n59_));
  NA2        u037(.A(men_men_n29_), .B(x02), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n60_), .B(men_men_n24_), .Y(men_men_n61_));
  OAI220     u039(.A0(men_men_n61_), .A1(men_men_n59_), .B0(men_men_n58_), .B1(men_men_n56_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n57_), .B(men_men_n48_), .Y(men_men_n63_));
  OAI210     u041(.A0(men_men_n30_), .A1(x11), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u042(.A0(men_men_n64_), .A1(men_men_n55_), .B0(men_men_n62_), .B1(men_men_n31_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n65_), .B(x05), .Y(men_men_n66_));
  NO2        u044(.A(men_men_n57_), .B(men_men_n23_), .Y(men_men_n67_));
  NA2        u045(.A(x09), .B(x05), .Y(men_men_n68_));
  NA2        u046(.A(x10), .B(x06), .Y(men_men_n69_));
  NA3        u047(.A(men_men_n69_), .B(men_men_n68_), .C(men_men_n28_), .Y(men_men_n70_));
  NO2        u048(.A(men_men_n57_), .B(men_men_n41_), .Y(men_men_n71_));
  OAI210     u049(.A0(men_men_n70_), .A1(men_men_n67_), .B0(x03), .Y(men_men_n72_));
  NOi31      u050(.An(x08), .B(x04), .C(x00), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n445_), .B(men_men_n24_), .Y(men_men_n74_));
  NO2        u052(.A(x09), .B(men_men_n41_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n75_), .B(men_men_n36_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n77_));
  AOI210     u055(.A0(men_men_n76_), .A1(men_men_n48_), .B0(men_men_n77_), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n36_), .B(x00), .Y(men_men_n79_));
  NO2        u057(.A(x08), .B(x01), .Y(men_men_n80_));
  OAI210     u058(.A0(men_men_n80_), .A1(men_men_n79_), .B0(men_men_n35_), .Y(men_men_n81_));
  NA2        u059(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n82_));
  NO3        u060(.A(men_men_n81_), .B(men_men_n78_), .C(men_men_n74_), .Y(men_men_n83_));
  AN2        u061(.A(men_men_n83_), .B(men_men_n72_), .Y(men_men_n84_));
  INV        u062(.A(men_men_n81_), .Y(men_men_n85_));
  NO2        u063(.A(x06), .B(x05), .Y(men_men_n86_));
  NA2        u064(.A(x11), .B(x00), .Y(men_men_n87_));
  NO2        u065(.A(x11), .B(men_men_n47_), .Y(men_men_n88_));
  NOi21      u066(.An(men_men_n87_), .B(men_men_n88_), .Y(men_men_n89_));
  AOI210     u067(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n89_), .Y(men_men_n90_));
  NOi21      u068(.An(x01), .B(x10), .Y(men_men_n91_));
  NO2        u069(.A(men_men_n29_), .B(men_men_n53_), .Y(men_men_n92_));
  NO3        u070(.A(men_men_n92_), .B(men_men_n91_), .C(x06), .Y(men_men_n93_));
  NA2        u071(.A(men_men_n93_), .B(men_men_n27_), .Y(men_men_n94_));
  OAI210     u072(.A0(men_men_n90_), .A1(x07), .B0(men_men_n94_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n84_), .C(men_men_n66_), .Y(men01));
  INV        u074(.A(x12), .Y(men_men_n97_));
  INV        u075(.A(x13), .Y(men_men_n98_));
  NA2        u076(.A(x08), .B(x04), .Y(men_men_n99_));
  NO2        u077(.A(men_men_n99_), .B(men_men_n53_), .Y(men_men_n100_));
  NA2        u078(.A(men_men_n100_), .B(men_men_n86_), .Y(men_men_n101_));
  NA2        u079(.A(men_men_n91_), .B(men_men_n28_), .Y(men_men_n102_));
  NO2        u080(.A(x10), .B(x01), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n29_), .B(x00), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n103_), .Y(men_men_n105_));
  NA2        u083(.A(x04), .B(men_men_n28_), .Y(men_men_n106_));
  NO3        u084(.A(men_men_n106_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n107_));
  NA2        u085(.A(men_men_n107_), .B(men_men_n105_), .Y(men_men_n108_));
  AOI210     u086(.A0(men_men_n108_), .A1(men_men_n101_), .B0(men_men_n98_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n52_), .B(x05), .Y(men_men_n110_));
  NOi21      u088(.An(men_men_n110_), .B(men_men_n54_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n35_), .B(x02), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n98_), .B(men_men_n36_), .Y(men_men_n113_));
  NA3        u091(.A(men_men_n113_), .B(men_men_n112_), .C(x06), .Y(men_men_n114_));
  INV        u092(.A(men_men_n114_), .Y(men_men_n115_));
  INV        u093(.A(x13), .Y(men_men_n116_));
  NA2        u094(.A(x09), .B(men_men_n35_), .Y(men_men_n117_));
  NA2        u095(.A(x13), .B(men_men_n35_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n118_), .B(x05), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n35_), .B(men_men_n53_), .Y(men_men_n120_));
  AOI210     u098(.A0(men_men_n53_), .A1(men_men_n76_), .B0(men_men_n111_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(men_men_n69_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n123_));
  NA2        u101(.A(x10), .B(men_men_n53_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n50_), .B(x05), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n36_), .B(x04), .Y(men_men_n127_));
  NA3        u105(.A(men_men_n127_), .B(men_men_n126_), .C(x13), .Y(men_men_n128_));
  NO3        u106(.A(men_men_n120_), .B(men_men_n75_), .C(men_men_n36_), .Y(men_men_n129_));
  NO2        u107(.A(men_men_n56_), .B(x05), .Y(men_men_n130_));
  NOi41      u108(.An(men_men_n128_), .B(men_men_n130_), .C(men_men_n129_), .D(men_men_n125_), .Y(men_men_n131_));
  NO3        u109(.A(men_men_n131_), .B(x06), .C(x03), .Y(men_men_n132_));
  NO4        u110(.A(men_men_n132_), .B(men_men_n122_), .C(men_men_n115_), .D(men_men_n109_), .Y(men_men_n133_));
  NA2        u111(.A(x13), .B(men_men_n36_), .Y(men_men_n134_));
  OAI210     u112(.A0(men_men_n80_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(men_men_n134_), .Y(men_men_n136_));
  NO2        u114(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n137_));
  AN2        u115(.A(men_men_n86_), .B(men_men_n137_), .Y(men_men_n138_));
  NO2        u116(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n29_), .B(x06), .Y(men_men_n140_));
  AOI210     u118(.A0(men_men_n140_), .A1(men_men_n49_), .B0(men_men_n139_), .Y(men_men_n141_));
  OA210      u119(.A0(men_men_n141_), .A1(men_men_n138_), .B0(men_men_n136_), .Y(men_men_n142_));
  NO2        u120(.A(x09), .B(x05), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n143_), .B(men_men_n47_), .Y(men_men_n144_));
  NO2        u122(.A(men_men_n105_), .B(men_men_n49_), .Y(men_men_n145_));
  NA2        u123(.A(x09), .B(x00), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n110_), .B(men_men_n146_), .Y(men_men_n147_));
  INV        u125(.A(men_men_n73_), .Y(men_men_n148_));
  NO2        u126(.A(men_men_n147_), .B(men_men_n140_), .Y(men_men_n149_));
  NO3        u127(.A(men_men_n149_), .B(men_men_n145_), .C(men_men_n142_), .Y(men_men_n150_));
  NO2        u128(.A(x03), .B(x02), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n81_), .B(men_men_n98_), .Y(men_men_n152_));
  OAI210     u130(.A0(men_men_n152_), .A1(men_men_n111_), .B0(men_men_n151_), .Y(men_men_n153_));
  OA210      u131(.A0(men_men_n150_), .A1(x11), .B0(men_men_n153_), .Y(men_men_n154_));
  OAI210     u132(.A0(men_men_n133_), .A1(men_men_n23_), .B0(men_men_n154_), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n105_), .B(men_men_n40_), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n157_));
  NAi21      u135(.An(x06), .B(x10), .Y(men_men_n158_));
  NOi21      u136(.An(x01), .B(x13), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  OR2        u138(.A(men_men_n160_), .B(men_men_n157_), .Y(men_men_n161_));
  AOI210     u139(.A0(men_men_n161_), .A1(men_men_n156_), .B0(men_men_n41_), .Y(men_men_n162_));
  NO2        u140(.A(men_men_n29_), .B(x03), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n98_), .B(x01), .Y(men_men_n164_));
  NO2        u142(.A(men_men_n164_), .B(x08), .Y(men_men_n165_));
  NO2        u143(.A(men_men_n163_), .B(men_men_n48_), .Y(men_men_n166_));
  AOI210     u144(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n167_));
  OAI210     u145(.A0(men_men_n166_), .A1(men_men_n162_), .B0(men_men_n167_), .Y(men_men_n168_));
  NA2        u146(.A(x04), .B(x02), .Y(men_men_n169_));
  NA2        u147(.A(x10), .B(x05), .Y(men_men_n170_));
  NA2        u148(.A(x09), .B(x06), .Y(men_men_n171_));
  AOI210     u149(.A0(men_men_n171_), .A1(men_men_n170_), .B0(men_men_n157_), .Y(men_men_n172_));
  NO2        u150(.A(x09), .B(x01), .Y(men_men_n173_));
  NO3        u151(.A(men_men_n173_), .B(men_men_n103_), .C(men_men_n31_), .Y(men_men_n174_));
  OAI210     u152(.A0(men_men_n174_), .A1(men_men_n172_), .B0(x00), .Y(men_men_n175_));
  NO2        u153(.A(men_men_n110_), .B(x08), .Y(men_men_n176_));
  NA3        u154(.A(men_men_n159_), .B(men_men_n158_), .C(men_men_n50_), .Y(men_men_n177_));
  NA2        u155(.A(men_men_n91_), .B(x05), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n178_), .A1(men_men_n113_), .B0(men_men_n177_), .Y(men_men_n179_));
  AOI210     u157(.A0(men_men_n176_), .A1(x06), .B0(men_men_n179_), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(x11), .B0(men_men_n175_), .Y(men_men_n181_));
  NAi21      u159(.An(men_men_n169_), .B(men_men_n181_), .Y(men_men_n182_));
  INV        u160(.A(men_men_n25_), .Y(men_men_n183_));
  NAi21      u161(.An(x13), .B(x00), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n184_), .Y(men_men_n185_));
  AOI220     u163(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n186_));
  OAI210     u164(.A0(men_men_n170_), .A1(men_men_n35_), .B0(men_men_n186_), .Y(men_men_n187_));
  AN2        u165(.A(men_men_n187_), .B(men_men_n185_), .Y(men_men_n188_));
  AN2        u166(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n189_));
  NO2        u167(.A(men_men_n92_), .B(x06), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n184_), .B(men_men_n36_), .Y(men_men_n191_));
  INV        u169(.A(men_men_n191_), .Y(men_men_n192_));
  OAI220     u170(.A0(men_men_n192_), .A1(men_men_n171_), .B0(men_men_n190_), .B1(men_men_n189_), .Y(men_men_n193_));
  OAI210     u171(.A0(men_men_n193_), .A1(men_men_n188_), .B0(men_men_n183_), .Y(men_men_n194_));
  NOi21      u172(.An(x09), .B(x00), .Y(men_men_n195_));
  NO3        u173(.A(men_men_n79_), .B(men_men_n195_), .C(men_men_n47_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n196_), .B(men_men_n124_), .Y(men_men_n197_));
  NA2        u175(.A(x10), .B(x08), .Y(men_men_n198_));
  INV        u176(.A(men_men_n198_), .Y(men_men_n199_));
  NA2        u177(.A(x06), .B(x05), .Y(men_men_n200_));
  OAI210     u178(.A0(men_men_n200_), .A1(men_men_n35_), .B0(men_men_n97_), .Y(men_men_n201_));
  AOI210     u179(.A0(men_men_n199_), .A1(men_men_n54_), .B0(men_men_n201_), .Y(men_men_n202_));
  NA2        u180(.A(men_men_n202_), .B(men_men_n197_), .Y(men_men_n203_));
  NO2        u181(.A(men_men_n98_), .B(x12), .Y(men_men_n204_));
  AOI210     u182(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n204_), .Y(men_men_n205_));
  NA2        u183(.A(men_men_n91_), .B(men_men_n50_), .Y(men_men_n206_));
  NO2        u184(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n207_), .B(x02), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n208_), .B(men_men_n206_), .Y(men_men_n209_));
  AOI210     u187(.A0(men_men_n205_), .A1(men_men_n203_), .B0(men_men_n209_), .Y(men_men_n210_));
  NA4        u188(.A(men_men_n210_), .B(men_men_n194_), .C(men_men_n182_), .D(men_men_n168_), .Y(men_men_n211_));
  AOI210     u189(.A0(men_men_n155_), .A1(men_men_n97_), .B0(men_men_n211_), .Y(men_men_n212_));
  INV        u190(.A(men_men_n70_), .Y(men_men_n213_));
  NA2        u191(.A(men_men_n213_), .B(men_men_n136_), .Y(men_men_n214_));
  NA2        u192(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(men_men_n135_), .Y(men_men_n216_));
  AOI210     u194(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n123_), .B(x06), .Y(men_men_n218_));
  AOI210     u196(.A0(men_men_n217_), .A1(men_men_n216_), .B0(men_men_n218_), .Y(men_men_n219_));
  AOI210     u197(.A0(men_men_n219_), .A1(men_men_n214_), .B0(x12), .Y(men_men_n220_));
  INV        u198(.A(men_men_n73_), .Y(men_men_n221_));
  NO2        u199(.A(x05), .B(men_men_n50_), .Y(men_men_n222_));
  OAI210     u200(.A0(men_men_n222_), .A1(men_men_n160_), .B0(men_men_n53_), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n223_), .B(men_men_n221_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n91_), .B(x06), .Y(men_men_n225_));
  AOI210     u203(.A0(men_men_n36_), .A1(x04), .B0(men_men_n50_), .Y(men_men_n226_));
  NO3        u204(.A(men_men_n226_), .B(men_men_n225_), .C(men_men_n41_), .Y(men_men_n227_));
  NA4        u205(.A(men_men_n158_), .B(men_men_n52_), .C(men_men_n36_), .D(x04), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n228_), .B(men_men_n140_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n229_), .A1(men_men_n227_), .B0(x02), .Y(men_men_n230_));
  AOI210     u208(.A0(men_men_n230_), .A1(men_men_n224_), .B0(men_men_n23_), .Y(men_men_n231_));
  OAI210     u209(.A0(men_men_n220_), .A1(men_men_n53_), .B0(men_men_n231_), .Y(men_men_n232_));
  INV        u210(.A(men_men_n140_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n50_), .B(x03), .Y(men_men_n234_));
  OAI210     u212(.A0(men_men_n75_), .A1(men_men_n36_), .B0(men_men_n117_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n98_), .B(x03), .Y(men_men_n236_));
  AOI220     u214(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n73_), .B1(men_men_n234_), .Y(men_men_n237_));
  NA2        u215(.A(men_men_n32_), .B(x06), .Y(men_men_n238_));
  INV        u216(.A(men_men_n158_), .Y(men_men_n239_));
  NOi21      u217(.An(x13), .B(x04), .Y(men_men_n240_));
  NO3        u218(.A(men_men_n240_), .B(men_men_n73_), .C(men_men_n195_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n241_), .B(x05), .Y(men_men_n242_));
  AOI220     u220(.A0(men_men_n242_), .A1(men_men_n238_), .B0(men_men_n239_), .B1(men_men_n53_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n237_), .A1(men_men_n233_), .B0(men_men_n243_), .Y(men_men_n244_));
  INV        u222(.A(men_men_n88_), .Y(men_men_n245_));
  NO2        u223(.A(men_men_n245_), .B(x12), .Y(men_men_n246_));
  NA2        u224(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n50_), .B(men_men_n36_), .Y(men_men_n248_));
  OAI210     u226(.A0(men_men_n248_), .A1(men_men_n187_), .B0(men_men_n185_), .Y(men_men_n249_));
  AOI210     u227(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n99_), .A1(men_men_n146_), .B0(men_men_n69_), .Y(men_men_n251_));
  INV        u229(.A(men_men_n251_), .Y(men_men_n252_));
  NA2        u230(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n253_), .B(x03), .Y(men_men_n254_));
  OA210      u232(.A0(men_men_n254_), .A1(men_men_n252_), .B0(men_men_n249_), .Y(men_men_n255_));
  NA2        u233(.A(x13), .B(men_men_n97_), .Y(men_men_n256_));
  NA3        u234(.A(men_men_n256_), .B(men_men_n201_), .C(men_men_n89_), .Y(men_men_n257_));
  OAI210     u235(.A0(men_men_n255_), .A1(men_men_n247_), .B0(men_men_n257_), .Y(men_men_n258_));
  AOI210     u236(.A0(men_men_n246_), .A1(men_men_n244_), .B0(men_men_n258_), .Y(men_men_n259_));
  AOI210     u237(.A0(men_men_n259_), .A1(men_men_n232_), .B0(x07), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n68_), .B(men_men_n29_), .Y(men_men_n261_));
  AOI210     u239(.A0(men_men_n134_), .A1(men_men_n148_), .B0(men_men_n261_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n98_), .B(x06), .Y(men_men_n263_));
  INV        u241(.A(men_men_n263_), .Y(men_men_n264_));
  NO2        u242(.A(x08), .B(x05), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n265_), .B(men_men_n250_), .Y(men_men_n266_));
  OAI210     u244(.A0(men_men_n73_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n267_));
  OAI210     u245(.A0(men_men_n266_), .A1(men_men_n264_), .B0(men_men_n267_), .Y(men_men_n268_));
  NO2        u246(.A(x12), .B(x02), .Y(men_men_n269_));
  INV        u247(.A(men_men_n269_), .Y(men_men_n270_));
  NO2        u248(.A(men_men_n270_), .B(men_men_n245_), .Y(men_men_n271_));
  OA210      u249(.A0(men_men_n268_), .A1(men_men_n262_), .B0(men_men_n271_), .Y(men_men_n272_));
  NA2        u250(.A(men_men_n50_), .B(men_men_n41_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n273_), .B(x01), .Y(men_men_n274_));
  NOi21      u252(.An(men_men_n80_), .B(men_men_n117_), .Y(men_men_n275_));
  NO2        u253(.A(men_men_n275_), .B(men_men_n274_), .Y(men_men_n276_));
  AOI210     u254(.A0(men_men_n276_), .A1(men_men_n128_), .B0(men_men_n29_), .Y(men_men_n277_));
  NA2        u255(.A(men_men_n263_), .B(men_men_n235_), .Y(men_men_n278_));
  NA2        u256(.A(men_men_n98_), .B(x04), .Y(men_men_n279_));
  OAI210     u257(.A0(x02), .A1(men_men_n116_), .B0(men_men_n278_), .Y(men_men_n280_));
  NO3        u258(.A(men_men_n87_), .B(x12), .C(x03), .Y(men_men_n281_));
  OAI210     u259(.A0(men_men_n280_), .A1(men_men_n277_), .B0(men_men_n281_), .Y(men_men_n282_));
  NOi21      u260(.An(men_men_n261_), .B(men_men_n225_), .Y(men_men_n283_));
  NO2        u261(.A(men_men_n25_), .B(x00), .Y(men_men_n284_));
  NA2        u262(.A(men_men_n283_), .B(men_men_n284_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n54_), .B(x05), .Y(men_men_n286_));
  NO3        u264(.A(men_men_n286_), .B(men_men_n226_), .C(men_men_n190_), .Y(men_men_n287_));
  NO2        u265(.A(men_men_n247_), .B(men_men_n28_), .Y(men_men_n288_));
  OAI210     u266(.A0(men_men_n287_), .A1(men_men_n233_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA3        u267(.A(men_men_n289_), .B(men_men_n285_), .C(men_men_n282_), .Y(men_men_n290_));
  NO3        u268(.A(men_men_n290_), .B(men_men_n272_), .C(men_men_n260_), .Y(men_men_n291_));
  OAI210     u269(.A0(men_men_n212_), .A1(men_men_n57_), .B0(men_men_n291_), .Y(men02));
  AOI210     u270(.A0(men_men_n134_), .A1(men_men_n81_), .B0(men_men_n126_), .Y(men_men_n293_));
  NOi21      u271(.An(men_men_n241_), .B(men_men_n173_), .Y(men_men_n294_));
  NO2        u272(.A(men_men_n98_), .B(men_men_n35_), .Y(men_men_n295_));
  NA3        u273(.A(men_men_n295_), .B(men_men_n199_), .C(men_men_n52_), .Y(men_men_n296_));
  OAI210     u274(.A0(men_men_n294_), .A1(men_men_n32_), .B0(men_men_n296_), .Y(men_men_n297_));
  OAI210     u275(.A0(men_men_n297_), .A1(men_men_n293_), .B0(men_men_n170_), .Y(men_men_n298_));
  INV        u276(.A(men_men_n170_), .Y(men_men_n299_));
  AOI210     u277(.A0(men_men_n112_), .A1(men_men_n82_), .B0(men_men_n226_), .Y(men_men_n300_));
  OAI220     u278(.A0(men_men_n300_), .A1(men_men_n98_), .B0(men_men_n81_), .B1(men_men_n50_), .Y(men_men_n301_));
  AOI220     u279(.A0(men_men_n301_), .A1(men_men_n299_), .B0(men_men_n152_), .B1(men_men_n151_), .Y(men_men_n302_));
  AOI210     u280(.A0(men_men_n302_), .A1(men_men_n298_), .B0(men_men_n48_), .Y(men_men_n303_));
  NO2        u281(.A(x05), .B(x02), .Y(men_men_n304_));
  OAI210     u282(.A0(men_men_n216_), .A1(men_men_n195_), .B0(men_men_n304_), .Y(men_men_n305_));
  AOI220     u283(.A0(men_men_n265_), .A1(men_men_n54_), .B0(men_men_n52_), .B1(men_men_n36_), .Y(men_men_n306_));
  NOi21      u284(.An(men_men_n295_), .B(men_men_n306_), .Y(men_men_n307_));
  AOI210     u285(.A0(men_men_n240_), .A1(men_men_n75_), .B0(men_men_n307_), .Y(men_men_n308_));
  AOI210     u286(.A0(men_men_n308_), .A1(men_men_n305_), .B0(men_men_n140_), .Y(men_men_n309_));
  NAi21      u287(.An(men_men_n242_), .B(men_men_n237_), .Y(men_men_n310_));
  NO2        u288(.A(men_men_n253_), .B(men_men_n47_), .Y(men_men_n311_));
  NA2        u289(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n312_));
  AN2        u290(.A(men_men_n236_), .B(men_men_n235_), .Y(men_men_n313_));
  OAI210     u291(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n314_));
  NA2        u292(.A(x13), .B(men_men_n28_), .Y(men_men_n315_));
  OA210      u293(.A0(men_men_n315_), .A1(x08), .B0(men_men_n144_), .Y(men_men_n316_));
  AOI210     u294(.A0(men_men_n316_), .A1(men_men_n135_), .B0(men_men_n314_), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n317_), .A1(men_men_n313_), .B0(men_men_n92_), .Y(men_men_n318_));
  NA3        u296(.A(men_men_n92_), .B(men_men_n80_), .C(men_men_n234_), .Y(men_men_n319_));
  NA3        u297(.A(men_men_n91_), .B(men_men_n79_), .C(men_men_n42_), .Y(men_men_n320_));
  AOI210     u298(.A0(men_men_n320_), .A1(men_men_n319_), .B0(x04), .Y(men_men_n321_));
  INV        u299(.A(men_men_n151_), .Y(men_men_n322_));
  OAI220     u300(.A0(men_men_n266_), .A1(men_men_n102_), .B0(men_men_n322_), .B1(men_men_n125_), .Y(men_men_n323_));
  AOI210     u301(.A0(men_men_n323_), .A1(x13), .B0(men_men_n321_), .Y(men_men_n324_));
  NA3        u302(.A(men_men_n324_), .B(men_men_n318_), .C(men_men_n312_), .Y(men_men_n325_));
  NO3        u303(.A(men_men_n325_), .B(men_men_n309_), .C(men_men_n303_), .Y(men_men_n326_));
  NA2        u304(.A(men_men_n139_), .B(x03), .Y(men_men_n327_));
  INV        u305(.A(men_men_n184_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n50_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n329_));
  AOI220     u307(.A0(men_men_n329_), .A1(men_men_n328_), .B0(men_men_n207_), .B1(x08), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n330_), .A1(men_men_n286_), .B0(men_men_n327_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n331_), .B(men_men_n103_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n169_), .B(men_men_n164_), .Y(men_men_n333_));
  AN2        u311(.A(men_men_n333_), .B(men_men_n176_), .Y(men_men_n334_));
  NO2        u312(.A(men_men_n126_), .B(men_men_n28_), .Y(men_men_n335_));
  OAI210     u313(.A0(men_men_n335_), .A1(men_men_n334_), .B0(men_men_n104_), .Y(men_men_n336_));
  NA2        u314(.A(men_men_n279_), .B(men_men_n97_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n97_), .B(men_men_n41_), .Y(men_men_n338_));
  NA3        u316(.A(men_men_n338_), .B(men_men_n337_), .C(men_men_n125_), .Y(men_men_n339_));
  NA4        u317(.A(men_men_n339_), .B(men_men_n336_), .C(men_men_n332_), .D(men_men_n48_), .Y(men_men_n340_));
  INV        u318(.A(men_men_n207_), .Y(men_men_n341_));
  NO2        u319(.A(men_men_n165_), .B(men_men_n40_), .Y(men_men_n342_));
  NA2        u320(.A(men_men_n32_), .B(x05), .Y(men_men_n343_));
  OAI220     u321(.A0(men_men_n343_), .A1(men_men_n342_), .B0(men_men_n341_), .B1(men_men_n55_), .Y(men_men_n344_));
  NA2        u322(.A(men_men_n344_), .B(x02), .Y(men_men_n345_));
  INV        u323(.A(men_men_n248_), .Y(men_men_n346_));
  NA2        u324(.A(men_men_n204_), .B(x04), .Y(men_men_n347_));
  NO3        u325(.A(men_men_n204_), .B(men_men_n163_), .C(men_men_n51_), .Y(men_men_n348_));
  OAI210     u326(.A0(men_men_n146_), .A1(men_men_n36_), .B0(men_men_n97_), .Y(men_men_n349_));
  OAI210     u327(.A0(men_men_n349_), .A1(men_men_n196_), .B0(men_men_n348_), .Y(men_men_n350_));
  NA3        u328(.A(men_men_n350_), .B(men_men_n345_), .C(x06), .Y(men_men_n351_));
  NA2        u329(.A(x09), .B(x03), .Y(men_men_n352_));
  OAI220     u330(.A0(men_men_n352_), .A1(men_men_n124_), .B0(men_men_n215_), .B1(men_men_n60_), .Y(men_men_n353_));
  OAI220     u331(.A0(men_men_n164_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n354_));
  NO3        u332(.A(men_men_n286_), .B(men_men_n123_), .C(x08), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n354_), .A1(men_men_n233_), .B0(men_men_n355_), .Y(men_men_n356_));
  NO2        u334(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n357_));
  NO3        u335(.A(men_men_n110_), .B(men_men_n124_), .C(men_men_n38_), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n348_), .A1(men_men_n357_), .B0(men_men_n358_), .Y(men_men_n359_));
  OAI210     u337(.A0(men_men_n356_), .A1(men_men_n28_), .B0(men_men_n359_), .Y(men_men_n360_));
  AO220      u338(.A0(men_men_n360_), .A1(x04), .B0(men_men_n353_), .B1(x05), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n351_), .A1(men_men_n340_), .B0(men_men_n361_), .Y(men_men_n362_));
  OAI210     u340(.A0(men_men_n326_), .A1(x12), .B0(men_men_n362_), .Y(men03));
  OR2        u341(.A(men_men_n42_), .B(men_men_n234_), .Y(men_men_n364_));
  AOI210     u342(.A0(men_men_n152_), .A1(men_men_n97_), .B0(men_men_n364_), .Y(men_men_n365_));
  AO210      u343(.A0(men_men_n346_), .A1(men_men_n82_), .B0(men_men_n347_), .Y(men_men_n366_));
  NA2        u344(.A(men_men_n204_), .B(men_men_n151_), .Y(men_men_n367_));
  NA3        u345(.A(men_men_n367_), .B(men_men_n366_), .C(men_men_n208_), .Y(men_men_n368_));
  OAI210     u346(.A0(men_men_n368_), .A1(men_men_n365_), .B0(x05), .Y(men_men_n369_));
  NA2        u347(.A(men_men_n364_), .B(x05), .Y(men_men_n370_));
  AOI210     u348(.A0(men_men_n135_), .A1(men_men_n221_), .B0(men_men_n370_), .Y(men_men_n371_));
  AOI210     u349(.A0(men_men_n236_), .A1(men_men_n76_), .B0(men_men_n119_), .Y(men_men_n372_));
  OAI220     u350(.A0(men_men_n372_), .A1(men_men_n55_), .B0(men_men_n315_), .B1(men_men_n306_), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n371_), .B0(men_men_n97_), .Y(men_men_n374_));
  AOI210     u352(.A0(men_men_n144_), .A1(men_men_n56_), .B0(men_men_n38_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n173_), .B(men_men_n130_), .Y(men_men_n376_));
  OAI220     u354(.A0(men_men_n376_), .A1(men_men_n37_), .B0(men_men_n147_), .B1(x13), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n377_), .A1(men_men_n375_), .B0(x04), .Y(men_men_n378_));
  NO3        u356(.A(men_men_n338_), .B(men_men_n81_), .C(men_men_n55_), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n192_), .A1(men_men_n97_), .B0(men_men_n144_), .Y(men_men_n380_));
  OA210      u358(.A0(men_men_n165_), .A1(x12), .B0(men_men_n130_), .Y(men_men_n381_));
  NO3        u359(.A(men_men_n381_), .B(men_men_n380_), .C(men_men_n379_), .Y(men_men_n382_));
  NA4        u360(.A(men_men_n382_), .B(men_men_n378_), .C(men_men_n374_), .D(men_men_n369_), .Y(men04));
  NO2        u361(.A(men_men_n85_), .B(men_men_n39_), .Y(men_men_n384_));
  XO2        u362(.A(men_men_n384_), .B(men_men_n256_), .Y(men05));
  NO2        u363(.A(men_men_n51_), .B(men_men_n218_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n386_), .A1(men_men_n314_), .B0(men_men_n25_), .Y(men_men_n387_));
  NO2        u365(.A(x06), .B(men_men_n24_), .Y(men_men_n388_));
  OAI210     u366(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n97_), .Y(men_men_n389_));
  NA2        u367(.A(x11), .B(men_men_n31_), .Y(men_men_n390_));
  NO2        u368(.A(men_men_n390_), .B(men_men_n77_), .Y(men_men_n391_));
  OAI210     u369(.A0(men_men_n26_), .A1(men_men_n97_), .B0(x07), .Y(men_men_n392_));
  AOI210     u370(.A0(men_men_n391_), .A1(x06), .B0(men_men_n392_), .Y(men_men_n393_));
  AOI220     u371(.A0(men_men_n77_), .A1(men_men_n31_), .B0(men_men_n51_), .B1(men_men_n50_), .Y(men_men_n394_));
  NO3        u372(.A(men_men_n394_), .B(men_men_n23_), .C(x00), .Y(men_men_n395_));
  NO2        u373(.A(men_men_n23_), .B(x10), .Y(men_men_n396_));
  OR3        u374(.A(x06), .B(men_men_n396_), .C(men_men_n44_), .Y(men_men_n397_));
  NA2        u375(.A(men_men_n397_), .B(men_men_n247_), .Y(men_men_n398_));
  OAI210     u376(.A0(men_men_n398_), .A1(men_men_n395_), .B0(men_men_n97_), .Y(men_men_n399_));
  NA2        u377(.A(men_men_n33_), .B(men_men_n97_), .Y(men_men_n400_));
  AOI210     u378(.A0(men_men_n400_), .A1(men_men_n88_), .B0(x07), .Y(men_men_n401_));
  AOI220     u379(.A0(men_men_n401_), .A1(men_men_n399_), .B0(men_men_n393_), .B1(men_men_n389_), .Y(men_men_n402_));
  OR2        u380(.A(men_men_n273_), .B(men_men_n270_), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n396_), .A1(men_men_n71_), .B0(men_men_n139_), .Y(men_men_n404_));
  OR2        u382(.A(men_men_n404_), .B(x03), .Y(men_men_n405_));
  NA2        u383(.A(men_men_n357_), .B(men_men_n57_), .Y(men_men_n406_));
  NO2        u384(.A(men_men_n406_), .B(x11), .Y(men_men_n407_));
  NO3        u385(.A(men_men_n407_), .B(men_men_n143_), .C(men_men_n28_), .Y(men_men_n408_));
  AOI220     u386(.A0(men_men_n408_), .A1(men_men_n405_), .B0(men_men_n403_), .B1(men_men_n47_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n409_), .B(men_men_n98_), .Y(men_men_n410_));
  AOI210     u388(.A0(men_men_n347_), .A1(men_men_n106_), .B0(men_men_n269_), .Y(men_men_n411_));
  NOi21      u389(.An(men_men_n327_), .B(men_men_n130_), .Y(men_men_n412_));
  NO2        u390(.A(men_men_n412_), .B(men_men_n270_), .Y(men_men_n413_));
  OAI210     u391(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n414_));
  AOI210     u392(.A0(men_men_n256_), .A1(men_men_n47_), .B0(men_men_n414_), .Y(men_men_n415_));
  NO4        u393(.A(men_men_n415_), .B(men_men_n413_), .C(men_men_n411_), .D(x08), .Y(men_men_n416_));
  NA2        u394(.A(x09), .B(men_men_n41_), .Y(men_men_n417_));
  OAI210     u395(.A0(men_men_n390_), .A1(men_men_n63_), .B0(men_men_n417_), .Y(men_men_n418_));
  NO2        u396(.A(x13), .B(x12), .Y(men_men_n419_));
  NO2        u397(.A(men_men_n126_), .B(men_men_n28_), .Y(men_men_n420_));
  NO2        u398(.A(men_men_n420_), .B(men_men_n274_), .Y(men_men_n421_));
  OR3        u399(.A(men_men_n421_), .B(x12), .C(x03), .Y(men_men_n422_));
  NA3        u400(.A(men_men_n341_), .B(men_men_n120_), .C(x12), .Y(men_men_n423_));
  AO210      u401(.A0(men_men_n341_), .A1(men_men_n120_), .B0(men_men_n256_), .Y(men_men_n424_));
  NA4        u402(.A(men_men_n424_), .B(men_men_n423_), .C(men_men_n422_), .D(x08), .Y(men_men_n425_));
  AOI210     u403(.A0(men_men_n419_), .A1(men_men_n418_), .B0(men_men_n425_), .Y(men_men_n426_));
  AOI210     u404(.A0(men_men_n416_), .A1(men_men_n410_), .B0(men_men_n426_), .Y(men_men_n427_));
  OAI210     u405(.A0(men_men_n406_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n428_));
  NO2        u406(.A(men_men_n170_), .B(x02), .Y(men_men_n429_));
  OAI210     u407(.A0(men_men_n429_), .A1(men_men_n428_), .B0(men_men_n191_), .Y(men_men_n430_));
  NA3        u408(.A(men_men_n421_), .B(men_men_n412_), .C(men_men_n337_), .Y(men_men_n431_));
  INV        u409(.A(x14), .Y(men_men_n432_));
  NO3        u410(.A(men_men_n327_), .B(men_men_n102_), .C(x11), .Y(men_men_n433_));
  NO3        u411(.A(men_men_n164_), .B(men_men_n71_), .C(men_men_n53_), .Y(men_men_n434_));
  NO3        u412(.A(men_men_n434_), .B(men_men_n433_), .C(men_men_n432_), .Y(men_men_n435_));
  NA3        u413(.A(men_men_n435_), .B(men_men_n431_), .C(men_men_n430_), .Y(men_men_n436_));
  NA2        u414(.A(men_men_n400_), .B(men_men_n57_), .Y(men_men_n437_));
  NOi21      u415(.An(men_men_n279_), .B(men_men_n147_), .Y(men_men_n438_));
  NO2        u416(.A(men_men_n44_), .B(x04), .Y(men_men_n439_));
  OAI210     u417(.A0(men_men_n439_), .A1(men_men_n438_), .B0(men_men_n97_), .Y(men_men_n440_));
  OAI210     u418(.A0(men_men_n437_), .A1(men_men_n87_), .B0(men_men_n440_), .Y(men_men_n441_));
  NO4        u419(.A(men_men_n441_), .B(men_men_n436_), .C(men_men_n427_), .D(men_men_n402_), .Y(men06));
  INV        u420(.A(x07), .Y(men_men_n445_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule