// Benchmark "top" written by ABC on Thu Jun 20 14:59:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n139_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1095_,
    new_new_n1096_, new_new_n1097_, new_new_n1098_, new_new_n1099_,
    new_new_n1100_, new_new_n1101_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  NA2        g0029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g0030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NO2        g0031(.A(new_new_n53_), .B(new_new_n52_), .Y(new_new_n54_));
  NA3        g0032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g0033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g0034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  INV        g0035(.A(new_new_n55_), .Y(new_new_n58_));
  NA2        g0036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g0037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g0038(.A(i_1_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g0040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n63_));
  NA2        g0041(.A(i_1_), .B(i_10_), .Y(new_new_n64_));
  NO2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NAi31      g0043(.An(new_new_n65_), .B(new_new_n63_), .C(new_new_n59_), .Y(new_new_n66_));
  NA2        g0044(.A(new_new_n51_), .B(i_2_), .Y(new_new_n67_));
  AOI210     g0045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n68_));
  NA2        g0046(.A(i_1_), .B(i_6_), .Y(new_new_n69_));
  NO2        g0047(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n70_));
  INV        g0048(.A(i_0_), .Y(new_new_n71_));
  NAi21      g0049(.An(i_5_), .B(i_10_), .Y(new_new_n72_));
  NA2        g0050(.A(i_5_), .B(i_9_), .Y(new_new_n73_));
  AOI210     g0051(.A0(new_new_n73_), .A1(new_new_n72_), .B0(new_new_n71_), .Y(new_new_n74_));
  NO2        g0052(.A(new_new_n74_), .B(new_new_n70_), .Y(new_new_n75_));
  OAI210     g0053(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n75_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n76_), .A1(new_new_n66_), .B0(i_0_), .Y(new_new_n77_));
  NA2        g0055(.A(i_12_), .B(i_5_), .Y(new_new_n78_));
  NA2        g0056(.A(i_2_), .B(i_8_), .Y(new_new_n79_));
  NO2        g0057(.A(i_3_), .B(i_9_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_7_), .Y(new_new_n81_));
  NO3        g0059(.A(new_new_n81_), .B(new_new_n80_), .C(new_new_n61_), .Y(new_new_n82_));
  INV        g0060(.A(i_6_), .Y(new_new_n83_));
  OR4        g0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  INV        g0062(.A(new_new_n84_), .Y(new_new_n85_));
  NO2        g0063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  NO2        g0064(.A(new_new_n85_), .B(new_new_n86_), .Y(new_new_n87_));
  NA2        g0065(.A(new_new_n82_), .B(new_new_n87_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n61_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g0070(.A(new_new_n92_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g0071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n88_), .B0(new_new_n78_), .Y(new_new_n95_));
  AN3        g0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g0074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g0075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g0076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g0077(.A0(new_new_n99_), .A1(new_new_n60_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g0078(.A(i_7_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n47_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g0080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(new_new_n83_), .Y(new_new_n104_));
  NA2        g0082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g0083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g0084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g0085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  NO3        g0086(.A(new_new_n108_), .B(new_new_n89_), .C(new_new_n52_), .Y(new_new_n109_));
  AN2        g0087(.A(i_2_), .B(i_10_), .Y(new_new_n110_));
  NO2        g0088(.A(new_new_n110_), .B(i_7_), .Y(new_new_n111_));
  OR2        g0089(.A(new_new_n78_), .B(new_new_n56_), .Y(new_new_n112_));
  NO2        g0090(.A(i_8_), .B(new_new_n101_), .Y(new_new_n113_));
  NO3        g0091(.A(new_new_n113_), .B(new_new_n112_), .C(new_new_n111_), .Y(new_new_n114_));
  NA2        g0092(.A(i_12_), .B(i_7_), .Y(new_new_n115_));
  NO2        g0093(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n116_));
  NA2        g0094(.A(new_new_n116_), .B(i_0_), .Y(new_new_n117_));
  NA2        g0095(.A(i_11_), .B(i_12_), .Y(new_new_n118_));
  OAI210     g0096(.A0(new_new_n117_), .A1(new_new_n115_), .B0(new_new_n118_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n119_), .B(new_new_n114_), .Y(new_new_n120_));
  NAi41      g0098(.An(new_new_n109_), .B(new_new_n120_), .C(new_new_n107_), .D(new_new_n100_), .Y(new_new_n121_));
  NOi21      g0099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g0102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g0104(.A(new_new_n126_), .B(new_new_n47_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n128_));
  NAi21      g0106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n60_), .Y(new_new_n130_));
  NOi21      g0108(.An(new_new_n130_), .B(new_new_n128_), .Y(new_new_n131_));
  NO2        g0109(.A(i_1_), .B(new_new_n83_), .Y(new_new_n132_));
  NO2        g0110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  AO210      g0112(.A0(new_new_n134_), .A1(new_new_n48_), .B0(new_new_n132_), .Y(new_new_n135_));
  OAI220     g0113(.A0(new_new_n135_), .A1(new_new_n108_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n136_));
  NO3        g0114(.A(new_new_n136_), .B(new_new_n121_), .C(new_new_n95_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(new_new_n77_), .Y(men2));
  NO2        g0116(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n139_));
  NA2        g0117(.A(i_6_), .B(new_new_n25_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(new_new_n139_), .Y(new_new_n141_));
  NA4        g0119(.A(new_new_n141_), .B(new_new_n75_), .C(new_new_n67_), .D(new_new_n30_), .Y(men0));
  AN2        g0120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g0122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g0123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g0124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g0125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g0126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  OR2        g0129(.A(new_new_n151_), .B(new_new_n25_), .Y(new_new_n152_));
  AN2        g0130(.A(new_new_n145_), .B(new_new_n80_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(new_new_n27_), .Y(new_new_n154_));
  NA2        g0132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n71_), .B(new_new_n47_), .Y(new_new_n156_));
  NA2        g0134(.A(new_new_n156_), .B(new_new_n36_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n158_));
  OR2        g0136(.A(i_0_), .B(i_1_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n78_), .C(i_13_), .Y(new_new_n160_));
  NAi32      g0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n161_));
  NAi21      g0139(.An(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NOi21      g0140(.An(i_4_), .B(i_10_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n40_), .Y(new_new_n164_));
  NO2        g0142(.A(i_3_), .B(i_5_), .Y(new_new_n165_));
  NO3        g0143(.A(new_new_n71_), .B(i_2_), .C(i_1_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  OAI210     g0145(.A0(new_new_n167_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n168_));
  NO2        g0146(.A(new_new_n168_), .B(new_new_n158_), .Y(new_new_n169_));
  AOI210     g0147(.A0(new_new_n169_), .A1(new_new_n152_), .B0(new_new_n144_), .Y(new_new_n170_));
  NA2        g0148(.A(i_3_), .B(new_new_n49_), .Y(new_new_n171_));
  NOi21      g0149(.An(i_4_), .B(i_9_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_11_), .B(i_13_), .Y(new_new_n173_));
  NA2        g0151(.A(new_new_n173_), .B(new_new_n172_), .Y(new_new_n174_));
  NO2        g0152(.A(i_4_), .B(i_5_), .Y(new_new_n175_));
  NAi21      g0153(.An(i_12_), .B(i_11_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n176_), .B(i_13_), .Y(new_new_n177_));
  NA3        g0155(.A(new_new_n177_), .B(new_new_n175_), .C(new_new_n80_), .Y(new_new_n178_));
  AOI210     g0156(.A0(new_new_n178_), .A1(new_new_n174_), .B0(i_2_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n71_), .B(new_new_n61_), .Y(new_new_n180_));
  NAi31      g0158(.An(new_new_n1101_), .B(new_new_n153_), .C(i_11_), .Y(new_new_n181_));
  NA2        g0159(.A(i_3_), .B(i_5_), .Y(new_new_n182_));
  AOI210     g0160(.A0(new_new_n174_), .A1(new_new_n181_), .B0(i_2_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n71_), .B(i_5_), .Y(new_new_n184_));
  NO2        g0162(.A(i_13_), .B(i_10_), .Y(new_new_n185_));
  NA3        g0163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n45_), .Y(new_new_n186_));
  NO2        g0164(.A(i_2_), .B(i_1_), .Y(new_new_n187_));
  NA2        g0165(.A(new_new_n187_), .B(i_3_), .Y(new_new_n188_));
  NAi21      g0166(.An(i_4_), .B(i_12_), .Y(new_new_n189_));
  NO4        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n186_), .D(new_new_n25_), .Y(new_new_n190_));
  NO3        g0168(.A(new_new_n190_), .B(new_new_n183_), .C(new_new_n179_), .Y(new_new_n191_));
  INV        g0169(.A(i_8_), .Y(new_new_n192_));
  NO2        g0170(.A(new_new_n192_), .B(i_7_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_6_), .Y(new_new_n194_));
  NO3        g0172(.A(i_3_), .B(new_new_n83_), .C(new_new_n49_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(new_new_n113_), .Y(new_new_n196_));
  NO3        g0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n197_));
  NA3        g0175(.A(new_new_n197_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n198_));
  NO3        g0176(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n199_));
  OAI210     g0177(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n199_), .Y(new_new_n200_));
  AOI210     g0178(.A0(new_new_n200_), .A1(new_new_n198_), .B0(new_new_n196_), .Y(new_new_n201_));
  NO2        g0179(.A(i_3_), .B(i_8_), .Y(new_new_n202_));
  NO3        g0180(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n202_), .C(new_new_n40_), .Y(new_new_n204_));
  NO2        g0182(.A(new_new_n103_), .B(new_new_n56_), .Y(new_new_n205_));
  NO2        g0183(.A(i_13_), .B(i_9_), .Y(new_new_n206_));
  NA3        g0184(.A(new_new_n206_), .B(i_6_), .C(new_new_n192_), .Y(new_new_n207_));
  NAi21      g0185(.An(i_12_), .B(i_3_), .Y(new_new_n208_));
  OR2        g0186(.A(new_new_n208_), .B(new_new_n207_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n45_), .B(i_5_), .Y(new_new_n210_));
  NO3        g0188(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n211_));
  NA2        g0189(.A(new_new_n211_), .B(i_10_), .Y(new_new_n212_));
  OAI220     g0190(.A0(new_new_n212_), .A1(new_new_n209_), .B0(new_new_n103_), .B1(new_new_n204_), .Y(new_new_n213_));
  AOI210     g0191(.A0(new_new_n213_), .A1(i_7_), .B0(new_new_n201_), .Y(new_new_n214_));
  OAI220     g0192(.A0(new_new_n214_), .A1(i_4_), .B0(new_new_n194_), .B1(new_new_n191_), .Y(new_new_n215_));
  NAi21      g0193(.An(i_12_), .B(i_7_), .Y(new_new_n216_));
  NA3        g0194(.A(i_13_), .B(new_new_n192_), .C(i_10_), .Y(new_new_n217_));
  NO2        g0195(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n218_));
  NA2        g0196(.A(i_0_), .B(i_5_), .Y(new_new_n219_));
  NA2        g0197(.A(new_new_n219_), .B(new_new_n104_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n220_), .A1(new_new_n188_), .B0(i_2_), .B1(new_new_n134_), .Y(new_new_n221_));
  NAi31      g0199(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n36_), .B(i_13_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n71_), .B(new_new_n26_), .Y(new_new_n224_));
  NO2        g0202(.A(new_new_n47_), .B(new_new_n61_), .Y(new_new_n225_));
  NA3        g0203(.A(new_new_n225_), .B(new_new_n224_), .C(new_new_n223_), .Y(new_new_n226_));
  INV        g0204(.A(i_13_), .Y(new_new_n227_));
  NO2        g0205(.A(i_12_), .B(new_new_n227_), .Y(new_new_n228_));
  NA3        g0206(.A(new_new_n228_), .B(new_new_n197_), .C(new_new_n195_), .Y(new_new_n229_));
  OAI210     g0207(.A0(new_new_n226_), .A1(new_new_n222_), .B0(new_new_n229_), .Y(new_new_n230_));
  AOI220     g0208(.A0(new_new_n230_), .A1(new_new_n143_), .B0(new_new_n221_), .B1(new_new_n218_), .Y(new_new_n231_));
  NO2        g0209(.A(i_12_), .B(new_new_n37_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n182_), .B(i_4_), .Y(new_new_n233_));
  NA2        g0211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  OR2        g0212(.A(i_8_), .B(i_7_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n235_), .B(new_new_n83_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n52_), .B(i_1_), .Y(new_new_n237_));
  NA2        g0215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  INV        g0216(.A(i_12_), .Y(new_new_n239_));
  NO3        g0217(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n240_));
  NA2        g0218(.A(i_2_), .B(i_1_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n238_), .B(new_new_n234_), .Y(new_new_n242_));
  NO3        g0220(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n243_));
  NAi21      g0221(.An(i_4_), .B(i_3_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n244_), .B(new_new_n73_), .Y(new_new_n245_));
  NO2        g0223(.A(i_0_), .B(i_6_), .Y(new_new_n246_));
  NOi41      g0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n247_), .B(new_new_n246_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n241_), .B(new_new_n182_), .Y(new_new_n249_));
  NA2        g0227(.A(new_new_n242_), .B(new_new_n206_), .Y(new_new_n250_));
  NO2        g0228(.A(i_11_), .B(new_new_n227_), .Y(new_new_n251_));
  NOi21      g0229(.An(i_1_), .B(i_6_), .Y(new_new_n252_));
  NAi21      g0230(.An(i_3_), .B(i_7_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n239_), .B(i_9_), .Y(new_new_n254_));
  OR4        g0232(.A(new_new_n254_), .B(new_new_n253_), .C(new_new_n252_), .D(new_new_n184_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n256_));
  NO2        g0234(.A(i_12_), .B(i_3_), .Y(new_new_n257_));
  NA2        g0235(.A(new_new_n71_), .B(i_5_), .Y(new_new_n258_));
  NA2        g0236(.A(i_3_), .B(i_9_), .Y(new_new_n259_));
  NAi21      g0237(.An(i_7_), .B(i_10_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n260_), .B(new_new_n259_), .Y(new_new_n261_));
  NA3        g0239(.A(new_new_n261_), .B(new_new_n258_), .C(new_new_n62_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n262_), .B(new_new_n255_), .Y(new_new_n263_));
  NA3        g0241(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n264_));
  NA2        g0242(.A(new_new_n263_), .B(new_new_n251_), .Y(new_new_n265_));
  NO2        g0243(.A(new_new_n235_), .B(new_new_n37_), .Y(new_new_n266_));
  NA2        g0244(.A(i_12_), .B(i_6_), .Y(new_new_n267_));
  OR2        g0245(.A(i_13_), .B(i_9_), .Y(new_new_n268_));
  NO3        g0246(.A(new_new_n268_), .B(new_new_n267_), .C(new_new_n49_), .Y(new_new_n269_));
  NO2        g0247(.A(new_new_n244_), .B(i_2_), .Y(new_new_n270_));
  NA3        g0248(.A(new_new_n270_), .B(new_new_n269_), .C(new_new_n45_), .Y(new_new_n271_));
  NA2        g0249(.A(new_new_n251_), .B(i_9_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n258_), .B(new_new_n62_), .Y(new_new_n273_));
  OAI210     g0251(.A0(new_new_n273_), .A1(new_new_n272_), .B0(new_new_n271_), .Y(new_new_n274_));
  NA2        g0252(.A(new_new_n156_), .B(new_new_n61_), .Y(new_new_n275_));
  NO3        g0253(.A(i_11_), .B(new_new_n227_), .C(new_new_n25_), .Y(new_new_n276_));
  NO2        g0254(.A(new_new_n253_), .B(i_8_), .Y(new_new_n277_));
  NO2        g0255(.A(i_6_), .B(new_new_n49_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n277_), .C(new_new_n276_), .Y(new_new_n279_));
  NO3        g0257(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n280_));
  NA3        g0258(.A(new_new_n280_), .B(new_new_n266_), .C(new_new_n228_), .Y(new_new_n281_));
  AOI210     g0259(.A0(new_new_n281_), .A1(new_new_n279_), .B0(new_new_n275_), .Y(new_new_n282_));
  AOI210     g0260(.A0(new_new_n274_), .A1(new_new_n266_), .B0(new_new_n282_), .Y(new_new_n283_));
  NA4        g0261(.A(new_new_n283_), .B(new_new_n265_), .C(new_new_n250_), .D(new_new_n231_), .Y(new_new_n284_));
  NO3        g0262(.A(i_12_), .B(new_new_n227_), .C(new_new_n37_), .Y(new_new_n285_));
  INV        g0263(.A(new_new_n285_), .Y(new_new_n286_));
  NA2        g0264(.A(i_8_), .B(new_new_n101_), .Y(new_new_n287_));
  NOi21      g0265(.An(new_new_n165_), .B(new_new_n83_), .Y(new_new_n288_));
  NO3        g0266(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n289_));
  AOI220     g0267(.A0(new_new_n289_), .A1(new_new_n195_), .B0(new_new_n288_), .B1(new_new_n237_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n290_), .B(new_new_n287_), .Y(new_new_n291_));
  NO3        g0269(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n241_), .B(i_0_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n193_), .B0(new_new_n292_), .B1(new_new_n143_), .Y(new_new_n294_));
  NA2        g0272(.A(new_new_n278_), .B(new_new_n26_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n295_), .B(new_new_n294_), .Y(new_new_n296_));
  NA2        g0274(.A(i_0_), .B(i_1_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(i_2_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n57_), .B(i_6_), .Y(new_new_n299_));
  NA3        g0277(.A(new_new_n299_), .B(new_new_n298_), .C(new_new_n165_), .Y(new_new_n300_));
  OAI210     g0278(.A0(new_new_n167_), .A1(new_new_n144_), .B0(new_new_n300_), .Y(new_new_n301_));
  NO3        g0279(.A(new_new_n301_), .B(new_new_n296_), .C(new_new_n291_), .Y(new_new_n302_));
  NO2        g0280(.A(i_3_), .B(i_10_), .Y(new_new_n303_));
  NA3        g0281(.A(new_new_n303_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n304_));
  NO2        g0282(.A(i_2_), .B(new_new_n101_), .Y(new_new_n305_));
  NOi21      g0283(.An(new_new_n219_), .B(new_new_n103_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(i_1_), .C(new_new_n305_), .Y(new_new_n307_));
  AN2        g0285(.A(i_3_), .B(i_10_), .Y(new_new_n308_));
  NA4        g0286(.A(new_new_n308_), .B(new_new_n197_), .C(new_new_n177_), .D(new_new_n175_), .Y(new_new_n309_));
  NO2        g0287(.A(i_5_), .B(new_new_n37_), .Y(new_new_n310_));
  NO2        g0288(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n311_));
  OR2        g0289(.A(new_new_n307_), .B(new_new_n304_), .Y(new_new_n312_));
  OAI220     g0290(.A0(new_new_n312_), .A1(i_6_), .B0(new_new_n302_), .B1(new_new_n286_), .Y(new_new_n313_));
  NO4        g0291(.A(new_new_n313_), .B(new_new_n284_), .C(new_new_n215_), .D(new_new_n170_), .Y(new_new_n314_));
  NO3        g0292(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n57_), .B(new_new_n83_), .Y(new_new_n316_));
  NA2        g0294(.A(new_new_n293_), .B(new_new_n316_), .Y(new_new_n317_));
  NO3        g0295(.A(i_6_), .B(new_new_n192_), .C(i_7_), .Y(new_new_n318_));
  NA2        g0296(.A(new_new_n318_), .B(new_new_n197_), .Y(new_new_n319_));
  AOI210     g0297(.A0(new_new_n319_), .A1(new_new_n317_), .B0(new_new_n171_), .Y(new_new_n320_));
  NO2        g0298(.A(i_2_), .B(i_3_), .Y(new_new_n321_));
  OR2        g0299(.A(i_0_), .B(i_5_), .Y(new_new_n322_));
  NA2        g0300(.A(new_new_n219_), .B(new_new_n322_), .Y(new_new_n323_));
  NA4        g0301(.A(new_new_n323_), .B(new_new_n236_), .C(new_new_n321_), .D(i_1_), .Y(new_new_n324_));
  NA3        g0302(.A(new_new_n293_), .B(new_new_n288_), .C(new_new_n113_), .Y(new_new_n325_));
  NO2        g0303(.A(new_new_n159_), .B(new_new_n47_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(i_7_), .C(new_new_n165_), .Y(new_new_n327_));
  NA3        g0305(.A(new_new_n327_), .B(new_new_n325_), .C(new_new_n324_), .Y(new_new_n328_));
  OAI210     g0306(.A0(new_new_n328_), .A1(new_new_n320_), .B0(i_4_), .Y(new_new_n329_));
  NO2        g0307(.A(i_12_), .B(i_10_), .Y(new_new_n330_));
  NOi21      g0308(.An(i_5_), .B(i_0_), .Y(new_new_n331_));
  AOI210     g0309(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n101_), .Y(new_new_n332_));
  NO3        g0310(.A(new_new_n332_), .B(i_4_), .C(new_new_n129_), .Y(new_new_n333_));
  NA4        g0311(.A(new_new_n81_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n334_));
  NA2        g0312(.A(new_new_n333_), .B(new_new_n330_), .Y(new_new_n335_));
  NO2        g0313(.A(i_6_), .B(i_8_), .Y(new_new_n336_));
  NOi21      g0314(.An(i_0_), .B(i_2_), .Y(new_new_n337_));
  AN2        g0315(.A(new_new_n337_), .B(new_new_n336_), .Y(new_new_n338_));
  NO2        g0316(.A(i_1_), .B(i_7_), .Y(new_new_n339_));
  NA3        g0317(.A(new_new_n336_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n340_));
  NA3        g0318(.A(new_new_n340_), .B(new_new_n335_), .C(new_new_n329_), .Y(new_new_n341_));
  NO2        g0319(.A(i_8_), .B(new_new_n323_), .Y(new_new_n342_));
  NOi21      g0320(.An(new_new_n155_), .B(new_new_n104_), .Y(new_new_n343_));
  NO2        g0321(.A(new_new_n343_), .B(new_new_n125_), .Y(new_new_n344_));
  OAI210     g0322(.A0(new_new_n344_), .A1(new_new_n342_), .B0(i_3_), .Y(new_new_n345_));
  INV        g0323(.A(new_new_n81_), .Y(new_new_n346_));
  NO2        g0324(.A(new_new_n297_), .B(new_new_n79_), .Y(new_new_n347_));
  NA2        g0325(.A(new_new_n347_), .B(new_new_n133_), .Y(new_new_n348_));
  NO2        g0326(.A(new_new_n92_), .B(new_new_n192_), .Y(new_new_n349_));
  NA3        g0327(.A(new_new_n306_), .B(new_new_n349_), .C(new_new_n61_), .Y(new_new_n350_));
  AOI210     g0328(.A0(new_new_n350_), .A1(new_new_n348_), .B0(new_new_n346_), .Y(new_new_n351_));
  NO2        g0329(.A(new_new_n192_), .B(i_9_), .Y(new_new_n352_));
  NA2        g0330(.A(new_new_n352_), .B(new_new_n205_), .Y(new_new_n353_));
  NO2        g0331(.A(new_new_n351_), .B(new_new_n296_), .Y(new_new_n354_));
  AOI210     g0332(.A0(new_new_n354_), .A1(new_new_n345_), .B0(new_new_n164_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n341_), .A1(new_new_n315_), .B0(new_new_n355_), .Y(new_new_n356_));
  NOi32      g0334(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n357_));
  INV        g0335(.A(new_new_n357_), .Y(new_new_n358_));
  NAi21      g0336(.An(i_0_), .B(i_6_), .Y(new_new_n359_));
  NAi21      g0337(.An(i_1_), .B(i_5_), .Y(new_new_n360_));
  NA2        g0338(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n25_), .Y(new_new_n362_));
  OAI210     g0340(.A0(new_new_n362_), .A1(new_new_n161_), .B0(new_new_n248_), .Y(new_new_n363_));
  NAi41      g0341(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n364_));
  OAI220     g0342(.A0(new_new_n364_), .A1(new_new_n360_), .B0(new_new_n222_), .B1(new_new_n161_), .Y(new_new_n365_));
  AOI210     g0343(.A0(new_new_n364_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n366_));
  NOi32      g0344(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n367_));
  NAi21      g0345(.An(i_6_), .B(i_1_), .Y(new_new_n368_));
  NA3        g0346(.A(new_new_n368_), .B(new_new_n367_), .C(new_new_n47_), .Y(new_new_n369_));
  NO2        g0347(.A(new_new_n369_), .B(i_0_), .Y(new_new_n370_));
  OR3        g0348(.A(new_new_n370_), .B(new_new_n366_), .C(new_new_n365_), .Y(new_new_n371_));
  NO2        g0349(.A(i_1_), .B(new_new_n101_), .Y(new_new_n372_));
  NAi21      g0350(.An(i_3_), .B(i_4_), .Y(new_new_n373_));
  NO2        g0351(.A(new_new_n373_), .B(i_9_), .Y(new_new_n374_));
  AN2        g0352(.A(i_6_), .B(i_7_), .Y(new_new_n375_));
  OAI210     g0353(.A0(new_new_n375_), .A1(new_new_n372_), .B0(new_new_n374_), .Y(new_new_n376_));
  NA2        g0354(.A(i_2_), .B(i_7_), .Y(new_new_n377_));
  NO2        g0355(.A(new_new_n373_), .B(i_10_), .Y(new_new_n378_));
  NA3        g0356(.A(new_new_n378_), .B(new_new_n377_), .C(new_new_n246_), .Y(new_new_n379_));
  AOI210     g0357(.A0(new_new_n379_), .A1(new_new_n376_), .B0(new_new_n184_), .Y(new_new_n380_));
  AOI210     g0358(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n381_));
  NA2        g0359(.A(new_new_n378_), .B(new_new_n339_), .Y(new_new_n382_));
  NO3        g0360(.A(new_new_n380_), .B(new_new_n371_), .C(new_new_n363_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n383_), .B(new_new_n358_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n385_));
  AN2        g0363(.A(i_12_), .B(i_5_), .Y(new_new_n386_));
  NO2        g0364(.A(i_4_), .B(new_new_n26_), .Y(new_new_n387_));
  NA2        g0365(.A(new_new_n387_), .B(new_new_n386_), .Y(new_new_n388_));
  NO2        g0366(.A(i_11_), .B(i_6_), .Y(new_new_n389_));
  NA3        g0367(.A(new_new_n389_), .B(new_new_n326_), .C(new_new_n227_), .Y(new_new_n390_));
  NO2        g0368(.A(new_new_n390_), .B(new_new_n388_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n244_), .B(i_5_), .Y(new_new_n392_));
  NO2        g0370(.A(i_5_), .B(i_10_), .Y(new_new_n393_));
  NA2        g0371(.A(new_new_n145_), .B(new_new_n46_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n394_), .B(new_new_n1100_), .Y(new_new_n395_));
  OAI210     g0373(.A0(new_new_n395_), .A1(new_new_n391_), .B0(new_new_n385_), .Y(new_new_n396_));
  NO2        g0374(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n397_));
  NO2        g0375(.A(new_new_n151_), .B(new_new_n83_), .Y(new_new_n398_));
  OAI210     g0376(.A0(new_new_n398_), .A1(new_new_n391_), .B0(new_new_n397_), .Y(new_new_n399_));
  NO3        g0377(.A(new_new_n83_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n400_));
  NO2        g0378(.A(i_3_), .B(new_new_n101_), .Y(new_new_n401_));
  NA3        g0379(.A(new_new_n303_), .B(new_new_n73_), .C(new_new_n53_), .Y(new_new_n402_));
  NO2        g0380(.A(i_11_), .B(i_12_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n403_), .B(new_new_n36_), .Y(new_new_n404_));
  NO2        g0382(.A(new_new_n402_), .B(new_new_n404_), .Y(new_new_n405_));
  NA2        g0383(.A(new_new_n393_), .B(new_new_n239_), .Y(new_new_n406_));
  NA3        g0384(.A(new_new_n113_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n222_), .Y(new_new_n408_));
  NAi21      g0386(.An(i_13_), .B(i_0_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n409_), .B(new_new_n241_), .Y(new_new_n410_));
  OAI210     g0388(.A0(new_new_n408_), .A1(new_new_n405_), .B0(new_new_n410_), .Y(new_new_n411_));
  NA3        g0389(.A(new_new_n411_), .B(new_new_n399_), .C(new_new_n396_), .Y(new_new_n412_));
  NO3        g0390(.A(i_1_), .B(i_12_), .C(new_new_n83_), .Y(new_new_n413_));
  NO2        g0391(.A(i_0_), .B(i_11_), .Y(new_new_n414_));
  AN2        g0392(.A(i_1_), .B(i_6_), .Y(new_new_n415_));
  NOi21      g0393(.An(i_2_), .B(i_12_), .Y(new_new_n416_));
  NA2        g0394(.A(new_new_n416_), .B(new_new_n415_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n417_), .B(new_new_n1096_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n143_), .B(i_9_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(i_4_), .Y(new_new_n420_));
  NA2        g0398(.A(new_new_n418_), .B(new_new_n420_), .Y(new_new_n421_));
  NAi21      g0399(.An(i_9_), .B(i_4_), .Y(new_new_n422_));
  OR2        g0400(.A(i_13_), .B(i_10_), .Y(new_new_n423_));
  NO3        g0401(.A(new_new_n423_), .B(new_new_n118_), .C(new_new_n422_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n174_), .B(new_new_n124_), .Y(new_new_n425_));
  BUFFER     g0403(.A(new_new_n217_), .Y(new_new_n426_));
  NO2        g0404(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n285_), .B(new_new_n427_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n278_), .B(new_new_n211_), .Y(new_new_n429_));
  OAI220     g0407(.A0(new_new_n429_), .A1(new_new_n426_), .B0(new_new_n428_), .B1(new_new_n343_), .Y(new_new_n430_));
  INV        g0408(.A(new_new_n430_), .Y(new_new_n431_));
  AOI210     g0409(.A0(new_new_n431_), .A1(new_new_n421_), .B0(new_new_n26_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n325_), .B(new_new_n324_), .Y(new_new_n433_));
  AOI220     g0411(.A0(new_new_n299_), .A1(new_new_n289_), .B0(new_new_n293_), .B1(new_new_n316_), .Y(new_new_n434_));
  NO2        g0412(.A(new_new_n434_), .B(new_new_n171_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n182_), .B(new_new_n83_), .Y(new_new_n436_));
  AOI220     g0414(.A0(new_new_n436_), .A1(new_new_n298_), .B0(new_new_n280_), .B1(new_new_n211_), .Y(new_new_n437_));
  NO2        g0415(.A(new_new_n437_), .B(new_new_n287_), .Y(new_new_n438_));
  NO3        g0416(.A(new_new_n438_), .B(new_new_n435_), .C(new_new_n433_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n195_), .B(new_new_n96_), .Y(new_new_n440_));
  NA3        g0418(.A(new_new_n326_), .B(new_new_n165_), .C(new_new_n83_), .Y(new_new_n441_));
  AOI210     g0419(.A0(new_new_n441_), .A1(new_new_n440_), .B0(i_8_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n192_), .B(i_10_), .Y(new_new_n443_));
  NA3        g0421(.A(new_new_n258_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n444_));
  NA2        g0422(.A(new_new_n299_), .B(new_new_n237_), .Y(new_new_n445_));
  OAI220     g0423(.A0(new_new_n445_), .A1(new_new_n182_), .B0(new_new_n444_), .B1(new_new_n443_), .Y(new_new_n446_));
  NO2        g0424(.A(i_3_), .B(new_new_n49_), .Y(new_new_n447_));
  NA3        g0425(.A(new_new_n339_), .B(new_new_n338_), .C(new_new_n447_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n318_), .B(new_new_n323_), .Y(new_new_n449_));
  OAI210     g0427(.A0(new_new_n449_), .A1(new_new_n188_), .B0(new_new_n448_), .Y(new_new_n450_));
  NO3        g0428(.A(new_new_n450_), .B(new_new_n446_), .C(new_new_n442_), .Y(new_new_n451_));
  AOI210     g0429(.A0(new_new_n451_), .A1(new_new_n439_), .B0(new_new_n272_), .Y(new_new_n452_));
  NO4        g0430(.A(new_new_n452_), .B(new_new_n432_), .C(new_new_n412_), .D(new_new_n384_), .Y(new_new_n453_));
  NO2        g0431(.A(new_new_n61_), .B(i_4_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n71_), .B(i_13_), .Y(new_new_n455_));
  NO2        g0433(.A(i_10_), .B(i_9_), .Y(new_new_n456_));
  NAi21      g0434(.An(i_12_), .B(i_8_), .Y(new_new_n457_));
  NO2        g0435(.A(new_new_n457_), .B(i_3_), .Y(new_new_n458_));
  NA2        g0436(.A(i_2_), .B(new_new_n104_), .Y(new_new_n459_));
  NO2        g0437(.A(new_new_n459_), .B(new_new_n204_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n311_), .B(i_0_), .Y(new_new_n461_));
  NO3        g0439(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n462_));
  NA2        g0440(.A(new_new_n267_), .B(new_new_n97_), .Y(new_new_n463_));
  NA2        g0441(.A(new_new_n463_), .B(new_new_n462_), .Y(new_new_n464_));
  NA2        g0442(.A(i_8_), .B(i_9_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n285_), .B(new_new_n205_), .Y(new_new_n466_));
  OAI220     g0444(.A0(new_new_n466_), .A1(new_new_n465_), .B0(new_new_n464_), .B1(new_new_n461_), .Y(new_new_n467_));
  NO3        g0445(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n468_));
  NA3        g0446(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n469_));
  NO2        g0447(.A(new_new_n467_), .B(new_new_n460_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n298_), .B(new_new_n108_), .Y(new_new_n471_));
  OR2        g0449(.A(new_new_n471_), .B(new_new_n207_), .Y(new_new_n472_));
  BUFFER     g0450(.A(new_new_n353_), .Y(new_new_n473_));
  OA220      g0451(.A0(new_new_n473_), .A1(new_new_n164_), .B0(new_new_n472_), .B1(new_new_n234_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n96_), .B(i_13_), .Y(new_new_n475_));
  NA2        g0453(.A(new_new_n436_), .B(new_new_n385_), .Y(new_new_n476_));
  NO2        g0454(.A(i_2_), .B(i_13_), .Y(new_new_n477_));
  NA3        g0455(.A(new_new_n477_), .B(new_new_n163_), .C(new_new_n99_), .Y(new_new_n478_));
  OAI220     g0456(.A0(new_new_n478_), .A1(new_new_n239_), .B0(new_new_n476_), .B1(new_new_n475_), .Y(new_new_n479_));
  NO3        g0457(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n480_));
  NO2        g0458(.A(i_6_), .B(i_7_), .Y(new_new_n481_));
  NO2        g0459(.A(i_11_), .B(i_1_), .Y(new_new_n482_));
  OR2        g0460(.A(i_11_), .B(i_8_), .Y(new_new_n483_));
  NOi21      g0461(.An(i_2_), .B(i_7_), .Y(new_new_n484_));
  NAi31      g0462(.An(new_new_n483_), .B(new_new_n484_), .C(new_new_n1098_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n423_), .B(i_6_), .Y(new_new_n486_));
  NA3        g0464(.A(new_new_n486_), .B(new_new_n454_), .C(new_new_n73_), .Y(new_new_n487_));
  NO2        g0465(.A(new_new_n487_), .B(new_new_n485_), .Y(new_new_n488_));
  NO2        g0466(.A(i_3_), .B(new_new_n192_), .Y(new_new_n489_));
  NO2        g0467(.A(i_6_), .B(i_10_), .Y(new_new_n490_));
  NA4        g0468(.A(new_new_n490_), .B(new_new_n315_), .C(new_new_n489_), .D(new_new_n239_), .Y(new_new_n491_));
  NO2        g0469(.A(new_new_n491_), .B(new_new_n157_), .Y(new_new_n492_));
  NA3        g0470(.A(new_new_n247_), .B(new_new_n173_), .C(new_new_n133_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n159_), .B(i_3_), .Y(new_new_n495_));
  NA3        g0473(.A(new_new_n397_), .B(new_new_n180_), .C(new_new_n150_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n496_), .B(new_new_n493_), .Y(new_new_n497_));
  NO4        g0475(.A(new_new_n497_), .B(new_new_n492_), .C(new_new_n488_), .D(new_new_n479_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n468_), .B(new_new_n393_), .Y(new_new_n499_));
  NO2        g0477(.A(new_new_n499_), .B(new_new_n226_), .Y(new_new_n500_));
  NAi21      g0478(.An(new_new_n217_), .B(new_new_n403_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n339_), .B(new_new_n219_), .Y(new_new_n502_));
  NO2        g0480(.A(new_new_n26_), .B(i_5_), .Y(new_new_n503_));
  NO2        g0481(.A(i_0_), .B(new_new_n83_), .Y(new_new_n504_));
  NA3        g0482(.A(new_new_n504_), .B(new_new_n503_), .C(new_new_n143_), .Y(new_new_n505_));
  OR3        g0483(.A(i_4_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n506_));
  OAI220     g0484(.A0(new_new_n506_), .A1(new_new_n505_), .B0(new_new_n502_), .B1(new_new_n501_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n27_), .B(i_10_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n315_), .B(new_new_n240_), .Y(new_new_n509_));
  OAI220     g0487(.A0(new_new_n509_), .A1(new_new_n444_), .B0(new_new_n508_), .B1(new_new_n475_), .Y(new_new_n510_));
  NO3        g0488(.A(new_new_n510_), .B(new_new_n507_), .C(new_new_n500_), .Y(new_new_n511_));
  NA4        g0489(.A(new_new_n511_), .B(new_new_n498_), .C(new_new_n474_), .D(new_new_n470_), .Y(new_new_n512_));
  NA3        g0490(.A(new_new_n308_), .B(new_new_n177_), .C(new_new_n175_), .Y(new_new_n513_));
  OAI210     g0491(.A0(new_new_n304_), .A1(new_new_n1101_), .B0(new_new_n513_), .Y(new_new_n514_));
  AN2        g0492(.A(new_new_n289_), .B(new_new_n236_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n515_), .B(new_new_n514_), .Y(new_new_n516_));
  NA2        g0494(.A(new_new_n123_), .B(new_new_n112_), .Y(new_new_n517_));
  AO220      g0495(.A0(new_new_n517_), .A1(new_new_n462_), .B0(new_new_n424_), .B1(i_6_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n315_), .B(new_new_n166_), .Y(new_new_n519_));
  OAI210     g0497(.A0(new_new_n519_), .A1(new_new_n234_), .B0(new_new_n309_), .Y(new_new_n520_));
  AOI220     g0498(.A0(new_new_n520_), .A1(i_7_), .B0(new_new_n518_), .B1(new_new_n311_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n386_), .B(new_new_n227_), .Y(new_new_n522_));
  NA2        g0500(.A(new_new_n357_), .B(new_new_n71_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n375_), .B(new_new_n367_), .Y(new_new_n524_));
  AO210      g0502(.A0(new_new_n523_), .A1(new_new_n522_), .B0(new_new_n524_), .Y(new_new_n525_));
  NO2        g0503(.A(new_new_n36_), .B(i_8_), .Y(new_new_n526_));
  AOI210     g0504(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n424_), .Y(new_new_n527_));
  NA2        g0505(.A(new_new_n527_), .B(new_new_n525_), .Y(new_new_n528_));
  INV        g0506(.A(new_new_n528_), .Y(new_new_n529_));
  OAI210     g0507(.A0(i_8_), .A1(i_5_), .B0(new_new_n135_), .Y(new_new_n530_));
  AOI210     g0508(.A0(new_new_n193_), .A1(i_9_), .B0(new_new_n266_), .Y(new_new_n531_));
  NO2        g0509(.A(new_new_n531_), .B(new_new_n198_), .Y(new_new_n532_));
  OR2        g0510(.A(new_new_n182_), .B(i_4_), .Y(new_new_n533_));
  INV        g0511(.A(new_new_n533_), .Y(new_new_n534_));
  AOI220     g0512(.A0(new_new_n534_), .A1(new_new_n532_), .B0(new_new_n530_), .B1(new_new_n425_), .Y(new_new_n535_));
  NA4        g0513(.A(new_new_n535_), .B(new_new_n529_), .C(new_new_n521_), .D(new_new_n516_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n392_), .B(new_new_n298_), .Y(new_new_n537_));
  OAI210     g0515(.A0(new_new_n388_), .A1(i_2_), .B0(new_new_n537_), .Y(new_new_n538_));
  NO2        g0516(.A(i_12_), .B(new_new_n192_), .Y(new_new_n539_));
  NA2        g0517(.A(new_new_n539_), .B(new_new_n227_), .Y(new_new_n540_));
  NO3        g0518(.A(i_10_), .B(new_new_n540_), .C(new_new_n471_), .Y(new_new_n541_));
  NOi31      g0519(.An(new_new_n318_), .B(new_new_n423_), .C(new_new_n38_), .Y(new_new_n542_));
  OAI210     g0520(.A0(new_new_n542_), .A1(new_new_n541_), .B0(new_new_n538_), .Y(new_new_n543_));
  NO2        g0521(.A(i_8_), .B(i_7_), .Y(new_new_n544_));
  OAI210     g0522(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n545_));
  NA2        g0523(.A(new_new_n545_), .B(new_new_n225_), .Y(new_new_n546_));
  AOI220     g0524(.A0(new_new_n326_), .A1(new_new_n40_), .B0(new_new_n237_), .B1(new_new_n206_), .Y(new_new_n547_));
  OAI220     g0525(.A0(new_new_n547_), .A1(new_new_n533_), .B0(new_new_n546_), .B1(new_new_n244_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n45_), .B(i_10_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n549_), .B(i_6_), .Y(new_new_n550_));
  NA3        g0528(.A(new_new_n550_), .B(new_new_n548_), .C(new_new_n544_), .Y(new_new_n551_));
  AOI220     g0529(.A0(new_new_n436_), .A1(new_new_n326_), .B0(new_new_n249_), .B1(new_new_n246_), .Y(new_new_n552_));
  OAI220     g0530(.A0(new_new_n552_), .A1(i_12_), .B0(new_new_n475_), .B1(new_new_n134_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n553_), .B(new_new_n266_), .Y(new_new_n554_));
  NOi31      g0532(.An(new_new_n293_), .B(new_new_n304_), .C(new_new_n1101_), .Y(new_new_n555_));
  NA3        g0533(.A(new_new_n308_), .B(new_new_n175_), .C(new_new_n96_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n223_), .B(new_new_n45_), .Y(new_new_n557_));
  NO2        g0535(.A(new_new_n159_), .B(i_5_), .Y(new_new_n558_));
  NA2        g0536(.A(new_new_n558_), .B(new_new_n321_), .Y(new_new_n559_));
  OAI210     g0537(.A0(new_new_n559_), .A1(new_new_n557_), .B0(new_new_n556_), .Y(new_new_n560_));
  OAI210     g0538(.A0(new_new_n560_), .A1(new_new_n555_), .B0(new_new_n468_), .Y(new_new_n561_));
  NA4        g0539(.A(new_new_n561_), .B(new_new_n554_), .C(new_new_n551_), .D(new_new_n543_), .Y(new_new_n562_));
  NA3        g0540(.A(new_new_n219_), .B(new_new_n69_), .C(new_new_n45_), .Y(new_new_n563_));
  NA2        g0541(.A(new_new_n285_), .B(new_new_n81_), .Y(new_new_n564_));
  AOI210     g0542(.A0(new_new_n563_), .A1(new_new_n348_), .B0(new_new_n564_), .Y(new_new_n565_));
  NA2        g0543(.A(new_new_n299_), .B(new_new_n289_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n566_), .B(new_new_n174_), .Y(new_new_n567_));
  NA2        g0545(.A(new_new_n225_), .B(new_new_n224_), .Y(new_new_n568_));
  NA2        g0546(.A(new_new_n456_), .B(new_new_n223_), .Y(new_new_n569_));
  NO2        g0547(.A(new_new_n568_), .B(new_new_n569_), .Y(new_new_n570_));
  AOI210     g0548(.A0(new_new_n368_), .A1(new_new_n47_), .B0(new_new_n372_), .Y(new_new_n571_));
  NA2        g0549(.A(i_0_), .B(new_new_n49_), .Y(new_new_n572_));
  NA3        g0550(.A(new_new_n539_), .B(new_new_n276_), .C(new_new_n572_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n571_), .B(new_new_n573_), .Y(new_new_n574_));
  NO4        g0552(.A(new_new_n574_), .B(new_new_n570_), .C(new_new_n567_), .D(new_new_n565_), .Y(new_new_n575_));
  NO4        g0553(.A(new_new_n252_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n576_));
  NO3        g0554(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n235_), .B(new_new_n36_), .Y(new_new_n578_));
  AN2        g0556(.A(new_new_n578_), .B(new_new_n577_), .Y(new_new_n579_));
  OA210      g0557(.A0(new_new_n579_), .A1(new_new_n576_), .B0(new_new_n357_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n423_), .B(i_1_), .Y(new_new_n581_));
  NOi31      g0559(.An(new_new_n581_), .B(new_new_n463_), .C(new_new_n71_), .Y(new_new_n582_));
  AN4        g0560(.A(new_new_n582_), .B(new_new_n420_), .C(new_new_n503_), .D(i_2_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n434_), .B(new_new_n178_), .Y(new_new_n584_));
  NO3        g0562(.A(new_new_n584_), .B(new_new_n583_), .C(new_new_n580_), .Y(new_new_n585_));
  NOi21      g0563(.An(i_10_), .B(i_6_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n587_));
  AOI220     g0565(.A0(new_new_n285_), .A1(new_new_n587_), .B0(new_new_n276_), .B1(new_new_n586_), .Y(new_new_n588_));
  NO2        g0566(.A(new_new_n588_), .B(new_new_n461_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n590_));
  NA2        g0568(.A(new_new_n318_), .B(new_new_n166_), .Y(new_new_n591_));
  AOI220     g0569(.A0(new_new_n591_), .A1(new_new_n445_), .B0(new_new_n174_), .B1(new_new_n181_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n197_), .B(new_new_n37_), .Y(new_new_n593_));
  NOi31      g0571(.An(new_new_n147_), .B(new_new_n593_), .C(new_new_n334_), .Y(new_new_n594_));
  NO3        g0572(.A(new_new_n594_), .B(new_new_n592_), .C(new_new_n589_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n523_), .B(new_new_n382_), .Y(new_new_n596_));
  INV        g0574(.A(new_new_n321_), .Y(new_new_n597_));
  NO2        g0575(.A(i_12_), .B(new_new_n83_), .Y(new_new_n598_));
  NA3        g0576(.A(new_new_n598_), .B(new_new_n276_), .C(new_new_n572_), .Y(new_new_n599_));
  NA3        g0577(.A(new_new_n389_), .B(new_new_n285_), .C(new_new_n219_), .Y(new_new_n600_));
  AOI210     g0578(.A0(new_new_n600_), .A1(new_new_n599_), .B0(new_new_n597_), .Y(new_new_n601_));
  NA2        g0579(.A(new_new_n175_), .B(i_0_), .Y(new_new_n602_));
  NO3        g0580(.A(new_new_n602_), .B(i_8_), .C(new_new_n304_), .Y(new_new_n603_));
  OR2        g0581(.A(i_2_), .B(i_5_), .Y(new_new_n604_));
  OR2        g0582(.A(new_new_n604_), .B(new_new_n415_), .Y(new_new_n605_));
  INV        g0583(.A(new_new_n197_), .Y(new_new_n606_));
  AOI210     g0584(.A0(new_new_n606_), .A1(new_new_n605_), .B0(new_new_n501_), .Y(new_new_n607_));
  NO4        g0585(.A(new_new_n607_), .B(new_new_n603_), .C(new_new_n601_), .D(new_new_n596_), .Y(new_new_n608_));
  NA4        g0586(.A(new_new_n608_), .B(new_new_n595_), .C(new_new_n585_), .D(new_new_n575_), .Y(new_new_n609_));
  NO4        g0587(.A(new_new_n609_), .B(new_new_n562_), .C(new_new_n536_), .D(new_new_n512_), .Y(new_new_n610_));
  NA4        g0588(.A(new_new_n610_), .B(new_new_n453_), .C(new_new_n356_), .D(new_new_n314_), .Y(men7));
  NO2        g0589(.A(new_new_n92_), .B(new_new_n53_), .Y(new_new_n612_));
  NO2        g0590(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n613_));
  NA2        g0591(.A(new_new_n387_), .B(new_new_n613_), .Y(new_new_n614_));
  NA2        g0592(.A(new_new_n490_), .B(new_new_n81_), .Y(new_new_n615_));
  NA2        g0593(.A(i_11_), .B(new_new_n192_), .Y(new_new_n616_));
  NA2        g0594(.A(new_new_n145_), .B(new_new_n616_), .Y(new_new_n617_));
  OAI210     g0595(.A0(new_new_n617_), .A1(new_new_n615_), .B0(new_new_n614_), .Y(new_new_n618_));
  NA3        g0596(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n239_), .B(i_4_), .Y(new_new_n620_));
  NA2        g0598(.A(new_new_n620_), .B(i_8_), .Y(new_new_n621_));
  NA2        g0599(.A(i_2_), .B(new_new_n83_), .Y(new_new_n622_));
  OAI210     g0600(.A0(new_new_n86_), .A1(new_new_n202_), .B0(new_new_n203_), .Y(new_new_n623_));
  NO2        g0601(.A(i_7_), .B(new_new_n37_), .Y(new_new_n624_));
  NA2        g0602(.A(i_4_), .B(i_8_), .Y(new_new_n625_));
  AOI210     g0603(.A0(new_new_n625_), .A1(new_new_n308_), .B0(new_new_n624_), .Y(new_new_n626_));
  OAI220     g0604(.A0(new_new_n626_), .A1(new_new_n622_), .B0(new_new_n623_), .B1(i_13_), .Y(new_new_n627_));
  NO3        g0605(.A(new_new_n627_), .B(new_new_n618_), .C(new_new_n612_), .Y(new_new_n628_));
  INV        g0606(.A(new_new_n163_), .Y(new_new_n629_));
  OR2        g0607(.A(i_6_), .B(i_10_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n630_), .B(new_new_n23_), .Y(new_new_n631_));
  OR3        g0609(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n632_));
  NO3        g0610(.A(new_new_n632_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n633_));
  INV        g0611(.A(new_new_n199_), .Y(new_new_n634_));
  NO2        g0612(.A(new_new_n633_), .B(new_new_n631_), .Y(new_new_n635_));
  OA220      g0613(.A0(new_new_n635_), .A1(new_new_n597_), .B0(new_new_n629_), .B1(new_new_n268_), .Y(new_new_n636_));
  AOI210     g0614(.A0(new_new_n636_), .A1(new_new_n628_), .B0(new_new_n61_), .Y(new_new_n637_));
  NOi21      g0615(.An(i_11_), .B(i_7_), .Y(new_new_n638_));
  AO210      g0616(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n639_));
  NO2        g0617(.A(new_new_n639_), .B(new_new_n638_), .Y(new_new_n640_));
  NA2        g0618(.A(new_new_n640_), .B(new_new_n206_), .Y(new_new_n641_));
  NA3        g0619(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n642_));
  NAi31      g0620(.An(new_new_n642_), .B(new_new_n216_), .C(i_11_), .Y(new_new_n643_));
  AOI210     g0621(.A0(new_new_n643_), .A1(new_new_n641_), .B0(new_new_n61_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n85_), .B(new_new_n61_), .Y(new_new_n645_));
  OR2        g0623(.A(new_new_n645_), .B(new_new_n41_), .Y(new_new_n646_));
  NO3        g0624(.A(new_new_n260_), .B(new_new_n208_), .C(new_new_n616_), .Y(new_new_n647_));
  OAI210     g0625(.A0(new_new_n647_), .A1(new_new_n228_), .B0(new_new_n61_), .Y(new_new_n648_));
  NA2        g0626(.A(new_new_n416_), .B(new_new_n31_), .Y(new_new_n649_));
  OR2        g0627(.A(new_new_n208_), .B(new_new_n108_), .Y(new_new_n650_));
  NA2        g0628(.A(new_new_n650_), .B(new_new_n649_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n61_), .B(i_9_), .Y(new_new_n652_));
  NO2        g0630(.A(new_new_n652_), .B(i_4_), .Y(new_new_n653_));
  NA2        g0631(.A(new_new_n653_), .B(new_new_n651_), .Y(new_new_n654_));
  NO2        g0632(.A(i_1_), .B(i_12_), .Y(new_new_n655_));
  NA3        g0633(.A(new_new_n655_), .B(new_new_n110_), .C(new_new_n24_), .Y(new_new_n656_));
  NA4        g0634(.A(new_new_n656_), .B(new_new_n654_), .C(new_new_n648_), .D(new_new_n646_), .Y(new_new_n657_));
  OAI210     g0635(.A0(new_new_n657_), .A1(new_new_n644_), .B0(i_6_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n642_), .B(new_new_n108_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n659_), .B(new_new_n598_), .Y(new_new_n660_));
  NO2        g0638(.A(i_6_), .B(i_11_), .Y(new_new_n661_));
  NA2        g0639(.A(new_new_n660_), .B(new_new_n464_), .Y(new_new_n662_));
  NO4        g0640(.A(new_new_n216_), .B(new_new_n129_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n663_), .B(new_new_n652_), .Y(new_new_n664_));
  NO3        g0642(.A(new_new_n630_), .B(new_new_n235_), .C(new_new_n23_), .Y(new_new_n665_));
  AOI210     g0643(.A0(i_1_), .A1(new_new_n261_), .B0(new_new_n665_), .Y(new_new_n666_));
  OAI210     g0644(.A0(new_new_n666_), .A1(new_new_n45_), .B0(new_new_n664_), .Y(new_new_n667_));
  NA3        g0645(.A(new_new_n544_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n668_));
  NA2        g0646(.A(new_new_n139_), .B(i_9_), .Y(new_new_n669_));
  NA3        g0647(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n670_));
  NO2        g0648(.A(new_new_n47_), .B(i_1_), .Y(new_new_n671_));
  NA3        g0649(.A(new_new_n671_), .B(new_new_n267_), .C(new_new_n45_), .Y(new_new_n672_));
  OAI220     g0650(.A0(new_new_n672_), .A1(new_new_n670_), .B0(new_new_n669_), .B1(new_new_n1095_), .Y(new_new_n673_));
  NA3        g0651(.A(new_new_n652_), .B(new_new_n321_), .C(i_6_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n23_), .Y(new_new_n675_));
  AOI210     g0653(.A0(new_new_n482_), .A1(new_new_n427_), .B0(new_new_n243_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n676_), .B(new_new_n622_), .Y(new_new_n677_));
  NAi21      g0655(.An(new_new_n668_), .B(new_new_n91_), .Y(new_new_n678_));
  NA2        g0656(.A(new_new_n671_), .B(new_new_n267_), .Y(new_new_n679_));
  NO2        g0657(.A(i_11_), .B(new_new_n37_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n680_), .B(new_new_n24_), .Y(new_new_n681_));
  OAI210     g0659(.A0(new_new_n681_), .A1(new_new_n679_), .B0(new_new_n678_), .Y(new_new_n682_));
  OR4        g0660(.A(new_new_n682_), .B(new_new_n677_), .C(new_new_n675_), .D(new_new_n673_), .Y(new_new_n683_));
  NO3        g0661(.A(new_new_n683_), .B(new_new_n667_), .C(new_new_n662_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n239_), .B(new_new_n101_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n685_), .B(new_new_n638_), .Y(new_new_n686_));
  NA2        g0664(.A(new_new_n686_), .B(i_1_), .Y(new_new_n687_));
  NO2        g0665(.A(new_new_n687_), .B(new_new_n632_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n422_), .B(new_new_n83_), .Y(new_new_n689_));
  NA2        g0667(.A(new_new_n688_), .B(new_new_n47_), .Y(new_new_n690_));
  NA2        g0668(.A(i_3_), .B(new_new_n192_), .Y(new_new_n691_));
  NO2        g0669(.A(new_new_n691_), .B(new_new_n115_), .Y(new_new_n692_));
  AN2        g0670(.A(new_new_n692_), .B(new_new_n550_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n118_), .B(new_new_n37_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n83_), .B(i_9_), .Y(new_new_n695_));
  NO2        g0673(.A(new_new_n695_), .B(new_new_n61_), .Y(new_new_n696_));
  NA2        g0674(.A(i_1_), .B(i_3_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n465_), .B(new_new_n92_), .Y(new_new_n698_));
  INV        g0676(.A(new_new_n698_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n699_), .B(new_new_n697_), .Y(new_new_n700_));
  NO2        g0678(.A(new_new_n700_), .B(new_new_n693_), .Y(new_new_n701_));
  NA4        g0679(.A(new_new_n701_), .B(new_new_n690_), .C(new_new_n684_), .D(new_new_n658_), .Y(new_new_n702_));
  NO3        g0680(.A(new_new_n483_), .B(i_3_), .C(i_7_), .Y(new_new_n703_));
  NOi21      g0681(.An(new_new_n703_), .B(i_10_), .Y(new_new_n704_));
  OA210      g0682(.A0(new_new_n704_), .A1(new_new_n247_), .B0(new_new_n83_), .Y(new_new_n705_));
  NA2        g0683(.A(new_new_n375_), .B(new_new_n374_), .Y(new_new_n706_));
  NA3        g0684(.A(new_new_n490_), .B(new_new_n526_), .C(new_new_n47_), .Y(new_new_n707_));
  NO3        g0685(.A(new_new_n484_), .B(new_new_n625_), .C(new_new_n83_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n708_), .B(new_new_n25_), .Y(new_new_n709_));
  NA3        g0687(.A(new_new_n163_), .B(new_new_n81_), .C(new_new_n83_), .Y(new_new_n710_));
  NA4        g0688(.A(new_new_n710_), .B(new_new_n709_), .C(new_new_n707_), .D(new_new_n706_), .Y(new_new_n711_));
  OAI210     g0689(.A0(new_new_n711_), .A1(new_new_n705_), .B0(i_1_), .Y(new_new_n712_));
  AOI210     g0690(.A0(new_new_n267_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n373_), .B(i_2_), .Y(new_new_n714_));
  NA2        g0692(.A(new_new_n714_), .B(new_new_n713_), .Y(new_new_n715_));
  OAI210     g0693(.A0(new_new_n674_), .A1(new_new_n457_), .B0(new_new_n715_), .Y(new_new_n716_));
  INV        g0694(.A(new_new_n716_), .Y(new_new_n717_));
  AOI210     g0695(.A0(new_new_n717_), .A1(new_new_n712_), .B0(i_13_), .Y(new_new_n718_));
  OR2        g0696(.A(i_11_), .B(i_7_), .Y(new_new_n719_));
  NA3        g0697(.A(new_new_n719_), .B(new_new_n106_), .C(new_new_n139_), .Y(new_new_n720_));
  AOI220     g0698(.A0(new_new_n477_), .A1(new_new_n163_), .B0(i_2_), .B1(new_new_n139_), .Y(new_new_n721_));
  OAI210     g0699(.A0(new_new_n721_), .A1(new_new_n45_), .B0(new_new_n720_), .Y(new_new_n722_));
  AOI210     g0700(.A0(new_new_n670_), .A1(new_new_n53_), .B0(i_12_), .Y(new_new_n723_));
  INV        g0701(.A(new_new_n723_), .Y(new_new_n724_));
  NO2        g0702(.A(new_new_n484_), .B(new_new_n24_), .Y(new_new_n725_));
  AOI220     g0703(.A0(new_new_n725_), .A1(new_new_n689_), .B0(new_new_n247_), .B1(new_new_n132_), .Y(new_new_n726_));
  OAI220     g0704(.A0(new_new_n726_), .A1(new_new_n41_), .B0(new_new_n724_), .B1(new_new_n92_), .Y(new_new_n727_));
  AOI210     g0705(.A0(new_new_n722_), .A1(new_new_n336_), .B0(new_new_n727_), .Y(new_new_n728_));
  AOI220     g0706(.A0(i_12_), .A1(new_new_n70_), .B0(new_new_n389_), .B1(new_new_n671_), .Y(new_new_n729_));
  NO2        g0707(.A(new_new_n729_), .B(new_new_n244_), .Y(new_new_n730_));
  AOI210     g0708(.A0(new_new_n457_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n731_));
  NOi31      g0709(.An(new_new_n731_), .B(new_new_n615_), .C(new_new_n45_), .Y(new_new_n732_));
  NA2        g0710(.A(new_new_n128_), .B(i_13_), .Y(new_new_n733_));
  NO2        g0711(.A(new_new_n670_), .B(new_new_n115_), .Y(new_new_n734_));
  INV        g0712(.A(new_new_n734_), .Y(new_new_n735_));
  OAI220     g0713(.A0(new_new_n735_), .A1(new_new_n69_), .B0(new_new_n733_), .B1(new_new_n713_), .Y(new_new_n736_));
  NO3        g0714(.A(new_new_n69_), .B(new_new_n32_), .C(new_new_n101_), .Y(new_new_n737_));
  NA2        g0715(.A(new_new_n26_), .B(new_new_n192_), .Y(new_new_n738_));
  NA2        g0716(.A(new_new_n738_), .B(i_7_), .Y(new_new_n739_));
  NO3        g0717(.A(new_new_n484_), .B(new_new_n239_), .C(new_new_n83_), .Y(new_new_n740_));
  AOI210     g0718(.A0(new_new_n740_), .A1(new_new_n739_), .B0(new_new_n737_), .Y(new_new_n741_));
  AOI220     g0719(.A0(new_new_n389_), .A1(new_new_n671_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n742_));
  OAI220     g0720(.A0(new_new_n742_), .A1(new_new_n621_), .B0(new_new_n741_), .B1(new_new_n634_), .Y(new_new_n743_));
  NO4        g0721(.A(new_new_n743_), .B(new_new_n736_), .C(new_new_n732_), .D(new_new_n730_), .Y(new_new_n744_));
  OR2        g0722(.A(i_11_), .B(i_6_), .Y(new_new_n745_));
  NA3        g0723(.A(new_new_n620_), .B(new_new_n738_), .C(i_7_), .Y(new_new_n746_));
  AOI210     g0724(.A0(new_new_n746_), .A1(new_new_n735_), .B0(new_new_n745_), .Y(new_new_n747_));
  NA3        g0725(.A(new_new_n416_), .B(new_new_n624_), .C(new_new_n97_), .Y(new_new_n748_));
  NA2        g0726(.A(new_new_n661_), .B(i_13_), .Y(new_new_n749_));
  NA2        g0727(.A(new_new_n102_), .B(new_new_n738_), .Y(new_new_n750_));
  NAi21      g0728(.An(i_11_), .B(i_12_), .Y(new_new_n751_));
  NOi41      g0729(.An(new_new_n111_), .B(new_new_n751_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n752_));
  NO3        g0730(.A(new_new_n484_), .B(new_new_n598_), .C(new_new_n625_), .Y(new_new_n753_));
  AOI220     g0731(.A0(new_new_n753_), .A1(new_new_n315_), .B0(new_new_n752_), .B1(new_new_n750_), .Y(new_new_n754_));
  NA3        g0732(.A(new_new_n754_), .B(new_new_n749_), .C(new_new_n748_), .Y(new_new_n755_));
  OAI210     g0733(.A0(new_new_n755_), .A1(new_new_n747_), .B0(new_new_n61_), .Y(new_new_n756_));
  NO2        g0734(.A(i_2_), .B(i_12_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n372_), .B(new_new_n757_), .Y(new_new_n758_));
  NA2        g0736(.A(i_8_), .B(new_new_n25_), .Y(new_new_n759_));
  NO3        g0737(.A(new_new_n759_), .B(new_new_n387_), .C(new_new_n620_), .Y(new_new_n760_));
  NA2        g0738(.A(new_new_n760_), .B(new_new_n372_), .Y(new_new_n761_));
  NO2        g0739(.A(new_new_n129_), .B(i_2_), .Y(new_new_n762_));
  NA2        g0740(.A(new_new_n762_), .B(new_new_n655_), .Y(new_new_n763_));
  NA3        g0741(.A(new_new_n763_), .B(new_new_n761_), .C(new_new_n758_), .Y(new_new_n764_));
  NA3        g0742(.A(new_new_n764_), .B(new_new_n46_), .C(new_new_n227_), .Y(new_new_n765_));
  NA4        g0743(.A(new_new_n765_), .B(new_new_n756_), .C(new_new_n744_), .D(new_new_n728_), .Y(new_new_n766_));
  OR4        g0744(.A(new_new_n766_), .B(new_new_n718_), .C(new_new_n702_), .D(new_new_n637_), .Y(men5));
  AOI210     g0745(.A0(new_new_n686_), .A1(new_new_n270_), .B0(new_new_n425_), .Y(new_new_n768_));
  AN2        g0746(.A(new_new_n24_), .B(i_10_), .Y(new_new_n769_));
  NA3        g0747(.A(new_new_n769_), .B(new_new_n757_), .C(new_new_n108_), .Y(new_new_n770_));
  NO2        g0748(.A(new_new_n621_), .B(i_11_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n86_), .B(new_new_n771_), .Y(new_new_n772_));
  NA3        g0750(.A(new_new_n772_), .B(new_new_n770_), .C(new_new_n768_), .Y(new_new_n773_));
  NO3        g0751(.A(i_11_), .B(new_new_n239_), .C(i_13_), .Y(new_new_n774_));
  NO2        g0752(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n775_));
  NA2        g0753(.A(i_12_), .B(i_8_), .Y(new_new_n776_));
  OAI210     g0754(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n776_), .Y(new_new_n777_));
  INV        g0755(.A(new_new_n456_), .Y(new_new_n778_));
  AOI220     g0756(.A0(new_new_n321_), .A1(new_new_n590_), .B0(new_new_n777_), .B1(new_new_n775_), .Y(new_new_n779_));
  INV        g0757(.A(new_new_n779_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n780_), .B(new_new_n773_), .Y(new_new_n781_));
  INV        g0759(.A(new_new_n173_), .Y(new_new_n782_));
  INV        g0760(.A(new_new_n247_), .Y(new_new_n783_));
  OAI210     g0761(.A0(new_new_n714_), .A1(new_new_n458_), .B0(new_new_n111_), .Y(new_new_n784_));
  AOI210     g0762(.A0(new_new_n784_), .A1(new_new_n783_), .B0(new_new_n782_), .Y(new_new_n785_));
  NO2        g0763(.A(new_new_n465_), .B(new_new_n26_), .Y(new_new_n786_));
  NO2        g0764(.A(new_new_n786_), .B(new_new_n427_), .Y(new_new_n787_));
  NA2        g0765(.A(new_new_n787_), .B(i_2_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n788_), .Y(new_new_n789_));
  AOI210     g0767(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n423_), .Y(new_new_n790_));
  AOI210     g0768(.A0(new_new_n790_), .A1(new_new_n789_), .B0(new_new_n785_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n189_), .B(new_new_n126_), .Y(new_new_n792_));
  OAI210     g0770(.A0(new_new_n792_), .A1(new_new_n775_), .B0(i_2_), .Y(new_new_n793_));
  NO2        g0771(.A(new_new_n793_), .B(new_new_n192_), .Y(new_new_n794_));
  OA210      g0772(.A0(new_new_n640_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n795_));
  NA2        g0773(.A(new_new_n199_), .B(new_new_n202_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n153_), .B(new_new_n616_), .Y(new_new_n797_));
  AOI210     g0775(.A0(new_new_n797_), .A1(new_new_n796_), .B0(new_new_n377_), .Y(new_new_n798_));
  AOI210     g0776(.A0(new_new_n208_), .A1(new_new_n149_), .B0(new_new_n526_), .Y(new_new_n799_));
  NA2        g0777(.A(new_new_n799_), .B(new_new_n427_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n102_), .B(new_new_n45_), .Y(new_new_n801_));
  INV        g0779(.A(new_new_n305_), .Y(new_new_n802_));
  NA4        g0780(.A(new_new_n802_), .B(new_new_n308_), .C(new_new_n125_), .D(new_new_n43_), .Y(new_new_n803_));
  OAI210     g0781(.A0(new_new_n803_), .A1(new_new_n801_), .B0(new_new_n800_), .Y(new_new_n804_));
  NO4        g0782(.A(new_new_n804_), .B(new_new_n798_), .C(new_new_n795_), .D(new_new_n794_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n590_), .B(new_new_n28_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n774_), .B(new_new_n277_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n807_), .B(new_new_n806_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n60_), .B(i_12_), .Y(new_new_n809_));
  NO2        g0787(.A(new_new_n809_), .B(new_new_n127_), .Y(new_new_n810_));
  NO2        g0788(.A(new_new_n810_), .B(new_new_n616_), .Y(new_new_n811_));
  AOI220     g0789(.A0(new_new_n811_), .A1(new_new_n36_), .B0(new_new_n808_), .B1(new_new_n47_), .Y(new_new_n812_));
  NA4        g0790(.A(new_new_n812_), .B(new_new_n805_), .C(new_new_n791_), .D(new_new_n781_), .Y(men6));
  NO3        g0791(.A(new_new_n256_), .B(new_new_n310_), .C(i_1_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n184_), .B(new_new_n140_), .Y(new_new_n815_));
  OAI210     g0793(.A0(new_new_n815_), .A1(new_new_n814_), .B0(new_new_n762_), .Y(new_new_n816_));
  NA3        g0794(.A(new_new_n393_), .B(new_new_n489_), .C(new_new_n69_), .Y(new_new_n817_));
  INV        g0795(.A(new_new_n817_), .Y(new_new_n818_));
  NO2        g0796(.A(new_new_n222_), .B(new_new_n494_), .Y(new_new_n819_));
  NO2        g0797(.A(i_11_), .B(i_9_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n818_), .B(new_new_n331_), .Y(new_new_n821_));
  AO210      g0799(.A0(new_new_n821_), .A1(new_new_n816_), .B0(i_12_), .Y(new_new_n822_));
  NA2        g0800(.A(new_new_n378_), .B(new_new_n339_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n598_), .B(new_new_n61_), .Y(new_new_n824_));
  NA2        g0802(.A(new_new_n704_), .B(new_new_n69_), .Y(new_new_n825_));
  NA4        g0803(.A(new_new_n645_), .B(new_new_n825_), .C(new_new_n824_), .D(new_new_n823_), .Y(new_new_n826_));
  INV        g0804(.A(new_new_n196_), .Y(new_new_n827_));
  AOI220     g0805(.A0(new_new_n827_), .A1(new_new_n820_), .B0(new_new_n826_), .B1(new_new_n71_), .Y(new_new_n828_));
  INV        g0806(.A(new_new_n330_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n73_), .B(new_new_n132_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n830_), .B(new_new_n829_), .Y(new_new_n831_));
  NO3        g0809(.A(new_new_n252_), .B(new_new_n133_), .C(i_9_), .Y(new_new_n832_));
  NA2        g0810(.A(new_new_n832_), .B(new_new_n809_), .Y(new_new_n833_));
  AOI210     g0811(.A0(new_new_n833_), .A1(new_new_n524_), .B0(new_new_n184_), .Y(new_new_n834_));
  NO2        g0812(.A(new_new_n32_), .B(i_11_), .Y(new_new_n835_));
  NA3        g0813(.A(new_new_n835_), .B(new_new_n481_), .C(new_new_n393_), .Y(new_new_n836_));
  NAi32      g0814(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n837_));
  AOI210     g0815(.A0(new_new_n745_), .A1(new_new_n84_), .B0(new_new_n837_), .Y(new_new_n838_));
  OAI210     g0816(.A0(new_new_n703_), .A1(new_new_n578_), .B0(new_new_n577_), .Y(new_new_n839_));
  NAi31      g0817(.An(new_new_n838_), .B(new_new_n839_), .C(new_new_n836_), .Y(new_new_n840_));
  OR3        g0818(.A(new_new_n840_), .B(new_new_n834_), .C(new_new_n831_), .Y(new_new_n841_));
  NO2        g0819(.A(new_new_n719_), .B(i_2_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n843_));
  OAI210     g0821(.A0(new_new_n843_), .A1(new_new_n415_), .B0(new_new_n362_), .Y(new_new_n844_));
  NA2        g0822(.A(new_new_n844_), .B(new_new_n842_), .Y(new_new_n845_));
  AO220      g0823(.A0(new_new_n361_), .A1(new_new_n352_), .B0(new_new_n400_), .B1(new_new_n616_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n846_), .B(new_new_n257_), .C(i_7_), .Y(new_new_n847_));
  OR2        g0825(.A(new_new_n640_), .B(new_new_n458_), .Y(new_new_n848_));
  NA3        g0826(.A(new_new_n848_), .B(new_new_n148_), .C(new_new_n67_), .Y(new_new_n849_));
  AO210      g0827(.A0(new_new_n499_), .A1(new_new_n778_), .B0(new_new_n36_), .Y(new_new_n850_));
  NA4        g0828(.A(new_new_n850_), .B(new_new_n849_), .C(new_new_n847_), .D(new_new_n845_), .Y(new_new_n851_));
  OAI210     g0829(.A0(i_6_), .A1(i_11_), .B0(new_new_n84_), .Y(new_new_n852_));
  AOI220     g0830(.A0(new_new_n852_), .A1(new_new_n577_), .B0(new_new_n819_), .B1(new_new_n739_), .Y(new_new_n853_));
  NA3        g0831(.A(new_new_n377_), .B(new_new_n240_), .C(new_new_n148_), .Y(new_new_n854_));
  NA2        g0832(.A(new_new_n400_), .B(new_new_n68_), .Y(new_new_n855_));
  NA4        g0833(.A(new_new_n855_), .B(new_new_n854_), .C(new_new_n853_), .D(new_new_n623_), .Y(new_new_n856_));
  AO210      g0834(.A0(new_new_n526_), .A1(new_new_n47_), .B0(new_new_n85_), .Y(new_new_n857_));
  NA3        g0835(.A(new_new_n857_), .B(new_new_n490_), .C(new_new_n219_), .Y(new_new_n858_));
  AOI210     g0836(.A0(new_new_n458_), .A1(new_new_n456_), .B0(new_new_n576_), .Y(new_new_n859_));
  NO2        g0837(.A(new_new_n630_), .B(new_new_n102_), .Y(new_new_n860_));
  OAI210     g0838(.A0(new_new_n860_), .A1(new_new_n112_), .B0(new_new_n414_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n246_), .B(new_new_n47_), .Y(new_new_n862_));
  INV        g0840(.A(new_new_n605_), .Y(new_new_n863_));
  NA3        g0841(.A(new_new_n863_), .B(new_new_n330_), .C(i_7_), .Y(new_new_n864_));
  NA4        g0842(.A(new_new_n864_), .B(new_new_n861_), .C(new_new_n859_), .D(new_new_n858_), .Y(new_new_n865_));
  NO4        g0843(.A(new_new_n865_), .B(new_new_n856_), .C(new_new_n851_), .D(new_new_n841_), .Y(new_new_n866_));
  NA4        g0844(.A(new_new_n866_), .B(new_new_n828_), .C(new_new_n822_), .D(new_new_n383_), .Y(men3));
  NA2        g0845(.A(i_12_), .B(i_10_), .Y(new_new_n868_));
  NA2        g0846(.A(i_6_), .B(i_7_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n869_), .B(i_0_), .Y(new_new_n870_));
  NO2        g0848(.A(i_11_), .B(new_new_n239_), .Y(new_new_n871_));
  OAI210     g0849(.A0(new_new_n870_), .A1(new_new_n293_), .B0(new_new_n871_), .Y(new_new_n872_));
  NO2        g0850(.A(new_new_n872_), .B(new_new_n192_), .Y(new_new_n873_));
  NO3        g0851(.A(new_new_n461_), .B(new_new_n89_), .C(new_new_n45_), .Y(new_new_n874_));
  OA210      g0852(.A0(new_new_n874_), .A1(new_new_n873_), .B0(new_new_n175_), .Y(new_new_n875_));
  NA3        g0853(.A(new_new_n854_), .B(new_new_n623_), .C(new_new_n376_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n876_), .B(new_new_n40_), .Y(new_new_n877_));
  NO3        g0855(.A(new_new_n650_), .B(new_new_n465_), .C(new_new_n132_), .Y(new_new_n878_));
  NA2        g0856(.A(new_new_n416_), .B(new_new_n46_), .Y(new_new_n879_));
  AN2        g0857(.A(new_new_n463_), .B(new_new_n54_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n880_), .B(new_new_n878_), .Y(new_new_n881_));
  AOI210     g0859(.A0(new_new_n881_), .A1(new_new_n877_), .B0(new_new_n49_), .Y(new_new_n882_));
  NO4        g0860(.A(new_new_n381_), .B(new_new_n386_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n883_));
  NA2        g0861(.A(new_new_n184_), .B(new_new_n586_), .Y(new_new_n884_));
  NOi21      g0862(.An(new_new_n884_), .B(new_new_n883_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n731_), .B(new_new_n695_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n337_), .B(new_new_n447_), .Y(new_new_n887_));
  OAI220     g0865(.A0(new_new_n887_), .A1(new_new_n886_), .B0(new_new_n885_), .B1(new_new_n61_), .Y(new_new_n888_));
  NOi21      g0866(.An(i_5_), .B(i_9_), .Y(new_new_n889_));
  NA2        g0867(.A(new_new_n889_), .B(new_new_n455_), .Y(new_new_n890_));
  AOI210     g0868(.A0(new_new_n267_), .A1(new_new_n482_), .B0(new_new_n708_), .Y(new_new_n891_));
  NO3        g0869(.A(new_new_n419_), .B(new_new_n267_), .C(new_new_n71_), .Y(new_new_n892_));
  INV        g0870(.A(new_new_n892_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n1101_), .B0(new_new_n891_), .B1(new_new_n890_), .Y(new_new_n894_));
  NO4        g0872(.A(new_new_n894_), .B(new_new_n888_), .C(new_new_n882_), .D(new_new_n875_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n184_), .B(new_new_n24_), .Y(new_new_n896_));
  NO2        g0874(.A(new_new_n694_), .B(new_new_n613_), .Y(new_new_n897_));
  NO2        g0875(.A(new_new_n897_), .B(new_new_n896_), .Y(new_new_n898_));
  NA2        g0876(.A(new_new_n315_), .B(new_new_n130_), .Y(new_new_n899_));
  NAi21      g0877(.An(new_new_n164_), .B(new_new_n447_), .Y(new_new_n900_));
  OAI220     g0878(.A0(new_new_n900_), .A1(new_new_n862_), .B0(new_new_n899_), .B1(new_new_n406_), .Y(new_new_n901_));
  NO2        g0879(.A(new_new_n901_), .B(new_new_n898_), .Y(new_new_n902_));
  NO2        g0880(.A(new_new_n393_), .B(new_new_n297_), .Y(new_new_n903_));
  NA2        g0881(.A(new_new_n903_), .B(new_new_n734_), .Y(new_new_n904_));
  NA2        g0882(.A(new_new_n587_), .B(i_0_), .Y(new_new_n905_));
  NO3        g0883(.A(new_new_n905_), .B(new_new_n388_), .C(new_new_n86_), .Y(new_new_n906_));
  NO4        g0884(.A(new_new_n604_), .B(new_new_n216_), .C(new_new_n423_), .D(new_new_n415_), .Y(new_new_n907_));
  AOI210     g0885(.A0(new_new_n907_), .A1(i_11_), .B0(new_new_n906_), .Y(new_new_n908_));
  INV        g0886(.A(new_new_n481_), .Y(new_new_n909_));
  AN2        g0887(.A(new_new_n96_), .B(new_new_n245_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n774_), .B(new_new_n331_), .Y(new_new_n911_));
  AOI210     g0889(.A0(new_new_n490_), .A1(new_new_n86_), .B0(new_new_n56_), .Y(new_new_n912_));
  OAI220     g0890(.A0(new_new_n912_), .A1(new_new_n911_), .B0(new_new_n681_), .B1(new_new_n546_), .Y(new_new_n913_));
  NO2        g0891(.A(new_new_n254_), .B(new_new_n155_), .Y(new_new_n914_));
  NA2        g0892(.A(i_0_), .B(i_10_), .Y(new_new_n915_));
  NO4        g0893(.A(new_new_n115_), .B(new_new_n56_), .C(new_new_n691_), .D(i_5_), .Y(new_new_n916_));
  AO220      g0894(.A0(new_new_n916_), .A1(new_new_n1097_), .B0(new_new_n914_), .B1(i_6_), .Y(new_new_n917_));
  AOI220     g0895(.A0(new_new_n337_), .A1(new_new_n98_), .B0(new_new_n184_), .B1(new_new_n81_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n581_), .B(i_4_), .Y(new_new_n919_));
  NA2        g0897(.A(new_new_n187_), .B(new_new_n202_), .Y(new_new_n920_));
  OAI220     g0898(.A0(new_new_n920_), .A1(new_new_n911_), .B0(new_new_n919_), .B1(new_new_n918_), .Y(new_new_n921_));
  NO4        g0899(.A(new_new_n921_), .B(new_new_n917_), .C(new_new_n913_), .D(new_new_n910_), .Y(new_new_n922_));
  NA4        g0900(.A(new_new_n922_), .B(new_new_n908_), .C(new_new_n904_), .D(new_new_n902_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n924_));
  NA2        g0902(.A(i_11_), .B(i_9_), .Y(new_new_n925_));
  NO3        g0903(.A(i_12_), .B(new_new_n925_), .C(new_new_n622_), .Y(new_new_n926_));
  AO220      g0904(.A0(new_new_n926_), .A1(new_new_n924_), .B0(new_new_n269_), .B1(new_new_n85_), .Y(new_new_n927_));
  NO2        g0905(.A(new_new_n49_), .B(i_7_), .Y(new_new_n928_));
  NA2        g0906(.A(new_new_n397_), .B(new_new_n180_), .Y(new_new_n929_));
  NA2        g0907(.A(new_new_n929_), .B(new_new_n162_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n925_), .B(new_new_n71_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n176_), .B(i_0_), .Y(new_new_n932_));
  INV        g0910(.A(new_new_n932_), .Y(new_new_n933_));
  NA2        g0911(.A(new_new_n481_), .B(new_new_n233_), .Y(new_new_n934_));
  AOI210     g0912(.A0(new_new_n375_), .A1(new_new_n42_), .B0(new_new_n413_), .Y(new_new_n935_));
  OAI220     g0913(.A0(new_new_n935_), .A1(new_new_n890_), .B0(new_new_n934_), .B1(new_new_n933_), .Y(new_new_n936_));
  NO3        g0914(.A(new_new_n936_), .B(new_new_n930_), .C(new_new_n927_), .Y(new_new_n937_));
  NA2        g0915(.A(new_new_n680_), .B(new_new_n122_), .Y(new_new_n938_));
  NO2        g0916(.A(i_6_), .B(new_new_n938_), .Y(new_new_n939_));
  AOI210     g0917(.A0(new_new_n457_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n173_), .B(new_new_n103_), .Y(new_new_n941_));
  NOi32      g0919(.An(new_new_n940_), .Bn(new_new_n187_), .C(new_new_n941_), .Y(new_new_n942_));
  NO2        g0920(.A(new_new_n1099_), .B(new_new_n879_), .Y(new_new_n943_));
  NO3        g0921(.A(new_new_n943_), .B(new_new_n942_), .C(new_new_n939_), .Y(new_new_n944_));
  NOi21      g0922(.An(i_7_), .B(i_5_), .Y(new_new_n945_));
  NOi31      g0923(.An(new_new_n945_), .B(i_0_), .C(new_new_n751_), .Y(new_new_n946_));
  NA3        g0924(.A(new_new_n946_), .B(new_new_n387_), .C(i_6_), .Y(new_new_n947_));
  OA210      g0925(.A0(new_new_n941_), .A1(new_new_n524_), .B0(new_new_n947_), .Y(new_new_n948_));
  NO3        g0926(.A(new_new_n409_), .B(new_new_n364_), .C(new_new_n360_), .Y(new_new_n949_));
  NO2        g0927(.A(new_new_n264_), .B(new_new_n322_), .Y(new_new_n950_));
  NO2        g0928(.A(new_new_n751_), .B(new_new_n259_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n951_), .A1(new_new_n950_), .B0(new_new_n949_), .Y(new_new_n952_));
  NA4        g0930(.A(new_new_n952_), .B(new_new_n948_), .C(new_new_n944_), .D(new_new_n937_), .Y(new_new_n953_));
  NO2        g0931(.A(new_new_n896_), .B(new_new_n241_), .Y(new_new_n954_));
  AN2        g0932(.A(new_new_n336_), .B(new_new_n331_), .Y(new_new_n955_));
  NA2        g0933(.A(new_new_n954_), .B(i_10_), .Y(new_new_n956_));
  INV        g0934(.A(new_new_n868_), .Y(new_new_n957_));
  OA210      g0935(.A0(new_new_n481_), .A1(new_new_n225_), .B0(new_new_n480_), .Y(new_new_n958_));
  NA2        g0936(.A(new_new_n957_), .B(new_new_n931_), .Y(new_new_n959_));
  NO2        g0937(.A(new_new_n900_), .B(new_new_n909_), .Y(new_new_n960_));
  NO2        g0938(.A(new_new_n257_), .B(new_new_n47_), .Y(new_new_n961_));
  NA2        g0939(.A(new_new_n931_), .B(new_new_n308_), .Y(new_new_n962_));
  OAI210     g0940(.A0(new_new_n961_), .A1(new_new_n186_), .B0(new_new_n962_), .Y(new_new_n963_));
  AOI220     g0941(.A0(new_new_n963_), .A1(new_new_n481_), .B0(new_new_n960_), .B1(new_new_n71_), .Y(new_new_n964_));
  NA2        g0942(.A(new_new_n92_), .B(new_new_n45_), .Y(new_new_n965_));
  NO2        g0943(.A(new_new_n73_), .B(new_new_n776_), .Y(new_new_n966_));
  AOI220     g0944(.A0(new_new_n966_), .A1(new_new_n965_), .B0(new_new_n175_), .B1(new_new_n613_), .Y(new_new_n967_));
  NO2        g0945(.A(new_new_n967_), .B(new_new_n48_), .Y(new_new_n968_));
  NO3        g0946(.A(new_new_n604_), .B(new_new_n359_), .C(new_new_n24_), .Y(new_new_n969_));
  AOI210     g0947(.A0(new_new_n725_), .A1(new_new_n558_), .B0(new_new_n969_), .Y(new_new_n970_));
  NAi21      g0948(.An(i_9_), .B(i_5_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n971_), .B(new_new_n409_), .Y(new_new_n972_));
  NO2        g0950(.A(new_new_n619_), .B(new_new_n105_), .Y(new_new_n973_));
  AOI220     g0951(.A0(new_new_n973_), .A1(i_0_), .B0(new_new_n972_), .B1(new_new_n640_), .Y(new_new_n974_));
  OAI220     g0952(.A0(new_new_n974_), .A1(new_new_n83_), .B0(new_new_n970_), .B1(new_new_n174_), .Y(new_new_n975_));
  NO3        g0953(.A(new_new_n975_), .B(new_new_n968_), .C(new_new_n528_), .Y(new_new_n976_));
  NA4        g0954(.A(new_new_n976_), .B(new_new_n964_), .C(new_new_n959_), .D(new_new_n956_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n977_), .B(new_new_n953_), .C(new_new_n923_), .Y(new_new_n978_));
  NO2        g0956(.A(i_0_), .B(new_new_n751_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n71_), .B(new_new_n45_), .Y(new_new_n980_));
  NA2        g0958(.A(new_new_n915_), .B(new_new_n980_), .Y(new_new_n981_));
  NO3        g0959(.A(new_new_n105_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n982_));
  AO220      g0960(.A0(new_new_n982_), .A1(new_new_n981_), .B0(new_new_n979_), .B1(new_new_n175_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n824_), .A1(new_new_n706_), .B0(new_new_n941_), .Y(new_new_n984_));
  AOI210     g0962(.A0(new_new_n983_), .A1(new_new_n349_), .B0(new_new_n984_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n762_), .B(new_new_n147_), .Y(new_new_n986_));
  INV        g0964(.A(new_new_n986_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n987_), .B(new_new_n695_), .C(new_new_n71_), .Y(new_new_n988_));
  NO2        g0966(.A(new_new_n839_), .B(new_new_n409_), .Y(new_new_n989_));
  NA3        g0967(.A(new_new_n870_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n990_));
  NA2        g0968(.A(new_new_n871_), .B(i_9_), .Y(new_new_n991_));
  AOI210     g0969(.A0(new_new_n990_), .A1(new_new_n505_), .B0(new_new_n991_), .Y(new_new_n992_));
  OAI210     g0970(.A0(new_new_n246_), .A1(i_9_), .B0(new_new_n232_), .Y(new_new_n993_));
  AOI210     g0971(.A0(new_new_n993_), .A1(new_new_n905_), .B0(new_new_n155_), .Y(new_new_n994_));
  NO3        g0972(.A(new_new_n994_), .B(new_new_n992_), .C(new_new_n989_), .Y(new_new_n995_));
  NA3        g0973(.A(new_new_n995_), .B(new_new_n988_), .C(new_new_n985_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n955_), .B(new_new_n377_), .Y(new_new_n997_));
  AOI210     g0975(.A0(new_new_n304_), .A1(new_new_n164_), .B0(new_new_n997_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n928_), .B(new_new_n495_), .Y(new_new_n1000_));
  AOI210     g0978(.A0(new_new_n999_), .A1(new_new_n164_), .B0(new_new_n1000_), .Y(new_new_n1001_));
  NO2        g0979(.A(new_new_n1001_), .B(new_new_n998_), .Y(new_new_n1002_));
  NA2        g0980(.A(new_new_n582_), .B(new_new_n73_), .Y(new_new_n1003_));
  NO3        g0981(.A(new_new_n210_), .B(new_new_n386_), .C(i_0_), .Y(new_new_n1004_));
  OAI210     g0982(.A0(new_new_n1004_), .A1(new_new_n74_), .B0(i_13_), .Y(new_new_n1005_));
  INV        g0983(.A(new_new_n219_), .Y(new_new_n1006_));
  OAI220     g0984(.A0(new_new_n540_), .A1(new_new_n140_), .B0(i_12_), .B1(new_new_n634_), .Y(new_new_n1007_));
  NA3        g0985(.A(new_new_n1007_), .B(new_new_n401_), .C(new_new_n1006_), .Y(new_new_n1008_));
  NA4        g0986(.A(new_new_n1008_), .B(new_new_n1005_), .C(new_new_n1003_), .D(new_new_n1002_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n244_), .B(new_new_n92_), .Y(new_new_n1010_));
  AOI210     g0988(.A0(new_new_n1010_), .A1(new_new_n979_), .B0(new_new_n109_), .Y(new_new_n1011_));
  AOI220     g0989(.A0(new_new_n945_), .A1(new_new_n495_), .B0(new_new_n870_), .B1(new_new_n165_), .Y(new_new_n1012_));
  NA2        g0990(.A(new_new_n352_), .B(new_new_n177_), .Y(new_new_n1013_));
  OA220      g0991(.A0(new_new_n1013_), .A1(new_new_n1012_), .B0(new_new_n1011_), .B1(i_5_), .Y(new_new_n1014_));
  AOI210     g0992(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n176_), .Y(new_new_n1015_));
  NA2        g0993(.A(new_new_n1015_), .B(new_new_n958_), .Y(new_new_n1016_));
  NA3        g0994(.A(new_new_n631_), .B(new_new_n184_), .C(new_new_n81_), .Y(new_new_n1017_));
  NA2        g0995(.A(new_new_n1017_), .B(new_new_n556_), .Y(new_new_n1018_));
  NA2        g0996(.A(new_new_n493_), .B(new_new_n478_), .Y(new_new_n1019_));
  NO2        g0997(.A(new_new_n1019_), .B(new_new_n1018_), .Y(new_new_n1020_));
  NA3        g0998(.A(new_new_n928_), .B(new_new_n293_), .C(new_new_n232_), .Y(new_new_n1021_));
  INV        g0999(.A(new_new_n1021_), .Y(new_new_n1022_));
  NA3        g1000(.A(new_new_n393_), .B(new_new_n338_), .C(new_new_n223_), .Y(new_new_n1023_));
  INV        g1001(.A(new_new_n1023_), .Y(new_new_n1024_));
  NOi31      g1002(.An(new_new_n392_), .B(new_new_n980_), .C(new_new_n241_), .Y(new_new_n1025_));
  NO3        g1003(.A(new_new_n1025_), .B(new_new_n1024_), .C(new_new_n1022_), .Y(new_new_n1026_));
  NA4        g1004(.A(new_new_n1026_), .B(new_new_n1020_), .C(new_new_n1016_), .D(new_new_n1014_), .Y(new_new_n1027_));
  INV        g1005(.A(new_new_n633_), .Y(new_new_n1028_));
  NO3        g1006(.A(new_new_n1028_), .B(new_new_n572_), .C(new_new_n346_), .Y(new_new_n1029_));
  INV        g1007(.A(new_new_n1029_), .Y(new_new_n1030_));
  NA3        g1008(.A(new_new_n308_), .B(i_5_), .C(new_new_n192_), .Y(new_new_n1031_));
  NAi31      g1009(.An(new_new_n243_), .B(new_new_n1031_), .C(new_new_n244_), .Y(new_new_n1032_));
  NO4        g1010(.A(new_new_n241_), .B(new_new_n210_), .C(i_0_), .D(i_12_), .Y(new_new_n1033_));
  AOI220     g1011(.A0(new_new_n1033_), .A1(new_new_n1032_), .B0(new_new_n818_), .B1(new_new_n177_), .Y(new_new_n1034_));
  AN2        g1012(.A(new_new_n915_), .B(new_new_n155_), .Y(new_new_n1035_));
  NO4        g1013(.A(new_new_n1035_), .B(i_12_), .C(new_new_n668_), .D(new_new_n132_), .Y(new_new_n1036_));
  NA2        g1014(.A(new_new_n1036_), .B(new_new_n219_), .Y(new_new_n1037_));
  NA3        g1015(.A(new_new_n98_), .B(new_new_n586_), .C(i_11_), .Y(new_new_n1038_));
  NO2        g1016(.A(new_new_n1038_), .B(new_new_n157_), .Y(new_new_n1039_));
  NA2        g1017(.A(new_new_n945_), .B(new_new_n477_), .Y(new_new_n1040_));
  OAI220     g1018(.A0(i_7_), .A1(new_new_n1031_), .B0(new_new_n1040_), .B1(new_new_n696_), .Y(new_new_n1041_));
  AOI210     g1019(.A0(new_new_n1041_), .A1(new_new_n932_), .B0(new_new_n1039_), .Y(new_new_n1042_));
  NA4        g1020(.A(new_new_n1042_), .B(new_new_n1037_), .C(new_new_n1034_), .D(new_new_n1030_), .Y(new_new_n1043_));
  NO4        g1021(.A(new_new_n1043_), .B(new_new_n1027_), .C(new_new_n1009_), .D(new_new_n996_), .Y(new_new_n1044_));
  NA2        g1022(.A(new_new_n835_), .B(new_new_n37_), .Y(new_new_n1045_));
  NA3        g1023(.A(new_new_n940_), .B(new_new_n372_), .C(i_5_), .Y(new_new_n1046_));
  NA3        g1024(.A(new_new_n1046_), .B(new_new_n1045_), .C(new_new_n629_), .Y(new_new_n1047_));
  NA2        g1025(.A(new_new_n1047_), .B(new_new_n206_), .Y(new_new_n1048_));
  AN2        g1026(.A(new_new_n719_), .B(new_new_n373_), .Y(new_new_n1049_));
  NA2        g1027(.A(new_new_n185_), .B(new_new_n187_), .Y(new_new_n1050_));
  AO210      g1028(.A0(new_new_n1049_), .A1(new_new_n33_), .B0(new_new_n1050_), .Y(new_new_n1051_));
  OAI210     g1029(.A0(new_new_n633_), .A1(new_new_n631_), .B0(new_new_n321_), .Y(new_new_n1052_));
  NAi31      g1030(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1053_));
  AOI210     g1031(.A0(new_new_n118_), .A1(new_new_n68_), .B0(new_new_n1053_), .Y(new_new_n1054_));
  NO2        g1032(.A(new_new_n1054_), .B(new_new_n665_), .Y(new_new_n1055_));
  NA3        g1033(.A(new_new_n1055_), .B(new_new_n1052_), .C(new_new_n1051_), .Y(new_new_n1056_));
  NO2        g1034(.A(new_new_n469_), .B(new_new_n267_), .Y(new_new_n1057_));
  NO4        g1035(.A(new_new_n235_), .B(new_new_n146_), .C(new_new_n697_), .D(new_new_n37_), .Y(new_new_n1058_));
  NO3        g1036(.A(new_new_n1058_), .B(new_new_n1057_), .C(new_new_n907_), .Y(new_new_n1059_));
  OAI210     g1037(.A0(new_new_n1038_), .A1(new_new_n149_), .B0(new_new_n1059_), .Y(new_new_n1060_));
  AOI210     g1038(.A0(new_new_n1056_), .A1(new_new_n49_), .B0(new_new_n1060_), .Y(new_new_n1061_));
  AOI210     g1039(.A0(new_new_n1061_), .A1(new_new_n1048_), .B0(new_new_n71_), .Y(new_new_n1062_));
  INV        g1040(.A(new_new_n579_), .Y(new_new_n1063_));
  NO2        g1041(.A(new_new_n1063_), .B(new_new_n782_), .Y(new_new_n1064_));
  OAI210     g1042(.A0(new_new_n78_), .A1(new_new_n53_), .B0(new_new_n108_), .Y(new_new_n1065_));
  NA2        g1043(.A(new_new_n1065_), .B(new_new_n74_), .Y(new_new_n1066_));
  AOI210     g1044(.A0(new_new_n1015_), .A1(new_new_n928_), .B0(new_new_n946_), .Y(new_new_n1067_));
  AOI210     g1045(.A0(new_new_n1067_), .A1(new_new_n1066_), .B0(new_new_n697_), .Y(new_new_n1068_));
  NA2        g1046(.A(new_new_n264_), .B(new_new_n55_), .Y(new_new_n1069_));
  AOI220     g1047(.A0(new_new_n1069_), .A1(new_new_n74_), .B0(new_new_n347_), .B1(new_new_n256_), .Y(new_new_n1070_));
  NO2        g1048(.A(new_new_n1070_), .B(new_new_n239_), .Y(new_new_n1071_));
  NA3        g1049(.A(new_new_n96_), .B(new_new_n310_), .C(new_new_n31_), .Y(new_new_n1072_));
  INV        g1050(.A(new_new_n1072_), .Y(new_new_n1073_));
  NO3        g1051(.A(new_new_n1073_), .B(new_new_n1071_), .C(new_new_n1068_), .Y(new_new_n1074_));
  OAI210     g1052(.A0(new_new_n269_), .A1(new_new_n160_), .B0(new_new_n86_), .Y(new_new_n1075_));
  NA3        g1053(.A(new_new_n786_), .B(new_new_n293_), .C(new_new_n78_), .Y(new_new_n1076_));
  AOI210     g1054(.A0(new_new_n1076_), .A1(new_new_n1075_), .B0(i_11_), .Y(new_new_n1077_));
  NA2        g1055(.A(new_new_n625_), .B(new_new_n216_), .Y(new_new_n1078_));
  OAI210     g1056(.A0(new_new_n1078_), .A1(new_new_n940_), .B0(new_new_n206_), .Y(new_new_n1079_));
  NA2        g1057(.A(new_new_n166_), .B(i_5_), .Y(new_new_n1080_));
  AOI210     g1058(.A0(new_new_n1079_), .A1(new_new_n796_), .B0(new_new_n1080_), .Y(new_new_n1081_));
  NO3        g1059(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n1082_));
  OAI210     g1060(.A0(new_new_n950_), .A1(new_new_n310_), .B0(new_new_n1082_), .Y(new_new_n1083_));
  NO2        g1061(.A(new_new_n1083_), .B(new_new_n751_), .Y(new_new_n1084_));
  NO4        g1062(.A(new_new_n971_), .B(new_new_n483_), .C(new_new_n253_), .D(new_new_n252_), .Y(new_new_n1085_));
  NO2        g1063(.A(new_new_n1085_), .B(new_new_n576_), .Y(new_new_n1086_));
  INV        g1064(.A(new_new_n365_), .Y(new_new_n1087_));
  AOI210     g1065(.A0(new_new_n1087_), .A1(new_new_n1086_), .B0(new_new_n41_), .Y(new_new_n1088_));
  NO4        g1066(.A(new_new_n1088_), .B(new_new_n1084_), .C(new_new_n1081_), .D(new_new_n1077_), .Y(new_new_n1089_));
  OAI210     g1067(.A0(new_new_n1074_), .A1(i_4_), .B0(new_new_n1089_), .Y(new_new_n1090_));
  NO3        g1068(.A(new_new_n1090_), .B(new_new_n1064_), .C(new_new_n1062_), .Y(new_new_n1091_));
  NA4        g1069(.A(new_new_n1091_), .B(new_new_n1044_), .C(new_new_n978_), .D(new_new_n895_), .Y(men4));
  INV        g1070(.A(i_2_), .Y(new_new_n1095_));
  INV        g1071(.A(i_5_), .Y(new_new_n1096_));
  INV        g1072(.A(new_new_n915_), .Y(new_new_n1097_));
  INV        g1073(.A(i_3_), .Y(new_new_n1098_));
  INV        g1074(.A(new_new_n331_), .Y(new_new_n1099_));
  INV        g1075(.A(new_new_n393_), .Y(new_new_n1100_));
  INV        g1076(.A(i_5_), .Y(new_new_n1101_));
endmodule


