// Benchmark "top" written by ABC on Fri Jun 21 17:49:22 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n139_,
    new_new_n140_, new_new_n141_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n608_,
    new_new_n609_, new_new_n610_, new_new_n611_, new_new_n612_,
    new_new_n613_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n751_, new_new_n752_, new_new_n753_,
    new_new_n754_, new_new_n755_, new_new_n756_, new_new_n757_,
    new_new_n758_, new_new_n759_, new_new_n760_, new_new_n761_,
    new_new_n762_, new_new_n763_, new_new_n764_, new_new_n765_,
    new_new_n766_, new_new_n767_, new_new_n768_, new_new_n769_,
    new_new_n770_, new_new_n771_, new_new_n772_, new_new_n773_,
    new_new_n774_, new_new_n775_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n797_, new_new_n798_,
    new_new_n799_, new_new_n800_, new_new_n801_, new_new_n802_,
    new_new_n803_, new_new_n804_, new_new_n805_, new_new_n806_,
    new_new_n807_, new_new_n808_, new_new_n809_, new_new_n810_,
    new_new_n811_, new_new_n812_, new_new_n813_, new_new_n814_,
    new_new_n815_, new_new_n816_, new_new_n817_, new_new_n818_,
    new_new_n819_, new_new_n820_, new_new_n821_, new_new_n822_,
    new_new_n823_, new_new_n824_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n848_, new_new_n849_, new_new_n850_, new_new_n851_,
    new_new_n852_, new_new_n853_, new_new_n854_, new_new_n855_,
    new_new_n856_, new_new_n857_, new_new_n858_, new_new_n859_,
    new_new_n860_, new_new_n861_, new_new_n862_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_,
    new_new_n872_, new_new_n873_, new_new_n874_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1074_, new_new_n1075_, new_new_n1076_,
    new_new_n1077_, new_new_n1078_, new_new_n1079_, new_new_n1080_,
    new_new_n1081_, new_new_n1082_, new_new_n1083_, new_new_n1084_,
    new_new_n1085_, new_new_n1086_, new_new_n1087_, new_new_n1088_,
    new_new_n1089_, new_new_n1090_, new_new_n1091_, new_new_n1092_,
    new_new_n1093_, new_new_n1094_, new_new_n1095_, new_new_n1096_,
    new_new_n1097_, new_new_n1098_, new_new_n1099_, new_new_n1103_,
    new_new_n1104_, new_new_n1105_, new_new_n1106_, new_new_n1107_,
    new_new_n1108_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  INV        g0062(.A(i_6_), .Y(new_new_n85_));
  OR4        g0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n86_));
  INV        g0064(.A(new_new_n86_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n63_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  NO3        g0070(.A(new_new_n92_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n93_));
  NO2        g0071(.A(new_new_n93_), .B(new_new_n91_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n1108_), .B0(new_new_n80_), .Y(new_new_n95_));
  AN3        g0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n96_));
  NAi21      g0074(.An(i_6_), .B(i_11_), .Y(new_new_n97_));
  NO2        g0075(.A(i_5_), .B(i_8_), .Y(new_new_n98_));
  NOi21      g0076(.An(new_new_n98_), .B(new_new_n97_), .Y(new_new_n99_));
  AOI220     g0077(.A0(new_new_n99_), .A1(new_new_n62_), .B0(new_new_n96_), .B1(new_new_n32_), .Y(new_new_n100_));
  INV        g0078(.A(i_7_), .Y(new_new_n101_));
  NA2        g0079(.A(new_new_n47_), .B(new_new_n101_), .Y(new_new_n102_));
  NO2        g0080(.A(i_0_), .B(i_5_), .Y(new_new_n103_));
  NO2        g0081(.A(new_new_n103_), .B(new_new_n85_), .Y(new_new_n104_));
  NA2        g0082(.A(i_12_), .B(i_3_), .Y(new_new_n105_));
  INV        g0083(.A(new_new_n105_), .Y(new_new_n106_));
  NA3        g0084(.A(new_new_n106_), .B(new_new_n104_), .C(new_new_n102_), .Y(new_new_n107_));
  NAi21      g0085(.An(i_7_), .B(i_11_), .Y(new_new_n108_));
  NO3        g0086(.A(new_new_n108_), .B(new_new_n89_), .C(new_new_n54_), .Y(new_new_n109_));
  AN2        g0087(.A(i_2_), .B(i_10_), .Y(new_new_n110_));
  NO2        g0088(.A(new_new_n110_), .B(i_7_), .Y(new_new_n111_));
  OR2        g0089(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n112_));
  NO2        g0090(.A(i_8_), .B(new_new_n101_), .Y(new_new_n113_));
  NO3        g0091(.A(new_new_n113_), .B(new_new_n112_), .C(new_new_n111_), .Y(new_new_n114_));
  NA2        g0092(.A(i_12_), .B(i_7_), .Y(new_new_n115_));
  NO2        g0093(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n116_));
  NA2        g0094(.A(new_new_n116_), .B(i_0_), .Y(new_new_n117_));
  NA2        g0095(.A(i_11_), .B(i_12_), .Y(new_new_n118_));
  OAI210     g0096(.A0(new_new_n117_), .A1(new_new_n115_), .B0(new_new_n118_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n119_), .B(new_new_n114_), .Y(new_new_n120_));
  NAi41      g0098(.An(new_new_n109_), .B(new_new_n120_), .C(new_new_n107_), .D(new_new_n100_), .Y(new_new_n121_));
  NOi21      g0099(.An(i_1_), .B(i_5_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(i_11_), .Y(new_new_n123_));
  NA2        g0101(.A(new_new_n101_), .B(new_new_n37_), .Y(new_new_n124_));
  NA2        g0102(.A(i_7_), .B(new_new_n25_), .Y(new_new_n125_));
  NA2        g0103(.A(new_new_n125_), .B(new_new_n124_), .Y(new_new_n126_));
  NO2        g0104(.A(new_new_n126_), .B(new_new_n47_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n128_));
  NAi21      g0106(.An(i_3_), .B(i_8_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n62_), .Y(new_new_n130_));
  NOi31      g0108(.An(new_new_n130_), .B(new_new_n128_), .C(new_new_n127_), .Y(new_new_n131_));
  NO2        g0109(.A(i_1_), .B(new_new_n85_), .Y(new_new_n132_));
  NO2        g0110(.A(i_6_), .B(i_5_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(i_3_), .Y(new_new_n134_));
  AO210      g0112(.A0(new_new_n134_), .A1(new_new_n48_), .B0(new_new_n132_), .Y(new_new_n135_));
  OAI220     g0113(.A0(new_new_n135_), .A1(new_new_n108_), .B0(new_new_n131_), .B1(new_new_n123_), .Y(new_new_n136_));
  NO3        g0114(.A(new_new_n136_), .B(new_new_n121_), .C(new_new_n95_), .Y(new_new_n137_));
  NA3        g0115(.A(new_new_n137_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0116(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n139_));
  NA2        g0117(.A(i_6_), .B(new_new_n25_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(new_new_n139_), .Y(new_new_n141_));
  NA4        g0119(.A(new_new_n141_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0120(.A(i_8_), .B(i_7_), .Y(new_new_n143_));
  NA2        g0121(.A(new_new_n143_), .B(i_6_), .Y(new_new_n144_));
  NO2        g0122(.A(i_12_), .B(i_13_), .Y(new_new_n145_));
  NAi21      g0123(.An(i_5_), .B(i_11_), .Y(new_new_n146_));
  NOi21      g0124(.An(new_new_n145_), .B(new_new_n146_), .Y(new_new_n147_));
  NO2        g0125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NA2        g0126(.A(i_2_), .B(i_3_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(i_4_), .Y(new_new_n150_));
  NA3        g0128(.A(new_new_n150_), .B(new_new_n148_), .C(new_new_n147_), .Y(new_new_n151_));
  OR2        g0129(.A(new_new_n151_), .B(new_new_n25_), .Y(new_new_n152_));
  AN2        g0130(.A(new_new_n145_), .B(new_new_n83_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(new_new_n27_), .Y(new_new_n154_));
  NA2        g0132(.A(i_1_), .B(i_5_), .Y(new_new_n155_));
  NO2        g0133(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n156_));
  NA2        g0134(.A(new_new_n156_), .B(new_new_n36_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n155_), .C(new_new_n154_), .Y(new_new_n158_));
  OR2        g0136(.A(i_0_), .B(i_1_), .Y(new_new_n159_));
  NO3        g0137(.A(new_new_n159_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n160_));
  NAi32      g0138(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n161_));
  NAi21      g0139(.An(new_new_n161_), .B(new_new_n160_), .Y(new_new_n162_));
  NOi21      g0140(.An(i_4_), .B(i_10_), .Y(new_new_n163_));
  NA2        g0141(.A(new_new_n163_), .B(new_new_n40_), .Y(new_new_n164_));
  NO2        g0142(.A(i_3_), .B(i_5_), .Y(new_new_n165_));
  NO3        g0143(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n166_));
  NA2        g0144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  OAI210     g0145(.A0(new_new_n167_), .A1(new_new_n164_), .B0(new_new_n162_), .Y(new_new_n168_));
  NO2        g0146(.A(new_new_n168_), .B(new_new_n158_), .Y(new_new_n169_));
  AOI210     g0147(.A0(new_new_n169_), .A1(new_new_n152_), .B0(new_new_n144_), .Y(new_new_n170_));
  NA3        g0148(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n171_));
  NA2        g0149(.A(i_3_), .B(new_new_n49_), .Y(new_new_n172_));
  NOi21      g0150(.An(i_4_), .B(i_9_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_11_), .B(i_13_), .Y(new_new_n174_));
  NA2        g0152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  OR2        g0153(.A(new_new_n175_), .B(new_new_n172_), .Y(new_new_n176_));
  NO2        g0154(.A(i_4_), .B(i_5_), .Y(new_new_n177_));
  NAi21      g0155(.An(i_12_), .B(i_11_), .Y(new_new_n178_));
  NO2        g0156(.A(new_new_n178_), .B(i_13_), .Y(new_new_n179_));
  NA3        g0157(.A(new_new_n179_), .B(new_new_n177_), .C(new_new_n83_), .Y(new_new_n180_));
  AOI210     g0158(.A0(new_new_n180_), .A1(new_new_n176_), .B0(new_new_n171_), .Y(new_new_n181_));
  NO2        g0159(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n182_));
  NA2        g0160(.A(new_new_n182_), .B(new_new_n47_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n36_), .B(i_5_), .Y(new_new_n184_));
  NAi31      g0162(.An(new_new_n184_), .B(new_new_n153_), .C(i_11_), .Y(new_new_n185_));
  NA2        g0163(.A(i_3_), .B(i_5_), .Y(new_new_n186_));
  OR2        g0164(.A(new_new_n186_), .B(new_new_n175_), .Y(new_new_n187_));
  AOI210     g0165(.A0(new_new_n187_), .A1(new_new_n185_), .B0(new_new_n183_), .Y(new_new_n188_));
  NO2        g0166(.A(new_new_n73_), .B(i_5_), .Y(new_new_n189_));
  NO2        g0167(.A(i_13_), .B(i_10_), .Y(new_new_n190_));
  NA3        g0168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n45_), .Y(new_new_n191_));
  NO2        g0169(.A(i_2_), .B(i_1_), .Y(new_new_n192_));
  NA2        g0170(.A(new_new_n192_), .B(i_3_), .Y(new_new_n193_));
  NAi21      g0171(.An(i_4_), .B(i_12_), .Y(new_new_n194_));
  NO4        g0172(.A(new_new_n194_), .B(new_new_n193_), .C(new_new_n191_), .D(new_new_n25_), .Y(new_new_n195_));
  NO3        g0173(.A(new_new_n195_), .B(new_new_n188_), .C(new_new_n181_), .Y(new_new_n196_));
  INV        g0174(.A(i_8_), .Y(new_new_n197_));
  NO2        g0175(.A(new_new_n197_), .B(i_7_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(i_6_), .Y(new_new_n199_));
  NO3        g0177(.A(i_3_), .B(new_new_n85_), .C(new_new_n49_), .Y(new_new_n200_));
  NA2        g0178(.A(new_new_n200_), .B(new_new_n113_), .Y(new_new_n201_));
  NO3        g0179(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n202_));
  NA3        g0180(.A(new_new_n202_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n203_));
  NO3        g0181(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n204_));
  OAI210     g0182(.A0(new_new_n96_), .A1(i_12_), .B0(new_new_n204_), .Y(new_new_n205_));
  AOI210     g0183(.A0(new_new_n205_), .A1(new_new_n203_), .B0(new_new_n201_), .Y(new_new_n206_));
  NO2        g0184(.A(i_3_), .B(i_8_), .Y(new_new_n207_));
  NO3        g0185(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n208_));
  NA3        g0186(.A(new_new_n208_), .B(new_new_n207_), .C(new_new_n40_), .Y(new_new_n209_));
  NO2        g0187(.A(new_new_n103_), .B(new_new_n58_), .Y(new_new_n210_));
  INV        g0188(.A(new_new_n210_), .Y(new_new_n211_));
  NO2        g0189(.A(i_13_), .B(i_9_), .Y(new_new_n212_));
  NA3        g0190(.A(new_new_n212_), .B(i_6_), .C(new_new_n197_), .Y(new_new_n213_));
  NAi21      g0191(.An(i_12_), .B(i_3_), .Y(new_new_n214_));
  OR2        g0192(.A(new_new_n214_), .B(new_new_n213_), .Y(new_new_n215_));
  NO2        g0193(.A(new_new_n45_), .B(i_5_), .Y(new_new_n216_));
  NO3        g0194(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n217_));
  NA2        g0195(.A(new_new_n217_), .B(i_10_), .Y(new_new_n218_));
  OAI220     g0196(.A0(new_new_n218_), .A1(new_new_n215_), .B0(new_new_n211_), .B1(new_new_n209_), .Y(new_new_n219_));
  AOI210     g0197(.A0(new_new_n219_), .A1(i_7_), .B0(new_new_n206_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n220_), .A1(i_4_), .B0(new_new_n199_), .B1(new_new_n196_), .Y(new_new_n221_));
  NAi21      g0199(.An(i_12_), .B(i_7_), .Y(new_new_n222_));
  NA3        g0200(.A(i_13_), .B(new_new_n197_), .C(i_10_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  NA2        g0202(.A(i_0_), .B(i_5_), .Y(new_new_n225_));
  OAI220     g0203(.A0(new_new_n85_), .A1(new_new_n193_), .B0(new_new_n183_), .B1(new_new_n134_), .Y(new_new_n226_));
  NAi31      g0204(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n36_), .B(i_13_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n229_));
  NA3        g0207(.A(new_new_n229_), .B(i_0_), .C(new_new_n228_), .Y(new_new_n230_));
  INV        g0208(.A(i_13_), .Y(new_new_n231_));
  NO2        g0209(.A(i_12_), .B(new_new_n231_), .Y(new_new_n232_));
  NA3        g0210(.A(new_new_n232_), .B(new_new_n202_), .C(new_new_n200_), .Y(new_new_n233_));
  OAI210     g0211(.A0(new_new_n230_), .A1(new_new_n227_), .B0(new_new_n233_), .Y(new_new_n234_));
  AOI220     g0212(.A0(new_new_n234_), .A1(new_new_n143_), .B0(new_new_n226_), .B1(new_new_n224_), .Y(new_new_n235_));
  NO2        g0213(.A(i_12_), .B(new_new_n37_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n186_), .B(i_4_), .Y(new_new_n237_));
  NA2        g0215(.A(new_new_n237_), .B(new_new_n236_), .Y(new_new_n238_));
  OR2        g0216(.A(i_8_), .B(i_7_), .Y(new_new_n239_));
  NO2        g0217(.A(new_new_n239_), .B(new_new_n85_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n54_), .B(i_1_), .Y(new_new_n241_));
  NA2        g0219(.A(new_new_n241_), .B(new_new_n240_), .Y(new_new_n242_));
  INV        g0220(.A(i_12_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n45_), .B(new_new_n243_), .Y(new_new_n244_));
  NO3        g0222(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n245_));
  NA2        g0223(.A(i_2_), .B(i_1_), .Y(new_new_n246_));
  NO2        g0224(.A(new_new_n242_), .B(new_new_n238_), .Y(new_new_n247_));
  NO3        g0225(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n248_));
  NAi21      g0226(.An(i_4_), .B(i_3_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n249_), .B(new_new_n75_), .Y(new_new_n250_));
  NO2        g0228(.A(i_0_), .B(i_6_), .Y(new_new_n251_));
  NOi41      g0229(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n252_));
  NA2        g0230(.A(new_new_n252_), .B(new_new_n251_), .Y(new_new_n253_));
  NO2        g0231(.A(new_new_n246_), .B(new_new_n186_), .Y(new_new_n254_));
  NAi21      g0232(.An(new_new_n253_), .B(new_new_n254_), .Y(new_new_n255_));
  INV        g0233(.A(new_new_n255_), .Y(new_new_n256_));
  AOI220     g0234(.A0(new_new_n256_), .A1(new_new_n40_), .B0(new_new_n247_), .B1(new_new_n212_), .Y(new_new_n257_));
  NO2        g0235(.A(i_11_), .B(new_new_n231_), .Y(new_new_n258_));
  NOi21      g0236(.An(i_1_), .B(i_6_), .Y(new_new_n259_));
  NAi21      g0237(.An(i_3_), .B(i_7_), .Y(new_new_n260_));
  NO2        g0238(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n261_));
  NO2        g0239(.A(i_12_), .B(i_3_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n73_), .B(i_5_), .Y(new_new_n263_));
  NA2        g0241(.A(i_3_), .B(i_9_), .Y(new_new_n264_));
  NAi21      g0242(.An(i_7_), .B(i_10_), .Y(new_new_n265_));
  NA3        g0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n266_));
  INV        g0244(.A(new_new_n144_), .Y(new_new_n267_));
  NA2        g0245(.A(new_new_n243_), .B(i_13_), .Y(new_new_n268_));
  NO2        g0246(.A(new_new_n268_), .B(new_new_n75_), .Y(new_new_n269_));
  NA2        g0247(.A(new_new_n269_), .B(new_new_n267_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n239_), .B(new_new_n37_), .Y(new_new_n271_));
  NA2        g0249(.A(i_12_), .B(i_6_), .Y(new_new_n272_));
  OR2        g0250(.A(i_13_), .B(i_9_), .Y(new_new_n273_));
  NO3        g0251(.A(new_new_n273_), .B(new_new_n272_), .C(new_new_n49_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n249_), .B(i_2_), .Y(new_new_n275_));
  NA3        g0253(.A(new_new_n275_), .B(new_new_n274_), .C(new_new_n45_), .Y(new_new_n276_));
  NA2        g0254(.A(new_new_n258_), .B(i_9_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n278_));
  OAI210     g0256(.A0(new_new_n278_), .A1(new_new_n277_), .B0(new_new_n276_), .Y(new_new_n279_));
  NA2        g0257(.A(new_new_n156_), .B(new_new_n63_), .Y(new_new_n280_));
  NO3        g0258(.A(i_11_), .B(new_new_n231_), .C(new_new_n25_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n260_), .B(i_8_), .Y(new_new_n282_));
  NO2        g0260(.A(i_6_), .B(new_new_n49_), .Y(new_new_n283_));
  NA3        g0261(.A(new_new_n283_), .B(new_new_n282_), .C(new_new_n281_), .Y(new_new_n284_));
  NO3        g0262(.A(new_new_n26_), .B(new_new_n85_), .C(i_5_), .Y(new_new_n285_));
  NA3        g0263(.A(new_new_n285_), .B(new_new_n271_), .C(new_new_n232_), .Y(new_new_n286_));
  AOI210     g0264(.A0(new_new_n286_), .A1(new_new_n284_), .B0(new_new_n280_), .Y(new_new_n287_));
  AOI210     g0265(.A0(new_new_n279_), .A1(new_new_n271_), .B0(new_new_n287_), .Y(new_new_n288_));
  NA4        g0266(.A(new_new_n288_), .B(new_new_n270_), .C(new_new_n257_), .D(new_new_n235_), .Y(new_new_n289_));
  NO3        g0267(.A(i_12_), .B(new_new_n231_), .C(new_new_n37_), .Y(new_new_n290_));
  INV        g0268(.A(new_new_n290_), .Y(new_new_n291_));
  NA2        g0269(.A(i_8_), .B(new_new_n101_), .Y(new_new_n292_));
  NO3        g0270(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n293_));
  AOI220     g0271(.A0(new_new_n293_), .A1(new_new_n200_), .B0(new_new_n165_), .B1(new_new_n241_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(new_new_n292_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n246_), .B(i_0_), .Y(new_new_n296_));
  AOI220     g0274(.A0(new_new_n296_), .A1(new_new_n198_), .B0(i_1_), .B1(new_new_n143_), .Y(new_new_n297_));
  NA2        g0275(.A(new_new_n283_), .B(new_new_n26_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n298_), .B(new_new_n297_), .Y(new_new_n299_));
  NA2        g0277(.A(i_0_), .B(i_1_), .Y(new_new_n300_));
  NO2        g0278(.A(new_new_n300_), .B(i_2_), .Y(new_new_n301_));
  NO2        g0279(.A(new_new_n59_), .B(i_6_), .Y(new_new_n302_));
  NA3        g0280(.A(new_new_n302_), .B(new_new_n301_), .C(new_new_n165_), .Y(new_new_n303_));
  OAI210     g0281(.A0(new_new_n167_), .A1(new_new_n144_), .B0(new_new_n303_), .Y(new_new_n304_));
  NO3        g0282(.A(new_new_n304_), .B(new_new_n299_), .C(new_new_n295_), .Y(new_new_n305_));
  NO2        g0283(.A(i_3_), .B(i_10_), .Y(new_new_n306_));
  NA3        g0284(.A(new_new_n306_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n307_));
  NO2        g0285(.A(i_2_), .B(new_new_n101_), .Y(new_new_n308_));
  NA2        g0286(.A(i_1_), .B(new_new_n36_), .Y(new_new_n309_));
  NOi21      g0287(.An(new_new_n225_), .B(new_new_n103_), .Y(new_new_n310_));
  NA3        g0288(.A(new_new_n310_), .B(i_1_), .C(new_new_n308_), .Y(new_new_n311_));
  AN2        g0289(.A(i_3_), .B(i_10_), .Y(new_new_n312_));
  NA4        g0290(.A(new_new_n312_), .B(new_new_n202_), .C(new_new_n179_), .D(new_new_n177_), .Y(new_new_n313_));
  NO2        g0291(.A(i_5_), .B(new_new_n37_), .Y(new_new_n314_));
  NO2        g0292(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n315_));
  OR2        g0293(.A(new_new_n311_), .B(new_new_n307_), .Y(new_new_n316_));
  OAI220     g0294(.A0(new_new_n316_), .A1(i_6_), .B0(new_new_n305_), .B1(new_new_n291_), .Y(new_new_n317_));
  NO4        g0295(.A(new_new_n317_), .B(new_new_n289_), .C(new_new_n221_), .D(new_new_n170_), .Y(new_new_n318_));
  NO3        g0296(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n319_));
  NO2        g0297(.A(new_new_n59_), .B(new_new_n85_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n296_), .B(new_new_n320_), .Y(new_new_n321_));
  NO3        g0299(.A(i_6_), .B(new_new_n197_), .C(i_7_), .Y(new_new_n322_));
  NA2        g0300(.A(new_new_n322_), .B(new_new_n202_), .Y(new_new_n323_));
  AOI210     g0301(.A0(new_new_n323_), .A1(new_new_n321_), .B0(new_new_n172_), .Y(new_new_n324_));
  NO2        g0302(.A(i_2_), .B(i_3_), .Y(new_new_n325_));
  OR2        g0303(.A(i_0_), .B(i_5_), .Y(new_new_n326_));
  NA2        g0304(.A(new_new_n225_), .B(new_new_n326_), .Y(new_new_n327_));
  NA4        g0305(.A(new_new_n327_), .B(new_new_n240_), .C(new_new_n325_), .D(i_1_), .Y(new_new_n328_));
  NA3        g0306(.A(new_new_n296_), .B(new_new_n165_), .C(new_new_n113_), .Y(new_new_n329_));
  NAi21      g0307(.An(i_8_), .B(i_7_), .Y(new_new_n330_));
  NO2        g0308(.A(new_new_n330_), .B(i_6_), .Y(new_new_n331_));
  NO2        g0309(.A(new_new_n159_), .B(new_new_n47_), .Y(new_new_n332_));
  NA3        g0310(.A(new_new_n332_), .B(new_new_n331_), .C(new_new_n165_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n333_), .B(new_new_n329_), .C(new_new_n328_), .Y(new_new_n334_));
  OAI210     g0312(.A0(new_new_n334_), .A1(new_new_n324_), .B0(i_4_), .Y(new_new_n335_));
  NO2        g0313(.A(i_12_), .B(i_10_), .Y(new_new_n336_));
  NOi21      g0314(.An(i_5_), .B(i_0_), .Y(new_new_n337_));
  AOI210     g0315(.A0(i_2_), .A1(new_new_n49_), .B0(new_new_n101_), .Y(new_new_n338_));
  NO4        g0316(.A(new_new_n338_), .B(new_new_n309_), .C(new_new_n337_), .D(new_new_n129_), .Y(new_new_n339_));
  NA4        g0317(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n85_), .D(i_8_), .Y(new_new_n340_));
  NA2        g0318(.A(new_new_n339_), .B(new_new_n336_), .Y(new_new_n341_));
  NO2        g0319(.A(i_6_), .B(i_8_), .Y(new_new_n342_));
  NOi21      g0320(.An(i_0_), .B(i_2_), .Y(new_new_n343_));
  AN2        g0321(.A(new_new_n343_), .B(new_new_n342_), .Y(new_new_n344_));
  NO2        g0322(.A(i_1_), .B(i_7_), .Y(new_new_n345_));
  AO220      g0323(.A0(new_new_n345_), .A1(new_new_n344_), .B0(new_new_n331_), .B1(new_new_n241_), .Y(new_new_n346_));
  NA2        g0324(.A(new_new_n346_), .B(new_new_n42_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n347_), .B(new_new_n341_), .C(new_new_n335_), .Y(new_new_n348_));
  NO3        g0326(.A(new_new_n239_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n349_));
  NO3        g0327(.A(new_new_n330_), .B(i_2_), .C(i_1_), .Y(new_new_n350_));
  OAI210     g0328(.A0(new_new_n350_), .A1(new_new_n349_), .B0(i_6_), .Y(new_new_n351_));
  NA3        g0329(.A(new_new_n259_), .B(new_new_n308_), .C(new_new_n197_), .Y(new_new_n352_));
  AOI210     g0330(.A0(new_new_n352_), .A1(new_new_n351_), .B0(new_new_n327_), .Y(new_new_n353_));
  NOi21      g0331(.An(new_new_n155_), .B(new_new_n104_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n354_), .B(new_new_n125_), .Y(new_new_n355_));
  OAI210     g0333(.A0(new_new_n355_), .A1(new_new_n353_), .B0(i_3_), .Y(new_new_n356_));
  INV        g0334(.A(new_new_n84_), .Y(new_new_n357_));
  NO2        g0335(.A(new_new_n300_), .B(new_new_n81_), .Y(new_new_n358_));
  NA2        g0336(.A(new_new_n358_), .B(new_new_n133_), .Y(new_new_n359_));
  NO2        g0337(.A(new_new_n92_), .B(new_new_n197_), .Y(new_new_n360_));
  NA3        g0338(.A(new_new_n310_), .B(new_new_n360_), .C(new_new_n63_), .Y(new_new_n361_));
  AOI210     g0339(.A0(new_new_n361_), .A1(new_new_n359_), .B0(new_new_n357_), .Y(new_new_n362_));
  NO2        g0340(.A(new_new_n197_), .B(i_9_), .Y(new_new_n363_));
  NA2        g0341(.A(new_new_n363_), .B(new_new_n210_), .Y(new_new_n364_));
  NO2        g0342(.A(new_new_n364_), .B(new_new_n47_), .Y(new_new_n365_));
  NO3        g0343(.A(new_new_n365_), .B(new_new_n362_), .C(new_new_n299_), .Y(new_new_n366_));
  AOI210     g0344(.A0(new_new_n366_), .A1(new_new_n356_), .B0(new_new_n164_), .Y(new_new_n367_));
  AOI210     g0345(.A0(new_new_n348_), .A1(new_new_n319_), .B0(new_new_n367_), .Y(new_new_n368_));
  NOi32      g0346(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n369_));
  INV        g0347(.A(new_new_n369_), .Y(new_new_n370_));
  NAi21      g0348(.An(i_0_), .B(i_6_), .Y(new_new_n371_));
  NAi21      g0349(.An(i_1_), .B(i_5_), .Y(new_new_n372_));
  NA2        g0350(.A(new_new_n372_), .B(new_new_n371_), .Y(new_new_n373_));
  NA2        g0351(.A(new_new_n373_), .B(new_new_n25_), .Y(new_new_n374_));
  OAI210     g0352(.A0(new_new_n374_), .A1(new_new_n161_), .B0(new_new_n253_), .Y(new_new_n375_));
  NAi41      g0353(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n376_));
  OAI220     g0354(.A0(new_new_n376_), .A1(new_new_n372_), .B0(new_new_n227_), .B1(new_new_n161_), .Y(new_new_n377_));
  AOI210     g0355(.A0(new_new_n376_), .A1(new_new_n161_), .B0(new_new_n159_), .Y(new_new_n378_));
  NOi32      g0356(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n379_));
  NAi21      g0357(.An(i_6_), .B(i_1_), .Y(new_new_n380_));
  NA3        g0358(.A(new_new_n380_), .B(new_new_n379_), .C(new_new_n47_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n381_), .B(i_0_), .Y(new_new_n382_));
  OR3        g0360(.A(new_new_n382_), .B(new_new_n378_), .C(new_new_n377_), .Y(new_new_n383_));
  NO2        g0361(.A(i_1_), .B(new_new_n101_), .Y(new_new_n384_));
  NAi21      g0362(.An(i_3_), .B(i_4_), .Y(new_new_n385_));
  NO2        g0363(.A(new_new_n385_), .B(i_9_), .Y(new_new_n386_));
  AN2        g0364(.A(i_6_), .B(i_7_), .Y(new_new_n387_));
  OAI210     g0365(.A0(new_new_n387_), .A1(new_new_n384_), .B0(new_new_n386_), .Y(new_new_n388_));
  NA2        g0366(.A(i_2_), .B(i_7_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n385_), .B(i_10_), .Y(new_new_n390_));
  NA3        g0368(.A(new_new_n390_), .B(new_new_n389_), .C(new_new_n251_), .Y(new_new_n391_));
  AOI210     g0369(.A0(new_new_n391_), .A1(new_new_n388_), .B0(new_new_n189_), .Y(new_new_n392_));
  AOI210     g0370(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n393_));
  OAI210     g0371(.A0(new_new_n393_), .A1(new_new_n192_), .B0(new_new_n390_), .Y(new_new_n394_));
  AOI220     g0372(.A0(new_new_n390_), .A1(new_new_n345_), .B0(new_new_n245_), .B1(new_new_n192_), .Y(new_new_n395_));
  AOI210     g0373(.A0(new_new_n395_), .A1(new_new_n394_), .B0(i_5_), .Y(new_new_n396_));
  NO4        g0374(.A(new_new_n396_), .B(new_new_n392_), .C(new_new_n383_), .D(new_new_n375_), .Y(new_new_n397_));
  NO2        g0375(.A(new_new_n397_), .B(new_new_n370_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n399_));
  AN2        g0377(.A(i_12_), .B(i_5_), .Y(new_new_n400_));
  NO2        g0378(.A(i_4_), .B(new_new_n26_), .Y(new_new_n401_));
  NA2        g0379(.A(new_new_n401_), .B(new_new_n400_), .Y(new_new_n402_));
  NO2        g0380(.A(i_11_), .B(i_6_), .Y(new_new_n403_));
  NA3        g0381(.A(new_new_n403_), .B(new_new_n332_), .C(new_new_n231_), .Y(new_new_n404_));
  NO2        g0382(.A(new_new_n404_), .B(new_new_n402_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n249_), .B(i_5_), .Y(new_new_n406_));
  NO2        g0384(.A(i_5_), .B(i_10_), .Y(new_new_n407_));
  AOI220     g0385(.A0(new_new_n407_), .A1(new_new_n275_), .B0(new_new_n406_), .B1(new_new_n202_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n145_), .B(new_new_n46_), .Y(new_new_n409_));
  NO2        g0387(.A(new_new_n409_), .B(new_new_n408_), .Y(new_new_n410_));
  OAI210     g0388(.A0(new_new_n410_), .A1(new_new_n405_), .B0(new_new_n399_), .Y(new_new_n411_));
  NO2        g0389(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n151_), .B(new_new_n85_), .Y(new_new_n413_));
  OAI210     g0391(.A0(new_new_n413_), .A1(new_new_n405_), .B0(new_new_n412_), .Y(new_new_n414_));
  NO3        g0392(.A(new_new_n85_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n415_));
  NO2        g0393(.A(i_11_), .B(i_12_), .Y(new_new_n416_));
  NA2        g0394(.A(new_new_n407_), .B(new_new_n243_), .Y(new_new_n417_));
  NA3        g0395(.A(new_new_n113_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n418_));
  OAI220     g0396(.A0(new_new_n418_), .A1(new_new_n227_), .B0(new_new_n417_), .B1(new_new_n340_), .Y(new_new_n419_));
  NAi21      g0397(.An(i_13_), .B(i_0_), .Y(new_new_n420_));
  NO2        g0398(.A(new_new_n420_), .B(new_new_n246_), .Y(new_new_n421_));
  NA2        g0399(.A(new_new_n419_), .B(new_new_n421_), .Y(new_new_n422_));
  NA3        g0400(.A(new_new_n422_), .B(new_new_n414_), .C(new_new_n411_), .Y(new_new_n423_));
  NA2        g0401(.A(new_new_n45_), .B(new_new_n231_), .Y(new_new_n424_));
  NO2        g0402(.A(i_0_), .B(i_11_), .Y(new_new_n425_));
  INV        g0403(.A(i_5_), .Y(new_new_n426_));
  NOi21      g0404(.An(i_2_), .B(i_12_), .Y(new_new_n427_));
  NA2        g0405(.A(new_new_n427_), .B(i_6_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n428_), .B(new_new_n426_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n143_), .B(i_9_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n430_), .B(i_4_), .Y(new_new_n431_));
  NA2        g0409(.A(new_new_n429_), .B(new_new_n431_), .Y(new_new_n432_));
  OR2        g0410(.A(i_13_), .B(i_10_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n175_), .B(new_new_n124_), .Y(new_new_n434_));
  OR2        g0412(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n101_), .B(new_new_n25_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n290_), .B(new_new_n436_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n283_), .B(new_new_n217_), .Y(new_new_n438_));
  OAI220     g0416(.A0(new_new_n438_), .A1(new_new_n435_), .B0(new_new_n437_), .B1(new_new_n354_), .Y(new_new_n439_));
  INV        g0417(.A(new_new_n439_), .Y(new_new_n440_));
  AOI210     g0418(.A0(new_new_n440_), .A1(new_new_n432_), .B0(new_new_n26_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n329_), .B(new_new_n328_), .Y(new_new_n442_));
  AOI220     g0420(.A0(new_new_n302_), .A1(new_new_n293_), .B0(new_new_n296_), .B1(new_new_n320_), .Y(new_new_n443_));
  NO2        g0421(.A(new_new_n443_), .B(new_new_n172_), .Y(new_new_n444_));
  NO2        g0422(.A(new_new_n186_), .B(new_new_n85_), .Y(new_new_n445_));
  AOI220     g0423(.A0(new_new_n445_), .A1(new_new_n301_), .B0(new_new_n285_), .B1(new_new_n217_), .Y(new_new_n446_));
  NO2        g0424(.A(new_new_n446_), .B(new_new_n292_), .Y(new_new_n447_));
  NO3        g0425(.A(new_new_n447_), .B(new_new_n444_), .C(new_new_n442_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n200_), .B(new_new_n96_), .Y(new_new_n449_));
  NA3        g0427(.A(new_new_n332_), .B(new_new_n165_), .C(new_new_n85_), .Y(new_new_n450_));
  AOI210     g0428(.A0(new_new_n450_), .A1(new_new_n449_), .B0(new_new_n330_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n302_), .B(new_new_n241_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n452_), .B(new_new_n186_), .Y(new_new_n453_));
  NO2        g0431(.A(i_3_), .B(new_new_n49_), .Y(new_new_n454_));
  NA3        g0432(.A(new_new_n345_), .B(new_new_n344_), .C(new_new_n454_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n322_), .B(new_new_n327_), .Y(new_new_n456_));
  OAI210     g0434(.A0(new_new_n456_), .A1(new_new_n193_), .B0(new_new_n455_), .Y(new_new_n457_));
  NO3        g0435(.A(new_new_n457_), .B(new_new_n453_), .C(new_new_n451_), .Y(new_new_n458_));
  AOI210     g0436(.A0(new_new_n458_), .A1(new_new_n448_), .B0(new_new_n277_), .Y(new_new_n459_));
  NO4        g0437(.A(new_new_n459_), .B(new_new_n441_), .C(new_new_n423_), .D(new_new_n398_), .Y(new_new_n460_));
  NO2        g0438(.A(new_new_n63_), .B(i_4_), .Y(new_new_n461_));
  NO2        g0439(.A(new_new_n73_), .B(i_13_), .Y(new_new_n462_));
  NA3        g0440(.A(new_new_n462_), .B(new_new_n461_), .C(i_2_), .Y(new_new_n463_));
  NO2        g0441(.A(i_10_), .B(i_9_), .Y(new_new_n464_));
  NAi21      g0442(.An(i_12_), .B(i_8_), .Y(new_new_n465_));
  NO2        g0443(.A(new_new_n465_), .B(i_3_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n466_), .B(new_new_n464_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n47_), .B(i_4_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n468_), .B(new_new_n104_), .Y(new_new_n469_));
  OAI220     g0447(.A0(new_new_n469_), .A1(new_new_n209_), .B0(new_new_n467_), .B1(new_new_n463_), .Y(new_new_n470_));
  NA2        g0448(.A(new_new_n315_), .B(i_0_), .Y(new_new_n471_));
  NO3        g0449(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n472_));
  NA2        g0450(.A(new_new_n272_), .B(new_new_n97_), .Y(new_new_n473_));
  NA2        g0451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NA2        g0452(.A(i_8_), .B(i_9_), .Y(new_new_n475_));
  NO2        g0453(.A(new_new_n474_), .B(new_new_n471_), .Y(new_new_n476_));
  NA2        g0454(.A(new_new_n258_), .B(new_new_n314_), .Y(new_new_n477_));
  NO3        g0455(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n478_));
  INV        g0456(.A(new_new_n478_), .Y(new_new_n479_));
  NA3        g0457(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n480_));
  NA4        g0458(.A(new_new_n146_), .B(new_new_n116_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n481_));
  OAI220     g0459(.A0(new_new_n481_), .A1(new_new_n480_), .B0(new_new_n479_), .B1(new_new_n477_), .Y(new_new_n482_));
  NO3        g0460(.A(new_new_n482_), .B(new_new_n476_), .C(new_new_n470_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n301_), .B(new_new_n108_), .Y(new_new_n484_));
  OR2        g0462(.A(new_new_n484_), .B(new_new_n213_), .Y(new_new_n485_));
  OR2        g0463(.A(new_new_n364_), .B(new_new_n101_), .Y(new_new_n486_));
  OA220      g0464(.A0(new_new_n486_), .A1(new_new_n164_), .B0(new_new_n485_), .B1(new_new_n238_), .Y(new_new_n487_));
  NA2        g0465(.A(new_new_n96_), .B(i_13_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n445_), .B(new_new_n399_), .Y(new_new_n489_));
  NO2        g0467(.A(i_2_), .B(i_13_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n491_));
  NO3        g0469(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n492_));
  NO2        g0470(.A(i_6_), .B(i_7_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n493_), .B(new_new_n492_), .Y(new_new_n494_));
  NO2        g0472(.A(i_11_), .B(i_1_), .Y(new_new_n495_));
  OR2        g0473(.A(i_11_), .B(i_8_), .Y(new_new_n496_));
  NOi21      g0474(.An(i_2_), .B(i_7_), .Y(new_new_n497_));
  NAi31      g0475(.An(new_new_n496_), .B(new_new_n497_), .C(i_0_), .Y(new_new_n498_));
  NO2        g0476(.A(new_new_n433_), .B(i_6_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n461_), .C(new_new_n75_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n500_), .B(new_new_n498_), .Y(new_new_n501_));
  NO2        g0479(.A(i_3_), .B(new_new_n197_), .Y(new_new_n502_));
  NO2        g0480(.A(i_6_), .B(i_10_), .Y(new_new_n503_));
  NA4        g0481(.A(new_new_n503_), .B(new_new_n319_), .C(new_new_n502_), .D(new_new_n243_), .Y(new_new_n504_));
  NO2        g0482(.A(new_new_n504_), .B(new_new_n157_), .Y(new_new_n505_));
  NA2        g0483(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n506_));
  NO2        g0484(.A(new_new_n159_), .B(i_3_), .Y(new_new_n507_));
  NAi31      g0485(.An(new_new_n506_), .B(new_new_n507_), .C(new_new_n232_), .Y(new_new_n508_));
  NA3        g0486(.A(new_new_n412_), .B(new_new_n182_), .C(new_new_n150_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n509_), .B(new_new_n508_), .Y(new_new_n510_));
  NO4        g0488(.A(new_new_n510_), .B(new_new_n505_), .C(new_new_n501_), .D(new_new_n491_), .Y(new_new_n511_));
  NA2        g0489(.A(new_new_n472_), .B(new_new_n400_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n478_), .B(new_new_n407_), .Y(new_new_n513_));
  NO2        g0491(.A(new_new_n513_), .B(new_new_n230_), .Y(new_new_n514_));
  NAi21      g0492(.An(new_new_n223_), .B(new_new_n416_), .Y(new_new_n515_));
  NA2        g0493(.A(new_new_n345_), .B(new_new_n225_), .Y(new_new_n516_));
  NO2        g0494(.A(new_new_n26_), .B(i_5_), .Y(new_new_n517_));
  NO2        g0495(.A(i_0_), .B(new_new_n85_), .Y(new_new_n518_));
  NA3        g0496(.A(new_new_n518_), .B(new_new_n517_), .C(new_new_n143_), .Y(new_new_n519_));
  OR3        g0497(.A(new_new_n309_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n520_));
  OAI220     g0498(.A0(new_new_n520_), .A1(new_new_n519_), .B0(new_new_n516_), .B1(new_new_n515_), .Y(new_new_n521_));
  NA4        g0499(.A(new_new_n312_), .B(new_new_n229_), .C(new_new_n73_), .D(new_new_n243_), .Y(new_new_n522_));
  NO2        g0500(.A(new_new_n522_), .B(new_new_n494_), .Y(new_new_n523_));
  NO3        g0501(.A(new_new_n523_), .B(new_new_n521_), .C(new_new_n514_), .Y(new_new_n524_));
  NA4        g0502(.A(new_new_n524_), .B(new_new_n511_), .C(new_new_n487_), .D(new_new_n483_), .Y(new_new_n525_));
  NA3        g0503(.A(new_new_n312_), .B(new_new_n179_), .C(new_new_n177_), .Y(new_new_n526_));
  OAI210     g0504(.A0(new_new_n307_), .A1(new_new_n184_), .B0(new_new_n526_), .Y(new_new_n527_));
  AN2        g0505(.A(new_new_n293_), .B(new_new_n240_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n528_), .B(new_new_n527_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n123_), .B(new_new_n112_), .Y(new_new_n530_));
  AN2        g0508(.A(new_new_n530_), .B(new_new_n472_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n319_), .B(new_new_n166_), .Y(new_new_n532_));
  OAI210     g0510(.A0(new_new_n532_), .A1(new_new_n238_), .B0(new_new_n313_), .Y(new_new_n533_));
  AOI220     g0511(.A0(new_new_n533_), .A1(new_new_n331_), .B0(new_new_n531_), .B1(new_new_n315_), .Y(new_new_n534_));
  NA4        g0512(.A(new_new_n462_), .B(new_new_n461_), .C(new_new_n207_), .D(i_2_), .Y(new_new_n535_));
  INV        g0513(.A(new_new_n535_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n369_), .B(new_new_n73_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n387_), .B(new_new_n379_), .Y(new_new_n538_));
  NO2        g0516(.A(new_new_n36_), .B(i_8_), .Y(new_new_n539_));
  NAi41      g0517(.An(new_new_n537_), .B(new_new_n503_), .C(new_new_n539_), .D(new_new_n47_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n39_), .B(i_13_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n541_), .B(new_new_n540_), .Y(new_new_n542_));
  AOI210     g0520(.A0(new_new_n536_), .A1(new_new_n208_), .B0(new_new_n542_), .Y(new_new_n543_));
  NA2        g0521(.A(new_new_n263_), .B(new_new_n64_), .Y(new_new_n544_));
  OAI210     g0522(.A0(i_8_), .A1(new_new_n544_), .B0(new_new_n135_), .Y(new_new_n545_));
  AOI210     g0523(.A0(new_new_n198_), .A1(i_9_), .B0(new_new_n271_), .Y(new_new_n546_));
  NO2        g0524(.A(new_new_n546_), .B(new_new_n203_), .Y(new_new_n547_));
  NO2        g0525(.A(new_new_n186_), .B(new_new_n85_), .Y(new_new_n548_));
  AOI220     g0526(.A0(new_new_n548_), .A1(new_new_n547_), .B0(new_new_n545_), .B1(new_new_n434_), .Y(new_new_n549_));
  NA4        g0527(.A(new_new_n549_), .B(new_new_n543_), .C(new_new_n534_), .D(new_new_n529_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n406_), .B(new_new_n301_), .Y(new_new_n551_));
  OAI210     g0529(.A0(new_new_n402_), .A1(new_new_n171_), .B0(new_new_n551_), .Y(new_new_n552_));
  NO2        g0530(.A(i_12_), .B(new_new_n197_), .Y(new_new_n553_));
  NA2        g0531(.A(new_new_n553_), .B(new_new_n231_), .Y(new_new_n554_));
  NO3        g0532(.A(new_new_n1105_), .B(new_new_n554_), .C(new_new_n484_), .Y(new_new_n555_));
  NOi31      g0533(.An(new_new_n322_), .B(new_new_n433_), .C(new_new_n38_), .Y(new_new_n556_));
  OAI210     g0534(.A0(new_new_n556_), .A1(new_new_n555_), .B0(new_new_n552_), .Y(new_new_n557_));
  NO2        g0535(.A(i_8_), .B(i_7_), .Y(new_new_n558_));
  OAI210     g0536(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n559_), .B(new_new_n229_), .Y(new_new_n560_));
  AOI220     g0538(.A0(new_new_n332_), .A1(new_new_n40_), .B0(new_new_n241_), .B1(new_new_n212_), .Y(new_new_n561_));
  OAI220     g0539(.A0(new_new_n561_), .A1(new_new_n186_), .B0(new_new_n560_), .B1(new_new_n249_), .Y(new_new_n562_));
  NA2        g0540(.A(new_new_n45_), .B(i_10_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n563_), .B(i_6_), .Y(new_new_n564_));
  NA3        g0542(.A(new_new_n564_), .B(new_new_n562_), .C(new_new_n558_), .Y(new_new_n565_));
  AOI220     g0543(.A0(new_new_n445_), .A1(new_new_n332_), .B0(new_new_n254_), .B1(new_new_n251_), .Y(new_new_n566_));
  OAI220     g0544(.A0(new_new_n566_), .A1(new_new_n268_), .B0(new_new_n488_), .B1(new_new_n134_), .Y(new_new_n567_));
  NA2        g0545(.A(new_new_n567_), .B(new_new_n271_), .Y(new_new_n568_));
  NOi31      g0546(.An(new_new_n296_), .B(new_new_n307_), .C(new_new_n184_), .Y(new_new_n569_));
  NA3        g0547(.A(new_new_n312_), .B(new_new_n177_), .C(new_new_n96_), .Y(new_new_n570_));
  NO2        g0548(.A(new_new_n228_), .B(new_new_n45_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n159_), .B(i_5_), .Y(new_new_n572_));
  NA3        g0550(.A(new_new_n572_), .B(new_new_n424_), .C(new_new_n325_), .Y(new_new_n573_));
  OAI210     g0551(.A0(new_new_n573_), .A1(new_new_n571_), .B0(new_new_n570_), .Y(new_new_n574_));
  OAI210     g0552(.A0(new_new_n574_), .A1(new_new_n569_), .B0(new_new_n478_), .Y(new_new_n575_));
  NA4        g0553(.A(new_new_n575_), .B(new_new_n568_), .C(new_new_n565_), .D(new_new_n557_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n290_), .B(new_new_n84_), .Y(new_new_n577_));
  NO2        g0555(.A(new_new_n359_), .B(new_new_n577_), .Y(new_new_n578_));
  NA2        g0556(.A(new_new_n302_), .B(new_new_n293_), .Y(new_new_n579_));
  NO2        g0557(.A(new_new_n579_), .B(new_new_n176_), .Y(new_new_n580_));
  AOI210     g0558(.A0(new_new_n380_), .A1(new_new_n47_), .B0(new_new_n384_), .Y(new_new_n581_));
  NA2        g0559(.A(i_0_), .B(new_new_n49_), .Y(new_new_n582_));
  NA3        g0560(.A(new_new_n553_), .B(new_new_n281_), .C(new_new_n582_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n581_), .B(new_new_n583_), .Y(new_new_n584_));
  NO3        g0562(.A(new_new_n584_), .B(new_new_n580_), .C(new_new_n578_), .Y(new_new_n585_));
  NO4        g0563(.A(new_new_n259_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n586_));
  NO3        g0564(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n239_), .B(new_new_n36_), .Y(new_new_n588_));
  AN2        g0566(.A(new_new_n588_), .B(new_new_n587_), .Y(new_new_n589_));
  OA210      g0567(.A0(new_new_n589_), .A1(new_new_n586_), .B0(new_new_n369_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n433_), .B(i_1_), .Y(new_new_n591_));
  NOi31      g0569(.An(new_new_n591_), .B(new_new_n473_), .C(new_new_n73_), .Y(new_new_n592_));
  AN4        g0570(.A(new_new_n592_), .B(new_new_n431_), .C(new_new_n517_), .D(i_2_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n443_), .B(new_new_n180_), .Y(new_new_n594_));
  NO3        g0572(.A(new_new_n594_), .B(new_new_n593_), .C(new_new_n590_), .Y(new_new_n595_));
  NOi21      g0573(.An(i_10_), .B(i_6_), .Y(new_new_n596_));
  NO2        g0574(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n597_));
  AOI220     g0575(.A0(new_new_n290_), .A1(new_new_n597_), .B0(new_new_n281_), .B1(new_new_n596_), .Y(new_new_n598_));
  NO2        g0576(.A(new_new_n598_), .B(new_new_n471_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n600_));
  NA2        g0578(.A(new_new_n322_), .B(new_new_n166_), .Y(new_new_n601_));
  AOI220     g0579(.A0(new_new_n601_), .A1(new_new_n452_), .B0(new_new_n187_), .B1(new_new_n185_), .Y(new_new_n602_));
  NO2        g0580(.A(new_new_n202_), .B(new_new_n37_), .Y(new_new_n603_));
  NOi31      g0581(.An(new_new_n147_), .B(new_new_n603_), .C(new_new_n340_), .Y(new_new_n604_));
  NO3        g0582(.A(new_new_n604_), .B(new_new_n602_), .C(new_new_n599_), .Y(new_new_n605_));
  NO2        g0583(.A(new_new_n537_), .B(new_new_n395_), .Y(new_new_n606_));
  INV        g0584(.A(new_new_n325_), .Y(new_new_n607_));
  NO2        g0585(.A(i_12_), .B(new_new_n85_), .Y(new_new_n608_));
  NA3        g0586(.A(new_new_n608_), .B(new_new_n281_), .C(new_new_n582_), .Y(new_new_n609_));
  NA3        g0587(.A(new_new_n403_), .B(new_new_n290_), .C(new_new_n225_), .Y(new_new_n610_));
  AOI210     g0588(.A0(new_new_n610_), .A1(new_new_n609_), .B0(new_new_n607_), .Y(new_new_n611_));
  NA2        g0589(.A(new_new_n177_), .B(i_0_), .Y(new_new_n612_));
  NO3        g0590(.A(new_new_n612_), .B(new_new_n351_), .C(new_new_n307_), .Y(new_new_n613_));
  OR2        g0591(.A(i_2_), .B(i_5_), .Y(new_new_n614_));
  OR2        g0592(.A(new_new_n614_), .B(i_6_), .Y(new_new_n615_));
  NO3        g0593(.A(new_new_n613_), .B(new_new_n611_), .C(new_new_n606_), .Y(new_new_n616_));
  NA4        g0594(.A(new_new_n616_), .B(new_new_n605_), .C(new_new_n595_), .D(new_new_n585_), .Y(new_new_n617_));
  NO4        g0595(.A(new_new_n617_), .B(new_new_n576_), .C(new_new_n550_), .D(new_new_n525_), .Y(new_new_n618_));
  NA4        g0596(.A(new_new_n618_), .B(new_new_n460_), .C(new_new_n368_), .D(new_new_n318_), .Y(men7));
  NO2        g0597(.A(new_new_n92_), .B(new_new_n55_), .Y(new_new_n620_));
  NO2        g0598(.A(new_new_n108_), .B(new_new_n89_), .Y(new_new_n621_));
  NA2        g0599(.A(new_new_n401_), .B(new_new_n621_), .Y(new_new_n622_));
  NA2        g0600(.A(new_new_n503_), .B(new_new_n84_), .Y(new_new_n623_));
  NA2        g0601(.A(i_11_), .B(new_new_n197_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n145_), .B(new_new_n624_), .Y(new_new_n625_));
  OAI210     g0603(.A0(new_new_n625_), .A1(new_new_n623_), .B0(new_new_n622_), .Y(new_new_n626_));
  NA3        g0604(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n243_), .B(i_4_), .Y(new_new_n628_));
  NA2        g0606(.A(new_new_n628_), .B(i_8_), .Y(new_new_n629_));
  NO2        g0607(.A(new_new_n105_), .B(new_new_n627_), .Y(new_new_n630_));
  NA2        g0608(.A(i_2_), .B(new_new_n85_), .Y(new_new_n631_));
  OAI210     g0609(.A0(new_new_n88_), .A1(new_new_n207_), .B0(new_new_n208_), .Y(new_new_n632_));
  NO2        g0610(.A(i_7_), .B(new_new_n37_), .Y(new_new_n633_));
  NA2        g0611(.A(i_4_), .B(i_8_), .Y(new_new_n634_));
  AOI210     g0612(.A0(new_new_n634_), .A1(new_new_n312_), .B0(new_new_n633_), .Y(new_new_n635_));
  OAI220     g0613(.A0(new_new_n635_), .A1(new_new_n631_), .B0(new_new_n632_), .B1(i_13_), .Y(new_new_n636_));
  NO4        g0614(.A(new_new_n636_), .B(new_new_n630_), .C(new_new_n626_), .D(new_new_n620_), .Y(new_new_n637_));
  AOI210     g0615(.A0(new_new_n129_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n638_));
  AOI210     g0616(.A0(new_new_n638_), .A1(new_new_n243_), .B0(new_new_n163_), .Y(new_new_n639_));
  OR2        g0617(.A(i_6_), .B(i_10_), .Y(new_new_n640_));
  NO2        g0618(.A(new_new_n640_), .B(new_new_n23_), .Y(new_new_n641_));
  OR3        g0619(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n642_));
  NO3        g0620(.A(new_new_n642_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n643_));
  INV        g0621(.A(new_new_n204_), .Y(new_new_n644_));
  NO2        g0622(.A(new_new_n643_), .B(new_new_n641_), .Y(new_new_n645_));
  OA220      g0623(.A0(new_new_n645_), .A1(new_new_n607_), .B0(new_new_n639_), .B1(new_new_n273_), .Y(new_new_n646_));
  AOI210     g0624(.A0(new_new_n646_), .A1(new_new_n637_), .B0(new_new_n63_), .Y(new_new_n647_));
  NOi21      g0625(.An(i_11_), .B(i_7_), .Y(new_new_n648_));
  AO210      g0626(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n649_));
  NO2        g0627(.A(new_new_n649_), .B(new_new_n648_), .Y(new_new_n650_));
  NA2        g0628(.A(new_new_n650_), .B(new_new_n212_), .Y(new_new_n651_));
  NA3        g0629(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n652_));
  NAi31      g0630(.An(new_new_n652_), .B(new_new_n222_), .C(i_11_), .Y(new_new_n653_));
  AOI210     g0631(.A0(new_new_n653_), .A1(new_new_n651_), .B0(new_new_n63_), .Y(new_new_n654_));
  NA2        g0632(.A(new_new_n87_), .B(new_new_n63_), .Y(new_new_n655_));
  AO210      g0633(.A0(new_new_n655_), .A1(new_new_n395_), .B0(new_new_n41_), .Y(new_new_n656_));
  NO3        g0634(.A(new_new_n265_), .B(new_new_n214_), .C(new_new_n624_), .Y(new_new_n657_));
  OAI210     g0635(.A0(new_new_n657_), .A1(new_new_n232_), .B0(new_new_n63_), .Y(new_new_n658_));
  NA2        g0636(.A(new_new_n427_), .B(new_new_n31_), .Y(new_new_n659_));
  OR2        g0637(.A(new_new_n214_), .B(new_new_n108_), .Y(new_new_n660_));
  NA2        g0638(.A(new_new_n660_), .B(new_new_n659_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n63_), .B(i_9_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n662_), .B(i_4_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n663_), .B(new_new_n661_), .Y(new_new_n664_));
  NO2        g0642(.A(i_1_), .B(i_12_), .Y(new_new_n665_));
  NA3        g0643(.A(new_new_n665_), .B(new_new_n110_), .C(new_new_n24_), .Y(new_new_n666_));
  NA4        g0644(.A(new_new_n666_), .B(new_new_n664_), .C(new_new_n658_), .D(new_new_n656_), .Y(new_new_n667_));
  OAI210     g0645(.A0(new_new_n667_), .A1(new_new_n654_), .B0(i_6_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n243_), .B(new_new_n85_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n669_), .B(i_11_), .Y(new_new_n670_));
  INV        g0648(.A(new_new_n474_), .Y(new_new_n671_));
  NO4        g0649(.A(new_new_n222_), .B(new_new_n129_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n672_));
  NA2        g0650(.A(new_new_n672_), .B(new_new_n662_), .Y(new_new_n673_));
  NA2        g0651(.A(new_new_n243_), .B(i_6_), .Y(new_new_n674_));
  INV        g0652(.A(new_new_n673_), .Y(new_new_n675_));
  NA3        g0653(.A(new_new_n558_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n676_));
  NA2        g0654(.A(new_new_n139_), .B(i_9_), .Y(new_new_n677_));
  NA3        g0655(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n47_), .B(i_1_), .Y(new_new_n679_));
  NA3        g0657(.A(new_new_n679_), .B(new_new_n272_), .C(new_new_n45_), .Y(new_new_n680_));
  OAI220     g0658(.A0(new_new_n680_), .A1(new_new_n678_), .B0(new_new_n677_), .B1(new_new_n1104_), .Y(new_new_n681_));
  NA3        g0659(.A(new_new_n662_), .B(new_new_n325_), .C(i_6_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n682_), .B(new_new_n23_), .Y(new_new_n683_));
  AOI210     g0661(.A0(new_new_n495_), .A1(new_new_n436_), .B0(new_new_n248_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n684_), .B(new_new_n631_), .Y(new_new_n685_));
  NA2        g0663(.A(new_new_n679_), .B(new_new_n272_), .Y(new_new_n686_));
  NO2        g0664(.A(i_11_), .B(new_new_n37_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n687_), .B(new_new_n24_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(new_new_n686_), .Y(new_new_n689_));
  OR4        g0667(.A(new_new_n689_), .B(new_new_n685_), .C(new_new_n683_), .D(new_new_n681_), .Y(new_new_n690_));
  NO3        g0668(.A(new_new_n690_), .B(new_new_n675_), .C(new_new_n671_), .Y(new_new_n691_));
  NO2        g0669(.A(new_new_n243_), .B(new_new_n101_), .Y(new_new_n692_));
  NO2        g0670(.A(new_new_n692_), .B(new_new_n648_), .Y(new_new_n693_));
  NA2        g0671(.A(new_new_n693_), .B(i_1_), .Y(new_new_n694_));
  NO2        g0672(.A(new_new_n694_), .B(new_new_n642_), .Y(new_new_n695_));
  NA2        g0673(.A(new_new_n695_), .B(new_new_n47_), .Y(new_new_n696_));
  NA2        g0674(.A(i_3_), .B(new_new_n197_), .Y(new_new_n697_));
  NO2        g0675(.A(new_new_n697_), .B(new_new_n115_), .Y(new_new_n698_));
  AN2        g0676(.A(new_new_n698_), .B(new_new_n564_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n239_), .B(new_new_n45_), .Y(new_new_n700_));
  NO3        g0678(.A(new_new_n700_), .B(new_new_n315_), .C(new_new_n244_), .Y(new_new_n701_));
  NO2        g0679(.A(new_new_n118_), .B(new_new_n37_), .Y(new_new_n702_));
  NO2        g0680(.A(new_new_n702_), .B(i_6_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n85_), .B(i_9_), .Y(new_new_n704_));
  NO2        g0682(.A(new_new_n704_), .B(new_new_n63_), .Y(new_new_n705_));
  NO2        g0683(.A(new_new_n705_), .B(new_new_n665_), .Y(new_new_n706_));
  NO4        g0684(.A(new_new_n706_), .B(new_new_n703_), .C(new_new_n701_), .D(i_4_), .Y(new_new_n707_));
  NA2        g0685(.A(i_1_), .B(i_3_), .Y(new_new_n708_));
  NO2        g0686(.A(new_new_n475_), .B(new_new_n92_), .Y(new_new_n709_));
  AOI210     g0687(.A0(new_new_n700_), .A1(new_new_n596_), .B0(new_new_n709_), .Y(new_new_n710_));
  NO2        g0688(.A(new_new_n710_), .B(new_new_n708_), .Y(new_new_n711_));
  NO3        g0689(.A(new_new_n711_), .B(new_new_n707_), .C(new_new_n699_), .Y(new_new_n712_));
  NA4        g0690(.A(new_new_n712_), .B(new_new_n696_), .C(new_new_n691_), .D(new_new_n668_), .Y(new_new_n713_));
  NO3        g0691(.A(new_new_n496_), .B(i_3_), .C(i_7_), .Y(new_new_n714_));
  NOi21      g0692(.An(new_new_n714_), .B(i_10_), .Y(new_new_n715_));
  OA210      g0693(.A0(new_new_n715_), .A1(new_new_n252_), .B0(new_new_n85_), .Y(new_new_n716_));
  NA2        g0694(.A(new_new_n387_), .B(new_new_n386_), .Y(new_new_n717_));
  NA3        g0695(.A(new_new_n503_), .B(new_new_n539_), .C(new_new_n47_), .Y(new_new_n718_));
  NO3        g0696(.A(new_new_n497_), .B(new_new_n634_), .C(new_new_n85_), .Y(new_new_n719_));
  NA2        g0697(.A(new_new_n719_), .B(new_new_n25_), .Y(new_new_n720_));
  NA3        g0698(.A(new_new_n163_), .B(new_new_n84_), .C(new_new_n85_), .Y(new_new_n721_));
  NA4        g0699(.A(new_new_n721_), .B(new_new_n720_), .C(new_new_n718_), .D(new_new_n717_), .Y(new_new_n722_));
  OAI210     g0700(.A0(new_new_n722_), .A1(new_new_n716_), .B0(i_1_), .Y(new_new_n723_));
  AOI210     g0701(.A0(new_new_n272_), .A1(new_new_n97_), .B0(i_1_), .Y(new_new_n724_));
  NO2        g0702(.A(new_new_n385_), .B(i_2_), .Y(new_new_n725_));
  NA2        g0703(.A(new_new_n725_), .B(new_new_n724_), .Y(new_new_n726_));
  OAI210     g0704(.A0(new_new_n682_), .A1(new_new_n465_), .B0(new_new_n726_), .Y(new_new_n727_));
  INV        g0705(.A(new_new_n727_), .Y(new_new_n728_));
  AOI210     g0706(.A0(new_new_n728_), .A1(new_new_n723_), .B0(i_13_), .Y(new_new_n729_));
  OR2        g0707(.A(i_11_), .B(i_7_), .Y(new_new_n730_));
  NA3        g0708(.A(new_new_n730_), .B(new_new_n106_), .C(new_new_n139_), .Y(new_new_n731_));
  AOI220     g0709(.A0(new_new_n490_), .A1(new_new_n163_), .B0(new_new_n468_), .B1(new_new_n139_), .Y(new_new_n732_));
  OAI210     g0710(.A0(new_new_n732_), .A1(new_new_n45_), .B0(new_new_n731_), .Y(new_new_n733_));
  AOI210     g0711(.A0(new_new_n678_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n734_));
  NO2        g0712(.A(new_new_n1103_), .B(new_new_n92_), .Y(new_new_n735_));
  AOI210     g0713(.A0(new_new_n733_), .A1(new_new_n342_), .B0(new_new_n735_), .Y(new_new_n736_));
  NA2        g0714(.A(new_new_n115_), .B(new_new_n108_), .Y(new_new_n737_));
  AOI220     g0715(.A0(new_new_n737_), .A1(new_new_n72_), .B0(new_new_n403_), .B1(new_new_n679_), .Y(new_new_n738_));
  NO2        g0716(.A(new_new_n738_), .B(new_new_n249_), .Y(new_new_n739_));
  AOI210     g0717(.A0(new_new_n465_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n740_));
  NOi31      g0718(.An(new_new_n740_), .B(new_new_n623_), .C(new_new_n45_), .Y(new_new_n741_));
  NA2        g0719(.A(new_new_n128_), .B(i_13_), .Y(new_new_n742_));
  NO2        g0720(.A(new_new_n678_), .B(new_new_n115_), .Y(new_new_n743_));
  INV        g0721(.A(new_new_n743_), .Y(new_new_n744_));
  OAI220     g0722(.A0(new_new_n744_), .A1(new_new_n71_), .B0(new_new_n742_), .B1(new_new_n724_), .Y(new_new_n745_));
  NO3        g0723(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n101_), .Y(new_new_n746_));
  NA2        g0724(.A(new_new_n26_), .B(new_new_n197_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n747_), .B(i_7_), .Y(new_new_n748_));
  NO3        g0726(.A(new_new_n497_), .B(new_new_n243_), .C(new_new_n85_), .Y(new_new_n749_));
  AOI210     g0727(.A0(new_new_n749_), .A1(new_new_n748_), .B0(new_new_n746_), .Y(new_new_n750_));
  AOI220     g0728(.A0(new_new_n403_), .A1(new_new_n679_), .B0(new_new_n91_), .B1(new_new_n102_), .Y(new_new_n751_));
  OAI220     g0729(.A0(new_new_n751_), .A1(new_new_n629_), .B0(new_new_n750_), .B1(new_new_n644_), .Y(new_new_n752_));
  NO4        g0730(.A(new_new_n752_), .B(new_new_n745_), .C(new_new_n741_), .D(new_new_n739_), .Y(new_new_n753_));
  OR2        g0731(.A(i_11_), .B(i_6_), .Y(new_new_n754_));
  NA3        g0732(.A(new_new_n628_), .B(new_new_n747_), .C(i_7_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n755_), .A1(new_new_n744_), .B0(new_new_n754_), .Y(new_new_n756_));
  NA3        g0734(.A(new_new_n427_), .B(new_new_n633_), .C(new_new_n97_), .Y(new_new_n757_));
  NA2        g0735(.A(new_new_n670_), .B(i_13_), .Y(new_new_n758_));
  NA2        g0736(.A(new_new_n102_), .B(new_new_n747_), .Y(new_new_n759_));
  NAi21      g0737(.An(i_11_), .B(i_12_), .Y(new_new_n760_));
  NOi41      g0738(.An(new_new_n111_), .B(new_new_n760_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n761_));
  NO3        g0739(.A(new_new_n497_), .B(new_new_n608_), .C(new_new_n634_), .Y(new_new_n762_));
  AOI220     g0740(.A0(new_new_n762_), .A1(new_new_n319_), .B0(new_new_n761_), .B1(new_new_n759_), .Y(new_new_n763_));
  NA3        g0741(.A(new_new_n763_), .B(new_new_n758_), .C(new_new_n757_), .Y(new_new_n764_));
  OAI210     g0742(.A0(new_new_n764_), .A1(new_new_n756_), .B0(new_new_n63_), .Y(new_new_n765_));
  NO2        g0743(.A(i_2_), .B(i_12_), .Y(new_new_n766_));
  NA2        g0744(.A(new_new_n384_), .B(new_new_n766_), .Y(new_new_n767_));
  NA2        g0745(.A(i_8_), .B(new_new_n25_), .Y(new_new_n768_));
  NO3        g0746(.A(new_new_n768_), .B(new_new_n401_), .C(new_new_n628_), .Y(new_new_n769_));
  OAI210     g0747(.A0(new_new_n769_), .A1(new_new_n386_), .B0(new_new_n384_), .Y(new_new_n770_));
  NO2        g0748(.A(new_new_n129_), .B(i_2_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(new_new_n665_), .Y(new_new_n772_));
  NA3        g0750(.A(new_new_n772_), .B(new_new_n770_), .C(new_new_n767_), .Y(new_new_n773_));
  NA3        g0751(.A(new_new_n773_), .B(new_new_n46_), .C(new_new_n231_), .Y(new_new_n774_));
  NA4        g0752(.A(new_new_n774_), .B(new_new_n765_), .C(new_new_n753_), .D(new_new_n736_), .Y(new_new_n775_));
  OR4        g0753(.A(new_new_n775_), .B(new_new_n729_), .C(new_new_n713_), .D(new_new_n647_), .Y(men5));
  AOI210     g0754(.A0(new_new_n693_), .A1(new_new_n275_), .B0(new_new_n434_), .Y(new_new_n777_));
  AN2        g0755(.A(new_new_n24_), .B(i_10_), .Y(new_new_n778_));
  NA3        g0756(.A(new_new_n778_), .B(new_new_n766_), .C(new_new_n108_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n629_), .B(i_11_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n88_), .B(new_new_n780_), .Y(new_new_n781_));
  NA3        g0759(.A(new_new_n781_), .B(new_new_n779_), .C(new_new_n777_), .Y(new_new_n782_));
  NO3        g0760(.A(i_11_), .B(new_new_n243_), .C(i_13_), .Y(new_new_n783_));
  NO2        g0761(.A(new_new_n125_), .B(new_new_n23_), .Y(new_new_n784_));
  NA2        g0762(.A(i_12_), .B(i_8_), .Y(new_new_n785_));
  OAI210     g0763(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n785_), .Y(new_new_n786_));
  INV        g0764(.A(new_new_n464_), .Y(new_new_n787_));
  AOI220     g0765(.A0(new_new_n325_), .A1(new_new_n600_), .B0(new_new_n786_), .B1(new_new_n784_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n788_), .Y(new_new_n789_));
  NO2        g0767(.A(new_new_n789_), .B(new_new_n782_), .Y(new_new_n790_));
  INV        g0768(.A(new_new_n174_), .Y(new_new_n791_));
  INV        g0769(.A(new_new_n252_), .Y(new_new_n792_));
  OAI210     g0770(.A0(new_new_n725_), .A1(new_new_n466_), .B0(new_new_n111_), .Y(new_new_n793_));
  AOI210     g0771(.A0(new_new_n793_), .A1(new_new_n792_), .B0(new_new_n791_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n475_), .B(new_new_n26_), .Y(new_new_n795_));
  NO2        g0773(.A(new_new_n795_), .B(new_new_n436_), .Y(new_new_n796_));
  NA2        g0774(.A(new_new_n796_), .B(i_2_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n797_), .Y(new_new_n798_));
  AOI210     g0776(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n433_), .Y(new_new_n799_));
  AOI210     g0777(.A0(new_new_n799_), .A1(new_new_n798_), .B0(new_new_n794_), .Y(new_new_n800_));
  NO2        g0778(.A(new_new_n194_), .B(new_new_n126_), .Y(new_new_n801_));
  OAI210     g0779(.A0(new_new_n801_), .A1(new_new_n784_), .B0(i_2_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n175_), .Y(new_new_n803_));
  NO3        g0781(.A(new_new_n649_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n804_));
  AOI210     g0782(.A0(new_new_n803_), .A1(new_new_n88_), .B0(new_new_n804_), .Y(new_new_n805_));
  AOI210     g0783(.A0(new_new_n805_), .A1(new_new_n802_), .B0(new_new_n197_), .Y(new_new_n806_));
  OA210      g0784(.A0(new_new_n650_), .A1(new_new_n127_), .B0(i_13_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n204_), .B(new_new_n207_), .Y(new_new_n808_));
  NA2        g0786(.A(new_new_n153_), .B(new_new_n624_), .Y(new_new_n809_));
  AOI210     g0787(.A0(new_new_n809_), .A1(new_new_n808_), .B0(new_new_n389_), .Y(new_new_n810_));
  AOI210     g0788(.A0(new_new_n214_), .A1(new_new_n149_), .B0(new_new_n539_), .Y(new_new_n811_));
  NA2        g0789(.A(new_new_n811_), .B(new_new_n436_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n102_), .B(new_new_n45_), .Y(new_new_n813_));
  INV        g0791(.A(new_new_n308_), .Y(new_new_n814_));
  NA4        g0792(.A(new_new_n814_), .B(new_new_n312_), .C(new_new_n125_), .D(new_new_n43_), .Y(new_new_n815_));
  OAI210     g0793(.A0(new_new_n815_), .A1(new_new_n813_), .B0(new_new_n812_), .Y(new_new_n816_));
  NO4        g0794(.A(new_new_n816_), .B(new_new_n810_), .C(new_new_n807_), .D(new_new_n806_), .Y(new_new_n817_));
  NA2        g0795(.A(new_new_n600_), .B(new_new_n28_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n783_), .B(new_new_n282_), .Y(new_new_n819_));
  NA2        g0797(.A(new_new_n819_), .B(new_new_n818_), .Y(new_new_n820_));
  NO2        g0798(.A(new_new_n62_), .B(i_12_), .Y(new_new_n821_));
  NO2        g0799(.A(new_new_n821_), .B(new_new_n127_), .Y(new_new_n822_));
  NO2        g0800(.A(new_new_n822_), .B(new_new_n624_), .Y(new_new_n823_));
  AOI220     g0801(.A0(new_new_n823_), .A1(new_new_n36_), .B0(new_new_n820_), .B1(new_new_n47_), .Y(new_new_n824_));
  NA4        g0802(.A(new_new_n824_), .B(new_new_n817_), .C(new_new_n800_), .D(new_new_n790_), .Y(men6));
  NO3        g0803(.A(new_new_n261_), .B(new_new_n314_), .C(i_1_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n189_), .B(new_new_n140_), .Y(new_new_n827_));
  OAI210     g0805(.A0(new_new_n827_), .A1(new_new_n826_), .B0(new_new_n771_), .Y(new_new_n828_));
  NA4        g0806(.A(new_new_n407_), .B(new_new_n502_), .C(new_new_n71_), .D(new_new_n101_), .Y(new_new_n829_));
  INV        g0807(.A(new_new_n829_), .Y(new_new_n830_));
  NO2        g0808(.A(new_new_n227_), .B(new_new_n506_), .Y(new_new_n831_));
  NO2        g0809(.A(i_11_), .B(i_9_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n830_), .B(new_new_n337_), .Y(new_new_n833_));
  AO210      g0811(.A0(new_new_n833_), .A1(new_new_n828_), .B0(i_12_), .Y(new_new_n834_));
  NA2        g0812(.A(new_new_n390_), .B(new_new_n345_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n608_), .B(new_new_n63_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n715_), .B(new_new_n71_), .Y(new_new_n837_));
  NA4        g0815(.A(new_new_n655_), .B(new_new_n837_), .C(new_new_n836_), .D(new_new_n835_), .Y(new_new_n838_));
  INV        g0816(.A(new_new_n201_), .Y(new_new_n839_));
  AOI220     g0817(.A0(new_new_n839_), .A1(new_new_n832_), .B0(new_new_n838_), .B1(new_new_n73_), .Y(new_new_n840_));
  INV        g0818(.A(new_new_n336_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n75_), .B(new_new_n132_), .Y(new_new_n842_));
  INV        g0820(.A(new_new_n125_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n843_), .B(new_new_n47_), .Y(new_new_n844_));
  AOI210     g0822(.A0(new_new_n844_), .A1(new_new_n842_), .B0(new_new_n841_), .Y(new_new_n845_));
  NO2        g0823(.A(new_new_n259_), .B(i_9_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n846_), .B(new_new_n821_), .Y(new_new_n847_));
  AOI210     g0825(.A0(new_new_n847_), .A1(new_new_n538_), .B0(new_new_n189_), .Y(new_new_n848_));
  NO2        g0826(.A(new_new_n32_), .B(i_11_), .Y(new_new_n849_));
  NA3        g0827(.A(new_new_n849_), .B(new_new_n493_), .C(new_new_n407_), .Y(new_new_n850_));
  NAi32      g0828(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n851_));
  AOI210     g0829(.A0(new_new_n754_), .A1(new_new_n86_), .B0(new_new_n851_), .Y(new_new_n852_));
  OAI210     g0830(.A0(new_new_n714_), .A1(new_new_n588_), .B0(new_new_n587_), .Y(new_new_n853_));
  NAi31      g0831(.An(new_new_n852_), .B(new_new_n853_), .C(new_new_n850_), .Y(new_new_n854_));
  OR3        g0832(.A(new_new_n854_), .B(new_new_n848_), .C(new_new_n845_), .Y(new_new_n855_));
  AO220      g0833(.A0(new_new_n373_), .A1(new_new_n363_), .B0(new_new_n415_), .B1(new_new_n624_), .Y(new_new_n856_));
  NA3        g0834(.A(new_new_n856_), .B(new_new_n262_), .C(i_7_), .Y(new_new_n857_));
  OR2        g0835(.A(new_new_n650_), .B(new_new_n466_), .Y(new_new_n858_));
  NA3        g0836(.A(new_new_n858_), .B(new_new_n148_), .C(new_new_n69_), .Y(new_new_n859_));
  AO210      g0837(.A0(new_new_n513_), .A1(new_new_n787_), .B0(new_new_n36_), .Y(new_new_n860_));
  NA3        g0838(.A(new_new_n860_), .B(new_new_n859_), .C(new_new_n857_), .Y(new_new_n861_));
  OAI210     g0839(.A0(new_new_n669_), .A1(i_11_), .B0(new_new_n86_), .Y(new_new_n862_));
  AOI220     g0840(.A0(new_new_n862_), .A1(new_new_n587_), .B0(new_new_n831_), .B1(new_new_n748_), .Y(new_new_n863_));
  NA3        g0841(.A(new_new_n389_), .B(new_new_n245_), .C(new_new_n148_), .Y(new_new_n864_));
  OAI210     g0842(.A0(new_new_n415_), .A1(new_new_n208_), .B0(new_new_n70_), .Y(new_new_n865_));
  NA4        g0843(.A(new_new_n865_), .B(new_new_n864_), .C(new_new_n863_), .D(new_new_n632_), .Y(new_new_n866_));
  AO210      g0844(.A0(new_new_n539_), .A1(new_new_n47_), .B0(new_new_n87_), .Y(new_new_n867_));
  NA3        g0845(.A(new_new_n867_), .B(new_new_n503_), .C(new_new_n225_), .Y(new_new_n868_));
  AOI210     g0846(.A0(new_new_n466_), .A1(new_new_n464_), .B0(new_new_n586_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n112_), .B(new_new_n425_), .Y(new_new_n870_));
  INV        g0848(.A(new_new_n615_), .Y(new_new_n871_));
  NA3        g0849(.A(new_new_n871_), .B(new_new_n336_), .C(i_7_), .Y(new_new_n872_));
  NA4        g0850(.A(new_new_n872_), .B(new_new_n870_), .C(new_new_n869_), .D(new_new_n868_), .Y(new_new_n873_));
  NO4        g0851(.A(new_new_n873_), .B(new_new_n866_), .C(new_new_n861_), .D(new_new_n855_), .Y(new_new_n874_));
  NA4        g0852(.A(new_new_n874_), .B(new_new_n840_), .C(new_new_n834_), .D(new_new_n397_), .Y(men3));
  NA2        g0853(.A(i_12_), .B(i_10_), .Y(new_new_n876_));
  NA2        g0854(.A(i_6_), .B(i_7_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n877_), .B(i_0_), .Y(new_new_n878_));
  NO2        g0856(.A(i_11_), .B(new_new_n243_), .Y(new_new_n879_));
  OAI210     g0857(.A0(new_new_n878_), .A1(new_new_n296_), .B0(new_new_n879_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n880_), .B(new_new_n197_), .Y(new_new_n881_));
  NO3        g0859(.A(new_new_n471_), .B(new_new_n89_), .C(new_new_n45_), .Y(new_new_n882_));
  OA210      g0860(.A0(new_new_n882_), .A1(new_new_n881_), .B0(new_new_n177_), .Y(new_new_n883_));
  NA3        g0861(.A(new_new_n864_), .B(new_new_n632_), .C(new_new_n388_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n884_), .B(new_new_n40_), .Y(new_new_n885_));
  NO3        g0863(.A(new_new_n660_), .B(new_new_n475_), .C(new_new_n132_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n427_), .B(new_new_n46_), .Y(new_new_n887_));
  AOI210     g0865(.A0(new_new_n1106_), .A1(new_new_n885_), .B0(new_new_n49_), .Y(new_new_n888_));
  NO4        g0866(.A(new_new_n393_), .B(new_new_n400_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n889_));
  NA2        g0867(.A(new_new_n189_), .B(new_new_n596_), .Y(new_new_n890_));
  NOi21      g0868(.An(new_new_n890_), .B(new_new_n889_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n740_), .B(new_new_n704_), .Y(new_new_n892_));
  NA2        g0870(.A(new_new_n343_), .B(new_new_n454_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n891_), .B1(new_new_n63_), .Y(new_new_n894_));
  NOi21      g0872(.An(i_5_), .B(i_9_), .Y(new_new_n895_));
  NA2        g0873(.A(new_new_n895_), .B(new_new_n462_), .Y(new_new_n896_));
  AOI210     g0874(.A0(new_new_n272_), .A1(new_new_n495_), .B0(new_new_n719_), .Y(new_new_n897_));
  NO3        g0875(.A(new_new_n430_), .B(new_new_n272_), .C(new_new_n73_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n178_), .B(new_new_n149_), .Y(new_new_n899_));
  AOI210     g0877(.A0(new_new_n899_), .A1(new_new_n251_), .B0(new_new_n898_), .Y(new_new_n900_));
  OAI220     g0878(.A0(new_new_n900_), .A1(new_new_n184_), .B0(new_new_n897_), .B1(new_new_n896_), .Y(new_new_n901_));
  NO4        g0879(.A(new_new_n901_), .B(new_new_n894_), .C(new_new_n888_), .D(new_new_n883_), .Y(new_new_n902_));
  NA2        g0880(.A(new_new_n189_), .B(new_new_n24_), .Y(new_new_n903_));
  NO2        g0881(.A(new_new_n702_), .B(new_new_n621_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n904_), .B(new_new_n903_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n319_), .B(new_new_n130_), .Y(new_new_n906_));
  NAi21      g0884(.An(new_new_n164_), .B(new_new_n454_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n906_), .B(new_new_n417_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n908_), .B(new_new_n905_), .Y(new_new_n909_));
  NO2        g0887(.A(new_new_n407_), .B(new_new_n300_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n910_), .B(new_new_n743_), .Y(new_new_n911_));
  NA2        g0889(.A(new_new_n597_), .B(i_0_), .Y(new_new_n912_));
  NO3        g0890(.A(new_new_n912_), .B(new_new_n402_), .C(new_new_n88_), .Y(new_new_n913_));
  NO4        g0891(.A(new_new_n614_), .B(new_new_n222_), .C(new_new_n433_), .D(i_6_), .Y(new_new_n914_));
  AOI210     g0892(.A0(new_new_n914_), .A1(i_11_), .B0(new_new_n913_), .Y(new_new_n915_));
  AN2        g0893(.A(new_new_n96_), .B(new_new_n250_), .Y(new_new_n916_));
  NA2        g0894(.A(new_new_n783_), .B(new_new_n337_), .Y(new_new_n917_));
  INV        g0895(.A(new_new_n58_), .Y(new_new_n918_));
  OAI220     g0896(.A0(new_new_n918_), .A1(new_new_n917_), .B0(new_new_n688_), .B1(new_new_n560_), .Y(new_new_n919_));
  NA2        g0897(.A(i_0_), .B(i_10_), .Y(new_new_n920_));
  OAI210     g0898(.A0(new_new_n920_), .A1(new_new_n85_), .B0(new_new_n563_), .Y(new_new_n921_));
  NO4        g0899(.A(new_new_n115_), .B(new_new_n58_), .C(new_new_n697_), .D(i_5_), .Y(new_new_n922_));
  AN2        g0900(.A(new_new_n922_), .B(new_new_n921_), .Y(new_new_n923_));
  AOI220     g0901(.A0(new_new_n343_), .A1(new_new_n98_), .B0(new_new_n189_), .B1(new_new_n84_), .Y(new_new_n924_));
  NA2        g0902(.A(new_new_n591_), .B(i_4_), .Y(new_new_n925_));
  NA2        g0903(.A(new_new_n192_), .B(new_new_n207_), .Y(new_new_n926_));
  OAI220     g0904(.A0(new_new_n926_), .A1(new_new_n917_), .B0(new_new_n925_), .B1(new_new_n924_), .Y(new_new_n927_));
  NO4        g0905(.A(new_new_n927_), .B(new_new_n923_), .C(new_new_n919_), .D(new_new_n916_), .Y(new_new_n928_));
  NA4        g0906(.A(new_new_n928_), .B(new_new_n915_), .C(new_new_n911_), .D(new_new_n909_), .Y(new_new_n929_));
  NO2        g0907(.A(new_new_n103_), .B(new_new_n37_), .Y(new_new_n930_));
  NA2        g0908(.A(i_11_), .B(i_9_), .Y(new_new_n931_));
  NO3        g0909(.A(i_12_), .B(new_new_n931_), .C(new_new_n631_), .Y(new_new_n932_));
  AO220      g0910(.A0(new_new_n932_), .A1(new_new_n930_), .B0(new_new_n274_), .B1(new_new_n87_), .Y(new_new_n933_));
  NO2        g0911(.A(new_new_n49_), .B(i_7_), .Y(new_new_n934_));
  NA2        g0912(.A(new_new_n412_), .B(new_new_n182_), .Y(new_new_n935_));
  NA2        g0913(.A(new_new_n935_), .B(new_new_n162_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n931_), .B(new_new_n73_), .Y(new_new_n937_));
  NO2        g0915(.A(new_new_n178_), .B(i_0_), .Y(new_new_n938_));
  INV        g0916(.A(new_new_n938_), .Y(new_new_n939_));
  NA2        g0917(.A(new_new_n493_), .B(new_new_n237_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n387_), .B(new_new_n42_), .Y(new_new_n941_));
  OAI220     g0919(.A0(new_new_n941_), .A1(new_new_n896_), .B0(new_new_n940_), .B1(new_new_n939_), .Y(new_new_n942_));
  NO3        g0920(.A(new_new_n942_), .B(new_new_n936_), .C(new_new_n933_), .Y(new_new_n943_));
  NA2        g0921(.A(new_new_n687_), .B(new_new_n122_), .Y(new_new_n944_));
  NO2        g0922(.A(i_6_), .B(new_new_n944_), .Y(new_new_n945_));
  AOI210     g0923(.A0(new_new_n465_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n946_));
  NA2        g0924(.A(new_new_n174_), .B(new_new_n103_), .Y(new_new_n947_));
  NOi32      g0925(.An(new_new_n946_), .Bn(new_new_n192_), .C(new_new_n947_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n633_), .B(new_new_n337_), .Y(new_new_n949_));
  NO2        g0927(.A(new_new_n949_), .B(new_new_n887_), .Y(new_new_n950_));
  NO3        g0928(.A(new_new_n950_), .B(new_new_n948_), .C(new_new_n945_), .Y(new_new_n951_));
  NOi21      g0929(.An(i_7_), .B(i_5_), .Y(new_new_n952_));
  NOi31      g0930(.An(new_new_n952_), .B(i_0_), .C(new_new_n760_), .Y(new_new_n953_));
  NA3        g0931(.A(new_new_n953_), .B(new_new_n401_), .C(i_6_), .Y(new_new_n954_));
  OA210      g0932(.A0(new_new_n947_), .A1(new_new_n538_), .B0(new_new_n954_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n420_), .B(new_new_n376_), .C(new_new_n372_), .Y(new_new_n956_));
  NO2        g0934(.A(new_new_n266_), .B(new_new_n326_), .Y(new_new_n957_));
  NO2        g0935(.A(new_new_n760_), .B(new_new_n264_), .Y(new_new_n958_));
  AOI210     g0936(.A0(new_new_n958_), .A1(new_new_n957_), .B0(new_new_n956_), .Y(new_new_n959_));
  NA4        g0937(.A(new_new_n959_), .B(new_new_n955_), .C(new_new_n951_), .D(new_new_n943_), .Y(new_new_n960_));
  NO2        g0938(.A(new_new_n903_), .B(new_new_n246_), .Y(new_new_n961_));
  AN2        g0939(.A(new_new_n342_), .B(new_new_n337_), .Y(new_new_n962_));
  AN2        g0940(.A(new_new_n962_), .B(new_new_n899_), .Y(new_new_n963_));
  OAI210     g0941(.A0(new_new_n963_), .A1(new_new_n961_), .B0(i_10_), .Y(new_new_n964_));
  NO2        g0942(.A(new_new_n876_), .B(new_new_n325_), .Y(new_new_n965_));
  OA210      g0943(.A0(new_new_n493_), .A1(new_new_n229_), .B0(new_new_n492_), .Y(new_new_n966_));
  NA2        g0944(.A(new_new_n965_), .B(new_new_n937_), .Y(new_new_n967_));
  NA3        g0945(.A(new_new_n492_), .B(new_new_n427_), .C(new_new_n46_), .Y(new_new_n968_));
  OAI210     g0946(.A0(new_new_n907_), .A1(i_6_), .B0(new_new_n968_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n937_), .B(new_new_n312_), .Y(new_new_n970_));
  NA2        g0948(.A(new_new_n191_), .B(new_new_n970_), .Y(new_new_n971_));
  AOI220     g0949(.A0(new_new_n971_), .A1(new_new_n493_), .B0(new_new_n969_), .B1(new_new_n73_), .Y(new_new_n972_));
  NA3        g0950(.A(i_5_), .B(new_new_n399_), .C(new_new_n669_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n92_), .B(new_new_n45_), .Y(new_new_n974_));
  NO2        g0952(.A(new_new_n75_), .B(new_new_n785_), .Y(new_new_n975_));
  AOI220     g0953(.A0(new_new_n975_), .A1(new_new_n974_), .B0(new_new_n177_), .B1(new_new_n621_), .Y(new_new_n976_));
  AOI210     g0954(.A0(new_new_n976_), .A1(new_new_n973_), .B0(new_new_n48_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n614_), .B(new_new_n371_), .C(new_new_n24_), .Y(new_new_n978_));
  INV        g0956(.A(new_new_n978_), .Y(new_new_n979_));
  NAi21      g0957(.An(i_9_), .B(i_5_), .Y(new_new_n980_));
  NO2        g0958(.A(new_new_n627_), .B(new_new_n105_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n981_), .B(i_0_), .Y(new_new_n982_));
  OAI220     g0960(.A0(new_new_n982_), .A1(new_new_n85_), .B0(new_new_n979_), .B1(new_new_n175_), .Y(new_new_n983_));
  NO3        g0961(.A(new_new_n983_), .B(new_new_n977_), .C(new_new_n542_), .Y(new_new_n984_));
  NA4        g0962(.A(new_new_n984_), .B(new_new_n972_), .C(new_new_n967_), .D(new_new_n964_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n985_), .B(new_new_n960_), .C(new_new_n929_), .Y(new_new_n986_));
  NO2        g0964(.A(i_0_), .B(new_new_n760_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n920_), .B(new_new_n988_), .Y(new_new_n989_));
  NO3        g0967(.A(new_new_n105_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n990_));
  AO220      g0968(.A0(new_new_n990_), .A1(new_new_n989_), .B0(new_new_n987_), .B1(new_new_n177_), .Y(new_new_n991_));
  AOI210     g0969(.A0(new_new_n836_), .A1(new_new_n717_), .B0(new_new_n947_), .Y(new_new_n992_));
  AOI210     g0970(.A0(new_new_n991_), .A1(new_new_n360_), .B0(new_new_n992_), .Y(new_new_n993_));
  NA2        g0971(.A(new_new_n771_), .B(new_new_n147_), .Y(new_new_n994_));
  INV        g0972(.A(new_new_n994_), .Y(new_new_n995_));
  NA3        g0973(.A(new_new_n995_), .B(new_new_n704_), .C(new_new_n73_), .Y(new_new_n996_));
  NO2        g0974(.A(new_new_n853_), .B(new_new_n420_), .Y(new_new_n997_));
  NA3        g0975(.A(new_new_n878_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n998_));
  NA2        g0976(.A(new_new_n879_), .B(i_9_), .Y(new_new_n999_));
  AOI210     g0977(.A0(new_new_n998_), .A1(new_new_n519_), .B0(new_new_n999_), .Y(new_new_n1000_));
  OAI210     g0978(.A0(new_new_n251_), .A1(i_9_), .B0(new_new_n236_), .Y(new_new_n1001_));
  AOI210     g0979(.A0(new_new_n1001_), .A1(new_new_n912_), .B0(new_new_n155_), .Y(new_new_n1002_));
  NO3        g0980(.A(new_new_n1002_), .B(new_new_n1000_), .C(new_new_n997_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n1003_), .B(new_new_n996_), .C(new_new_n993_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n962_), .B(new_new_n389_), .Y(new_new_n1005_));
  AOI210     g0983(.A0(new_new_n307_), .A1(new_new_n164_), .B0(new_new_n1005_), .Y(new_new_n1006_));
  NA3        g0984(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n1007_));
  NA2        g0985(.A(new_new_n934_), .B(new_new_n507_), .Y(new_new_n1008_));
  AOI210     g0986(.A0(new_new_n1007_), .A1(new_new_n164_), .B0(new_new_n1008_), .Y(new_new_n1009_));
  NO2        g0987(.A(new_new_n1009_), .B(new_new_n1006_), .Y(new_new_n1010_));
  NO3        g0988(.A(new_new_n920_), .B(new_new_n895_), .C(new_new_n194_), .Y(new_new_n1011_));
  AOI220     g0989(.A0(new_new_n1011_), .A1(i_11_), .B0(new_new_n592_), .B1(new_new_n75_), .Y(new_new_n1012_));
  NO3        g0990(.A(new_new_n216_), .B(new_new_n400_), .C(i_0_), .Y(new_new_n1013_));
  OAI210     g0991(.A0(new_new_n1013_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n1014_));
  INV        g0992(.A(new_new_n225_), .Y(new_new_n1015_));
  OAI220     g0993(.A0(new_new_n554_), .A1(new_new_n140_), .B0(new_new_n674_), .B1(new_new_n644_), .Y(new_new_n1016_));
  NA3        g0994(.A(new_new_n1016_), .B(i_7_), .C(new_new_n1015_), .Y(new_new_n1017_));
  NA4        g0995(.A(new_new_n1017_), .B(new_new_n1014_), .C(new_new_n1012_), .D(new_new_n1010_), .Y(new_new_n1018_));
  NO2        g0996(.A(new_new_n249_), .B(new_new_n92_), .Y(new_new_n1019_));
  AOI210     g0997(.A0(new_new_n1019_), .A1(new_new_n987_), .B0(new_new_n109_), .Y(new_new_n1020_));
  AOI220     g0998(.A0(new_new_n952_), .A1(new_new_n507_), .B0(new_new_n878_), .B1(new_new_n165_), .Y(new_new_n1021_));
  NA2        g0999(.A(new_new_n363_), .B(new_new_n179_), .Y(new_new_n1022_));
  OA220      g1000(.A0(new_new_n1022_), .A1(new_new_n1021_), .B0(new_new_n1020_), .B1(i_5_), .Y(new_new_n1023_));
  AOI210     g1001(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n178_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n1024_), .B(new_new_n966_), .Y(new_new_n1025_));
  INV        g1003(.A(new_new_n570_), .Y(new_new_n1026_));
  NO3        g1004(.A(new_new_n887_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1027_));
  INV        g1005(.A(new_new_n512_), .Y(new_new_n1028_));
  NO3        g1006(.A(new_new_n1028_), .B(new_new_n1027_), .C(new_new_n1026_), .Y(new_new_n1029_));
  NA3        g1007(.A(new_new_n407_), .B(new_new_n174_), .C(new_new_n173_), .Y(new_new_n1030_));
  NA3        g1008(.A(new_new_n934_), .B(new_new_n296_), .C(new_new_n236_), .Y(new_new_n1031_));
  NA2        g1009(.A(new_new_n1031_), .B(new_new_n1030_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n407_), .B(new_new_n344_), .C(new_new_n228_), .Y(new_new_n1033_));
  INV        g1011(.A(new_new_n1033_), .Y(new_new_n1034_));
  NOi31      g1012(.An(new_new_n406_), .B(new_new_n988_), .C(new_new_n246_), .Y(new_new_n1035_));
  NO3        g1013(.A(new_new_n931_), .B(new_new_n225_), .C(new_new_n194_), .Y(new_new_n1036_));
  NO4        g1014(.A(new_new_n1036_), .B(new_new_n1035_), .C(new_new_n1034_), .D(new_new_n1032_), .Y(new_new_n1037_));
  NA4        g1015(.A(new_new_n1037_), .B(new_new_n1029_), .C(new_new_n1025_), .D(new_new_n1023_), .Y(new_new_n1038_));
  NO2        g1016(.A(new_new_n85_), .B(i_5_), .Y(new_new_n1039_));
  NA3        g1017(.A(new_new_n879_), .B(new_new_n110_), .C(new_new_n125_), .Y(new_new_n1040_));
  INV        g1018(.A(new_new_n1040_), .Y(new_new_n1041_));
  NA2        g1019(.A(new_new_n1041_), .B(new_new_n1039_), .Y(new_new_n1042_));
  NA3        g1020(.A(new_new_n312_), .B(i_5_), .C(new_new_n197_), .Y(new_new_n1043_));
  NAi31      g1021(.An(new_new_n248_), .B(new_new_n1043_), .C(new_new_n249_), .Y(new_new_n1044_));
  NO4        g1022(.A(new_new_n246_), .B(new_new_n216_), .C(i_0_), .D(i_12_), .Y(new_new_n1045_));
  AOI220     g1023(.A0(new_new_n1045_), .A1(new_new_n1044_), .B0(new_new_n830_), .B1(new_new_n179_), .Y(new_new_n1046_));
  AN2        g1024(.A(new_new_n920_), .B(new_new_n155_), .Y(new_new_n1047_));
  NO4        g1025(.A(new_new_n1047_), .B(i_12_), .C(new_new_n676_), .D(new_new_n132_), .Y(new_new_n1048_));
  NA2        g1026(.A(new_new_n1048_), .B(new_new_n225_), .Y(new_new_n1049_));
  NA3        g1027(.A(new_new_n98_), .B(new_new_n596_), .C(i_11_), .Y(new_new_n1050_));
  NO2        g1028(.A(new_new_n1050_), .B(new_new_n157_), .Y(new_new_n1051_));
  NA2        g1029(.A(new_new_n64_), .B(new_new_n101_), .Y(new_new_n1052_));
  NO2        g1030(.A(new_new_n1052_), .B(new_new_n1043_), .Y(new_new_n1053_));
  AOI210     g1031(.A0(new_new_n1053_), .A1(new_new_n938_), .B0(new_new_n1051_), .Y(new_new_n1054_));
  NA4        g1032(.A(new_new_n1054_), .B(new_new_n1049_), .C(new_new_n1046_), .D(new_new_n1042_), .Y(new_new_n1055_));
  NO4        g1033(.A(new_new_n1055_), .B(new_new_n1038_), .C(new_new_n1018_), .D(new_new_n1004_), .Y(new_new_n1056_));
  NA2        g1034(.A(new_new_n849_), .B(new_new_n37_), .Y(new_new_n1057_));
  NA3        g1035(.A(new_new_n946_), .B(new_new_n384_), .C(i_5_), .Y(new_new_n1058_));
  NA3        g1036(.A(new_new_n1058_), .B(new_new_n1057_), .C(new_new_n639_), .Y(new_new_n1059_));
  NA2        g1037(.A(new_new_n1059_), .B(new_new_n212_), .Y(new_new_n1060_));
  AN2        g1038(.A(new_new_n730_), .B(new_new_n385_), .Y(new_new_n1061_));
  NA2        g1039(.A(new_new_n190_), .B(new_new_n192_), .Y(new_new_n1062_));
  AO210      g1040(.A0(new_new_n1061_), .A1(new_new_n33_), .B0(new_new_n1062_), .Y(new_new_n1063_));
  OAI210     g1041(.A0(new_new_n643_), .A1(new_new_n641_), .B0(new_new_n325_), .Y(new_new_n1064_));
  NA2        g1042(.A(new_new_n1064_), .B(new_new_n1063_), .Y(new_new_n1065_));
  NO2        g1043(.A(new_new_n480_), .B(new_new_n272_), .Y(new_new_n1066_));
  NO4        g1044(.A(new_new_n239_), .B(new_new_n146_), .C(new_new_n708_), .D(new_new_n37_), .Y(new_new_n1067_));
  NO3        g1045(.A(new_new_n1067_), .B(new_new_n1066_), .C(new_new_n914_), .Y(new_new_n1068_));
  OAI210     g1046(.A0(new_new_n1050_), .A1(new_new_n149_), .B0(new_new_n1068_), .Y(new_new_n1069_));
  AOI210     g1047(.A0(new_new_n1065_), .A1(new_new_n49_), .B0(new_new_n1069_), .Y(new_new_n1070_));
  AOI210     g1048(.A0(new_new_n1070_), .A1(new_new_n1060_), .B0(new_new_n73_), .Y(new_new_n1071_));
  NO2        g1049(.A(new_new_n589_), .B(new_new_n396_), .Y(new_new_n1072_));
  NO2        g1050(.A(new_new_n1072_), .B(new_new_n791_), .Y(new_new_n1073_));
  OAI210     g1051(.A0(new_new_n80_), .A1(new_new_n55_), .B0(new_new_n108_), .Y(new_new_n1074_));
  NA2        g1052(.A(new_new_n1074_), .B(new_new_n76_), .Y(new_new_n1075_));
  AOI210     g1053(.A0(new_new_n1024_), .A1(new_new_n934_), .B0(new_new_n953_), .Y(new_new_n1076_));
  AOI210     g1054(.A0(new_new_n1076_), .A1(new_new_n1075_), .B0(new_new_n708_), .Y(new_new_n1077_));
  NA2        g1055(.A(new_new_n266_), .B(new_new_n57_), .Y(new_new_n1078_));
  AOI220     g1056(.A0(new_new_n1078_), .A1(new_new_n76_), .B0(new_new_n358_), .B1(new_new_n261_), .Y(new_new_n1079_));
  NO2        g1057(.A(new_new_n1079_), .B(new_new_n243_), .Y(new_new_n1080_));
  NA3        g1058(.A(new_new_n96_), .B(new_new_n314_), .C(new_new_n31_), .Y(new_new_n1081_));
  INV        g1059(.A(new_new_n1081_), .Y(new_new_n1082_));
  NO3        g1060(.A(new_new_n1082_), .B(new_new_n1080_), .C(new_new_n1077_), .Y(new_new_n1083_));
  OAI210     g1061(.A0(new_new_n274_), .A1(new_new_n160_), .B0(new_new_n88_), .Y(new_new_n1084_));
  NA3        g1062(.A(new_new_n795_), .B(new_new_n296_), .C(new_new_n80_), .Y(new_new_n1085_));
  AOI210     g1063(.A0(new_new_n1085_), .A1(new_new_n1084_), .B0(i_11_), .Y(new_new_n1086_));
  OAI210     g1064(.A0(new_new_n1107_), .A1(new_new_n946_), .B0(new_new_n212_), .Y(new_new_n1087_));
  NA2        g1065(.A(new_new_n166_), .B(i_5_), .Y(new_new_n1088_));
  AOI210     g1066(.A0(new_new_n1087_), .A1(new_new_n808_), .B0(new_new_n1088_), .Y(new_new_n1089_));
  NO3        g1067(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1090_));
  OAI210     g1068(.A0(new_new_n957_), .A1(new_new_n314_), .B0(new_new_n1090_), .Y(new_new_n1091_));
  NO2        g1069(.A(new_new_n1091_), .B(new_new_n760_), .Y(new_new_n1092_));
  NO4        g1070(.A(new_new_n980_), .B(new_new_n496_), .C(new_new_n260_), .D(new_new_n259_), .Y(new_new_n1093_));
  NO2        g1071(.A(new_new_n1093_), .B(new_new_n586_), .Y(new_new_n1094_));
  INV        g1072(.A(new_new_n377_), .Y(new_new_n1095_));
  AOI210     g1073(.A0(new_new_n1095_), .A1(new_new_n1094_), .B0(new_new_n41_), .Y(new_new_n1096_));
  NO4        g1074(.A(new_new_n1096_), .B(new_new_n1092_), .C(new_new_n1089_), .D(new_new_n1086_), .Y(new_new_n1097_));
  OAI210     g1075(.A0(new_new_n1083_), .A1(i_4_), .B0(new_new_n1097_), .Y(new_new_n1098_));
  NO3        g1076(.A(new_new_n1098_), .B(new_new_n1073_), .C(new_new_n1071_), .Y(new_new_n1099_));
  NA4        g1077(.A(new_new_n1099_), .B(new_new_n1056_), .C(new_new_n986_), .D(new_new_n902_), .Y(men4));
  INV        g1078(.A(new_new_n734_), .Y(new_new_n1103_));
  INV        g1079(.A(i_2_), .Y(new_new_n1104_));
  INV        g1080(.A(new_new_n503_), .Y(new_new_n1105_));
  INV        g1081(.A(new_new_n886_), .Y(new_new_n1106_));
  INV        g1082(.A(i_12_), .Y(new_new_n1107_));
  INV        g1083(.A(new_new_n82_), .Y(new_new_n1108_));
endmodule


