library verilog;
use verilog.vl_types.all;
entity mux4bits4x1_vlg_vec_tst is
end mux4bits4x1_vlg_vec_tst;
