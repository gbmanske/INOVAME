//Benchmark atmr_misex3_1774_0.0625

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1042_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1061_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1072_, ori_ori_n1073_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1122_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1172_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  INV        o0001(.A(d), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  INV        o0010(.A(h), .Y(ori_ori_n39_));
  NAi21      o0011(.An(j), .B(l), .Y(ori_ori_n40_));
  NAi32      o0012(.An(n), .Bn(g), .C(m), .Y(ori_ori_n41_));
  NO3        o0013(.A(ori_ori_n41_), .B(ori_ori_n40_), .C(ori_ori_n39_), .Y(ori_ori_n42_));
  NAi31      o0014(.An(n), .B(m), .C(l), .Y(ori_ori_n43_));
  INV        o0015(.A(i), .Y(ori_ori_n44_));
  AN2        o0016(.A(h), .B(g), .Y(ori_ori_n45_));
  NA2        o0017(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori_ori_n46_));
  NO2        o0018(.A(ori_ori_n46_), .B(ori_ori_n43_), .Y(ori_ori_n47_));
  NAi21      o0019(.An(n), .B(m), .Y(ori_ori_n48_));
  NOi32      o0020(.An(k), .Bn(h), .C(l), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(g), .Y(ori_ori_n50_));
  INV        o0022(.A(ori_ori_n50_), .Y(ori_ori_n51_));
  NO2        o0023(.A(ori_ori_n51_), .B(ori_ori_n48_), .Y(ori_ori_n52_));
  NO3        o0024(.A(ori_ori_n52_), .B(ori_ori_n47_), .C(ori_ori_n42_), .Y(ori_ori_n53_));
  AOI210     o0025(.A0(ori_ori_n53_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n54_));
  INV        o0026(.A(c), .Y(ori_ori_n55_));
  NA2        o0027(.A(e), .B(b), .Y(ori_ori_n56_));
  NO2        o0028(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  INV        o0029(.A(d), .Y(ori_ori_n58_));
  NAi21      o0030(.An(i), .B(h), .Y(ori_ori_n59_));
  NAi41      o0031(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n60_));
  NA2        o0032(.A(g), .B(f), .Y(ori_ori_n61_));
  NO2        o0033(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n62_));
  NAi32      o0034(.An(n), .Bn(k), .C(m), .Y(ori_ori_n63_));
  NAi31      o0035(.An(l), .B(m), .C(k), .Y(ori_ori_n64_));
  NAi21      o0036(.An(e), .B(h), .Y(ori_ori_n65_));
  NAi41      o0037(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n66_));
  INV        o0038(.A(m), .Y(ori_ori_n67_));
  NOi21      o0039(.An(k), .B(l), .Y(ori_ori_n68_));
  NA2        o0040(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n69_));
  AN4        o0041(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n70_));
  NOi21      o0042(.An(h), .B(f), .Y(ori_ori_n71_));
  NA2        o0043(.A(ori_ori_n71_), .B(ori_ori_n70_), .Y(ori_ori_n72_));
  NAi32      o0044(.An(m), .Bn(k), .C(j), .Y(ori_ori_n73_));
  NOi32      o0045(.An(h), .Bn(g), .C(f), .Y(ori_ori_n74_));
  INV        o0046(.A(n), .Y(ori_ori_n75_));
  NOi32      o0047(.An(e), .Bn(b), .C(d), .Y(ori_ori_n76_));
  NA2        o0048(.A(ori_ori_n76_), .B(ori_ori_n75_), .Y(ori_ori_n77_));
  INV        o0049(.A(j), .Y(ori_ori_n78_));
  AN3        o0050(.A(m), .B(k), .C(i), .Y(ori_ori_n79_));
  NA3        o0051(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .Y(ori_ori_n80_));
  NO2        o0052(.A(ori_ori_n80_), .B(f), .Y(ori_ori_n81_));
  NAi32      o0053(.An(g), .Bn(f), .C(h), .Y(ori_ori_n82_));
  NAi31      o0054(.An(j), .B(m), .C(l), .Y(ori_ori_n83_));
  NO2        o0055(.A(ori_ori_n83_), .B(ori_ori_n82_), .Y(ori_ori_n84_));
  NA2        o0056(.A(m), .B(l), .Y(ori_ori_n85_));
  NAi31      o0057(.An(k), .B(j), .C(g), .Y(ori_ori_n86_));
  NO3        o0058(.A(ori_ori_n86_), .B(ori_ori_n85_), .C(f), .Y(ori_ori_n87_));
  AN2        o0059(.A(j), .B(g), .Y(ori_ori_n88_));
  NOi32      o0060(.An(m), .Bn(l), .C(i), .Y(ori_ori_n89_));
  NOi32      o0061(.An(m), .Bn(j), .C(k), .Y(ori_ori_n90_));
  AOI220     o0062(.A0(ori_ori_n90_), .A1(g), .B0(ori_ori_n89_), .B1(ori_ori_n88_), .Y(ori_ori_n91_));
  NO2        o0063(.A(ori_ori_n91_), .B(f), .Y(ori_ori_n92_));
  NO3        o0064(.A(ori_ori_n92_), .B(ori_ori_n84_), .C(ori_ori_n81_), .Y(ori_ori_n93_));
  NAi41      o0065(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n94_));
  AN2        o0066(.A(e), .B(b), .Y(ori_ori_n95_));
  NOi31      o0067(.An(c), .B(h), .C(f), .Y(ori_ori_n96_));
  NA2        o0068(.A(ori_ori_n96_), .B(ori_ori_n95_), .Y(ori_ori_n97_));
  NO2        o0069(.A(ori_ori_n97_), .B(ori_ori_n94_), .Y(ori_ori_n98_));
  NOi21      o0070(.An(i), .B(h), .Y(ori_ori_n99_));
  INV        o0071(.A(a), .Y(ori_ori_n100_));
  NA2        o0072(.A(ori_ori_n95_), .B(ori_ori_n100_), .Y(ori_ori_n101_));
  INV        o0073(.A(l), .Y(ori_ori_n102_));
  NOi21      o0074(.An(m), .B(n), .Y(ori_ori_n103_));
  AN2        o0075(.A(k), .B(h), .Y(ori_ori_n104_));
  INV        o0076(.A(b), .Y(ori_ori_n105_));
  NA2        o0077(.A(l), .B(j), .Y(ori_ori_n106_));
  AN2        o0078(.A(k), .B(i), .Y(ori_ori_n107_));
  NA2        o0079(.A(ori_ori_n107_), .B(ori_ori_n106_), .Y(ori_ori_n108_));
  NA2        o0080(.A(g), .B(e), .Y(ori_ori_n109_));
  NOi32      o0081(.An(c), .Bn(a), .C(d), .Y(ori_ori_n110_));
  NA2        o0082(.A(ori_ori_n110_), .B(ori_ori_n103_), .Y(ori_ori_n111_));
  INV        o0083(.A(ori_ori_n98_), .Y(ori_ori_n112_));
  OAI210     o0084(.A0(ori_ori_n93_), .A1(ori_ori_n77_), .B0(ori_ori_n112_), .Y(ori_ori_n113_));
  NOi31      o0085(.An(k), .B(m), .C(j), .Y(ori_ori_n114_));
  NA3        o0086(.A(ori_ori_n114_), .B(ori_ori_n71_), .C(ori_ori_n70_), .Y(ori_ori_n115_));
  NOi31      o0087(.An(k), .B(m), .C(i), .Y(ori_ori_n116_));
  NA3        o0088(.A(ori_ori_n116_), .B(ori_ori_n74_), .C(ori_ori_n70_), .Y(ori_ori_n117_));
  NA2        o0089(.A(ori_ori_n117_), .B(ori_ori_n115_), .Y(ori_ori_n118_));
  NOi32      o0090(.An(f), .Bn(b), .C(e), .Y(ori_ori_n119_));
  NAi21      o0091(.An(g), .B(h), .Y(ori_ori_n120_));
  NAi21      o0092(.An(m), .B(n), .Y(ori_ori_n121_));
  NAi41      o0093(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n122_));
  NAi31      o0094(.An(j), .B(k), .C(h), .Y(ori_ori_n123_));
  NO3        o0095(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(ori_ori_n121_), .Y(ori_ori_n124_));
  INV        o0096(.A(ori_ori_n124_), .Y(ori_ori_n125_));
  NO2        o0097(.A(k), .B(j), .Y(ori_ori_n126_));
  NO2        o0098(.A(ori_ori_n126_), .B(ori_ori_n121_), .Y(ori_ori_n127_));
  AN2        o0099(.A(k), .B(j), .Y(ori_ori_n128_));
  NAi21      o0100(.An(c), .B(b), .Y(ori_ori_n129_));
  NA2        o0101(.A(f), .B(d), .Y(ori_ori_n130_));
  NO4        o0102(.A(ori_ori_n130_), .B(ori_ori_n129_), .C(ori_ori_n128_), .D(ori_ori_n120_), .Y(ori_ori_n131_));
  NA2        o0103(.A(h), .B(c), .Y(ori_ori_n132_));
  NAi31      o0104(.An(f), .B(e), .C(b), .Y(ori_ori_n133_));
  NA2        o0105(.A(ori_ori_n131_), .B(ori_ori_n127_), .Y(ori_ori_n134_));
  NA2        o0106(.A(d), .B(b), .Y(ori_ori_n135_));
  NAi21      o0107(.An(e), .B(f), .Y(ori_ori_n136_));
  NO2        o0108(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n137_));
  NA2        o0109(.A(b), .B(a), .Y(ori_ori_n138_));
  NAi21      o0110(.An(e), .B(g), .Y(ori_ori_n139_));
  NAi21      o0111(.An(c), .B(d), .Y(ori_ori_n140_));
  NAi31      o0112(.An(l), .B(k), .C(h), .Y(ori_ori_n141_));
  NO2        o0113(.A(ori_ori_n121_), .B(ori_ori_n141_), .Y(ori_ori_n142_));
  NA2        o0114(.A(ori_ori_n142_), .B(ori_ori_n137_), .Y(ori_ori_n143_));
  NAi41      o0115(.An(ori_ori_n118_), .B(ori_ori_n143_), .C(ori_ori_n134_), .D(ori_ori_n125_), .Y(ori_ori_n144_));
  NAi31      o0116(.An(e), .B(f), .C(b), .Y(ori_ori_n145_));
  NOi21      o0117(.An(g), .B(d), .Y(ori_ori_n146_));
  NO2        o0118(.A(ori_ori_n146_), .B(ori_ori_n145_), .Y(ori_ori_n147_));
  NOi21      o0119(.An(h), .B(i), .Y(ori_ori_n148_));
  NOi21      o0120(.An(k), .B(m), .Y(ori_ori_n149_));
  NA3        o0121(.A(ori_ori_n149_), .B(ori_ori_n148_), .C(n), .Y(ori_ori_n150_));
  NOi21      o0122(.An(ori_ori_n147_), .B(ori_ori_n150_), .Y(ori_ori_n151_));
  NOi21      o0123(.An(h), .B(g), .Y(ori_ori_n152_));
  NO2        o0124(.A(ori_ori_n130_), .B(ori_ori_n129_), .Y(ori_ori_n153_));
  NAi31      o0125(.An(l), .B(j), .C(h), .Y(ori_ori_n154_));
  INV        o0126(.A(ori_ori_n48_), .Y(ori_ori_n155_));
  NA2        o0127(.A(ori_ori_n155_), .B(ori_ori_n62_), .Y(ori_ori_n156_));
  NOi32      o0128(.An(n), .Bn(k), .C(m), .Y(ori_ori_n157_));
  INV        o0129(.A(ori_ori_n156_), .Y(ori_ori_n158_));
  NAi31      o0130(.An(d), .B(f), .C(c), .Y(ori_ori_n159_));
  NAi31      o0131(.An(e), .B(f), .C(c), .Y(ori_ori_n160_));
  NA2        o0132(.A(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NA2        o0133(.A(j), .B(h), .Y(ori_ori_n162_));
  OR3        o0134(.A(n), .B(m), .C(k), .Y(ori_ori_n163_));
  NO2        o0135(.A(ori_ori_n163_), .B(ori_ori_n162_), .Y(ori_ori_n164_));
  NAi32      o0136(.An(m), .Bn(k), .C(n), .Y(ori_ori_n165_));
  NO2        o0137(.A(ori_ori_n165_), .B(ori_ori_n162_), .Y(ori_ori_n166_));
  AOI220     o0138(.A0(ori_ori_n166_), .A1(ori_ori_n147_), .B0(ori_ori_n164_), .B1(ori_ori_n161_), .Y(ori_ori_n167_));
  NO2        o0139(.A(n), .B(m), .Y(ori_ori_n168_));
  NA2        o0140(.A(ori_ori_n168_), .B(ori_ori_n49_), .Y(ori_ori_n169_));
  NAi21      o0141(.An(f), .B(e), .Y(ori_ori_n170_));
  NA2        o0142(.A(d), .B(c), .Y(ori_ori_n171_));
  NO2        o0143(.A(ori_ori_n171_), .B(ori_ori_n170_), .Y(ori_ori_n172_));
  NOi21      o0144(.An(ori_ori_n172_), .B(ori_ori_n169_), .Y(ori_ori_n173_));
  NAi31      o0145(.An(m), .B(n), .C(b), .Y(ori_ori_n174_));
  NAi21      o0146(.An(h), .B(f), .Y(ori_ori_n175_));
  NO2        o0147(.A(ori_ori_n174_), .B(ori_ori_n140_), .Y(ori_ori_n176_));
  NOi32      o0148(.An(f), .Bn(c), .C(d), .Y(ori_ori_n177_));
  NOi32      o0149(.An(f), .Bn(c), .C(e), .Y(ori_ori_n178_));
  NO2        o0150(.A(ori_ori_n178_), .B(ori_ori_n177_), .Y(ori_ori_n179_));
  NO3        o0151(.A(n), .B(m), .C(j), .Y(ori_ori_n180_));
  NA2        o0152(.A(ori_ori_n180_), .B(ori_ori_n104_), .Y(ori_ori_n181_));
  AO210      o0153(.A0(ori_ori_n181_), .A1(ori_ori_n169_), .B0(ori_ori_n179_), .Y(ori_ori_n182_));
  NAi31      o0154(.An(ori_ori_n173_), .B(ori_ori_n182_), .C(ori_ori_n167_), .Y(ori_ori_n183_));
  OR4        o0155(.A(ori_ori_n183_), .B(ori_ori_n158_), .C(ori_ori_n151_), .D(ori_ori_n144_), .Y(ori_ori_n184_));
  NO3        o0156(.A(ori_ori_n184_), .B(ori_ori_n113_), .C(ori_ori_n54_), .Y(ori_ori_n185_));
  NA3        o0157(.A(m), .B(ori_ori_n102_), .C(j), .Y(ori_ori_n186_));
  NAi31      o0158(.An(n), .B(h), .C(g), .Y(ori_ori_n187_));
  NO2        o0159(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NOi32      o0160(.An(m), .Bn(k), .C(l), .Y(ori_ori_n189_));
  NA3        o0161(.A(ori_ori_n189_), .B(ori_ori_n78_), .C(g), .Y(ori_ori_n190_));
  NO2        o0162(.A(ori_ori_n190_), .B(n), .Y(ori_ori_n191_));
  NOi21      o0163(.An(k), .B(j), .Y(ori_ori_n192_));
  NA4        o0164(.A(ori_ori_n192_), .B(ori_ori_n103_), .C(i), .D(g), .Y(ori_ori_n193_));
  AN2        o0165(.A(i), .B(g), .Y(ori_ori_n194_));
  NA3        o0166(.A(ori_ori_n68_), .B(ori_ori_n194_), .C(ori_ori_n103_), .Y(ori_ori_n195_));
  NA2        o0167(.A(ori_ori_n195_), .B(ori_ori_n193_), .Y(ori_ori_n196_));
  NO3        o0168(.A(ori_ori_n196_), .B(ori_ori_n191_), .C(ori_ori_n188_), .Y(ori_ori_n197_));
  NAi41      o0169(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n198_));
  INV        o0170(.A(ori_ori_n198_), .Y(ori_ori_n199_));
  INV        o0171(.A(f), .Y(ori_ori_n200_));
  INV        o0172(.A(g), .Y(ori_ori_n201_));
  NOi31      o0173(.An(i), .B(j), .C(h), .Y(ori_ori_n202_));
  NOi21      o0174(.An(l), .B(m), .Y(ori_ori_n203_));
  NA2        o0175(.A(ori_ori_n203_), .B(ori_ori_n202_), .Y(ori_ori_n204_));
  NO3        o0176(.A(ori_ori_n204_), .B(ori_ori_n201_), .C(ori_ori_n200_), .Y(ori_ori_n205_));
  NA2        o0177(.A(ori_ori_n205_), .B(ori_ori_n199_), .Y(ori_ori_n206_));
  OAI210     o0178(.A0(ori_ori_n197_), .A1(ori_ori_n32_), .B0(ori_ori_n206_), .Y(ori_ori_n207_));
  NOi21      o0179(.An(n), .B(m), .Y(ori_ori_n208_));
  NOi32      o0180(.An(l), .Bn(i), .C(j), .Y(ori_ori_n209_));
  NA2        o0181(.A(ori_ori_n209_), .B(ori_ori_n208_), .Y(ori_ori_n210_));
  OA220      o0182(.A0(ori_ori_n210_), .A1(ori_ori_n97_), .B0(ori_ori_n73_), .B1(ori_ori_n72_), .Y(ori_ori_n211_));
  NAi21      o0183(.An(j), .B(h), .Y(ori_ori_n212_));
  XN2        o0184(.A(i), .B(h), .Y(ori_ori_n213_));
  NA2        o0185(.A(ori_ori_n213_), .B(ori_ori_n212_), .Y(ori_ori_n214_));
  NOi31      o0186(.An(k), .B(n), .C(m), .Y(ori_ori_n215_));
  NOi31      o0187(.An(ori_ori_n215_), .B(ori_ori_n171_), .C(ori_ori_n170_), .Y(ori_ori_n216_));
  NA2        o0188(.A(ori_ori_n216_), .B(ori_ori_n214_), .Y(ori_ori_n217_));
  NAi31      o0189(.An(f), .B(e), .C(c), .Y(ori_ori_n218_));
  NO4        o0190(.A(ori_ori_n218_), .B(ori_ori_n163_), .C(ori_ori_n162_), .D(ori_ori_n58_), .Y(ori_ori_n219_));
  NA4        o0191(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n220_));
  NAi32      o0192(.An(m), .Bn(i), .C(k), .Y(ori_ori_n221_));
  INV        o0193(.A(k), .Y(ori_ori_n222_));
  INV        o0194(.A(ori_ori_n219_), .Y(ori_ori_n223_));
  NAi21      o0195(.An(n), .B(a), .Y(ori_ori_n224_));
  NO2        o0196(.A(ori_ori_n224_), .B(ori_ori_n135_), .Y(ori_ori_n225_));
  NAi41      o0197(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n226_));
  NO2        o0198(.A(ori_ori_n226_), .B(e), .Y(ori_ori_n227_));
  NA2        o0199(.A(ori_ori_n227_), .B(ori_ori_n225_), .Y(ori_ori_n228_));
  AN4        o0200(.A(ori_ori_n228_), .B(ori_ori_n223_), .C(ori_ori_n217_), .D(ori_ori_n211_), .Y(ori_ori_n229_));
  NO2        o0201(.A(h), .B(ori_ori_n94_), .Y(ori_ori_n230_));
  NA2        o0202(.A(ori_ori_n230_), .B(ori_ori_n119_), .Y(ori_ori_n231_));
  NAi41      o0203(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n232_));
  NO2        o0204(.A(ori_ori_n232_), .B(ori_ori_n200_), .Y(ori_ori_n233_));
  NA2        o0205(.A(ori_ori_n149_), .B(ori_ori_n99_), .Y(ori_ori_n234_));
  NO2        o0206(.A(n), .B(a), .Y(ori_ori_n235_));
  NAi31      o0207(.An(ori_ori_n226_), .B(ori_ori_n235_), .C(ori_ori_n95_), .Y(ori_ori_n236_));
  NAi21      o0208(.An(h), .B(i), .Y(ori_ori_n237_));
  NA2        o0209(.A(ori_ori_n168_), .B(k), .Y(ori_ori_n238_));
  NO2        o0210(.A(ori_ori_n238_), .B(ori_ori_n237_), .Y(ori_ori_n239_));
  NA2        o0211(.A(ori_ori_n239_), .B(ori_ori_n177_), .Y(ori_ori_n240_));
  NA3        o0212(.A(ori_ori_n240_), .B(ori_ori_n236_), .C(ori_ori_n231_), .Y(ori_ori_n241_));
  NOi21      o0213(.An(g), .B(e), .Y(ori_ori_n242_));
  NO2        o0214(.A(ori_ori_n66_), .B(ori_ori_n67_), .Y(ori_ori_n243_));
  NOi32      o0215(.An(l), .Bn(j), .C(i), .Y(ori_ori_n244_));
  AOI210     o0216(.A0(ori_ori_n68_), .A1(ori_ori_n78_), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NO2        o0217(.A(ori_ori_n237_), .B(ori_ori_n43_), .Y(ori_ori_n246_));
  NAi21      o0218(.An(f), .B(g), .Y(ori_ori_n247_));
  NO2        o0219(.A(ori_ori_n247_), .B(ori_ori_n60_), .Y(ori_ori_n248_));
  NO2        o0220(.A(ori_ori_n63_), .B(ori_ori_n106_), .Y(ori_ori_n249_));
  AOI220     o0221(.A0(ori_ori_n249_), .A1(ori_ori_n248_), .B0(ori_ori_n246_), .B1(ori_ori_n62_), .Y(ori_ori_n250_));
  INV        o0222(.A(ori_ori_n250_), .Y(ori_ori_n251_));
  NOi41      o0223(.An(ori_ori_n229_), .B(ori_ori_n251_), .C(ori_ori_n241_), .D(ori_ori_n207_), .Y(ori_ori_n252_));
  NO3        o0224(.A(ori_ori_n188_), .B(ori_ori_n47_), .C(ori_ori_n42_), .Y(ori_ori_n253_));
  NO2        o0225(.A(ori_ori_n253_), .B(ori_ori_n101_), .Y(ori_ori_n254_));
  NA3        o0226(.A(ori_ori_n58_), .B(c), .C(b), .Y(ori_ori_n255_));
  OR4        o0227(.A(h), .B(ori_ori_n255_), .C(ori_ori_n210_), .D(e), .Y(ori_ori_n256_));
  NO2        o0228(.A(ori_ori_n234_), .B(ori_ori_n247_), .Y(ori_ori_n257_));
  NAi31      o0229(.An(g), .B(k), .C(h), .Y(ori_ori_n258_));
  NO3        o0230(.A(ori_ori_n121_), .B(ori_ori_n258_), .C(l), .Y(ori_ori_n259_));
  NAi31      o0231(.An(e), .B(d), .C(a), .Y(ori_ori_n260_));
  NA2        o0232(.A(ori_ori_n259_), .B(ori_ori_n119_), .Y(ori_ori_n261_));
  NA2        o0233(.A(ori_ori_n261_), .B(ori_ori_n256_), .Y(ori_ori_n262_));
  NA3        o0234(.A(ori_ori_n149_), .B(ori_ori_n148_), .C(ori_ori_n75_), .Y(ori_ori_n263_));
  NO2        o0235(.A(ori_ori_n263_), .B(ori_ori_n179_), .Y(ori_ori_n264_));
  INV        o0236(.A(ori_ori_n264_), .Y(ori_ori_n265_));
  NA3        o0237(.A(e), .B(c), .C(b), .Y(ori_ori_n266_));
  NAi32      o0238(.An(k), .Bn(i), .C(j), .Y(ori_ori_n267_));
  INV        o0239(.A(ori_ori_n48_), .Y(ori_ori_n268_));
  NA2        o0240(.A(ori_ori_n248_), .B(ori_ori_n268_), .Y(ori_ori_n269_));
  NAi21      o0241(.An(l), .B(k), .Y(ori_ori_n270_));
  NOi21      o0242(.An(l), .B(j), .Y(ori_ori_n271_));
  NA2        o0243(.A(ori_ori_n152_), .B(ori_ori_n271_), .Y(ori_ori_n272_));
  NAi32      o0244(.An(j), .Bn(h), .C(i), .Y(ori_ori_n273_));
  NAi21      o0245(.An(m), .B(l), .Y(ori_ori_n274_));
  NO3        o0246(.A(ori_ori_n274_), .B(ori_ori_n273_), .C(ori_ori_n75_), .Y(ori_ori_n275_));
  NA2        o0247(.A(h), .B(g), .Y(ori_ori_n276_));
  NA2        o0248(.A(ori_ori_n157_), .B(ori_ori_n44_), .Y(ori_ori_n277_));
  NO2        o0249(.A(ori_ori_n277_), .B(ori_ori_n276_), .Y(ori_ori_n278_));
  OAI210     o0250(.A0(ori_ori_n278_), .A1(ori_ori_n275_), .B0(ori_ori_n153_), .Y(ori_ori_n279_));
  NA3        o0251(.A(ori_ori_n279_), .B(ori_ori_n269_), .C(ori_ori_n265_), .Y(ori_ori_n280_));
  NO2        o0252(.A(ori_ori_n133_), .B(d), .Y(ori_ori_n281_));
  NO2        o0253(.A(ori_ori_n97_), .B(ori_ori_n94_), .Y(ori_ori_n282_));
  NAi32      o0254(.An(n), .Bn(m), .C(l), .Y(ori_ori_n283_));
  NO2        o0255(.A(ori_ori_n283_), .B(ori_ori_n273_), .Y(ori_ori_n284_));
  NA2        o0256(.A(ori_ori_n284_), .B(ori_ori_n172_), .Y(ori_ori_n285_));
  NAi31      o0257(.An(k), .B(l), .C(j), .Y(ori_ori_n286_));
  OAI210     o0258(.A0(ori_ori_n270_), .A1(j), .B0(ori_ori_n286_), .Y(ori_ori_n287_));
  NOi21      o0259(.An(ori_ori_n287_), .B(ori_ori_n109_), .Y(ori_ori_n288_));
  INV        o0260(.A(ori_ori_n285_), .Y(ori_ori_n289_));
  NO4        o0261(.A(ori_ori_n289_), .B(ori_ori_n280_), .C(ori_ori_n262_), .D(ori_ori_n254_), .Y(ori_ori_n290_));
  NA2        o0262(.A(ori_ori_n239_), .B(ori_ori_n178_), .Y(ori_ori_n291_));
  NAi21      o0263(.An(m), .B(k), .Y(ori_ori_n292_));
  NO2        o0264(.A(ori_ori_n213_), .B(ori_ori_n292_), .Y(ori_ori_n293_));
  NAi41      o0265(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n294_));
  NO2        o0266(.A(ori_ori_n294_), .B(ori_ori_n139_), .Y(ori_ori_n295_));
  NA2        o0267(.A(ori_ori_n295_), .B(ori_ori_n293_), .Y(ori_ori_n296_));
  NO4        o0268(.A(i), .B(ori_ori_n139_), .C(ori_ori_n66_), .D(ori_ori_n67_), .Y(ori_ori_n297_));
  NA2        o0269(.A(e), .B(c), .Y(ori_ori_n298_));
  NO3        o0270(.A(ori_ori_n298_), .B(n), .C(d), .Y(ori_ori_n299_));
  NAi31      o0271(.An(d), .B(e), .C(b), .Y(ori_ori_n300_));
  NAi31      o0272(.An(ori_ori_n297_), .B(ori_ori_n296_), .C(ori_ori_n291_), .Y(ori_ori_n301_));
  NO4        o0273(.A(ori_ori_n294_), .B(ori_ori_n73_), .C(ori_ori_n65_), .D(ori_ori_n201_), .Y(ori_ori_n302_));
  NA2        o0274(.A(ori_ori_n235_), .B(ori_ori_n95_), .Y(ori_ori_n303_));
  NOi31      o0275(.An(l), .B(n), .C(m), .Y(ori_ori_n304_));
  NAi32      o0276(.An(m), .Bn(j), .C(k), .Y(ori_ori_n305_));
  NAi41      o0277(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n306_));
  NOi31      o0278(.An(j), .B(m), .C(k), .Y(ori_ori_n307_));
  NO2        o0279(.A(ori_ori_n114_), .B(ori_ori_n307_), .Y(ori_ori_n308_));
  AN3        o0280(.A(h), .B(g), .C(f), .Y(ori_ori_n309_));
  NOi32      o0281(.An(m), .Bn(j), .C(l), .Y(ori_ori_n310_));
  NO2        o0282(.A(ori_ori_n310_), .B(ori_ori_n89_), .Y(ori_ori_n311_));
  NAi32      o0283(.An(ori_ori_n311_), .Bn(ori_ori_n187_), .C(ori_ori_n281_), .Y(ori_ori_n312_));
  NO2        o0284(.A(ori_ori_n274_), .B(ori_ori_n273_), .Y(ori_ori_n313_));
  NO2        o0285(.A(ori_ori_n204_), .B(g), .Y(ori_ori_n314_));
  NO2        o0286(.A(ori_ori_n145_), .B(ori_ori_n75_), .Y(ori_ori_n315_));
  AOI220     o0287(.A0(ori_ori_n315_), .A1(ori_ori_n314_), .B0(ori_ori_n233_), .B1(ori_ori_n313_), .Y(ori_ori_n316_));
  INV        o0288(.A(ori_ori_n221_), .Y(ori_ori_n317_));
  NA3        o0289(.A(ori_ori_n317_), .B(ori_ori_n309_), .C(ori_ori_n199_), .Y(ori_ori_n318_));
  NA3        o0290(.A(ori_ori_n318_), .B(ori_ori_n316_), .C(ori_ori_n312_), .Y(ori_ori_n319_));
  NA3        o0291(.A(h), .B(g), .C(f), .Y(ori_ori_n320_));
  NO2        o0292(.A(ori_ori_n320_), .B(ori_ori_n69_), .Y(ori_ori_n321_));
  NA2        o0293(.A(ori_ori_n152_), .B(e), .Y(ori_ori_n322_));
  NO2        o0294(.A(ori_ori_n322_), .B(ori_ori_n40_), .Y(ori_ori_n323_));
  NOi32      o0295(.An(j), .Bn(g), .C(i), .Y(ori_ori_n324_));
  NA3        o0296(.A(ori_ori_n324_), .B(ori_ori_n270_), .C(ori_ori_n103_), .Y(ori_ori_n325_));
  AO210      o0297(.A0(ori_ori_n101_), .A1(ori_ori_n32_), .B0(ori_ori_n325_), .Y(ori_ori_n326_));
  NOi32      o0298(.An(e), .Bn(b), .C(a), .Y(ori_ori_n327_));
  AN2        o0299(.A(l), .B(j), .Y(ori_ori_n328_));
  NO2        o0300(.A(ori_ori_n292_), .B(ori_ori_n328_), .Y(ori_ori_n329_));
  NO3        o0301(.A(ori_ori_n294_), .B(ori_ori_n65_), .C(ori_ori_n201_), .Y(ori_ori_n330_));
  NA3        o0302(.A(ori_ori_n195_), .B(ori_ori_n193_), .C(ori_ori_n35_), .Y(ori_ori_n331_));
  AOI220     o0303(.A0(ori_ori_n331_), .A1(ori_ori_n327_), .B0(ori_ori_n330_), .B1(ori_ori_n329_), .Y(ori_ori_n332_));
  NO2        o0304(.A(ori_ori_n300_), .B(n), .Y(ori_ori_n333_));
  NA2        o0305(.A(ori_ori_n194_), .B(k), .Y(ori_ori_n334_));
  NA3        o0306(.A(m), .B(ori_ori_n102_), .C(ori_ori_n200_), .Y(ori_ori_n335_));
  NA4        o0307(.A(ori_ori_n189_), .B(ori_ori_n78_), .C(g), .D(ori_ori_n200_), .Y(ori_ori_n336_));
  OAI210     o0308(.A0(ori_ori_n335_), .A1(ori_ori_n334_), .B0(ori_ori_n336_), .Y(ori_ori_n337_));
  NAi41      o0309(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n338_));
  NA2        o0310(.A(ori_ori_n50_), .B(ori_ori_n103_), .Y(ori_ori_n339_));
  NO2        o0311(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  NA2        o0312(.A(ori_ori_n337_), .B(ori_ori_n333_), .Y(ori_ori_n341_));
  NA3        o0313(.A(ori_ori_n341_), .B(ori_ori_n332_), .C(ori_ori_n326_), .Y(ori_ori_n342_));
  NO4        o0314(.A(ori_ori_n342_), .B(ori_ori_n319_), .C(ori_ori_n302_), .D(ori_ori_n301_), .Y(ori_ori_n343_));
  NA4        o0315(.A(ori_ori_n343_), .B(ori_ori_n290_), .C(ori_ori_n252_), .D(ori_ori_n185_), .Y(ori10));
  NA3        o0316(.A(m), .B(k), .C(i), .Y(ori_ori_n345_));
  NO3        o0317(.A(ori_ori_n345_), .B(j), .C(ori_ori_n201_), .Y(ori_ori_n346_));
  NOi21      o0318(.An(e), .B(f), .Y(ori_ori_n347_));
  NO4        o0319(.A(ori_ori_n140_), .B(ori_ori_n347_), .C(n), .D(ori_ori_n100_), .Y(ori_ori_n348_));
  NAi31      o0320(.An(b), .B(f), .C(c), .Y(ori_ori_n349_));
  INV        o0321(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NOi32      o0322(.An(k), .Bn(h), .C(j), .Y(ori_ori_n351_));
  NA2        o0323(.A(ori_ori_n351_), .B(ori_ori_n208_), .Y(ori_ori_n352_));
  NA2        o0324(.A(ori_ori_n150_), .B(ori_ori_n352_), .Y(ori_ori_n353_));
  AOI220     o0325(.A0(ori_ori_n353_), .A1(ori_ori_n350_), .B0(ori_ori_n348_), .B1(ori_ori_n346_), .Y(ori_ori_n354_));
  AN2        o0326(.A(j), .B(h), .Y(ori_ori_n355_));
  NO3        o0327(.A(n), .B(m), .C(k), .Y(ori_ori_n356_));
  NA2        o0328(.A(ori_ori_n356_), .B(ori_ori_n355_), .Y(ori_ori_n357_));
  NO3        o0329(.A(ori_ori_n357_), .B(ori_ori_n140_), .C(ori_ori_n200_), .Y(ori_ori_n358_));
  OR2        o0330(.A(m), .B(k), .Y(ori_ori_n359_));
  NO2        o0331(.A(ori_ori_n162_), .B(ori_ori_n359_), .Y(ori_ori_n360_));
  NA4        o0332(.A(n), .B(f), .C(c), .D(ori_ori_n105_), .Y(ori_ori_n361_));
  NOi21      o0333(.An(ori_ori_n360_), .B(ori_ori_n361_), .Y(ori_ori_n362_));
  NOi32      o0334(.An(d), .Bn(a), .C(c), .Y(ori_ori_n363_));
  NA2        o0335(.A(ori_ori_n363_), .B(ori_ori_n170_), .Y(ori_ori_n364_));
  NAi21      o0336(.An(i), .B(g), .Y(ori_ori_n365_));
  NAi31      o0337(.An(k), .B(m), .C(j), .Y(ori_ori_n366_));
  NO3        o0338(.A(ori_ori_n366_), .B(ori_ori_n365_), .C(n), .Y(ori_ori_n367_));
  NOi21      o0339(.An(ori_ori_n367_), .B(ori_ori_n364_), .Y(ori_ori_n368_));
  NO3        o0340(.A(ori_ori_n368_), .B(ori_ori_n362_), .C(ori_ori_n358_), .Y(ori_ori_n369_));
  NO2        o0341(.A(ori_ori_n361_), .B(ori_ori_n274_), .Y(ori_ori_n370_));
  NOi32      o0342(.An(f), .Bn(d), .C(c), .Y(ori_ori_n371_));
  AOI220     o0343(.A0(ori_ori_n371_), .A1(ori_ori_n284_), .B0(ori_ori_n370_), .B1(ori_ori_n202_), .Y(ori_ori_n372_));
  NA3        o0344(.A(ori_ori_n372_), .B(ori_ori_n369_), .C(ori_ori_n354_), .Y(ori_ori_n373_));
  NO2        o0345(.A(ori_ori_n58_), .B(ori_ori_n105_), .Y(ori_ori_n374_));
  NA2        o0346(.A(ori_ori_n235_), .B(ori_ori_n374_), .Y(ori_ori_n375_));
  INV        o0347(.A(e), .Y(ori_ori_n376_));
  NA2        o0348(.A(ori_ori_n45_), .B(e), .Y(ori_ori_n377_));
  OAI220     o0349(.A0(ori_ori_n377_), .A1(ori_ori_n186_), .B0(ori_ori_n190_), .B1(ori_ori_n376_), .Y(ori_ori_n378_));
  NO2        o0350(.A(ori_ori_n80_), .B(ori_ori_n376_), .Y(ori_ori_n379_));
  NO2        o0351(.A(ori_ori_n91_), .B(ori_ori_n376_), .Y(ori_ori_n380_));
  NO3        o0352(.A(ori_ori_n380_), .B(ori_ori_n379_), .C(ori_ori_n378_), .Y(ori_ori_n381_));
  NOi32      o0353(.An(h), .Bn(e), .C(g), .Y(ori_ori_n382_));
  AN3        o0354(.A(h), .B(g), .C(e), .Y(ori_ori_n383_));
  NO2        o0355(.A(ori_ori_n381_), .B(ori_ori_n375_), .Y(ori_ori_n384_));
  NAi31      o0356(.An(b), .B(c), .C(a), .Y(ori_ori_n385_));
  NO2        o0357(.A(ori_ori_n385_), .B(n), .Y(ori_ori_n386_));
  NA2        o0358(.A(ori_ori_n50_), .B(m), .Y(ori_ori_n387_));
  NO2        o0359(.A(ori_ori_n387_), .B(ori_ori_n136_), .Y(ori_ori_n388_));
  NA2        o0360(.A(ori_ori_n388_), .B(ori_ori_n386_), .Y(ori_ori_n389_));
  INV        o0361(.A(ori_ori_n389_), .Y(ori_ori_n390_));
  NO3        o0362(.A(ori_ori_n390_), .B(ori_ori_n384_), .C(ori_ori_n373_), .Y(ori_ori_n391_));
  NA2        o0363(.A(i), .B(g), .Y(ori_ori_n392_));
  NOi21      o0364(.An(a), .B(n), .Y(ori_ori_n393_));
  NOi21      o0365(.An(d), .B(c), .Y(ori_ori_n394_));
  NA2        o0366(.A(ori_ori_n394_), .B(ori_ori_n393_), .Y(ori_ori_n395_));
  NA3        o0367(.A(i), .B(g), .C(f), .Y(ori_ori_n396_));
  OR2        o0368(.A(n), .B(m), .Y(ori_ori_n397_));
  NO2        o0369(.A(ori_ori_n397_), .B(ori_ori_n141_), .Y(ori_ori_n398_));
  NO2        o0370(.A(ori_ori_n171_), .B(ori_ori_n136_), .Y(ori_ori_n399_));
  OAI210     o0371(.A0(ori_ori_n398_), .A1(ori_ori_n164_), .B0(ori_ori_n399_), .Y(ori_ori_n400_));
  INV        o0372(.A(ori_ori_n339_), .Y(ori_ori_n401_));
  NA3        o0373(.A(ori_ori_n401_), .B(ori_ori_n327_), .C(d), .Y(ori_ori_n402_));
  NO2        o0374(.A(ori_ori_n385_), .B(ori_ori_n48_), .Y(ori_ori_n403_));
  NAi21      o0375(.An(k), .B(j), .Y(ori_ori_n404_));
  NAi21      o0376(.An(e), .B(d), .Y(ori_ori_n405_));
  INV        o0377(.A(ori_ori_n405_), .Y(ori_ori_n406_));
  NO2        o0378(.A(ori_ori_n238_), .B(ori_ori_n200_), .Y(ori_ori_n407_));
  NA3        o0379(.A(ori_ori_n407_), .B(ori_ori_n406_), .C(ori_ori_n214_), .Y(ori_ori_n408_));
  NA3        o0380(.A(ori_ori_n408_), .B(ori_ori_n402_), .C(ori_ori_n400_), .Y(ori_ori_n409_));
  NOi31      o0381(.An(n), .B(m), .C(k), .Y(ori_ori_n410_));
  AOI220     o0382(.A0(ori_ori_n410_), .A1(ori_ori_n355_), .B0(ori_ori_n208_), .B1(ori_ori_n49_), .Y(ori_ori_n411_));
  NAi31      o0383(.An(g), .B(f), .C(c), .Y(ori_ori_n412_));
  OR3        o0384(.A(ori_ori_n412_), .B(ori_ori_n411_), .C(e), .Y(ori_ori_n413_));
  NA2        o0385(.A(ori_ori_n413_), .B(ori_ori_n285_), .Y(ori_ori_n414_));
  NO3        o0386(.A(ori_ori_n414_), .B(ori_ori_n409_), .C(ori_ori_n251_), .Y(ori_ori_n415_));
  NOi32      o0387(.An(c), .Bn(a), .C(b), .Y(ori_ori_n416_));
  NA2        o0388(.A(ori_ori_n416_), .B(ori_ori_n103_), .Y(ori_ori_n417_));
  AN2        o0389(.A(e), .B(d), .Y(ori_ori_n418_));
  INV        o0390(.A(ori_ori_n136_), .Y(ori_ori_n419_));
  NO2        o0391(.A(ori_ori_n120_), .B(ori_ori_n40_), .Y(ori_ori_n420_));
  NO2        o0392(.A(ori_ori_n61_), .B(e), .Y(ori_ori_n421_));
  NOi31      o0393(.An(j), .B(k), .C(i), .Y(ori_ori_n422_));
  NOi21      o0394(.An(ori_ori_n154_), .B(ori_ori_n422_), .Y(ori_ori_n423_));
  NA3        o0395(.A(ori_ori_n423_), .B(ori_ori_n245_), .C(ori_ori_n108_), .Y(ori_ori_n424_));
  AOI220     o0396(.A0(ori_ori_n424_), .A1(ori_ori_n421_), .B0(ori_ori_n420_), .B1(ori_ori_n419_), .Y(ori_ori_n425_));
  NO2        o0397(.A(ori_ori_n425_), .B(ori_ori_n417_), .Y(ori_ori_n426_));
  NO2        o0398(.A(ori_ori_n196_), .B(ori_ori_n191_), .Y(ori_ori_n427_));
  NOi21      o0399(.An(a), .B(b), .Y(ori_ori_n428_));
  NA3        o0400(.A(e), .B(d), .C(c), .Y(ori_ori_n429_));
  NAi21      o0401(.An(ori_ori_n429_), .B(ori_ori_n428_), .Y(ori_ori_n430_));
  AOI210     o0402(.A0(ori_ori_n253_), .A1(ori_ori_n427_), .B0(ori_ori_n430_), .Y(ori_ori_n431_));
  NO4        o0403(.A(ori_ori_n175_), .B(ori_ori_n94_), .C(ori_ori_n55_), .D(b), .Y(ori_ori_n432_));
  NA2        o0404(.A(ori_ori_n350_), .B(ori_ori_n142_), .Y(ori_ori_n433_));
  OR2        o0405(.A(k), .B(j), .Y(ori_ori_n434_));
  NA2        o0406(.A(l), .B(k), .Y(ori_ori_n435_));
  NA3        o0407(.A(ori_ori_n435_), .B(ori_ori_n434_), .C(ori_ori_n208_), .Y(ori_ori_n436_));
  AOI210     o0408(.A0(ori_ori_n221_), .A1(ori_ori_n305_), .B0(ori_ori_n75_), .Y(ori_ori_n437_));
  NOi21      o0409(.An(ori_ori_n436_), .B(ori_ori_n437_), .Y(ori_ori_n438_));
  OR3        o0410(.A(ori_ori_n438_), .B(ori_ori_n132_), .C(ori_ori_n122_), .Y(ori_ori_n439_));
  NA2        o0411(.A(ori_ori_n117_), .B(ori_ori_n115_), .Y(ori_ori_n440_));
  NO2        o0412(.A(ori_ori_n440_), .B(ori_ori_n297_), .Y(ori_ori_n441_));
  NA3        o0413(.A(ori_ori_n441_), .B(ori_ori_n439_), .C(ori_ori_n433_), .Y(ori_ori_n442_));
  NO4        o0414(.A(ori_ori_n442_), .B(ori_ori_n432_), .C(ori_ori_n431_), .D(ori_ori_n426_), .Y(ori_ori_n443_));
  INV        o0415(.A(e), .Y(ori_ori_n444_));
  NO2        o0416(.A(ori_ori_n175_), .B(ori_ori_n55_), .Y(ori_ori_n445_));
  NAi31      o0417(.An(j), .B(l), .C(i), .Y(ori_ori_n446_));
  OAI210     o0418(.A0(ori_ori_n446_), .A1(ori_ori_n121_), .B0(ori_ori_n94_), .Y(ori_ori_n447_));
  NA3        o0419(.A(ori_ori_n447_), .B(ori_ori_n445_), .C(ori_ori_n444_), .Y(ori_ori_n448_));
  NO3        o0420(.A(ori_ori_n364_), .B(ori_ori_n311_), .C(ori_ori_n187_), .Y(ori_ori_n449_));
  NO2        o0421(.A(ori_ori_n364_), .B(ori_ori_n339_), .Y(ori_ori_n450_));
  NO4        o0422(.A(ori_ori_n450_), .B(ori_ori_n449_), .C(ori_ori_n173_), .D(ori_ori_n282_), .Y(ori_ori_n451_));
  NA3        o0423(.A(ori_ori_n451_), .B(ori_ori_n448_), .C(ori_ori_n229_), .Y(ori_ori_n452_));
  OAI210     o0424(.A0(ori_ori_n116_), .A1(ori_ori_n114_), .B0(n), .Y(ori_ori_n453_));
  NO2        o0425(.A(ori_ori_n453_), .B(ori_ori_n120_), .Y(ori_ori_n454_));
  XO2        o0426(.A(i), .B(h), .Y(ori_ori_n455_));
  NA3        o0427(.A(ori_ori_n455_), .B(ori_ori_n149_), .C(n), .Y(ori_ori_n456_));
  NAi41      o0428(.An(ori_ori_n275_), .B(ori_ori_n456_), .C(ori_ori_n411_), .D(ori_ori_n352_), .Y(ori_ori_n457_));
  NOi32      o0429(.An(ori_ori_n457_), .Bn(ori_ori_n421_), .C(ori_ori_n255_), .Y(ori_ori_n458_));
  NAi31      o0430(.An(c), .B(f), .C(d), .Y(ori_ori_n459_));
  AOI210     o0431(.A0(ori_ori_n263_), .A1(ori_ori_n181_), .B0(ori_ori_n459_), .Y(ori_ori_n460_));
  INV        o0432(.A(ori_ori_n460_), .Y(ori_ori_n461_));
  NA2        o0433(.A(ori_ori_n215_), .B(ori_ori_n99_), .Y(ori_ori_n462_));
  AOI210     o0434(.A0(ori_ori_n462_), .A1(ori_ori_n169_), .B0(ori_ori_n459_), .Y(ori_ori_n463_));
  NO2        o0435(.A(ori_ori_n325_), .B(ori_ori_n430_), .Y(ori_ori_n464_));
  NO2        o0436(.A(ori_ori_n464_), .B(ori_ori_n463_), .Y(ori_ori_n465_));
  AO220      o0437(.A0(ori_ori_n268_), .A1(ori_ori_n248_), .B0(ori_ori_n155_), .B1(ori_ori_n62_), .Y(ori_ori_n466_));
  NA3        o0438(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n467_));
  NO2        o0439(.A(ori_ori_n467_), .B(ori_ori_n395_), .Y(ori_ori_n468_));
  INV        o0440(.A(ori_ori_n468_), .Y(ori_ori_n469_));
  NAi41      o0441(.An(ori_ori_n466_), .B(ori_ori_n469_), .C(ori_ori_n465_), .D(ori_ori_n461_), .Y(ori_ori_n470_));
  NO3        o0442(.A(ori_ori_n470_), .B(ori_ori_n458_), .C(ori_ori_n452_), .Y(ori_ori_n471_));
  NA4        o0443(.A(ori_ori_n471_), .B(ori_ori_n443_), .C(ori_ori_n415_), .D(ori_ori_n391_), .Y(ori11));
  NO2        o0444(.A(ori_ori_n66_), .B(f), .Y(ori_ori_n473_));
  NA2        o0445(.A(j), .B(g), .Y(ori_ori_n474_));
  NAi31      o0446(.An(i), .B(m), .C(l), .Y(ori_ori_n475_));
  NA3        o0447(.A(m), .B(k), .C(j), .Y(ori_ori_n476_));
  OAI220     o0448(.A0(ori_ori_n476_), .A1(ori_ori_n120_), .B0(ori_ori_n475_), .B1(ori_ori_n474_), .Y(ori_ori_n477_));
  NA2        o0449(.A(ori_ori_n477_), .B(ori_ori_n473_), .Y(ori_ori_n478_));
  NOi32      o0450(.An(e), .Bn(b), .C(f), .Y(ori_ori_n479_));
  NA2        o0451(.A(ori_ori_n45_), .B(j), .Y(ori_ori_n480_));
  NO2        o0452(.A(ori_ori_n480_), .B(ori_ori_n277_), .Y(ori_ori_n481_));
  NAi31      o0453(.An(d), .B(e), .C(a), .Y(ori_ori_n482_));
  NO2        o0454(.A(ori_ori_n482_), .B(n), .Y(ori_ori_n483_));
  AOI220     o0455(.A0(ori_ori_n483_), .A1(ori_ori_n92_), .B0(ori_ori_n481_), .B1(ori_ori_n479_), .Y(ori_ori_n484_));
  NAi31      o0456(.An(f), .B(e), .C(a), .Y(ori_ori_n485_));
  AN2        o0457(.A(ori_ori_n485_), .B(ori_ori_n338_), .Y(ori_ori_n486_));
  NA2        o0458(.A(j), .B(i), .Y(ori_ori_n487_));
  NAi31      o0459(.An(n), .B(m), .C(k), .Y(ori_ori_n488_));
  NO3        o0460(.A(ori_ori_n488_), .B(ori_ori_n487_), .C(ori_ori_n102_), .Y(ori_ori_n489_));
  NO4        o0461(.A(n), .B(d), .C(ori_ori_n105_), .D(a), .Y(ori_ori_n490_));
  OR2        o0462(.A(n), .B(c), .Y(ori_ori_n491_));
  NO2        o0463(.A(ori_ori_n491_), .B(ori_ori_n138_), .Y(ori_ori_n492_));
  NO2        o0464(.A(ori_ori_n492_), .B(ori_ori_n490_), .Y(ori_ori_n493_));
  NOi32      o0465(.An(g), .Bn(f), .C(i), .Y(ori_ori_n494_));
  AOI220     o0466(.A0(ori_ori_n494_), .A1(ori_ori_n90_), .B0(ori_ori_n477_), .B1(f), .Y(ori_ori_n495_));
  NO2        o0467(.A(ori_ori_n258_), .B(ori_ori_n48_), .Y(ori_ori_n496_));
  NO2        o0468(.A(ori_ori_n495_), .B(ori_ori_n493_), .Y(ori_ori_n497_));
  INV        o0469(.A(ori_ori_n497_), .Y(ori_ori_n498_));
  NA2        o0470(.A(ori_ori_n128_), .B(ori_ori_n34_), .Y(ori_ori_n499_));
  OAI220     o0471(.A0(ori_ori_n499_), .A1(m), .B0(ori_ori_n480_), .B1(ori_ori_n221_), .Y(ori_ori_n500_));
  NOi41      o0472(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n501_));
  NAi32      o0473(.An(e), .Bn(b), .C(c), .Y(ori_ori_n502_));
  OR2        o0474(.A(ori_ori_n502_), .B(ori_ori_n75_), .Y(ori_ori_n503_));
  AN2        o0475(.A(ori_ori_n306_), .B(ori_ori_n294_), .Y(ori_ori_n504_));
  NA2        o0476(.A(ori_ori_n504_), .B(ori_ori_n503_), .Y(ori_ori_n505_));
  AN2        o0477(.A(ori_ori_n505_), .B(ori_ori_n500_), .Y(ori_ori_n506_));
  OAI220     o0478(.A0(ori_ori_n366_), .A1(ori_ori_n365_), .B0(ori_ori_n475_), .B1(ori_ori_n474_), .Y(ori_ori_n507_));
  NAi31      o0479(.An(d), .B(c), .C(a), .Y(ori_ori_n508_));
  NO2        o0480(.A(ori_ori_n508_), .B(n), .Y(ori_ori_n509_));
  NO2        o0481(.A(ori_ori_n218_), .B(ori_ori_n100_), .Y(ori_ori_n510_));
  NA2        o0482(.A(ori_ori_n367_), .B(ori_ori_n510_), .Y(ori_ori_n511_));
  INV        o0483(.A(ori_ori_n511_), .Y(ori_ori_n512_));
  NO2        o0484(.A(ori_ori_n260_), .B(n), .Y(ori_ori_n513_));
  NO2        o0485(.A(ori_ori_n386_), .B(ori_ori_n513_), .Y(ori_ori_n514_));
  NA2        o0486(.A(ori_ori_n507_), .B(f), .Y(ori_ori_n515_));
  NAi32      o0487(.An(d), .Bn(a), .C(b), .Y(ori_ori_n516_));
  NO2        o0488(.A(ori_ori_n516_), .B(ori_ori_n48_), .Y(ori_ori_n517_));
  NA2        o0489(.A(h), .B(f), .Y(ori_ori_n518_));
  NO2        o0490(.A(ori_ori_n518_), .B(ori_ori_n86_), .Y(ori_ori_n519_));
  NO3        o0491(.A(ori_ori_n165_), .B(ori_ori_n162_), .C(g), .Y(ori_ori_n520_));
  AOI220     o0492(.A0(ori_ori_n520_), .A1(ori_ori_n57_), .B0(ori_ori_n519_), .B1(ori_ori_n517_), .Y(ori_ori_n521_));
  OAI210     o0493(.A0(ori_ori_n515_), .A1(ori_ori_n514_), .B0(ori_ori_n521_), .Y(ori_ori_n522_));
  AN3        o0494(.A(j), .B(h), .C(g), .Y(ori_ori_n523_));
  NO2        o0495(.A(ori_ori_n135_), .B(c), .Y(ori_ori_n524_));
  NA3        o0496(.A(ori_ori_n524_), .B(ori_ori_n523_), .C(ori_ori_n410_), .Y(ori_ori_n525_));
  NA3        o0497(.A(f), .B(d), .C(b), .Y(ori_ori_n526_));
  NO4        o0498(.A(ori_ori_n526_), .B(ori_ori_n165_), .C(ori_ori_n162_), .D(g), .Y(ori_ori_n527_));
  NAi21      o0499(.An(ori_ori_n527_), .B(ori_ori_n525_), .Y(ori_ori_n528_));
  NO4        o0500(.A(ori_ori_n528_), .B(ori_ori_n522_), .C(ori_ori_n512_), .D(ori_ori_n506_), .Y(ori_ori_n529_));
  AN4        o0501(.A(ori_ori_n529_), .B(ori_ori_n498_), .C(ori_ori_n484_), .D(ori_ori_n478_), .Y(ori_ori_n530_));
  INV        o0502(.A(k), .Y(ori_ori_n531_));
  NA3        o0503(.A(l), .B(ori_ori_n531_), .C(i), .Y(ori_ori_n532_));
  INV        o0504(.A(ori_ori_n532_), .Y(ori_ori_n533_));
  NAi32      o0505(.An(h), .Bn(f), .C(g), .Y(ori_ori_n534_));
  NAi41      o0506(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n535_));
  OAI210     o0507(.A0(ori_ori_n482_), .A1(n), .B0(ori_ori_n535_), .Y(ori_ori_n536_));
  NA2        o0508(.A(ori_ori_n536_), .B(m), .Y(ori_ori_n537_));
  NAi31      o0509(.An(h), .B(g), .C(f), .Y(ori_ori_n538_));
  NO3        o0510(.A(ori_ori_n534_), .B(ori_ori_n66_), .C(ori_ori_n67_), .Y(ori_ori_n539_));
  NO4        o0511(.A(ori_ori_n538_), .B(ori_ori_n491_), .C(ori_ori_n138_), .D(ori_ori_n67_), .Y(ori_ori_n540_));
  OR2        o0512(.A(ori_ori_n540_), .B(ori_ori_n539_), .Y(ori_ori_n541_));
  NAi31      o0513(.An(f), .B(h), .C(g), .Y(ori_ori_n542_));
  NOi32      o0514(.An(b), .Bn(a), .C(c), .Y(ori_ori_n543_));
  NOi32      o0515(.An(d), .Bn(a), .C(e), .Y(ori_ori_n544_));
  NA2        o0516(.A(ori_ori_n544_), .B(ori_ori_n103_), .Y(ori_ori_n545_));
  NO2        o0517(.A(n), .B(c), .Y(ori_ori_n546_));
  NA3        o0518(.A(ori_ori_n546_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n547_));
  NA2        o0519(.A(ori_ori_n547_), .B(ori_ori_n545_), .Y(ori_ori_n548_));
  NOi32      o0520(.An(e), .Bn(a), .C(d), .Y(ori_ori_n549_));
  AOI210     o0521(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n549_), .Y(ori_ori_n550_));
  INV        o0522(.A(ori_ori_n499_), .Y(ori_ori_n551_));
  NA2        o0523(.A(ori_ori_n551_), .B(ori_ori_n548_), .Y(ori_ori_n552_));
  INV        o0524(.A(ori_ori_n552_), .Y(ori_ori_n553_));
  AOI210     o0525(.A0(ori_ori_n541_), .A1(ori_ori_n533_), .B0(ori_ori_n553_), .Y(ori_ori_n554_));
  NO3        o0526(.A(ori_ori_n292_), .B(ori_ori_n59_), .C(n), .Y(ori_ori_n555_));
  NA3        o0527(.A(ori_ori_n459_), .B(ori_ori_n160_), .C(ori_ori_n159_), .Y(ori_ori_n556_));
  NA2        o0528(.A(ori_ori_n412_), .B(ori_ori_n218_), .Y(ori_ori_n557_));
  OR2        o0529(.A(ori_ori_n557_), .B(ori_ori_n556_), .Y(ori_ori_n558_));
  NA2        o0530(.A(ori_ori_n558_), .B(ori_ori_n555_), .Y(ori_ori_n559_));
  NO2        o0531(.A(ori_ori_n559_), .B(ori_ori_n78_), .Y(ori_ori_n560_));
  NA3        o0532(.A(ori_ori_n501_), .B(ori_ori_n307_), .C(ori_ori_n45_), .Y(ori_ori_n561_));
  NOi32      o0533(.An(e), .Bn(c), .C(f), .Y(ori_ori_n562_));
  INV        o0534(.A(ori_ori_n198_), .Y(ori_ori_n563_));
  NA2        o0535(.A(ori_ori_n562_), .B(ori_ori_n164_), .Y(ori_ori_n564_));
  NA3        o0536(.A(ori_ori_n564_), .B(ori_ori_n561_), .C(ori_ori_n167_), .Y(ori_ori_n565_));
  AOI210     o0537(.A0(ori_ori_n486_), .A1(ori_ori_n364_), .B0(ori_ori_n276_), .Y(ori_ori_n566_));
  NA2        o0538(.A(ori_ori_n566_), .B(ori_ori_n249_), .Y(ori_ori_n567_));
  NOi21      o0539(.An(j), .B(l), .Y(ori_ori_n568_));
  NAi21      o0540(.An(k), .B(h), .Y(ori_ori_n569_));
  NO2        o0541(.A(ori_ori_n569_), .B(ori_ori_n247_), .Y(ori_ori_n570_));
  NA2        o0542(.A(ori_ori_n570_), .B(ori_ori_n568_), .Y(ori_ori_n571_));
  OR2        o0543(.A(ori_ori_n571_), .B(ori_ori_n537_), .Y(ori_ori_n572_));
  NOi31      o0544(.An(m), .B(n), .C(k), .Y(ori_ori_n573_));
  NA2        o0545(.A(ori_ori_n568_), .B(ori_ori_n573_), .Y(ori_ori_n574_));
  AOI210     o0546(.A0(ori_ori_n364_), .A1(ori_ori_n338_), .B0(ori_ori_n276_), .Y(ori_ori_n575_));
  NAi21      o0547(.An(ori_ori_n574_), .B(ori_ori_n575_), .Y(ori_ori_n576_));
  NO2        o0548(.A(ori_ori_n260_), .B(ori_ori_n48_), .Y(ori_ori_n577_));
  NA2        o0549(.A(ori_ori_n577_), .B(ori_ori_n519_), .Y(ori_ori_n578_));
  NA4        o0550(.A(ori_ori_n578_), .B(ori_ori_n576_), .C(ori_ori_n572_), .D(ori_ori_n567_), .Y(ori_ori_n579_));
  NA2        o0551(.A(ori_ori_n99_), .B(ori_ori_n36_), .Y(ori_ori_n580_));
  INV        o0552(.A(ori_ori_n327_), .Y(ori_ori_n581_));
  NO2        o0553(.A(ori_ori_n581_), .B(n), .Y(ori_ori_n582_));
  NO2        o0554(.A(ori_ori_n480_), .B(ori_ori_n165_), .Y(ori_ori_n583_));
  NA3        o0555(.A(ori_ori_n502_), .B(ori_ori_n255_), .C(ori_ori_n133_), .Y(ori_ori_n584_));
  NA2        o0556(.A(ori_ori_n455_), .B(ori_ori_n149_), .Y(ori_ori_n585_));
  NO3        o0557(.A(ori_ori_n361_), .B(ori_ori_n585_), .C(ori_ori_n78_), .Y(ori_ori_n586_));
  AOI210     o0558(.A0(ori_ori_n584_), .A1(ori_ori_n583_), .B0(ori_ori_n586_), .Y(ori_ori_n587_));
  AN3        o0559(.A(f), .B(d), .C(b), .Y(ori_ori_n588_));
  NA2        o0560(.A(ori_ori_n119_), .B(n), .Y(ori_ori_n589_));
  NA3        o0561(.A(ori_ori_n455_), .B(ori_ori_n149_), .C(ori_ori_n201_), .Y(ori_ori_n590_));
  AOI210     o0562(.A0(ori_ori_n589_), .A1(ori_ori_n220_), .B0(ori_ori_n590_), .Y(ori_ori_n591_));
  NAi31      o0563(.An(m), .B(n), .C(k), .Y(ori_ori_n592_));
  OR2        o0564(.A(ori_ori_n122_), .B(ori_ori_n59_), .Y(ori_ori_n593_));
  OAI210     o0565(.A0(ori_ori_n593_), .A1(ori_ori_n592_), .B0(ori_ori_n236_), .Y(ori_ori_n594_));
  OAI210     o0566(.A0(ori_ori_n594_), .A1(ori_ori_n591_), .B0(j), .Y(ori_ori_n595_));
  NA2        o0567(.A(ori_ori_n595_), .B(ori_ori_n587_), .Y(ori_ori_n596_));
  NO4        o0568(.A(ori_ori_n596_), .B(ori_ori_n579_), .C(ori_ori_n565_), .D(ori_ori_n560_), .Y(ori_ori_n597_));
  NA2        o0569(.A(ori_ori_n348_), .B(ori_ori_n152_), .Y(ori_ori_n598_));
  NAi31      o0570(.An(g), .B(h), .C(f), .Y(ori_ori_n599_));
  OR3        o0571(.A(ori_ori_n599_), .B(ori_ori_n260_), .C(n), .Y(ori_ori_n600_));
  OA210      o0572(.A0(ori_ori_n482_), .A1(n), .B0(ori_ori_n535_), .Y(ori_ori_n601_));
  NA3        o0573(.A(ori_ori_n382_), .B(ori_ori_n110_), .C(ori_ori_n75_), .Y(ori_ori_n602_));
  OAI210     o0574(.A0(ori_ori_n601_), .A1(ori_ori_n82_), .B0(ori_ori_n602_), .Y(ori_ori_n603_));
  NOi21      o0575(.An(ori_ori_n600_), .B(ori_ori_n603_), .Y(ori_ori_n604_));
  AOI210     o0576(.A0(ori_ori_n604_), .A1(ori_ori_n598_), .B0(ori_ori_n476_), .Y(ori_ori_n605_));
  OR2        o0577(.A(ori_ori_n66_), .B(ori_ori_n67_), .Y(ori_ori_n606_));
  NA2        o0578(.A(ori_ori_n543_), .B(ori_ori_n309_), .Y(ori_ori_n607_));
  OA220      o0579(.A0(ori_ori_n574_), .A1(ori_ori_n607_), .B0(ori_ori_n571_), .B1(ori_ori_n606_), .Y(ori_ori_n608_));
  NA3        o0580(.A(ori_ori_n473_), .B(ori_ori_n90_), .C(g), .Y(ori_ori_n609_));
  AN2        o0581(.A(h), .B(f), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n610_), .B(ori_ori_n37_), .Y(ori_ori_n611_));
  NA2        o0583(.A(ori_ori_n90_), .B(ori_ori_n45_), .Y(ori_ori_n612_));
  OAI220     o0584(.A0(ori_ori_n612_), .A1(ori_ori_n303_), .B0(ori_ori_n611_), .B1(ori_ori_n417_), .Y(ori_ori_n613_));
  AOI210     o0585(.A0(ori_ori_n516_), .A1(ori_ori_n385_), .B0(ori_ori_n48_), .Y(ori_ori_n614_));
  INV        o0586(.A(ori_ori_n613_), .Y(ori_ori_n615_));
  NA3        o0587(.A(ori_ori_n615_), .B(ori_ori_n609_), .C(ori_ori_n608_), .Y(ori_ori_n616_));
  NA2        o0588(.A(ori_ori_n121_), .B(ori_ori_n48_), .Y(ori_ori_n617_));
  AOI220     o0589(.A0(ori_ori_n617_), .A1(ori_ori_n479_), .B0(ori_ori_n327_), .B1(ori_ori_n103_), .Y(ori_ori_n618_));
  OA220      o0590(.A0(ori_ori_n618_), .A1(ori_ori_n499_), .B0(ori_ori_n325_), .B1(ori_ori_n101_), .Y(ori_ori_n619_));
  INV        o0591(.A(ori_ori_n619_), .Y(ori_ori_n620_));
  NO3        o0592(.A(ori_ori_n371_), .B(ori_ori_n178_), .C(ori_ori_n177_), .Y(ori_ori_n621_));
  NA2        o0593(.A(ori_ori_n621_), .B(ori_ori_n218_), .Y(ori_ori_n622_));
  NA3        o0594(.A(ori_ori_n622_), .B(ori_ori_n239_), .C(j), .Y(ori_ori_n623_));
  NO3        o0595(.A(ori_ori_n412_), .B(ori_ori_n162_), .C(i), .Y(ori_ori_n624_));
  NA2        o0596(.A(ori_ori_n416_), .B(ori_ori_n75_), .Y(ori_ori_n625_));
  NA2        o0597(.A(ori_ori_n623_), .B(ori_ori_n369_), .Y(ori_ori_n626_));
  NO4        o0598(.A(ori_ori_n626_), .B(ori_ori_n620_), .C(ori_ori_n616_), .D(ori_ori_n605_), .Y(ori_ori_n627_));
  NA4        o0599(.A(ori_ori_n627_), .B(ori_ori_n597_), .C(ori_ori_n554_), .D(ori_ori_n530_), .Y(ori08));
  NO2        o0600(.A(k), .B(h), .Y(ori_ori_n629_));
  AO210      o0601(.A0(ori_ori_n237_), .A1(ori_ori_n404_), .B0(ori_ori_n629_), .Y(ori_ori_n630_));
  NO2        o0602(.A(ori_ori_n630_), .B(ori_ori_n274_), .Y(ori_ori_n631_));
  NA2        o0603(.A(ori_ori_n562_), .B(ori_ori_n75_), .Y(ori_ori_n632_));
  INV        o0604(.A(ori_ori_n632_), .Y(ori_ori_n633_));
  NA2        o0605(.A(ori_ori_n633_), .B(ori_ori_n631_), .Y(ori_ori_n634_));
  NA2        o0606(.A(ori_ori_n75_), .B(ori_ori_n100_), .Y(ori_ori_n635_));
  NO2        o0607(.A(ori_ori_n635_), .B(ori_ori_n56_), .Y(ori_ori_n636_));
  NO4        o0608(.A(ori_ori_n345_), .B(ori_ori_n102_), .C(j), .D(ori_ori_n201_), .Y(ori_ori_n637_));
  NA2        o0609(.A(ori_ori_n526_), .B(ori_ori_n220_), .Y(ori_ori_n638_));
  AOI220     o0610(.A0(ori_ori_n638_), .A1(ori_ori_n314_), .B0(ori_ori_n637_), .B1(ori_ori_n636_), .Y(ori_ori_n639_));
  AOI210     o0611(.A0(ori_ori_n526_), .A1(ori_ori_n145_), .B0(ori_ori_n75_), .Y(ori_ori_n640_));
  NA4        o0612(.A(ori_ori_n203_), .B(ori_ori_n128_), .C(ori_ori_n44_), .D(h), .Y(ori_ori_n641_));
  AN2        o0613(.A(l), .B(k), .Y(ori_ori_n642_));
  NA3        o0614(.A(ori_ori_n642_), .B(ori_ori_n99_), .C(ori_ori_n67_), .Y(ori_ori_n643_));
  OAI210     o0615(.A0(ori_ori_n641_), .A1(g), .B0(ori_ori_n643_), .Y(ori_ori_n644_));
  NA2        o0616(.A(ori_ori_n644_), .B(ori_ori_n640_), .Y(ori_ori_n645_));
  NA4        o0617(.A(ori_ori_n645_), .B(ori_ori_n639_), .C(ori_ori_n634_), .D(ori_ori_n316_), .Y(ori_ori_n646_));
  AN2        o0618(.A(ori_ori_n483_), .B(ori_ori_n87_), .Y(ori_ori_n647_));
  NO4        o0619(.A(ori_ori_n162_), .B(ori_ori_n359_), .C(ori_ori_n102_), .D(g), .Y(ori_ori_n648_));
  AOI210     o0620(.A0(ori_ori_n648_), .A1(ori_ori_n638_), .B0(ori_ori_n468_), .Y(ori_ori_n649_));
  NO2        o0621(.A(ori_ori_n38_), .B(ori_ori_n200_), .Y(ori_ori_n650_));
  AOI220     o0622(.A0(ori_ori_n563_), .A1(ori_ori_n313_), .B0(ori_ori_n650_), .B1(ori_ori_n513_), .Y(ori_ori_n651_));
  NAi31      o0623(.An(ori_ori_n647_), .B(ori_ori_n651_), .C(ori_ori_n649_), .Y(ori_ori_n652_));
  OAI210     o0624(.A0(ori_ori_n502_), .A1(ori_ori_n46_), .B0(ori_ori_n593_), .Y(ori_ori_n653_));
  NO2        o0625(.A(ori_ori_n435_), .B(ori_ori_n121_), .Y(ori_ori_n654_));
  NA2        o0626(.A(ori_ori_n654_), .B(ori_ori_n653_), .Y(ori_ori_n655_));
  NO3        o0627(.A(ori_ori_n292_), .B(ori_ori_n120_), .C(ori_ori_n40_), .Y(ori_ori_n656_));
  NAi21      o0628(.An(ori_ori_n656_), .B(ori_ori_n643_), .Y(ori_ori_n657_));
  NA2        o0629(.A(ori_ori_n630_), .B(ori_ori_n123_), .Y(ori_ori_n658_));
  AOI220     o0630(.A0(ori_ori_n658_), .A1(ori_ori_n370_), .B0(ori_ori_n657_), .B1(ori_ori_n70_), .Y(ori_ori_n659_));
  NA2        o0631(.A(ori_ori_n655_), .B(ori_ori_n659_), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n327_), .B(ori_ori_n42_), .Y(ori_ori_n661_));
  NA3        o0633(.A(ori_ori_n622_), .B(ori_ori_n304_), .C(ori_ori_n351_), .Y(ori_ori_n662_));
  NA3        o0634(.A(m), .B(l), .C(k), .Y(ori_ori_n663_));
  AOI210     o0635(.A0(ori_ori_n602_), .A1(ori_ori_n600_), .B0(ori_ori_n663_), .Y(ori_ori_n664_));
  INV        o0636(.A(ori_ori_n664_), .Y(ori_ori_n665_));
  NA3        o0637(.A(ori_ori_n665_), .B(ori_ori_n662_), .C(ori_ori_n661_), .Y(ori_ori_n666_));
  NO4        o0638(.A(ori_ori_n666_), .B(ori_ori_n660_), .C(ori_ori_n652_), .D(ori_ori_n646_), .Y(ori_ori_n667_));
  INV        o0639(.A(ori_ori_n450_), .Y(ori_ori_n668_));
  NA2        o0640(.A(ori_ori_n668_), .B(ori_ori_n236_), .Y(ori_ori_n669_));
  NA2        o0641(.A(ori_ori_n642_), .B(ori_ori_n67_), .Y(ori_ori_n670_));
  NO4        o0642(.A(ori_ori_n621_), .B(ori_ori_n162_), .C(n), .D(i), .Y(ori_ori_n671_));
  NOi21      o0643(.An(h), .B(j), .Y(ori_ori_n672_));
  NA2        o0644(.A(ori_ori_n672_), .B(f), .Y(ori_ori_n673_));
  NO2        o0645(.A(ori_ori_n671_), .B(ori_ori_n624_), .Y(ori_ori_n674_));
  NO2        o0646(.A(ori_ori_n674_), .B(ori_ori_n670_), .Y(ori_ori_n675_));
  AOI210     o0647(.A0(ori_ori_n669_), .A1(l), .B0(ori_ori_n675_), .Y(ori_ori_n676_));
  NO2        o0648(.A(j), .B(i), .Y(ori_ori_n677_));
  NA3        o0649(.A(ori_ori_n677_), .B(ori_ori_n74_), .C(l), .Y(ori_ori_n678_));
  NA2        o0650(.A(ori_ori_n677_), .B(ori_ori_n33_), .Y(ori_ori_n679_));
  OR2        o0651(.A(ori_ori_n678_), .B(ori_ori_n537_), .Y(ori_ori_n680_));
  NO3        o0652(.A(ori_ori_n140_), .B(ori_ori_n48_), .C(ori_ori_n100_), .Y(ori_ori_n681_));
  NO3        o0653(.A(ori_ori_n491_), .B(ori_ori_n138_), .C(ori_ori_n67_), .Y(ori_ori_n682_));
  NO3        o0654(.A(ori_ori_n435_), .B(ori_ori_n396_), .C(j), .Y(ori_ori_n683_));
  AOI210     o0655(.A0(ori_ori_n479_), .A1(n), .B0(ori_ori_n501_), .Y(ori_ori_n684_));
  NA2        o0656(.A(ori_ori_n684_), .B(ori_ori_n504_), .Y(ori_ori_n685_));
  NO3        o0657(.A(ori_ori_n162_), .B(ori_ori_n359_), .C(ori_ori_n102_), .Y(ori_ori_n686_));
  AOI220     o0658(.A0(ori_ori_n686_), .A1(ori_ori_n233_), .B0(ori_ori_n557_), .B1(ori_ori_n284_), .Y(ori_ori_n687_));
  NAi31      o0659(.An(ori_ori_n550_), .B(ori_ori_n84_), .C(ori_ori_n75_), .Y(ori_ori_n688_));
  NA2        o0660(.A(ori_ori_n688_), .B(ori_ori_n687_), .Y(ori_ori_n689_));
  NA2        o0661(.A(ori_ori_n656_), .B(ori_ori_n640_), .Y(ori_ori_n690_));
  NO2        o0662(.A(ori_ori_n663_), .B(ori_ori_n82_), .Y(ori_ori_n691_));
  NO2        o0663(.A(ori_ori_n538_), .B(ori_ori_n106_), .Y(ori_ori_n692_));
  OAI210     o0664(.A0(ori_ori_n692_), .A1(ori_ori_n683_), .B0(ori_ori_n614_), .Y(ori_ori_n693_));
  NA2        o0665(.A(ori_ori_n693_), .B(ori_ori_n690_), .Y(ori_ori_n694_));
  OR2        o0666(.A(ori_ori_n694_), .B(ori_ori_n689_), .Y(ori_ori_n695_));
  NA3        o0667(.A(ori_ori_n684_), .B(ori_ori_n504_), .C(ori_ori_n503_), .Y(ori_ori_n696_));
  NA4        o0668(.A(ori_ori_n696_), .B(ori_ori_n203_), .C(ori_ori_n404_), .D(ori_ori_n34_), .Y(ori_ori_n697_));
  NO4        o0669(.A(ori_ori_n435_), .B(ori_ori_n392_), .C(j), .D(f), .Y(ori_ori_n698_));
  OAI220     o0670(.A0(ori_ori_n641_), .A1(ori_ori_n632_), .B0(ori_ori_n303_), .B1(ori_ori_n38_), .Y(ori_ori_n699_));
  AOI210     o0671(.A0(ori_ori_n698_), .A1(ori_ori_n243_), .B0(ori_ori_n699_), .Y(ori_ori_n700_));
  NA3        o0672(.A(ori_ori_n494_), .B(ori_ori_n271_), .C(h), .Y(ori_ori_n701_));
  OAI220     o0673(.A0(ori_ori_n701_), .A1(ori_ori_n547_), .B0(ori_ori_n678_), .B1(ori_ori_n606_), .Y(ori_ori_n702_));
  INV        o0674(.A(ori_ori_n702_), .Y(ori_ori_n703_));
  NA3        o0675(.A(ori_ori_n703_), .B(ori_ori_n700_), .C(ori_ori_n697_), .Y(ori_ori_n704_));
  OR2        o0676(.A(ori_ori_n691_), .B(ori_ori_n87_), .Y(ori_ori_n705_));
  AOI220     o0677(.A0(ori_ori_n705_), .A1(ori_ori_n225_), .B0(ori_ori_n683_), .B1(ori_ori_n577_), .Y(ori_ori_n706_));
  NO2        o0678(.A(ori_ori_n601_), .B(ori_ori_n67_), .Y(ori_ori_n707_));
  NA2        o0679(.A(ori_ori_n698_), .B(ori_ori_n707_), .Y(ori_ori_n708_));
  NA3        o0680(.A(ori_ori_n235_), .B(ori_ori_n58_), .C(b), .Y(ori_ori_n709_));
  AOI220     o0681(.A0(ori_ori_n546_), .A1(ori_ori_n29_), .B0(ori_ori_n416_), .B1(ori_ori_n75_), .Y(ori_ori_n710_));
  NA2        o0682(.A(ori_ori_n708_), .B(ori_ori_n706_), .Y(ori_ori_n711_));
  NOi41      o0683(.An(ori_ori_n680_), .B(ori_ori_n711_), .C(ori_ori_n704_), .D(ori_ori_n695_), .Y(ori_ori_n712_));
  NO3        o0684(.A(ori_ori_n308_), .B(ori_ori_n276_), .C(ori_ori_n102_), .Y(ori_ori_n713_));
  NA2        o0685(.A(ori_ori_n713_), .B(ori_ori_n685_), .Y(ori_ori_n714_));
  NA2        o0686(.A(ori_ori_n714_), .B(ori_ori_n372_), .Y(ori_ori_n715_));
  OR2        o0687(.A(ori_ori_n599_), .B(ori_ori_n83_), .Y(ori_ori_n716_));
  NOi31      o0688(.An(b), .B(d), .C(a), .Y(ori_ori_n717_));
  NO2        o0689(.A(ori_ori_n717_), .B(ori_ori_n544_), .Y(ori_ori_n718_));
  NO2        o0690(.A(ori_ori_n718_), .B(n), .Y(ori_ori_n719_));
  NOi21      o0691(.An(ori_ori_n710_), .B(ori_ori_n719_), .Y(ori_ori_n720_));
  OAI220     o0692(.A0(ori_ori_n720_), .A1(ori_ori_n716_), .B0(ori_ori_n701_), .B1(ori_ori_n545_), .Y(ori_ori_n721_));
  NO2        o0693(.A(ori_ori_n502_), .B(ori_ori_n75_), .Y(ori_ori_n722_));
  NO2        o0694(.A(ori_ori_n300_), .B(ori_ori_n106_), .Y(ori_ori_n723_));
  NOi21      o0695(.An(ori_ori_n723_), .B(ori_ori_n150_), .Y(ori_ori_n724_));
  AOI210     o0696(.A0(ori_ori_n713_), .A1(ori_ori_n722_), .B0(ori_ori_n724_), .Y(ori_ori_n725_));
  INV        o0697(.A(ori_ori_n725_), .Y(ori_ori_n726_));
  NO2        o0698(.A(ori_ori_n621_), .B(n), .Y(ori_ori_n727_));
  NA2        o0699(.A(ori_ori_n727_), .B(ori_ori_n631_), .Y(ori_ori_n728_));
  NO2        o0700(.A(ori_ori_n298_), .B(ori_ori_n224_), .Y(ori_ori_n729_));
  OAI210     o0701(.A0(ori_ori_n87_), .A1(ori_ori_n84_), .B0(ori_ori_n729_), .Y(ori_ori_n730_));
  INV        o0702(.A(ori_ori_n730_), .Y(ori_ori_n731_));
  OAI210     o0703(.A0(ori_ori_n540_), .A1(ori_ori_n539_), .B0(ori_ori_n328_), .Y(ori_ori_n732_));
  NAi31      o0704(.An(ori_ori_n731_), .B(ori_ori_n732_), .C(ori_ori_n728_), .Y(ori_ori_n733_));
  NO4        o0705(.A(ori_ori_n733_), .B(ori_ori_n726_), .C(ori_ori_n721_), .D(ori_ori_n715_), .Y(ori_ori_n734_));
  NA4        o0706(.A(ori_ori_n734_), .B(ori_ori_n712_), .C(ori_ori_n676_), .D(ori_ori_n667_), .Y(ori09));
  INV        o0707(.A(ori_ori_n111_), .Y(ori_ori_n736_));
  NA2        o0708(.A(f), .B(e), .Y(ori_ori_n737_));
  NO2        o0709(.A(ori_ori_n213_), .B(ori_ori_n102_), .Y(ori_ori_n738_));
  NA4        o0710(.A(ori_ori_n286_), .B(ori_ori_n423_), .C(ori_ori_n245_), .D(ori_ori_n108_), .Y(ori_ori_n739_));
  AOI210     o0711(.A0(ori_ori_n739_), .A1(g), .B0(ori_ori_n420_), .Y(ori_ori_n740_));
  NO2        o0712(.A(ori_ori_n740_), .B(ori_ori_n737_), .Y(ori_ori_n741_));
  NA2        o0713(.A(ori_ori_n398_), .B(e), .Y(ori_ori_n742_));
  NO2        o0714(.A(ori_ori_n742_), .B(ori_ori_n459_), .Y(ori_ori_n743_));
  AOI210     o0715(.A0(ori_ori_n741_), .A1(ori_ori_n736_), .B0(ori_ori_n743_), .Y(ori_ori_n744_));
  NO2        o0716(.A(ori_ori_n190_), .B(ori_ori_n200_), .Y(ori_ori_n745_));
  NA3        o0717(.A(m), .B(l), .C(i), .Y(ori_ori_n746_));
  NA4        o0718(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .D(f), .Y(ori_ori_n747_));
  INV        o0719(.A(ori_ori_n747_), .Y(ori_ori_n748_));
  OR2        o0720(.A(ori_ori_n748_), .B(ori_ori_n745_), .Y(ori_ori_n749_));
  NA2        o0721(.A(ori_ori_n716_), .B(ori_ori_n515_), .Y(ori_ori_n750_));
  OA210      o0722(.A0(ori_ori_n750_), .A1(ori_ori_n749_), .B0(ori_ori_n719_), .Y(ori_ori_n751_));
  INV        o0723(.A(ori_ori_n306_), .Y(ori_ori_n752_));
  NO2        o0724(.A(ori_ori_n116_), .B(ori_ori_n114_), .Y(ori_ori_n753_));
  INV        o0725(.A(ori_ori_n307_), .Y(ori_ori_n754_));
  AOI210     o0726(.A0(ori_ori_n754_), .A1(ori_ori_n753_), .B0(ori_ori_n542_), .Y(ori_ori_n755_));
  NA2        o0727(.A(ori_ori_n709_), .B(ori_ori_n303_), .Y(ori_ori_n756_));
  NA2        o0728(.A(ori_ori_n309_), .B(ori_ori_n310_), .Y(ori_ori_n757_));
  OAI210     o0729(.A0(ori_ori_n190_), .A1(ori_ori_n200_), .B0(ori_ori_n757_), .Y(ori_ori_n758_));
  AOI220     o0730(.A0(ori_ori_n758_), .A1(ori_ori_n756_), .B0(ori_ori_n755_), .B1(ori_ori_n752_), .Y(ori_ori_n759_));
  NA2        o0731(.A(ori_ori_n630_), .B(ori_ori_n123_), .Y(ori_ori_n760_));
  NA3        o0732(.A(ori_ori_n760_), .B(ori_ori_n176_), .C(ori_ori_n31_), .Y(ori_ori_n761_));
  NA3        o0733(.A(ori_ori_n761_), .B(ori_ori_n759_), .C(ori_ori_n564_), .Y(ori_ori_n762_));
  NO2        o0734(.A(ori_ori_n534_), .B(ori_ori_n446_), .Y(ori_ori_n763_));
  NA2        o0735(.A(ori_ori_n763_), .B(ori_ori_n176_), .Y(ori_ori_n764_));
  NOi21      o0736(.An(f), .B(d), .Y(ori_ori_n765_));
  NA2        o0737(.A(ori_ori_n765_), .B(m), .Y(ori_ori_n766_));
  NOi32      o0738(.An(g), .Bn(f), .C(d), .Y(ori_ori_n767_));
  NA4        o0739(.A(ori_ori_n767_), .B(ori_ori_n546_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n768_));
  NOi21      o0740(.An(ori_ori_n287_), .B(ori_ori_n768_), .Y(ori_ori_n769_));
  INV        o0741(.A(ori_ori_n769_), .Y(ori_ori_n770_));
  NA3        o0742(.A(ori_ori_n286_), .B(ori_ori_n245_), .C(ori_ori_n108_), .Y(ori_ori_n771_));
  AN2        o0743(.A(f), .B(d), .Y(ori_ori_n772_));
  NA3        o0744(.A(ori_ori_n428_), .B(ori_ori_n772_), .C(ori_ori_n75_), .Y(ori_ori_n773_));
  NO3        o0745(.A(ori_ori_n773_), .B(ori_ori_n67_), .C(ori_ori_n201_), .Y(ori_ori_n774_));
  NA2        o0746(.A(ori_ori_n771_), .B(ori_ori_n774_), .Y(ori_ori_n775_));
  NAi41      o0747(.An(ori_ori_n440_), .B(ori_ori_n775_), .C(ori_ori_n770_), .D(ori_ori_n764_), .Y(ori_ori_n776_));
  NA2        o0748(.A(ori_ori_n544_), .B(ori_ori_n75_), .Y(ori_ori_n777_));
  NO2        o0749(.A(ori_ori_n757_), .B(ori_ori_n777_), .Y(ori_ori_n778_));
  NO2        o0750(.A(ori_ori_n773_), .B(ori_ori_n387_), .Y(ori_ori_n779_));
  NOi41      o0751(.An(ori_ori_n211_), .B(ori_ori_n779_), .C(ori_ori_n778_), .D(ori_ori_n282_), .Y(ori_ori_n780_));
  NA2        o0752(.A(c), .B(ori_ori_n105_), .Y(ori_ori_n781_));
  NO2        o0753(.A(ori_ori_n781_), .B(ori_ori_n376_), .Y(ori_ori_n782_));
  NA3        o0754(.A(ori_ori_n782_), .B(ori_ori_n457_), .C(f), .Y(ori_ori_n783_));
  OR2        o0755(.A(ori_ori_n599_), .B(ori_ori_n488_), .Y(ori_ori_n784_));
  INV        o0756(.A(ori_ori_n784_), .Y(ori_ori_n785_));
  NA2        o0757(.A(ori_ori_n718_), .B(ori_ori_n101_), .Y(ori_ori_n786_));
  NA2        o0758(.A(ori_ori_n786_), .B(ori_ori_n785_), .Y(ori_ori_n787_));
  NA3        o0759(.A(ori_ori_n787_), .B(ori_ori_n783_), .C(ori_ori_n780_), .Y(ori_ori_n788_));
  NO4        o0760(.A(ori_ori_n788_), .B(ori_ori_n776_), .C(ori_ori_n762_), .D(ori_ori_n751_), .Y(ori_ori_n789_));
  NA2        o0761(.A(ori_ori_n102_), .B(j), .Y(ori_ori_n790_));
  NO2        o0762(.A(ori_ori_n303_), .B(ori_ori_n747_), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n123_), .B(ori_ori_n121_), .Y(ori_ori_n792_));
  NO2        o0764(.A(ori_ori_n218_), .B(ori_ori_n212_), .Y(ori_ori_n793_));
  AOI220     o0765(.A0(ori_ori_n793_), .A1(ori_ori_n215_), .B0(ori_ori_n281_), .B1(ori_ori_n792_), .Y(ori_ori_n794_));
  NO2        o0766(.A(ori_ori_n387_), .B(ori_ori_n737_), .Y(ori_ori_n795_));
  NA2        o0767(.A(ori_ori_n795_), .B(ori_ori_n509_), .Y(ori_ori_n796_));
  NA2        o0768(.A(ori_ori_n796_), .B(ori_ori_n794_), .Y(ori_ori_n797_));
  NA2        o0769(.A(e), .B(d), .Y(ori_ori_n798_));
  OAI220     o0770(.A0(ori_ori_n798_), .A1(c), .B0(ori_ori_n298_), .B1(d), .Y(ori_ori_n799_));
  NA3        o0771(.A(ori_ori_n799_), .B(ori_ori_n407_), .C(ori_ori_n455_), .Y(ori_ori_n800_));
  AOI210     o0772(.A0(ori_ori_n462_), .A1(ori_ori_n169_), .B0(ori_ori_n218_), .Y(ori_ori_n801_));
  AOI210     o0773(.A0(ori_ori_n563_), .A1(ori_ori_n313_), .B0(ori_ori_n801_), .Y(ori_ori_n802_));
  NA2        o0774(.A(ori_ori_n267_), .B(ori_ori_n154_), .Y(ori_ori_n803_));
  NA2        o0775(.A(ori_ori_n774_), .B(ori_ori_n803_), .Y(ori_ori_n804_));
  NA3        o0776(.A(ori_ori_n804_), .B(ori_ori_n802_), .C(ori_ori_n800_), .Y(ori_ori_n805_));
  NO3        o0777(.A(ori_ori_n805_), .B(ori_ori_n797_), .C(ori_ori_n791_), .Y(ori_ori_n806_));
  NA2        o0778(.A(ori_ori_n752_), .B(ori_ori_n31_), .Y(ori_ori_n807_));
  AO210      o0779(.A0(ori_ori_n807_), .A1(ori_ori_n632_), .B0(ori_ori_n204_), .Y(ori_ori_n808_));
  NA2        o0780(.A(ori_ori_n555_), .B(ori_ori_n562_), .Y(ori_ori_n809_));
  OAI210     o0781(.A0(ori_ori_n742_), .A1(ori_ori_n159_), .B0(ori_ori_n809_), .Y(ori_ori_n810_));
  OAI210     o0782(.A0(ori_ori_n738_), .A1(ori_ori_n803_), .B0(ori_ori_n767_), .Y(ori_ori_n811_));
  NO2        o0783(.A(ori_ori_n811_), .B(ori_ori_n547_), .Y(ori_ori_n812_));
  AOI210     o0784(.A0(ori_ori_n107_), .A1(ori_ori_n106_), .B0(ori_ori_n244_), .Y(ori_ori_n813_));
  NOi31      o0785(.An(ori_ori_n492_), .B(ori_ori_n766_), .C(ori_ori_n272_), .Y(ori_ori_n814_));
  NO3        o0786(.A(ori_ori_n814_), .B(ori_ori_n812_), .C(ori_ori_n810_), .Y(ori_ori_n815_));
  AO220      o0787(.A0(ori_ori_n407_), .A1(ori_ori_n672_), .B0(ori_ori_n164_), .B1(f), .Y(ori_ori_n816_));
  NA2        o0788(.A(ori_ori_n816_), .B(ori_ori_n799_), .Y(ori_ori_n817_));
  NO2        o0789(.A(ori_ori_n396_), .B(ori_ori_n64_), .Y(ori_ori_n818_));
  OAI210     o0790(.A0(ori_ori_n750_), .A1(ori_ori_n818_), .B0(ori_ori_n636_), .Y(ori_ori_n819_));
  AN4        o0791(.A(ori_ori_n819_), .B(ori_ori_n817_), .C(ori_ori_n815_), .D(ori_ori_n808_), .Y(ori_ori_n820_));
  NA4        o0792(.A(ori_ori_n820_), .B(ori_ori_n806_), .C(ori_ori_n789_), .D(ori_ori_n744_), .Y(ori12));
  NO4        o0793(.A(ori_ori_n397_), .B(ori_ori_n237_), .C(ori_ori_n531_), .D(ori_ori_n201_), .Y(ori_ori_n822_));
  NA2        o0794(.A(ori_ori_n492_), .B(ori_ori_n818_), .Y(ori_ori_n823_));
  NO2        o0795(.A(ori_ori_n405_), .B(ori_ori_n105_), .Y(ori_ori_n824_));
  NO2        o0796(.A(ori_ori_n753_), .B(ori_ori_n320_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n599_), .B(ori_ori_n345_), .Y(ori_ori_n826_));
  NA2        o0798(.A(ori_ori_n825_), .B(ori_ori_n824_), .Y(ori_ori_n827_));
  NA2        o0799(.A(ori_ori_n827_), .B(ori_ori_n823_), .Y(ori_ori_n828_));
  AOI210     o0800(.A0(ori_ori_n221_), .A1(ori_ori_n305_), .B0(ori_ori_n187_), .Y(ori_ori_n829_));
  OR2        o0801(.A(ori_ori_n829_), .B(ori_ori_n822_), .Y(ori_ori_n830_));
  NO2        o0802(.A(ori_ori_n357_), .B(ori_ori_n201_), .Y(ori_ori_n831_));
  OAI210     o0803(.A0(ori_ori_n831_), .A1(ori_ori_n830_), .B0(ori_ori_n371_), .Y(ori_ori_n832_));
  NO2        o0804(.A(ori_ori_n580_), .B(ori_ori_n247_), .Y(ori_ori_n833_));
  NO2        o0805(.A(ori_ori_n538_), .B(ori_ori_n746_), .Y(ori_ori_n834_));
  AOI220     o0806(.A0(ori_ori_n834_), .A1(ori_ori_n513_), .B0(ori_ori_n729_), .B1(ori_ori_n833_), .Y(ori_ori_n835_));
  NO2        o0807(.A(ori_ori_n140_), .B(ori_ori_n224_), .Y(ori_ori_n836_));
  NA3        o0808(.A(ori_ori_n836_), .B(ori_ori_n227_), .C(i), .Y(ori_ori_n837_));
  NA3        o0809(.A(ori_ori_n837_), .B(ori_ori_n835_), .C(ori_ori_n832_), .Y(ori_ori_n838_));
  OR2        o0810(.A(ori_ori_n299_), .B(ori_ori_n824_), .Y(ori_ori_n839_));
  NA2        o0811(.A(ori_ori_n839_), .B(ori_ori_n321_), .Y(ori_ori_n840_));
  NA4        o0812(.A(ori_ori_n398_), .B(ori_ori_n394_), .C(ori_ori_n170_), .D(g), .Y(ori_ori_n841_));
  NA2        o0813(.A(ori_ori_n841_), .B(ori_ori_n840_), .Y(ori_ori_n842_));
  NO3        o0814(.A(ori_ori_n604_), .B(ori_ori_n83_), .C(ori_ori_n44_), .Y(ori_ori_n843_));
  NO4        o0815(.A(ori_ori_n843_), .B(ori_ori_n842_), .C(ori_ori_n838_), .D(ori_ori_n828_), .Y(ori_ori_n844_));
  NO2        o0816(.A(ori_ori_n335_), .B(ori_ori_n334_), .Y(ori_ori_n845_));
  INV        o0817(.A(ori_ori_n66_), .Y(ori_ori_n846_));
  NA2        o0818(.A(ori_ori_n502_), .B(ori_ori_n133_), .Y(ori_ori_n847_));
  NOi21      o0819(.An(ori_ori_n34_), .B(ori_ori_n592_), .Y(ori_ori_n848_));
  AOI220     o0820(.A0(ori_ori_n848_), .A1(ori_ori_n847_), .B0(ori_ori_n846_), .B1(ori_ori_n845_), .Y(ori_ori_n849_));
  OAI210     o0821(.A0(ori_ori_n236_), .A1(ori_ori_n44_), .B0(ori_ori_n849_), .Y(ori_ori_n850_));
  INV        o0822(.A(ori_ori_n296_), .Y(ori_ori_n851_));
  NO2        o0823(.A(ori_ori_n48_), .B(ori_ori_n44_), .Y(ori_ori_n852_));
  NO2        o0824(.A(ori_ori_n453_), .B(ori_ori_n276_), .Y(ori_ori_n853_));
  INV        o0825(.A(ori_ori_n853_), .Y(ori_ori_n854_));
  NO2        o0826(.A(ori_ori_n854_), .B(ori_ori_n133_), .Y(ori_ori_n855_));
  INV        o0827(.A(ori_ori_n332_), .Y(ori_ori_n856_));
  NO4        o0828(.A(ori_ori_n856_), .B(ori_ori_n855_), .C(ori_ori_n851_), .D(ori_ori_n850_), .Y(ori_ori_n857_));
  NA2        o0829(.A(ori_ori_n313_), .B(g), .Y(ori_ori_n858_));
  NA2        o0830(.A(ori_ori_n152_), .B(i), .Y(ori_ori_n859_));
  NA2        o0831(.A(ori_ori_n45_), .B(i), .Y(ori_ori_n860_));
  OAI220     o0832(.A0(ori_ori_n860_), .A1(ori_ori_n186_), .B0(ori_ori_n859_), .B1(ori_ori_n83_), .Y(ori_ori_n861_));
  INV        o0833(.A(ori_ori_n861_), .Y(ori_ori_n862_));
  NO2        o0834(.A(ori_ori_n133_), .B(ori_ori_n75_), .Y(ori_ori_n863_));
  OR2        o0835(.A(ori_ori_n863_), .B(ori_ori_n501_), .Y(ori_ori_n864_));
  NA2        o0836(.A(ori_ori_n502_), .B(ori_ori_n349_), .Y(ori_ori_n865_));
  AOI210     o0837(.A0(ori_ori_n865_), .A1(n), .B0(ori_ori_n864_), .Y(ori_ori_n866_));
  OAI220     o0838(.A0(ori_ori_n866_), .A1(ori_ori_n858_), .B0(ori_ori_n862_), .B1(ori_ori_n303_), .Y(ori_ori_n867_));
  NO2        o0839(.A(ori_ori_n599_), .B(ori_ori_n446_), .Y(ori_ori_n868_));
  NA3        o0840(.A(ori_ori_n309_), .B(ori_ori_n568_), .C(i), .Y(ori_ori_n869_));
  OAI210     o0841(.A0(ori_ori_n396_), .A1(ori_ori_n286_), .B0(ori_ori_n869_), .Y(ori_ori_n870_));
  OAI220     o0842(.A0(ori_ori_n870_), .A1(ori_ori_n868_), .B0(ori_ori_n614_), .B1(ori_ori_n682_), .Y(ori_ori_n871_));
  NA2        o0843(.A(ori_ori_n549_), .B(ori_ori_n103_), .Y(ori_ori_n872_));
  OR3        o0844(.A(ori_ori_n286_), .B(ori_ori_n392_), .C(f), .Y(ori_ori_n873_));
  NA2        o0845(.A(ori_ori_n74_), .B(i), .Y(ori_ori_n874_));
  OR2        o0846(.A(ori_ori_n873_), .B(ori_ori_n537_), .Y(ori_ori_n875_));
  NO2        o0847(.A(ori_ori_n611_), .B(m), .Y(ori_ori_n876_));
  OAI210     o0848(.A0(ori_ori_n876_), .A1(ori_ori_n825_), .B0(ori_ori_n299_), .Y(ori_ori_n877_));
  NA2        o0849(.A(ori_ori_n625_), .B(ori_ori_n777_), .Y(ori_ori_n878_));
  INV        o0850(.A(ori_ori_n747_), .Y(ori_ori_n879_));
  NA2        o0851(.A(ori_ori_n209_), .B(ori_ori_n71_), .Y(ori_ori_n880_));
  NA2        o0852(.A(ori_ori_n880_), .B(ori_ori_n874_), .Y(ori_ori_n881_));
  AOI220     o0853(.A0(ori_ori_n881_), .A1(ori_ori_n243_), .B0(ori_ori_n879_), .B1(ori_ori_n878_), .Y(ori_ori_n882_));
  NA4        o0854(.A(ori_ori_n882_), .B(ori_ori_n877_), .C(ori_ori_n875_), .D(ori_ori_n871_), .Y(ori_ori_n883_));
  NO2        o0855(.A(ori_ori_n345_), .B(ori_ori_n82_), .Y(ori_ori_n884_));
  OAI210     o0856(.A0(ori_ori_n884_), .A1(ori_ori_n833_), .B0(ori_ori_n225_), .Y(ori_ori_n885_));
  NA2        o0857(.A(ori_ori_n603_), .B(ori_ori_n79_), .Y(ori_ori_n886_));
  NO2        o0858(.A(ori_ori_n411_), .B(ori_ori_n201_), .Y(ori_ori_n887_));
  AOI220     o0859(.A0(ori_ori_n887_), .A1(ori_ori_n350_), .B0(ori_ori_n839_), .B1(ori_ori_n205_), .Y(ori_ori_n888_));
  AOI220     o0860(.A0(ori_ori_n826_), .A1(ori_ori_n836_), .B0(ori_ori_n536_), .B1(ori_ori_n81_), .Y(ori_ori_n889_));
  NA4        o0861(.A(ori_ori_n889_), .B(ori_ori_n888_), .C(ori_ori_n886_), .D(ori_ori_n885_), .Y(ori_ori_n890_));
  OAI210     o0862(.A0(ori_ori_n879_), .A1(ori_ori_n834_), .B0(ori_ori_n490_), .Y(ori_ori_n891_));
  NA2        o0863(.A(ori_ori_n876_), .B(ori_ori_n824_), .Y(ori_ori_n892_));
  NO3        o0864(.A(ori_ori_n790_), .B(ori_ori_n48_), .C(ori_ori_n44_), .Y(ori_ori_n893_));
  AOI220     o0865(.A0(ori_ori_n893_), .A1(ori_ori_n566_), .B0(ori_ori_n583_), .B1(ori_ori_n479_), .Y(ori_ori_n894_));
  NA3        o0866(.A(ori_ori_n894_), .B(ori_ori_n892_), .C(ori_ori_n891_), .Y(ori_ori_n895_));
  NO4        o0867(.A(ori_ori_n895_), .B(ori_ori_n890_), .C(ori_ori_n883_), .D(ori_ori_n867_), .Y(ori_ori_n896_));
  NAi31      o0868(.An(ori_ori_n129_), .B(ori_ori_n383_), .C(n), .Y(ori_ori_n897_));
  NO2        o0869(.A(ori_ori_n114_), .B(ori_ori_n307_), .Y(ori_ori_n898_));
  NO2        o0870(.A(ori_ori_n898_), .B(ori_ori_n897_), .Y(ori_ori_n899_));
  NA2        o0871(.A(ori_ori_n218_), .B(ori_ori_n160_), .Y(ori_ori_n900_));
  NO3        o0872(.A(ori_ori_n284_), .B(ori_ori_n398_), .C(ori_ori_n164_), .Y(ori_ori_n901_));
  NOi31      o0873(.An(ori_ori_n900_), .B(ori_ori_n901_), .C(ori_ori_n201_), .Y(ori_ori_n902_));
  NAi21      o0874(.An(ori_ori_n502_), .B(ori_ori_n887_), .Y(ori_ori_n903_));
  NA2        o0875(.A(ori_ori_n432_), .B(g), .Y(ori_ori_n904_));
  NA2        o0876(.A(ori_ori_n904_), .B(ori_ori_n903_), .Y(ori_ori_n905_));
  OAI220     o0877(.A0(ori_ori_n897_), .A1(ori_ori_n221_), .B0(ori_ori_n869_), .B1(ori_ori_n545_), .Y(ori_ori_n906_));
  NO2        o0878(.A(ori_ori_n600_), .B(ori_ori_n345_), .Y(ori_ori_n907_));
  INV        o0879(.A(ori_ori_n561_), .Y(ori_ori_n908_));
  OAI210     o0880(.A0(ori_ori_n829_), .A1(ori_ori_n822_), .B0(ori_ori_n900_), .Y(ori_ori_n909_));
  NA3        o0881(.A(ori_ori_n865_), .B(ori_ori_n437_), .C(ori_ori_n45_), .Y(ori_ori_n910_));
  AOI210     o0882(.A0(ori_ori_n348_), .A1(ori_ori_n346_), .B0(ori_ori_n302_), .Y(ori_ori_n911_));
  NA4        o0883(.A(ori_ori_n911_), .B(ori_ori_n910_), .C(ori_ori_n909_), .D(ori_ori_n256_), .Y(ori_ori_n912_));
  OR4        o0884(.A(ori_ori_n912_), .B(ori_ori_n908_), .C(ori_ori_n907_), .D(ori_ori_n906_), .Y(ori_ori_n913_));
  NO4        o0885(.A(ori_ori_n913_), .B(ori_ori_n905_), .C(ori_ori_n902_), .D(ori_ori_n899_), .Y(ori_ori_n914_));
  NA4        o0886(.A(ori_ori_n914_), .B(ori_ori_n896_), .C(ori_ori_n857_), .D(ori_ori_n844_), .Y(ori13));
  AN2        o0887(.A(c), .B(b), .Y(ori_ori_n916_));
  NA3        o0888(.A(ori_ori_n235_), .B(ori_ori_n916_), .C(m), .Y(ori_ori_n917_));
  AN2        o0889(.A(d), .B(c), .Y(ori_ori_n918_));
  NA2        o0890(.A(ori_ori_n918_), .B(ori_ori_n105_), .Y(ori_ori_n919_));
  NAi32      o0891(.An(f), .Bn(e), .C(c), .Y(ori_ori_n920_));
  NO3        o0892(.A(m), .B(i), .C(h), .Y(ori_ori_n921_));
  NA3        o0893(.A(k), .B(j), .C(i), .Y(ori_ori_n922_));
  NO2        o0894(.A(f), .B(c), .Y(ori_ori_n923_));
  NOi21      o0895(.An(ori_ori_n923_), .B(ori_ori_n397_), .Y(ori_ori_n924_));
  AN3        o0896(.A(g), .B(f), .C(c), .Y(ori_ori_n925_));
  NA3        o0897(.A(l), .B(k), .C(j), .Y(ori_ori_n926_));
  NA2        o0898(.A(i), .B(h), .Y(ori_ori_n927_));
  NO3        o0899(.A(ori_ori_n927_), .B(ori_ori_n926_), .C(ori_ori_n121_), .Y(ori_ori_n928_));
  NO3        o0900(.A(ori_ori_n130_), .B(ori_ori_n266_), .C(ori_ori_n201_), .Y(ori_ori_n929_));
  NA3        o0901(.A(c), .B(b), .C(a), .Y(ori_ori_n930_));
  NO2        o0902(.A(ori_ori_n475_), .B(ori_ori_n542_), .Y(ori_ori_n931_));
  NA4        o0903(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(g), .D(ori_ori_n200_), .Y(ori_ori_n932_));
  NA4        o0904(.A(ori_ori_n523_), .B(m), .C(ori_ori_n102_), .D(ori_ori_n200_), .Y(ori_ori_n933_));
  NA3        o0905(.A(ori_ori_n933_), .B(ori_ori_n336_), .C(ori_ori_n932_), .Y(ori_ori_n934_));
  NO2        o0906(.A(ori_ori_n934_), .B(ori_ori_n931_), .Y(ori_ori_n935_));
  NOi41      o0907(.An(ori_ori_n716_), .B(ori_ori_n758_), .C(ori_ori_n748_), .D(ori_ori_n650_), .Y(ori_ori_n936_));
  OAI220     o0908(.A0(ori_ori_n936_), .A1(ori_ori_n625_), .B0(ori_ori_n935_), .B1(ori_ori_n535_), .Y(ori_ori_n937_));
  NOi31      o0909(.An(m), .B(n), .C(f), .Y(ori_ori_n938_));
  NA2        o0910(.A(ori_ori_n938_), .B(ori_ori_n50_), .Y(ori_ori_n939_));
  NA2        o0911(.A(ori_ori_n455_), .B(l), .Y(ori_ori_n940_));
  NOi31      o0912(.An(ori_ori_n767_), .B(ori_ori_n917_), .C(ori_ori_n940_), .Y(ori_ori_n941_));
  NO2        o0913(.A(ori_ori_n266_), .B(a), .Y(ori_ori_n942_));
  NO2        o0914(.A(ori_ori_n78_), .B(g), .Y(ori_ori_n943_));
  NO4        o0915(.A(ori_ori_n941_), .B(ori_ori_n937_), .C(ori_ori_n731_), .D(ori_ori_n512_), .Y(ori_ori_n944_));
  NA2        o0916(.A(c), .B(b), .Y(ori_ori_n945_));
  NO2        o0917(.A(ori_ori_n635_), .B(ori_ori_n945_), .Y(ori_ori_n946_));
  OAI210     o0918(.A0(ori_ori_n766_), .A1(ori_ori_n740_), .B0(ori_ori_n381_), .Y(ori_ori_n947_));
  NA2        o0919(.A(ori_ori_n947_), .B(ori_ori_n946_), .Y(ori_ori_n948_));
  NA3        o0920(.A(ori_ori_n386_), .B(ori_ori_n507_), .C(f), .Y(ori_ori_n949_));
  NA2        o0921(.A(ori_ori_n496_), .B(ori_ori_n942_), .Y(ori_ori_n950_));
  NA2        o0922(.A(ori_ori_n950_), .B(ori_ori_n949_), .Y(ori_ori_n951_));
  INV        o0923(.A(g), .Y(ori_ori_n952_));
  NAi21      o0924(.An(f), .B(d), .Y(ori_ori_n953_));
  NO2        o0925(.A(ori_ori_n953_), .B(ori_ori_n930_), .Y(ori_ori_n954_));
  INV        o0926(.A(ori_ori_n954_), .Y(ori_ori_n955_));
  AOI210     o0927(.A0(ori_ori_n952_), .A1(ori_ori_n272_), .B0(ori_ori_n955_), .Y(ori_ori_n956_));
  AOI210     o0928(.A0(ori_ori_n956_), .A1(ori_ori_n103_), .B0(ori_ori_n951_), .Y(ori_ori_n957_));
  NA2        o0929(.A(ori_ori_n420_), .B(ori_ori_n419_), .Y(ori_ori_n958_));
  NO2        o0930(.A(ori_ori_n171_), .B(ori_ori_n224_), .Y(ori_ori_n959_));
  NA2        o0931(.A(ori_ori_n959_), .B(m), .Y(ori_ori_n960_));
  NA3        o0932(.A(ori_ori_n813_), .B(ori_ori_n940_), .C(ori_ori_n423_), .Y(ori_ori_n961_));
  OAI210     o0933(.A0(ori_ori_n961_), .A1(ori_ori_n287_), .B0(ori_ori_n421_), .Y(ori_ori_n962_));
  AOI210     o0934(.A0(ori_ori_n962_), .A1(ori_ori_n958_), .B0(ori_ori_n960_), .Y(ori_ori_n963_));
  NA2        o0935(.A(ori_ori_n509_), .B(ori_ori_n378_), .Y(ori_ori_n964_));
  NA2        o0936(.A(ori_ori_n401_), .B(ori_ori_n954_), .Y(ori_ori_n965_));
  NO2        o0937(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n966_));
  NA2        o0938(.A(ori_ori_n959_), .B(ori_ori_n388_), .Y(ori_ori_n967_));
  NAi41      o0939(.An(ori_ori_n966_), .B(ori_ori_n967_), .C(ori_ori_n965_), .D(ori_ori_n964_), .Y(ori_ori_n968_));
  NO2        o0940(.A(ori_ori_n968_), .B(ori_ori_n963_), .Y(ori_ori_n969_));
  NA4        o0941(.A(ori_ori_n969_), .B(ori_ori_n957_), .C(ori_ori_n948_), .D(ori_ori_n944_), .Y(ori00));
  NO2        o0942(.A(ori_ori_n275_), .B(ori_ori_n259_), .Y(ori_ori_n971_));
  NO2        o0943(.A(ori_ori_n971_), .B(ori_ori_n526_), .Y(ori_ori_n972_));
  NA2        o0944(.A(ori_ori_n795_), .B(ori_ori_n836_), .Y(ori_ori_n973_));
  INV        o0945(.A(ori_ori_n973_), .Y(ori_ori_n974_));
  NA2        o0946(.A(ori_ori_n457_), .B(f), .Y(ori_ori_n975_));
  OAI210     o0947(.A0(ori_ori_n898_), .A1(ori_ori_n39_), .B0(ori_ori_n585_), .Y(ori_ori_n976_));
  NA3        o0948(.A(ori_ori_n976_), .B(ori_ori_n242_), .C(n), .Y(ori_ori_n977_));
  AOI210     o0949(.A0(ori_ori_n977_), .A1(ori_ori_n975_), .B0(ori_ori_n919_), .Y(ori_ori_n978_));
  NO3        o0950(.A(ori_ori_n978_), .B(ori_ori_n974_), .C(ori_ori_n972_), .Y(ori_ori_n979_));
  NA3        o0951(.A(d), .B(ori_ori_n55_), .C(b), .Y(ori_ori_n980_));
  INV        o0952(.A(ori_ori_n525_), .Y(ori_ori_n981_));
  NO3        o0953(.A(ori_ori_n981_), .B(ori_ori_n966_), .C(ori_ori_n814_), .Y(ori_ori_n982_));
  NO4        o0954(.A(ori_ori_n438_), .B(ori_ori_n322_), .C(ori_ori_n945_), .D(ori_ori_n58_), .Y(ori_ori_n983_));
  NA3        o0955(.A(ori_ori_n351_), .B(ori_ori_n208_), .C(g), .Y(ori_ori_n984_));
  OA220      o0956(.A0(ori_ori_n984_), .A1(ori_ori_n980_), .B0(ori_ori_n352_), .B1(ori_ori_n122_), .Y(ori_ori_n985_));
  NO2        o0957(.A(h), .B(g), .Y(ori_ori_n986_));
  NA4        o0958(.A(ori_ori_n447_), .B(ori_ori_n418_), .C(ori_ori_n986_), .D(ori_ori_n916_), .Y(ori_ori_n987_));
  OAI220     o0959(.A0(ori_ori_n475_), .A1(ori_ori_n542_), .B0(ori_ori_n83_), .B1(ori_ori_n82_), .Y(ori_ori_n988_));
  NA2        o0960(.A(ori_ori_n988_), .B(ori_ori_n483_), .Y(ori_ori_n989_));
  AOI220     o0961(.A0(ori_ori_n293_), .A1(ori_ori_n233_), .B0(ori_ori_n166_), .B1(ori_ori_n137_), .Y(ori_ori_n990_));
  NA4        o0962(.A(ori_ori_n990_), .B(ori_ori_n989_), .C(ori_ori_n987_), .D(ori_ori_n985_), .Y(ori_ori_n991_));
  NO3        o0963(.A(ori_ori_n991_), .B(ori_ori_n983_), .C(ori_ori_n251_), .Y(ori_ori_n992_));
  INV        o0964(.A(ori_ori_n297_), .Y(ori_ori_n993_));
  AOI210     o0965(.A0(ori_ori_n233_), .A1(ori_ori_n313_), .B0(ori_ori_n527_), .Y(ori_ori_n994_));
  NA3        o0966(.A(ori_ori_n994_), .B(ori_ori_n993_), .C(ori_ori_n143_), .Y(ori_ori_n995_));
  NO2        o0967(.A(ori_ori_n995_), .B(ori_ori_n466_), .Y(ori_ori_n996_));
  AN3        o0968(.A(ori_ori_n996_), .B(ori_ori_n992_), .C(ori_ori_n982_), .Y(ori_ori_n997_));
  NA2        o0969(.A(ori_ori_n483_), .B(ori_ori_n92_), .Y(ori_ori_n998_));
  NA2        o0970(.A(ori_ori_n998_), .B(ori_ori_n228_), .Y(ori_ori_n999_));
  NA2        o0971(.A(ori_ori_n934_), .B(ori_ori_n483_), .Y(ori_ori_n1000_));
  NA4        o0972(.A(ori_ori_n588_), .B(ori_ori_n192_), .C(ori_ori_n208_), .D(ori_ori_n152_), .Y(ori_ori_n1001_));
  NA2        o0973(.A(ori_ori_n1001_), .B(ori_ori_n1000_), .Y(ori_ori_n1002_));
  OAI210     o0974(.A0(ori_ori_n417_), .A1(ori_ori_n109_), .B0(ori_ori_n768_), .Y(ori_ori_n1003_));
  AOI220     o0975(.A0(ori_ori_n1003_), .A1(ori_ori_n961_), .B0(ori_ori_n509_), .B1(ori_ori_n378_), .Y(ori_ori_n1004_));
  NO2        o0976(.A(ori_ori_n204_), .B(ori_ori_n201_), .Y(ori_ori_n1005_));
  NA2        o0977(.A(n), .B(e), .Y(ori_ori_n1006_));
  NO2        o0978(.A(ori_ori_n1006_), .B(ori_ori_n135_), .Y(ori_ori_n1007_));
  AOI220     o0979(.A0(ori_ori_n1007_), .A1(ori_ori_n257_), .B0(ori_ori_n752_), .B1(ori_ori_n1005_), .Y(ori_ori_n1008_));
  OAI210     o0980(.A0(ori_ori_n323_), .A1(ori_ori_n288_), .B0(ori_ori_n403_), .Y(ori_ori_n1009_));
  NA3        o0981(.A(ori_ori_n1009_), .B(ori_ori_n1008_), .C(ori_ori_n1004_), .Y(ori_ori_n1010_));
  NA2        o0982(.A(ori_ori_n1007_), .B(ori_ori_n755_), .Y(ori_ori_n1011_));
  NA2        o0983(.A(ori_ori_n1011_), .B(ori_ori_n770_), .Y(ori_ori_n1012_));
  NO4        o0984(.A(ori_ori_n1012_), .B(ori_ori_n1010_), .C(ori_ori_n1002_), .D(ori_ori_n999_), .Y(ori_ori_n1013_));
  NA2        o0985(.A(ori_ori_n741_), .B(ori_ori_n681_), .Y(ori_ori_n1014_));
  NA4        o0986(.A(ori_ori_n1014_), .B(ori_ori_n1013_), .C(ori_ori_n997_), .D(ori_ori_n979_), .Y(ori01));
  INV        o0987(.A(ori_ori_n264_), .Y(ori_ori_n1016_));
  NA2        o0988(.A(ori_ori_n362_), .B(i), .Y(ori_ori_n1017_));
  NA2        o0989(.A(ori_ori_n1017_), .B(ori_ori_n1016_), .Y(ori_ori_n1018_));
  NA2        o0990(.A(ori_ori_n536_), .B(ori_ori_n81_), .Y(ori_ori_n1019_));
  NA2        o0991(.A(ori_ori_n502_), .B(ori_ori_n255_), .Y(ori_ori_n1020_));
  NA2        o0992(.A(ori_ori_n853_), .B(ori_ori_n1020_), .Y(ori_ori_n1021_));
  NA3        o0993(.A(ori_ori_n1021_), .B(ori_ori_n1019_), .C(ori_ori_n809_), .Y(ori_ori_n1022_));
  NA2        o0994(.A(ori_ori_n642_), .B(ori_ori_n88_), .Y(ori_ori_n1023_));
  NO2        o0995(.A(ori_ori_n1023_), .B(i), .Y(ori_ori_n1024_));
  OAI210     o0996(.A0(ori_ori_n701_), .A1(ori_ori_n545_), .B0(ori_ori_n1001_), .Y(ori_ori_n1025_));
  AOI210     o0997(.A0(ori_ori_n1024_), .A1(ori_ori_n577_), .B0(ori_ori_n1025_), .Y(ori_ori_n1026_));
  OR2        o0998(.A(ori_ori_n601_), .B(ori_ori_n336_), .Y(ori_ori_n1027_));
  NAi41      o0999(.An(ori_ori_n151_), .B(ori_ori_n1027_), .C(ori_ori_n1026_), .D(ori_ori_n794_), .Y(ori_ori_n1028_));
  NO2        o1000(.A(ori_ori_n613_), .B(ori_ori_n460_), .Y(ori_ori_n1029_));
  NA4        o1001(.A(ori_ori_n642_), .B(ori_ori_n88_), .C(ori_ori_n44_), .D(ori_ori_n200_), .Y(ori_ori_n1030_));
  OA220      o1002(.A0(ori_ori_n1030_), .A1(ori_ori_n606_), .B0(ori_ori_n181_), .B1(ori_ori_n179_), .Y(ori_ori_n1031_));
  NA3        o1003(.A(ori_ori_n1031_), .B(ori_ori_n1029_), .C(ori_ori_n125_), .Y(ori_ori_n1032_));
  NO4        o1004(.A(ori_ori_n1032_), .B(ori_ori_n1028_), .C(ori_ori_n1022_), .D(ori_ori_n1018_), .Y(ori_ori_n1033_));
  INV        o1005(.A(ori_ori_n984_), .Y(ori_ori_n1034_));
  OAI210     o1006(.A0(ori_ori_n1034_), .A1(ori_ori_n278_), .B0(ori_ori_n479_), .Y(ori_ori_n1035_));
  AOI210     o1007(.A0(ori_ori_n190_), .A1(ori_ori_n80_), .B0(ori_ori_n200_), .Y(ori_ori_n1036_));
  OAI210     o1008(.A0(ori_ori_n719_), .A1(ori_ori_n386_), .B0(ori_ori_n1036_), .Y(ori_ori_n1037_));
  NA2        o1009(.A(ori_ori_n1037_), .B(ori_ori_n1035_), .Y(ori_ori_n1038_));
  NA2        o1010(.A(ori_ori_n541_), .B(ori_ori_n107_), .Y(ori_ori_n1039_));
  INV        o1011(.A(ori_ori_n1039_), .Y(ori_ori_n1040_));
  NA2        o1012(.A(ori_ori_n1024_), .B(ori_ori_n614_), .Y(ori_ori_n1041_));
  NA2        o1013(.A(ori_ori_n1041_), .B(ori_ori_n703_), .Y(ori_ori_n1042_));
  NO3        o1014(.A(ori_ori_n1042_), .B(ori_ori_n1040_), .C(ori_ori_n1038_), .Y(ori_ori_n1043_));
  NA3        o1015(.A(ori_ori_n546_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1044_));
  NO2        o1016(.A(ori_ori_n1044_), .B(ori_ori_n190_), .Y(ori_ori_n1045_));
  AOI210     o1017(.A0(ori_ori_n454_), .A1(ori_ori_n57_), .B0(ori_ori_n1045_), .Y(ori_ori_n1046_));
  NO2        o1018(.A(ori_ori_n1030_), .B(ori_ori_n872_), .Y(ori_ori_n1047_));
  NO2        o1019(.A(ori_ori_n193_), .B(ori_ori_n101_), .Y(ori_ori_n1048_));
  NO2        o1020(.A(ori_ori_n1048_), .B(ori_ori_n1047_), .Y(ori_ori_n1049_));
  NA3        o1021(.A(ori_ori_n1049_), .B(ori_ori_n1046_), .C(ori_ori_n680_), .Y(ori_ori_n1050_));
  NO2        o1022(.A(ori_ori_n859_), .B(ori_ori_n220_), .Y(ori_ori_n1051_));
  NO2        o1023(.A(ori_ori_n860_), .B(ori_ori_n504_), .Y(ori_ori_n1052_));
  OAI210     o1024(.A0(ori_ori_n1052_), .A1(ori_ori_n1051_), .B0(ori_ori_n307_), .Y(ori_ori_n1053_));
  NA2        o1025(.A(ori_ori_n519_), .B(ori_ori_n517_), .Y(ori_ori_n1054_));
  NO3        o1026(.A(ori_ori_n73_), .B(ori_ori_n276_), .C(ori_ori_n44_), .Y(ori_ori_n1055_));
  NA2        o1027(.A(ori_ori_n1055_), .B(ori_ori_n501_), .Y(ori_ori_n1056_));
  NA3        o1028(.A(ori_ori_n1056_), .B(ori_ori_n1054_), .C(ori_ori_n608_), .Y(ori_ori_n1057_));
  OR2        o1029(.A(ori_ori_n984_), .B(ori_ori_n980_), .Y(ori_ori_n1058_));
  NO2        o1030(.A(ori_ori_n336_), .B(ori_ori_n66_), .Y(ori_ori_n1059_));
  INV        o1031(.A(ori_ori_n1059_), .Y(ori_ori_n1060_));
  NA2        o1032(.A(ori_ori_n1055_), .B(ori_ori_n722_), .Y(ori_ori_n1061_));
  NA4        o1033(.A(ori_ori_n1061_), .B(ori_ori_n1060_), .C(ori_ori_n1058_), .D(ori_ori_n354_), .Y(ori_ori_n1062_));
  NOi41      o1034(.An(ori_ori_n1053_), .B(ori_ori_n1062_), .C(ori_ori_n1057_), .D(ori_ori_n1050_), .Y(ori_ori_n1063_));
  INV        o1035(.A(ori_ori_n122_), .Y(ori_ori_n1064_));
  NO3        o1036(.A(ori_ori_n927_), .B(ori_ori_n165_), .C(ori_ori_n78_), .Y(ori_ori_n1065_));
  AOI220     o1037(.A0(ori_ori_n1065_), .A1(ori_ori_n1064_), .B0(ori_ori_n1055_), .B1(ori_ori_n863_), .Y(ori_ori_n1066_));
  INV        o1038(.A(ori_ori_n1066_), .Y(ori_ori_n1067_));
  NO2        o1039(.A(ori_ori_n557_), .B(ori_ori_n556_), .Y(ori_ori_n1068_));
  NO4        o1040(.A(ori_ori_n927_), .B(ori_ori_n1068_), .C(ori_ori_n163_), .D(ori_ori_n78_), .Y(ori_ori_n1069_));
  NO3        o1041(.A(ori_ori_n1069_), .B(ori_ori_n1067_), .C(ori_ori_n579_), .Y(ori_ori_n1070_));
  NA4        o1042(.A(ori_ori_n1070_), .B(ori_ori_n1063_), .C(ori_ori_n1043_), .D(ori_ori_n1033_), .Y(ori06));
  NO2        o1043(.A(ori_ori_n212_), .B(ori_ori_n94_), .Y(ori_ori_n1072_));
  OAI210     o1044(.A0(ori_ori_n1072_), .A1(ori_ori_n1065_), .B0(ori_ori_n350_), .Y(ori_ori_n1073_));
  NO3        o1045(.A(ori_ori_n543_), .B(ori_ori_n717_), .C(ori_ori_n544_), .Y(ori_ori_n1074_));
  OR2        o1046(.A(ori_ori_n1074_), .B(ori_ori_n784_), .Y(ori_ori_n1075_));
  NA3        o1047(.A(ori_ori_n1075_), .B(ori_ori_n1073_), .C(ori_ori_n1053_), .Y(ori_ori_n1076_));
  NO3        o1048(.A(ori_ori_n1076_), .B(ori_ori_n1057_), .C(ori_ori_n241_), .Y(ori_ori_n1077_));
  NO2        o1049(.A(ori_ori_n276_), .B(ori_ori_n44_), .Y(ori_ori_n1078_));
  AOI210     o1050(.A0(ori_ori_n1078_), .A1(ori_ori_n864_), .B0(ori_ori_n1051_), .Y(ori_ori_n1079_));
  NA2        o1051(.A(ori_ori_n1078_), .B(ori_ori_n505_), .Y(ori_ori_n1080_));
  AOI210     o1052(.A0(ori_ori_n1080_), .A1(ori_ori_n1079_), .B0(ori_ori_n305_), .Y(ori_ori_n1081_));
  OAI210     o1053(.A0(ori_ori_n80_), .A1(ori_ori_n39_), .B0(ori_ori_n612_), .Y(ori_ori_n1082_));
  NA2        o1054(.A(ori_ori_n1082_), .B(ori_ori_n582_), .Y(ori_ori_n1083_));
  NO2        o1055(.A(ori_ori_n462_), .B(ori_ori_n160_), .Y(ori_ori_n1084_));
  NOi21      o1056(.An(ori_ori_n124_), .B(ori_ori_n44_), .Y(ori_ori_n1085_));
  NO2        o1057(.A(ori_ori_n550_), .B(ori_ori_n939_), .Y(ori_ori_n1086_));
  NO3        o1058(.A(ori_ori_n1086_), .B(ori_ori_n1085_), .C(ori_ori_n1084_), .Y(ori_ori_n1087_));
  NA2        o1059(.A(ori_ori_n1087_), .B(ori_ori_n1083_), .Y(ori_ori_n1088_));
  NO2        o1060(.A(ori_ori_n673_), .B(ori_ori_n334_), .Y(ori_ori_n1089_));
  NO2        o1061(.A(ori_ori_n614_), .B(ori_ori_n577_), .Y(ori_ori_n1090_));
  NOi21      o1062(.An(ori_ori_n1089_), .B(ori_ori_n1090_), .Y(ori_ori_n1091_));
  AN2        o1063(.A(ori_ori_n848_), .B(ori_ori_n584_), .Y(ori_ori_n1092_));
  NO4        o1064(.A(ori_ori_n1092_), .B(ori_ori_n1091_), .C(ori_ori_n1088_), .D(ori_ori_n1081_), .Y(ori_ori_n1093_));
  NO3        o1065(.A(h), .B(ori_ori_n94_), .C(ori_ori_n266_), .Y(ori_ori_n1094_));
  OAI220     o1066(.A0(ori_ori_n632_), .A1(ori_ori_n234_), .B0(ori_ori_n459_), .B1(ori_ori_n462_), .Y(ori_ori_n1095_));
  INV        o1067(.A(k), .Y(ori_ori_n1096_));
  NO3        o1068(.A(ori_ori_n1096_), .B(ori_ori_n542_), .C(j), .Y(ori_ori_n1097_));
  NOi21      o1069(.An(ori_ori_n1097_), .B(ori_ori_n606_), .Y(ori_ori_n1098_));
  NO3        o1070(.A(ori_ori_n1098_), .B(ori_ori_n1095_), .C(ori_ori_n1094_), .Y(ori_ori_n1099_));
  NA4        o1071(.A(ori_ori_n710_), .B(ori_ori_n709_), .C(ori_ori_n395_), .D(ori_ori_n777_), .Y(ori_ori_n1100_));
  NAi31      o1072(.An(ori_ori_n673_), .B(ori_ori_n1100_), .C(ori_ori_n189_), .Y(ori_ori_n1101_));
  NA2        o1073(.A(ori_ori_n1101_), .B(ori_ori_n1099_), .Y(ori_ori_n1102_));
  AOI210     o1074(.A0(ori_ori_n519_), .A1(ori_ori_n403_), .B0(ori_ori_n340_), .Y(ori_ori_n1103_));
  NA2        o1075(.A(ori_ori_n1097_), .B(ori_ori_n707_), .Y(ori_ori_n1104_));
  NA2        o1076(.A(ori_ori_n1104_), .B(ori_ori_n1103_), .Y(ori_ori_n1105_));
  NO2        o1077(.A(ori_ori_n450_), .B(ori_ori_n432_), .Y(ori_ori_n1106_));
  NA2        o1078(.A(ori_ori_n1106_), .B(ori_ori_n1061_), .Y(ori_ori_n1107_));
  NAi21      o1079(.An(j), .B(i), .Y(ori_ori_n1108_));
  NO4        o1080(.A(ori_ori_n1068_), .B(ori_ori_n1108_), .C(ori_ori_n397_), .D(ori_ori_n222_), .Y(ori_ori_n1109_));
  NO4        o1081(.A(ori_ori_n1109_), .B(ori_ori_n1107_), .C(ori_ori_n1105_), .D(ori_ori_n1102_), .Y(ori_ori_n1110_));
  NA4        o1082(.A(ori_ori_n1110_), .B(ori_ori_n1093_), .C(ori_ori_n1077_), .D(ori_ori_n1070_), .Y(ori07));
  NAi32      o1083(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1112_));
  NO3        o1084(.A(ori_ori_n1112_), .B(g), .C(f), .Y(ori_ori_n1113_));
  OR2        o1085(.A(e), .B(d), .Y(ori_ori_n1114_));
  NOi31      o1086(.An(n), .B(m), .C(b), .Y(ori_ori_n1115_));
  NO3        o1087(.A(ori_ori_n121_), .B(ori_ori_n404_), .C(h), .Y(ori_ori_n1116_));
  NO3        o1088(.A(n), .B(m), .C(h), .Y(ori_ori_n1117_));
  NO2        o1089(.A(ori_ori_n920_), .B(ori_ori_n397_), .Y(ori_ori_n1118_));
  INV        o1090(.A(ori_ori_n1118_), .Y(ori_ori_n1119_));
  NO2        o1091(.A(ori_ori_n922_), .B(ori_ori_n283_), .Y(ori_ori_n1120_));
  NA2        o1092(.A(ori_ori_n489_), .B(ori_ori_n74_), .Y(ori_ori_n1121_));
  NA2        o1093(.A(ori_ori_n1121_), .B(ori_ori_n1119_), .Y(ori_ori_n1122_));
  NO2        o1094(.A(ori_ori_n1122_), .B(ori_ori_n1113_), .Y(ori_ori_n1123_));
  NO3        o1095(.A(e), .B(d), .C(c), .Y(ori_ori_n1124_));
  NO2        o1096(.A(ori_ori_n121_), .B(ori_ori_n201_), .Y(ori_ori_n1125_));
  NA2        o1097(.A(ori_ori_n1125_), .B(ori_ori_n1124_), .Y(ori_ori_n1126_));
  INV        o1098(.A(ori_ori_n1126_), .Y(ori_ori_n1127_));
  NA3        o1099(.A(ori_ori_n629_), .B(ori_ori_n617_), .C(ori_ori_n102_), .Y(ori_ori_n1128_));
  NO2        o1100(.A(ori_ori_n1128_), .B(ori_ori_n44_), .Y(ori_ori_n1129_));
  NO2        o1101(.A(l), .B(k), .Y(ori_ori_n1130_));
  NO3        o1102(.A(ori_ori_n397_), .B(d), .C(c), .Y(ori_ori_n1131_));
  NO2        o1103(.A(ori_ori_n1129_), .B(ori_ori_n1127_), .Y(ori_ori_n1132_));
  NO2        o1104(.A(g), .B(c), .Y(ori_ori_n1133_));
  NO2        o1105(.A(ori_ori_n405_), .B(a), .Y(ori_ori_n1134_));
  NA2        o1106(.A(ori_ori_n1134_), .B(ori_ori_n103_), .Y(ori_ori_n1135_));
  NO2        o1107(.A(ori_ori_n679_), .B(ori_ori_n175_), .Y(ori_ori_n1136_));
  NOi31      o1108(.An(m), .B(n), .C(b), .Y(ori_ori_n1137_));
  NOi31      o1109(.An(f), .B(d), .C(c), .Y(ori_ori_n1138_));
  NA2        o1110(.A(ori_ori_n1138_), .B(ori_ori_n1137_), .Y(ori_ori_n1139_));
  INV        o1111(.A(ori_ori_n1139_), .Y(ori_ori_n1140_));
  NO2        o1112(.A(ori_ori_n1140_), .B(ori_ori_n1136_), .Y(ori_ori_n1141_));
  NA2        o1113(.A(ori_ori_n925_), .B(ori_ori_n418_), .Y(ori_ori_n1142_));
  NO2        o1114(.A(ori_ori_n1142_), .B(ori_ori_n397_), .Y(ori_ori_n1143_));
  NO3        o1115(.A(ori_ori_n40_), .B(i), .C(h), .Y(ori_ori_n1144_));
  NO2        o1116(.A(ori_ori_n921_), .B(ori_ori_n1143_), .Y(ori_ori_n1145_));
  AN3        o1117(.A(ori_ori_n1145_), .B(ori_ori_n1141_), .C(ori_ori_n1135_), .Y(ori_ori_n1146_));
  NA2        o1118(.A(ori_ori_n1115_), .B(ori_ori_n347_), .Y(ori_ori_n1147_));
  INV        o1119(.A(ori_ori_n1147_), .Y(ori_ori_n1148_));
  INV        o1120(.A(ori_ori_n928_), .Y(ori_ori_n1149_));
  NAi21      o1121(.An(ori_ori_n1148_), .B(ori_ori_n1149_), .Y(ori_ori_n1150_));
  NO4        o1122(.A(ori_ori_n121_), .B(g), .C(f), .D(e), .Y(ori_ori_n1151_));
  NA2        o1123(.A(ori_ori_n1117_), .B(ori_ori_n1130_), .Y(ori_ori_n1152_));
  INV        o1124(.A(ori_ori_n1152_), .Y(ori_ori_n1153_));
  OR3        o1125(.A(ori_ori_n488_), .B(ori_ori_n487_), .C(ori_ori_n102_), .Y(ori_ori_n1154_));
  NA2        o1126(.A(ori_ori_n938_), .B(ori_ori_n376_), .Y(ori_ori_n1155_));
  NO2        o1127(.A(ori_ori_n1155_), .B(ori_ori_n394_), .Y(ori_ori_n1156_));
  AO210      o1128(.A0(ori_ori_n1156_), .A1(ori_ori_n105_), .B0(ori_ori_n1153_), .Y(ori_ori_n1157_));
  NO2        o1129(.A(ori_ori_n1157_), .B(ori_ori_n1150_), .Y(ori_ori_n1158_));
  NA4        o1130(.A(ori_ori_n1158_), .B(ori_ori_n1146_), .C(ori_ori_n1132_), .D(ori_ori_n1123_), .Y(ori_ori_n1159_));
  NO2        o1131(.A(ori_ori_n945_), .B(ori_ori_n100_), .Y(ori_ori_n1160_));
  NO2        o1132(.A(ori_ori_n359_), .B(j), .Y(ori_ori_n1161_));
  NA2        o1133(.A(ori_ori_n1144_), .B(ori_ori_n938_), .Y(ori_ori_n1162_));
  NA2        o1134(.A(ori_ori_n924_), .B(ori_ori_n139_), .Y(ori_ori_n1163_));
  NA2        o1135(.A(ori_ori_n1163_), .B(ori_ori_n1162_), .Y(ori_ori_n1164_));
  NA2        o1136(.A(ori_ori_n1161_), .B(ori_ori_n148_), .Y(ori_ori_n1165_));
  INV        o1137(.A(ori_ori_n1165_), .Y(ori_ori_n1166_));
  NO2        o1138(.A(ori_ori_n1166_), .B(ori_ori_n1164_), .Y(ori_ori_n1167_));
  INV        o1139(.A(ori_ori_n48_), .Y(ori_ori_n1168_));
  NA2        o1140(.A(ori_ori_n1168_), .B(ori_ori_n986_), .Y(ori_ori_n1169_));
  INV        o1141(.A(ori_ori_n1169_), .Y(ori_ori_n1170_));
  NO2        o1142(.A(ori_ori_n212_), .B(ori_ori_n165_), .Y(ori_ori_n1171_));
  NO2        o1143(.A(ori_ori_n1154_), .B(ori_ori_n320_), .Y(ori_ori_n1172_));
  NO3        o1144(.A(ori_ori_n1172_), .B(ori_ori_n1171_), .C(ori_ori_n1170_), .Y(ori_ori_n1173_));
  NO3        o1145(.A(ori_ori_n930_), .B(ori_ori_n1114_), .C(ori_ori_n48_), .Y(ori_ori_n1174_));
  NA3        o1146(.A(ori_ori_n1160_), .B(ori_ori_n418_), .C(f), .Y(ori_ori_n1175_));
  NO2        o1147(.A(ori_ori_n1210_), .B(ori_ori_n1175_), .Y(ori_ori_n1176_));
  NO2        o1148(.A(ori_ori_n1108_), .B(ori_ori_n163_), .Y(ori_ori_n1177_));
  NOi21      o1149(.An(d), .B(f), .Y(ori_ori_n1178_));
  NA2        o1150(.A(h), .B(ori_ori_n1177_), .Y(ori_ori_n1179_));
  INV        o1151(.A(ori_ori_n1179_), .Y(ori_ori_n1180_));
  NO2        o1152(.A(ori_ori_n1180_), .B(ori_ori_n1176_), .Y(ori_ori_n1181_));
  NA3        o1153(.A(ori_ori_n1181_), .B(ori_ori_n1173_), .C(ori_ori_n1167_), .Y(ori_ori_n1182_));
  NA2        o1154(.A(h), .B(ori_ori_n1120_), .Y(ori_ori_n1183_));
  OAI210     o1155(.A0(ori_ori_n1151_), .A1(ori_ori_n1115_), .B0(ori_ori_n781_), .Y(ori_ori_n1184_));
  NA2        o1156(.A(ori_ori_n1184_), .B(ori_ori_n1183_), .Y(ori_ori_n1185_));
  NA2        o1157(.A(ori_ori_n1133_), .B(ori_ori_n1178_), .Y(ori_ori_n1186_));
  NO2        o1158(.A(ori_ori_n1186_), .B(m), .Y(ori_ori_n1187_));
  NA2        o1159(.A(ori_ori_n929_), .B(ori_ori_n208_), .Y(ori_ori_n1188_));
  NO2        o1160(.A(ori_ori_n140_), .B(ori_ori_n170_), .Y(ori_ori_n1189_));
  OAI210     o1161(.A0(ori_ori_n1189_), .A1(ori_ori_n100_), .B0(ori_ori_n1137_), .Y(ori_ori_n1190_));
  NA2        o1162(.A(ori_ori_n1190_), .B(ori_ori_n1188_), .Y(ori_ori_n1191_));
  NO3        o1163(.A(ori_ori_n1191_), .B(ori_ori_n1187_), .C(ori_ori_n1185_), .Y(ori_ori_n1192_));
  NO2        o1164(.A(ori_ori_n1131_), .B(ori_ori_n1174_), .Y(ori_ori_n1193_));
  INV        o1165(.A(ori_ori_n943_), .Y(ori_ori_n1194_));
  OAI210     o1166(.A0(ori_ori_n1194_), .A1(ori_ori_n63_), .B0(ori_ori_n1193_), .Y(ori_ori_n1195_));
  OR2        o1167(.A(h), .B(ori_ori_n487_), .Y(ori_ori_n1196_));
  NO2        o1168(.A(ori_ori_n1196_), .B(ori_ori_n163_), .Y(ori_ori_n1197_));
  NO2        o1169(.A(ori_ori_n48_), .B(l), .Y(ori_ori_n1198_));
  INV        o1170(.A(ori_ori_n434_), .Y(ori_ori_n1199_));
  NA2        o1171(.A(ori_ori_n1199_), .B(ori_ori_n1198_), .Y(ori_ori_n1200_));
  INV        o1172(.A(ori_ori_n1200_), .Y(ori_ori_n1201_));
  NO3        o1173(.A(ori_ori_n1201_), .B(ori_ori_n1197_), .C(ori_ori_n1195_), .Y(ori_ori_n1202_));
  NA2        o1174(.A(ori_ori_n1202_), .B(ori_ori_n1192_), .Y(ori_ori_n1203_));
  NA3        o1175(.A(ori_ori_n852_), .B(ori_ori_n126_), .C(ori_ori_n45_), .Y(ori_ori_n1204_));
  NO2        o1176(.A(ori_ori_n1155_), .B(d), .Y(ori_ori_n1205_));
  NA3        o1177(.A(ori_ori_n1211_), .B(ori_ori_n1212_), .C(ori_ori_n1204_), .Y(ori_ori_n1206_));
  OR4        o1178(.A(ori_ori_n1206_), .B(ori_ori_n1203_), .C(ori_ori_n1182_), .D(ori_ori_n1159_), .Y(ori04));
  INV        o1179(.A(ori_ori_n103_), .Y(ori_ori_n1210_));
  INV        o1180(.A(ori_ori_n1205_), .Y(ori_ori_n1211_));
  INV        o1181(.A(ori_ori_n1116_), .Y(ori_ori_n1212_));
  ZERO       o1182(.Y(ori02));
  ZERO       o1183(.Y(ori03));
  ZERO       o1184(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  INV        m0015(.A(i), .Y(mai_mai_n44_));
  AN2        m0016(.A(h), .B(g), .Y(mai_mai_n45_));
  NA2        m0017(.A(mai_mai_n45_), .B(mai_mai_n44_), .Y(mai_mai_n46_));
  NAi21      m0018(.An(n), .B(m), .Y(mai_mai_n47_));
  NOi32      m0019(.An(k), .Bn(h), .C(l), .Y(mai_mai_n48_));
  NOi32      m0020(.An(k), .Bn(h), .C(g), .Y(mai_mai_n49_));
  INV        m0021(.A(mai_mai_n49_), .Y(mai_mai_n50_));
  NO2        m0022(.A(mai_mai_n50_), .B(mai_mai_n47_), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n43_), .B(mai_mai_n39_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n32_), .Y(mai_mai_n53_));
  INV        m0025(.A(c), .Y(mai_mai_n54_));
  NA2        m0026(.A(e), .B(b), .Y(mai_mai_n55_));
  NO2        m0027(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  INV        m0028(.A(d), .Y(mai_mai_n57_));
  NAi21      m0029(.An(i), .B(h), .Y(mai_mai_n58_));
  NAi31      m0030(.An(i), .B(l), .C(j), .Y(mai_mai_n59_));
  NAi41      m0031(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n60_));
  NA2        m0032(.A(g), .B(f), .Y(mai_mai_n61_));
  NO2        m0033(.A(mai_mai_n61_), .B(mai_mai_n60_), .Y(mai_mai_n62_));
  NAi21      m0034(.An(i), .B(j), .Y(mai_mai_n63_));
  NAi32      m0035(.An(n), .Bn(k), .C(m), .Y(mai_mai_n64_));
  NO2        m0036(.A(mai_mai_n64_), .B(mai_mai_n63_), .Y(mai_mai_n65_));
  NAi31      m0037(.An(l), .B(m), .C(k), .Y(mai_mai_n66_));
  NAi41      m0038(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n67_));
  NA2        m0039(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n68_));
  INV        m0040(.A(m), .Y(mai_mai_n69_));
  NOi21      m0041(.An(k), .B(l), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n70_), .B(mai_mai_n69_), .Y(mai_mai_n71_));
  AN4        m0043(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n72_));
  NOi31      m0044(.An(h), .B(g), .C(f), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  NAi32      m0046(.An(m), .Bn(k), .C(j), .Y(mai_mai_n75_));
  NOi32      m0047(.An(h), .Bn(g), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n72_), .Y(mai_mai_n77_));
  OA220      m0049(.A0(mai_mai_n77_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .B1(mai_mai_n71_), .Y(mai_mai_n78_));
  NA2        m0050(.A(mai_mai_n78_), .B(mai_mai_n68_), .Y(mai_mai_n79_));
  INV        m0051(.A(n), .Y(mai_mai_n80_));
  NOi32      m0052(.An(e), .Bn(b), .C(d), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n80_), .Y(mai_mai_n82_));
  INV        m0054(.A(j), .Y(mai_mai_n83_));
  AN3        m0055(.A(m), .B(k), .C(i), .Y(mai_mai_n84_));
  NA3        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n85_));
  NAi32      m0057(.An(g), .Bn(f), .C(h), .Y(mai_mai_n86_));
  NAi31      m0058(.An(j), .B(m), .C(l), .Y(mai_mai_n87_));
  NA2        m0059(.A(m), .B(l), .Y(mai_mai_n88_));
  NAi31      m0060(.An(k), .B(j), .C(g), .Y(mai_mai_n89_));
  AN2        m0061(.A(j), .B(g), .Y(mai_mai_n90_));
  NOi32      m0062(.An(m), .Bn(l), .C(i), .Y(mai_mai_n91_));
  NOi21      m0063(.An(g), .B(i), .Y(mai_mai_n92_));
  NAi41      m0064(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n93_));
  AN2        m0065(.A(e), .B(b), .Y(mai_mai_n94_));
  NOi31      m0066(.An(c), .B(h), .C(f), .Y(mai_mai_n95_));
  NA2        m0067(.A(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  NO2        m0068(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n97_));
  NOi21      m0069(.An(i), .B(h), .Y(mai_mai_n98_));
  NA3        m0070(.A(mai_mai_n98_), .B(g), .C(mai_mai_n36_), .Y(mai_mai_n99_));
  INV        m0071(.A(a), .Y(mai_mai_n100_));
  NA2        m0072(.A(mai_mai_n94_), .B(mai_mai_n100_), .Y(mai_mai_n101_));
  INV        m0073(.A(l), .Y(mai_mai_n102_));
  NOi21      m0074(.An(m), .B(n), .Y(mai_mai_n103_));
  AN2        m0075(.A(k), .B(h), .Y(mai_mai_n104_));
  NO2        m0076(.A(mai_mai_n99_), .B(mai_mai_n82_), .Y(mai_mai_n105_));
  INV        m0077(.A(b), .Y(mai_mai_n106_));
  NA2        m0078(.A(l), .B(j), .Y(mai_mai_n107_));
  AN2        m0079(.A(k), .B(i), .Y(mai_mai_n108_));
  NA2        m0080(.A(g), .B(e), .Y(mai_mai_n109_));
  NOi32      m0081(.An(c), .Bn(a), .C(d), .Y(mai_mai_n110_));
  NA2        m0082(.A(mai_mai_n110_), .B(mai_mai_n103_), .Y(mai_mai_n111_));
  NO4        m0083(.A(mai_mai_n111_), .B(mai_mai_n109_), .C(mai_mai_n1430_), .D(mai_mai_n106_), .Y(mai_mai_n112_));
  NO3        m0084(.A(mai_mai_n112_), .B(mai_mai_n105_), .C(mai_mai_n97_), .Y(mai_mai_n113_));
  INV        m0085(.A(mai_mai_n113_), .Y(mai_mai_n114_));
  NOi31      m0086(.An(k), .B(m), .C(j), .Y(mai_mai_n115_));
  NOi31      m0087(.An(k), .B(m), .C(i), .Y(mai_mai_n116_));
  NOi32      m0088(.An(f), .Bn(b), .C(e), .Y(mai_mai_n117_));
  NAi21      m0089(.An(g), .B(h), .Y(mai_mai_n118_));
  NAi21      m0090(.An(m), .B(n), .Y(mai_mai_n119_));
  NAi21      m0091(.An(j), .B(k), .Y(mai_mai_n120_));
  NO3        m0092(.A(mai_mai_n120_), .B(mai_mai_n119_), .C(mai_mai_n118_), .Y(mai_mai_n121_));
  NAi41      m0093(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n122_));
  NAi31      m0094(.An(j), .B(k), .C(h), .Y(mai_mai_n123_));
  NA2        m0095(.A(mai_mai_n121_), .B(mai_mai_n117_), .Y(mai_mai_n124_));
  NO2        m0096(.A(k), .B(j), .Y(mai_mai_n125_));
  AN2        m0097(.A(k), .B(j), .Y(mai_mai_n126_));
  NAi21      m0098(.An(c), .B(b), .Y(mai_mai_n127_));
  NA2        m0099(.A(f), .B(d), .Y(mai_mai_n128_));
  NA2        m0100(.A(h), .B(c), .Y(mai_mai_n129_));
  NAi31      m0101(.An(f), .B(e), .C(b), .Y(mai_mai_n130_));
  NA2        m0102(.A(d), .B(b), .Y(mai_mai_n131_));
  NAi21      m0103(.An(e), .B(f), .Y(mai_mai_n132_));
  NO2        m0104(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n133_));
  NA2        m0105(.A(b), .B(a), .Y(mai_mai_n134_));
  NAi21      m0106(.An(e), .B(g), .Y(mai_mai_n135_));
  NAi21      m0107(.An(c), .B(d), .Y(mai_mai_n136_));
  NAi31      m0108(.An(l), .B(k), .C(h), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n119_), .B(mai_mai_n137_), .Y(mai_mai_n138_));
  INV        m0110(.A(mai_mai_n124_), .Y(mai_mai_n139_));
  NAi31      m0111(.An(e), .B(f), .C(b), .Y(mai_mai_n140_));
  NOi21      m0112(.An(g), .B(d), .Y(mai_mai_n141_));
  NO2        m0113(.A(mai_mai_n141_), .B(mai_mai_n140_), .Y(mai_mai_n142_));
  NOi21      m0114(.An(h), .B(i), .Y(mai_mai_n143_));
  NOi21      m0115(.An(k), .B(m), .Y(mai_mai_n144_));
  NA3        m0116(.A(mai_mai_n144_), .B(mai_mai_n143_), .C(n), .Y(mai_mai_n145_));
  NOi21      m0117(.An(mai_mai_n142_), .B(mai_mai_n145_), .Y(mai_mai_n146_));
  NOi21      m0118(.An(h), .B(g), .Y(mai_mai_n147_));
  NO2        m0119(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n148_));
  NA2        m0120(.A(mai_mai_n148_), .B(mai_mai_n147_), .Y(mai_mai_n149_));
  NOi32      m0121(.An(n), .Bn(k), .C(m), .Y(mai_mai_n150_));
  NA2        m0122(.A(l), .B(i), .Y(mai_mai_n151_));
  NA2        m0123(.A(mai_mai_n151_), .B(mai_mai_n150_), .Y(mai_mai_n152_));
  NO2        m0124(.A(mai_mai_n152_), .B(mai_mai_n149_), .Y(mai_mai_n153_));
  NAi31      m0125(.An(d), .B(f), .C(c), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(c), .Y(mai_mai_n155_));
  NA2        m0127(.A(mai_mai_n155_), .B(mai_mai_n154_), .Y(mai_mai_n156_));
  NA2        m0128(.A(j), .B(h), .Y(mai_mai_n157_));
  OR3        m0129(.A(n), .B(m), .C(k), .Y(mai_mai_n158_));
  NO2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NAi32      m0131(.An(m), .Bn(k), .C(n), .Y(mai_mai_n160_));
  NO2        m0132(.A(mai_mai_n160_), .B(mai_mai_n157_), .Y(mai_mai_n161_));
  AOI220     m0133(.A0(mai_mai_n161_), .A1(mai_mai_n142_), .B0(mai_mai_n159_), .B1(mai_mai_n156_), .Y(mai_mai_n162_));
  NO2        m0134(.A(n), .B(m), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n48_), .Y(mai_mai_n164_));
  NAi21      m0136(.An(f), .B(e), .Y(mai_mai_n165_));
  NA2        m0137(.A(d), .B(c), .Y(mai_mai_n166_));
  NO2        m0138(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  NOi21      m0139(.An(mai_mai_n167_), .B(mai_mai_n164_), .Y(mai_mai_n168_));
  NAi21      m0140(.An(d), .B(c), .Y(mai_mai_n169_));
  NAi31      m0141(.An(m), .B(n), .C(b), .Y(mai_mai_n170_));
  NA2        m0142(.A(k), .B(i), .Y(mai_mai_n171_));
  NAi21      m0143(.An(h), .B(f), .Y(mai_mai_n172_));
  NO2        m0144(.A(mai_mai_n172_), .B(mai_mai_n171_), .Y(mai_mai_n173_));
  NO2        m0145(.A(mai_mai_n170_), .B(mai_mai_n136_), .Y(mai_mai_n174_));
  NA2        m0146(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NOi32      m0147(.An(f), .Bn(c), .C(d), .Y(mai_mai_n176_));
  NOi32      m0148(.An(f), .Bn(c), .C(e), .Y(mai_mai_n177_));
  NO2        m0149(.A(mai_mai_n177_), .B(mai_mai_n176_), .Y(mai_mai_n178_));
  NO3        m0150(.A(n), .B(m), .C(j), .Y(mai_mai_n179_));
  NA2        m0151(.A(mai_mai_n179_), .B(mai_mai_n104_), .Y(mai_mai_n180_));
  AO210      m0152(.A0(mai_mai_n180_), .A1(mai_mai_n164_), .B0(mai_mai_n178_), .Y(mai_mai_n181_));
  NAi41      m0153(.An(mai_mai_n168_), .B(mai_mai_n181_), .C(mai_mai_n175_), .D(mai_mai_n162_), .Y(mai_mai_n182_));
  OR4        m0154(.A(mai_mai_n182_), .B(mai_mai_n153_), .C(mai_mai_n146_), .D(mai_mai_n139_), .Y(mai_mai_n183_));
  NO4        m0155(.A(mai_mai_n183_), .B(mai_mai_n114_), .C(mai_mai_n79_), .D(mai_mai_n53_), .Y(mai_mai_n184_));
  NAi31      m0156(.An(n), .B(h), .C(g), .Y(mai_mai_n185_));
  NOi32      m0157(.An(m), .Bn(k), .C(l), .Y(mai_mai_n186_));
  NA3        m0158(.A(mai_mai_n186_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n187_), .B(n), .Y(mai_mai_n188_));
  NOi21      m0160(.An(k), .B(j), .Y(mai_mai_n189_));
  NA4        m0161(.A(mai_mai_n189_), .B(mai_mai_n103_), .C(i), .D(g), .Y(mai_mai_n190_));
  AN2        m0162(.A(i), .B(g), .Y(mai_mai_n191_));
  NA3        m0163(.A(mai_mai_n70_), .B(mai_mai_n191_), .C(mai_mai_n103_), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n190_), .Y(mai_mai_n193_));
  INV        m0165(.A(mai_mai_n193_), .Y(mai_mai_n194_));
  NAi41      m0166(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n195_));
  INV        m0167(.A(f), .Y(mai_mai_n196_));
  INV        m0168(.A(g), .Y(mai_mai_n197_));
  NOi31      m0169(.An(i), .B(j), .C(h), .Y(mai_mai_n198_));
  NOi21      m0170(.An(l), .B(m), .Y(mai_mai_n199_));
  NA2        m0171(.A(mai_mai_n199_), .B(mai_mai_n198_), .Y(mai_mai_n200_));
  NO2        m0172(.A(mai_mai_n194_), .B(mai_mai_n32_), .Y(mai_mai_n201_));
  NOi21      m0173(.An(n), .B(m), .Y(mai_mai_n202_));
  NOi32      m0174(.An(l), .Bn(i), .C(j), .Y(mai_mai_n203_));
  NA2        m0175(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  OA220      m0176(.A0(mai_mai_n204_), .A1(mai_mai_n96_), .B0(mai_mai_n75_), .B1(mai_mai_n74_), .Y(mai_mai_n205_));
  NAi21      m0177(.An(j), .B(h), .Y(mai_mai_n206_));
  XN2        m0178(.A(i), .B(h), .Y(mai_mai_n207_));
  NA2        m0179(.A(mai_mai_n207_), .B(mai_mai_n206_), .Y(mai_mai_n208_));
  NOi31      m0180(.An(k), .B(n), .C(m), .Y(mai_mai_n209_));
  NOi31      m0181(.An(mai_mai_n209_), .B(mai_mai_n166_), .C(mai_mai_n165_), .Y(mai_mai_n210_));
  NA2        m0182(.A(mai_mai_n210_), .B(mai_mai_n208_), .Y(mai_mai_n211_));
  NAi31      m0183(.An(f), .B(e), .C(c), .Y(mai_mai_n212_));
  NO4        m0184(.A(mai_mai_n212_), .B(mai_mai_n158_), .C(mai_mai_n157_), .D(mai_mai_n57_), .Y(mai_mai_n213_));
  NA4        m0185(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n214_));
  NAi32      m0186(.An(m), .Bn(i), .C(k), .Y(mai_mai_n215_));
  NO3        m0187(.A(mai_mai_n215_), .B(mai_mai_n86_), .C(mai_mai_n214_), .Y(mai_mai_n216_));
  INV        m0188(.A(k), .Y(mai_mai_n217_));
  NO2        m0189(.A(mai_mai_n216_), .B(mai_mai_n213_), .Y(mai_mai_n218_));
  NAi21      m0190(.An(n), .B(a), .Y(mai_mai_n219_));
  NO2        m0191(.A(mai_mai_n219_), .B(mai_mai_n131_), .Y(mai_mai_n220_));
  NAi41      m0192(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n221_));
  NO2        m0193(.A(mai_mai_n221_), .B(e), .Y(mai_mai_n222_));
  NO2        m0194(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n223_));
  OAI210     m0195(.A0(mai_mai_n223_), .A1(mai_mai_n222_), .B0(mai_mai_n220_), .Y(mai_mai_n224_));
  AN4        m0196(.A(mai_mai_n224_), .B(mai_mai_n218_), .C(mai_mai_n211_), .D(mai_mai_n205_), .Y(mai_mai_n225_));
  OR2        m0197(.A(h), .B(g), .Y(mai_mai_n226_));
  NO2        m0198(.A(mai_mai_n226_), .B(mai_mai_n93_), .Y(mai_mai_n227_));
  NA2        m0199(.A(mai_mai_n227_), .B(mai_mai_n117_), .Y(mai_mai_n228_));
  NAi41      m0200(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n229_));
  NO2        m0201(.A(mai_mai_n229_), .B(mai_mai_n196_), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n144_), .B(mai_mai_n98_), .Y(mai_mai_n231_));
  NAi21      m0203(.An(mai_mai_n231_), .B(mai_mai_n230_), .Y(mai_mai_n232_));
  NO2        m0204(.A(n), .B(a), .Y(mai_mai_n233_));
  NAi31      m0205(.An(mai_mai_n221_), .B(mai_mai_n233_), .C(mai_mai_n94_), .Y(mai_mai_n234_));
  AN2        m0206(.A(mai_mai_n234_), .B(mai_mai_n232_), .Y(mai_mai_n235_));
  NAi21      m0207(.An(h), .B(i), .Y(mai_mai_n236_));
  NA2        m0208(.A(mai_mai_n163_), .B(k), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  NA2        m0210(.A(mai_mai_n238_), .B(mai_mai_n176_), .Y(mai_mai_n239_));
  NA3        m0211(.A(mai_mai_n239_), .B(mai_mai_n235_), .C(mai_mai_n228_), .Y(mai_mai_n240_));
  NOi21      m0212(.An(g), .B(e), .Y(mai_mai_n241_));
  NAi21      m0213(.An(f), .B(g), .Y(mai_mai_n242_));
  NO2        m0214(.A(mai_mai_n64_), .B(mai_mai_n107_), .Y(mai_mai_n243_));
  NO3        m0215(.A(mai_mai_n120_), .B(mai_mai_n47_), .C(mai_mai_n44_), .Y(mai_mai_n244_));
  NOi31      m0216(.An(mai_mai_n225_), .B(mai_mai_n240_), .C(mai_mai_n201_), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n43_), .B(mai_mai_n39_), .Y(mai_mai_n246_));
  NO2        m0218(.A(mai_mai_n246_), .B(mai_mai_n101_), .Y(mai_mai_n247_));
  NA3        m0219(.A(mai_mai_n57_), .B(c), .C(b), .Y(mai_mai_n248_));
  NAi21      m0220(.An(h), .B(g), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n231_), .B(mai_mai_n242_), .Y(mai_mai_n250_));
  NAi31      m0222(.An(g), .B(k), .C(h), .Y(mai_mai_n251_));
  NO3        m0223(.A(mai_mai_n119_), .B(mai_mai_n251_), .C(l), .Y(mai_mai_n252_));
  NAi31      m0224(.An(e), .B(d), .C(a), .Y(mai_mai_n253_));
  NA2        m0225(.A(mai_mai_n252_), .B(mai_mai_n117_), .Y(mai_mai_n254_));
  INV        m0226(.A(mai_mai_n254_), .Y(mai_mai_n255_));
  NA4        m0227(.A(mai_mai_n144_), .B(mai_mai_n76_), .C(mai_mai_n72_), .D(mai_mai_n107_), .Y(mai_mai_n256_));
  NA3        m0228(.A(mai_mai_n144_), .B(mai_mai_n143_), .C(mai_mai_n80_), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n257_), .B(mai_mai_n178_), .Y(mai_mai_n258_));
  NOi21      m0230(.An(mai_mai_n256_), .B(mai_mai_n258_), .Y(mai_mai_n259_));
  NA3        m0231(.A(e), .B(c), .C(b), .Y(mai_mai_n260_));
  NAi21      m0232(.An(l), .B(k), .Y(mai_mai_n261_));
  NO2        m0233(.A(mai_mai_n261_), .B(mai_mai_n47_), .Y(mai_mai_n262_));
  NOi21      m0234(.An(l), .B(j), .Y(mai_mai_n263_));
  NA2        m0235(.A(mai_mai_n147_), .B(mai_mai_n263_), .Y(mai_mai_n264_));
  NA3        m0236(.A(mai_mai_n108_), .B(mai_mai_n107_), .C(g), .Y(mai_mai_n265_));
  OR3        m0237(.A(mai_mai_n67_), .B(mai_mai_n69_), .C(e), .Y(mai_mai_n266_));
  AOI210     m0238(.A0(mai_mai_n265_), .A1(mai_mai_n264_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  INV        m0239(.A(mai_mai_n267_), .Y(mai_mai_n268_));
  NAi32      m0240(.An(j), .Bn(h), .C(i), .Y(mai_mai_n269_));
  NAi21      m0241(.An(m), .B(l), .Y(mai_mai_n270_));
  NO3        m0242(.A(mai_mai_n270_), .B(mai_mai_n269_), .C(mai_mai_n80_), .Y(mai_mai_n271_));
  NA2        m0243(.A(h), .B(g), .Y(mai_mai_n272_));
  NA2        m0244(.A(mai_mai_n271_), .B(mai_mai_n148_), .Y(mai_mai_n273_));
  NA3        m0245(.A(mai_mai_n273_), .B(mai_mai_n268_), .C(mai_mai_n259_), .Y(mai_mai_n274_));
  NO2        m0246(.A(mai_mai_n130_), .B(d), .Y(mai_mai_n275_));
  NA2        m0247(.A(mai_mai_n275_), .B(mai_mai_n51_), .Y(mai_mai_n276_));
  NO2        m0248(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n277_));
  NAi32      m0249(.An(n), .Bn(m), .C(l), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n278_), .B(mai_mai_n269_), .Y(mai_mai_n279_));
  NA2        m0251(.A(mai_mai_n279_), .B(mai_mai_n167_), .Y(mai_mai_n280_));
  NO2        m0252(.A(mai_mai_n111_), .B(mai_mai_n106_), .Y(mai_mai_n281_));
  NAi31      m0253(.An(k), .B(l), .C(j), .Y(mai_mai_n282_));
  NA2        m0254(.A(mai_mai_n261_), .B(mai_mai_n282_), .Y(mai_mai_n283_));
  NOi21      m0255(.An(mai_mai_n283_), .B(mai_mai_n109_), .Y(mai_mai_n284_));
  NA2        m0256(.A(mai_mai_n284_), .B(mai_mai_n281_), .Y(mai_mai_n285_));
  NA3        m0257(.A(mai_mai_n285_), .B(mai_mai_n280_), .C(mai_mai_n276_), .Y(mai_mai_n286_));
  NO4        m0258(.A(mai_mai_n286_), .B(mai_mai_n274_), .C(mai_mai_n255_), .D(mai_mai_n247_), .Y(mai_mai_n287_));
  NA2        m0259(.A(mai_mai_n238_), .B(mai_mai_n177_), .Y(mai_mai_n288_));
  NAi21      m0260(.An(m), .B(k), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n207_), .B(mai_mai_n289_), .Y(mai_mai_n290_));
  NAi41      m0262(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n291_));
  NO2        m0263(.A(mai_mai_n291_), .B(mai_mai_n135_), .Y(mai_mai_n292_));
  NA2        m0264(.A(mai_mai_n292_), .B(mai_mai_n290_), .Y(mai_mai_n293_));
  NA2        m0265(.A(e), .B(c), .Y(mai_mai_n294_));
  NO3        m0266(.A(mai_mai_n294_), .B(n), .C(d), .Y(mai_mai_n295_));
  NOi21      m0267(.An(f), .B(h), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n296_), .B(mai_mai_n108_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n297_), .B(mai_mai_n197_), .Y(mai_mai_n298_));
  NAi31      m0270(.An(d), .B(e), .C(b), .Y(mai_mai_n299_));
  NO2        m0271(.A(mai_mai_n119_), .B(mai_mai_n299_), .Y(mai_mai_n300_));
  NA2        m0272(.A(mai_mai_n300_), .B(mai_mai_n298_), .Y(mai_mai_n301_));
  NA3        m0273(.A(mai_mai_n301_), .B(mai_mai_n293_), .C(mai_mai_n288_), .Y(mai_mai_n302_));
  NA2        m0274(.A(mai_mai_n233_), .B(mai_mai_n94_), .Y(mai_mai_n303_));
  OR2        m0275(.A(mai_mai_n303_), .B(mai_mai_n187_), .Y(mai_mai_n304_));
  NOi31      m0276(.An(l), .B(n), .C(m), .Y(mai_mai_n305_));
  NA2        m0277(.A(mai_mai_n305_), .B(mai_mai_n198_), .Y(mai_mai_n306_));
  NO2        m0278(.A(mai_mai_n306_), .B(mai_mai_n178_), .Y(mai_mai_n307_));
  NAi21      m0279(.An(mai_mai_n307_), .B(mai_mai_n304_), .Y(mai_mai_n308_));
  NAi32      m0280(.An(m), .Bn(j), .C(k), .Y(mai_mai_n309_));
  NAi41      m0281(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n195_), .B(mai_mai_n310_), .Y(mai_mai_n311_));
  NOi31      m0283(.An(j), .B(m), .C(k), .Y(mai_mai_n312_));
  NO2        m0284(.A(mai_mai_n115_), .B(mai_mai_n312_), .Y(mai_mai_n313_));
  AN3        m0285(.A(h), .B(g), .C(f), .Y(mai_mai_n314_));
  NAi31      m0286(.An(mai_mai_n313_), .B(mai_mai_n314_), .C(mai_mai_n311_), .Y(mai_mai_n315_));
  NOi32      m0287(.An(m), .Bn(j), .C(l), .Y(mai_mai_n316_));
  NO2        m0288(.A(mai_mai_n316_), .B(mai_mai_n91_), .Y(mai_mai_n317_));
  NAi32      m0289(.An(mai_mai_n317_), .Bn(mai_mai_n185_), .C(mai_mai_n275_), .Y(mai_mai_n318_));
  NO2        m0290(.A(mai_mai_n270_), .B(mai_mai_n269_), .Y(mai_mai_n319_));
  NO2        m0291(.A(mai_mai_n200_), .B(g), .Y(mai_mai_n320_));
  NO2        m0292(.A(mai_mai_n140_), .B(mai_mai_n80_), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n318_), .B(mai_mai_n315_), .Y(mai_mai_n322_));
  NA3        m0294(.A(h), .B(g), .C(f), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n323_), .B(mai_mai_n71_), .Y(mai_mai_n324_));
  NA2        m0296(.A(mai_mai_n310_), .B(mai_mai_n195_), .Y(mai_mai_n325_));
  NA2        m0297(.A(mai_mai_n147_), .B(e), .Y(mai_mai_n326_));
  NO2        m0298(.A(mai_mai_n326_), .B(mai_mai_n41_), .Y(mai_mai_n327_));
  AOI220     m0299(.A0(mai_mai_n327_), .A1(mai_mai_n281_), .B0(mai_mai_n325_), .B1(mai_mai_n324_), .Y(mai_mai_n328_));
  NOi32      m0300(.An(j), .Bn(g), .C(i), .Y(mai_mai_n329_));
  NA3        m0301(.A(mai_mai_n329_), .B(mai_mai_n261_), .C(mai_mai_n103_), .Y(mai_mai_n330_));
  NOi32      m0302(.An(e), .Bn(b), .C(a), .Y(mai_mai_n331_));
  AN2        m0303(.A(l), .B(j), .Y(mai_mai_n332_));
  NA3        m0304(.A(mai_mai_n192_), .B(mai_mai_n190_), .C(mai_mai_n35_), .Y(mai_mai_n333_));
  NA2        m0305(.A(mai_mai_n333_), .B(mai_mai_n331_), .Y(mai_mai_n334_));
  NO2        m0306(.A(mai_mai_n299_), .B(n), .Y(mai_mai_n335_));
  NA2        m0307(.A(mai_mai_n191_), .B(k), .Y(mai_mai_n336_));
  NA3        m0308(.A(m), .B(mai_mai_n102_), .C(mai_mai_n196_), .Y(mai_mai_n337_));
  NA3        m0309(.A(mai_mai_n186_), .B(mai_mai_n83_), .C(g), .Y(mai_mai_n338_));
  INV        m0310(.A(mai_mai_n338_), .Y(mai_mai_n339_));
  NAi41      m0311(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n340_));
  NA2        m0312(.A(mai_mai_n49_), .B(mai_mai_n103_), .Y(mai_mai_n341_));
  NO2        m0313(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n342_));
  AOI220     m0314(.A0(mai_mai_n342_), .A1(b), .B0(mai_mai_n339_), .B1(mai_mai_n335_), .Y(mai_mai_n343_));
  NA3        m0315(.A(mai_mai_n343_), .B(mai_mai_n334_), .C(mai_mai_n328_), .Y(mai_mai_n344_));
  NO4        m0316(.A(mai_mai_n344_), .B(mai_mai_n322_), .C(mai_mai_n308_), .D(mai_mai_n302_), .Y(mai_mai_n345_));
  NA4        m0317(.A(mai_mai_n345_), .B(mai_mai_n287_), .C(mai_mai_n245_), .D(mai_mai_n184_), .Y(mai10));
  NA3        m0318(.A(m), .B(k), .C(i), .Y(mai_mai_n347_));
  NO3        m0319(.A(mai_mai_n347_), .B(j), .C(mai_mai_n197_), .Y(mai_mai_n348_));
  NOi21      m0320(.An(e), .B(f), .Y(mai_mai_n349_));
  NO4        m0321(.A(mai_mai_n136_), .B(mai_mai_n349_), .C(n), .D(mai_mai_n100_), .Y(mai_mai_n350_));
  NAi31      m0322(.An(b), .B(f), .C(c), .Y(mai_mai_n351_));
  INV        m0323(.A(mai_mai_n351_), .Y(mai_mai_n352_));
  NOi32      m0324(.An(k), .Bn(h), .C(j), .Y(mai_mai_n353_));
  NA2        m0325(.A(mai_mai_n353_), .B(mai_mai_n202_), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n145_), .B(mai_mai_n354_), .Y(mai_mai_n355_));
  NA2        m0327(.A(mai_mai_n355_), .B(mai_mai_n352_), .Y(mai_mai_n356_));
  AN2        m0328(.A(j), .B(h), .Y(mai_mai_n357_));
  NO3        m0329(.A(n), .B(m), .C(k), .Y(mai_mai_n358_));
  NA2        m0330(.A(mai_mai_n358_), .B(mai_mai_n357_), .Y(mai_mai_n359_));
  NO3        m0331(.A(mai_mai_n359_), .B(mai_mai_n136_), .C(mai_mai_n196_), .Y(mai_mai_n360_));
  OR2        m0332(.A(m), .B(k), .Y(mai_mai_n361_));
  NO2        m0333(.A(mai_mai_n157_), .B(mai_mai_n361_), .Y(mai_mai_n362_));
  NA4        m0334(.A(n), .B(f), .C(c), .D(mai_mai_n106_), .Y(mai_mai_n363_));
  NOi21      m0335(.An(mai_mai_n362_), .B(mai_mai_n363_), .Y(mai_mai_n364_));
  NOi32      m0336(.An(d), .Bn(a), .C(c), .Y(mai_mai_n365_));
  NA2        m0337(.A(mai_mai_n365_), .B(mai_mai_n165_), .Y(mai_mai_n366_));
  NAi21      m0338(.An(i), .B(g), .Y(mai_mai_n367_));
  NAi31      m0339(.An(k), .B(m), .C(j), .Y(mai_mai_n368_));
  NO3        m0340(.A(mai_mai_n368_), .B(mai_mai_n367_), .C(n), .Y(mai_mai_n369_));
  NOi21      m0341(.An(mai_mai_n369_), .B(mai_mai_n366_), .Y(mai_mai_n370_));
  NO3        m0342(.A(mai_mai_n370_), .B(mai_mai_n364_), .C(mai_mai_n360_), .Y(mai_mai_n371_));
  NO2        m0343(.A(mai_mai_n363_), .B(mai_mai_n270_), .Y(mai_mai_n372_));
  NOi32      m0344(.An(f), .Bn(d), .C(c), .Y(mai_mai_n373_));
  AOI220     m0345(.A0(mai_mai_n373_), .A1(mai_mai_n279_), .B0(mai_mai_n372_), .B1(mai_mai_n198_), .Y(mai_mai_n374_));
  NA3        m0346(.A(mai_mai_n374_), .B(mai_mai_n371_), .C(mai_mai_n356_), .Y(mai_mai_n375_));
  NO2        m0347(.A(mai_mai_n57_), .B(mai_mai_n106_), .Y(mai_mai_n376_));
  NA2        m0348(.A(mai_mai_n233_), .B(mai_mai_n376_), .Y(mai_mai_n377_));
  INV        m0349(.A(e), .Y(mai_mai_n378_));
  NA2        m0350(.A(mai_mai_n45_), .B(e), .Y(mai_mai_n379_));
  AN2        m0351(.A(g), .B(e), .Y(mai_mai_n380_));
  NA3        m0352(.A(mai_mai_n380_), .B(mai_mai_n186_), .C(i), .Y(mai_mai_n381_));
  OAI210     m0353(.A0(mai_mai_n85_), .A1(mai_mai_n378_), .B0(mai_mai_n381_), .Y(mai_mai_n382_));
  INV        m0354(.A(mai_mai_n382_), .Y(mai_mai_n383_));
  NOi32      m0355(.An(h), .Bn(e), .C(g), .Y(mai_mai_n384_));
  NA3        m0356(.A(mai_mai_n384_), .B(mai_mai_n263_), .C(m), .Y(mai_mai_n385_));
  NOi21      m0357(.An(g), .B(h), .Y(mai_mai_n386_));
  AN3        m0358(.A(m), .B(l), .C(i), .Y(mai_mai_n387_));
  NA3        m0359(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(e), .Y(mai_mai_n388_));
  AN3        m0360(.A(h), .B(g), .C(e), .Y(mai_mai_n389_));
  NA2        m0361(.A(mai_mai_n389_), .B(mai_mai_n91_), .Y(mai_mai_n390_));
  AN3        m0362(.A(mai_mai_n390_), .B(mai_mai_n388_), .C(mai_mai_n385_), .Y(mai_mai_n391_));
  AOI210     m0363(.A0(mai_mai_n391_), .A1(mai_mai_n383_), .B0(mai_mai_n377_), .Y(mai_mai_n392_));
  NA3        m0364(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n393_));
  NO2        m0365(.A(mai_mai_n393_), .B(mai_mai_n377_), .Y(mai_mai_n394_));
  NA3        m0366(.A(mai_mai_n365_), .B(mai_mai_n165_), .C(mai_mai_n80_), .Y(mai_mai_n395_));
  NAi31      m0367(.An(b), .B(c), .C(a), .Y(mai_mai_n396_));
  NO2        m0368(.A(mai_mai_n396_), .B(n), .Y(mai_mai_n397_));
  NA2        m0369(.A(mai_mai_n49_), .B(m), .Y(mai_mai_n398_));
  NO2        m0370(.A(mai_mai_n398_), .B(mai_mai_n132_), .Y(mai_mai_n399_));
  NA2        m0371(.A(mai_mai_n399_), .B(mai_mai_n397_), .Y(mai_mai_n400_));
  INV        m0372(.A(mai_mai_n400_), .Y(mai_mai_n401_));
  NO4        m0373(.A(mai_mai_n401_), .B(mai_mai_n394_), .C(mai_mai_n392_), .D(mai_mai_n375_), .Y(mai_mai_n402_));
  NA2        m0374(.A(i), .B(g), .Y(mai_mai_n403_));
  NO3        m0375(.A(mai_mai_n253_), .B(mai_mai_n403_), .C(c), .Y(mai_mai_n404_));
  NOi21      m0376(.An(a), .B(n), .Y(mai_mai_n405_));
  NOi21      m0377(.An(d), .B(c), .Y(mai_mai_n406_));
  NA2        m0378(.A(mai_mai_n406_), .B(mai_mai_n405_), .Y(mai_mai_n407_));
  NA3        m0379(.A(i), .B(g), .C(f), .Y(mai_mai_n408_));
  OR2        m0380(.A(mai_mai_n408_), .B(mai_mai_n66_), .Y(mai_mai_n409_));
  NA3        m0381(.A(mai_mai_n387_), .B(mai_mai_n386_), .C(mai_mai_n165_), .Y(mai_mai_n410_));
  AOI210     m0382(.A0(mai_mai_n410_), .A1(mai_mai_n409_), .B0(mai_mai_n407_), .Y(mai_mai_n411_));
  AOI210     m0383(.A0(mai_mai_n404_), .A1(mai_mai_n262_), .B0(mai_mai_n411_), .Y(mai_mai_n412_));
  OR2        m0384(.A(n), .B(m), .Y(mai_mai_n413_));
  NO2        m0385(.A(mai_mai_n413_), .B(mai_mai_n137_), .Y(mai_mai_n414_));
  NO2        m0386(.A(mai_mai_n166_), .B(mai_mai_n132_), .Y(mai_mai_n415_));
  OAI210     m0387(.A0(mai_mai_n414_), .A1(mai_mai_n159_), .B0(mai_mai_n415_), .Y(mai_mai_n416_));
  INV        m0388(.A(mai_mai_n341_), .Y(mai_mai_n417_));
  NA3        m0389(.A(mai_mai_n417_), .B(mai_mai_n331_), .C(d), .Y(mai_mai_n418_));
  NO2        m0390(.A(mai_mai_n396_), .B(mai_mai_n47_), .Y(mai_mai_n419_));
  NO3        m0391(.A(mai_mai_n61_), .B(mai_mai_n102_), .C(e), .Y(mai_mai_n420_));
  NAi21      m0392(.An(k), .B(j), .Y(mai_mai_n421_));
  NA2        m0393(.A(mai_mai_n420_), .B(mai_mai_n419_), .Y(mai_mai_n422_));
  NAi21      m0394(.An(e), .B(d), .Y(mai_mai_n423_));
  INV        m0395(.A(mai_mai_n423_), .Y(mai_mai_n424_));
  NO2        m0396(.A(mai_mai_n237_), .B(mai_mai_n196_), .Y(mai_mai_n425_));
  NA3        m0397(.A(mai_mai_n425_), .B(mai_mai_n424_), .C(mai_mai_n208_), .Y(mai_mai_n426_));
  NA4        m0398(.A(mai_mai_n426_), .B(mai_mai_n422_), .C(mai_mai_n418_), .D(mai_mai_n416_), .Y(mai_mai_n427_));
  NO2        m0399(.A(mai_mai_n306_), .B(mai_mai_n196_), .Y(mai_mai_n428_));
  NA2        m0400(.A(mai_mai_n428_), .B(mai_mai_n424_), .Y(mai_mai_n429_));
  NOi31      m0401(.An(n), .B(m), .C(k), .Y(mai_mai_n430_));
  AOI220     m0402(.A0(mai_mai_n430_), .A1(mai_mai_n357_), .B0(mai_mai_n202_), .B1(mai_mai_n48_), .Y(mai_mai_n431_));
  NAi31      m0403(.An(g), .B(f), .C(c), .Y(mai_mai_n432_));
  NA2        m0404(.A(mai_mai_n429_), .B(mai_mai_n280_), .Y(mai_mai_n433_));
  NOi31      m0405(.An(mai_mai_n412_), .B(mai_mai_n433_), .C(mai_mai_n427_), .Y(mai_mai_n434_));
  NOi32      m0406(.An(c), .Bn(a), .C(b), .Y(mai_mai_n435_));
  NA2        m0407(.A(mai_mai_n435_), .B(mai_mai_n103_), .Y(mai_mai_n436_));
  INV        m0408(.A(mai_mai_n251_), .Y(mai_mai_n437_));
  AN2        m0409(.A(e), .B(d), .Y(mai_mai_n438_));
  NA2        m0410(.A(mai_mai_n438_), .B(mai_mai_n437_), .Y(mai_mai_n439_));
  INV        m0411(.A(mai_mai_n132_), .Y(mai_mai_n440_));
  NO2        m0412(.A(mai_mai_n118_), .B(mai_mai_n41_), .Y(mai_mai_n441_));
  NO2        m0413(.A(mai_mai_n61_), .B(e), .Y(mai_mai_n442_));
  NA2        m0414(.A(k), .B(mai_mai_n442_), .Y(mai_mai_n443_));
  AOI210     m0415(.A0(mai_mai_n443_), .A1(mai_mai_n439_), .B0(mai_mai_n436_), .Y(mai_mai_n444_));
  NO2        m0416(.A(mai_mai_n193_), .B(mai_mai_n188_), .Y(mai_mai_n445_));
  NOi21      m0417(.An(a), .B(b), .Y(mai_mai_n446_));
  NA3        m0418(.A(e), .B(d), .C(c), .Y(mai_mai_n447_));
  NAi21      m0419(.An(mai_mai_n447_), .B(mai_mai_n446_), .Y(mai_mai_n448_));
  NO2        m0420(.A(mai_mai_n395_), .B(mai_mai_n187_), .Y(mai_mai_n449_));
  NOi21      m0421(.An(mai_mai_n448_), .B(mai_mai_n449_), .Y(mai_mai_n450_));
  AOI210     m0422(.A0(mai_mai_n246_), .A1(mai_mai_n445_), .B0(mai_mai_n450_), .Y(mai_mai_n451_));
  NO4        m0423(.A(mai_mai_n172_), .B(mai_mai_n93_), .C(mai_mai_n54_), .D(b), .Y(mai_mai_n452_));
  NA2        m0424(.A(mai_mai_n352_), .B(mai_mai_n138_), .Y(mai_mai_n453_));
  OR2        m0425(.A(k), .B(j), .Y(mai_mai_n454_));
  NA2        m0426(.A(l), .B(k), .Y(mai_mai_n455_));
  NA3        m0427(.A(mai_mai_n455_), .B(mai_mai_n454_), .C(mai_mai_n202_), .Y(mai_mai_n456_));
  AOI210     m0428(.A0(mai_mai_n215_), .A1(mai_mai_n309_), .B0(mai_mai_n80_), .Y(mai_mai_n457_));
  NOi21      m0429(.An(mai_mai_n456_), .B(mai_mai_n457_), .Y(mai_mai_n458_));
  OR3        m0430(.A(mai_mai_n458_), .B(mai_mai_n129_), .C(mai_mai_n122_), .Y(mai_mai_n459_));
  INV        m0431(.A(mai_mai_n256_), .Y(mai_mai_n460_));
  NA2        m0432(.A(mai_mai_n365_), .B(mai_mai_n103_), .Y(mai_mai_n461_));
  NO4        m0433(.A(mai_mai_n461_), .B(mai_mai_n89_), .C(mai_mai_n102_), .D(e), .Y(mai_mai_n462_));
  NO3        m0434(.A(mai_mai_n395_), .B(mai_mai_n87_), .C(mai_mai_n118_), .Y(mai_mai_n463_));
  NO3        m0435(.A(mai_mai_n463_), .B(mai_mai_n462_), .C(mai_mai_n460_), .Y(mai_mai_n464_));
  NA3        m0436(.A(mai_mai_n464_), .B(mai_mai_n459_), .C(mai_mai_n453_), .Y(mai_mai_n465_));
  NO4        m0437(.A(mai_mai_n465_), .B(mai_mai_n452_), .C(mai_mai_n451_), .D(mai_mai_n444_), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n65_), .B(mai_mai_n62_), .Y(mai_mai_n467_));
  NOi21      m0439(.An(d), .B(e), .Y(mai_mai_n468_));
  NO2        m0440(.A(mai_mai_n172_), .B(mai_mai_n54_), .Y(mai_mai_n469_));
  NAi31      m0441(.An(j), .B(l), .C(i), .Y(mai_mai_n470_));
  OAI210     m0442(.A0(mai_mai_n470_), .A1(mai_mai_n119_), .B0(mai_mai_n93_), .Y(mai_mai_n471_));
  NA3        m0443(.A(mai_mai_n471_), .B(mai_mai_n469_), .C(mai_mai_n468_), .Y(mai_mai_n472_));
  NO3        m0444(.A(mai_mai_n366_), .B(mai_mai_n317_), .C(mai_mai_n185_), .Y(mai_mai_n473_));
  NO2        m0445(.A(mai_mai_n366_), .B(mai_mai_n341_), .Y(mai_mai_n474_));
  NO4        m0446(.A(mai_mai_n474_), .B(mai_mai_n473_), .C(mai_mai_n168_), .D(mai_mai_n277_), .Y(mai_mai_n475_));
  NA4        m0447(.A(mai_mai_n475_), .B(mai_mai_n472_), .C(mai_mai_n467_), .D(mai_mai_n225_), .Y(mai_mai_n476_));
  OAI210     m0448(.A0(mai_mai_n116_), .A1(mai_mai_n115_), .B0(n), .Y(mai_mai_n477_));
  NO2        m0449(.A(mai_mai_n477_), .B(mai_mai_n118_), .Y(mai_mai_n478_));
  BUFFER     m0450(.A(mai_mai_n227_), .Y(mai_mai_n479_));
  OA210      m0451(.A0(mai_mai_n479_), .A1(mai_mai_n478_), .B0(mai_mai_n177_), .Y(mai_mai_n480_));
  XO2        m0452(.A(i), .B(h), .Y(mai_mai_n481_));
  NA3        m0453(.A(mai_mai_n481_), .B(mai_mai_n144_), .C(n), .Y(mai_mai_n482_));
  NAi41      m0454(.An(mai_mai_n271_), .B(mai_mai_n482_), .C(mai_mai_n431_), .D(mai_mai_n354_), .Y(mai_mai_n483_));
  NAi31      m0455(.An(c), .B(f), .C(d), .Y(mai_mai_n484_));
  AOI210     m0456(.A0(mai_mai_n257_), .A1(mai_mai_n180_), .B0(mai_mai_n484_), .Y(mai_mai_n485_));
  NOi21      m0457(.An(mai_mai_n78_), .B(mai_mai_n485_), .Y(mai_mai_n486_));
  NA3        m0458(.A(mai_mai_n350_), .B(mai_mai_n91_), .C(mai_mai_n90_), .Y(mai_mai_n487_));
  NA2        m0459(.A(mai_mai_n209_), .B(mai_mai_n98_), .Y(mai_mai_n488_));
  AOI210     m0460(.A0(mai_mai_n488_), .A1(mai_mai_n164_), .B0(mai_mai_n484_), .Y(mai_mai_n489_));
  AOI210     m0461(.A0(mai_mai_n330_), .A1(mai_mai_n35_), .B0(mai_mai_n448_), .Y(mai_mai_n490_));
  NOi31      m0462(.An(mai_mai_n487_), .B(mai_mai_n490_), .C(mai_mai_n489_), .Y(mai_mai_n491_));
  NA3        m0463(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n492_));
  NO2        m0464(.A(mai_mai_n492_), .B(mai_mai_n407_), .Y(mai_mai_n493_));
  NO2        m0465(.A(mai_mai_n493_), .B(mai_mai_n267_), .Y(mai_mai_n494_));
  NA3        m0466(.A(mai_mai_n494_), .B(mai_mai_n491_), .C(mai_mai_n486_), .Y(mai_mai_n495_));
  NO3        m0467(.A(mai_mai_n495_), .B(mai_mai_n480_), .C(mai_mai_n476_), .Y(mai_mai_n496_));
  NA4        m0468(.A(mai_mai_n496_), .B(mai_mai_n466_), .C(mai_mai_n434_), .D(mai_mai_n402_), .Y(mai11));
  NO2        m0469(.A(mai_mai_n67_), .B(f), .Y(mai_mai_n498_));
  NA2        m0470(.A(j), .B(g), .Y(mai_mai_n499_));
  NAi31      m0471(.An(i), .B(m), .C(l), .Y(mai_mai_n500_));
  NA3        m0472(.A(m), .B(k), .C(j), .Y(mai_mai_n501_));
  NOi32      m0473(.An(e), .Bn(b), .C(f), .Y(mai_mai_n502_));
  NA2        m0474(.A(l), .B(mai_mai_n103_), .Y(mai_mai_n503_));
  NA2        m0475(.A(mai_mai_n45_), .B(j), .Y(mai_mai_n504_));
  NAi31      m0476(.An(d), .B(e), .C(a), .Y(mai_mai_n505_));
  NO2        m0477(.A(mai_mai_n505_), .B(n), .Y(mai_mai_n506_));
  NAi41      m0478(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n507_));
  AN2        m0479(.A(mai_mai_n507_), .B(mai_mai_n340_), .Y(mai_mai_n508_));
  AOI210     m0480(.A0(mai_mai_n508_), .A1(mai_mai_n366_), .B0(mai_mai_n249_), .Y(mai_mai_n509_));
  NA2        m0481(.A(j), .B(i), .Y(mai_mai_n510_));
  NAi31      m0482(.An(n), .B(m), .C(k), .Y(mai_mai_n511_));
  NO3        m0483(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n102_), .Y(mai_mai_n512_));
  NO4        m0484(.A(n), .B(d), .C(mai_mai_n106_), .D(a), .Y(mai_mai_n513_));
  OR2        m0485(.A(n), .B(c), .Y(mai_mai_n514_));
  NO2        m0486(.A(mai_mai_n514_), .B(mai_mai_n134_), .Y(mai_mai_n515_));
  NOi32      m0487(.An(g), .Bn(f), .C(i), .Y(mai_mai_n516_));
  NO2        m0488(.A(mai_mai_n251_), .B(mai_mai_n47_), .Y(mai_mai_n517_));
  NA2        m0489(.A(mai_mai_n512_), .B(mai_mai_n509_), .Y(mai_mai_n518_));
  NA2        m0490(.A(mai_mai_n126_), .B(mai_mai_n34_), .Y(mai_mai_n519_));
  OAI220     m0491(.A0(mai_mai_n519_), .A1(m), .B0(mai_mai_n504_), .B1(mai_mai_n215_), .Y(mai_mai_n520_));
  NOi41      m0492(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n521_));
  NAi32      m0493(.An(e), .Bn(b), .C(c), .Y(mai_mai_n522_));
  OR2        m0494(.A(mai_mai_n522_), .B(mai_mai_n80_), .Y(mai_mai_n523_));
  AN2        m0495(.A(mai_mai_n310_), .B(mai_mai_n291_), .Y(mai_mai_n524_));
  NA2        m0496(.A(mai_mai_n524_), .B(mai_mai_n523_), .Y(mai_mai_n525_));
  OA210      m0497(.A0(mai_mai_n525_), .A1(mai_mai_n521_), .B0(mai_mai_n520_), .Y(mai_mai_n526_));
  OAI220     m0498(.A0(mai_mai_n368_), .A1(mai_mai_n367_), .B0(mai_mai_n500_), .B1(mai_mai_n499_), .Y(mai_mai_n527_));
  NAi31      m0499(.An(d), .B(c), .C(a), .Y(mai_mai_n528_));
  NO2        m0500(.A(mai_mai_n528_), .B(n), .Y(mai_mai_n529_));
  NA3        m0501(.A(mai_mai_n529_), .B(mai_mai_n527_), .C(e), .Y(mai_mai_n530_));
  NO3        m0502(.A(mai_mai_n59_), .B(mai_mai_n47_), .C(mai_mai_n197_), .Y(mai_mai_n531_));
  NO2        m0503(.A(mai_mai_n212_), .B(mai_mai_n100_), .Y(mai_mai_n532_));
  OAI210     m0504(.A0(mai_mai_n531_), .A1(mai_mai_n369_), .B0(mai_mai_n532_), .Y(mai_mai_n533_));
  NA2        m0505(.A(mai_mai_n533_), .B(mai_mai_n530_), .Y(mai_mai_n534_));
  NAi32      m0506(.An(d), .Bn(a), .C(b), .Y(mai_mai_n535_));
  AN3        m0507(.A(j), .B(h), .C(g), .Y(mai_mai_n536_));
  NO2        m0508(.A(mai_mai_n131_), .B(c), .Y(mai_mai_n537_));
  NA3        m0509(.A(f), .B(d), .C(b), .Y(mai_mai_n538_));
  NO2        m0510(.A(mai_mai_n534_), .B(mai_mai_n526_), .Y(mai_mai_n539_));
  AN2        m0511(.A(mai_mai_n539_), .B(mai_mai_n518_), .Y(mai_mai_n540_));
  INV        m0512(.A(k), .Y(mai_mai_n541_));
  NA3        m0513(.A(l), .B(mai_mai_n541_), .C(i), .Y(mai_mai_n542_));
  INV        m0514(.A(mai_mai_n542_), .Y(mai_mai_n543_));
  NA4        m0515(.A(mai_mai_n365_), .B(mai_mai_n386_), .C(mai_mai_n165_), .D(mai_mai_n103_), .Y(mai_mai_n544_));
  NAi32      m0516(.An(h), .Bn(f), .C(g), .Y(mai_mai_n545_));
  NAi41      m0517(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n546_));
  OAI210     m0518(.A0(mai_mai_n505_), .A1(n), .B0(mai_mai_n546_), .Y(mai_mai_n547_));
  NA2        m0519(.A(mai_mai_n547_), .B(m), .Y(mai_mai_n548_));
  NAi31      m0520(.An(h), .B(g), .C(f), .Y(mai_mai_n549_));
  OR3        m0521(.A(mai_mai_n549_), .B(mai_mai_n253_), .C(mai_mai_n47_), .Y(mai_mai_n550_));
  NA4        m0522(.A(mai_mai_n386_), .B(mai_mai_n110_), .C(mai_mai_n103_), .D(e), .Y(mai_mai_n551_));
  AN2        m0523(.A(mai_mai_n551_), .B(mai_mai_n550_), .Y(mai_mai_n552_));
  OA210      m0524(.A0(mai_mai_n548_), .A1(mai_mai_n545_), .B0(mai_mai_n552_), .Y(mai_mai_n553_));
  NA2        m0525(.A(mai_mai_n553_), .B(mai_mai_n544_), .Y(mai_mai_n554_));
  NAi31      m0526(.An(f), .B(h), .C(g), .Y(mai_mai_n555_));
  NO4        m0527(.A(mai_mai_n282_), .B(mai_mai_n555_), .C(mai_mai_n67_), .D(mai_mai_n69_), .Y(mai_mai_n556_));
  NOi41      m0528(.An(b), .B(mai_mai_n323_), .C(mai_mai_n64_), .D(mai_mai_n107_), .Y(mai_mai_n557_));
  OR2        m0529(.A(mai_mai_n557_), .B(mai_mai_n556_), .Y(mai_mai_n558_));
  NOi32      m0530(.An(d), .Bn(a), .C(e), .Y(mai_mai_n559_));
  NO2        m0531(.A(n), .B(c), .Y(mai_mai_n560_));
  NA3        m0532(.A(mai_mai_n560_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n561_));
  INV        m0533(.A(n), .Y(mai_mai_n562_));
  NOi32      m0534(.An(e), .Bn(a), .C(d), .Y(mai_mai_n563_));
  AOI210     m0535(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n563_), .Y(mai_mai_n564_));
  NO2        m0536(.A(mai_mai_n564_), .B(mai_mai_n519_), .Y(mai_mai_n565_));
  AOI210     m0537(.A0(mai_mai_n565_), .A1(mai_mai_n562_), .B0(mai_mai_n558_), .Y(mai_mai_n566_));
  OAI210     m0538(.A0(mai_mai_n232_), .A1(mai_mai_n83_), .B0(mai_mai_n566_), .Y(mai_mai_n567_));
  AOI210     m0539(.A0(mai_mai_n554_), .A1(mai_mai_n543_), .B0(mai_mai_n567_), .Y(mai_mai_n568_));
  NO3        m0540(.A(mai_mai_n289_), .B(mai_mai_n58_), .C(n), .Y(mai_mai_n569_));
  NA3        m0541(.A(mai_mai_n484_), .B(mai_mai_n155_), .C(mai_mai_n154_), .Y(mai_mai_n570_));
  NA2        m0542(.A(mai_mai_n432_), .B(mai_mai_n212_), .Y(mai_mai_n571_));
  OR2        m0543(.A(mai_mai_n571_), .B(mai_mai_n570_), .Y(mai_mai_n572_));
  NA2        m0544(.A(mai_mai_n70_), .B(mai_mai_n103_), .Y(mai_mai_n573_));
  NO2        m0545(.A(mai_mai_n573_), .B(mai_mai_n44_), .Y(mai_mai_n574_));
  AOI220     m0546(.A0(mai_mai_n574_), .A1(mai_mai_n509_), .B0(mai_mai_n572_), .B1(mai_mai_n569_), .Y(mai_mai_n575_));
  NO2        m0547(.A(mai_mai_n575_), .B(mai_mai_n83_), .Y(mai_mai_n576_));
  NOi32      m0548(.An(e), .Bn(c), .C(f), .Y(mai_mai_n577_));
  NOi21      m0549(.An(f), .B(g), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n578_), .B(mai_mai_n195_), .Y(mai_mai_n579_));
  AOI220     m0551(.A0(mai_mai_n579_), .A1(mai_mai_n362_), .B0(mai_mai_n577_), .B1(mai_mai_n159_), .Y(mai_mai_n580_));
  NA2        m0552(.A(mai_mai_n580_), .B(mai_mai_n162_), .Y(mai_mai_n581_));
  AOI210     m0553(.A0(mai_mai_n508_), .A1(mai_mai_n366_), .B0(mai_mai_n272_), .Y(mai_mai_n582_));
  NAi21      m0554(.An(k), .B(h), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n583_), .B(mai_mai_n242_), .Y(mai_mai_n584_));
  NOi31      m0556(.An(m), .B(n), .C(k), .Y(mai_mai_n585_));
  NA2        m0557(.A(j), .B(mai_mai_n585_), .Y(mai_mai_n586_));
  AOI210     m0558(.A0(mai_mai_n366_), .A1(mai_mai_n340_), .B0(mai_mai_n272_), .Y(mai_mai_n587_));
  NAi21      m0559(.An(mai_mai_n586_), .B(mai_mai_n587_), .Y(mai_mai_n588_));
  NO2        m0560(.A(mai_mai_n505_), .B(mai_mai_n47_), .Y(mai_mai_n589_));
  INV        m0561(.A(mai_mai_n588_), .Y(mai_mai_n590_));
  NA2        m0562(.A(mai_mai_n98_), .B(mai_mai_n36_), .Y(mai_mai_n591_));
  NO2        m0563(.A(k), .B(mai_mai_n197_), .Y(mai_mai_n592_));
  INV        m0564(.A(mai_mai_n331_), .Y(mai_mai_n593_));
  NO2        m0565(.A(mai_mai_n593_), .B(n), .Y(mai_mai_n594_));
  NAi31      m0566(.An(mai_mai_n591_), .B(mai_mai_n594_), .C(mai_mai_n592_), .Y(mai_mai_n595_));
  NO2        m0567(.A(mai_mai_n504_), .B(mai_mai_n160_), .Y(mai_mai_n596_));
  NA3        m0568(.A(mai_mai_n522_), .B(mai_mai_n248_), .C(mai_mai_n130_), .Y(mai_mai_n597_));
  NA2        m0569(.A(mai_mai_n481_), .B(mai_mai_n144_), .Y(mai_mai_n598_));
  NO3        m0570(.A(mai_mai_n363_), .B(mai_mai_n598_), .C(mai_mai_n83_), .Y(mai_mai_n599_));
  AOI210     m0571(.A0(mai_mai_n597_), .A1(mai_mai_n596_), .B0(mai_mai_n599_), .Y(mai_mai_n600_));
  AN3        m0572(.A(f), .B(d), .C(b), .Y(mai_mai_n601_));
  OAI210     m0573(.A0(mai_mai_n601_), .A1(mai_mai_n117_), .B0(n), .Y(mai_mai_n602_));
  NA3        m0574(.A(mai_mai_n481_), .B(mai_mai_n144_), .C(mai_mai_n197_), .Y(mai_mai_n603_));
  AOI210     m0575(.A0(mai_mai_n602_), .A1(mai_mai_n214_), .B0(mai_mai_n603_), .Y(mai_mai_n604_));
  NAi31      m0576(.An(m), .B(n), .C(k), .Y(mai_mai_n605_));
  OR2        m0577(.A(mai_mai_n122_), .B(mai_mai_n58_), .Y(mai_mai_n606_));
  OAI210     m0578(.A0(mai_mai_n606_), .A1(mai_mai_n605_), .B0(mai_mai_n234_), .Y(mai_mai_n607_));
  OAI210     m0579(.A0(mai_mai_n607_), .A1(mai_mai_n604_), .B0(j), .Y(mai_mai_n608_));
  NA3        m0580(.A(mai_mai_n608_), .B(mai_mai_n600_), .C(mai_mai_n595_), .Y(mai_mai_n609_));
  NO4        m0581(.A(mai_mai_n609_), .B(mai_mai_n590_), .C(mai_mai_n581_), .D(mai_mai_n576_), .Y(mai_mai_n610_));
  NA2        m0582(.A(mai_mai_n350_), .B(mai_mai_n147_), .Y(mai_mai_n611_));
  NAi31      m0583(.An(g), .B(h), .C(f), .Y(mai_mai_n612_));
  OR3        m0584(.A(mai_mai_n612_), .B(mai_mai_n253_), .C(n), .Y(mai_mai_n613_));
  OA210      m0585(.A0(mai_mai_n505_), .A1(n), .B0(mai_mai_n546_), .Y(mai_mai_n614_));
  NA3        m0586(.A(mai_mai_n384_), .B(mai_mai_n110_), .C(mai_mai_n80_), .Y(mai_mai_n615_));
  OAI210     m0587(.A0(mai_mai_n614_), .A1(mai_mai_n86_), .B0(mai_mai_n615_), .Y(mai_mai_n616_));
  NOi21      m0588(.An(mai_mai_n613_), .B(mai_mai_n616_), .Y(mai_mai_n617_));
  AOI210     m0589(.A0(mai_mai_n617_), .A1(mai_mai_n611_), .B0(mai_mai_n501_), .Y(mai_mai_n618_));
  NO3        m0590(.A(g), .B(mai_mai_n196_), .C(mai_mai_n54_), .Y(mai_mai_n619_));
  NO2        m0591(.A(mai_mai_n488_), .B(mai_mai_n83_), .Y(mai_mai_n620_));
  OAI210     m0592(.A0(mai_mai_n620_), .A1(mai_mai_n362_), .B0(mai_mai_n619_), .Y(mai_mai_n621_));
  AN2        m0593(.A(h), .B(f), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n622_), .B(mai_mai_n37_), .Y(mai_mai_n623_));
  AOI210     m0595(.A0(mai_mai_n535_), .A1(mai_mai_n396_), .B0(mai_mai_n47_), .Y(mai_mai_n624_));
  OAI220     m0596(.A0(mai_mai_n549_), .A1(mai_mai_n542_), .B0(mai_mai_n297_), .B1(mai_mai_n499_), .Y(mai_mai_n625_));
  NA2        m0597(.A(mai_mai_n625_), .B(mai_mai_n624_), .Y(mai_mai_n626_));
  NA2        m0598(.A(mai_mai_n626_), .B(mai_mai_n621_), .Y(mai_mai_n627_));
  NO2        m0599(.A(mai_mai_n236_), .B(f), .Y(mai_mai_n628_));
  NO2        m0600(.A(mai_mai_n578_), .B(mai_mai_n58_), .Y(mai_mai_n629_));
  NO3        m0601(.A(mai_mai_n629_), .B(mai_mai_n628_), .C(mai_mai_n34_), .Y(mai_mai_n630_));
  NA2        m0602(.A(mai_mai_n300_), .B(mai_mai_n126_), .Y(mai_mai_n631_));
  NA2        m0603(.A(mai_mai_n119_), .B(mai_mai_n47_), .Y(mai_mai_n632_));
  NA2        m0604(.A(mai_mai_n331_), .B(mai_mai_n103_), .Y(mai_mai_n633_));
  OA220      m0605(.A0(mai_mai_n633_), .A1(mai_mai_n519_), .B0(mai_mai_n330_), .B1(mai_mai_n101_), .Y(mai_mai_n634_));
  OAI210     m0606(.A0(mai_mai_n631_), .A1(mai_mai_n630_), .B0(mai_mai_n634_), .Y(mai_mai_n635_));
  NO3        m0607(.A(mai_mai_n373_), .B(mai_mai_n177_), .C(mai_mai_n176_), .Y(mai_mai_n636_));
  NA2        m0608(.A(mai_mai_n636_), .B(mai_mai_n212_), .Y(mai_mai_n637_));
  NA3        m0609(.A(mai_mai_n637_), .B(mai_mai_n238_), .C(j), .Y(mai_mai_n638_));
  NA2        m0610(.A(mai_mai_n435_), .B(mai_mai_n80_), .Y(mai_mai_n639_));
  NO4        m0611(.A(mai_mai_n501_), .B(mai_mai_n639_), .C(mai_mai_n118_), .D(mai_mai_n196_), .Y(mai_mai_n640_));
  INV        m0612(.A(mai_mai_n640_), .Y(mai_mai_n641_));
  NA4        m0613(.A(mai_mai_n641_), .B(mai_mai_n638_), .C(mai_mai_n487_), .D(mai_mai_n371_), .Y(mai_mai_n642_));
  NO4        m0614(.A(mai_mai_n642_), .B(mai_mai_n635_), .C(mai_mai_n627_), .D(mai_mai_n618_), .Y(mai_mai_n643_));
  NA4        m0615(.A(mai_mai_n643_), .B(mai_mai_n610_), .C(mai_mai_n568_), .D(mai_mai_n540_), .Y(mai08));
  NO2        m0616(.A(k), .B(h), .Y(mai_mai_n645_));
  AO210      m0617(.A0(mai_mai_n236_), .A1(mai_mai_n421_), .B0(mai_mai_n645_), .Y(mai_mai_n646_));
  NO2        m0618(.A(mai_mai_n646_), .B(mai_mai_n270_), .Y(mai_mai_n647_));
  NA2        m0619(.A(mai_mai_n577_), .B(mai_mai_n80_), .Y(mai_mai_n648_));
  NA2        m0620(.A(mai_mai_n648_), .B(mai_mai_n432_), .Y(mai_mai_n649_));
  AOI210     m0621(.A0(mai_mai_n649_), .A1(mai_mai_n647_), .B0(mai_mai_n463_), .Y(mai_mai_n650_));
  NA2        m0622(.A(mai_mai_n80_), .B(mai_mai_n100_), .Y(mai_mai_n651_));
  NO2        m0623(.A(mai_mai_n651_), .B(mai_mai_n55_), .Y(mai_mai_n652_));
  NO4        m0624(.A(mai_mai_n347_), .B(mai_mai_n102_), .C(j), .D(mai_mai_n197_), .Y(mai_mai_n653_));
  NA2        m0625(.A(mai_mai_n538_), .B(mai_mai_n214_), .Y(mai_mai_n654_));
  AOI220     m0626(.A0(mai_mai_n654_), .A1(mai_mai_n320_), .B0(mai_mai_n653_), .B1(mai_mai_n652_), .Y(mai_mai_n655_));
  AOI210     m0627(.A0(mai_mai_n538_), .A1(mai_mai_n140_), .B0(mai_mai_n80_), .Y(mai_mai_n656_));
  NA4        m0628(.A(mai_mai_n199_), .B(mai_mai_n126_), .C(mai_mai_n44_), .D(h), .Y(mai_mai_n657_));
  AN2        m0629(.A(l), .B(k), .Y(mai_mai_n658_));
  NA4        m0630(.A(mai_mai_n658_), .B(mai_mai_n98_), .C(mai_mai_n69_), .D(mai_mai_n197_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n657_), .B(mai_mai_n659_), .Y(mai_mai_n660_));
  NA2        m0632(.A(mai_mai_n660_), .B(mai_mai_n656_), .Y(mai_mai_n661_));
  NA3        m0633(.A(mai_mai_n661_), .B(mai_mai_n655_), .C(mai_mai_n650_), .Y(mai_mai_n662_));
  NO4        m0634(.A(mai_mai_n157_), .B(mai_mai_n361_), .C(mai_mai_n102_), .D(g), .Y(mai_mai_n663_));
  NO2        m0635(.A(mai_mai_n508_), .B(mai_mai_n35_), .Y(mai_mai_n664_));
  OAI210     m0636(.A0(mai_mai_n522_), .A1(mai_mai_n46_), .B0(mai_mai_n606_), .Y(mai_mai_n665_));
  NO2        m0637(.A(mai_mai_n455_), .B(mai_mai_n119_), .Y(mai_mai_n666_));
  AOI210     m0638(.A0(mai_mai_n666_), .A1(mai_mai_n665_), .B0(mai_mai_n664_), .Y(mai_mai_n667_));
  INV        m0639(.A(mai_mai_n659_), .Y(mai_mai_n668_));
  NA2        m0640(.A(mai_mai_n646_), .B(mai_mai_n123_), .Y(mai_mai_n669_));
  AOI220     m0641(.A0(mai_mai_n669_), .A1(mai_mai_n372_), .B0(mai_mai_n668_), .B1(mai_mai_n72_), .Y(mai_mai_n670_));
  NA2        m0642(.A(mai_mai_n667_), .B(mai_mai_n670_), .Y(mai_mai_n671_));
  NA2        m0643(.A(mai_mai_n331_), .B(mai_mai_n43_), .Y(mai_mai_n672_));
  NA3        m0644(.A(mai_mai_n637_), .B(mai_mai_n305_), .C(mai_mai_n353_), .Y(mai_mai_n673_));
  NA2        m0645(.A(mai_mai_n658_), .B(mai_mai_n202_), .Y(mai_mai_n674_));
  NO2        m0646(.A(mai_mai_n674_), .B(mai_mai_n299_), .Y(mai_mai_n675_));
  AOI210     m0647(.A0(mai_mai_n675_), .A1(mai_mai_n628_), .B0(mai_mai_n462_), .Y(mai_mai_n676_));
  NA3        m0648(.A(m), .B(l), .C(k), .Y(mai_mai_n677_));
  AOI210     m0649(.A0(mai_mai_n615_), .A1(mai_mai_n613_), .B0(mai_mai_n677_), .Y(mai_mai_n678_));
  NO2        m0650(.A(mai_mai_n507_), .B(mai_mai_n249_), .Y(mai_mai_n679_));
  NOi21      m0651(.An(mai_mai_n679_), .B(mai_mai_n503_), .Y(mai_mai_n680_));
  NA4        m0652(.A(mai_mai_n103_), .B(l), .C(k), .D(mai_mai_n83_), .Y(mai_mai_n681_));
  NA3        m0653(.A(mai_mai_n110_), .B(mai_mai_n380_), .C(i), .Y(mai_mai_n682_));
  NO2        m0654(.A(mai_mai_n682_), .B(mai_mai_n681_), .Y(mai_mai_n683_));
  NO3        m0655(.A(mai_mai_n683_), .B(mai_mai_n680_), .C(mai_mai_n678_), .Y(mai_mai_n684_));
  NA4        m0656(.A(mai_mai_n684_), .B(mai_mai_n676_), .C(mai_mai_n673_), .D(mai_mai_n672_), .Y(mai_mai_n685_));
  NO4        m0657(.A(mai_mai_n685_), .B(mai_mai_n671_), .C(mai_mai_n493_), .D(mai_mai_n662_), .Y(mai_mai_n686_));
  NA2        m0658(.A(mai_mai_n579_), .B(mai_mai_n362_), .Y(mai_mai_n687_));
  NOi31      m0659(.An(g), .B(h), .C(f), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n589_), .B(mai_mai_n688_), .Y(mai_mai_n689_));
  AO210      m0661(.A0(mai_mai_n689_), .A1(mai_mai_n550_), .B0(mai_mai_n510_), .Y(mai_mai_n690_));
  NO3        m0662(.A(mai_mai_n366_), .B(mai_mai_n499_), .C(h), .Y(mai_mai_n691_));
  AOI210     m0663(.A0(mai_mai_n691_), .A1(mai_mai_n103_), .B0(mai_mai_n474_), .Y(mai_mai_n692_));
  NA4        m0664(.A(mai_mai_n692_), .B(mai_mai_n690_), .C(mai_mai_n687_), .D(mai_mai_n235_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n658_), .B(mai_mai_n69_), .Y(mai_mai_n694_));
  NO4        m0666(.A(mai_mai_n636_), .B(mai_mai_n157_), .C(n), .D(i), .Y(mai_mai_n695_));
  NOi21      m0667(.An(h), .B(j), .Y(mai_mai_n696_));
  NA2        m0668(.A(mai_mai_n696_), .B(f), .Y(mai_mai_n697_));
  NO2        m0669(.A(mai_mai_n697_), .B(mai_mai_n229_), .Y(mai_mai_n698_));
  NO2        m0670(.A(mai_mai_n698_), .B(mai_mai_n695_), .Y(mai_mai_n699_));
  OAI220     m0671(.A0(mai_mai_n699_), .A1(mai_mai_n694_), .B0(mai_mai_n552_), .B1(mai_mai_n59_), .Y(mai_mai_n700_));
  AOI210     m0672(.A0(mai_mai_n693_), .A1(l), .B0(mai_mai_n700_), .Y(mai_mai_n701_));
  NO2        m0673(.A(j), .B(i), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n702_), .B(mai_mai_n33_), .Y(mai_mai_n703_));
  NA2        m0675(.A(mai_mai_n389_), .B(mai_mai_n110_), .Y(mai_mai_n704_));
  OR2        m0676(.A(mai_mai_n704_), .B(mai_mai_n703_), .Y(mai_mai_n705_));
  NO3        m0677(.A(mai_mai_n136_), .B(mai_mai_n47_), .C(mai_mai_n100_), .Y(mai_mai_n706_));
  NO3        m0678(.A(mai_mai_n514_), .B(mai_mai_n134_), .C(mai_mai_n69_), .Y(mai_mai_n707_));
  NO3        m0679(.A(mai_mai_n455_), .B(mai_mai_n408_), .C(j), .Y(mai_mai_n708_));
  OAI210     m0680(.A0(mai_mai_n707_), .A1(mai_mai_n706_), .B0(mai_mai_n708_), .Y(mai_mai_n709_));
  OAI210     m0681(.A0(mai_mai_n689_), .A1(mai_mai_n59_), .B0(mai_mai_n709_), .Y(mai_mai_n710_));
  NA2        m0682(.A(k), .B(j), .Y(mai_mai_n711_));
  NO3        m0683(.A(mai_mai_n270_), .B(mai_mai_n711_), .C(mai_mai_n40_), .Y(mai_mai_n712_));
  AOI210     m0684(.A0(mai_mai_n502_), .A1(n), .B0(mai_mai_n521_), .Y(mai_mai_n713_));
  NA2        m0685(.A(mai_mai_n713_), .B(mai_mai_n524_), .Y(mai_mai_n714_));
  AN3        m0686(.A(mai_mai_n714_), .B(mai_mai_n712_), .C(mai_mai_n92_), .Y(mai_mai_n715_));
  NO3        m0687(.A(mai_mai_n157_), .B(mai_mai_n361_), .C(mai_mai_n102_), .Y(mai_mai_n716_));
  AOI220     m0688(.A0(mai_mai_n716_), .A1(mai_mai_n230_), .B0(mai_mai_n571_), .B1(mai_mai_n279_), .Y(mai_mai_n717_));
  INV        m0689(.A(mai_mai_n717_), .Y(mai_mai_n718_));
  NO2        m0690(.A(mai_mai_n270_), .B(mai_mai_n123_), .Y(mai_mai_n719_));
  NA2        m0691(.A(mai_mai_n719_), .B(mai_mai_n579_), .Y(mai_mai_n720_));
  NO2        m0692(.A(mai_mai_n677_), .B(mai_mai_n86_), .Y(mai_mai_n721_));
  NA2        m0693(.A(mai_mai_n721_), .B(mai_mai_n547_), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n549_), .B(mai_mai_n107_), .Y(mai_mai_n723_));
  OAI210     m0695(.A0(mai_mai_n723_), .A1(mai_mai_n708_), .B0(mai_mai_n624_), .Y(mai_mai_n724_));
  NA3        m0696(.A(mai_mai_n724_), .B(mai_mai_n722_), .C(mai_mai_n720_), .Y(mai_mai_n725_));
  OR4        m0697(.A(mai_mai_n725_), .B(mai_mai_n718_), .C(mai_mai_n715_), .D(mai_mai_n710_), .Y(mai_mai_n726_));
  NA3        m0698(.A(mai_mai_n713_), .B(mai_mai_n524_), .C(mai_mai_n523_), .Y(mai_mai_n727_));
  NA4        m0699(.A(mai_mai_n727_), .B(mai_mai_n199_), .C(mai_mai_n421_), .D(mai_mai_n34_), .Y(mai_mai_n728_));
  OAI220     m0700(.A0(mai_mai_n657_), .A1(mai_mai_n648_), .B0(mai_mai_n303_), .B1(mai_mai_n38_), .Y(mai_mai_n729_));
  INV        m0701(.A(mai_mai_n729_), .Y(mai_mai_n730_));
  NA3        m0702(.A(mai_mai_n516_), .B(mai_mai_n263_), .C(h), .Y(mai_mai_n731_));
  NOi21      m0703(.An(mai_mai_n624_), .B(mai_mai_n731_), .Y(mai_mai_n732_));
  NO2        m0704(.A(mai_mai_n87_), .B(mai_mai_n46_), .Y(mai_mai_n733_));
  NA2        m0705(.A(mai_mai_n733_), .B(mai_mai_n594_), .Y(mai_mai_n734_));
  NAi41      m0706(.An(mai_mai_n732_), .B(mai_mai_n734_), .C(mai_mai_n730_), .D(mai_mai_n728_), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n721_), .B(mai_mai_n220_), .Y(mai_mai_n736_));
  INV        m0708(.A(mai_mai_n307_), .Y(mai_mai_n737_));
  OAI210     m0709(.A0(mai_mai_n677_), .A1(mai_mai_n612_), .B0(mai_mai_n492_), .Y(mai_mai_n738_));
  NA3        m0710(.A(mai_mai_n233_), .B(mai_mai_n57_), .C(b), .Y(mai_mai_n739_));
  AOI220     m0711(.A0(mai_mai_n560_), .A1(mai_mai_n29_), .B0(mai_mai_n435_), .B1(mai_mai_n80_), .Y(mai_mai_n740_));
  NA2        m0712(.A(mai_mai_n740_), .B(mai_mai_n739_), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n731_), .B(mai_mai_n461_), .Y(mai_mai_n742_));
  AOI210     m0714(.A0(mai_mai_n741_), .A1(mai_mai_n738_), .B0(mai_mai_n742_), .Y(mai_mai_n743_));
  NA3        m0715(.A(mai_mai_n743_), .B(mai_mai_n737_), .C(mai_mai_n736_), .Y(mai_mai_n744_));
  NOi41      m0716(.An(mai_mai_n705_), .B(mai_mai_n744_), .C(mai_mai_n735_), .D(mai_mai_n726_), .Y(mai_mai_n745_));
  OR2        m0717(.A(mai_mai_n657_), .B(mai_mai_n214_), .Y(mai_mai_n746_));
  NO3        m0718(.A(mai_mai_n313_), .B(mai_mai_n272_), .C(mai_mai_n102_), .Y(mai_mai_n747_));
  NA2        m0719(.A(mai_mai_n747_), .B(mai_mai_n714_), .Y(mai_mai_n748_));
  NA2        m0720(.A(mai_mai_n45_), .B(mai_mai_n54_), .Y(mai_mai_n749_));
  NO3        m0721(.A(mai_mai_n749_), .B(mai_mai_n703_), .C(mai_mai_n253_), .Y(mai_mai_n750_));
  NO3        m0722(.A(mai_mai_n499_), .B(mai_mai_n88_), .C(h), .Y(mai_mai_n751_));
  AOI210     m0723(.A0(mai_mai_n751_), .A1(mai_mai_n652_), .B0(mai_mai_n750_), .Y(mai_mai_n752_));
  NA4        m0724(.A(mai_mai_n752_), .B(mai_mai_n748_), .C(mai_mai_n746_), .D(mai_mai_n374_), .Y(mai_mai_n753_));
  NOi31      m0725(.An(b), .B(d), .C(a), .Y(mai_mai_n754_));
  NO2        m0726(.A(mai_mai_n754_), .B(mai_mai_n559_), .Y(mai_mai_n755_));
  NO2        m0727(.A(mai_mai_n755_), .B(n), .Y(mai_mai_n756_));
  NO2        m0728(.A(mai_mai_n522_), .B(mai_mai_n80_), .Y(mai_mai_n757_));
  NA2        m0729(.A(mai_mai_n747_), .B(mai_mai_n757_), .Y(mai_mai_n758_));
  OAI210     m0730(.A0(mai_mai_n657_), .A1(mai_mai_n363_), .B0(mai_mai_n758_), .Y(mai_mai_n759_));
  NO2        m0731(.A(mai_mai_n636_), .B(n), .Y(mai_mai_n760_));
  BUFFER     m0732(.A(mai_mai_n719_), .Y(mai_mai_n761_));
  AOI220     m0733(.A0(mai_mai_n761_), .A1(mai_mai_n619_), .B0(mai_mai_n760_), .B1(mai_mai_n647_), .Y(mai_mai_n762_));
  NA2        m0734(.A(mai_mai_n110_), .B(mai_mai_n80_), .Y(mai_mai_n763_));
  AOI210     m0735(.A0(mai_mai_n393_), .A1(mai_mai_n385_), .B0(mai_mai_n763_), .Y(mai_mai_n764_));
  NA2        m0736(.A(mai_mai_n675_), .B(mai_mai_n34_), .Y(mai_mai_n765_));
  NAi21      m0737(.An(mai_mai_n681_), .B(mai_mai_n404_), .Y(mai_mai_n766_));
  NO2        m0738(.A(mai_mai_n249_), .B(i), .Y(mai_mai_n767_));
  NA2        m0739(.A(mai_mai_n663_), .B(mai_mai_n321_), .Y(mai_mai_n768_));
  AN2        m0740(.A(mai_mai_n768_), .B(mai_mai_n766_), .Y(mai_mai_n769_));
  NAi41      m0741(.An(mai_mai_n764_), .B(mai_mai_n769_), .C(mai_mai_n765_), .D(mai_mai_n762_), .Y(mai_mai_n770_));
  NO3        m0742(.A(mai_mai_n770_), .B(mai_mai_n759_), .C(mai_mai_n753_), .Y(mai_mai_n771_));
  NA4        m0743(.A(mai_mai_n771_), .B(mai_mai_n745_), .C(mai_mai_n701_), .D(mai_mai_n686_), .Y(mai09));
  INV        m0744(.A(mai_mai_n111_), .Y(mai_mai_n773_));
  NA2        m0745(.A(f), .B(e), .Y(mai_mai_n774_));
  NO2        m0746(.A(mai_mai_n207_), .B(mai_mai_n102_), .Y(mai_mai_n775_));
  NA2        m0747(.A(mai_mai_n775_), .B(g), .Y(mai_mai_n776_));
  AOI210     m0748(.A0(mai_mai_n70_), .A1(g), .B0(mai_mai_n441_), .Y(mai_mai_n777_));
  AOI210     m0749(.A0(mai_mai_n777_), .A1(mai_mai_n776_), .B0(mai_mai_n774_), .Y(mai_mai_n778_));
  NA2        m0750(.A(mai_mai_n414_), .B(e), .Y(mai_mai_n779_));
  NO2        m0751(.A(mai_mai_n779_), .B(mai_mai_n484_), .Y(mai_mai_n780_));
  AOI210     m0752(.A0(mai_mai_n778_), .A1(mai_mai_n773_), .B0(mai_mai_n780_), .Y(mai_mai_n781_));
  NO2        m0753(.A(mai_mai_n187_), .B(mai_mai_n196_), .Y(mai_mai_n782_));
  NA3        m0754(.A(m), .B(l), .C(i), .Y(mai_mai_n783_));
  OAI220     m0755(.A0(mai_mai_n549_), .A1(mai_mai_n783_), .B0(mai_mai_n323_), .B1(mai_mai_n500_), .Y(mai_mai_n784_));
  NA4        m0756(.A(mai_mai_n84_), .B(mai_mai_n83_), .C(g), .D(f), .Y(mai_mai_n785_));
  NAi31      m0757(.An(mai_mai_n784_), .B(mai_mai_n785_), .C(mai_mai_n409_), .Y(mai_mai_n786_));
  OR2        m0758(.A(mai_mai_n786_), .B(mai_mai_n782_), .Y(mai_mai_n787_));
  INV        m0759(.A(mai_mai_n492_), .Y(mai_mai_n788_));
  OA210      m0760(.A0(mai_mai_n788_), .A1(mai_mai_n787_), .B0(mai_mai_n756_), .Y(mai_mai_n789_));
  INV        m0761(.A(mai_mai_n310_), .Y(mai_mai_n790_));
  NO2        m0762(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n791_));
  NOi31      m0763(.An(k), .B(m), .C(l), .Y(mai_mai_n792_));
  NO2        m0764(.A(mai_mai_n312_), .B(mai_mai_n792_), .Y(mai_mai_n793_));
  AOI210     m0765(.A0(mai_mai_n793_), .A1(mai_mai_n791_), .B0(mai_mai_n555_), .Y(mai_mai_n794_));
  INV        m0766(.A(mai_mai_n303_), .Y(mai_mai_n795_));
  NA2        m0767(.A(mai_mai_n794_), .B(mai_mai_n790_), .Y(mai_mai_n796_));
  NA3        m0768(.A(mai_mai_n104_), .B(mai_mai_n174_), .C(mai_mai_n31_), .Y(mai_mai_n797_));
  NA4        m0769(.A(mai_mai_n797_), .B(mai_mai_n796_), .C(mai_mai_n580_), .D(mai_mai_n78_), .Y(mai_mai_n798_));
  NO2        m0770(.A(mai_mai_n545_), .B(mai_mai_n470_), .Y(mai_mai_n799_));
  NA2        m0771(.A(mai_mai_n799_), .B(mai_mai_n174_), .Y(mai_mai_n800_));
  NOi21      m0772(.An(f), .B(d), .Y(mai_mai_n801_));
  NA2        m0773(.A(mai_mai_n801_), .B(m), .Y(mai_mai_n802_));
  NO2        m0774(.A(mai_mai_n802_), .B(mai_mai_n50_), .Y(mai_mai_n803_));
  NOi32      m0775(.An(g), .Bn(f), .C(d), .Y(mai_mai_n804_));
  NA4        m0776(.A(mai_mai_n804_), .B(mai_mai_n560_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n805_));
  NOi21      m0777(.An(mai_mai_n283_), .B(mai_mai_n805_), .Y(mai_mai_n806_));
  AOI210     m0778(.A0(mai_mai_n803_), .A1(mai_mai_n515_), .B0(mai_mai_n806_), .Y(mai_mai_n807_));
  AN2        m0779(.A(f), .B(d), .Y(mai_mai_n808_));
  NA3        m0780(.A(mai_mai_n446_), .B(mai_mai_n808_), .C(mai_mai_n80_), .Y(mai_mai_n809_));
  NO3        m0781(.A(mai_mai_n809_), .B(mai_mai_n69_), .C(mai_mai_n197_), .Y(mai_mai_n810_));
  NO2        m0782(.A(k), .B(mai_mai_n54_), .Y(mai_mai_n811_));
  NAi31      m0783(.An(mai_mai_n460_), .B(mai_mai_n807_), .C(mai_mai_n800_), .Y(mai_mai_n812_));
  NO4        m0784(.A(mai_mai_n578_), .B(mai_mai_n119_), .C(mai_mai_n299_), .D(mai_mai_n137_), .Y(mai_mai_n813_));
  NO2        m0785(.A(mai_mai_n605_), .B(mai_mai_n299_), .Y(mai_mai_n814_));
  AN2        m0786(.A(mai_mai_n814_), .B(mai_mai_n628_), .Y(mai_mai_n815_));
  NO3        m0787(.A(mai_mai_n815_), .B(mai_mai_n813_), .C(mai_mai_n216_), .Y(mai_mai_n816_));
  NA2        m0788(.A(mai_mai_n559_), .B(mai_mai_n80_), .Y(mai_mai_n817_));
  NA3        m0789(.A(mai_mai_n144_), .B(mai_mai_n98_), .C(g), .Y(mai_mai_n818_));
  OAI220     m0790(.A0(mai_mai_n809_), .A1(mai_mai_n398_), .B0(mai_mai_n310_), .B1(mai_mai_n818_), .Y(mai_mai_n819_));
  NOi31      m0791(.An(mai_mai_n205_), .B(mai_mai_n819_), .C(mai_mai_n277_), .Y(mai_mai_n820_));
  NA2        m0792(.A(c), .B(mai_mai_n106_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n821_), .B(mai_mai_n378_), .Y(mai_mai_n822_));
  NA3        m0794(.A(mai_mai_n822_), .B(mai_mai_n483_), .C(f), .Y(mai_mai_n823_));
  OR2        m0795(.A(mai_mai_n612_), .B(mai_mai_n511_), .Y(mai_mai_n824_));
  INV        m0796(.A(mai_mai_n824_), .Y(mai_mai_n825_));
  NA2        m0797(.A(mai_mai_n755_), .B(mai_mai_n101_), .Y(mai_mai_n826_));
  NA2        m0798(.A(mai_mai_n826_), .B(mai_mai_n825_), .Y(mai_mai_n827_));
  NA4        m0799(.A(mai_mai_n827_), .B(mai_mai_n823_), .C(mai_mai_n820_), .D(mai_mai_n816_), .Y(mai_mai_n828_));
  NO4        m0800(.A(mai_mai_n828_), .B(mai_mai_n812_), .C(mai_mai_n798_), .D(mai_mai_n789_), .Y(mai_mai_n829_));
  OR2        m0801(.A(mai_mai_n809_), .B(mai_mai_n69_), .Y(mai_mai_n830_));
  NA2        m0802(.A(mai_mai_n102_), .B(j), .Y(mai_mai_n831_));
  NA2        m0803(.A(mai_mai_n775_), .B(g), .Y(mai_mai_n832_));
  AOI210     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n264_), .B0(mai_mai_n830_), .Y(mai_mai_n833_));
  NO2        m0805(.A(mai_mai_n303_), .B(mai_mai_n785_), .Y(mai_mai_n834_));
  NO2        m0806(.A(mai_mai_n212_), .B(mai_mai_n206_), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n835_), .B(mai_mai_n209_), .Y(mai_mai_n836_));
  NO2        m0808(.A(mai_mai_n398_), .B(mai_mai_n774_), .Y(mai_mai_n837_));
  NA2        m0809(.A(mai_mai_n837_), .B(mai_mai_n529_), .Y(mai_mai_n838_));
  NA2        m0810(.A(mai_mai_n838_), .B(mai_mai_n836_), .Y(mai_mai_n839_));
  NA2        m0811(.A(e), .B(d), .Y(mai_mai_n840_));
  OAI220     m0812(.A0(mai_mai_n840_), .A1(c), .B0(mai_mai_n294_), .B1(d), .Y(mai_mai_n841_));
  NA3        m0813(.A(mai_mai_n841_), .B(mai_mai_n425_), .C(mai_mai_n481_), .Y(mai_mai_n842_));
  AOI210     m0814(.A0(mai_mai_n488_), .A1(mai_mai_n164_), .B0(mai_mai_n212_), .Y(mai_mai_n843_));
  INV        m0815(.A(mai_mai_n843_), .Y(mai_mai_n844_));
  NA2        m0816(.A(mai_mai_n810_), .B(j), .Y(mai_mai_n845_));
  NA3        m0817(.A(mai_mai_n150_), .B(mai_mai_n81_), .C(mai_mai_n34_), .Y(mai_mai_n846_));
  NA4        m0818(.A(mai_mai_n846_), .B(mai_mai_n845_), .C(mai_mai_n844_), .D(mai_mai_n842_), .Y(mai_mai_n847_));
  NO4        m0819(.A(mai_mai_n847_), .B(mai_mai_n839_), .C(mai_mai_n834_), .D(mai_mai_n833_), .Y(mai_mai_n848_));
  NA2        m0820(.A(mai_mai_n790_), .B(mai_mai_n31_), .Y(mai_mai_n849_));
  AO210      m0821(.A0(mai_mai_n849_), .A1(mai_mai_n648_), .B0(mai_mai_n200_), .Y(mai_mai_n850_));
  OAI220     m0822(.A0(mai_mai_n578_), .A1(mai_mai_n58_), .B0(mai_mai_n272_), .B1(j), .Y(mai_mai_n851_));
  AOI220     m0823(.A0(mai_mai_n851_), .A1(mai_mai_n814_), .B0(mai_mai_n569_), .B1(mai_mai_n577_), .Y(mai_mai_n852_));
  OAI210     m0824(.A0(mai_mai_n779_), .A1(mai_mai_n154_), .B0(mai_mai_n852_), .Y(mai_mai_n853_));
  NO2        m0825(.A(mai_mai_n1428_), .B(mai_mai_n805_), .Y(mai_mai_n854_));
  AO210      m0826(.A0(mai_mai_n795_), .A1(mai_mai_n784_), .B0(mai_mai_n854_), .Y(mai_mai_n855_));
  NOi31      m0827(.An(mai_mai_n515_), .B(mai_mai_n802_), .C(mai_mai_n264_), .Y(mai_mai_n856_));
  NO3        m0828(.A(mai_mai_n856_), .B(mai_mai_n855_), .C(mai_mai_n853_), .Y(mai_mai_n857_));
  AO220      m0829(.A0(mai_mai_n425_), .A1(mai_mai_n696_), .B0(mai_mai_n159_), .B1(f), .Y(mai_mai_n858_));
  OAI210     m0830(.A0(mai_mai_n858_), .A1(mai_mai_n428_), .B0(mai_mai_n841_), .Y(mai_mai_n859_));
  NO2        m0831(.A(mai_mai_n408_), .B(mai_mai_n66_), .Y(mai_mai_n860_));
  OAI210     m0832(.A0(mai_mai_n788_), .A1(mai_mai_n860_), .B0(mai_mai_n652_), .Y(mai_mai_n861_));
  AN4        m0833(.A(mai_mai_n861_), .B(mai_mai_n859_), .C(mai_mai_n857_), .D(mai_mai_n850_), .Y(mai_mai_n862_));
  NA4        m0834(.A(mai_mai_n862_), .B(mai_mai_n848_), .C(mai_mai_n829_), .D(mai_mai_n781_), .Y(mai12));
  NO2        m0835(.A(mai_mai_n423_), .B(c), .Y(mai_mai_n864_));
  NO4        m0836(.A(mai_mai_n413_), .B(mai_mai_n236_), .C(mai_mai_n541_), .D(mai_mai_n197_), .Y(mai_mai_n865_));
  NA2        m0837(.A(mai_mai_n865_), .B(mai_mai_n864_), .Y(mai_mai_n866_));
  NA2        m0838(.A(mai_mai_n515_), .B(mai_mai_n860_), .Y(mai_mai_n867_));
  NO2        m0839(.A(mai_mai_n423_), .B(mai_mai_n106_), .Y(mai_mai_n868_));
  NO2        m0840(.A(mai_mai_n791_), .B(mai_mai_n323_), .Y(mai_mai_n869_));
  NO2        m0841(.A(mai_mai_n612_), .B(mai_mai_n347_), .Y(mai_mai_n870_));
  AOI220     m0842(.A0(mai_mai_n870_), .A1(mai_mai_n513_), .B0(mai_mai_n869_), .B1(mai_mai_n868_), .Y(mai_mai_n871_));
  NA4        m0843(.A(mai_mai_n871_), .B(mai_mai_n867_), .C(mai_mai_n866_), .D(mai_mai_n412_), .Y(mai_mai_n872_));
  AOI210     m0844(.A0(mai_mai_n215_), .A1(mai_mai_n309_), .B0(mai_mai_n185_), .Y(mai_mai_n873_));
  OR2        m0845(.A(mai_mai_n873_), .B(mai_mai_n865_), .Y(mai_mai_n874_));
  AOI210     m0846(.A0(mai_mai_n306_), .A1(mai_mai_n359_), .B0(mai_mai_n197_), .Y(mai_mai_n875_));
  OAI210     m0847(.A0(mai_mai_n875_), .A1(mai_mai_n874_), .B0(mai_mai_n373_), .Y(mai_mai_n876_));
  NO2        m0848(.A(mai_mai_n549_), .B(mai_mai_n783_), .Y(mai_mai_n877_));
  NO2        m0849(.A(mai_mai_n136_), .B(mai_mai_n219_), .Y(mai_mai_n878_));
  NA3        m0850(.A(mai_mai_n878_), .B(mai_mai_n222_), .C(i), .Y(mai_mai_n879_));
  NA2        m0851(.A(mai_mai_n879_), .B(mai_mai_n876_), .Y(mai_mai_n880_));
  NO3        m0852(.A(mai_mai_n119_), .B(mai_mai_n137_), .C(mai_mai_n197_), .Y(mai_mai_n881_));
  NA2        m0853(.A(mai_mai_n881_), .B(mai_mai_n502_), .Y(mai_mai_n882_));
  NA4        m0854(.A(mai_mai_n414_), .B(mai_mai_n406_), .C(mai_mai_n165_), .D(g), .Y(mai_mai_n883_));
  NA2        m0855(.A(mai_mai_n883_), .B(mai_mai_n882_), .Y(mai_mai_n884_));
  NO3        m0856(.A(mai_mai_n617_), .B(mai_mai_n87_), .C(mai_mai_n44_), .Y(mai_mai_n885_));
  NO4        m0857(.A(mai_mai_n885_), .B(mai_mai_n884_), .C(mai_mai_n880_), .D(mai_mai_n872_), .Y(mai_mai_n886_));
  NO2        m0858(.A(mai_mai_n337_), .B(mai_mai_n336_), .Y(mai_mai_n887_));
  INV        m0859(.A(mai_mai_n546_), .Y(mai_mai_n888_));
  NA2        m0860(.A(mai_mai_n522_), .B(mai_mai_n130_), .Y(mai_mai_n889_));
  NOi21      m0861(.An(mai_mai_n34_), .B(mai_mai_n605_), .Y(mai_mai_n890_));
  AOI220     m0862(.A0(mai_mai_n890_), .A1(mai_mai_n889_), .B0(mai_mai_n888_), .B1(mai_mai_n887_), .Y(mai_mai_n891_));
  OAI210     m0863(.A0(mai_mai_n234_), .A1(mai_mai_n44_), .B0(mai_mai_n891_), .Y(mai_mai_n892_));
  NA2        m0864(.A(mai_mai_n404_), .B(mai_mai_n243_), .Y(mai_mai_n893_));
  NO3        m0865(.A(mai_mai_n763_), .B(mai_mai_n85_), .C(mai_mai_n378_), .Y(mai_mai_n894_));
  NAi31      m0866(.An(mai_mai_n894_), .B(mai_mai_n893_), .C(mai_mai_n293_), .Y(mai_mai_n895_));
  NO2        m0867(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n896_));
  NO2        m0868(.A(mai_mai_n477_), .B(mai_mai_n272_), .Y(mai_mai_n897_));
  INV        m0869(.A(mai_mai_n897_), .Y(mai_mai_n898_));
  NO2        m0870(.A(mai_mai_n898_), .B(mai_mai_n130_), .Y(mai_mai_n899_));
  NA2        m0871(.A(mai_mai_n585_), .B(mai_mai_n332_), .Y(mai_mai_n900_));
  INV        m0872(.A(mai_mai_n334_), .Y(mai_mai_n901_));
  NO4        m0873(.A(mai_mai_n901_), .B(mai_mai_n899_), .C(mai_mai_n895_), .D(mai_mai_n892_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n319_), .B(g), .Y(mai_mai_n903_));
  NA2        m0875(.A(mai_mai_n147_), .B(i), .Y(mai_mai_n904_));
  NO2        m0876(.A(mai_mai_n904_), .B(mai_mai_n87_), .Y(mai_mai_n905_));
  AOI210     m0877(.A0(mai_mai_n387_), .A1(mai_mai_n37_), .B0(mai_mai_n905_), .Y(mai_mai_n906_));
  NO2        m0878(.A(mai_mai_n130_), .B(mai_mai_n80_), .Y(mai_mai_n907_));
  OR2        m0879(.A(mai_mai_n907_), .B(mai_mai_n521_), .Y(mai_mai_n908_));
  NA2        m0880(.A(mai_mai_n522_), .B(mai_mai_n351_), .Y(mai_mai_n909_));
  AOI210     m0881(.A0(mai_mai_n909_), .A1(n), .B0(mai_mai_n908_), .Y(mai_mai_n910_));
  OAI220     m0882(.A0(mai_mai_n910_), .A1(mai_mai_n903_), .B0(mai_mai_n906_), .B1(mai_mai_n303_), .Y(mai_mai_n911_));
  NA3        m0883(.A(mai_mai_n296_), .B(mai_mai_n108_), .C(g), .Y(mai_mai_n912_));
  AOI210     m0884(.A0(mai_mai_n623_), .A1(mai_mai_n912_), .B0(m), .Y(mai_mai_n913_));
  OAI210     m0885(.A0(mai_mai_n913_), .A1(mai_mai_n869_), .B0(mai_mai_n295_), .Y(mai_mai_n914_));
  NA2        m0886(.A(mai_mai_n639_), .B(mai_mai_n817_), .Y(mai_mai_n915_));
  NA2        m0887(.A(mai_mai_n785_), .B(mai_mai_n409_), .Y(mai_mai_n916_));
  NA2        m0888(.A(mai_mai_n916_), .B(mai_mai_n915_), .Y(mai_mai_n917_));
  NA2        m0889(.A(mai_mai_n917_), .B(mai_mai_n914_), .Y(mai_mai_n918_));
  NA2        m0890(.A(mai_mai_n616_), .B(mai_mai_n84_), .Y(mai_mai_n919_));
  NO2        m0891(.A(mai_mai_n431_), .B(mai_mai_n197_), .Y(mai_mai_n920_));
  NA2        m0892(.A(mai_mai_n920_), .B(mai_mai_n352_), .Y(mai_mai_n921_));
  NA2        m0893(.A(mai_mai_n921_), .B(mai_mai_n919_), .Y(mai_mai_n922_));
  OAI210     m0894(.A0(mai_mai_n916_), .A1(mai_mai_n877_), .B0(mai_mai_n513_), .Y(mai_mai_n923_));
  AOI210     m0895(.A0(mai_mai_n388_), .A1(mai_mai_n381_), .B0(mai_mai_n763_), .Y(mai_mai_n924_));
  OAI210     m0896(.A0(mai_mai_n337_), .A1(mai_mai_n336_), .B0(mai_mai_n99_), .Y(mai_mai_n925_));
  AOI210     m0897(.A0(mai_mai_n925_), .A1(mai_mai_n506_), .B0(mai_mai_n924_), .Y(mai_mai_n926_));
  NA2        m0898(.A(mai_mai_n913_), .B(mai_mai_n868_), .Y(mai_mai_n927_));
  NO3        m0899(.A(mai_mai_n831_), .B(mai_mai_n47_), .C(mai_mai_n44_), .Y(mai_mai_n928_));
  AOI220     m0900(.A0(mai_mai_n928_), .A1(mai_mai_n582_), .B0(mai_mai_n596_), .B1(mai_mai_n502_), .Y(mai_mai_n929_));
  NA4        m0901(.A(mai_mai_n929_), .B(mai_mai_n927_), .C(mai_mai_n926_), .D(mai_mai_n923_), .Y(mai_mai_n930_));
  NO4        m0902(.A(mai_mai_n930_), .B(mai_mai_n922_), .C(mai_mai_n918_), .D(mai_mai_n911_), .Y(mai_mai_n931_));
  NAi31      m0903(.An(mai_mai_n127_), .B(mai_mai_n389_), .C(n), .Y(mai_mai_n932_));
  NO3        m0904(.A(mai_mai_n115_), .B(mai_mai_n312_), .C(mai_mai_n792_), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n933_), .B(mai_mai_n932_), .Y(mai_mai_n934_));
  NO3        m0906(.A(mai_mai_n249_), .B(mai_mai_n127_), .C(mai_mai_n378_), .Y(mai_mai_n935_));
  AOI210     m0907(.A0(mai_mai_n935_), .A1(mai_mai_n471_), .B0(mai_mai_n934_), .Y(mai_mai_n936_));
  NA2        m0908(.A(mai_mai_n463_), .B(i), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n937_), .B(mai_mai_n936_), .Y(mai_mai_n938_));
  NA2        m0910(.A(mai_mai_n212_), .B(mai_mai_n155_), .Y(mai_mai_n939_));
  NO3        m0911(.A(mai_mai_n279_), .B(mai_mai_n414_), .C(mai_mai_n159_), .Y(mai_mai_n940_));
  NOi31      m0912(.An(mai_mai_n939_), .B(mai_mai_n940_), .C(mai_mai_n197_), .Y(mai_mai_n941_));
  NAi21      m0913(.An(mai_mai_n522_), .B(mai_mai_n920_), .Y(mai_mai_n942_));
  NO3        m0914(.A(mai_mai_n408_), .B(mai_mai_n282_), .C(mai_mai_n69_), .Y(mai_mai_n943_));
  AOI220     m0915(.A0(mai_mai_n943_), .A1(mai_mai_n405_), .B0(mai_mai_n452_), .B1(g), .Y(mai_mai_n944_));
  NA2        m0916(.A(mai_mai_n944_), .B(mai_mai_n942_), .Y(mai_mai_n945_));
  NO2        m0917(.A(mai_mai_n613_), .B(mai_mai_n347_), .Y(mai_mai_n946_));
  NA2        m0918(.A(mai_mai_n873_), .B(mai_mai_n864_), .Y(mai_mai_n947_));
  NO3        m0919(.A(mai_mai_n514_), .B(mai_mai_n134_), .C(mai_mai_n196_), .Y(mai_mai_n948_));
  OAI210     m0920(.A0(mai_mai_n948_), .A1(mai_mai_n498_), .B0(mai_mai_n348_), .Y(mai_mai_n949_));
  OAI220     m0921(.A0(mai_mai_n870_), .A1(mai_mai_n877_), .B0(mai_mai_n515_), .B1(mai_mai_n397_), .Y(mai_mai_n950_));
  NA3        m0922(.A(mai_mai_n950_), .B(mai_mai_n949_), .C(mai_mai_n947_), .Y(mai_mai_n951_));
  OAI210     m0923(.A0(mai_mai_n873_), .A1(mai_mai_n865_), .B0(mai_mai_n939_), .Y(mai_mai_n952_));
  NA3        m0924(.A(mai_mai_n909_), .B(mai_mai_n457_), .C(mai_mai_n45_), .Y(mai_mai_n953_));
  NA2        m0925(.A(mai_mai_n953_), .B(mai_mai_n952_), .Y(mai_mai_n954_));
  OR3        m0926(.A(mai_mai_n954_), .B(mai_mai_n951_), .C(mai_mai_n946_), .Y(mai_mai_n955_));
  NO4        m0927(.A(mai_mai_n955_), .B(mai_mai_n945_), .C(mai_mai_n941_), .D(mai_mai_n938_), .Y(mai_mai_n956_));
  NA4        m0928(.A(mai_mai_n956_), .B(mai_mai_n931_), .C(mai_mai_n902_), .D(mai_mai_n886_), .Y(mai13));
  INV        m0929(.A(mai_mai_n45_), .Y(mai_mai_n958_));
  AN2        m0930(.A(c), .B(b), .Y(mai_mai_n959_));
  NA3        m0931(.A(mai_mai_n233_), .B(mai_mai_n959_), .C(m), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n468_), .B(f), .Y(mai_mai_n961_));
  NO4        m0933(.A(mai_mai_n961_), .B(mai_mai_n960_), .C(mai_mai_n958_), .D(mai_mai_n542_), .Y(mai_mai_n962_));
  NA2        m0934(.A(mai_mai_n243_), .B(mai_mai_n959_), .Y(mai_mai_n963_));
  NO3        m0935(.A(mai_mai_n963_), .B(mai_mai_n961_), .C(mai_mai_n904_), .Y(mai_mai_n964_));
  NAi32      m0936(.An(d), .Bn(c), .C(e), .Y(mai_mai_n965_));
  NA2        m0937(.A(mai_mai_n126_), .B(mai_mai_n44_), .Y(mai_mai_n966_));
  NO4        m0938(.A(mai_mai_n966_), .B(mai_mai_n965_), .C(mai_mai_n549_), .D(mai_mai_n278_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n380_), .B(mai_mai_n196_), .Y(mai_mai_n968_));
  AN2        m0940(.A(d), .B(c), .Y(mai_mai_n969_));
  NA2        m0941(.A(mai_mai_n969_), .B(mai_mai_n106_), .Y(mai_mai_n970_));
  NO4        m0942(.A(mai_mai_n970_), .B(mai_mai_n968_), .C(mai_mai_n160_), .D(mai_mai_n151_), .Y(mai_mai_n971_));
  NA2        m0943(.A(mai_mai_n468_), .B(c), .Y(mai_mai_n972_));
  NO4        m0944(.A(mai_mai_n966_), .B(mai_mai_n545_), .C(mai_mai_n972_), .D(mai_mai_n278_), .Y(mai_mai_n973_));
  OR2        m0945(.A(mai_mai_n971_), .B(mai_mai_n973_), .Y(mai_mai_n974_));
  OR4        m0946(.A(mai_mai_n974_), .B(mai_mai_n967_), .C(mai_mai_n964_), .D(mai_mai_n962_), .Y(mai_mai_n975_));
  NAi32      m0947(.An(f), .Bn(e), .C(c), .Y(mai_mai_n976_));
  NO2        m0948(.A(mai_mai_n976_), .B(mai_mai_n131_), .Y(mai_mai_n977_));
  NA2        m0949(.A(mai_mai_n977_), .B(g), .Y(mai_mai_n978_));
  OR3        m0950(.A(mai_mai_n206_), .B(mai_mai_n160_), .C(mai_mai_n151_), .Y(mai_mai_n979_));
  NO2        m0951(.A(mai_mai_n979_), .B(mai_mai_n978_), .Y(mai_mai_n980_));
  NO2        m0952(.A(mai_mai_n972_), .B(mai_mai_n278_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n584_), .B(mai_mai_n1426_), .Y(mai_mai_n982_));
  NOi21      m0954(.An(mai_mai_n981_), .B(mai_mai_n982_), .Y(mai_mai_n983_));
  NO2        m0955(.A(mai_mai_n711_), .B(mai_mai_n102_), .Y(mai_mai_n984_));
  NOi41      m0956(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n985_));
  NA2        m0957(.A(mai_mai_n985_), .B(mai_mai_n984_), .Y(mai_mai_n986_));
  NO2        m0958(.A(mai_mai_n986_), .B(mai_mai_n978_), .Y(mai_mai_n987_));
  OR3        m0959(.A(e), .B(d), .C(c), .Y(mai_mai_n988_));
  NA3        m0960(.A(k), .B(j), .C(i), .Y(mai_mai_n989_));
  NO3        m0961(.A(mai_mai_n989_), .B(mai_mai_n278_), .C(mai_mai_n86_), .Y(mai_mai_n990_));
  NOi21      m0962(.An(mai_mai_n990_), .B(mai_mai_n988_), .Y(mai_mai_n991_));
  OR4        m0963(.A(mai_mai_n991_), .B(mai_mai_n987_), .C(mai_mai_n983_), .D(mai_mai_n980_), .Y(mai_mai_n992_));
  NA3        m0964(.A(mai_mai_n438_), .B(mai_mai_n305_), .C(mai_mai_n54_), .Y(mai_mai_n993_));
  NO2        m0965(.A(mai_mai_n993_), .B(mai_mai_n982_), .Y(mai_mai_n994_));
  NO3        m0966(.A(mai_mai_n993_), .B(mai_mai_n545_), .C(mai_mai_n421_), .Y(mai_mai_n995_));
  NO2        m0967(.A(f), .B(c), .Y(mai_mai_n996_));
  NOi21      m0968(.An(mai_mai_n996_), .B(mai_mai_n413_), .Y(mai_mai_n997_));
  NA2        m0969(.A(mai_mai_n997_), .B(mai_mai_n57_), .Y(mai_mai_n998_));
  OR2        m0970(.A(k), .B(i), .Y(mai_mai_n999_));
  NO3        m0971(.A(mai_mai_n999_), .B(mai_mai_n226_), .C(l), .Y(mai_mai_n1000_));
  NOi31      m0972(.An(mai_mai_n1000_), .B(mai_mai_n998_), .C(j), .Y(mai_mai_n1001_));
  OR3        m0973(.A(mai_mai_n1001_), .B(mai_mai_n995_), .C(mai_mai_n994_), .Y(mai_mai_n1002_));
  OR3        m0974(.A(mai_mai_n1002_), .B(mai_mai_n992_), .C(mai_mai_n975_), .Y(mai02));
  OR2        m0975(.A(l), .B(k), .Y(mai_mai_n1004_));
  OR3        m0976(.A(h), .B(g), .C(f), .Y(mai_mai_n1005_));
  OR3        m0977(.A(n), .B(m), .C(i), .Y(mai_mai_n1006_));
  NO4        m0978(.A(mai_mai_n1006_), .B(mai_mai_n1005_), .C(mai_mai_n1004_), .D(mai_mai_n988_), .Y(mai_mai_n1007_));
  NOi31      m0979(.An(e), .B(d), .C(c), .Y(mai_mai_n1008_));
  AOI210     m0980(.A0(mai_mai_n990_), .A1(mai_mai_n1008_), .B0(mai_mai_n967_), .Y(mai_mai_n1009_));
  AN3        m0981(.A(g), .B(f), .C(c), .Y(mai_mai_n1010_));
  NA3        m0982(.A(mai_mai_n1010_), .B(mai_mai_n438_), .C(h), .Y(mai_mai_n1011_));
  OR2        m0983(.A(mai_mai_n989_), .B(mai_mai_n278_), .Y(mai_mai_n1012_));
  OR2        m0984(.A(mai_mai_n1012_), .B(mai_mai_n1011_), .Y(mai_mai_n1013_));
  NO3        m0985(.A(mai_mai_n993_), .B(mai_mai_n966_), .C(mai_mai_n545_), .Y(mai_mai_n1014_));
  NO2        m0986(.A(mai_mai_n1014_), .B(mai_mai_n980_), .Y(mai_mai_n1015_));
  NA3        m0987(.A(l), .B(k), .C(j), .Y(mai_mai_n1016_));
  NA2        m0988(.A(i), .B(h), .Y(mai_mai_n1017_));
  NO3        m0989(.A(mai_mai_n1017_), .B(mai_mai_n1016_), .C(mai_mai_n119_), .Y(mai_mai_n1018_));
  NO3        m0990(.A(mai_mai_n128_), .B(mai_mai_n260_), .C(mai_mai_n197_), .Y(mai_mai_n1019_));
  AOI210     m0991(.A0(mai_mai_n1019_), .A1(mai_mai_n1018_), .B0(mai_mai_n983_), .Y(mai_mai_n1020_));
  NA3        m0992(.A(c), .B(b), .C(a), .Y(mai_mai_n1021_));
  NO3        m0993(.A(mai_mai_n1021_), .B(mai_mai_n840_), .C(mai_mai_n196_), .Y(mai_mai_n1022_));
  NO3        m0994(.A(mai_mai_n989_), .B(mai_mai_n272_), .C(mai_mai_n47_), .Y(mai_mai_n1023_));
  AOI210     m0995(.A0(mai_mai_n1023_), .A1(mai_mai_n1022_), .B0(mai_mai_n994_), .Y(mai_mai_n1024_));
  AN4        m0996(.A(mai_mai_n1024_), .B(mai_mai_n1020_), .C(mai_mai_n1015_), .D(mai_mai_n1013_), .Y(mai_mai_n1025_));
  NO2        m0997(.A(mai_mai_n970_), .B(mai_mai_n968_), .Y(mai_mai_n1026_));
  NA2        m0998(.A(mai_mai_n986_), .B(mai_mai_n979_), .Y(mai_mai_n1027_));
  AOI210     m0999(.A0(mai_mai_n1027_), .A1(mai_mai_n1026_), .B0(mai_mai_n962_), .Y(mai_mai_n1028_));
  NAi41      m1000(.An(mai_mai_n1007_), .B(mai_mai_n1028_), .C(mai_mai_n1025_), .D(mai_mai_n1009_), .Y(mai03));
  NA4        m1001(.A(mai_mai_n536_), .B(m), .C(mai_mai_n102_), .D(mai_mai_n196_), .Y(mai_mai_n1030_));
  NA2        m1002(.A(mai_mai_n1030_), .B(mai_mai_n338_), .Y(mai_mai_n1031_));
  NO2        m1003(.A(mai_mai_n1031_), .B(mai_mai_n925_), .Y(mai_mai_n1032_));
  INV        m1004(.A(mai_mai_n786_), .Y(mai_mai_n1033_));
  OAI220     m1005(.A0(mai_mai_n1033_), .A1(mai_mai_n639_), .B0(mai_mai_n1032_), .B1(mai_mai_n546_), .Y(mai_mai_n1034_));
  NOi31      m1006(.An(i), .B(k), .C(j), .Y(mai_mai_n1035_));
  NA4        m1007(.A(mai_mai_n1035_), .B(mai_mai_n1008_), .C(mai_mai_n314_), .D(mai_mai_n305_), .Y(mai_mai_n1036_));
  OAI210     m1008(.A0(mai_mai_n763_), .A1(mai_mai_n390_), .B0(mai_mai_n1036_), .Y(mai_mai_n1037_));
  NOi31      m1009(.An(m), .B(n), .C(f), .Y(mai_mai_n1038_));
  NA2        m1010(.A(mai_mai_n1038_), .B(mai_mai_n49_), .Y(mai_mai_n1039_));
  AN2        m1011(.A(e), .B(c), .Y(mai_mai_n1040_));
  NA2        m1012(.A(mai_mai_n1040_), .B(a), .Y(mai_mai_n1041_));
  OAI220     m1013(.A0(mai_mai_n1041_), .A1(mai_mai_n1039_), .B0(mai_mai_n824_), .B1(mai_mai_n396_), .Y(mai_mai_n1042_));
  NA2        m1014(.A(mai_mai_n481_), .B(l), .Y(mai_mai_n1043_));
  NOi31      m1015(.An(mai_mai_n804_), .B(mai_mai_n960_), .C(mai_mai_n1043_), .Y(mai_mai_n1044_));
  NO4        m1016(.A(mai_mai_n1044_), .B(mai_mai_n1042_), .C(mai_mai_n1037_), .D(mai_mai_n924_), .Y(mai_mai_n1045_));
  NO2        m1017(.A(mai_mai_n260_), .B(a), .Y(mai_mai_n1046_));
  INV        m1018(.A(mai_mai_n967_), .Y(mai_mai_n1047_));
  NO2        m1019(.A(mai_mai_n1017_), .B(mai_mai_n455_), .Y(mai_mai_n1048_));
  NO2        m1020(.A(mai_mai_n83_), .B(g), .Y(mai_mai_n1049_));
  AOI210     m1021(.A0(mai_mai_n1049_), .A1(mai_mai_n1048_), .B0(mai_mai_n1000_), .Y(mai_mai_n1050_));
  OR2        m1022(.A(mai_mai_n1050_), .B(mai_mai_n998_), .Y(mai_mai_n1051_));
  NA3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1047_), .C(mai_mai_n1045_), .Y(mai_mai_n1052_));
  NO4        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1034_), .C(mai_mai_n764_), .D(mai_mai_n534_), .Y(mai_mai_n1053_));
  NA2        m1025(.A(c), .B(b), .Y(mai_mai_n1054_));
  NO2        m1026(.A(mai_mai_n651_), .B(mai_mai_n1054_), .Y(mai_mai_n1055_));
  OAI210     m1027(.A0(mai_mai_n382_), .A1(mai_mai_n803_), .B0(mai_mai_n1055_), .Y(mai_mai_n1056_));
  NAi21      m1028(.An(mai_mai_n391_), .B(mai_mai_n1055_), .Y(mai_mai_n1057_));
  NA3        m1029(.A(mai_mai_n397_), .B(mai_mai_n527_), .C(f), .Y(mai_mai_n1058_));
  OAI210     m1030(.A0(mai_mai_n517_), .A1(mai_mai_n39_), .B0(mai_mai_n1046_), .Y(mai_mai_n1059_));
  NA3        m1031(.A(mai_mai_n1059_), .B(mai_mai_n1058_), .C(mai_mai_n1057_), .Y(mai_mai_n1060_));
  NAi21      m1032(.An(f), .B(d), .Y(mai_mai_n1061_));
  NO2        m1033(.A(mai_mai_n1061_), .B(mai_mai_n1021_), .Y(mai_mai_n1062_));
  INV        m1034(.A(mai_mai_n1060_), .Y(mai_mai_n1063_));
  NA2        m1035(.A(mai_mai_n441_), .B(mai_mai_n440_), .Y(mai_mai_n1064_));
  NO2        m1036(.A(mai_mai_n166_), .B(mai_mai_n219_), .Y(mai_mai_n1065_));
  NA2        m1037(.A(mai_mai_n1065_), .B(m), .Y(mai_mai_n1066_));
  NA2        m1038(.A(mai_mai_n283_), .B(mai_mai_n442_), .Y(mai_mai_n1067_));
  AOI210     m1039(.A0(mai_mai_n1067_), .A1(mai_mai_n1064_), .B0(mai_mai_n1066_), .Y(mai_mai_n1068_));
  NA2        m1040(.A(mai_mai_n143_), .B(mai_mai_n33_), .Y(mai_mai_n1069_));
  AOI210     m1041(.A0(mai_mai_n900_), .A1(mai_mai_n1069_), .B0(mai_mai_n197_), .Y(mai_mai_n1070_));
  NA2        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1062_), .Y(mai_mai_n1071_));
  NO2        m1043(.A(mai_mai_n341_), .B(mai_mai_n340_), .Y(mai_mai_n1072_));
  AOI210     m1044(.A0(mai_mai_n1065_), .A1(mai_mai_n399_), .B0(mai_mai_n894_), .Y(mai_mai_n1073_));
  NAi31      m1045(.An(mai_mai_n1072_), .B(mai_mai_n1073_), .C(mai_mai_n1071_), .Y(mai_mai_n1074_));
  NO2        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1068_), .Y(mai_mai_n1075_));
  NA4        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1063_), .C(mai_mai_n1056_), .D(mai_mai_n1053_), .Y(mai00));
  AOI210     m1048(.A0(mai_mai_n271_), .A1(mai_mai_n197_), .B0(mai_mai_n252_), .Y(mai_mai_n1077_));
  NO2        m1049(.A(mai_mai_n1077_), .B(mai_mai_n538_), .Y(mai_mai_n1078_));
  AOI210     m1050(.A0(mai_mai_n837_), .A1(mai_mai_n878_), .B0(mai_mai_n1037_), .Y(mai_mai_n1079_));
  NO2        m1051(.A(mai_mai_n1014_), .B(mai_mai_n894_), .Y(mai_mai_n1080_));
  NA3        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1079_), .C(mai_mai_n926_), .Y(mai_mai_n1081_));
  NA2        m1053(.A(mai_mai_n483_), .B(f), .Y(mai_mai_n1082_));
  OAI210     m1054(.A0(mai_mai_n933_), .A1(mai_mai_n40_), .B0(mai_mai_n598_), .Y(mai_mai_n1083_));
  NA3        m1055(.A(mai_mai_n1083_), .B(mai_mai_n241_), .C(n), .Y(mai_mai_n1084_));
  AOI210     m1056(.A0(mai_mai_n1084_), .A1(mai_mai_n1082_), .B0(mai_mai_n970_), .Y(mai_mai_n1085_));
  NO4        m1057(.A(mai_mai_n1085_), .B(mai_mai_n1081_), .C(mai_mai_n1078_), .D(mai_mai_n992_), .Y(mai_mai_n1086_));
  NA3        m1058(.A(mai_mai_n150_), .B(mai_mai_n45_), .C(mai_mai_n44_), .Y(mai_mai_n1087_));
  NA3        m1059(.A(d), .B(mai_mai_n54_), .C(b), .Y(mai_mai_n1088_));
  NOi31      m1060(.An(n), .B(m), .C(i), .Y(mai_mai_n1089_));
  NA3        m1061(.A(mai_mai_n1089_), .B(mai_mai_n601_), .C(mai_mai_n49_), .Y(mai_mai_n1090_));
  OAI210     m1062(.A0(mai_mai_n1088_), .A1(mai_mai_n1087_), .B0(mai_mai_n1090_), .Y(mai_mai_n1091_));
  NO3        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1072_), .C(mai_mai_n856_), .Y(mai_mai_n1092_));
  NO4        m1064(.A(mai_mai_n458_), .B(mai_mai_n326_), .C(mai_mai_n1054_), .D(mai_mai_n57_), .Y(mai_mai_n1093_));
  NA3        m1065(.A(mai_mai_n353_), .B(mai_mai_n202_), .C(g), .Y(mai_mai_n1094_));
  OR2        m1066(.A(mai_mai_n1094_), .B(mai_mai_n1088_), .Y(mai_mai_n1095_));
  NO2        m1067(.A(h), .B(g), .Y(mai_mai_n1096_));
  NA4        m1068(.A(mai_mai_n471_), .B(mai_mai_n438_), .C(mai_mai_n1096_), .D(mai_mai_n959_), .Y(mai_mai_n1097_));
  NA2        m1069(.A(mai_mai_n881_), .B(mai_mai_n537_), .Y(mai_mai_n1098_));
  AOI220     m1070(.A0(mai_mai_n290_), .A1(mai_mai_n230_), .B0(mai_mai_n161_), .B1(mai_mai_n133_), .Y(mai_mai_n1099_));
  NA4        m1071(.A(mai_mai_n1099_), .B(mai_mai_n1098_), .C(mai_mai_n1097_), .D(mai_mai_n1095_), .Y(mai_mai_n1100_));
  NO2        m1072(.A(mai_mai_n1100_), .B(mai_mai_n1093_), .Y(mai_mai_n1101_));
  NO2        m1073(.A(mai_mai_n221_), .B(mai_mai_n165_), .Y(mai_mai_n1102_));
  NA2        m1074(.A(mai_mai_n1102_), .B(mai_mai_n397_), .Y(mai_mai_n1103_));
  NA3        m1075(.A(mai_mai_n163_), .B(mai_mai_n102_), .C(g), .Y(mai_mai_n1104_));
  NA3        m1076(.A(mai_mai_n438_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1105_));
  NOi31      m1077(.An(mai_mai_n811_), .B(mai_mai_n1105_), .C(mai_mai_n1104_), .Y(mai_mai_n1106_));
  NAi31      m1078(.An(mai_mai_n170_), .B(mai_mai_n799_), .C(mai_mai_n438_), .Y(mai_mai_n1107_));
  NAi31      m1079(.An(mai_mai_n1106_), .B(mai_mai_n1107_), .C(mai_mai_n1103_), .Y(mai_mai_n1108_));
  NO2        m1080(.A(mai_mai_n251_), .B(mai_mai_n69_), .Y(mai_mai_n1109_));
  NO3        m1081(.A(mai_mai_n396_), .B(mai_mai_n774_), .C(n), .Y(mai_mai_n1110_));
  AOI210     m1082(.A0(mai_mai_n1110_), .A1(mai_mai_n1109_), .B0(mai_mai_n1007_), .Y(mai_mai_n1111_));
  NAi31      m1083(.An(mai_mai_n973_), .B(mai_mai_n1111_), .C(mai_mai_n68_), .Y(mai_mai_n1112_));
  NO2        m1084(.A(mai_mai_n1112_), .B(mai_mai_n1108_), .Y(mai_mai_n1113_));
  AN3        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1101_), .C(mai_mai_n1092_), .Y(mai_mai_n1114_));
  NA3        m1086(.A(mai_mai_n1038_), .B(mai_mai_n563_), .C(mai_mai_n437_), .Y(mai_mai_n1115_));
  NA3        m1087(.A(mai_mai_n1115_), .B(mai_mai_n530_), .C(mai_mai_n224_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(mai_mai_n1031_), .B(mai_mai_n506_), .Y(mai_mai_n1117_));
  NA4        m1089(.A(mai_mai_n601_), .B(mai_mai_n189_), .C(mai_mai_n202_), .D(mai_mai_n147_), .Y(mai_mai_n1118_));
  NA3        m1090(.A(mai_mai_n1118_), .B(mai_mai_n1117_), .C(mai_mai_n268_), .Y(mai_mai_n1119_));
  OR3        m1091(.A(mai_mai_n970_), .B(mai_mai_n249_), .C(mai_mai_n204_), .Y(mai_mai_n1120_));
  NO2        m1092(.A(mai_mai_n200_), .B(mai_mai_n197_), .Y(mai_mai_n1121_));
  NA2        m1093(.A(n), .B(e), .Y(mai_mai_n1122_));
  NO2        m1094(.A(mai_mai_n1122_), .B(mai_mai_n131_), .Y(mai_mai_n1123_));
  AOI220     m1095(.A0(mai_mai_n1123_), .A1(mai_mai_n250_), .B0(mai_mai_n790_), .B1(mai_mai_n1121_), .Y(mai_mai_n1124_));
  OAI210     m1096(.A0(mai_mai_n327_), .A1(mai_mai_n284_), .B0(mai_mai_n419_), .Y(mai_mai_n1125_));
  NA3        m1097(.A(mai_mai_n1125_), .B(mai_mai_n1124_), .C(mai_mai_n1120_), .Y(mai_mai_n1126_));
  AOI210     m1098(.A0(mai_mai_n1123_), .A1(mai_mai_n794_), .B0(mai_mai_n764_), .Y(mai_mai_n1127_));
  AOI220     m1099(.A0(mai_mai_n890_), .A1(mai_mai_n537_), .B0(mai_mai_n601_), .B1(mai_mai_n227_), .Y(mai_mai_n1128_));
  NO2        m1100(.A(mai_mai_n63_), .B(h), .Y(mai_mai_n1129_));
  NO3        m1101(.A(mai_mai_n970_), .B(mai_mai_n968_), .C(mai_mai_n674_), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n1004_), .B(mai_mai_n119_), .Y(mai_mai_n1131_));
  AN2        m1103(.A(mai_mai_n1131_), .B(mai_mai_n1019_), .Y(mai_mai_n1132_));
  OAI210     m1104(.A0(mai_mai_n1132_), .A1(mai_mai_n1130_), .B0(mai_mai_n1129_), .Y(mai_mai_n1133_));
  NA4        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1128_), .C(mai_mai_n1127_), .D(mai_mai_n807_), .Y(mai_mai_n1134_));
  NO4        m1106(.A(mai_mai_n1134_), .B(mai_mai_n1126_), .C(mai_mai_n1119_), .D(mai_mai_n1116_), .Y(mai_mai_n1135_));
  NA2        m1107(.A(mai_mai_n778_), .B(mai_mai_n706_), .Y(mai_mai_n1136_));
  NA4        m1108(.A(mai_mai_n1136_), .B(mai_mai_n1135_), .C(mai_mai_n1114_), .D(mai_mai_n1086_), .Y(mai01));
  AN2        m1109(.A(mai_mai_n949_), .B(mai_mai_n947_), .Y(mai_mai_n1138_));
  NO4        m1110(.A(mai_mai_n750_), .B(mai_mai_n742_), .C(mai_mai_n449_), .D(mai_mai_n258_), .Y(mai_mai_n1139_));
  NA2        m1111(.A(mai_mai_n364_), .B(i), .Y(mai_mai_n1140_));
  NA3        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1139_), .C(mai_mai_n1138_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(mai_mai_n522_), .B(mai_mai_n248_), .Y(mai_mai_n1142_));
  NA2        m1114(.A(mai_mai_n897_), .B(mai_mai_n1142_), .Y(mai_mai_n1143_));
  NA3        m1115(.A(mai_mai_n1143_), .B(mai_mai_n852_), .C(mai_mai_n304_), .Y(mai_mai_n1144_));
  NA2        m1116(.A(mai_mai_n658_), .B(mai_mai_n90_), .Y(mai_mai_n1145_));
  INV        m1117(.A(mai_mai_n108_), .Y(mai_mai_n1146_));
  OA220      m1118(.A0(mai_mai_n1146_), .A1(mai_mai_n544_), .B0(mai_mai_n614_), .B1(mai_mai_n338_), .Y(mai_mai_n1147_));
  NAi41      m1119(.An(mai_mai_n146_), .B(mai_mai_n1147_), .C(mai_mai_n1118_), .D(mai_mai_n836_), .Y(mai_mai_n1148_));
  NO2        m1120(.A(mai_mai_n732_), .B(mai_mai_n485_), .Y(mai_mai_n1149_));
  OR2        m1121(.A(mai_mai_n180_), .B(mai_mai_n178_), .Y(mai_mai_n1150_));
  NA3        m1122(.A(mai_mai_n1150_), .B(mai_mai_n1149_), .C(mai_mai_n124_), .Y(mai_mai_n1151_));
  NO4        m1123(.A(mai_mai_n1151_), .B(mai_mai_n1148_), .C(mai_mai_n1144_), .D(mai_mai_n1141_), .Y(mai_mai_n1152_));
  INV        m1124(.A(mai_mai_n1094_), .Y(mai_mai_n1153_));
  NA2        m1125(.A(mai_mai_n1153_), .B(mai_mai_n502_), .Y(mai_mai_n1154_));
  NA2        m1126(.A(mai_mai_n508_), .B(mai_mai_n366_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(mai_mai_n531_), .B(mai_mai_n1155_), .Y(mai_mai_n1156_));
  AOI210     m1128(.A0(mai_mai_n187_), .A1(mai_mai_n85_), .B0(mai_mai_n196_), .Y(mai_mai_n1157_));
  OAI210     m1129(.A0(mai_mai_n756_), .A1(mai_mai_n397_), .B0(mai_mai_n1157_), .Y(mai_mai_n1158_));
  AN3        m1130(.A(m), .B(l), .C(k), .Y(mai_mai_n1159_));
  OAI210     m1131(.A0(mai_mai_n329_), .A1(mai_mai_n34_), .B0(mai_mai_n1159_), .Y(mai_mai_n1160_));
  NA2        m1132(.A(mai_mai_n186_), .B(mai_mai_n34_), .Y(mai_mai_n1161_));
  AO210      m1133(.A0(mai_mai_n1161_), .A1(mai_mai_n1160_), .B0(mai_mai_n303_), .Y(mai_mai_n1162_));
  NA4        m1134(.A(mai_mai_n1162_), .B(mai_mai_n1158_), .C(mai_mai_n1156_), .D(mai_mai_n1154_), .Y(mai_mai_n1163_));
  INV        m1135(.A(mai_mai_n558_), .Y(mai_mai_n1164_));
  OAI210     m1136(.A0(mai_mai_n1146_), .A1(mai_mai_n553_), .B0(mai_mai_n1164_), .Y(mai_mai_n1165_));
  NA2        m1137(.A(mai_mai_n257_), .B(mai_mai_n180_), .Y(mai_mai_n1166_));
  NA2        m1138(.A(mai_mai_n1166_), .B(mai_mai_n619_), .Y(mai_mai_n1167_));
  NO3        m1139(.A(mai_mai_n763_), .B(mai_mai_n187_), .C(mai_mai_n378_), .Y(mai_mai_n1168_));
  NO2        m1140(.A(mai_mai_n1168_), .B(mai_mai_n894_), .Y(mai_mai_n1169_));
  NA2        m1141(.A(mai_mai_n298_), .B(mai_mai_n624_), .Y(mai_mai_n1170_));
  NA4        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1169_), .C(mai_mai_n1167_), .D(mai_mai_n734_), .Y(mai_mai_n1171_));
  NO3        m1143(.A(mai_mai_n1171_), .B(mai_mai_n1165_), .C(mai_mai_n1163_), .Y(mai_mai_n1172_));
  NA3        m1144(.A(mai_mai_n560_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1173_));
  NO2        m1145(.A(mai_mai_n1173_), .B(mai_mai_n187_), .Y(mai_mai_n1174_));
  AOI210     m1146(.A0(mai_mai_n478_), .A1(mai_mai_n56_), .B0(mai_mai_n1174_), .Y(mai_mai_n1175_));
  OR3        m1147(.A(mai_mai_n1145_), .B(mai_mai_n561_), .C(i), .Y(mai_mai_n1176_));
  NO2        m1148(.A(mai_mai_n190_), .B(mai_mai_n101_), .Y(mai_mai_n1177_));
  NO2        m1149(.A(mai_mai_n1177_), .B(mai_mai_n1091_), .Y(mai_mai_n1178_));
  NA4        m1150(.A(mai_mai_n1178_), .B(mai_mai_n1176_), .C(mai_mai_n1175_), .D(mai_mai_n705_), .Y(mai_mai_n1179_));
  NO3        m1151(.A(mai_mai_n75_), .B(mai_mai_n272_), .C(mai_mai_n44_), .Y(mai_mai_n1180_));
  OR2        m1152(.A(mai_mai_n1094_), .B(mai_mai_n1088_), .Y(mai_mai_n1181_));
  NO2        m1153(.A(mai_mai_n338_), .B(mai_mai_n67_), .Y(mai_mai_n1182_));
  INV        m1154(.A(mai_mai_n1182_), .Y(mai_mai_n1183_));
  NA2        m1155(.A(mai_mai_n1180_), .B(mai_mai_n757_), .Y(mai_mai_n1184_));
  NA4        m1156(.A(mai_mai_n1184_), .B(mai_mai_n1183_), .C(mai_mai_n1181_), .D(mai_mai_n356_), .Y(mai_mai_n1185_));
  NO2        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1179_), .Y(mai_mai_n1186_));
  NO2        m1158(.A(mai_mai_n118_), .B(mai_mai_n44_), .Y(mai_mai_n1187_));
  NO2        m1159(.A(mai_mai_n44_), .B(mai_mai_n40_), .Y(mai_mai_n1188_));
  AO220      m1160(.A0(mai_mai_n1188_), .A1(mai_mai_n579_), .B0(mai_mai_n1187_), .B1(mai_mai_n656_), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n1189_), .B(mai_mai_n312_), .Y(mai_mai_n1190_));
  INV        m1162(.A(mai_mai_n122_), .Y(mai_mai_n1191_));
  NO3        m1163(.A(mai_mai_n1017_), .B(mai_mai_n160_), .C(mai_mai_n83_), .Y(mai_mai_n1192_));
  AOI220     m1164(.A0(mai_mai_n1192_), .A1(mai_mai_n1191_), .B0(mai_mai_n1180_), .B1(mai_mai_n907_), .Y(mai_mai_n1193_));
  NA2        m1165(.A(mai_mai_n1193_), .B(mai_mai_n1190_), .Y(mai_mai_n1194_));
  NO2        m1166(.A(mai_mai_n571_), .B(mai_mai_n570_), .Y(mai_mai_n1195_));
  NO4        m1167(.A(mai_mai_n1017_), .B(mai_mai_n1195_), .C(mai_mai_n158_), .D(mai_mai_n83_), .Y(mai_mai_n1196_));
  NO3        m1168(.A(mai_mai_n1196_), .B(mai_mai_n1194_), .C(mai_mai_n590_), .Y(mai_mai_n1197_));
  NA4        m1169(.A(mai_mai_n1197_), .B(mai_mai_n1186_), .C(mai_mai_n1172_), .D(mai_mai_n1152_), .Y(mai06));
  NO2        m1170(.A(mai_mai_n379_), .B(mai_mai_n528_), .Y(mai_mai_n1199_));
  INV        m1171(.A(mai_mai_n681_), .Y(mai_mai_n1200_));
  NA2        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1199_), .Y(mai_mai_n1201_));
  NO2        m1173(.A(mai_mai_n206_), .B(mai_mai_n93_), .Y(mai_mai_n1202_));
  OAI210     m1174(.A0(mai_mai_n1202_), .A1(mai_mai_n1192_), .B0(mai_mai_n352_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n1203_), .B(mai_mai_n1201_), .Y(mai_mai_n1204_));
  NO2        m1176(.A(mai_mai_n1204_), .B(mai_mai_n240_), .Y(mai_mai_n1205_));
  NO2        m1177(.A(mai_mai_n272_), .B(mai_mai_n44_), .Y(mai_mai_n1206_));
  NA2        m1178(.A(mai_mai_n1206_), .B(mai_mai_n908_), .Y(mai_mai_n1207_));
  AOI210     m1179(.A0(mai_mai_n1206_), .A1(mai_mai_n525_), .B0(mai_mai_n1189_), .Y(mai_mai_n1208_));
  AOI210     m1180(.A0(mai_mai_n1208_), .A1(mai_mai_n1207_), .B0(mai_mai_n309_), .Y(mai_mai_n1209_));
  NO2        m1181(.A(mai_mai_n85_), .B(mai_mai_n40_), .Y(mai_mai_n1210_));
  NA2        m1182(.A(mai_mai_n1210_), .B(mai_mai_n594_), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n488_), .B(mai_mai_n155_), .Y(mai_mai_n1212_));
  NO2        m1184(.A(mai_mai_n564_), .B(mai_mai_n1039_), .Y(mai_mai_n1213_));
  OAI210     m1185(.A0(mai_mai_n432_), .A1(mai_mai_n231_), .B0(mai_mai_n846_), .Y(mai_mai_n1214_));
  NO3        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1213_), .C(mai_mai_n1212_), .Y(mai_mai_n1215_));
  OR2        m1187(.A(mai_mai_n557_), .B(mai_mai_n556_), .Y(mai_mai_n1216_));
  NO2        m1188(.A(mai_mai_n337_), .B(mai_mai_n123_), .Y(mai_mai_n1217_));
  AOI210     m1189(.A0(mai_mai_n1217_), .A1(mai_mai_n547_), .B0(mai_mai_n1216_), .Y(mai_mai_n1218_));
  NA3        m1190(.A(mai_mai_n1218_), .B(mai_mai_n1215_), .C(mai_mai_n1211_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n697_), .B(mai_mai_n336_), .Y(mai_mai_n1220_));
  INV        m1192(.A(mai_mai_n707_), .Y(mai_mai_n1221_));
  NOi21      m1193(.An(mai_mai_n1220_), .B(mai_mai_n1221_), .Y(mai_mai_n1222_));
  AN2        m1194(.A(mai_mai_n890_), .B(mai_mai_n597_), .Y(mai_mai_n1223_));
  NO4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n1222_), .C(mai_mai_n1219_), .D(mai_mai_n1209_), .Y(mai_mai_n1224_));
  NO2        m1196(.A(mai_mai_n749_), .B(mai_mai_n253_), .Y(mai_mai_n1225_));
  OAI220     m1197(.A0(mai_mai_n681_), .A1(mai_mai_n46_), .B0(mai_mai_n206_), .B1(mai_mai_n573_), .Y(mai_mai_n1226_));
  OAI210     m1198(.A0(mai_mai_n253_), .A1(c), .B0(mai_mai_n593_), .Y(mai_mai_n1227_));
  AOI220     m1199(.A0(mai_mai_n1227_), .A1(mai_mai_n1226_), .B0(mai_mai_n1225_), .B1(mai_mai_n244_), .Y(mai_mai_n1228_));
  NO3        m1200(.A(mai_mai_n226_), .B(mai_mai_n93_), .C(mai_mai_n260_), .Y(mai_mai_n1229_));
  OAI220     m1201(.A0(mai_mai_n648_), .A1(mai_mai_n231_), .B0(mai_mai_n484_), .B1(mai_mai_n488_), .Y(mai_mai_n1230_));
  NO3        m1202(.A(mai_mai_n1230_), .B(mai_mai_n1229_), .C(mai_mai_n1042_), .Y(mai_mai_n1231_));
  NA4        m1203(.A(mai_mai_n740_), .B(mai_mai_n739_), .C(mai_mai_n407_), .D(mai_mai_n817_), .Y(mai_mai_n1232_));
  NAi31      m1204(.An(mai_mai_n697_), .B(mai_mai_n1232_), .C(mai_mai_n186_), .Y(mai_mai_n1233_));
  NA4        m1205(.A(mai_mai_n1233_), .B(mai_mai_n1231_), .C(mai_mai_n1228_), .D(mai_mai_n1128_), .Y(mai_mai_n1234_));
  OR2        m1206(.A(mai_mai_n731_), .B(mai_mai_n511_), .Y(mai_mai_n1235_));
  OR3        m1207(.A(mai_mai_n340_), .B(mai_mai_n206_), .C(mai_mai_n573_), .Y(mai_mai_n1236_));
  INV        m1208(.A(mai_mai_n342_), .Y(mai_mai_n1237_));
  NA3        m1209(.A(mai_mai_n1237_), .B(mai_mai_n1236_), .C(mai_mai_n1235_), .Y(mai_mai_n1238_));
  AOI220     m1210(.A0(mai_mai_n1220_), .A1(mai_mai_n706_), .B0(mai_mai_n1217_), .B1(mai_mai_n220_), .Y(mai_mai_n1239_));
  AN2        m1211(.A(mai_mai_n865_), .B(mai_mai_n864_), .Y(mai_mai_n1240_));
  NO4        m1212(.A(mai_mai_n1240_), .B(mai_mai_n815_), .C(mai_mai_n474_), .D(mai_mai_n452_), .Y(mai_mai_n1241_));
  NA3        m1213(.A(mai_mai_n1241_), .B(mai_mai_n1239_), .C(mai_mai_n1184_), .Y(mai_mai_n1242_));
  NAi21      m1214(.An(j), .B(i), .Y(mai_mai_n1243_));
  NO4        m1215(.A(mai_mai_n1195_), .B(mai_mai_n1243_), .C(mai_mai_n413_), .D(mai_mai_n217_), .Y(mai_mai_n1244_));
  NO4        m1216(.A(mai_mai_n1244_), .B(mai_mai_n1242_), .C(mai_mai_n1238_), .D(mai_mai_n1234_), .Y(mai_mai_n1245_));
  NA4        m1217(.A(mai_mai_n1245_), .B(mai_mai_n1224_), .C(mai_mai_n1205_), .D(mai_mai_n1197_), .Y(mai07));
  NOi21      m1218(.An(j), .B(k), .Y(mai_mai_n1247_));
  NA4        m1219(.A(mai_mai_n163_), .B(mai_mai_n98_), .C(mai_mai_n1247_), .D(f), .Y(mai_mai_n1248_));
  NAi32      m1220(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1249_));
  NO3        m1221(.A(mai_mai_n1249_), .B(g), .C(f), .Y(mai_mai_n1250_));
  OAI210     m1222(.A0(i), .A1(mai_mai_n454_), .B0(mai_mai_n1250_), .Y(mai_mai_n1251_));
  NAi21      m1223(.An(f), .B(c), .Y(mai_mai_n1252_));
  OR2        m1224(.A(e), .B(d), .Y(mai_mai_n1253_));
  OAI220     m1225(.A0(mai_mai_n1253_), .A1(mai_mai_n1252_), .B0(mai_mai_n583_), .B1(mai_mai_n294_), .Y(mai_mai_n1254_));
  NA3        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1426_), .C(mai_mai_n163_), .Y(mai_mai_n1255_));
  NOi31      m1227(.An(n), .B(m), .C(b), .Y(mai_mai_n1256_));
  NO3        m1228(.A(mai_mai_n119_), .B(mai_mai_n421_), .C(h), .Y(mai_mai_n1257_));
  NA3        m1229(.A(mai_mai_n1255_), .B(mai_mai_n1251_), .C(mai_mai_n1248_), .Y(mai_mai_n1258_));
  NOi41      m1230(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1259_));
  NA3        m1231(.A(mai_mai_n1259_), .B(mai_mai_n808_), .C(mai_mai_n380_), .Y(mai_mai_n1260_));
  NO2        m1232(.A(mai_mai_n1260_), .B(mai_mai_n54_), .Y(mai_mai_n1261_));
  NO2        m1233(.A(k), .B(i), .Y(mai_mai_n1262_));
  NA2        m1234(.A(mai_mai_n83_), .B(mai_mai_n44_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n976_), .B(mai_mai_n413_), .Y(mai_mai_n1264_));
  NA3        m1236(.A(mai_mai_n1264_), .B(mai_mai_n1263_), .C(mai_mai_n197_), .Y(mai_mai_n1265_));
  NO2        m1237(.A(mai_mai_n989_), .B(mai_mai_n278_), .Y(mai_mai_n1266_));
  NA2        m1238(.A(mai_mai_n512_), .B(mai_mai_n76_), .Y(mai_mai_n1267_));
  NA2        m1239(.A(mai_mai_n1129_), .B(mai_mai_n262_), .Y(mai_mai_n1268_));
  NA3        m1240(.A(mai_mai_n1268_), .B(mai_mai_n1267_), .C(mai_mai_n1265_), .Y(mai_mai_n1269_));
  NO3        m1241(.A(mai_mai_n1269_), .B(mai_mai_n1261_), .C(mai_mai_n1258_), .Y(mai_mai_n1270_));
  NO3        m1242(.A(e), .B(d), .C(c), .Y(mai_mai_n1271_));
  NA2        m1243(.A(mai_mai_n1424_), .B(mai_mai_n1271_), .Y(mai_mai_n1272_));
  NO2        m1244(.A(mai_mai_n1272_), .B(mai_mai_n197_), .Y(mai_mai_n1273_));
  NA3        m1245(.A(mai_mai_n645_), .B(mai_mai_n632_), .C(mai_mai_n102_), .Y(mai_mai_n1274_));
  NO2        m1246(.A(mai_mai_n1274_), .B(mai_mai_n44_), .Y(mai_mai_n1275_));
  NO2        m1247(.A(l), .B(k), .Y(mai_mai_n1276_));
  NOi41      m1248(.An(mai_mai_n516_), .B(mai_mai_n1276_), .C(mai_mai_n447_), .D(mai_mai_n413_), .Y(mai_mai_n1277_));
  NO3        m1249(.A(mai_mai_n413_), .B(d), .C(c), .Y(mai_mai_n1278_));
  NO3        m1250(.A(mai_mai_n1277_), .B(mai_mai_n1275_), .C(mai_mai_n1273_), .Y(mai_mai_n1279_));
  NO2        m1251(.A(mai_mai_n132_), .B(h), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n999_), .B(l), .Y(mai_mai_n1281_));
  NO2        m1253(.A(g), .B(c), .Y(mai_mai_n1282_));
  NA3        m1254(.A(mai_mai_n1282_), .B(mai_mai_n128_), .C(mai_mai_n171_), .Y(mai_mai_n1283_));
  NO2        m1255(.A(mai_mai_n1283_), .B(mai_mai_n1281_), .Y(mai_mai_n1284_));
  NA2        m1256(.A(mai_mai_n1284_), .B(mai_mai_n163_), .Y(mai_mai_n1285_));
  NO2        m1257(.A(mai_mai_n423_), .B(a), .Y(mai_mai_n1286_));
  NA3        m1258(.A(mai_mai_n1286_), .B(mai_mai_n1427_), .C(mai_mai_n103_), .Y(mai_mai_n1287_));
  NO2        m1259(.A(i), .B(h), .Y(mai_mai_n1288_));
  NA2        m1260(.A(mai_mai_n1061_), .B(h), .Y(mai_mai_n1289_));
  NA2        m1261(.A(mai_mai_n125_), .B(mai_mai_n202_), .Y(mai_mai_n1290_));
  NO2        m1262(.A(mai_mai_n1290_), .B(mai_mai_n1289_), .Y(mai_mai_n1291_));
  NO2        m1263(.A(mai_mai_n703_), .B(mai_mai_n172_), .Y(mai_mai_n1292_));
  NOi31      m1264(.An(m), .B(n), .C(b), .Y(mai_mai_n1293_));
  NOi31      m1265(.An(f), .B(d), .C(c), .Y(mai_mai_n1294_));
  NA2        m1266(.A(mai_mai_n1294_), .B(mai_mai_n1293_), .Y(mai_mai_n1295_));
  INV        m1267(.A(mai_mai_n1295_), .Y(mai_mai_n1296_));
  NO3        m1268(.A(mai_mai_n1296_), .B(mai_mai_n1292_), .C(mai_mai_n1291_), .Y(mai_mai_n1297_));
  NA2        m1269(.A(mai_mai_n1010_), .B(mai_mai_n438_), .Y(mai_mai_n1298_));
  OAI210     m1270(.A0(mai_mai_n166_), .A1(mai_mai_n499_), .B0(mai_mai_n985_), .Y(mai_mai_n1299_));
  AN4        m1271(.A(mai_mai_n1299_), .B(mai_mai_n1297_), .C(mai_mai_n1287_), .D(mai_mai_n1285_), .Y(mai_mai_n1300_));
  NA2        m1272(.A(mai_mai_n1256_), .B(mai_mai_n349_), .Y(mai_mai_n1301_));
  NA2        m1273(.A(mai_mai_n1018_), .B(mai_mai_n1298_), .Y(mai_mai_n1302_));
  INV        m1274(.A(mai_mai_n1302_), .Y(mai_mai_n1303_));
  NO4        m1275(.A(mai_mai_n119_), .B(g), .C(f), .D(e), .Y(mai_mai_n1304_));
  NA3        m1276(.A(mai_mai_n1262_), .B(mai_mai_n263_), .C(h), .Y(mai_mai_n1305_));
  NA2        m1277(.A(mai_mai_n179_), .B(mai_mai_n92_), .Y(mai_mai_n1306_));
  OR2        m1278(.A(e), .B(a), .Y(mai_mai_n1307_));
  NOi41      m1279(.An(h), .B(f), .C(e), .D(a), .Y(mai_mai_n1308_));
  NA2        m1280(.A(mai_mai_n1308_), .B(mai_mai_n103_), .Y(mai_mai_n1309_));
  NA2        m1281(.A(mai_mai_n1259_), .B(mai_mai_n1276_), .Y(mai_mai_n1310_));
  NA2        m1282(.A(mai_mai_n1310_), .B(mai_mai_n1309_), .Y(mai_mai_n1311_));
  OR3        m1283(.A(mai_mai_n511_), .B(mai_mai_n510_), .C(mai_mai_n102_), .Y(mai_mai_n1312_));
  NA2        m1284(.A(mai_mai_n1038_), .B(mai_mai_n378_), .Y(mai_mai_n1313_));
  NO2        m1285(.A(mai_mai_n1313_), .B(mai_mai_n406_), .Y(mai_mai_n1314_));
  AO210      m1286(.A0(mai_mai_n1314_), .A1(mai_mai_n106_), .B0(mai_mai_n1311_), .Y(mai_mai_n1315_));
  NO2        m1287(.A(mai_mai_n1315_), .B(mai_mai_n1303_), .Y(mai_mai_n1316_));
  NA4        m1288(.A(mai_mai_n1316_), .B(mai_mai_n1300_), .C(mai_mai_n1279_), .D(mai_mai_n1270_), .Y(mai_mai_n1317_));
  NO2        m1289(.A(mai_mai_n1054_), .B(mai_mai_n100_), .Y(mai_mai_n1318_));
  NA2        m1290(.A(mai_mai_n349_), .B(mai_mai_n54_), .Y(mai_mai_n1319_));
  NA2        m1291(.A(mai_mai_n198_), .B(mai_mai_n163_), .Y(mai_mai_n1320_));
  AOI210     m1292(.A0(mai_mai_n1320_), .A1(mai_mai_n1104_), .B0(mai_mai_n1319_), .Y(mai_mai_n1321_));
  NO2        m1293(.A(mai_mai_n361_), .B(j), .Y(mai_mai_n1322_));
  NAi41      m1294(.An(mai_mai_n1288_), .B(mai_mai_n997_), .C(mai_mai_n151_), .D(mai_mai_n135_), .Y(mai_mai_n1323_));
  INV        m1295(.A(mai_mai_n1323_), .Y(mai_mai_n1324_));
  NA3        m1296(.A(g), .B(mai_mai_n1322_), .C(mai_mai_n143_), .Y(mai_mai_n1325_));
  INV        m1297(.A(mai_mai_n1325_), .Y(mai_mai_n1326_));
  NO3        m1298(.A(mai_mai_n697_), .B(mai_mai_n158_), .C(mai_mai_n380_), .Y(mai_mai_n1327_));
  NO3        m1299(.A(mai_mai_n1327_), .B(mai_mai_n1326_), .C(mai_mai_n1324_), .Y(mai_mai_n1328_));
  NO3        m1300(.A(mai_mai_n1006_), .B(mai_mai_n541_), .C(g), .Y(mai_mai_n1329_));
  NOi21      m1301(.An(mai_mai_n1320_), .B(mai_mai_n1329_), .Y(mai_mai_n1330_));
  AOI210     m1302(.A0(mai_mai_n1330_), .A1(mai_mai_n1306_), .B0(mai_mai_n976_), .Y(mai_mai_n1331_));
  OR2        m1303(.A(n), .B(i), .Y(mai_mai_n1332_));
  OAI210     m1304(.A0(mai_mai_n1332_), .A1(mai_mai_n996_), .B0(mai_mai_n47_), .Y(mai_mai_n1333_));
  AOI220     m1305(.A0(mai_mai_n1333_), .A1(mai_mai_n1096_), .B0(mai_mai_n767_), .B1(mai_mai_n179_), .Y(mai_mai_n1334_));
  INV        m1306(.A(mai_mai_n1334_), .Y(mai_mai_n1335_));
  NO2        m1307(.A(mai_mai_n119_), .B(l), .Y(mai_mai_n1336_));
  NO2        m1308(.A(mai_mai_n206_), .B(k), .Y(mai_mai_n1337_));
  OAI210     m1309(.A0(mai_mai_n1337_), .A1(mai_mai_n1288_), .B0(mai_mai_n1336_), .Y(mai_mai_n1338_));
  NO2        m1310(.A(mai_mai_n1338_), .B(mai_mai_n31_), .Y(mai_mai_n1339_));
  NO3        m1311(.A(mai_mai_n1312_), .B(mai_mai_n438_), .C(mai_mai_n323_), .Y(mai_mai_n1340_));
  NO4        m1312(.A(mai_mai_n1340_), .B(mai_mai_n1339_), .C(mai_mai_n1335_), .D(mai_mai_n1331_), .Y(mai_mai_n1341_));
  NO3        m1313(.A(mai_mai_n1021_), .B(mai_mai_n1253_), .C(mai_mai_n47_), .Y(mai_mai_n1342_));
  NO2        m1314(.A(mai_mai_n1006_), .B(h), .Y(mai_mai_n1343_));
  NA3        m1315(.A(mai_mai_n1343_), .B(d), .C(mai_mai_n968_), .Y(mai_mai_n1344_));
  NO2        m1316(.A(mai_mai_n1344_), .B(c), .Y(mai_mai_n1345_));
  NA3        m1317(.A(mai_mai_n1318_), .B(mai_mai_n438_), .C(f), .Y(mai_mai_n1346_));
  NO2        m1318(.A(mai_mai_n1247_), .B(mai_mai_n42_), .Y(mai_mai_n1347_));
  AOI210     m1319(.A0(mai_mai_n103_), .A1(mai_mai_n40_), .B0(mai_mai_n1347_), .Y(mai_mai_n1348_));
  NO2        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1346_), .Y(mai_mai_n1349_));
  NOi21      m1321(.An(d), .B(f), .Y(mai_mai_n1350_));
  NA2        m1322(.A(mai_mai_n1286_), .B(mai_mai_n1347_), .Y(mai_mai_n1351_));
  INV        m1323(.A(mai_mai_n1351_), .Y(mai_mai_n1352_));
  NO3        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1349_), .C(mai_mai_n1345_), .Y(mai_mai_n1353_));
  NA4        m1325(.A(mai_mai_n1353_), .B(mai_mai_n1341_), .C(mai_mai_n1328_), .D(mai_mai_n1425_), .Y(mai_mai_n1354_));
  NO3        m1326(.A(mai_mai_n1010_), .B(mai_mai_n996_), .C(mai_mai_n40_), .Y(mai_mai_n1355_));
  NO2        m1327(.A(mai_mai_n438_), .B(mai_mai_n272_), .Y(mai_mai_n1356_));
  OAI210     m1328(.A0(mai_mai_n1356_), .A1(mai_mai_n1355_), .B0(mai_mai_n1266_), .Y(mai_mai_n1357_));
  OAI210     m1329(.A0(mai_mai_n1304_), .A1(mai_mai_n1256_), .B0(mai_mai_n821_), .Y(mai_mai_n1358_));
  NO2        m1330(.A(mai_mai_n965_), .B(mai_mai_n119_), .Y(mai_mai_n1359_));
  NA2        m1331(.A(mai_mai_n1359_), .B(mai_mai_n578_), .Y(mai_mai_n1360_));
  NA3        m1332(.A(mai_mai_n1360_), .B(mai_mai_n1358_), .C(mai_mai_n1357_), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n1282_), .B(mai_mai_n1350_), .Y(mai_mai_n1362_));
  NO2        m1334(.A(mai_mai_n1362_), .B(m), .Y(mai_mai_n1363_));
  NO2        m1335(.A(mai_mai_n136_), .B(mai_mai_n165_), .Y(mai_mai_n1364_));
  OAI210     m1336(.A0(mai_mai_n1364_), .A1(mai_mai_n100_), .B0(mai_mai_n1293_), .Y(mai_mai_n1365_));
  INV        m1337(.A(mai_mai_n1365_), .Y(mai_mai_n1366_));
  NO3        m1338(.A(mai_mai_n1366_), .B(mai_mai_n1363_), .C(mai_mai_n1361_), .Y(mai_mai_n1367_));
  NO2        m1339(.A(mai_mai_n1252_), .B(e), .Y(mai_mai_n1368_));
  NA2        m1340(.A(mai_mai_n1368_), .B(mai_mai_n376_), .Y(mai_mai_n1369_));
  NA2        m1341(.A(mai_mai_n1049_), .B(mai_mai_n585_), .Y(mai_mai_n1370_));
  OR3        m1342(.A(mai_mai_n1337_), .B(mai_mai_n1129_), .C(mai_mai_n119_), .Y(mai_mai_n1371_));
  OAI220     m1343(.A0(mai_mai_n1371_), .A1(mai_mai_n1369_), .B0(mai_mai_n1370_), .B1(mai_mai_n415_), .Y(mai_mai_n1372_));
  INV        m1344(.A(mai_mai_n1372_), .Y(mai_mai_n1373_));
  NO2        m1345(.A(mai_mai_n165_), .B(c), .Y(mai_mai_n1374_));
  OAI210     m1346(.A0(mai_mai_n1374_), .A1(mai_mai_n1368_), .B0(mai_mai_n163_), .Y(mai_mai_n1375_));
  AOI220     m1347(.A0(mai_mai_n1375_), .A1(mai_mai_n998_), .B0(mai_mai_n504_), .B1(mai_mai_n336_), .Y(mai_mai_n1376_));
  NA2        m1348(.A(mai_mai_n510_), .B(g), .Y(mai_mai_n1377_));
  AOI210     m1349(.A0(mai_mai_n1377_), .A1(mai_mai_n1278_), .B0(mai_mai_n1342_), .Y(mai_mai_n1378_));
  NO2        m1350(.A(mai_mai_n1307_), .B(f), .Y(mai_mai_n1379_));
  NO2        m1351(.A(mai_mai_n1378_), .B(mai_mai_n196_), .Y(mai_mai_n1380_));
  NA2        m1352(.A(mai_mai_n1379_), .B(mai_mai_n1263_), .Y(mai_mai_n1381_));
  OAI220     m1353(.A0(mai_mai_n1381_), .A1(mai_mai_n47_), .B0(mai_mai_n1429_), .B1(mai_mai_n158_), .Y(mai_mai_n1382_));
  NA4        m1354(.A(mai_mai_n1019_), .B(mai_mai_n1016_), .C(mai_mai_n202_), .D(mai_mai_n63_), .Y(mai_mai_n1383_));
  NA2        m1355(.A(mai_mai_n1257_), .B(mai_mai_n166_), .Y(mai_mai_n1384_));
  NO2        m1356(.A(mai_mai_n47_), .B(l), .Y(mai_mai_n1385_));
  OAI210     m1357(.A0(mai_mai_n1307_), .A1(mai_mai_n801_), .B0(mai_mai_n454_), .Y(mai_mai_n1386_));
  OAI210     m1358(.A0(mai_mai_n1386_), .A1(mai_mai_n1022_), .B0(mai_mai_n1385_), .Y(mai_mai_n1387_));
  NO2        m1359(.A(mai_mai_n236_), .B(g), .Y(mai_mai_n1388_));
  NO2        m1360(.A(m), .B(i), .Y(mai_mai_n1389_));
  BUFFER     m1361(.A(mai_mai_n1389_), .Y(mai_mai_n1390_));
  AOI220     m1362(.A0(mai_mai_n1390_), .A1(mai_mai_n1280_), .B0(mai_mai_n997_), .B1(mai_mai_n1388_), .Y(mai_mai_n1391_));
  NA4        m1363(.A(mai_mai_n1391_), .B(mai_mai_n1387_), .C(mai_mai_n1384_), .D(mai_mai_n1383_), .Y(mai_mai_n1392_));
  NO4        m1364(.A(mai_mai_n1392_), .B(mai_mai_n1382_), .C(mai_mai_n1380_), .D(mai_mai_n1376_), .Y(mai_mai_n1393_));
  NA3        m1365(.A(mai_mai_n1393_), .B(mai_mai_n1373_), .C(mai_mai_n1367_), .Y(mai_mai_n1394_));
  NA3        m1366(.A(mai_mai_n896_), .B(mai_mai_n125_), .C(mai_mai_n45_), .Y(mai_mai_n1395_));
  AOI210     m1367(.A0(mai_mai_n133_), .A1(c), .B0(mai_mai_n1395_), .Y(mai_mai_n1396_));
  INV        m1368(.A(mai_mai_n169_), .Y(mai_mai_n1397_));
  NA2        m1369(.A(mai_mai_n1397_), .B(mai_mai_n1343_), .Y(mai_mai_n1398_));
  INV        m1370(.A(mai_mai_n1398_), .Y(mai_mai_n1399_));
  NO2        m1371(.A(mai_mai_n1399_), .B(mai_mai_n1396_), .Y(mai_mai_n1400_));
  NOi21      m1372(.An(mai_mai_n1257_), .B(e), .Y(mai_mai_n1401_));
  AN2        m1373(.A(mai_mai_n1019_), .B(mai_mai_n1004_), .Y(mai_mai_n1402_));
  AOI220     m1374(.A0(mai_mai_n1389_), .A1(mai_mai_n592_), .B0(mai_mai_n1426_), .B1(mai_mai_n144_), .Y(mai_mai_n1403_));
  NOi31      m1375(.An(mai_mai_n30_), .B(mai_mai_n1403_), .C(n), .Y(mai_mai_n1404_));
  AOI210     m1376(.A0(mai_mai_n1402_), .A1(mai_mai_n1089_), .B0(mai_mai_n1404_), .Y(mai_mai_n1405_));
  NO2        m1377(.A(mai_mai_n1346_), .B(mai_mai_n64_), .Y(mai_mai_n1406_));
  NA2        m1378(.A(mai_mai_n57_), .B(a), .Y(mai_mai_n1407_));
  NO2        m1379(.A(mai_mai_n1262_), .B(mai_mai_n108_), .Y(mai_mai_n1408_));
  OAI220     m1380(.A0(mai_mai_n1408_), .A1(mai_mai_n1301_), .B0(mai_mai_n1313_), .B1(mai_mai_n1407_), .Y(mai_mai_n1409_));
  NO2        m1381(.A(mai_mai_n1409_), .B(mai_mai_n1406_), .Y(mai_mai_n1410_));
  NA4        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1405_), .C(mai_mai_n1431_), .D(mai_mai_n1400_), .Y(mai_mai_n1411_));
  OR4        m1383(.A(mai_mai_n1411_), .B(mai_mai_n1394_), .C(mai_mai_n1354_), .D(mai_mai_n1317_), .Y(mai04));
  NOi31      m1384(.An(mai_mai_n1304_), .B(mai_mai_n1305_), .C(mai_mai_n970_), .Y(mai_mai_n1413_));
  INV        m1385(.A(mai_mai_n767_), .Y(mai_mai_n1414_));
  NO3        m1386(.A(mai_mai_n1414_), .B(mai_mai_n960_), .C(mai_mai_n455_), .Y(mai_mai_n1415_));
  OR3        m1387(.A(mai_mai_n1415_), .B(mai_mai_n1413_), .C(mai_mai_n987_), .Y(mai_mai_n1416_));
  NO3        m1388(.A(mai_mai_n1263_), .B(mai_mai_n86_), .C(k), .Y(mai_mai_n1417_));
  AOI210     m1389(.A0(mai_mai_n1417_), .A1(mai_mai_n981_), .B0(mai_mai_n1106_), .Y(mai_mai_n1418_));
  NA2        m1390(.A(mai_mai_n1418_), .B(mai_mai_n1133_), .Y(mai_mai_n1419_));
  NO4        m1391(.A(mai_mai_n1419_), .B(mai_mai_n1416_), .C(mai_mai_n995_), .D(mai_mai_n975_), .Y(mai_mai_n1420_));
  NA4        m1392(.A(mai_mai_n1420_), .B(mai_mai_n1051_), .C(mai_mai_n1036_), .D(mai_mai_n1025_), .Y(mai05));
  INV        m1393(.A(m), .Y(mai_mai_n1424_));
  INV        m1394(.A(mai_mai_n1321_), .Y(mai_mai_n1425_));
  INV        m1395(.A(j), .Y(mai_mai_n1426_));
  INV        m1396(.A(i), .Y(mai_mai_n1427_));
  INV        m1397(.A(k), .Y(mai_mai_n1428_));
  INV        m1398(.A(mai_mai_n95_), .Y(mai_mai_n1429_));
  INV        m1399(.A(k), .Y(mai_mai_n1430_));
  INV        m1400(.A(mai_mai_n1401_), .Y(mai_mai_n1431_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi31      u0013(.An(n), .B(m), .C(l), .Y(men_men_n42_));
  INV        u0014(.A(i), .Y(men_men_n43_));
  AN2        u0015(.A(h), .B(g), .Y(men_men_n44_));
  NA2        u0016(.A(men_men_n44_), .B(men_men_n43_), .Y(men_men_n45_));
  NO2        u0017(.A(men_men_n45_), .B(men_men_n42_), .Y(men_men_n46_));
  NAi21      u0018(.An(n), .B(m), .Y(men_men_n47_));
  NOi32      u0019(.An(k), .Bn(h), .C(l), .Y(men_men_n48_));
  NOi32      u0020(.An(k), .Bn(h), .C(g), .Y(men_men_n49_));
  INV        u0021(.A(men_men_n49_), .Y(men_men_n50_));
  NO2        u0022(.A(men_men_n50_), .B(men_men_n47_), .Y(men_men_n51_));
  NO3        u0023(.A(men_men_n51_), .B(men_men_n46_), .C(men_men_n39_), .Y(men_men_n52_));
  AOI210     u0024(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n53_));
  INV        u0025(.A(c), .Y(men_men_n54_));
  NA2        u0026(.A(e), .B(b), .Y(men_men_n55_));
  NO2        u0027(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  INV        u0028(.A(d), .Y(men_men_n57_));
  NA3        u0029(.A(g), .B(men_men_n57_), .C(a), .Y(men_men_n58_));
  NAi21      u0030(.An(i), .B(h), .Y(men_men_n59_));
  NAi31      u0031(.An(i), .B(l), .C(j), .Y(men_men_n60_));
  NO2        u0032(.A(men_men_n59_), .B(men_men_n42_), .Y(men_men_n61_));
  NAi31      u0033(.An(men_men_n58_), .B(men_men_n61_), .C(men_men_n56_), .Y(men_men_n62_));
  NAi41      u0034(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n63_));
  NA2        u0035(.A(g), .B(f), .Y(men_men_n64_));
  NO2        u0036(.A(men_men_n64_), .B(men_men_n63_), .Y(men_men_n65_));
  NAi21      u0037(.An(i), .B(j), .Y(men_men_n66_));
  NAi32      u0038(.An(n), .Bn(k), .C(m), .Y(men_men_n67_));
  NO2        u0039(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n68_));
  NAi31      u0040(.An(l), .B(m), .C(k), .Y(men_men_n69_));
  NAi21      u0041(.An(e), .B(h), .Y(men_men_n70_));
  NAi41      u0042(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n71_));
  NA2        u0043(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n72_));
  INV        u0044(.A(m), .Y(men_men_n73_));
  NOi21      u0045(.An(k), .B(l), .Y(men_men_n74_));
  NA2        u0046(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n75_));
  AN4        u0047(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n76_));
  NOi31      u0048(.An(h), .B(g), .C(f), .Y(men_men_n77_));
  NA2        u0049(.A(men_men_n77_), .B(men_men_n76_), .Y(men_men_n78_));
  NAi32      u0050(.An(m), .Bn(k), .C(j), .Y(men_men_n79_));
  NOi32      u0051(.An(h), .Bn(g), .C(f), .Y(men_men_n80_));
  OR2        u0052(.A(men_men_n78_), .B(men_men_n75_), .Y(men_men_n81_));
  NA3        u0053(.A(men_men_n81_), .B(men_men_n72_), .C(men_men_n62_), .Y(men_men_n82_));
  INV        u0054(.A(n), .Y(men_men_n83_));
  NOi32      u0055(.An(e), .Bn(b), .C(d), .Y(men_men_n84_));
  NA2        u0056(.A(men_men_n84_), .B(men_men_n83_), .Y(men_men_n85_));
  INV        u0057(.A(j), .Y(men_men_n86_));
  AN3        u0058(.A(m), .B(k), .C(i), .Y(men_men_n87_));
  NA3        u0059(.A(men_men_n87_), .B(men_men_n86_), .C(g), .Y(men_men_n88_));
  NO2        u0060(.A(men_men_n88_), .B(f), .Y(men_men_n89_));
  NAi32      u0061(.An(g), .Bn(f), .C(h), .Y(men_men_n90_));
  NAi31      u0062(.An(j), .B(m), .C(l), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  NA2        u0064(.A(m), .B(l), .Y(men_men_n93_));
  NAi31      u0065(.An(k), .B(j), .C(g), .Y(men_men_n94_));
  NO3        u0066(.A(men_men_n94_), .B(men_men_n93_), .C(f), .Y(men_men_n95_));
  AN2        u0067(.A(j), .B(g), .Y(men_men_n96_));
  NOi32      u0068(.An(m), .Bn(l), .C(i), .Y(men_men_n97_));
  NOi21      u0069(.An(g), .B(i), .Y(men_men_n98_));
  NOi32      u0070(.An(m), .Bn(j), .C(k), .Y(men_men_n99_));
  AOI220     u0071(.A0(men_men_n99_), .A1(men_men_n98_), .B0(men_men_n97_), .B1(men_men_n96_), .Y(men_men_n100_));
  NO2        u0072(.A(men_men_n100_), .B(f), .Y(men_men_n101_));
  NO4        u0073(.A(men_men_n101_), .B(men_men_n95_), .C(men_men_n92_), .D(men_men_n89_), .Y(men_men_n102_));
  NAi41      u0074(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n103_));
  AN2        u0075(.A(e), .B(b), .Y(men_men_n104_));
  NOi21      u0076(.An(g), .B(f), .Y(men_men_n105_));
  NOi21      u0077(.An(i), .B(h), .Y(men_men_n106_));
  NA3        u0078(.A(men_men_n106_), .B(men_men_n105_), .C(men_men_n36_), .Y(men_men_n107_));
  INV        u0079(.A(a), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n104_), .B(men_men_n108_), .Y(men_men_n109_));
  INV        u0081(.A(l), .Y(men_men_n110_));
  NOi21      u0082(.An(m), .B(n), .Y(men_men_n111_));
  AN2        u0083(.A(k), .B(h), .Y(men_men_n112_));
  NO2        u0084(.A(men_men_n107_), .B(men_men_n85_), .Y(men_men_n113_));
  INV        u0085(.A(b), .Y(men_men_n114_));
  NA2        u0086(.A(l), .B(j), .Y(men_men_n115_));
  AN2        u0087(.A(k), .B(i), .Y(men_men_n116_));
  NA2        u0088(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NA2        u0089(.A(g), .B(e), .Y(men_men_n118_));
  NOi32      u0090(.An(c), .Bn(a), .C(d), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n111_), .Y(men_men_n120_));
  INV        u0092(.A(men_men_n113_), .Y(men_men_n121_));
  OAI210     u0093(.A0(men_men_n102_), .A1(men_men_n85_), .B0(men_men_n121_), .Y(men_men_n122_));
  NOi31      u0094(.An(k), .B(m), .C(j), .Y(men_men_n123_));
  NA3        u0095(.A(men_men_n123_), .B(men_men_n77_), .C(men_men_n76_), .Y(men_men_n124_));
  NOi31      u0096(.An(k), .B(m), .C(i), .Y(men_men_n125_));
  NA3        u0097(.A(men_men_n125_), .B(men_men_n80_), .C(men_men_n76_), .Y(men_men_n126_));
  NA2        u0098(.A(men_men_n126_), .B(men_men_n124_), .Y(men_men_n127_));
  NOi32      u0099(.An(f), .Bn(b), .C(e), .Y(men_men_n128_));
  NAi21      u0100(.An(g), .B(h), .Y(men_men_n129_));
  NAi21      u0101(.An(m), .B(n), .Y(men_men_n130_));
  NAi21      u0102(.An(j), .B(k), .Y(men_men_n131_));
  NO3        u0103(.A(men_men_n131_), .B(men_men_n130_), .C(men_men_n129_), .Y(men_men_n132_));
  NAi41      u0104(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n133_));
  NAi31      u0105(.An(j), .B(k), .C(h), .Y(men_men_n134_));
  NO3        u0106(.A(men_men_n134_), .B(men_men_n133_), .C(men_men_n130_), .Y(men_men_n135_));
  AOI210     u0107(.A0(men_men_n132_), .A1(men_men_n128_), .B0(men_men_n135_), .Y(men_men_n136_));
  NO2        u0108(.A(k), .B(j), .Y(men_men_n137_));
  NO2        u0109(.A(men_men_n137_), .B(men_men_n130_), .Y(men_men_n138_));
  AN2        u0110(.A(k), .B(j), .Y(men_men_n139_));
  NAi21      u0111(.An(c), .B(b), .Y(men_men_n140_));
  NA2        u0112(.A(f), .B(d), .Y(men_men_n141_));
  NO3        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n129_), .Y(men_men_n142_));
  NAi31      u0114(.An(f), .B(e), .C(b), .Y(men_men_n143_));
  NA2        u0115(.A(men_men_n142_), .B(men_men_n138_), .Y(men_men_n144_));
  NA2        u0116(.A(d), .B(b), .Y(men_men_n145_));
  NAi21      u0117(.An(e), .B(f), .Y(men_men_n146_));
  NO2        u0118(.A(men_men_n146_), .B(men_men_n145_), .Y(men_men_n147_));
  NA2        u0119(.A(b), .B(a), .Y(men_men_n148_));
  NAi21      u0120(.An(e), .B(g), .Y(men_men_n149_));
  NAi21      u0121(.An(c), .B(d), .Y(men_men_n150_));
  NAi31      u0122(.An(l), .B(k), .C(h), .Y(men_men_n151_));
  NO2        u0123(.A(men_men_n130_), .B(men_men_n151_), .Y(men_men_n152_));
  NA2        u0124(.A(men_men_n152_), .B(men_men_n147_), .Y(men_men_n153_));
  NAi41      u0125(.An(men_men_n127_), .B(men_men_n153_), .C(men_men_n144_), .D(men_men_n136_), .Y(men_men_n154_));
  NAi31      u0126(.An(e), .B(f), .C(b), .Y(men_men_n155_));
  NOi21      u0127(.An(g), .B(d), .Y(men_men_n156_));
  NO2        u0128(.A(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  NOi21      u0129(.An(h), .B(i), .Y(men_men_n158_));
  NOi21      u0130(.An(k), .B(m), .Y(men_men_n159_));
  NA3        u0131(.A(men_men_n159_), .B(men_men_n158_), .C(n), .Y(men_men_n160_));
  NOi21      u0132(.An(h), .B(g), .Y(men_men_n161_));
  NO2        u0133(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n162_));
  NAi31      u0134(.An(l), .B(j), .C(h), .Y(men_men_n163_));
  NO2        u0135(.A(men_men_n163_), .B(men_men_n47_), .Y(men_men_n164_));
  NA2        u0136(.A(men_men_n164_), .B(men_men_n65_), .Y(men_men_n165_));
  NOi32      u0137(.An(n), .Bn(k), .C(m), .Y(men_men_n166_));
  NA2        u0138(.A(l), .B(i), .Y(men_men_n167_));
  INV        u0139(.A(men_men_n165_), .Y(men_men_n168_));
  NAi31      u0140(.An(d), .B(f), .C(c), .Y(men_men_n169_));
  NAi31      u0141(.An(e), .B(f), .C(c), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NA2        u0143(.A(j), .B(h), .Y(men_men_n172_));
  OR3        u0144(.A(n), .B(m), .C(k), .Y(men_men_n173_));
  NO2        u0145(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NAi32      u0146(.An(m), .Bn(k), .C(n), .Y(men_men_n175_));
  NO2        u0147(.A(men_men_n175_), .B(men_men_n172_), .Y(men_men_n176_));
  AOI220     u0148(.A0(men_men_n176_), .A1(men_men_n157_), .B0(men_men_n174_), .B1(men_men_n171_), .Y(men_men_n177_));
  NO2        u0149(.A(n), .B(m), .Y(men_men_n178_));
  NA2        u0150(.A(men_men_n178_), .B(men_men_n48_), .Y(men_men_n179_));
  NAi21      u0151(.An(f), .B(e), .Y(men_men_n180_));
  NA2        u0152(.A(d), .B(c), .Y(men_men_n181_));
  NAi31      u0153(.An(m), .B(n), .C(b), .Y(men_men_n182_));
  NA2        u0154(.A(k), .B(i), .Y(men_men_n183_));
  NAi21      u0155(.An(h), .B(f), .Y(men_men_n184_));
  NO2        u0156(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  NO2        u0157(.A(men_men_n182_), .B(men_men_n150_), .Y(men_men_n186_));
  NA2        u0158(.A(men_men_n186_), .B(men_men_n185_), .Y(men_men_n187_));
  NOi32      u0159(.An(f), .Bn(c), .C(d), .Y(men_men_n188_));
  NOi32      u0160(.An(f), .Bn(c), .C(e), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NO3        u0162(.A(n), .B(m), .C(j), .Y(men_men_n191_));
  NA2        u0163(.A(men_men_n191_), .B(men_men_n112_), .Y(men_men_n192_));
  AO210      u0164(.A0(men_men_n192_), .A1(men_men_n179_), .B0(men_men_n190_), .Y(men_men_n193_));
  NA3        u0165(.A(men_men_n193_), .B(men_men_n187_), .C(men_men_n177_), .Y(men_men_n194_));
  OR3        u0166(.A(men_men_n194_), .B(men_men_n168_), .C(men_men_n154_), .Y(men_men_n195_));
  NO4        u0167(.A(men_men_n195_), .B(men_men_n122_), .C(men_men_n82_), .D(men_men_n53_), .Y(men_men_n196_));
  NA3        u0168(.A(m), .B(men_men_n110_), .C(j), .Y(men_men_n197_));
  NAi31      u0169(.An(n), .B(h), .C(g), .Y(men_men_n198_));
  NO2        u0170(.A(men_men_n198_), .B(men_men_n197_), .Y(men_men_n199_));
  NOi32      u0171(.An(m), .Bn(k), .C(l), .Y(men_men_n200_));
  NA3        u0172(.A(men_men_n200_), .B(men_men_n86_), .C(g), .Y(men_men_n201_));
  AN2        u0173(.A(i), .B(g), .Y(men_men_n202_));
  NA3        u0174(.A(men_men_n74_), .B(men_men_n202_), .C(men_men_n111_), .Y(men_men_n203_));
  INV        u0175(.A(men_men_n199_), .Y(men_men_n204_));
  NAi41      u0176(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n205_));
  INV        u0177(.A(men_men_n205_), .Y(men_men_n206_));
  INV        u0178(.A(f), .Y(men_men_n207_));
  INV        u0179(.A(g), .Y(men_men_n208_));
  NOi31      u0180(.An(i), .B(j), .C(h), .Y(men_men_n209_));
  NOi21      u0181(.An(l), .B(m), .Y(men_men_n210_));
  NA2        u0182(.A(men_men_n210_), .B(men_men_n209_), .Y(men_men_n211_));
  NO3        u0183(.A(men_men_n211_), .B(men_men_n208_), .C(men_men_n207_), .Y(men_men_n212_));
  NA2        u0184(.A(men_men_n212_), .B(men_men_n206_), .Y(men_men_n213_));
  OAI210     u0185(.A0(men_men_n204_), .A1(men_men_n32_), .B0(men_men_n213_), .Y(men_men_n214_));
  NOi21      u0186(.An(n), .B(m), .Y(men_men_n215_));
  NOi32      u0187(.An(l), .Bn(i), .C(j), .Y(men_men_n216_));
  NA2        u0188(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NAi21      u0189(.An(j), .B(h), .Y(men_men_n218_));
  XN2        u0190(.A(i), .B(h), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n220_));
  NOi31      u0192(.An(k), .B(n), .C(m), .Y(men_men_n221_));
  NOi31      u0193(.An(men_men_n221_), .B(men_men_n181_), .C(men_men_n180_), .Y(men_men_n222_));
  NA2        u0194(.A(men_men_n222_), .B(men_men_n220_), .Y(men_men_n223_));
  NAi31      u0195(.An(f), .B(e), .C(c), .Y(men_men_n224_));
  NO4        u0196(.A(men_men_n224_), .B(men_men_n173_), .C(men_men_n172_), .D(men_men_n57_), .Y(men_men_n225_));
  NA4        u0197(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n226_));
  NAi32      u0198(.An(m), .Bn(i), .C(k), .Y(men_men_n227_));
  NO3        u0199(.A(men_men_n227_), .B(men_men_n90_), .C(men_men_n226_), .Y(men_men_n228_));
  INV        u0200(.A(k), .Y(men_men_n229_));
  NO2        u0201(.A(men_men_n228_), .B(men_men_n225_), .Y(men_men_n230_));
  NAi21      u0202(.An(n), .B(a), .Y(men_men_n231_));
  NO2        u0203(.A(men_men_n231_), .B(men_men_n145_), .Y(men_men_n232_));
  NAi41      u0204(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n233_));
  NO2        u0205(.A(men_men_n233_), .B(e), .Y(men_men_n234_));
  NO3        u0206(.A(men_men_n146_), .B(men_men_n94_), .C(men_men_n93_), .Y(men_men_n235_));
  OAI210     u0207(.A0(men_men_n235_), .A1(men_men_n234_), .B0(men_men_n232_), .Y(men_men_n236_));
  AN3        u0208(.A(men_men_n236_), .B(men_men_n230_), .C(men_men_n223_), .Y(men_men_n237_));
  OR2        u0209(.A(h), .B(g), .Y(men_men_n238_));
  NO2        u0210(.A(men_men_n238_), .B(men_men_n103_), .Y(men_men_n239_));
  NA2        u0211(.A(men_men_n239_), .B(men_men_n128_), .Y(men_men_n240_));
  NAi41      u0212(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n207_), .Y(men_men_n242_));
  NA2        u0214(.A(men_men_n159_), .B(men_men_n106_), .Y(men_men_n243_));
  NAi21      u0215(.An(men_men_n243_), .B(men_men_n242_), .Y(men_men_n244_));
  NO2        u0216(.A(n), .B(a), .Y(men_men_n245_));
  NAi31      u0217(.An(men_men_n233_), .B(men_men_n245_), .C(men_men_n104_), .Y(men_men_n246_));
  AN2        u0218(.A(men_men_n246_), .B(men_men_n244_), .Y(men_men_n247_));
  NAi21      u0219(.An(h), .B(i), .Y(men_men_n248_));
  NA2        u0220(.A(men_men_n178_), .B(k), .Y(men_men_n249_));
  NO2        u0221(.A(men_men_n249_), .B(men_men_n248_), .Y(men_men_n250_));
  NA2        u0222(.A(men_men_n250_), .B(men_men_n188_), .Y(men_men_n251_));
  NA3        u0223(.A(men_men_n251_), .B(men_men_n247_), .C(men_men_n240_), .Y(men_men_n252_));
  NOi21      u0224(.An(g), .B(e), .Y(men_men_n253_));
  NO2        u0225(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n254_));
  NA2        u0226(.A(men_men_n254_), .B(men_men_n253_), .Y(men_men_n255_));
  NOi32      u0227(.An(l), .Bn(j), .C(i), .Y(men_men_n256_));
  AOI210     u0228(.A0(men_men_n74_), .A1(men_men_n86_), .B0(men_men_n256_), .Y(men_men_n257_));
  NO2        u0229(.A(men_men_n248_), .B(men_men_n42_), .Y(men_men_n258_));
  NAi21      u0230(.An(f), .B(g), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n63_), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n67_), .B(men_men_n115_), .Y(men_men_n261_));
  AOI220     u0233(.A0(men_men_n261_), .A1(men_men_n260_), .B0(men_men_n258_), .B1(men_men_n65_), .Y(men_men_n262_));
  OAI210     u0234(.A0(men_men_n257_), .A1(men_men_n255_), .B0(men_men_n262_), .Y(men_men_n263_));
  NO3        u0235(.A(men_men_n131_), .B(men_men_n47_), .C(men_men_n43_), .Y(men_men_n264_));
  NOi41      u0236(.An(men_men_n237_), .B(men_men_n263_), .C(men_men_n252_), .D(men_men_n214_), .Y(men_men_n265_));
  NO3        u0237(.A(men_men_n199_), .B(men_men_n46_), .C(men_men_n39_), .Y(men_men_n266_));
  NO2        u0238(.A(men_men_n266_), .B(men_men_n109_), .Y(men_men_n267_));
  NAi21      u0239(.An(h), .B(g), .Y(men_men_n268_));
  OR4        u0240(.A(men_men_n268_), .B(men_men_n1484_), .C(men_men_n217_), .D(e), .Y(men_men_n269_));
  NAi31      u0241(.An(g), .B(k), .C(h), .Y(men_men_n270_));
  NAi31      u0242(.An(e), .B(d), .C(a), .Y(men_men_n271_));
  NA4        u0243(.A(men_men_n159_), .B(men_men_n80_), .C(men_men_n76_), .D(men_men_n115_), .Y(men_men_n272_));
  NA3        u0244(.A(men_men_n159_), .B(men_men_n158_), .C(men_men_n83_), .Y(men_men_n273_));
  NO2        u0245(.A(men_men_n273_), .B(men_men_n190_), .Y(men_men_n274_));
  NOi21      u0246(.An(men_men_n272_), .B(men_men_n274_), .Y(men_men_n275_));
  NA3        u0247(.A(e), .B(c), .C(b), .Y(men_men_n276_));
  NO2        u0248(.A(men_men_n58_), .B(men_men_n276_), .Y(men_men_n277_));
  NAi32      u0249(.An(k), .Bn(i), .C(j), .Y(men_men_n278_));
  NAi31      u0250(.An(h), .B(l), .C(i), .Y(men_men_n279_));
  NA3        u0251(.A(men_men_n279_), .B(men_men_n278_), .C(men_men_n163_), .Y(men_men_n280_));
  NOi21      u0252(.An(men_men_n280_), .B(men_men_n47_), .Y(men_men_n281_));
  OAI210     u0253(.A0(men_men_n260_), .A1(men_men_n277_), .B0(men_men_n281_), .Y(men_men_n282_));
  NAi21      u0254(.An(l), .B(k), .Y(men_men_n283_));
  NO2        u0255(.A(men_men_n283_), .B(men_men_n47_), .Y(men_men_n284_));
  NOi21      u0256(.An(l), .B(j), .Y(men_men_n285_));
  NA2        u0257(.A(men_men_n161_), .B(men_men_n285_), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n116_), .B(men_men_n115_), .C(g), .Y(men_men_n287_));
  OR3        u0259(.A(men_men_n71_), .B(men_men_n73_), .C(e), .Y(men_men_n288_));
  AOI210     u0260(.A0(men_men_n287_), .A1(men_men_n286_), .B0(men_men_n288_), .Y(men_men_n289_));
  INV        u0261(.A(men_men_n289_), .Y(men_men_n290_));
  NAi32      u0262(.An(j), .Bn(h), .C(i), .Y(men_men_n291_));
  NAi21      u0263(.An(m), .B(l), .Y(men_men_n292_));
  NO3        u0264(.A(men_men_n292_), .B(men_men_n291_), .C(men_men_n83_), .Y(men_men_n293_));
  NA2        u0265(.A(h), .B(g), .Y(men_men_n294_));
  NA2        u0266(.A(men_men_n166_), .B(men_men_n43_), .Y(men_men_n295_));
  NO2        u0267(.A(men_men_n295_), .B(men_men_n294_), .Y(men_men_n296_));
  NA2        u0268(.A(men_men_n296_), .B(men_men_n162_), .Y(men_men_n297_));
  NA4        u0269(.A(men_men_n297_), .B(men_men_n290_), .C(men_men_n282_), .D(men_men_n275_), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n143_), .B(d), .Y(men_men_n299_));
  NA2        u0271(.A(men_men_n299_), .B(men_men_n51_), .Y(men_men_n300_));
  NAi32      u0272(.An(n), .Bn(m), .C(l), .Y(men_men_n301_));
  NO2        u0273(.A(men_men_n120_), .B(men_men_n114_), .Y(men_men_n302_));
  NAi31      u0274(.An(k), .B(l), .C(j), .Y(men_men_n303_));
  OAI210     u0275(.A0(men_men_n283_), .A1(j), .B0(men_men_n303_), .Y(men_men_n304_));
  NOi21      u0276(.An(men_men_n304_), .B(men_men_n118_), .Y(men_men_n305_));
  NA2        u0277(.A(men_men_n305_), .B(men_men_n302_), .Y(men_men_n306_));
  NA2        u0278(.A(men_men_n306_), .B(men_men_n300_), .Y(men_men_n307_));
  NO4        u0279(.A(men_men_n307_), .B(men_men_n298_), .C(men_men_n1482_), .D(men_men_n267_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n250_), .B(men_men_n189_), .Y(men_men_n309_));
  NAi21      u0281(.An(m), .B(k), .Y(men_men_n310_));
  NAi41      u0282(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n311_));
  NAi31      u0283(.An(i), .B(l), .C(h), .Y(men_men_n312_));
  NO4        u0284(.A(men_men_n312_), .B(men_men_n149_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n313_));
  NA2        u0285(.A(e), .B(c), .Y(men_men_n314_));
  NO3        u0286(.A(men_men_n314_), .B(n), .C(d), .Y(men_men_n315_));
  NOi21      u0287(.An(f), .B(h), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n316_), .B(men_men_n116_), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n317_), .B(men_men_n208_), .Y(men_men_n318_));
  NAi31      u0290(.An(d), .B(e), .C(b), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n130_), .B(men_men_n319_), .Y(men_men_n320_));
  NA2        u0292(.A(men_men_n320_), .B(men_men_n318_), .Y(men_men_n321_));
  NAi31      u0293(.An(men_men_n313_), .B(men_men_n321_), .C(men_men_n309_), .Y(men_men_n322_));
  NO4        u0294(.A(men_men_n311_), .B(men_men_n79_), .C(men_men_n70_), .D(men_men_n208_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n245_), .B(men_men_n104_), .Y(men_men_n324_));
  OR2        u0296(.A(men_men_n324_), .B(men_men_n201_), .Y(men_men_n325_));
  NOi31      u0297(.An(l), .B(n), .C(m), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n326_), .B(men_men_n209_), .Y(men_men_n327_));
  NO2        u0299(.A(men_men_n327_), .B(men_men_n190_), .Y(men_men_n328_));
  NAi32      u0300(.An(men_men_n328_), .Bn(men_men_n323_), .C(men_men_n325_), .Y(men_men_n329_));
  NAi32      u0301(.An(m), .Bn(j), .C(k), .Y(men_men_n330_));
  NAi41      u0302(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n205_), .B(men_men_n331_), .Y(men_men_n332_));
  NOi31      u0304(.An(j), .B(m), .C(k), .Y(men_men_n333_));
  NO2        u0305(.A(men_men_n123_), .B(men_men_n333_), .Y(men_men_n334_));
  AN3        u0306(.A(h), .B(g), .C(f), .Y(men_men_n335_));
  NAi31      u0307(.An(men_men_n334_), .B(men_men_n335_), .C(men_men_n332_), .Y(men_men_n336_));
  NOi32      u0308(.An(m), .Bn(j), .C(l), .Y(men_men_n337_));
  NO2        u0309(.A(men_men_n292_), .B(men_men_n291_), .Y(men_men_n338_));
  NO2        u0310(.A(men_men_n211_), .B(g), .Y(men_men_n339_));
  NO2        u0311(.A(men_men_n155_), .B(men_men_n83_), .Y(men_men_n340_));
  AOI220     u0312(.A0(men_men_n340_), .A1(men_men_n339_), .B0(men_men_n242_), .B1(men_men_n338_), .Y(men_men_n341_));
  INV        u0313(.A(men_men_n227_), .Y(men_men_n342_));
  NA3        u0314(.A(men_men_n342_), .B(men_men_n335_), .C(men_men_n206_), .Y(men_men_n343_));
  NA3        u0315(.A(men_men_n343_), .B(men_men_n341_), .C(men_men_n336_), .Y(men_men_n344_));
  NA3        u0316(.A(h), .B(g), .C(f), .Y(men_men_n345_));
  NO2        u0317(.A(men_men_n345_), .B(men_men_n75_), .Y(men_men_n346_));
  NA2        u0318(.A(men_men_n331_), .B(men_men_n205_), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NOi32      u0320(.An(j), .Bn(g), .C(i), .Y(men_men_n349_));
  NA3        u0321(.A(men_men_n349_), .B(men_men_n283_), .C(men_men_n111_), .Y(men_men_n350_));
  AO210      u0322(.A0(men_men_n109_), .A1(men_men_n32_), .B0(men_men_n350_), .Y(men_men_n351_));
  NOi32      u0323(.An(e), .Bn(b), .C(a), .Y(men_men_n352_));
  AN2        u0324(.A(l), .B(j), .Y(men_men_n353_));
  INV        u0325(.A(men_men_n310_), .Y(men_men_n354_));
  NO3        u0326(.A(men_men_n311_), .B(men_men_n70_), .C(men_men_n208_), .Y(men_men_n355_));
  NA2        u0327(.A(men_men_n203_), .B(men_men_n35_), .Y(men_men_n356_));
  AOI220     u0328(.A0(men_men_n356_), .A1(men_men_n352_), .B0(men_men_n355_), .B1(men_men_n354_), .Y(men_men_n357_));
  NO2        u0329(.A(men_men_n319_), .B(n), .Y(men_men_n358_));
  NA2        u0330(.A(men_men_n202_), .B(k), .Y(men_men_n359_));
  NA3        u0331(.A(m), .B(men_men_n110_), .C(men_men_n207_), .Y(men_men_n360_));
  NO2        u0332(.A(men_men_n360_), .B(men_men_n359_), .Y(men_men_n361_));
  NAi41      u0333(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n362_));
  NA2        u0334(.A(men_men_n49_), .B(men_men_n111_), .Y(men_men_n363_));
  NA2        u0335(.A(men_men_n361_), .B(men_men_n358_), .Y(men_men_n364_));
  NA4        u0336(.A(men_men_n364_), .B(men_men_n357_), .C(men_men_n351_), .D(men_men_n348_), .Y(men_men_n365_));
  NO4        u0337(.A(men_men_n365_), .B(men_men_n344_), .C(men_men_n329_), .D(men_men_n322_), .Y(men_men_n366_));
  NA4        u0338(.A(men_men_n366_), .B(men_men_n308_), .C(men_men_n265_), .D(men_men_n196_), .Y(men10));
  NA3        u0339(.A(m), .B(k), .C(i), .Y(men_men_n368_));
  NO3        u0340(.A(men_men_n368_), .B(j), .C(men_men_n208_), .Y(men_men_n369_));
  NOi21      u0341(.An(e), .B(f), .Y(men_men_n370_));
  NO4        u0342(.A(men_men_n150_), .B(men_men_n370_), .C(n), .D(men_men_n108_), .Y(men_men_n371_));
  NAi31      u0343(.An(b), .B(f), .C(c), .Y(men_men_n372_));
  INV        u0344(.A(men_men_n372_), .Y(men_men_n373_));
  NOi32      u0345(.An(k), .Bn(h), .C(j), .Y(men_men_n374_));
  NA2        u0346(.A(men_men_n374_), .B(men_men_n215_), .Y(men_men_n375_));
  NA2        u0347(.A(men_men_n160_), .B(men_men_n375_), .Y(men_men_n376_));
  AOI220     u0348(.A0(men_men_n376_), .A1(men_men_n373_), .B0(men_men_n371_), .B1(men_men_n369_), .Y(men_men_n377_));
  AN2        u0349(.A(j), .B(h), .Y(men_men_n378_));
  NO3        u0350(.A(n), .B(m), .C(k), .Y(men_men_n379_));
  NA2        u0351(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n380_));
  NO3        u0352(.A(men_men_n380_), .B(men_men_n150_), .C(men_men_n207_), .Y(men_men_n381_));
  OR2        u0353(.A(m), .B(k), .Y(men_men_n382_));
  NO2        u0354(.A(men_men_n172_), .B(men_men_n382_), .Y(men_men_n383_));
  NA4        u0355(.A(n), .B(f), .C(c), .D(men_men_n114_), .Y(men_men_n384_));
  NOi21      u0356(.An(men_men_n383_), .B(men_men_n384_), .Y(men_men_n385_));
  NOi32      u0357(.An(d), .Bn(a), .C(c), .Y(men_men_n386_));
  NA2        u0358(.A(men_men_n386_), .B(men_men_n180_), .Y(men_men_n387_));
  NAi21      u0359(.An(i), .B(g), .Y(men_men_n388_));
  NAi31      u0360(.An(k), .B(m), .C(j), .Y(men_men_n389_));
  NO2        u0361(.A(men_men_n385_), .B(men_men_n381_), .Y(men_men_n390_));
  NO2        u0362(.A(men_men_n384_), .B(men_men_n292_), .Y(men_men_n391_));
  NOi32      u0363(.An(f), .Bn(d), .C(c), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n390_), .B(men_men_n377_), .Y(men_men_n393_));
  NO2        u0365(.A(men_men_n57_), .B(men_men_n114_), .Y(men_men_n394_));
  NA2        u0366(.A(men_men_n245_), .B(men_men_n394_), .Y(men_men_n395_));
  INV        u0367(.A(e), .Y(men_men_n396_));
  NA2        u0368(.A(men_men_n44_), .B(e), .Y(men_men_n397_));
  OAI220     u0369(.A0(men_men_n397_), .A1(men_men_n197_), .B0(men_men_n201_), .B1(men_men_n396_), .Y(men_men_n398_));
  AN2        u0370(.A(g), .B(e), .Y(men_men_n399_));
  NA3        u0371(.A(men_men_n399_), .B(men_men_n200_), .C(i), .Y(men_men_n400_));
  INV        u0372(.A(men_men_n400_), .Y(men_men_n401_));
  NO2        u0373(.A(men_men_n100_), .B(men_men_n396_), .Y(men_men_n402_));
  NO3        u0374(.A(men_men_n402_), .B(men_men_n401_), .C(men_men_n398_), .Y(men_men_n403_));
  NOi32      u0375(.An(h), .Bn(e), .C(g), .Y(men_men_n404_));
  NA3        u0376(.A(men_men_n404_), .B(men_men_n285_), .C(m), .Y(men_men_n405_));
  NOi21      u0377(.An(g), .B(h), .Y(men_men_n406_));
  AN3        u0378(.A(m), .B(l), .C(i), .Y(men_men_n407_));
  NA3        u0379(.A(men_men_n407_), .B(men_men_n406_), .C(e), .Y(men_men_n408_));
  AN3        u0380(.A(h), .B(g), .C(e), .Y(men_men_n409_));
  NA2        u0381(.A(men_men_n409_), .B(men_men_n97_), .Y(men_men_n410_));
  AN3        u0382(.A(men_men_n410_), .B(men_men_n408_), .C(men_men_n405_), .Y(men_men_n411_));
  AOI210     u0383(.A0(men_men_n411_), .A1(men_men_n403_), .B0(men_men_n395_), .Y(men_men_n412_));
  NA3        u0384(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n413_));
  NO2        u0385(.A(men_men_n413_), .B(men_men_n395_), .Y(men_men_n414_));
  NA3        u0386(.A(men_men_n386_), .B(men_men_n180_), .C(men_men_n83_), .Y(men_men_n415_));
  NAi31      u0387(.An(b), .B(c), .C(a), .Y(men_men_n416_));
  NO2        u0388(.A(men_men_n416_), .B(n), .Y(men_men_n417_));
  NO3        u0389(.A(men_men_n414_), .B(men_men_n412_), .C(men_men_n393_), .Y(men_men_n418_));
  NA2        u0390(.A(i), .B(g), .Y(men_men_n419_));
  NO3        u0391(.A(men_men_n271_), .B(men_men_n419_), .C(c), .Y(men_men_n420_));
  NOi21      u0392(.An(a), .B(n), .Y(men_men_n421_));
  NOi21      u0393(.An(d), .B(c), .Y(men_men_n422_));
  NA2        u0394(.A(men_men_n422_), .B(men_men_n421_), .Y(men_men_n423_));
  NA3        u0395(.A(i), .B(g), .C(f), .Y(men_men_n424_));
  OR2        u0396(.A(men_men_n424_), .B(men_men_n69_), .Y(men_men_n425_));
  NA3        u0397(.A(men_men_n407_), .B(men_men_n406_), .C(men_men_n180_), .Y(men_men_n426_));
  AOI210     u0398(.A0(men_men_n426_), .A1(men_men_n425_), .B0(men_men_n423_), .Y(men_men_n427_));
  AOI210     u0399(.A0(men_men_n420_), .A1(men_men_n284_), .B0(men_men_n427_), .Y(men_men_n428_));
  OR2        u0400(.A(n), .B(m), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n429_), .B(men_men_n151_), .Y(men_men_n430_));
  NO2        u0402(.A(men_men_n181_), .B(men_men_n146_), .Y(men_men_n431_));
  OAI210     u0403(.A0(men_men_n430_), .A1(men_men_n174_), .B0(men_men_n431_), .Y(men_men_n432_));
  INV        u0404(.A(men_men_n363_), .Y(men_men_n433_));
  NA3        u0405(.A(men_men_n433_), .B(men_men_n352_), .C(d), .Y(men_men_n434_));
  NO2        u0406(.A(men_men_n416_), .B(men_men_n47_), .Y(men_men_n435_));
  NO3        u0407(.A(men_men_n64_), .B(men_men_n110_), .C(e), .Y(men_men_n436_));
  NAi21      u0408(.An(k), .B(j), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n248_), .B(men_men_n437_), .Y(men_men_n438_));
  NA3        u0410(.A(men_men_n438_), .B(men_men_n436_), .C(men_men_n435_), .Y(men_men_n439_));
  NAi21      u0411(.An(e), .B(d), .Y(men_men_n440_));
  INV        u0412(.A(men_men_n440_), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n249_), .B(men_men_n207_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n442_), .B(men_men_n441_), .C(men_men_n220_), .Y(men_men_n443_));
  NA4        u0415(.A(men_men_n443_), .B(men_men_n439_), .C(men_men_n434_), .D(men_men_n432_), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n327_), .B(men_men_n207_), .Y(men_men_n445_));
  NA2        u0417(.A(men_men_n445_), .B(men_men_n441_), .Y(men_men_n446_));
  NOi31      u0418(.An(n), .B(m), .C(k), .Y(men_men_n447_));
  AOI220     u0419(.A0(men_men_n447_), .A1(men_men_n378_), .B0(men_men_n215_), .B1(men_men_n48_), .Y(men_men_n448_));
  NAi31      u0420(.An(g), .B(f), .C(c), .Y(men_men_n449_));
  OR3        u0421(.A(men_men_n449_), .B(men_men_n448_), .C(e), .Y(men_men_n450_));
  NA2        u0422(.A(men_men_n450_), .B(men_men_n446_), .Y(men_men_n451_));
  NOi41      u0423(.An(men_men_n428_), .B(men_men_n451_), .C(men_men_n444_), .D(men_men_n263_), .Y(men_men_n452_));
  NOi32      u0424(.An(c), .Bn(a), .C(b), .Y(men_men_n453_));
  NA2        u0425(.A(men_men_n453_), .B(men_men_n111_), .Y(men_men_n454_));
  INV        u0426(.A(men_men_n270_), .Y(men_men_n455_));
  AN2        u0427(.A(e), .B(d), .Y(men_men_n456_));
  NA2        u0428(.A(men_men_n456_), .B(men_men_n455_), .Y(men_men_n457_));
  INV        u0429(.A(men_men_n146_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n129_), .B(men_men_n41_), .Y(men_men_n459_));
  NO2        u0431(.A(men_men_n64_), .B(e), .Y(men_men_n460_));
  NOi31      u0432(.An(j), .B(k), .C(i), .Y(men_men_n461_));
  NOi21      u0433(.An(men_men_n163_), .B(men_men_n461_), .Y(men_men_n462_));
  NA3        u0434(.A(men_men_n312_), .B(men_men_n462_), .C(men_men_n117_), .Y(men_men_n463_));
  AOI220     u0435(.A0(men_men_n463_), .A1(men_men_n460_), .B0(men_men_n459_), .B1(men_men_n458_), .Y(men_men_n464_));
  AOI210     u0436(.A0(men_men_n464_), .A1(men_men_n457_), .B0(men_men_n454_), .Y(men_men_n465_));
  NOi21      u0437(.An(a), .B(b), .Y(men_men_n466_));
  NA3        u0438(.A(e), .B(d), .C(c), .Y(men_men_n467_));
  NAi21      u0439(.An(men_men_n467_), .B(men_men_n466_), .Y(men_men_n468_));
  NO2        u0440(.A(men_men_n415_), .B(men_men_n201_), .Y(men_men_n469_));
  NOi21      u0441(.An(men_men_n468_), .B(men_men_n469_), .Y(men_men_n470_));
  AOI210     u0442(.A0(men_men_n266_), .A1(men_men_n201_), .B0(men_men_n470_), .Y(men_men_n471_));
  NO4        u0443(.A(men_men_n184_), .B(men_men_n103_), .C(men_men_n54_), .D(b), .Y(men_men_n472_));
  OR2        u0444(.A(k), .B(j), .Y(men_men_n473_));
  NA2        u0445(.A(l), .B(k), .Y(men_men_n474_));
  NA3        u0446(.A(men_men_n272_), .B(men_men_n126_), .C(men_men_n124_), .Y(men_men_n475_));
  NA2        u0447(.A(men_men_n386_), .B(men_men_n111_), .Y(men_men_n476_));
  NO4        u0448(.A(men_men_n476_), .B(men_men_n94_), .C(men_men_n110_), .D(e), .Y(men_men_n477_));
  NO3        u0449(.A(men_men_n415_), .B(men_men_n91_), .C(men_men_n129_), .Y(men_men_n478_));
  NO4        u0450(.A(men_men_n478_), .B(men_men_n477_), .C(men_men_n475_), .D(men_men_n313_), .Y(men_men_n479_));
  INV        u0451(.A(men_men_n479_), .Y(men_men_n480_));
  NO4        u0452(.A(men_men_n480_), .B(men_men_n472_), .C(men_men_n471_), .D(men_men_n465_), .Y(men_men_n481_));
  NA2        u0453(.A(men_men_n68_), .B(men_men_n65_), .Y(men_men_n482_));
  NOi21      u0454(.An(d), .B(e), .Y(men_men_n483_));
  NAi31      u0455(.An(j), .B(l), .C(i), .Y(men_men_n484_));
  OAI210     u0456(.A0(men_men_n484_), .A1(men_men_n130_), .B0(men_men_n103_), .Y(men_men_n485_));
  NA2        u0457(.A(men_men_n482_), .B(men_men_n237_), .Y(men_men_n486_));
  OAI210     u0458(.A0(men_men_n125_), .A1(men_men_n123_), .B0(n), .Y(men_men_n487_));
  NO2        u0459(.A(men_men_n487_), .B(men_men_n129_), .Y(men_men_n488_));
  OR2        u0460(.A(men_men_n293_), .B(men_men_n239_), .Y(men_men_n489_));
  OA210      u0461(.A0(men_men_n489_), .A1(men_men_n488_), .B0(men_men_n189_), .Y(men_men_n490_));
  XO2        u0462(.A(i), .B(h), .Y(men_men_n491_));
  NA3        u0463(.A(men_men_n491_), .B(men_men_n159_), .C(n), .Y(men_men_n492_));
  NAi41      u0464(.An(men_men_n293_), .B(men_men_n492_), .C(men_men_n448_), .D(men_men_n375_), .Y(men_men_n493_));
  NOi32      u0465(.An(men_men_n493_), .Bn(men_men_n460_), .C(men_men_n1484_), .Y(men_men_n494_));
  NAi31      u0466(.An(c), .B(f), .C(d), .Y(men_men_n495_));
  AOI210     u0467(.A0(men_men_n273_), .A1(men_men_n192_), .B0(men_men_n495_), .Y(men_men_n496_));
  NOi21      u0468(.An(men_men_n81_), .B(men_men_n496_), .Y(men_men_n497_));
  NA3        u0469(.A(men_men_n371_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n498_));
  NA2        u0470(.A(men_men_n221_), .B(men_men_n106_), .Y(men_men_n499_));
  AOI210     u0471(.A0(men_men_n499_), .A1(men_men_n179_), .B0(men_men_n495_), .Y(men_men_n500_));
  NO2        u0472(.A(men_men_n35_), .B(men_men_n468_), .Y(men_men_n501_));
  NOi31      u0473(.An(men_men_n498_), .B(men_men_n501_), .C(men_men_n500_), .Y(men_men_n502_));
  AO220      u0474(.A0(men_men_n281_), .A1(men_men_n260_), .B0(men_men_n164_), .B1(men_men_n65_), .Y(men_men_n503_));
  NA3        u0475(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n504_));
  INV        u0476(.A(men_men_n289_), .Y(men_men_n505_));
  NAi41      u0477(.An(men_men_n503_), .B(men_men_n505_), .C(men_men_n502_), .D(men_men_n497_), .Y(men_men_n506_));
  NO4        u0478(.A(men_men_n506_), .B(men_men_n494_), .C(men_men_n490_), .D(men_men_n486_), .Y(men_men_n507_));
  NA4        u0479(.A(men_men_n507_), .B(men_men_n481_), .C(men_men_n452_), .D(men_men_n418_), .Y(men11));
  NO2        u0480(.A(men_men_n71_), .B(f), .Y(men_men_n509_));
  NA2        u0481(.A(j), .B(g), .Y(men_men_n510_));
  NAi31      u0482(.An(i), .B(m), .C(l), .Y(men_men_n511_));
  NA3        u0483(.A(m), .B(k), .C(j), .Y(men_men_n512_));
  OAI220     u0484(.A0(men_men_n512_), .A1(men_men_n129_), .B0(men_men_n511_), .B1(men_men_n510_), .Y(men_men_n513_));
  NA2        u0485(.A(men_men_n513_), .B(men_men_n509_), .Y(men_men_n514_));
  NOi32      u0486(.An(e), .Bn(b), .C(f), .Y(men_men_n515_));
  NA2        u0487(.A(men_men_n256_), .B(men_men_n111_), .Y(men_men_n516_));
  NA2        u0488(.A(men_men_n44_), .B(j), .Y(men_men_n517_));
  NO2        u0489(.A(men_men_n517_), .B(men_men_n295_), .Y(men_men_n518_));
  NAi31      u0490(.An(d), .B(e), .C(a), .Y(men_men_n519_));
  NO2        u0491(.A(men_men_n519_), .B(n), .Y(men_men_n520_));
  AOI220     u0492(.A0(men_men_n520_), .A1(men_men_n101_), .B0(men_men_n518_), .B1(men_men_n515_), .Y(men_men_n521_));
  NAi41      u0493(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n522_));
  AN2        u0494(.A(men_men_n522_), .B(men_men_n362_), .Y(men_men_n523_));
  AOI210     u0495(.A0(men_men_n523_), .A1(men_men_n387_), .B0(men_men_n268_), .Y(men_men_n524_));
  NA2        u0496(.A(j), .B(i), .Y(men_men_n525_));
  NAi31      u0497(.An(n), .B(m), .C(k), .Y(men_men_n526_));
  NO3        u0498(.A(men_men_n526_), .B(men_men_n525_), .C(men_men_n110_), .Y(men_men_n527_));
  NO4        u0499(.A(n), .B(d), .C(men_men_n114_), .D(a), .Y(men_men_n528_));
  OR2        u0500(.A(n), .B(c), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n148_), .Y(men_men_n530_));
  NO2        u0502(.A(men_men_n530_), .B(men_men_n528_), .Y(men_men_n531_));
  NOi32      u0503(.An(g), .Bn(f), .C(i), .Y(men_men_n532_));
  AOI220     u0504(.A0(men_men_n532_), .A1(men_men_n99_), .B0(men_men_n513_), .B1(f), .Y(men_men_n533_));
  NO2        u0505(.A(men_men_n270_), .B(men_men_n47_), .Y(men_men_n534_));
  NO2        u0506(.A(men_men_n533_), .B(men_men_n531_), .Y(men_men_n535_));
  AOI210     u0507(.A0(men_men_n527_), .A1(men_men_n524_), .B0(men_men_n535_), .Y(men_men_n536_));
  NA2        u0508(.A(men_men_n139_), .B(men_men_n34_), .Y(men_men_n537_));
  OAI220     u0509(.A0(men_men_n537_), .A1(m), .B0(men_men_n517_), .B1(men_men_n227_), .Y(men_men_n538_));
  NOi41      u0510(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n539_));
  AN2        u0511(.A(men_men_n331_), .B(men_men_n311_), .Y(men_men_n540_));
  INV        u0512(.A(men_men_n540_), .Y(men_men_n541_));
  OA210      u0513(.A0(men_men_n541_), .A1(men_men_n539_), .B0(men_men_n538_), .Y(men_men_n542_));
  OAI220     u0514(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n511_), .B1(men_men_n510_), .Y(men_men_n543_));
  NAi31      u0515(.An(d), .B(c), .C(a), .Y(men_men_n544_));
  NO2        u0516(.A(men_men_n544_), .B(n), .Y(men_men_n545_));
  NA3        u0517(.A(men_men_n545_), .B(men_men_n543_), .C(e), .Y(men_men_n546_));
  NO3        u0518(.A(men_men_n60_), .B(men_men_n47_), .C(men_men_n208_), .Y(men_men_n547_));
  NO2        u0519(.A(men_men_n224_), .B(men_men_n108_), .Y(men_men_n548_));
  NA2        u0520(.A(men_men_n547_), .B(men_men_n548_), .Y(men_men_n549_));
  NA2        u0521(.A(men_men_n549_), .B(men_men_n546_), .Y(men_men_n550_));
  NO2        u0522(.A(men_men_n271_), .B(n), .Y(men_men_n551_));
  NO2        u0523(.A(men_men_n417_), .B(men_men_n551_), .Y(men_men_n552_));
  NA2        u0524(.A(men_men_n543_), .B(f), .Y(men_men_n553_));
  NAi32      u0525(.An(d), .Bn(a), .C(b), .Y(men_men_n554_));
  NO2        u0526(.A(men_men_n554_), .B(men_men_n47_), .Y(men_men_n555_));
  NA2        u0527(.A(h), .B(f), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n556_), .B(men_men_n94_), .Y(men_men_n557_));
  NO3        u0529(.A(men_men_n175_), .B(men_men_n172_), .C(g), .Y(men_men_n558_));
  AOI220     u0530(.A0(men_men_n558_), .A1(men_men_n56_), .B0(men_men_n557_), .B1(men_men_n555_), .Y(men_men_n559_));
  OAI210     u0531(.A0(men_men_n553_), .A1(men_men_n552_), .B0(men_men_n559_), .Y(men_men_n560_));
  AN3        u0532(.A(j), .B(h), .C(g), .Y(men_men_n561_));
  NO2        u0533(.A(men_men_n145_), .B(c), .Y(men_men_n562_));
  NA3        u0534(.A(men_men_n562_), .B(men_men_n561_), .C(men_men_n447_), .Y(men_men_n563_));
  NA3        u0535(.A(f), .B(d), .C(b), .Y(men_men_n564_));
  NO4        u0536(.A(men_men_n564_), .B(men_men_n175_), .C(men_men_n172_), .D(g), .Y(men_men_n565_));
  NAi21      u0537(.An(men_men_n565_), .B(men_men_n563_), .Y(men_men_n566_));
  NO4        u0538(.A(men_men_n566_), .B(men_men_n560_), .C(men_men_n550_), .D(men_men_n542_), .Y(men_men_n567_));
  AN4        u0539(.A(men_men_n567_), .B(men_men_n536_), .C(men_men_n521_), .D(men_men_n514_), .Y(men_men_n568_));
  INV        u0540(.A(k), .Y(men_men_n569_));
  NA3        u0541(.A(l), .B(men_men_n569_), .C(i), .Y(men_men_n570_));
  INV        u0542(.A(men_men_n570_), .Y(men_men_n571_));
  NA4        u0543(.A(men_men_n386_), .B(men_men_n406_), .C(men_men_n180_), .D(men_men_n111_), .Y(men_men_n572_));
  NAi32      u0544(.An(h), .Bn(f), .C(g), .Y(men_men_n573_));
  NAi41      u0545(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n574_));
  OAI210     u0546(.A0(men_men_n519_), .A1(n), .B0(men_men_n574_), .Y(men_men_n575_));
  NA2        u0547(.A(men_men_n575_), .B(m), .Y(men_men_n576_));
  NAi31      u0548(.An(h), .B(g), .C(f), .Y(men_men_n577_));
  OR3        u0549(.A(men_men_n577_), .B(men_men_n271_), .C(men_men_n47_), .Y(men_men_n578_));
  NA4        u0550(.A(men_men_n406_), .B(men_men_n119_), .C(men_men_n111_), .D(e), .Y(men_men_n579_));
  AN2        u0551(.A(men_men_n579_), .B(men_men_n578_), .Y(men_men_n580_));
  OA210      u0552(.A0(men_men_n576_), .A1(men_men_n573_), .B0(men_men_n580_), .Y(men_men_n581_));
  NO3        u0553(.A(men_men_n573_), .B(men_men_n71_), .C(men_men_n73_), .Y(men_men_n582_));
  NO4        u0554(.A(men_men_n577_), .B(men_men_n529_), .C(men_men_n148_), .D(men_men_n73_), .Y(men_men_n583_));
  OR2        u0555(.A(men_men_n583_), .B(men_men_n582_), .Y(men_men_n584_));
  NAi31      u0556(.An(men_men_n584_), .B(men_men_n581_), .C(men_men_n572_), .Y(men_men_n585_));
  NAi31      u0557(.An(f), .B(h), .C(g), .Y(men_men_n586_));
  NO4        u0558(.A(men_men_n303_), .B(men_men_n586_), .C(men_men_n71_), .D(men_men_n73_), .Y(men_men_n587_));
  NOi32      u0559(.An(b), .Bn(a), .C(c), .Y(men_men_n588_));
  NOi41      u0560(.An(men_men_n588_), .B(men_men_n345_), .C(men_men_n67_), .D(men_men_n115_), .Y(men_men_n589_));
  OR2        u0561(.A(men_men_n589_), .B(men_men_n587_), .Y(men_men_n590_));
  NOi32      u0562(.An(d), .Bn(a), .C(e), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n111_), .Y(men_men_n592_));
  NO2        u0564(.A(n), .B(c), .Y(men_men_n593_));
  NA3        u0565(.A(men_men_n593_), .B(men_men_n29_), .C(m), .Y(men_men_n594_));
  NAi32      u0566(.An(n), .Bn(f), .C(m), .Y(men_men_n595_));
  NA3        u0567(.A(men_men_n595_), .B(men_men_n594_), .C(men_men_n592_), .Y(men_men_n596_));
  NOi32      u0568(.An(e), .Bn(a), .C(d), .Y(men_men_n597_));
  AOI210     u0569(.A0(men_men_n29_), .A1(d), .B0(men_men_n597_), .Y(men_men_n598_));
  AOI210     u0570(.A0(men_men_n598_), .A1(men_men_n207_), .B0(men_men_n537_), .Y(men_men_n599_));
  AOI210     u0571(.A0(men_men_n599_), .A1(men_men_n596_), .B0(men_men_n590_), .Y(men_men_n600_));
  OAI210     u0572(.A0(men_men_n244_), .A1(men_men_n86_), .B0(men_men_n600_), .Y(men_men_n601_));
  AOI210     u0573(.A0(men_men_n585_), .A1(men_men_n571_), .B0(men_men_n601_), .Y(men_men_n602_));
  NO3        u0574(.A(men_men_n310_), .B(men_men_n59_), .C(n), .Y(men_men_n603_));
  NA3        u0575(.A(men_men_n495_), .B(men_men_n170_), .C(men_men_n169_), .Y(men_men_n604_));
  NA2        u0576(.A(men_men_n449_), .B(men_men_n224_), .Y(men_men_n605_));
  OR2        u0577(.A(men_men_n605_), .B(men_men_n604_), .Y(men_men_n606_));
  NA2        u0578(.A(men_men_n74_), .B(men_men_n111_), .Y(men_men_n607_));
  NO2        u0579(.A(men_men_n607_), .B(men_men_n43_), .Y(men_men_n608_));
  AOI220     u0580(.A0(men_men_n608_), .A1(men_men_n524_), .B0(men_men_n606_), .B1(men_men_n603_), .Y(men_men_n609_));
  NO2        u0581(.A(men_men_n609_), .B(men_men_n86_), .Y(men_men_n610_));
  NA3        u0582(.A(men_men_n539_), .B(men_men_n333_), .C(men_men_n44_), .Y(men_men_n611_));
  NOi32      u0583(.An(e), .Bn(c), .C(f), .Y(men_men_n612_));
  NOi21      u0584(.An(f), .B(g), .Y(men_men_n613_));
  NO2        u0585(.A(men_men_n613_), .B(men_men_n205_), .Y(men_men_n614_));
  AOI220     u0586(.A0(men_men_n614_), .A1(men_men_n383_), .B0(men_men_n612_), .B1(men_men_n174_), .Y(men_men_n615_));
  NA3        u0587(.A(men_men_n615_), .B(men_men_n611_), .C(men_men_n177_), .Y(men_men_n616_));
  AOI210     u0588(.A0(men_men_n523_), .A1(men_men_n387_), .B0(men_men_n294_), .Y(men_men_n617_));
  NA2        u0589(.A(men_men_n617_), .B(men_men_n261_), .Y(men_men_n618_));
  NOi21      u0590(.An(j), .B(l), .Y(men_men_n619_));
  NAi21      u0591(.An(k), .B(h), .Y(men_men_n620_));
  NO2        u0592(.A(men_men_n620_), .B(men_men_n259_), .Y(men_men_n621_));
  NA2        u0593(.A(men_men_n621_), .B(men_men_n619_), .Y(men_men_n622_));
  OR2        u0594(.A(men_men_n622_), .B(men_men_n576_), .Y(men_men_n623_));
  NOi31      u0595(.An(m), .B(n), .C(k), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n619_), .B(men_men_n624_), .Y(men_men_n625_));
  NO2        u0597(.A(men_men_n271_), .B(men_men_n47_), .Y(men_men_n626_));
  NO2        u0598(.A(men_men_n303_), .B(men_men_n586_), .Y(men_men_n627_));
  NO2        u0599(.A(men_men_n519_), .B(men_men_n47_), .Y(men_men_n628_));
  AOI220     u0600(.A0(men_men_n628_), .A1(men_men_n627_), .B0(men_men_n626_), .B1(men_men_n557_), .Y(men_men_n629_));
  NA3        u0601(.A(men_men_n629_), .B(men_men_n623_), .C(men_men_n618_), .Y(men_men_n630_));
  NA2        u0602(.A(men_men_n106_), .B(men_men_n36_), .Y(men_men_n631_));
  NO2        u0603(.A(k), .B(men_men_n208_), .Y(men_men_n632_));
  NO2        u0604(.A(men_men_n515_), .B(men_men_n352_), .Y(men_men_n633_));
  NO2        u0605(.A(men_men_n633_), .B(n), .Y(men_men_n634_));
  NAi31      u0606(.An(men_men_n631_), .B(men_men_n634_), .C(men_men_n632_), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n491_), .B(men_men_n159_), .Y(men_men_n636_));
  NO3        u0608(.A(men_men_n384_), .B(men_men_n636_), .C(men_men_n86_), .Y(men_men_n637_));
  INV        u0609(.A(men_men_n637_), .Y(men_men_n638_));
  AN3        u0610(.A(f), .B(d), .C(b), .Y(men_men_n639_));
  OAI210     u0611(.A0(men_men_n639_), .A1(men_men_n128_), .B0(n), .Y(men_men_n640_));
  NA3        u0612(.A(men_men_n491_), .B(men_men_n159_), .C(men_men_n208_), .Y(men_men_n641_));
  AOI210     u0613(.A0(men_men_n640_), .A1(men_men_n226_), .B0(men_men_n641_), .Y(men_men_n642_));
  NAi31      u0614(.An(m), .B(n), .C(k), .Y(men_men_n643_));
  INV        u0615(.A(men_men_n246_), .Y(men_men_n644_));
  OAI210     u0616(.A0(men_men_n644_), .A1(men_men_n642_), .B0(j), .Y(men_men_n645_));
  NA3        u0617(.A(men_men_n645_), .B(men_men_n638_), .C(men_men_n635_), .Y(men_men_n646_));
  NO4        u0618(.A(men_men_n646_), .B(men_men_n630_), .C(men_men_n616_), .D(men_men_n610_), .Y(men_men_n647_));
  NAi31      u0619(.An(g), .B(h), .C(f), .Y(men_men_n648_));
  OA210      u0620(.A0(men_men_n519_), .A1(n), .B0(men_men_n574_), .Y(men_men_n649_));
  NO3        u0621(.A(g), .B(men_men_n207_), .C(men_men_n54_), .Y(men_men_n650_));
  NAi21      u0622(.An(h), .B(j), .Y(men_men_n651_));
  NO2        u0623(.A(men_men_n499_), .B(men_men_n86_), .Y(men_men_n652_));
  OAI210     u0624(.A0(men_men_n652_), .A1(men_men_n383_), .B0(men_men_n650_), .Y(men_men_n653_));
  OR2        u0625(.A(men_men_n71_), .B(men_men_n73_), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n588_), .B(men_men_n335_), .Y(men_men_n655_));
  OA220      u0627(.A0(men_men_n625_), .A1(men_men_n655_), .B0(men_men_n622_), .B1(men_men_n654_), .Y(men_men_n656_));
  NA3        u0628(.A(men_men_n509_), .B(men_men_n99_), .C(men_men_n98_), .Y(men_men_n657_));
  AN2        u0629(.A(h), .B(f), .Y(men_men_n658_));
  NA2        u0630(.A(men_men_n658_), .B(men_men_n37_), .Y(men_men_n659_));
  NA2        u0631(.A(men_men_n99_), .B(men_men_n44_), .Y(men_men_n660_));
  OAI220     u0632(.A0(men_men_n660_), .A1(men_men_n324_), .B0(men_men_n659_), .B1(men_men_n454_), .Y(men_men_n661_));
  AOI210     u0633(.A0(men_men_n554_), .A1(men_men_n416_), .B0(men_men_n47_), .Y(men_men_n662_));
  OAI220     u0634(.A0(men_men_n577_), .A1(men_men_n570_), .B0(men_men_n317_), .B1(men_men_n510_), .Y(men_men_n663_));
  AOI210     u0635(.A0(men_men_n663_), .A1(men_men_n662_), .B0(men_men_n661_), .Y(men_men_n664_));
  NA4        u0636(.A(men_men_n664_), .B(men_men_n657_), .C(men_men_n656_), .D(men_men_n653_), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n248_), .B(f), .Y(men_men_n666_));
  NO2        u0638(.A(men_men_n613_), .B(men_men_n59_), .Y(men_men_n667_));
  NO3        u0639(.A(men_men_n667_), .B(men_men_n666_), .C(men_men_n34_), .Y(men_men_n668_));
  NA2        u0640(.A(men_men_n320_), .B(men_men_n139_), .Y(men_men_n669_));
  NA2        u0641(.A(men_men_n130_), .B(men_men_n47_), .Y(men_men_n670_));
  NA2        u0642(.A(men_men_n670_), .B(men_men_n515_), .Y(men_men_n671_));
  OA220      u0643(.A0(men_men_n671_), .A1(men_men_n537_), .B0(men_men_n350_), .B1(men_men_n109_), .Y(men_men_n672_));
  OAI210     u0644(.A0(men_men_n669_), .A1(men_men_n668_), .B0(men_men_n672_), .Y(men_men_n673_));
  NO3        u0645(.A(men_men_n392_), .B(men_men_n189_), .C(men_men_n188_), .Y(men_men_n674_));
  NA2        u0646(.A(men_men_n674_), .B(men_men_n224_), .Y(men_men_n675_));
  NA3        u0647(.A(men_men_n675_), .B(men_men_n250_), .C(j), .Y(men_men_n676_));
  NO3        u0648(.A(men_men_n449_), .B(men_men_n172_), .C(i), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n453_), .B(men_men_n83_), .Y(men_men_n678_));
  NO4        u0650(.A(men_men_n512_), .B(men_men_n678_), .C(men_men_n129_), .D(men_men_n207_), .Y(men_men_n679_));
  INV        u0651(.A(men_men_n679_), .Y(men_men_n680_));
  NA4        u0652(.A(men_men_n680_), .B(men_men_n676_), .C(men_men_n498_), .D(men_men_n390_), .Y(men_men_n681_));
  NO3        u0653(.A(men_men_n681_), .B(men_men_n673_), .C(men_men_n665_), .Y(men_men_n682_));
  NA4        u0654(.A(men_men_n682_), .B(men_men_n647_), .C(men_men_n602_), .D(men_men_n568_), .Y(men08));
  NO2        u0655(.A(k), .B(h), .Y(men_men_n684_));
  AO210      u0656(.A0(men_men_n248_), .A1(men_men_n437_), .B0(men_men_n684_), .Y(men_men_n685_));
  NO2        u0657(.A(men_men_n685_), .B(men_men_n292_), .Y(men_men_n686_));
  NA2        u0658(.A(men_men_n612_), .B(men_men_n83_), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n687_), .B(men_men_n449_), .Y(men_men_n688_));
  AOI210     u0660(.A0(men_men_n688_), .A1(men_men_n686_), .B0(men_men_n478_), .Y(men_men_n689_));
  NA2        u0661(.A(men_men_n83_), .B(men_men_n108_), .Y(men_men_n690_));
  NO2        u0662(.A(men_men_n690_), .B(men_men_n55_), .Y(men_men_n691_));
  NA2        u0663(.A(men_men_n564_), .B(men_men_n226_), .Y(men_men_n692_));
  AOI210     u0664(.A0(men_men_n564_), .A1(men_men_n155_), .B0(men_men_n83_), .Y(men_men_n693_));
  NA4        u0665(.A(men_men_n210_), .B(men_men_n139_), .C(men_men_n43_), .D(h), .Y(men_men_n694_));
  AN2        u0666(.A(l), .B(k), .Y(men_men_n695_));
  NA2        u0667(.A(men_men_n689_), .B(men_men_n341_), .Y(men_men_n696_));
  AN2        u0668(.A(men_men_n520_), .B(men_men_n95_), .Y(men_men_n697_));
  NO4        u0669(.A(men_men_n172_), .B(men_men_n382_), .C(men_men_n110_), .D(g), .Y(men_men_n698_));
  NA2        u0670(.A(men_men_n698_), .B(men_men_n692_), .Y(men_men_n699_));
  NO2        u0671(.A(men_men_n38_), .B(men_men_n207_), .Y(men_men_n700_));
  AOI220     u0672(.A0(men_men_n614_), .A1(men_men_n338_), .B0(men_men_n700_), .B1(men_men_n551_), .Y(men_men_n701_));
  NAi31      u0673(.An(men_men_n697_), .B(men_men_n701_), .C(men_men_n699_), .Y(men_men_n702_));
  NO2        u0674(.A(men_men_n523_), .B(men_men_n35_), .Y(men_men_n703_));
  INV        u0675(.A(men_men_n703_), .Y(men_men_n704_));
  NO3        u0676(.A(men_men_n310_), .B(men_men_n129_), .C(men_men_n41_), .Y(men_men_n705_));
  BUFFER     u0677(.A(men_men_n705_), .Y(men_men_n706_));
  INV        u0678(.A(men_men_n685_), .Y(men_men_n707_));
  AOI220     u0679(.A0(men_men_n707_), .A1(men_men_n391_), .B0(men_men_n706_), .B1(men_men_n76_), .Y(men_men_n708_));
  OAI210     u0680(.A0(men_men_n704_), .A1(men_men_n86_), .B0(men_men_n708_), .Y(men_men_n709_));
  NA3        u0681(.A(men_men_n675_), .B(men_men_n326_), .C(men_men_n374_), .Y(men_men_n710_));
  NA2        u0682(.A(men_men_n695_), .B(men_men_n215_), .Y(men_men_n711_));
  NO2        u0683(.A(men_men_n711_), .B(men_men_n319_), .Y(men_men_n712_));
  AOI210     u0684(.A0(men_men_n712_), .A1(men_men_n666_), .B0(men_men_n477_), .Y(men_men_n713_));
  NA3        u0685(.A(m), .B(l), .C(k), .Y(men_men_n714_));
  NO2        u0686(.A(men_men_n522_), .B(men_men_n268_), .Y(men_men_n715_));
  NOi21      u0687(.An(men_men_n715_), .B(men_men_n516_), .Y(men_men_n716_));
  NA4        u0688(.A(men_men_n111_), .B(l), .C(k), .D(men_men_n86_), .Y(men_men_n717_));
  NA3        u0689(.A(men_men_n119_), .B(men_men_n399_), .C(i), .Y(men_men_n718_));
  NO2        u0690(.A(men_men_n718_), .B(men_men_n717_), .Y(men_men_n719_));
  NO2        u0691(.A(men_men_n719_), .B(men_men_n716_), .Y(men_men_n720_));
  NA3        u0692(.A(men_men_n720_), .B(men_men_n713_), .C(men_men_n710_), .Y(men_men_n721_));
  NO4        u0693(.A(men_men_n721_), .B(men_men_n709_), .C(men_men_n702_), .D(men_men_n696_), .Y(men_men_n722_));
  NA2        u0694(.A(men_men_n614_), .B(men_men_n383_), .Y(men_men_n723_));
  NOi31      u0695(.An(g), .B(h), .C(f), .Y(men_men_n724_));
  NA2        u0696(.A(men_men_n628_), .B(men_men_n724_), .Y(men_men_n725_));
  AO210      u0697(.A0(men_men_n725_), .A1(men_men_n578_), .B0(men_men_n525_), .Y(men_men_n726_));
  NO3        u0698(.A(men_men_n387_), .B(men_men_n510_), .C(h), .Y(men_men_n727_));
  NA2        u0699(.A(men_men_n727_), .B(men_men_n111_), .Y(men_men_n728_));
  NA4        u0700(.A(men_men_n728_), .B(men_men_n726_), .C(men_men_n723_), .D(men_men_n247_), .Y(men_men_n729_));
  NA2        u0701(.A(men_men_n695_), .B(men_men_n73_), .Y(men_men_n730_));
  NO4        u0702(.A(men_men_n674_), .B(men_men_n172_), .C(n), .D(i), .Y(men_men_n731_));
  NOi21      u0703(.An(h), .B(j), .Y(men_men_n732_));
  NA2        u0704(.A(men_men_n732_), .B(f), .Y(men_men_n733_));
  NO2        u0705(.A(men_men_n733_), .B(men_men_n241_), .Y(men_men_n734_));
  NO3        u0706(.A(men_men_n734_), .B(men_men_n731_), .C(men_men_n677_), .Y(men_men_n735_));
  OAI220     u0707(.A0(men_men_n735_), .A1(men_men_n730_), .B0(men_men_n580_), .B1(men_men_n60_), .Y(men_men_n736_));
  AOI210     u0708(.A0(men_men_n729_), .A1(l), .B0(men_men_n736_), .Y(men_men_n737_));
  NO2        u0709(.A(j), .B(i), .Y(men_men_n738_));
  NA3        u0710(.A(men_men_n738_), .B(men_men_n80_), .C(l), .Y(men_men_n739_));
  NA2        u0711(.A(men_men_n738_), .B(men_men_n33_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n409_), .B(men_men_n119_), .Y(men_men_n741_));
  OA220      u0713(.A0(men_men_n741_), .A1(men_men_n740_), .B0(men_men_n739_), .B1(men_men_n576_), .Y(men_men_n742_));
  NO3        u0714(.A(men_men_n150_), .B(men_men_n47_), .C(men_men_n108_), .Y(men_men_n743_));
  NO3        u0715(.A(men_men_n529_), .B(men_men_n148_), .C(men_men_n73_), .Y(men_men_n744_));
  NO3        u0716(.A(men_men_n474_), .B(men_men_n424_), .C(j), .Y(men_men_n745_));
  OAI210     u0717(.A0(men_men_n744_), .A1(men_men_n743_), .B0(men_men_n745_), .Y(men_men_n746_));
  OAI210     u0718(.A0(men_men_n725_), .A1(men_men_n60_), .B0(men_men_n746_), .Y(men_men_n747_));
  NA2        u0719(.A(k), .B(j), .Y(men_men_n748_));
  NO3        u0720(.A(men_men_n292_), .B(men_men_n748_), .C(men_men_n40_), .Y(men_men_n749_));
  AOI210     u0721(.A0(men_men_n515_), .A1(n), .B0(men_men_n539_), .Y(men_men_n750_));
  NA2        u0722(.A(men_men_n750_), .B(men_men_n540_), .Y(men_men_n751_));
  AN3        u0723(.A(men_men_n751_), .B(men_men_n749_), .C(men_men_n98_), .Y(men_men_n752_));
  NAi31      u0724(.An(men_men_n598_), .B(men_men_n92_), .C(men_men_n83_), .Y(men_men_n753_));
  INV        u0725(.A(men_men_n753_), .Y(men_men_n754_));
  NO2        u0726(.A(men_men_n292_), .B(men_men_n134_), .Y(men_men_n755_));
  AOI220     u0727(.A0(men_men_n755_), .A1(men_men_n614_), .B0(men_men_n705_), .B1(men_men_n693_), .Y(men_men_n756_));
  NO2        u0728(.A(men_men_n714_), .B(men_men_n90_), .Y(men_men_n757_));
  NA2        u0729(.A(men_men_n757_), .B(men_men_n575_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n758_), .B(men_men_n756_), .Y(men_men_n759_));
  OR4        u0731(.A(men_men_n759_), .B(men_men_n754_), .C(men_men_n752_), .D(men_men_n747_), .Y(men_men_n760_));
  NA2        u0732(.A(men_men_n750_), .B(men_men_n540_), .Y(men_men_n761_));
  NA4        u0733(.A(men_men_n761_), .B(men_men_n210_), .C(men_men_n437_), .D(men_men_n34_), .Y(men_men_n762_));
  NO4        u0734(.A(men_men_n474_), .B(men_men_n419_), .C(j), .D(f), .Y(men_men_n763_));
  OAI220     u0735(.A0(men_men_n694_), .A1(men_men_n687_), .B0(men_men_n324_), .B1(men_men_n38_), .Y(men_men_n764_));
  AOI210     u0736(.A0(men_men_n763_), .A1(men_men_n254_), .B0(men_men_n764_), .Y(men_men_n765_));
  NA3        u0737(.A(men_men_n532_), .B(men_men_n285_), .C(h), .Y(men_men_n766_));
  NOi21      u0738(.An(men_men_n662_), .B(men_men_n766_), .Y(men_men_n767_));
  NO2        u0739(.A(men_men_n91_), .B(men_men_n45_), .Y(men_men_n768_));
  OAI220     u0740(.A0(men_men_n766_), .A1(men_men_n594_), .B0(men_men_n739_), .B1(men_men_n654_), .Y(men_men_n769_));
  AOI210     u0741(.A0(men_men_n768_), .A1(men_men_n634_), .B0(men_men_n769_), .Y(men_men_n770_));
  NAi41      u0742(.An(men_men_n767_), .B(men_men_n770_), .C(men_men_n765_), .D(men_men_n762_), .Y(men_men_n771_));
  BUFFER     u0743(.A(men_men_n95_), .Y(men_men_n772_));
  AOI220     u0744(.A0(men_men_n772_), .A1(men_men_n232_), .B0(men_men_n745_), .B1(men_men_n626_), .Y(men_men_n773_));
  NO2        u0745(.A(men_men_n649_), .B(men_men_n73_), .Y(men_men_n774_));
  AOI210     u0746(.A0(men_men_n763_), .A1(men_men_n774_), .B0(men_men_n328_), .Y(men_men_n775_));
  OAI210     u0747(.A0(men_men_n714_), .A1(men_men_n648_), .B0(men_men_n504_), .Y(men_men_n776_));
  NA3        u0748(.A(men_men_n245_), .B(men_men_n57_), .C(b), .Y(men_men_n777_));
  AOI220     u0749(.A0(men_men_n593_), .A1(men_men_n29_), .B0(men_men_n453_), .B1(men_men_n83_), .Y(men_men_n778_));
  NA2        u0750(.A(men_men_n778_), .B(men_men_n777_), .Y(men_men_n779_));
  NO2        u0751(.A(men_men_n766_), .B(men_men_n476_), .Y(men_men_n780_));
  AOI210     u0752(.A0(men_men_n779_), .A1(men_men_n776_), .B0(men_men_n780_), .Y(men_men_n781_));
  NA3        u0753(.A(men_men_n781_), .B(men_men_n775_), .C(men_men_n773_), .Y(men_men_n782_));
  NOi41      u0754(.An(men_men_n742_), .B(men_men_n782_), .C(men_men_n771_), .D(men_men_n760_), .Y(men_men_n783_));
  OR3        u0755(.A(men_men_n694_), .B(men_men_n226_), .C(g), .Y(men_men_n784_));
  NO3        u0756(.A(men_men_n334_), .B(men_men_n294_), .C(men_men_n110_), .Y(men_men_n785_));
  NA2        u0757(.A(men_men_n785_), .B(men_men_n751_), .Y(men_men_n786_));
  NA2        u0758(.A(men_men_n44_), .B(men_men_n54_), .Y(men_men_n787_));
  NO3        u0759(.A(men_men_n787_), .B(men_men_n740_), .C(men_men_n271_), .Y(men_men_n788_));
  NO3        u0760(.A(men_men_n510_), .B(men_men_n93_), .C(h), .Y(men_men_n789_));
  AOI210     u0761(.A0(men_men_n789_), .A1(men_men_n691_), .B0(men_men_n788_), .Y(men_men_n790_));
  NA3        u0762(.A(men_men_n790_), .B(men_men_n786_), .C(men_men_n784_), .Y(men_men_n791_));
  OR2        u0763(.A(men_men_n648_), .B(men_men_n91_), .Y(men_men_n792_));
  NOi31      u0764(.An(b), .B(d), .C(a), .Y(men_men_n793_));
  NO2        u0765(.A(men_men_n793_), .B(men_men_n591_), .Y(men_men_n794_));
  NO2        u0766(.A(men_men_n794_), .B(n), .Y(men_men_n795_));
  NOi21      u0767(.An(men_men_n778_), .B(men_men_n795_), .Y(men_men_n796_));
  OAI220     u0768(.A0(men_men_n796_), .A1(men_men_n792_), .B0(men_men_n766_), .B1(men_men_n592_), .Y(men_men_n797_));
  NO3        u0769(.A(men_men_n613_), .B(men_men_n319_), .C(men_men_n115_), .Y(men_men_n798_));
  NOi21      u0770(.An(men_men_n798_), .B(men_men_n160_), .Y(men_men_n799_));
  INV        u0771(.A(men_men_n799_), .Y(men_men_n800_));
  OAI210     u0772(.A0(men_men_n694_), .A1(men_men_n384_), .B0(men_men_n800_), .Y(men_men_n801_));
  NO2        u0773(.A(men_men_n674_), .B(n), .Y(men_men_n802_));
  AOI220     u0774(.A0(men_men_n755_), .A1(men_men_n650_), .B0(men_men_n802_), .B1(men_men_n686_), .Y(men_men_n803_));
  NO2        u0775(.A(men_men_n314_), .B(men_men_n231_), .Y(men_men_n804_));
  OAI210     u0776(.A0(men_men_n95_), .A1(men_men_n92_), .B0(men_men_n804_), .Y(men_men_n805_));
  NA2        u0777(.A(men_men_n119_), .B(men_men_n83_), .Y(men_men_n806_));
  AOI210     u0778(.A0(men_men_n413_), .A1(men_men_n405_), .B0(men_men_n806_), .Y(men_men_n807_));
  NAi21      u0779(.An(men_men_n807_), .B(men_men_n805_), .Y(men_men_n808_));
  NA2        u0780(.A(men_men_n712_), .B(men_men_n34_), .Y(men_men_n809_));
  NAi21      u0781(.An(men_men_n717_), .B(men_men_n420_), .Y(men_men_n810_));
  NO2        u0782(.A(men_men_n268_), .B(i), .Y(men_men_n811_));
  NA2        u0783(.A(men_men_n698_), .B(men_men_n340_), .Y(men_men_n812_));
  OAI210     u0784(.A0(men_men_n583_), .A1(men_men_n582_), .B0(men_men_n353_), .Y(men_men_n813_));
  AN3        u0785(.A(men_men_n813_), .B(men_men_n812_), .C(men_men_n810_), .Y(men_men_n814_));
  NAi41      u0786(.An(men_men_n808_), .B(men_men_n814_), .C(men_men_n809_), .D(men_men_n803_), .Y(men_men_n815_));
  NO4        u0787(.A(men_men_n815_), .B(men_men_n801_), .C(men_men_n797_), .D(men_men_n791_), .Y(men_men_n816_));
  NA4        u0788(.A(men_men_n816_), .B(men_men_n783_), .C(men_men_n737_), .D(men_men_n722_), .Y(men09));
  INV        u0789(.A(men_men_n120_), .Y(men_men_n818_));
  NA2        u0790(.A(f), .B(e), .Y(men_men_n819_));
  NO2        u0791(.A(men_men_n219_), .B(men_men_n110_), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n820_), .B(g), .Y(men_men_n821_));
  NA4        u0793(.A(men_men_n303_), .B(men_men_n462_), .C(men_men_n257_), .D(men_men_n117_), .Y(men_men_n822_));
  AOI210     u0794(.A0(men_men_n822_), .A1(g), .B0(men_men_n459_), .Y(men_men_n823_));
  AOI210     u0795(.A0(men_men_n823_), .A1(men_men_n821_), .B0(men_men_n819_), .Y(men_men_n824_));
  NA2        u0796(.A(men_men_n824_), .B(men_men_n818_), .Y(men_men_n825_));
  NA3        u0797(.A(m), .B(l), .C(i), .Y(men_men_n826_));
  OAI220     u0798(.A0(men_men_n577_), .A1(men_men_n826_), .B0(men_men_n345_), .B1(men_men_n511_), .Y(men_men_n827_));
  NAi21      u0799(.An(men_men_n827_), .B(men_men_n425_), .Y(men_men_n828_));
  NA3        u0800(.A(men_men_n792_), .B(men_men_n553_), .C(men_men_n504_), .Y(men_men_n829_));
  OA210      u0801(.A0(men_men_n829_), .A1(men_men_n828_), .B0(men_men_n795_), .Y(men_men_n830_));
  INV        u0802(.A(men_men_n331_), .Y(men_men_n831_));
  NOi31      u0803(.An(k), .B(m), .C(l), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n333_), .B(men_men_n832_), .Y(men_men_n833_));
  NO2        u0805(.A(men_men_n833_), .B(men_men_n586_), .Y(men_men_n834_));
  NA2        u0806(.A(men_men_n777_), .B(men_men_n324_), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n335_), .B(men_men_n337_), .Y(men_men_n836_));
  OAI210     u0808(.A0(men_men_n201_), .A1(men_men_n207_), .B0(men_men_n836_), .Y(men_men_n837_));
  AOI220     u0809(.A0(men_men_n837_), .A1(men_men_n835_), .B0(men_men_n834_), .B1(men_men_n831_), .Y(men_men_n838_));
  NA2        u0810(.A(men_men_n167_), .B(men_men_n112_), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n839_), .B(men_men_n685_), .Y(men_men_n840_));
  NA3        u0812(.A(men_men_n840_), .B(men_men_n186_), .C(men_men_n31_), .Y(men_men_n841_));
  NA4        u0813(.A(men_men_n841_), .B(men_men_n838_), .C(men_men_n615_), .D(men_men_n81_), .Y(men_men_n842_));
  NO2        u0814(.A(men_men_n573_), .B(men_men_n484_), .Y(men_men_n843_));
  NOi21      u0815(.An(f), .B(d), .Y(men_men_n844_));
  NA2        u0816(.A(men_men_n844_), .B(m), .Y(men_men_n845_));
  NO2        u0817(.A(men_men_n845_), .B(men_men_n50_), .Y(men_men_n846_));
  NOi32      u0818(.An(g), .Bn(f), .C(d), .Y(men_men_n847_));
  NA4        u0819(.A(men_men_n847_), .B(men_men_n593_), .C(men_men_n29_), .D(m), .Y(men_men_n848_));
  NA2        u0820(.A(men_men_n846_), .B(men_men_n530_), .Y(men_men_n849_));
  NA3        u0821(.A(men_men_n303_), .B(men_men_n257_), .C(men_men_n117_), .Y(men_men_n850_));
  AN2        u0822(.A(f), .B(d), .Y(men_men_n851_));
  NA3        u0823(.A(men_men_n466_), .B(men_men_n851_), .C(men_men_n83_), .Y(men_men_n852_));
  NO3        u0824(.A(men_men_n852_), .B(men_men_n73_), .C(men_men_n208_), .Y(men_men_n853_));
  NO2        u0825(.A(men_men_n278_), .B(men_men_n54_), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n850_), .B(men_men_n853_), .Y(men_men_n855_));
  NAi31      u0827(.An(men_men_n475_), .B(men_men_n855_), .C(men_men_n849_), .Y(men_men_n856_));
  NO4        u0828(.A(men_men_n613_), .B(men_men_n130_), .C(men_men_n319_), .D(men_men_n151_), .Y(men_men_n857_));
  NO2        u0829(.A(men_men_n643_), .B(men_men_n319_), .Y(men_men_n858_));
  AN2        u0830(.A(men_men_n858_), .B(men_men_n666_), .Y(men_men_n859_));
  NO3        u0831(.A(men_men_n859_), .B(men_men_n857_), .C(men_men_n228_), .Y(men_men_n860_));
  NA2        u0832(.A(men_men_n591_), .B(men_men_n83_), .Y(men_men_n861_));
  NO2        u0833(.A(men_men_n836_), .B(men_men_n861_), .Y(men_men_n862_));
  NA3        u0834(.A(men_men_n159_), .B(men_men_n106_), .C(men_men_n105_), .Y(men_men_n863_));
  NO2        u0835(.A(men_men_n331_), .B(men_men_n863_), .Y(men_men_n864_));
  NO2        u0836(.A(men_men_n864_), .B(men_men_n862_), .Y(men_men_n865_));
  NA2        u0837(.A(c), .B(men_men_n114_), .Y(men_men_n866_));
  NO2        u0838(.A(men_men_n866_), .B(men_men_n396_), .Y(men_men_n867_));
  NA3        u0839(.A(men_men_n867_), .B(men_men_n493_), .C(f), .Y(men_men_n868_));
  OR2        u0840(.A(men_men_n648_), .B(men_men_n526_), .Y(men_men_n869_));
  INV        u0841(.A(men_men_n869_), .Y(men_men_n870_));
  NA2        u0842(.A(men_men_n794_), .B(men_men_n109_), .Y(men_men_n871_));
  NA2        u0843(.A(men_men_n871_), .B(men_men_n870_), .Y(men_men_n872_));
  NA4        u0844(.A(men_men_n872_), .B(men_men_n868_), .C(men_men_n865_), .D(men_men_n860_), .Y(men_men_n873_));
  NO4        u0845(.A(men_men_n873_), .B(men_men_n856_), .C(men_men_n842_), .D(men_men_n830_), .Y(men_men_n874_));
  OR2        u0846(.A(men_men_n852_), .B(men_men_n73_), .Y(men_men_n875_));
  NA2        u0847(.A(men_men_n820_), .B(g), .Y(men_men_n876_));
  AOI210     u0848(.A0(men_men_n876_), .A1(men_men_n286_), .B0(men_men_n875_), .Y(men_men_n877_));
  NO2        u0849(.A(men_men_n134_), .B(men_men_n130_), .Y(men_men_n878_));
  NO2        u0850(.A(men_men_n224_), .B(men_men_n218_), .Y(men_men_n879_));
  AOI220     u0851(.A0(men_men_n879_), .A1(men_men_n221_), .B0(men_men_n299_), .B1(men_men_n878_), .Y(men_men_n880_));
  NA2        u0852(.A(e), .B(d), .Y(men_men_n881_));
  OAI220     u0853(.A0(men_men_n881_), .A1(c), .B0(men_men_n314_), .B1(d), .Y(men_men_n882_));
  NA3        u0854(.A(men_men_n882_), .B(men_men_n442_), .C(men_men_n491_), .Y(men_men_n883_));
  AOI210     u0855(.A0(men_men_n499_), .A1(men_men_n179_), .B0(men_men_n224_), .Y(men_men_n884_));
  AOI210     u0856(.A0(men_men_n614_), .A1(men_men_n338_), .B0(men_men_n884_), .Y(men_men_n885_));
  NA2        u0857(.A(men_men_n278_), .B(men_men_n163_), .Y(men_men_n886_));
  NA3        u0858(.A(men_men_n166_), .B(men_men_n84_), .C(men_men_n34_), .Y(men_men_n887_));
  NA3        u0859(.A(men_men_n887_), .B(men_men_n885_), .C(men_men_n883_), .Y(men_men_n888_));
  NO3        u0860(.A(men_men_n888_), .B(men_men_n1483_), .C(men_men_n877_), .Y(men_men_n889_));
  OAI220     u0861(.A0(men_men_n613_), .A1(men_men_n59_), .B0(men_men_n294_), .B1(j), .Y(men_men_n890_));
  AOI220     u0862(.A0(men_men_n890_), .A1(men_men_n858_), .B0(men_men_n603_), .B1(men_men_n612_), .Y(men_men_n891_));
  INV        u0863(.A(men_men_n891_), .Y(men_men_n892_));
  OAI210     u0864(.A0(men_men_n820_), .A1(men_men_n886_), .B0(men_men_n847_), .Y(men_men_n893_));
  NO2        u0865(.A(men_men_n893_), .B(men_men_n594_), .Y(men_men_n894_));
  AOI210     u0866(.A0(men_men_n116_), .A1(men_men_n115_), .B0(men_men_n256_), .Y(men_men_n895_));
  NO2        u0867(.A(men_men_n895_), .B(men_men_n848_), .Y(men_men_n896_));
  AO210      u0868(.A0(men_men_n835_), .A1(men_men_n827_), .B0(men_men_n896_), .Y(men_men_n897_));
  NO3        u0869(.A(men_men_n897_), .B(men_men_n894_), .C(men_men_n892_), .Y(men_men_n898_));
  AO220      u0870(.A0(men_men_n442_), .A1(men_men_n732_), .B0(men_men_n174_), .B1(f), .Y(men_men_n899_));
  OAI210     u0871(.A0(men_men_n899_), .A1(men_men_n445_), .B0(men_men_n882_), .Y(men_men_n900_));
  NA2        u0872(.A(men_men_n829_), .B(men_men_n691_), .Y(men_men_n901_));
  AN3        u0873(.A(men_men_n901_), .B(men_men_n900_), .C(men_men_n898_), .Y(men_men_n902_));
  NA4        u0874(.A(men_men_n902_), .B(men_men_n889_), .C(men_men_n874_), .D(men_men_n825_), .Y(men12));
  NO2        u0875(.A(men_men_n440_), .B(c), .Y(men_men_n904_));
  NO4        u0876(.A(men_men_n429_), .B(men_men_n248_), .C(men_men_n569_), .D(men_men_n208_), .Y(men_men_n905_));
  NA2        u0877(.A(men_men_n905_), .B(men_men_n904_), .Y(men_men_n906_));
  NO2        u0878(.A(men_men_n440_), .B(men_men_n114_), .Y(men_men_n907_));
  NO2        u0879(.A(men_men_n648_), .B(men_men_n368_), .Y(men_men_n908_));
  NA2        u0880(.A(men_men_n908_), .B(men_men_n528_), .Y(men_men_n909_));
  NA3        u0881(.A(men_men_n909_), .B(men_men_n906_), .C(men_men_n428_), .Y(men_men_n910_));
  AOI210     u0882(.A0(men_men_n227_), .A1(men_men_n330_), .B0(men_men_n198_), .Y(men_men_n911_));
  OR2        u0883(.A(men_men_n911_), .B(men_men_n905_), .Y(men_men_n912_));
  AOI210     u0884(.A0(men_men_n327_), .A1(men_men_n380_), .B0(men_men_n208_), .Y(men_men_n913_));
  OAI210     u0885(.A0(men_men_n913_), .A1(men_men_n912_), .B0(men_men_n392_), .Y(men_men_n914_));
  NO2        u0886(.A(men_men_n631_), .B(men_men_n259_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n577_), .B(men_men_n826_), .Y(men_men_n916_));
  AOI220     u0888(.A0(men_men_n916_), .A1(men_men_n551_), .B0(men_men_n804_), .B1(men_men_n915_), .Y(men_men_n917_));
  NO2        u0889(.A(men_men_n150_), .B(men_men_n231_), .Y(men_men_n918_));
  NA2        u0890(.A(men_men_n917_), .B(men_men_n914_), .Y(men_men_n919_));
  OR2        u0891(.A(men_men_n315_), .B(men_men_n907_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n920_), .B(men_men_n346_), .Y(men_men_n921_));
  NO3        u0893(.A(men_men_n130_), .B(men_men_n151_), .C(men_men_n208_), .Y(men_men_n922_));
  NA2        u0894(.A(men_men_n922_), .B(men_men_n515_), .Y(men_men_n923_));
  NA2        u0895(.A(men_men_n923_), .B(men_men_n921_), .Y(men_men_n924_));
  NO3        u0896(.A(men_men_n924_), .B(men_men_n919_), .C(men_men_n910_), .Y(men_men_n925_));
  NO2        u0897(.A(men_men_n360_), .B(men_men_n359_), .Y(men_men_n926_));
  NA2        u0898(.A(men_men_n574_), .B(men_men_n71_), .Y(men_men_n927_));
  NOi21      u0899(.An(men_men_n34_), .B(men_men_n643_), .Y(men_men_n928_));
  NA2        u0900(.A(men_men_n927_), .B(men_men_n926_), .Y(men_men_n929_));
  OAI210     u0901(.A0(men_men_n246_), .A1(men_men_n43_), .B0(men_men_n929_), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n420_), .B(men_men_n261_), .Y(men_men_n931_));
  NO3        u0903(.A(men_men_n806_), .B(men_men_n88_), .C(men_men_n396_), .Y(men_men_n932_));
  NAi21      u0904(.An(men_men_n932_), .B(men_men_n931_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n47_), .B(men_men_n43_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n624_), .B(men_men_n353_), .Y(men_men_n935_));
  OAI210     u0907(.A0(men_men_n718_), .A1(men_men_n935_), .B0(men_men_n357_), .Y(men_men_n936_));
  NO3        u0908(.A(men_men_n936_), .B(men_men_n933_), .C(men_men_n930_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n161_), .B(i), .Y(men_men_n938_));
  NA2        u0910(.A(men_men_n44_), .B(i), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n939_), .B(men_men_n197_), .Y(men_men_n940_));
  AOI210     u0912(.A0(men_men_n407_), .A1(men_men_n37_), .B0(men_men_n940_), .Y(men_men_n941_));
  NO2        u0913(.A(men_men_n941_), .B(men_men_n324_), .Y(men_men_n942_));
  NO2        u0914(.A(men_men_n648_), .B(men_men_n484_), .Y(men_men_n943_));
  NA3        u0915(.A(men_men_n335_), .B(men_men_n619_), .C(i), .Y(men_men_n944_));
  OAI210     u0916(.A0(men_men_n424_), .A1(men_men_n303_), .B0(men_men_n944_), .Y(men_men_n945_));
  OAI220     u0917(.A0(men_men_n945_), .A1(men_men_n943_), .B0(men_men_n662_), .B1(men_men_n744_), .Y(men_men_n946_));
  NA2        u0918(.A(men_men_n597_), .B(men_men_n111_), .Y(men_men_n947_));
  OR3        u0919(.A(men_men_n303_), .B(men_men_n419_), .C(f), .Y(men_men_n948_));
  NA3        u0920(.A(men_men_n619_), .B(men_men_n80_), .C(i), .Y(men_men_n949_));
  OA220      u0921(.A0(men_men_n949_), .A1(men_men_n947_), .B0(men_men_n948_), .B1(men_men_n576_), .Y(men_men_n950_));
  NA3        u0922(.A(men_men_n316_), .B(men_men_n116_), .C(g), .Y(men_men_n951_));
  AOI210     u0923(.A0(men_men_n659_), .A1(men_men_n951_), .B0(m), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n952_), .B(men_men_n315_), .Y(men_men_n953_));
  NA2        u0925(.A(men_men_n678_), .B(men_men_n861_), .Y(men_men_n954_));
  INV        u0926(.A(men_men_n425_), .Y(men_men_n955_));
  NA2        u0927(.A(men_men_n216_), .B(men_men_n77_), .Y(men_men_n956_));
  NA3        u0928(.A(men_men_n956_), .B(men_men_n949_), .C(men_men_n948_), .Y(men_men_n957_));
  AOI220     u0929(.A0(men_men_n957_), .A1(men_men_n254_), .B0(men_men_n955_), .B1(men_men_n954_), .Y(men_men_n958_));
  NA4        u0930(.A(men_men_n958_), .B(men_men_n953_), .C(men_men_n950_), .D(men_men_n946_), .Y(men_men_n959_));
  NO2        u0931(.A(men_men_n368_), .B(men_men_n90_), .Y(men_men_n960_));
  OAI210     u0932(.A0(men_men_n960_), .A1(men_men_n915_), .B0(men_men_n232_), .Y(men_men_n961_));
  NO2        u0933(.A(men_men_n448_), .B(men_men_n208_), .Y(men_men_n962_));
  AOI220     u0934(.A0(men_men_n962_), .A1(men_men_n373_), .B0(men_men_n920_), .B1(men_men_n212_), .Y(men_men_n963_));
  AOI220     u0935(.A0(men_men_n908_), .A1(men_men_n918_), .B0(men_men_n575_), .B1(men_men_n89_), .Y(men_men_n964_));
  NA3        u0936(.A(men_men_n964_), .B(men_men_n963_), .C(men_men_n961_), .Y(men_men_n965_));
  NA2        u0937(.A(men_men_n955_), .B(men_men_n528_), .Y(men_men_n966_));
  AOI210     u0938(.A0(men_men_n408_), .A1(men_men_n400_), .B0(men_men_n806_), .Y(men_men_n967_));
  OAI210     u0939(.A0(men_men_n360_), .A1(men_men_n359_), .B0(men_men_n107_), .Y(men_men_n968_));
  AOI210     u0940(.A0(men_men_n968_), .A1(men_men_n520_), .B0(men_men_n967_), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n952_), .B(men_men_n907_), .Y(men_men_n970_));
  NA3        u0942(.A(men_men_n970_), .B(men_men_n969_), .C(men_men_n966_), .Y(men_men_n971_));
  NO4        u0943(.A(men_men_n971_), .B(men_men_n965_), .C(men_men_n959_), .D(men_men_n942_), .Y(men_men_n972_));
  NAi31      u0944(.An(men_men_n140_), .B(men_men_n409_), .C(n), .Y(men_men_n973_));
  NO2        u0945(.A(men_men_n333_), .B(men_men_n832_), .Y(men_men_n974_));
  NO2        u0946(.A(men_men_n974_), .B(men_men_n973_), .Y(men_men_n975_));
  NO3        u0947(.A(men_men_n268_), .B(men_men_n140_), .C(men_men_n396_), .Y(men_men_n976_));
  AOI210     u0948(.A0(men_men_n976_), .A1(men_men_n485_), .B0(men_men_n975_), .Y(men_men_n977_));
  NA2        u0949(.A(men_men_n478_), .B(i), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n978_), .B(men_men_n977_), .Y(men_men_n979_));
  NA2        u0951(.A(men_men_n224_), .B(men_men_n170_), .Y(men_men_n980_));
  NO2        u0952(.A(men_men_n430_), .B(men_men_n174_), .Y(men_men_n981_));
  NOi31      u0953(.An(men_men_n980_), .B(men_men_n981_), .C(men_men_n208_), .Y(men_men_n982_));
  NA2        u0954(.A(men_men_n423_), .B(men_men_n861_), .Y(men_men_n983_));
  NO3        u0955(.A(men_men_n424_), .B(men_men_n303_), .C(men_men_n73_), .Y(men_men_n984_));
  AOI220     u0956(.A0(men_men_n984_), .A1(men_men_n983_), .B0(men_men_n472_), .B1(g), .Y(men_men_n985_));
  INV        u0957(.A(men_men_n985_), .Y(men_men_n986_));
  OAI220     u0958(.A0(men_men_n973_), .A1(men_men_n227_), .B0(men_men_n944_), .B1(men_men_n592_), .Y(men_men_n987_));
  NA2        u0959(.A(men_men_n911_), .B(men_men_n904_), .Y(men_men_n988_));
  NO3        u0960(.A(men_men_n529_), .B(men_men_n148_), .C(men_men_n207_), .Y(men_men_n989_));
  OAI210     u0961(.A0(men_men_n989_), .A1(men_men_n509_), .B0(men_men_n369_), .Y(men_men_n990_));
  OAI220     u0962(.A0(men_men_n908_), .A1(men_men_n916_), .B0(men_men_n530_), .B1(men_men_n417_), .Y(men_men_n991_));
  NA4        u0963(.A(men_men_n991_), .B(men_men_n990_), .C(men_men_n988_), .D(men_men_n611_), .Y(men_men_n992_));
  OAI210     u0964(.A0(men_men_n911_), .A1(men_men_n905_), .B0(men_men_n980_), .Y(men_men_n993_));
  AOI210     u0965(.A0(men_men_n371_), .A1(men_men_n369_), .B0(men_men_n323_), .Y(men_men_n994_));
  NA3        u0966(.A(men_men_n994_), .B(men_men_n993_), .C(men_men_n269_), .Y(men_men_n995_));
  OR3        u0967(.A(men_men_n995_), .B(men_men_n992_), .C(men_men_n987_), .Y(men_men_n996_));
  NO4        u0968(.A(men_men_n996_), .B(men_men_n986_), .C(men_men_n982_), .D(men_men_n979_), .Y(men_men_n997_));
  NA4        u0969(.A(men_men_n997_), .B(men_men_n972_), .C(men_men_n937_), .D(men_men_n925_), .Y(men13));
  NA3        u0970(.A(men_men_n245_), .B(b), .C(m), .Y(men_men_n999_));
  NA2        u0971(.A(men_men_n483_), .B(f), .Y(men_men_n1000_));
  NO4        u0972(.A(men_men_n1000_), .B(men_men_n999_), .C(j), .D(men_men_n570_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n261_), .B(b), .Y(men_men_n1002_));
  NO4        u0974(.A(men_men_n1002_), .B(men_men_n1000_), .C(men_men_n938_), .D(a), .Y(men_men_n1003_));
  NAi32      u0975(.An(d), .Bn(c), .C(e), .Y(men_men_n1004_));
  NA2        u0976(.A(men_men_n139_), .B(men_men_n43_), .Y(men_men_n1005_));
  NO4        u0977(.A(men_men_n1005_), .B(men_men_n1004_), .C(men_men_n577_), .D(men_men_n301_), .Y(men_men_n1006_));
  NA2        u0978(.A(men_men_n651_), .B(men_men_n218_), .Y(men_men_n1007_));
  NA2        u0979(.A(men_men_n399_), .B(men_men_n207_), .Y(men_men_n1008_));
  AN2        u0980(.A(d), .B(c), .Y(men_men_n1009_));
  NA2        u0981(.A(men_men_n1009_), .B(men_men_n114_), .Y(men_men_n1010_));
  NO4        u0982(.A(men_men_n1010_), .B(men_men_n1008_), .C(men_men_n175_), .D(men_men_n167_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n483_), .B(c), .Y(men_men_n1012_));
  NO4        u0984(.A(men_men_n1005_), .B(men_men_n573_), .C(men_men_n1012_), .D(men_men_n301_), .Y(men_men_n1013_));
  AO210      u0985(.A0(men_men_n1011_), .A1(men_men_n1007_), .B0(men_men_n1013_), .Y(men_men_n1014_));
  OR4        u0986(.A(men_men_n1014_), .B(men_men_n1006_), .C(men_men_n1003_), .D(men_men_n1001_), .Y(men_men_n1015_));
  NAi32      u0987(.An(f), .Bn(e), .C(c), .Y(men_men_n1016_));
  NO2        u0988(.A(men_men_n1016_), .B(men_men_n145_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n1017_), .B(g), .Y(men_men_n1018_));
  OR3        u0990(.A(men_men_n218_), .B(men_men_n175_), .C(men_men_n167_), .Y(men_men_n1019_));
  NO2        u0991(.A(men_men_n1019_), .B(men_men_n1018_), .Y(men_men_n1020_));
  NO2        u0992(.A(men_men_n1012_), .B(men_men_n301_), .Y(men_men_n1021_));
  NO2        u0993(.A(j), .B(men_men_n43_), .Y(men_men_n1022_));
  NA2        u0994(.A(men_men_n621_), .B(men_men_n1022_), .Y(men_men_n1023_));
  NOi21      u0995(.An(men_men_n1021_), .B(men_men_n1023_), .Y(men_men_n1024_));
  NO2        u0996(.A(men_men_n748_), .B(men_men_n110_), .Y(men_men_n1025_));
  NOi41      u0997(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1026_));
  NA2        u0998(.A(men_men_n1026_), .B(men_men_n1025_), .Y(men_men_n1027_));
  NO2        u0999(.A(men_men_n1027_), .B(men_men_n1018_), .Y(men_men_n1028_));
  OR3        u1000(.A(e), .B(d), .C(c), .Y(men_men_n1029_));
  NA3        u1001(.A(k), .B(j), .C(i), .Y(men_men_n1030_));
  NO3        u1002(.A(men_men_n1030_), .B(men_men_n301_), .C(men_men_n90_), .Y(men_men_n1031_));
  NOi21      u1003(.An(men_men_n1031_), .B(men_men_n1029_), .Y(men_men_n1032_));
  OR4        u1004(.A(men_men_n1032_), .B(men_men_n1028_), .C(men_men_n1024_), .D(men_men_n1020_), .Y(men_men_n1033_));
  NA3        u1005(.A(men_men_n456_), .B(men_men_n326_), .C(men_men_n54_), .Y(men_men_n1034_));
  NO2        u1006(.A(men_men_n1034_), .B(men_men_n1023_), .Y(men_men_n1035_));
  NO4        u1007(.A(men_men_n1034_), .B(men_men_n573_), .C(men_men_n437_), .D(men_men_n43_), .Y(men_men_n1036_));
  NO2        u1008(.A(f), .B(c), .Y(men_men_n1037_));
  NOi21      u1009(.An(men_men_n1037_), .B(men_men_n429_), .Y(men_men_n1038_));
  NA2        u1010(.A(men_men_n1038_), .B(men_men_n57_), .Y(men_men_n1039_));
  NO3        u1011(.A(i), .B(men_men_n238_), .C(l), .Y(men_men_n1040_));
  NOi31      u1012(.An(men_men_n1040_), .B(men_men_n1039_), .C(j), .Y(men_men_n1041_));
  OR3        u1013(.A(men_men_n1041_), .B(men_men_n1036_), .C(men_men_n1035_), .Y(men_men_n1042_));
  OR3        u1014(.A(men_men_n1042_), .B(men_men_n1033_), .C(men_men_n1015_), .Y(men02));
  OR3        u1015(.A(h), .B(g), .C(f), .Y(men_men_n1044_));
  OR3        u1016(.A(n), .B(m), .C(i), .Y(men_men_n1045_));
  NO4        u1017(.A(men_men_n1045_), .B(men_men_n1044_), .C(l), .D(men_men_n1029_), .Y(men_men_n1046_));
  NOi31      u1018(.An(e), .B(d), .C(c), .Y(men_men_n1047_));
  AOI210     u1019(.A0(men_men_n1031_), .A1(men_men_n1047_), .B0(men_men_n1006_), .Y(men_men_n1048_));
  AN3        u1020(.A(g), .B(f), .C(c), .Y(men_men_n1049_));
  NA3        u1021(.A(men_men_n1049_), .B(men_men_n456_), .C(h), .Y(men_men_n1050_));
  OR2        u1022(.A(men_men_n1030_), .B(men_men_n301_), .Y(men_men_n1051_));
  OR2        u1023(.A(men_men_n1051_), .B(men_men_n1050_), .Y(men_men_n1052_));
  NO3        u1024(.A(men_men_n1034_), .B(men_men_n1005_), .C(men_men_n573_), .Y(men_men_n1053_));
  NO2        u1025(.A(men_men_n1053_), .B(men_men_n1020_), .Y(men_men_n1054_));
  NA3        u1026(.A(l), .B(k), .C(j), .Y(men_men_n1055_));
  NA2        u1027(.A(i), .B(h), .Y(men_men_n1056_));
  NO3        u1028(.A(men_men_n1056_), .B(men_men_n1055_), .C(men_men_n130_), .Y(men_men_n1057_));
  NO3        u1029(.A(men_men_n141_), .B(men_men_n276_), .C(men_men_n208_), .Y(men_men_n1058_));
  AOI210     u1030(.A0(men_men_n1058_), .A1(men_men_n1057_), .B0(men_men_n1024_), .Y(men_men_n1059_));
  NA3        u1031(.A(c), .B(b), .C(a), .Y(men_men_n1060_));
  NO3        u1032(.A(men_men_n1060_), .B(men_men_n881_), .C(men_men_n207_), .Y(men_men_n1061_));
  NO3        u1033(.A(men_men_n1030_), .B(men_men_n47_), .C(men_men_n110_), .Y(men_men_n1062_));
  AOI210     u1034(.A0(men_men_n1062_), .A1(men_men_n1061_), .B0(men_men_n1035_), .Y(men_men_n1063_));
  AN4        u1035(.A(men_men_n1063_), .B(men_men_n1059_), .C(men_men_n1054_), .D(men_men_n1052_), .Y(men_men_n1064_));
  NO2        u1036(.A(men_men_n1010_), .B(men_men_n1008_), .Y(men_men_n1065_));
  NA2        u1037(.A(men_men_n1027_), .B(men_men_n1019_), .Y(men_men_n1066_));
  AOI210     u1038(.A0(men_men_n1066_), .A1(men_men_n1065_), .B0(men_men_n1001_), .Y(men_men_n1067_));
  NAi41      u1039(.An(men_men_n1046_), .B(men_men_n1067_), .C(men_men_n1064_), .D(men_men_n1048_), .Y(men03));
  NO2        u1040(.A(men_men_n511_), .B(men_men_n586_), .Y(men_men_n1069_));
  NA4        u1041(.A(men_men_n87_), .B(men_men_n86_), .C(g), .D(men_men_n207_), .Y(men_men_n1070_));
  INV        u1042(.A(men_men_n1070_), .Y(men_men_n1071_));
  NO3        u1043(.A(men_men_n1071_), .B(men_men_n1069_), .C(men_men_n968_), .Y(men_men_n1072_));
  NOi41      u1044(.An(men_men_n792_), .B(men_men_n837_), .C(men_men_n828_), .D(men_men_n700_), .Y(men_men_n1073_));
  OAI220     u1045(.A0(men_men_n1073_), .A1(men_men_n678_), .B0(men_men_n1072_), .B1(men_men_n574_), .Y(men_men_n1074_));
  NA4        u1046(.A(i), .B(men_men_n1047_), .C(men_men_n335_), .D(men_men_n326_), .Y(men_men_n1075_));
  OAI210     u1047(.A0(men_men_n806_), .A1(men_men_n410_), .B0(men_men_n1075_), .Y(men_men_n1076_));
  NOi31      u1048(.An(m), .B(n), .C(f), .Y(men_men_n1077_));
  NA2        u1049(.A(men_men_n1077_), .B(men_men_n49_), .Y(men_men_n1078_));
  AN2        u1050(.A(e), .B(c), .Y(men_men_n1079_));
  NA2        u1051(.A(men_men_n1079_), .B(a), .Y(men_men_n1080_));
  OAI220     u1052(.A0(men_men_n1080_), .A1(men_men_n1078_), .B0(men_men_n869_), .B1(men_men_n416_), .Y(men_men_n1081_));
  NA2        u1053(.A(men_men_n491_), .B(l), .Y(men_men_n1082_));
  NO3        u1054(.A(men_men_n1081_), .B(men_men_n1076_), .C(men_men_n967_), .Y(men_men_n1083_));
  NO2        u1055(.A(men_men_n276_), .B(a), .Y(men_men_n1084_));
  INV        u1056(.A(men_men_n1006_), .Y(men_men_n1085_));
  NO2        u1057(.A(men_men_n1056_), .B(men_men_n474_), .Y(men_men_n1086_));
  NO2        u1058(.A(men_men_n86_), .B(g), .Y(men_men_n1087_));
  AOI210     u1059(.A0(men_men_n1087_), .A1(men_men_n1086_), .B0(men_men_n1040_), .Y(men_men_n1088_));
  OR2        u1060(.A(men_men_n1088_), .B(men_men_n1039_), .Y(men_men_n1089_));
  NA3        u1061(.A(men_men_n1089_), .B(men_men_n1085_), .C(men_men_n1083_), .Y(men_men_n1090_));
  NO4        u1062(.A(men_men_n1090_), .B(men_men_n1074_), .C(men_men_n808_), .D(men_men_n550_), .Y(men_men_n1091_));
  NA2        u1063(.A(c), .B(b), .Y(men_men_n1092_));
  NO2        u1064(.A(men_men_n690_), .B(men_men_n1092_), .Y(men_men_n1093_));
  OAI210     u1065(.A0(men_men_n845_), .A1(men_men_n823_), .B0(men_men_n403_), .Y(men_men_n1094_));
  OAI210     u1066(.A0(men_men_n1094_), .A1(men_men_n846_), .B0(men_men_n1093_), .Y(men_men_n1095_));
  NAi21      u1067(.An(men_men_n411_), .B(men_men_n1093_), .Y(men_men_n1096_));
  OAI210     u1068(.A0(men_men_n534_), .A1(men_men_n39_), .B0(men_men_n1084_), .Y(men_men_n1097_));
  NA2        u1069(.A(men_men_n1097_), .B(men_men_n1096_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n257_), .B(men_men_n117_), .Y(men_men_n1099_));
  OAI210     u1071(.A0(men_men_n1099_), .A1(men_men_n280_), .B0(g), .Y(men_men_n1100_));
  NAi21      u1072(.An(f), .B(d), .Y(men_men_n1101_));
  NO2        u1073(.A(men_men_n1101_), .B(men_men_n1060_), .Y(men_men_n1102_));
  INV        u1074(.A(men_men_n1102_), .Y(men_men_n1103_));
  AOI210     u1075(.A0(men_men_n1100_), .A1(men_men_n286_), .B0(men_men_n1103_), .Y(men_men_n1104_));
  AOI210     u1076(.A0(men_men_n1104_), .A1(men_men_n111_), .B0(men_men_n1098_), .Y(men_men_n1105_));
  NO2        u1077(.A(men_men_n181_), .B(men_men_n231_), .Y(men_men_n1106_));
  NA2        u1078(.A(men_men_n1106_), .B(m), .Y(men_men_n1107_));
  NA3        u1079(.A(men_men_n895_), .B(men_men_n1082_), .C(men_men_n462_), .Y(men_men_n1108_));
  NA2        u1080(.A(men_men_n1108_), .B(men_men_n460_), .Y(men_men_n1109_));
  NO2        u1081(.A(men_men_n1109_), .B(men_men_n1107_), .Y(men_men_n1110_));
  NA2        u1082(.A(men_men_n545_), .B(men_men_n398_), .Y(men_men_n1111_));
  NA2        u1083(.A(men_men_n158_), .B(men_men_n33_), .Y(men_men_n1112_));
  AOI210     u1084(.A0(men_men_n935_), .A1(men_men_n1112_), .B0(men_men_n208_), .Y(men_men_n1113_));
  OAI210     u1085(.A0(men_men_n1113_), .A1(men_men_n433_), .B0(men_men_n1102_), .Y(men_men_n1114_));
  INV        u1086(.A(men_men_n932_), .Y(men_men_n1115_));
  NA3        u1087(.A(men_men_n1115_), .B(men_men_n1114_), .C(men_men_n1111_), .Y(men_men_n1116_));
  NO2        u1088(.A(men_men_n1116_), .B(men_men_n1110_), .Y(men_men_n1117_));
  NA4        u1089(.A(men_men_n1117_), .B(men_men_n1105_), .C(men_men_n1095_), .D(men_men_n1091_), .Y(men00));
  INV        u1090(.A(men_men_n1076_), .Y(men_men_n1119_));
  NO3        u1091(.A(men_men_n1053_), .B(men_men_n932_), .C(men_men_n697_), .Y(men_men_n1120_));
  NA3        u1092(.A(men_men_n1120_), .B(men_men_n1119_), .C(men_men_n969_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n493_), .B(f), .Y(men_men_n1122_));
  NO2        u1094(.A(men_men_n974_), .B(men_men_n40_), .Y(men_men_n1123_));
  NA3        u1095(.A(men_men_n1123_), .B(men_men_n253_), .C(n), .Y(men_men_n1124_));
  AOI210     u1096(.A0(men_men_n1124_), .A1(men_men_n1122_), .B0(men_men_n1010_), .Y(men_men_n1125_));
  NO3        u1097(.A(men_men_n1125_), .B(men_men_n1121_), .C(men_men_n1033_), .Y(men_men_n1126_));
  NA3        u1098(.A(men_men_n166_), .B(men_men_n44_), .C(men_men_n43_), .Y(men_men_n1127_));
  NA3        u1099(.A(d), .B(men_men_n54_), .C(b), .Y(men_men_n1128_));
  NOi31      u1100(.An(n), .B(m), .C(i), .Y(men_men_n1129_));
  NA3        u1101(.A(men_men_n1129_), .B(men_men_n639_), .C(men_men_n49_), .Y(men_men_n1130_));
  OAI210     u1102(.A0(men_men_n1128_), .A1(men_men_n1127_), .B0(men_men_n1130_), .Y(men_men_n1131_));
  INV        u1103(.A(men_men_n563_), .Y(men_men_n1132_));
  NO2        u1104(.A(men_men_n1132_), .B(men_men_n1131_), .Y(men_men_n1133_));
  OR2        u1105(.A(men_men_n375_), .B(men_men_n133_), .Y(men_men_n1134_));
  NO2        u1106(.A(h), .B(g), .Y(men_men_n1135_));
  OAI220     u1107(.A0(men_men_n511_), .A1(men_men_n586_), .B0(men_men_n91_), .B1(men_men_n90_), .Y(men_men_n1136_));
  AOI220     u1108(.A0(men_men_n1136_), .A1(men_men_n520_), .B0(men_men_n922_), .B1(men_men_n562_), .Y(men_men_n1137_));
  NA2        u1109(.A(men_men_n1137_), .B(men_men_n1134_), .Y(men_men_n1138_));
  NO2        u1110(.A(men_men_n1138_), .B(men_men_n263_), .Y(men_men_n1139_));
  INV        u1111(.A(men_men_n313_), .Y(men_men_n1140_));
  AOI210     u1112(.A0(men_men_n242_), .A1(men_men_n338_), .B0(men_men_n565_), .Y(men_men_n1141_));
  NA3        u1113(.A(men_men_n1141_), .B(men_men_n1140_), .C(men_men_n153_), .Y(men_men_n1142_));
  NO2        u1114(.A(men_men_n233_), .B(men_men_n180_), .Y(men_men_n1143_));
  NA2        u1115(.A(men_men_n1143_), .B(men_men_n417_), .Y(men_men_n1144_));
  NA3        u1116(.A(men_men_n178_), .B(men_men_n110_), .C(g), .Y(men_men_n1145_));
  NA3        u1117(.A(men_men_n456_), .B(men_men_n40_), .C(f), .Y(men_men_n1146_));
  NOi31      u1118(.An(men_men_n854_), .B(men_men_n1146_), .C(men_men_n1145_), .Y(men_men_n1147_));
  NAi31      u1119(.An(men_men_n182_), .B(men_men_n843_), .C(men_men_n456_), .Y(men_men_n1148_));
  NAi31      u1120(.An(men_men_n1147_), .B(men_men_n1148_), .C(men_men_n1144_), .Y(men_men_n1149_));
  NO2        u1121(.A(men_men_n270_), .B(men_men_n73_), .Y(men_men_n1150_));
  NO3        u1122(.A(men_men_n416_), .B(men_men_n819_), .C(n), .Y(men_men_n1151_));
  AOI210     u1123(.A0(men_men_n1151_), .A1(men_men_n1150_), .B0(men_men_n1046_), .Y(men_men_n1152_));
  NAi31      u1124(.An(men_men_n1013_), .B(men_men_n1152_), .C(men_men_n72_), .Y(men_men_n1153_));
  NO4        u1125(.A(men_men_n1153_), .B(men_men_n1149_), .C(men_men_n1142_), .D(men_men_n503_), .Y(men_men_n1154_));
  AN3        u1126(.A(men_men_n1154_), .B(men_men_n1139_), .C(men_men_n1133_), .Y(men_men_n1155_));
  NA2        u1127(.A(men_men_n520_), .B(men_men_n101_), .Y(men_men_n1156_));
  NA3        u1128(.A(men_men_n1077_), .B(men_men_n597_), .C(men_men_n455_), .Y(men_men_n1157_));
  NA4        u1129(.A(men_men_n1157_), .B(men_men_n546_), .C(men_men_n1156_), .D(men_men_n236_), .Y(men_men_n1158_));
  NA2        u1130(.A(men_men_n1071_), .B(men_men_n520_), .Y(men_men_n1159_));
  NA2        u1131(.A(men_men_n1159_), .B(men_men_n290_), .Y(men_men_n1160_));
  OAI210     u1132(.A0(men_men_n454_), .A1(men_men_n118_), .B0(men_men_n848_), .Y(men_men_n1161_));
  AOI220     u1133(.A0(men_men_n1161_), .A1(men_men_n1108_), .B0(men_men_n545_), .B1(men_men_n398_), .Y(men_men_n1162_));
  OR4        u1134(.A(men_men_n1010_), .B(men_men_n268_), .C(men_men_n217_), .D(e), .Y(men_men_n1163_));
  NA2        u1135(.A(n), .B(e), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n1164_), .B(men_men_n145_), .Y(men_men_n1165_));
  NA2        u1137(.A(men_men_n1163_), .B(men_men_n1162_), .Y(men_men_n1166_));
  AOI210     u1138(.A0(men_men_n1165_), .A1(men_men_n834_), .B0(men_men_n807_), .Y(men_men_n1167_));
  AOI220     u1139(.A0(men_men_n928_), .A1(men_men_n562_), .B0(men_men_n639_), .B1(men_men_n239_), .Y(men_men_n1168_));
  NO2        u1140(.A(men_men_n66_), .B(h), .Y(men_men_n1169_));
  NO3        u1141(.A(men_men_n1010_), .B(men_men_n1008_), .C(men_men_n711_), .Y(men_men_n1170_));
  INV        u1142(.A(men_men_n130_), .Y(men_men_n1171_));
  AN2        u1143(.A(men_men_n1171_), .B(men_men_n1058_), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n1172_), .A1(men_men_n1170_), .B0(men_men_n1169_), .Y(men_men_n1173_));
  NA4        u1145(.A(men_men_n1173_), .B(men_men_n1168_), .C(men_men_n1167_), .D(men_men_n849_), .Y(men_men_n1174_));
  NO4        u1146(.A(men_men_n1174_), .B(men_men_n1166_), .C(men_men_n1160_), .D(men_men_n1158_), .Y(men_men_n1175_));
  NA2        u1147(.A(men_men_n824_), .B(men_men_n743_), .Y(men_men_n1176_));
  NA4        u1148(.A(men_men_n1176_), .B(men_men_n1175_), .C(men_men_n1155_), .D(men_men_n1126_), .Y(men01));
  AN2        u1149(.A(men_men_n990_), .B(men_men_n988_), .Y(men_men_n1178_));
  NO4        u1150(.A(men_men_n788_), .B(men_men_n780_), .C(men_men_n469_), .D(men_men_n274_), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n579_), .B(men_men_n283_), .Y(men_men_n1180_));
  OAI210     u1152(.A0(men_men_n1180_), .A1(men_men_n385_), .B0(i), .Y(men_men_n1181_));
  NA3        u1153(.A(men_men_n1181_), .B(men_men_n1179_), .C(men_men_n1178_), .Y(men_men_n1182_));
  NA2        u1154(.A(men_men_n575_), .B(men_men_n89_), .Y(men_men_n1183_));
  NA3        u1155(.A(men_men_n1183_), .B(men_men_n891_), .C(men_men_n325_), .Y(men_men_n1184_));
  NA2        u1156(.A(men_men_n43_), .B(f), .Y(men_men_n1185_));
  NA2        u1157(.A(men_men_n695_), .B(men_men_n96_), .Y(men_men_n1186_));
  NO2        u1158(.A(men_men_n1186_), .B(men_men_n1185_), .Y(men_men_n1187_));
  NO2        u1159(.A(men_men_n766_), .B(men_men_n592_), .Y(men_men_n1188_));
  AOI210     u1160(.A0(men_men_n1187_), .A1(men_men_n626_), .B0(men_men_n1188_), .Y(men_men_n1189_));
  INV        u1161(.A(men_men_n116_), .Y(men_men_n1190_));
  OR2        u1162(.A(men_men_n1190_), .B(men_men_n572_), .Y(men_men_n1191_));
  NA3        u1163(.A(men_men_n1191_), .B(men_men_n1189_), .C(men_men_n880_), .Y(men_men_n1192_));
  NO3        u1164(.A(men_men_n767_), .B(men_men_n661_), .C(men_men_n496_), .Y(men_men_n1193_));
  NA4        u1165(.A(men_men_n695_), .B(men_men_n96_), .C(men_men_n43_), .D(men_men_n207_), .Y(men_men_n1194_));
  OA220      u1166(.A0(men_men_n1194_), .A1(men_men_n654_), .B0(men_men_n192_), .B1(men_men_n190_), .Y(men_men_n1195_));
  NA3        u1167(.A(men_men_n1195_), .B(men_men_n1193_), .C(men_men_n136_), .Y(men_men_n1196_));
  NO4        u1168(.A(men_men_n1196_), .B(men_men_n1192_), .C(men_men_n1184_), .D(men_men_n1182_), .Y(men_men_n1197_));
  NA2        u1169(.A(men_men_n296_), .B(men_men_n515_), .Y(men_men_n1198_));
  NA2        u1170(.A(men_men_n523_), .B(men_men_n387_), .Y(men_men_n1199_));
  NOi21      u1171(.An(men_men_n547_), .B(men_men_n569_), .Y(men_men_n1200_));
  NA2        u1172(.A(men_men_n1200_), .B(men_men_n1199_), .Y(men_men_n1201_));
  AN3        u1173(.A(m), .B(l), .C(k), .Y(men_men_n1202_));
  OAI210     u1174(.A0(men_men_n349_), .A1(men_men_n34_), .B0(men_men_n1202_), .Y(men_men_n1203_));
  NA2        u1175(.A(men_men_n200_), .B(men_men_n34_), .Y(men_men_n1204_));
  AO210      u1176(.A0(men_men_n1204_), .A1(men_men_n1203_), .B0(men_men_n324_), .Y(men_men_n1205_));
  NA3        u1177(.A(men_men_n1205_), .B(men_men_n1201_), .C(men_men_n1198_), .Y(men_men_n1206_));
  AOI210     u1178(.A0(men_men_n584_), .A1(men_men_n116_), .B0(men_men_n590_), .Y(men_men_n1207_));
  OAI210     u1179(.A0(men_men_n1190_), .A1(men_men_n581_), .B0(men_men_n1207_), .Y(men_men_n1208_));
  NA2        u1180(.A(men_men_n273_), .B(men_men_n192_), .Y(men_men_n1209_));
  NA2        u1181(.A(men_men_n1209_), .B(men_men_n650_), .Y(men_men_n1210_));
  NO3        u1182(.A(men_men_n806_), .B(men_men_n201_), .C(men_men_n396_), .Y(men_men_n1211_));
  NO2        u1183(.A(men_men_n1211_), .B(men_men_n932_), .Y(men_men_n1212_));
  OAI210     u1184(.A0(men_men_n1187_), .A1(men_men_n318_), .B0(men_men_n662_), .Y(men_men_n1213_));
  NA4        u1185(.A(men_men_n1213_), .B(men_men_n1212_), .C(men_men_n1210_), .D(men_men_n770_), .Y(men_men_n1214_));
  NO3        u1186(.A(men_men_n1214_), .B(men_men_n1208_), .C(men_men_n1206_), .Y(men_men_n1215_));
  NA2        u1187(.A(men_men_n488_), .B(men_men_n56_), .Y(men_men_n1216_));
  OR3        u1188(.A(men_men_n1186_), .B(men_men_n594_), .C(men_men_n1185_), .Y(men_men_n1217_));
  NO2        u1189(.A(men_men_n1194_), .B(men_men_n947_), .Y(men_men_n1218_));
  NO2        u1190(.A(men_men_n1218_), .B(men_men_n1131_), .Y(men_men_n1219_));
  NA4        u1191(.A(men_men_n1219_), .B(men_men_n1217_), .C(men_men_n1216_), .D(men_men_n742_), .Y(men_men_n1220_));
  NO2        u1192(.A(men_men_n938_), .B(men_men_n226_), .Y(men_men_n1221_));
  NO2        u1193(.A(men_men_n939_), .B(men_men_n540_), .Y(men_men_n1222_));
  OAI210     u1194(.A0(men_men_n1222_), .A1(men_men_n1221_), .B0(men_men_n333_), .Y(men_men_n1223_));
  NA2        u1195(.A(men_men_n557_), .B(men_men_n555_), .Y(men_men_n1224_));
  NO3        u1196(.A(men_men_n79_), .B(men_men_n294_), .C(men_men_n43_), .Y(men_men_n1225_));
  NA2        u1197(.A(men_men_n1225_), .B(men_men_n539_), .Y(men_men_n1226_));
  NA3        u1198(.A(men_men_n1226_), .B(men_men_n1224_), .C(men_men_n656_), .Y(men_men_n1227_));
  INV        u1199(.A(men_men_n377_), .Y(men_men_n1228_));
  NOi41      u1200(.An(men_men_n1223_), .B(men_men_n1228_), .C(men_men_n1227_), .D(men_men_n1220_), .Y(men_men_n1229_));
  NO2        u1201(.A(men_men_n129_), .B(men_men_n43_), .Y(men_men_n1230_));
  NO2        u1202(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n1231_));
  AO220      u1203(.A0(men_men_n1231_), .A1(men_men_n614_), .B0(men_men_n1230_), .B1(men_men_n693_), .Y(men_men_n1232_));
  NA2        u1204(.A(men_men_n1232_), .B(men_men_n333_), .Y(men_men_n1233_));
  NO3        u1205(.A(men_men_n1056_), .B(men_men_n175_), .C(men_men_n86_), .Y(men_men_n1234_));
  INV        u1206(.A(men_men_n1233_), .Y(men_men_n1235_));
  NO2        u1207(.A(men_men_n605_), .B(men_men_n604_), .Y(men_men_n1236_));
  NO4        u1208(.A(men_men_n1056_), .B(men_men_n1236_), .C(men_men_n173_), .D(men_men_n86_), .Y(men_men_n1237_));
  NO3        u1209(.A(men_men_n1237_), .B(men_men_n1235_), .C(men_men_n630_), .Y(men_men_n1238_));
  NA4        u1210(.A(men_men_n1238_), .B(men_men_n1229_), .C(men_men_n1215_), .D(men_men_n1197_), .Y(men06));
  NO2        u1211(.A(men_men_n397_), .B(men_men_n544_), .Y(men_men_n1240_));
  INV        u1212(.A(men_men_n717_), .Y(men_men_n1241_));
  OAI210     u1213(.A0(men_men_n1241_), .A1(men_men_n264_), .B0(men_men_n1240_), .Y(men_men_n1242_));
  NO2        u1214(.A(men_men_n218_), .B(men_men_n103_), .Y(men_men_n1243_));
  OAI210     u1215(.A0(men_men_n1243_), .A1(men_men_n1234_), .B0(men_men_n373_), .Y(men_men_n1244_));
  NO3        u1216(.A(men_men_n588_), .B(men_men_n793_), .C(men_men_n591_), .Y(men_men_n1245_));
  OR2        u1217(.A(men_men_n1245_), .B(men_men_n869_), .Y(men_men_n1246_));
  NA4        u1218(.A(men_men_n1246_), .B(men_men_n1244_), .C(men_men_n1242_), .D(men_men_n1223_), .Y(men_men_n1247_));
  NO3        u1219(.A(men_men_n1247_), .B(men_men_n1227_), .C(men_men_n252_), .Y(men_men_n1248_));
  INV        u1220(.A(men_men_n1221_), .Y(men_men_n1249_));
  INV        u1221(.A(men_men_n1232_), .Y(men_men_n1250_));
  AOI210     u1222(.A0(men_men_n1250_), .A1(men_men_n1249_), .B0(men_men_n330_), .Y(men_men_n1251_));
  INV        u1223(.A(men_men_n660_), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n1252_), .B(men_men_n634_), .Y(men_men_n1253_));
  NOi21      u1225(.An(men_men_n135_), .B(men_men_n43_), .Y(men_men_n1254_));
  NO2        u1226(.A(men_men_n598_), .B(men_men_n1078_), .Y(men_men_n1255_));
  OAI210     u1227(.A0(men_men_n449_), .A1(men_men_n243_), .B0(men_men_n887_), .Y(men_men_n1256_));
  NO3        u1228(.A(men_men_n1256_), .B(men_men_n1255_), .C(men_men_n1254_), .Y(men_men_n1257_));
  OR2        u1229(.A(men_men_n589_), .B(men_men_n587_), .Y(men_men_n1258_));
  INV        u1230(.A(men_men_n1258_), .Y(men_men_n1259_));
  NA3        u1231(.A(men_men_n1259_), .B(men_men_n1257_), .C(men_men_n1253_), .Y(men_men_n1260_));
  NO2        u1232(.A(men_men_n733_), .B(men_men_n359_), .Y(men_men_n1261_));
  NO3        u1233(.A(men_men_n662_), .B(men_men_n744_), .C(men_men_n626_), .Y(men_men_n1262_));
  NOi21      u1234(.An(men_men_n1261_), .B(men_men_n1262_), .Y(men_men_n1263_));
  NO3        u1235(.A(men_men_n1263_), .B(men_men_n1260_), .C(men_men_n1251_), .Y(men_men_n1264_));
  NO2        u1236(.A(men_men_n787_), .B(men_men_n271_), .Y(men_men_n1265_));
  OAI220     u1237(.A0(men_men_n717_), .A1(men_men_n45_), .B0(men_men_n218_), .B1(men_men_n607_), .Y(men_men_n1266_));
  OAI210     u1238(.A0(men_men_n271_), .A1(c), .B0(men_men_n633_), .Y(men_men_n1267_));
  AOI220     u1239(.A0(men_men_n1267_), .A1(men_men_n1266_), .B0(men_men_n1265_), .B1(men_men_n264_), .Y(men_men_n1268_));
  OAI220     u1240(.A0(men_men_n687_), .A1(men_men_n243_), .B0(men_men_n495_), .B1(men_men_n499_), .Y(men_men_n1269_));
  OAI210     u1241(.A0(l), .A1(i), .B0(k), .Y(men_men_n1270_));
  NO3        u1242(.A(men_men_n1270_), .B(men_men_n586_), .C(j), .Y(men_men_n1271_));
  NOi21      u1243(.An(men_men_n1271_), .B(men_men_n654_), .Y(men_men_n1272_));
  NO3        u1244(.A(men_men_n1272_), .B(men_men_n1269_), .C(men_men_n1081_), .Y(men_men_n1273_));
  NA3        u1245(.A(men_men_n1273_), .B(men_men_n1268_), .C(men_men_n1168_), .Y(men_men_n1274_));
  NOi31      u1246(.An(men_men_n1245_), .B(men_men_n453_), .C(men_men_n386_), .Y(men_men_n1275_));
  OR3        u1247(.A(men_men_n1275_), .B(men_men_n766_), .C(men_men_n526_), .Y(men_men_n1276_));
  OR3        u1248(.A(men_men_n362_), .B(men_men_n218_), .C(men_men_n607_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n557_), .B(men_men_n435_), .Y(men_men_n1278_));
  NA2        u1250(.A(men_men_n1271_), .B(men_men_n774_), .Y(men_men_n1279_));
  NA4        u1251(.A(men_men_n1279_), .B(men_men_n1278_), .C(men_men_n1277_), .D(men_men_n1276_), .Y(men_men_n1280_));
  NA2        u1252(.A(men_men_n1261_), .B(men_men_n743_), .Y(men_men_n1281_));
  AN2        u1253(.A(men_men_n905_), .B(men_men_n904_), .Y(men_men_n1282_));
  NO3        u1254(.A(men_men_n1282_), .B(men_men_n859_), .C(men_men_n472_), .Y(men_men_n1283_));
  NA2        u1255(.A(men_men_n1283_), .B(men_men_n1281_), .Y(men_men_n1284_));
  NAi21      u1256(.An(j), .B(i), .Y(men_men_n1285_));
  NO4        u1257(.A(men_men_n1236_), .B(men_men_n1285_), .C(men_men_n429_), .D(men_men_n229_), .Y(men_men_n1286_));
  NO4        u1258(.A(men_men_n1286_), .B(men_men_n1284_), .C(men_men_n1280_), .D(men_men_n1274_), .Y(men_men_n1287_));
  NA4        u1259(.A(men_men_n1287_), .B(men_men_n1264_), .C(men_men_n1248_), .D(men_men_n1238_), .Y(men07));
  NAi32      u1260(.An(m), .Bn(b), .C(n), .Y(men_men_n1289_));
  NO3        u1261(.A(men_men_n1289_), .B(g), .C(f), .Y(men_men_n1290_));
  OAI210     u1262(.A0(men_men_n312_), .A1(men_men_n473_), .B0(men_men_n1290_), .Y(men_men_n1291_));
  NAi21      u1263(.An(f), .B(c), .Y(men_men_n1292_));
  OR2        u1264(.A(e), .B(d), .Y(men_men_n1293_));
  NOi31      u1265(.An(n), .B(m), .C(b), .Y(men_men_n1294_));
  INV        u1266(.A(men_men_n1291_), .Y(men_men_n1295_));
  NOi41      u1267(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1296_));
  NA2        u1268(.A(men_men_n1058_), .B(men_men_n215_), .Y(men_men_n1297_));
  NO2        u1269(.A(men_men_n1297_), .B(men_men_n59_), .Y(men_men_n1298_));
  NO2        u1270(.A(k), .B(i), .Y(men_men_n1299_));
  NA2        u1271(.A(men_men_n86_), .B(men_men_n43_), .Y(men_men_n1300_));
  NO2        u1272(.A(men_men_n1016_), .B(men_men_n429_), .Y(men_men_n1301_));
  NA3        u1273(.A(men_men_n1301_), .B(men_men_n1300_), .C(men_men_n208_), .Y(men_men_n1302_));
  NO2        u1274(.A(men_men_n1030_), .B(men_men_n301_), .Y(men_men_n1303_));
  NA2        u1275(.A(men_men_n1169_), .B(men_men_n284_), .Y(men_men_n1304_));
  NA2        u1276(.A(men_men_n1304_), .B(men_men_n1302_), .Y(men_men_n1305_));
  NO3        u1277(.A(men_men_n1305_), .B(men_men_n1298_), .C(men_men_n1295_), .Y(men_men_n1306_));
  NO3        u1278(.A(e), .B(d), .C(c), .Y(men_men_n1307_));
  OAI210     u1279(.A0(men_men_n130_), .A1(men_men_n208_), .B0(men_men_n595_), .Y(men_men_n1308_));
  NA2        u1280(.A(men_men_n1308_), .B(men_men_n1307_), .Y(men_men_n1309_));
  INV        u1281(.A(men_men_n1309_), .Y(men_men_n1310_));
  OR2        u1282(.A(h), .B(f), .Y(men_men_n1311_));
  NO3        u1283(.A(n), .B(m), .C(i), .Y(men_men_n1312_));
  OAI210     u1284(.A0(men_men_n1079_), .A1(men_men_n156_), .B0(men_men_n1312_), .Y(men_men_n1313_));
  NO2        u1285(.A(i), .B(g), .Y(men_men_n1314_));
  OR3        u1286(.A(men_men_n1314_), .B(men_men_n1289_), .C(men_men_n70_), .Y(men_men_n1315_));
  OAI220     u1287(.A0(men_men_n1315_), .A1(men_men_n473_), .B0(men_men_n1313_), .B1(men_men_n1311_), .Y(men_men_n1316_));
  NA3        u1288(.A(men_men_n684_), .B(men_men_n670_), .C(men_men_n110_), .Y(men_men_n1317_));
  NA3        u1289(.A(men_men_n1294_), .B(men_men_n1025_), .C(men_men_n658_), .Y(men_men_n1318_));
  AOI210     u1290(.A0(men_men_n1318_), .A1(men_men_n1317_), .B0(men_men_n43_), .Y(men_men_n1319_));
  NA2        u1291(.A(men_men_n1312_), .B(men_men_n632_), .Y(men_men_n1320_));
  NO2        u1292(.A(l), .B(k), .Y(men_men_n1321_));
  NO3        u1293(.A(men_men_n429_), .B(d), .C(c), .Y(men_men_n1322_));
  NO3        u1294(.A(men_men_n1319_), .B(men_men_n1316_), .C(men_men_n1310_), .Y(men_men_n1323_));
  NO2        u1295(.A(men_men_n146_), .B(h), .Y(men_men_n1324_));
  NO2        u1296(.A(i), .B(l), .Y(men_men_n1325_));
  NO2        u1297(.A(g), .B(c), .Y(men_men_n1326_));
  NA3        u1298(.A(men_men_n1326_), .B(men_men_n141_), .C(men_men_n183_), .Y(men_men_n1327_));
  NO2        u1299(.A(men_men_n1327_), .B(men_men_n1325_), .Y(men_men_n1328_));
  NA2        u1300(.A(men_men_n1328_), .B(men_men_n178_), .Y(men_men_n1329_));
  NO2        u1301(.A(men_men_n440_), .B(a), .Y(men_men_n1330_));
  NA3        u1302(.A(men_men_n1330_), .B(k), .C(men_men_n111_), .Y(men_men_n1331_));
  NO2        u1303(.A(i), .B(h), .Y(men_men_n1332_));
  NA2        u1304(.A(men_men_n1332_), .B(men_men_n215_), .Y(men_men_n1333_));
  NA2        u1305(.A(men_men_n1101_), .B(h), .Y(men_men_n1334_));
  NA2        u1306(.A(men_men_n137_), .B(men_men_n215_), .Y(men_men_n1335_));
  AOI210     u1307(.A0(men_men_n253_), .A1(men_men_n114_), .B0(men_men_n515_), .Y(men_men_n1336_));
  OAI220     u1308(.A0(men_men_n1336_), .A1(men_men_n1333_), .B0(men_men_n1335_), .B1(men_men_n1334_), .Y(men_men_n1337_));
  NO2        u1309(.A(men_men_n740_), .B(men_men_n184_), .Y(men_men_n1338_));
  NOi31      u1310(.An(m), .B(n), .C(b), .Y(men_men_n1339_));
  NOi31      u1311(.An(f), .B(d), .C(c), .Y(men_men_n1340_));
  NA2        u1312(.A(men_men_n1340_), .B(men_men_n1339_), .Y(men_men_n1341_));
  INV        u1313(.A(men_men_n1341_), .Y(men_men_n1342_));
  NO3        u1314(.A(men_men_n1342_), .B(men_men_n1338_), .C(men_men_n1337_), .Y(men_men_n1343_));
  NA2        u1315(.A(men_men_n1049_), .B(men_men_n456_), .Y(men_men_n1344_));
  NO4        u1316(.A(men_men_n1344_), .B(men_men_n1025_), .C(men_men_n429_), .D(men_men_n43_), .Y(men_men_n1345_));
  OAI210     u1317(.A0(men_men_n181_), .A1(men_men_n510_), .B0(men_men_n1026_), .Y(men_men_n1346_));
  NO3        u1318(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1347_));
  INV        u1319(.A(men_men_n1346_), .Y(men_men_n1348_));
  NO2        u1320(.A(men_men_n1348_), .B(men_men_n1345_), .Y(men_men_n1349_));
  AN4        u1321(.A(men_men_n1349_), .B(men_men_n1343_), .C(men_men_n1331_), .D(men_men_n1329_), .Y(men_men_n1350_));
  NA2        u1322(.A(men_men_n1294_), .B(men_men_n370_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n1351_), .B(men_men_n1007_), .Y(men_men_n1352_));
  NA2        u1324(.A(men_men_n1322_), .B(men_men_n209_), .Y(men_men_n1353_));
  NO2        u1325(.A(men_men_n184_), .B(b), .Y(men_men_n1354_));
  AOI220     u1326(.A0(men_men_n1129_), .A1(men_men_n1354_), .B0(men_men_n1057_), .B1(men_men_n1344_), .Y(men_men_n1355_));
  NO2        u1327(.A(i), .B(men_men_n207_), .Y(men_men_n1356_));
  NA4        u1328(.A(men_men_n1106_), .B(men_men_n1356_), .C(men_men_n104_), .D(m), .Y(men_men_n1357_));
  NAi41      u1329(.An(men_men_n1352_), .B(men_men_n1357_), .C(men_men_n1355_), .D(men_men_n1353_), .Y(men_men_n1358_));
  NO4        u1330(.A(men_men_n130_), .B(g), .C(f), .D(e), .Y(men_men_n1359_));
  NA3        u1331(.A(men_men_n1299_), .B(men_men_n285_), .C(h), .Y(men_men_n1360_));
  OR2        u1332(.A(e), .B(a), .Y(men_men_n1361_));
  NO2        u1333(.A(men_men_n1293_), .B(men_men_n1292_), .Y(men_men_n1362_));
  AOI210     u1334(.A0(men_men_n30_), .A1(h), .B0(men_men_n1362_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n1363_), .B(men_men_n1045_), .Y(men_men_n1364_));
  NA2        u1336(.A(men_men_n1296_), .B(men_men_n1321_), .Y(men_men_n1365_));
  INV        u1337(.A(men_men_n1365_), .Y(men_men_n1366_));
  OR3        u1338(.A(men_men_n526_), .B(men_men_n525_), .C(men_men_n110_), .Y(men_men_n1367_));
  NA2        u1339(.A(men_men_n1077_), .B(men_men_n396_), .Y(men_men_n1368_));
  OAI220     u1340(.A0(men_men_n1368_), .A1(men_men_n422_), .B0(men_men_n1367_), .B1(men_men_n294_), .Y(men_men_n1369_));
  AO210      u1341(.A0(men_men_n1369_), .A1(men_men_n114_), .B0(men_men_n1366_), .Y(men_men_n1370_));
  NO3        u1342(.A(men_men_n1370_), .B(men_men_n1364_), .C(men_men_n1358_), .Y(men_men_n1371_));
  NA4        u1343(.A(men_men_n1371_), .B(men_men_n1350_), .C(men_men_n1323_), .D(men_men_n1306_), .Y(men_men_n1372_));
  NA2        u1344(.A(men_men_n370_), .B(men_men_n54_), .Y(men_men_n1373_));
  AOI210     u1345(.A0(men_men_n1373_), .A1(men_men_n1016_), .B0(men_men_n1320_), .Y(men_men_n1374_));
  NO2        u1346(.A(men_men_n1050_), .B(men_men_n1045_), .Y(men_men_n1375_));
  NO2        u1347(.A(men_men_n1375_), .B(men_men_n1374_), .Y(men_men_n1376_));
  NO2        u1348(.A(men_men_n382_), .B(j), .Y(men_men_n1377_));
  NA3        u1349(.A(men_men_n1347_), .B(men_men_n1293_), .C(men_men_n1077_), .Y(men_men_n1378_));
  NAi41      u1350(.An(men_men_n1332_), .B(men_men_n1038_), .C(men_men_n167_), .D(men_men_n149_), .Y(men_men_n1379_));
  NA2        u1351(.A(men_men_n1379_), .B(men_men_n1378_), .Y(men_men_n1380_));
  NA3        u1352(.A(g), .B(men_men_n1377_), .C(men_men_n158_), .Y(men_men_n1381_));
  INV        u1353(.A(men_men_n1381_), .Y(men_men_n1382_));
  NO3        u1354(.A(men_men_n733_), .B(men_men_n173_), .C(men_men_n399_), .Y(men_men_n1383_));
  NO3        u1355(.A(men_men_n1383_), .B(men_men_n1382_), .C(men_men_n1380_), .Y(men_men_n1384_));
  OR2        u1356(.A(n), .B(i), .Y(men_men_n1385_));
  OAI210     u1357(.A0(men_men_n1385_), .A1(men_men_n1037_), .B0(men_men_n47_), .Y(men_men_n1386_));
  AOI220     u1358(.A0(men_men_n1386_), .A1(men_men_n1135_), .B0(men_men_n811_), .B1(men_men_n191_), .Y(men_men_n1387_));
  INV        u1359(.A(men_men_n1387_), .Y(men_men_n1388_));
  OAI220     u1360(.A0(men_men_n651_), .A1(g), .B0(men_men_n218_), .B1(c), .Y(men_men_n1389_));
  AOI210     u1361(.A0(men_men_n1354_), .A1(men_men_n41_), .B0(men_men_n1389_), .Y(men_men_n1390_));
  NO2        u1362(.A(men_men_n218_), .B(k), .Y(men_men_n1391_));
  NO2        u1363(.A(men_men_n1390_), .B(men_men_n175_), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n1392_), .B(men_men_n1388_), .Y(men_men_n1393_));
  INV        u1365(.A(men_men_n47_), .Y(men_men_n1394_));
  NO3        u1366(.A(men_men_n1060_), .B(men_men_n1293_), .C(men_men_n47_), .Y(men_men_n1395_));
  NA2        u1367(.A(men_men_n1061_), .B(men_men_n1394_), .Y(men_men_n1396_));
  NO2        u1368(.A(men_men_n1045_), .B(h), .Y(men_men_n1397_));
  NA3        u1369(.A(men_men_n1397_), .B(d), .C(men_men_n1008_), .Y(men_men_n1398_));
  OAI220     u1370(.A0(men_men_n1398_), .A1(c), .B0(men_men_n1396_), .B1(j), .Y(men_men_n1399_));
  NA2        u1371(.A(men_men_n178_), .B(men_men_n110_), .Y(men_men_n1400_));
  AOI210     u1372(.A0(men_men_n510_), .A1(h), .B0(men_men_n67_), .Y(men_men_n1401_));
  NA2        u1373(.A(men_men_n1401_), .B(men_men_n1330_), .Y(men_men_n1402_));
  NO2        u1374(.A(men_men_n1285_), .B(men_men_n173_), .Y(men_men_n1403_));
  NOi21      u1375(.An(d), .B(f), .Y(men_men_n1404_));
  NO3        u1376(.A(men_men_n1340_), .B(men_men_n1404_), .C(men_men_n40_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1405_), .B(men_men_n1403_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1293_), .B(f), .Y(men_men_n1407_));
  NO2        u1379(.A(men_men_n294_), .B(c), .Y(men_men_n1408_));
  NA2        u1380(.A(men_men_n1408_), .B(men_men_n527_), .Y(men_men_n1409_));
  NA3        u1381(.A(men_men_n1409_), .B(men_men_n1406_), .C(men_men_n1402_), .Y(men_men_n1410_));
  NO2        u1382(.A(men_men_n1410_), .B(men_men_n1399_), .Y(men_men_n1411_));
  NA4        u1383(.A(men_men_n1411_), .B(men_men_n1393_), .C(men_men_n1384_), .D(men_men_n1376_), .Y(men_men_n1412_));
  NO3        u1384(.A(men_men_n1049_), .B(men_men_n1037_), .C(men_men_n40_), .Y(men_men_n1413_));
  NO2        u1385(.A(men_men_n456_), .B(men_men_n294_), .Y(men_men_n1414_));
  OAI210     u1386(.A0(men_men_n1414_), .A1(men_men_n1413_), .B0(men_men_n1303_), .Y(men_men_n1415_));
  OAI210     u1387(.A0(men_men_n1359_), .A1(men_men_n1294_), .B0(men_men_n866_), .Y(men_men_n1416_));
  OAI220     u1388(.A0(men_men_n1004_), .A1(men_men_n130_), .B0(men_men_n651_), .B1(men_men_n173_), .Y(men_men_n1417_));
  NA2        u1389(.A(men_men_n1417_), .B(men_men_n613_), .Y(men_men_n1418_));
  NA3        u1390(.A(men_men_n1418_), .B(men_men_n1416_), .C(men_men_n1415_), .Y(men_men_n1419_));
  NA2        u1391(.A(men_men_n1326_), .B(men_men_n1404_), .Y(men_men_n1420_));
  NO2        u1392(.A(men_men_n1420_), .B(m), .Y(men_men_n1421_));
  NA3        u1393(.A(men_men_n1058_), .B(men_men_n106_), .C(men_men_n215_), .Y(men_men_n1422_));
  NO2        u1394(.A(men_men_n150_), .B(men_men_n180_), .Y(men_men_n1423_));
  OAI210     u1395(.A0(men_men_n1423_), .A1(men_men_n108_), .B0(men_men_n1339_), .Y(men_men_n1424_));
  NA2        u1396(.A(men_men_n1424_), .B(men_men_n1422_), .Y(men_men_n1425_));
  NO3        u1397(.A(men_men_n1425_), .B(men_men_n1421_), .C(men_men_n1419_), .Y(men_men_n1426_));
  NO2        u1398(.A(men_men_n1292_), .B(e), .Y(men_men_n1427_));
  NA2        u1399(.A(men_men_n1427_), .B(men_men_n394_), .Y(men_men_n1428_));
  NA2        u1400(.A(men_men_n1087_), .B(men_men_n624_), .Y(men_men_n1429_));
  OR3        u1401(.A(men_men_n1391_), .B(men_men_n1169_), .C(men_men_n130_), .Y(men_men_n1430_));
  OAI220     u1402(.A0(men_men_n1430_), .A1(men_men_n1428_), .B0(men_men_n1429_), .B1(men_men_n431_), .Y(men_men_n1431_));
  NO3        u1403(.A(men_men_n1367_), .B(men_men_n345_), .C(a), .Y(men_men_n1432_));
  NO2        u1404(.A(men_men_n1432_), .B(men_men_n1431_), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n180_), .B(c), .Y(men_men_n1434_));
  OAI210     u1406(.A0(men_men_n1434_), .A1(men_men_n1427_), .B0(men_men_n178_), .Y(men_men_n1435_));
  AOI220     u1407(.A0(men_men_n1435_), .A1(men_men_n1039_), .B0(men_men_n517_), .B1(men_men_n359_), .Y(men_men_n1436_));
  NA2        u1408(.A(men_men_n525_), .B(g), .Y(men_men_n1437_));
  AOI210     u1409(.A0(men_men_n1437_), .A1(men_men_n1322_), .B0(men_men_n1395_), .Y(men_men_n1438_));
  NO2        u1410(.A(men_men_n1361_), .B(f), .Y(men_men_n1439_));
  AOI210     u1411(.A0(men_men_n1087_), .A1(a), .B0(men_men_n1439_), .Y(men_men_n1440_));
  OAI220     u1412(.A0(men_men_n1440_), .A1(men_men_n67_), .B0(men_men_n1438_), .B1(men_men_n207_), .Y(men_men_n1441_));
  NA2        u1413(.A(men_men_n881_), .B(men_men_n406_), .Y(men_men_n1442_));
  OR2        u1414(.A(men_men_n1442_), .B(men_men_n525_), .Y(men_men_n1443_));
  NO2        u1415(.A(men_men_n1443_), .B(men_men_n173_), .Y(men_men_n1444_));
  NO2        u1416(.A(men_men_n47_), .B(l), .Y(men_men_n1445_));
  OAI210     u1417(.A0(men_men_n1361_), .A1(men_men_n844_), .B0(men_men_n473_), .Y(men_men_n1446_));
  OAI210     u1418(.A0(men_men_n1446_), .A1(men_men_n1061_), .B0(men_men_n1445_), .Y(men_men_n1447_));
  NO2        u1419(.A(m), .B(i), .Y(men_men_n1448_));
  BUFFER     u1420(.A(men_men_n1448_), .Y(men_men_n1449_));
  NA2        u1421(.A(men_men_n1449_), .B(men_men_n1324_), .Y(men_men_n1450_));
  NA2        u1422(.A(men_men_n1450_), .B(men_men_n1447_), .Y(men_men_n1451_));
  NO4        u1423(.A(men_men_n1451_), .B(men_men_n1444_), .C(men_men_n1441_), .D(men_men_n1436_), .Y(men_men_n1452_));
  NA3        u1424(.A(men_men_n1452_), .B(men_men_n1433_), .C(men_men_n1426_), .Y(men_men_n1453_));
  NA3        u1425(.A(men_men_n934_), .B(men_men_n137_), .C(men_men_n44_), .Y(men_men_n1454_));
  AO210      u1426(.A0(men_men_n131_), .A1(l), .B0(men_men_n1351_), .Y(men_men_n1455_));
  NO2        u1427(.A(men_men_n70_), .B(c), .Y(men_men_n1456_));
  NO4        u1428(.A(men_men_n1311_), .B(men_men_n182_), .C(men_men_n437_), .D(men_men_n43_), .Y(men_men_n1457_));
  AOI210     u1429(.A0(men_men_n1403_), .A1(men_men_n1456_), .B0(men_men_n1457_), .Y(men_men_n1458_));
  NA2        u1430(.A(men_men_n1458_), .B(men_men_n1455_), .Y(men_men_n1459_));
  INV        u1431(.A(men_men_n1459_), .Y(men_men_n1460_));
  NO4        u1432(.A(men_men_n218_), .B(men_men_n182_), .C(men_men_n253_), .D(k), .Y(men_men_n1461_));
  AOI210     u1433(.A0(men_men_n156_), .A1(men_men_n54_), .B0(men_men_n1427_), .Y(men_men_n1462_));
  NO2        u1434(.A(men_men_n1462_), .B(men_men_n1400_), .Y(men_men_n1463_));
  NO2        u1435(.A(men_men_n1454_), .B(men_men_n108_), .Y(men_men_n1464_));
  NO3        u1436(.A(men_men_n1464_), .B(men_men_n1463_), .C(men_men_n1461_), .Y(men_men_n1465_));
  NA2        u1437(.A(men_men_n57_), .B(a), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n1368_), .B(men_men_n1466_), .Y(men_men_n1467_));
  NA3        u1439(.A(men_men_n1481_), .B(men_men_n1465_), .C(men_men_n1460_), .Y(men_men_n1468_));
  OR4        u1440(.A(men_men_n1468_), .B(men_men_n1453_), .C(men_men_n1412_), .D(men_men_n1372_), .Y(men04));
  NOi31      u1441(.An(men_men_n1359_), .B(men_men_n1360_), .C(men_men_n1010_), .Y(men_men_n1470_));
  NA2        u1442(.A(men_men_n1407_), .B(men_men_n811_), .Y(men_men_n1471_));
  NO4        u1443(.A(men_men_n1471_), .B(men_men_n999_), .C(men_men_n474_), .D(j), .Y(men_men_n1472_));
  OR3        u1444(.A(men_men_n1472_), .B(men_men_n1470_), .C(men_men_n1028_), .Y(men_men_n1473_));
  NO3        u1445(.A(men_men_n1300_), .B(men_men_n90_), .C(k), .Y(men_men_n1474_));
  AOI210     u1446(.A0(men_men_n1474_), .A1(men_men_n1021_), .B0(men_men_n1147_), .Y(men_men_n1475_));
  NA2        u1447(.A(men_men_n1475_), .B(men_men_n1173_), .Y(men_men_n1476_));
  NO4        u1448(.A(men_men_n1476_), .B(men_men_n1473_), .C(men_men_n1036_), .D(men_men_n1015_), .Y(men_men_n1477_));
  NA4        u1449(.A(men_men_n1477_), .B(men_men_n1089_), .C(men_men_n1075_), .D(men_men_n1064_), .Y(men05));
  INV        u1450(.A(men_men_n1467_), .Y(men_men_n1481_));
  INV        u1451(.A(men_men_n269_), .Y(men_men_n1482_));
  INV        u1452(.A(men_men_n880_), .Y(men_men_n1483_));
  INV        u1453(.A(c), .Y(men_men_n1484_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule