library verilog;
use verilog.vl_types.all;
entity demux14_vlg_vec_tst is
end demux14_vlg_vec_tst;
