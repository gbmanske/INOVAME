//Benchmark atmr_5xp1_76_0.125

module atmr_5xp1(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n61_, ori_ori_n65_, ori_ori_n66_, ori_ori_n68_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n64_, mai_mai_n65_, mai_mai_n67_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n62_, men_men_n63_, men_men_n65_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n88_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09;
  INV        o00(.A(i_5_), .Y(ori_ori_n18_));
  NO3        o01(.A(i_4_), .B(i_6_), .C(ori_ori_n18_), .Y(ori_ori_n19_));
  INV        o02(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o03(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n21_));
  INV        o04(.A(i_1_), .Y(ori_ori_n22_));
  AOI210     o05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(ori_ori_n23_));
  NA2        o06(.A(ori_ori_n23_), .B(ori_ori_n22_), .Y(ori_ori_n24_));
  NO2        o07(.A(ori_ori_n24_), .B(ori_ori_n21_), .Y(ori_ori_n25_));
  INV        o08(.A(i_6_), .Y(ori_ori_n26_));
  NO2        o09(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n27_));
  INV        o10(.A(i_0_), .Y(ori_ori_n28_));
  NO2        o11(.A(i_2_), .B(i_1_), .Y(ori_ori_n29_));
  OAI210     o12(.A0(ori_ori_n29_), .A1(ori_ori_n28_), .B0(ori_ori_n20_), .Y(ori_ori_n30_));
  NO2        o13(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n31_));
  NO2        o14(.A(i_2_), .B(i_3_), .Y(ori_ori_n32_));
  NO3        o15(.A(ori_ori_n32_), .B(ori_ori_n28_), .C(ori_ori_n22_), .Y(ori_ori_n33_));
  AO220      o16(.A0(ori_ori_n33_), .A1(ori_ori_n31_), .B0(ori_ori_n30_), .B1(ori_ori_n27_), .Y(ori_ori_n34_));
  NA2        o17(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n35_));
  NA2        o18(.A(i_2_), .B(i_3_), .Y(ori_ori_n36_));
  NO2        o19(.A(ori_ori_n36_), .B(ori_ori_n22_), .Y(ori_ori_n37_));
  NO3        o20(.A(ori_ori_n37_), .B(ori_ori_n35_), .C(i_0_), .Y(ori_ori_n38_));
  OR3        o21(.A(ori_ori_n34_), .B(ori_ori_n25_), .C(ori_ori_n19_), .Y(ori01));
  NA2        o22(.A(i_0_), .B(i_1_), .Y(ori_ori_n40_));
  NA2        o23(.A(ori_ori_n28_), .B(ori_ori_n18_), .Y(ori_ori_n41_));
  AOI210     o24(.A0(ori_ori_n23_), .A1(ori_ori_n22_), .B0(ori_ori_n26_), .Y(ori_ori_n42_));
  AOI220     o25(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n40_), .B1(ori_ori_n26_), .Y(ori_ori_n43_));
  NA2        o26(.A(ori_ori_n29_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  OAI220     o27(.A0(ori_ori_n44_), .A1(ori_ori_n26_), .B0(ori_ori_n35_), .B1(ori_ori_n28_), .Y(ori_ori_n45_));
  NO3        o28(.A(ori_ori_n45_), .B(ori_ori_n43_), .C(i_4_), .Y(ori_ori_n46_));
  NA2        o29(.A(i_0_), .B(i_6_), .Y(ori_ori_n47_));
  OAI210     o30(.A0(i_0_), .A1(i_1_), .B0(ori_ori_n47_), .Y(ori_ori_n48_));
  NOi31      o31(.An(ori_ori_n48_), .B(ori_ori_n23_), .C(ori_ori_n18_), .Y(ori_ori_n49_));
  NA3        o32(.A(i_1_), .B(i_6_), .C(i_5_), .Y(ori_ori_n50_));
  AOI210     o33(.A0(ori_ori_n50_), .A1(ori_ori_n47_), .B0(ori_ori_n29_), .Y(ori_ori_n51_));
  NO3        o34(.A(ori_ori_n51_), .B(ori_ori_n49_), .C(ori_ori_n20_), .Y(ori_ori_n52_));
  AOI210     o35(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(ori_ori_n53_));
  AO220      o36(.A0(ori_ori_n53_), .A1(ori_ori_n31_), .B0(ori_ori_n37_), .B1(ori_ori_n19_), .Y(ori_ori_n54_));
  INV        o37(.A(ori_ori_n54_), .Y(ori_ori_n55_));
  OAI210     o38(.A0(ori_ori_n52_), .A1(ori_ori_n46_), .B0(ori_ori_n55_), .Y(ori02));
  NAi21      o39(.An(ori_ori_n21_), .B(ori_ori_n42_), .Y(ori_ori_n57_));
  NA3        o40(.A(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n58_));
  INV        o41(.A(ori_ori_n31_), .Y(ori_ori_n59_));
  NA2        o42(.A(ori_ori_n59_), .B(ori_ori_n57_), .Y(ori00));
  INV        o43(.A(i_5_), .Y(ori_ori_n61_));
  NO2        o44(.A(ori_ori_n61_), .B(ori_ori_n20_), .Y(ori09));
  NOi21      o45(.An(ori_ori_n36_), .B(ori_ori_n32_), .Y(ori07));
  INV        o46(.A(i_3_), .Y(ori08));
  INV        o47(.A(ori_ori_n29_), .Y(ori_ori_n65_));
  NA2        o48(.A(ori07), .B(ori_ori_n65_), .Y(ori_ori_n66_));
  XO2        o49(.A(ori_ori_n66_), .B(ori_ori_n28_), .Y(ori05));
  NO2        o50(.A(i_2_), .B(ori08), .Y(ori_ori_n68_));
  XO2        o51(.A(ori_ori_n68_), .B(i_1_), .Y(ori06));
  INV        o52(.A(ori_ori_n44_), .Y(ori_ori_n70_));
  NA2        o53(.A(ori_ori_n70_), .B(i_0_), .Y(ori_ori_n71_));
  NO2        o54(.A(i_1_), .B(i_6_), .Y(ori_ori_n72_));
  NO3        o55(.A(ori_ori_n72_), .B(ori_ori_n41_), .C(ori_ori_n36_), .Y(ori_ori_n73_));
  NO2        o56(.A(ori_ori_n73_), .B(ori_ori_n38_), .Y(ori_ori_n74_));
  AO210      o57(.A0(ori_ori_n40_), .A1(ori_ori_n24_), .B0(ori_ori_n18_), .Y(ori_ori_n75_));
  OAI210     o58(.A0(ori_ori_n22_), .A1(i_6_), .B0(ori_ori_n18_), .Y(ori_ori_n76_));
  NO2        o59(.A(ori_ori_n76_), .B(ori_ori_n48_), .Y(ori_ori_n77_));
  INV        o60(.A(ori_ori_n77_), .Y(ori_ori_n78_));
  NA4        o61(.A(ori_ori_n78_), .B(ori_ori_n75_), .C(ori_ori_n74_), .D(ori_ori_n71_), .Y(ori03));
  NA2        o62(.A(ori_ori_n28_), .B(ori08), .Y(ori_ori_n80_));
  OAI210     o63(.A0(ori_ori_n80_), .A1(i_1_), .B0(ori_ori_n58_), .Y(ori_ori_n81_));
  OAI210     o64(.A0(ori_ori_n81_), .A1(ori_ori_n33_), .B0(i_6_), .Y(ori_ori_n82_));
  AOI210     o65(.A0(ori_ori_n32_), .A1(ori_ori_n26_), .B0(ori_ori_n29_), .Y(ori_ori_n83_));
  OR2        o66(.A(ori_ori_n83_), .B(ori_ori_n72_), .Y(ori_ori_n84_));
  NA3        o67(.A(ori_ori_n80_), .B(ori_ori_n72_), .C(i_2_), .Y(ori_ori_n85_));
  NA3        o68(.A(ori_ori_n23_), .B(i_1_), .C(ori_ori_n26_), .Y(ori_ori_n86_));
  NA4        o69(.A(ori_ori_n86_), .B(ori_ori_n85_), .C(ori_ori_n84_), .D(ori_ori_n82_), .Y(ori04));
  INV        m00(.A(i_5_), .Y(mai_mai_n18_));
  NO3        m01(.A(i_4_), .B(i_6_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m02(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m03(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n21_));
  INV        m04(.A(i_1_), .Y(mai_mai_n22_));
  AOI210     m05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(mai_mai_n23_));
  NA2        m06(.A(mai_mai_n23_), .B(mai_mai_n22_), .Y(mai_mai_n24_));
  NO2        m07(.A(mai_mai_n24_), .B(mai_mai_n21_), .Y(mai_mai_n25_));
  INV        m08(.A(i_6_), .Y(mai_mai_n26_));
  NO2        m09(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n27_));
  INV        m10(.A(i_0_), .Y(mai_mai_n28_));
  NO2        m11(.A(i_2_), .B(i_1_), .Y(mai_mai_n29_));
  OAI210     m12(.A0(mai_mai_n29_), .A1(mai_mai_n28_), .B0(mai_mai_n20_), .Y(mai_mai_n30_));
  NO2        m13(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n31_));
  NO2        m14(.A(i_2_), .B(i_3_), .Y(mai_mai_n32_));
  NO3        m15(.A(mai_mai_n32_), .B(mai_mai_n28_), .C(mai_mai_n22_), .Y(mai_mai_n33_));
  AN2        m16(.A(mai_mai_n30_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  NA2        m17(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n35_));
  NA2        m18(.A(i_2_), .B(i_3_), .Y(mai_mai_n36_));
  NO2        m19(.A(mai_mai_n35_), .B(i_0_), .Y(mai_mai_n37_));
  OR4        m20(.A(mai_mai_n37_), .B(mai_mai_n34_), .C(mai_mai_n25_), .D(mai_mai_n19_), .Y(mai01));
  NA2        m21(.A(mai_mai_n28_), .B(mai_mai_n18_), .Y(mai_mai_n39_));
  AOI210     m22(.A0(mai_mai_n23_), .A1(mai_mai_n22_), .B0(mai_mai_n26_), .Y(mai_mai_n40_));
  AOI210     m23(.A0(mai_mai_n40_), .A1(mai_mai_n39_), .B0(mai_mai_n26_), .Y(mai_mai_n41_));
  NA2        m24(.A(mai_mai_n29_), .B(mai_mai_n18_), .Y(mai_mai_n42_));
  OAI220     m25(.A0(mai_mai_n42_), .A1(mai_mai_n26_), .B0(mai_mai_n35_), .B1(mai_mai_n28_), .Y(mai_mai_n43_));
  NO3        m26(.A(mai_mai_n43_), .B(mai_mai_n41_), .C(i_4_), .Y(mai_mai_n44_));
  NA2        m27(.A(i_0_), .B(i_6_), .Y(mai_mai_n45_));
  OAI210     m28(.A0(i_0_), .A1(i_1_), .B0(mai_mai_n45_), .Y(mai_mai_n46_));
  NOi31      m29(.An(mai_mai_n46_), .B(mai_mai_n23_), .C(mai_mai_n18_), .Y(mai_mai_n47_));
  NA3        m30(.A(i_1_), .B(i_6_), .C(i_5_), .Y(mai_mai_n48_));
  AOI210     m31(.A0(mai_mai_n48_), .A1(mai_mai_n45_), .B0(mai_mai_n29_), .Y(mai_mai_n49_));
  NO2        m32(.A(i_6_), .B(i_5_), .Y(mai_mai_n50_));
  NO4        m33(.A(mai_mai_n50_), .B(mai_mai_n49_), .C(mai_mai_n47_), .D(mai_mai_n20_), .Y(mai_mai_n51_));
  NA2        m34(.A(mai_mai_n28_), .B(mai_mai_n26_), .Y(mai_mai_n52_));
  NO2        m35(.A(mai_mai_n52_), .B(mai_mai_n20_), .Y(mai_mai_n53_));
  INV        m36(.A(mai_mai_n53_), .Y(mai_mai_n54_));
  OAI210     m37(.A0(mai_mai_n51_), .A1(mai_mai_n44_), .B0(mai_mai_n54_), .Y(mai02));
  NAi21      m38(.An(mai_mai_n21_), .B(mai_mai_n40_), .Y(mai_mai_n56_));
  NA3        m39(.A(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n57_));
  NO2        m40(.A(mai_mai_n53_), .B(mai_mai_n31_), .Y(mai_mai_n58_));
  NA2        m41(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai00));
  NA2        m42(.A(mai_mai_n52_), .B(i_5_), .Y(mai_mai_n60_));
  NO2        m43(.A(mai_mai_n60_), .B(mai_mai_n20_), .Y(mai09));
  NOi21      m44(.An(mai_mai_n36_), .B(mai_mai_n32_), .Y(mai07));
  INV        m45(.A(i_3_), .Y(mai08));
  INV        m46(.A(mai_mai_n29_), .Y(mai_mai_n64_));
  NA2        m47(.A(mai07), .B(mai_mai_n64_), .Y(mai_mai_n65_));
  XO2        m48(.A(mai_mai_n65_), .B(mai_mai_n28_), .Y(mai05));
  NO2        m49(.A(i_2_), .B(mai08), .Y(mai_mai_n67_));
  XO2        m50(.A(mai_mai_n67_), .B(i_1_), .Y(mai06));
  NAi21      m51(.An(mai_mai_n50_), .B(mai_mai_n42_), .Y(mai_mai_n69_));
  NA2        m52(.A(mai_mai_n69_), .B(i_0_), .Y(mai_mai_n70_));
  NO2        m53(.A(i_1_), .B(i_6_), .Y(mai_mai_n71_));
  NO3        m54(.A(mai_mai_n71_), .B(mai_mai_n39_), .C(mai_mai_n36_), .Y(mai_mai_n72_));
  NO2        m55(.A(mai_mai_n72_), .B(mai_mai_n37_), .Y(mai_mai_n73_));
  OR2        m56(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n74_));
  NO2        m57(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n75_));
  NO2        m58(.A(mai_mai_n26_), .B(mai_mai_n18_), .Y(mai_mai_n76_));
  OAI210     m59(.A0(mai_mai_n22_), .A1(i_6_), .B0(mai_mai_n18_), .Y(mai_mai_n77_));
  NO2        m60(.A(mai_mai_n77_), .B(mai_mai_n46_), .Y(mai_mai_n78_));
  AOI210     m61(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  NA4        m62(.A(mai_mai_n79_), .B(mai_mai_n74_), .C(mai_mai_n73_), .D(mai_mai_n70_), .Y(mai03));
  NA2        m63(.A(mai_mai_n28_), .B(mai08), .Y(mai_mai_n81_));
  OAI210     m64(.A0(mai_mai_n81_), .A1(i_1_), .B0(mai_mai_n57_), .Y(mai_mai_n82_));
  OAI210     m65(.A0(mai_mai_n82_), .A1(mai_mai_n33_), .B0(i_6_), .Y(mai_mai_n83_));
  NO2        m66(.A(mai_mai_n26_), .B(mai_mai_n29_), .Y(mai_mai_n84_));
  OR2        m67(.A(mai_mai_n84_), .B(mai_mai_n71_), .Y(mai_mai_n85_));
  NA3        m68(.A(mai_mai_n81_), .B(mai_mai_n71_), .C(i_2_), .Y(mai_mai_n86_));
  NA3        m69(.A(mai_mai_n86_), .B(mai_mai_n85_), .C(mai_mai_n83_), .Y(mai04));
  INV        u00(.A(i_5_), .Y(men_men_n18_));
  NO3        u01(.A(i_4_), .B(i_6_), .C(men_men_n18_), .Y(men_men_n19_));
  INV        u02(.A(i_4_), .Y(men_men_n20_));
  NA2        u03(.A(men_men_n20_), .B(i_5_), .Y(men_men_n21_));
  INV        u04(.A(i_1_), .Y(men_men_n22_));
  AOI210     u05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(men_men_n23_));
  INV        u06(.A(i_6_), .Y(men_men_n24_));
  NO2        u07(.A(men_men_n24_), .B(i_5_), .Y(men_men_n25_));
  INV        u08(.A(i_0_), .Y(men_men_n26_));
  NO2        u09(.A(i_2_), .B(i_1_), .Y(men_men_n27_));
  OAI210     u10(.A0(men_men_n27_), .A1(men_men_n26_), .B0(men_men_n20_), .Y(men_men_n28_));
  NO2        u11(.A(men_men_n20_), .B(i_5_), .Y(men_men_n29_));
  NO2        u12(.A(i_2_), .B(i_3_), .Y(men_men_n30_));
  NO3        u13(.A(men_men_n30_), .B(men_men_n26_), .C(men_men_n22_), .Y(men_men_n31_));
  AO220      u14(.A0(men_men_n31_), .A1(men_men_n29_), .B0(men_men_n28_), .B1(men_men_n25_), .Y(men_men_n32_));
  NA2        u15(.A(men_men_n24_), .B(i_5_), .Y(men_men_n33_));
  NA2        u16(.A(i_2_), .B(i_3_), .Y(men_men_n34_));
  NO2        u17(.A(men_men_n34_), .B(men_men_n22_), .Y(men_men_n35_));
  NO3        u18(.A(men_men_n35_), .B(men_men_n33_), .C(i_0_), .Y(men_men_n36_));
  OR3        u19(.A(men_men_n36_), .B(men_men_n32_), .C(men_men_n19_), .Y(men01));
  OR2        u20(.A(i_2_), .B(i_3_), .Y(men_men_n38_));
  NA3        u21(.A(men_men_n38_), .B(i_0_), .C(i_1_), .Y(men_men_n39_));
  NA2        u22(.A(men_men_n26_), .B(men_men_n18_), .Y(men_men_n40_));
  AOI220     u23(.A0(i_6_), .A1(men_men_n40_), .B0(men_men_n39_), .B1(men_men_n24_), .Y(men_men_n41_));
  NO2        u24(.A(men_men_n33_), .B(men_men_n26_), .Y(men_men_n42_));
  NO3        u25(.A(men_men_n42_), .B(men_men_n41_), .C(i_4_), .Y(men_men_n43_));
  NA2        u26(.A(i_0_), .B(i_6_), .Y(men_men_n44_));
  OAI210     u27(.A0(i_0_), .A1(i_1_), .B0(men_men_n44_), .Y(men_men_n45_));
  NO3        u28(.A(men_men_n38_), .B(i_6_), .C(i_5_), .Y(men_men_n46_));
  NO3        u29(.A(men_men_n46_), .B(men_men_n88_), .C(men_men_n20_), .Y(men_men_n47_));
  NA2        u30(.A(men_men_n26_), .B(men_men_n24_), .Y(men_men_n48_));
  NO2        u31(.A(men_men_n48_), .B(men_men_n20_), .Y(men_men_n49_));
  AOI210     u32(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(men_men_n50_));
  AO220      u33(.A0(men_men_n50_), .A1(men_men_n29_), .B0(men_men_n35_), .B1(men_men_n19_), .Y(men_men_n51_));
  AOI210     u34(.A0(men_men_n49_), .A1(men_men_n34_), .B0(men_men_n51_), .Y(men_men_n52_));
  OAI210     u35(.A0(men_men_n47_), .A1(men_men_n43_), .B0(men_men_n52_), .Y(men02));
  NAi21      u36(.An(men_men_n21_), .B(i_6_), .Y(men_men_n54_));
  NA3        u37(.A(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n55_));
  AOI210     u38(.A0(men_men_n49_), .A1(men_men_n55_), .B0(men_men_n29_), .Y(men_men_n56_));
  NA2        u39(.A(men_men_n56_), .B(men_men_n54_), .Y(men00));
  OAI210     u40(.A0(men_men_n48_), .A1(men_men_n35_), .B0(i_5_), .Y(men_men_n58_));
  NO2        u41(.A(men_men_n58_), .B(men_men_n20_), .Y(men09));
  NOi21      u42(.An(men_men_n34_), .B(men_men_n30_), .Y(men07));
  INV        u43(.A(i_3_), .Y(men08));
  INV        u44(.A(men_men_n27_), .Y(men_men_n62_));
  NA2        u45(.A(men07), .B(men_men_n62_), .Y(men_men_n63_));
  XO2        u46(.A(men_men_n63_), .B(men_men_n26_), .Y(men05));
  NO2        u47(.A(i_2_), .B(men08), .Y(men_men_n65_));
  XO2        u48(.A(men_men_n65_), .B(i_1_), .Y(men06));
  NA2        u49(.A(men_men_n46_), .B(i_0_), .Y(men_men_n67_));
  NO2        u50(.A(i_1_), .B(i_6_), .Y(men_men_n68_));
  NO3        u51(.A(men_men_n68_), .B(men_men_n40_), .C(men_men_n34_), .Y(men_men_n69_));
  NO2        u52(.A(men_men_n69_), .B(men_men_n36_), .Y(men_men_n70_));
  OR2        u53(.A(men_men_n39_), .B(men_men_n18_), .Y(men_men_n71_));
  NO2        u54(.A(men_men_n27_), .B(men_men_n26_), .Y(men_men_n72_));
  NO2        u55(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n73_));
  OAI210     u56(.A0(men_men_n22_), .A1(i_6_), .B0(men_men_n18_), .Y(men_men_n74_));
  NO2        u57(.A(men_men_n74_), .B(men_men_n45_), .Y(men_men_n75_));
  AOI210     u58(.A0(men_men_n73_), .A1(men_men_n72_), .B0(men_men_n75_), .Y(men_men_n76_));
  NA4        u59(.A(men_men_n76_), .B(men_men_n71_), .C(men_men_n70_), .D(men_men_n67_), .Y(men03));
  NA2        u60(.A(men_men_n26_), .B(men08), .Y(men_men_n78_));
  OAI210     u61(.A0(men_men_n78_), .A1(i_1_), .B0(men_men_n55_), .Y(men_men_n79_));
  OAI210     u62(.A0(men_men_n79_), .A1(men_men_n31_), .B0(i_6_), .Y(men_men_n80_));
  AOI210     u63(.A0(men_men_n30_), .A1(men_men_n24_), .B0(men_men_n27_), .Y(men_men_n81_));
  OR2        u64(.A(men_men_n81_), .B(men_men_n68_), .Y(men_men_n82_));
  NA3        u65(.A(men_men_n78_), .B(men_men_n68_), .C(i_2_), .Y(men_men_n83_));
  NA3        u66(.A(men_men_n23_), .B(i_1_), .C(men_men_n24_), .Y(men_men_n84_));
  NA4        u67(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n82_), .D(men_men_n80_), .Y(men04));
  INV        u68(.A(men_men_n44_), .Y(men_men_n88_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
endmodule