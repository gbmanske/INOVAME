library verilog;
use verilog.vl_types.all;
entity testeflecha_vlg_check_tst is
    port(
        q1              : in     vl_logic;
        q2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end testeflecha_vlg_check_tst;
