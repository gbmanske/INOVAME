//Benchmark atmr_5xp1_76_0.5

module atmr_5xp1(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n51_, ori_ori_n52_, ori_ori_n54_, ori_ori_n56_, ori_ori_n57_, ori_ori_n59_, ori_ori_n60_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n51_, mai_mai_n55_, mai_mai_n56_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n63_, men_men_n67_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n88_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09;
  INV        o00(.A(i_5_), .Y(ori_ori_n18_));
  NO3        o01(.A(i_4_), .B(i_6_), .C(ori_ori_n18_), .Y(ori_ori_n19_));
  INV        o02(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o03(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n21_));
  INV        o04(.A(i_1_), .Y(ori_ori_n22_));
  AOI210     o05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(ori_ori_n23_));
  INV        o06(.A(i_6_), .Y(ori_ori_n24_));
  NO2        o07(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n25_));
  INV        o08(.A(i_0_), .Y(ori_ori_n26_));
  NO2        o09(.A(i_2_), .B(i_1_), .Y(ori_ori_n27_));
  NO2        o10(.A(ori_ori_n20_), .B(i_5_), .Y(ori_ori_n28_));
  NO2        o11(.A(i_2_), .B(i_3_), .Y(ori_ori_n29_));
  NO3        o12(.A(ori_ori_n29_), .B(ori_ori_n26_), .C(ori_ori_n22_), .Y(ori_ori_n30_));
  NA2        o13(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n31_));
  NA2        o14(.A(i_2_), .B(i_3_), .Y(ori_ori_n32_));
  NO2        o15(.A(ori_ori_n31_), .B(i_0_), .Y(ori_ori_n33_));
  OR3        o16(.A(ori_ori_n33_), .B(ori_ori_n25_), .C(ori_ori_n19_), .Y(ori01));
  NA2        o17(.A(i_0_), .B(i_1_), .Y(ori_ori_n35_));
  NO2        o18(.A(ori_ori_n35_), .B(i_6_), .Y(ori_ori_n36_));
  NO2        o19(.A(ori_ori_n31_), .B(ori_ori_n26_), .Y(ori_ori_n37_));
  NO3        o20(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(i_4_), .Y(ori_ori_n38_));
  NO2        o21(.A(i_6_), .B(ori_ori_n20_), .Y(ori_ori_n39_));
  NA2        o22(.A(ori_ori_n26_), .B(ori_ori_n24_), .Y(ori_ori_n40_));
  NO2        o23(.A(ori_ori_n40_), .B(ori_ori_n20_), .Y(ori_ori_n41_));
  INV        o24(.A(ori_ori_n41_), .Y(ori_ori_n42_));
  OAI210     o25(.A0(ori_ori_n39_), .A1(ori_ori_n38_), .B0(ori_ori_n42_), .Y(ori02));
  NAi21      o26(.An(ori_ori_n21_), .B(i_6_), .Y(ori_ori_n44_));
  NO2        o27(.A(ori_ori_n41_), .B(ori_ori_n28_), .Y(ori_ori_n45_));
  NA2        o28(.A(ori_ori_n45_), .B(ori_ori_n44_), .Y(ori00));
  NA2        o29(.A(ori_ori_n40_), .B(i_5_), .Y(ori_ori_n47_));
  NO2        o30(.A(ori_ori_n47_), .B(ori_ori_n20_), .Y(ori09));
  NOi21      o31(.An(ori_ori_n32_), .B(ori_ori_n29_), .Y(ori07));
  INV        o32(.A(i_3_), .Y(ori08));
  INV        o33(.A(ori_ori_n27_), .Y(ori_ori_n51_));
  NA2        o34(.A(ori07), .B(ori_ori_n51_), .Y(ori_ori_n52_));
  XO2        o35(.A(ori_ori_n52_), .B(ori_ori_n26_), .Y(ori05));
  NO2        o36(.A(i_2_), .B(ori08), .Y(ori_ori_n54_));
  XO2        o37(.A(ori_ori_n54_), .B(i_1_), .Y(ori06));
  INV        o38(.A(ori_ori_n33_), .Y(ori_ori_n56_));
  OR2        o39(.A(ori_ori_n35_), .B(ori_ori_n18_), .Y(ori_ori_n57_));
  NA2        o40(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori03));
  NA2        o41(.A(ori_ori_n30_), .B(i_6_), .Y(ori_ori_n59_));
  NA3        o42(.A(ori_ori_n23_), .B(i_1_), .C(ori_ori_n24_), .Y(ori_ori_n60_));
  NA2        o43(.A(ori_ori_n60_), .B(ori_ori_n59_), .Y(ori04));
  INV        m00(.A(i_5_), .Y(mai_mai_n18_));
  NO3        m01(.A(i_4_), .B(i_6_), .C(mai_mai_n18_), .Y(mai_mai_n19_));
  INV        m02(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m03(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n21_));
  INV        m04(.A(i_1_), .Y(mai_mai_n22_));
  AOI210     m05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(mai_mai_n23_));
  NA2        m06(.A(mai_mai_n23_), .B(mai_mai_n22_), .Y(mai_mai_n24_));
  NO2        m07(.A(mai_mai_n24_), .B(mai_mai_n21_), .Y(mai_mai_n25_));
  INV        m08(.A(i_6_), .Y(mai_mai_n26_));
  INV        m09(.A(i_0_), .Y(mai_mai_n27_));
  NO2        m10(.A(i_2_), .B(i_1_), .Y(mai_mai_n28_));
  NO2        m11(.A(mai_mai_n20_), .B(i_5_), .Y(mai_mai_n29_));
  NO2        m12(.A(i_2_), .B(i_3_), .Y(mai_mai_n30_));
  NO3        m13(.A(mai_mai_n30_), .B(mai_mai_n27_), .C(mai_mai_n22_), .Y(mai_mai_n31_));
  NA2        m14(.A(i_2_), .B(i_3_), .Y(mai_mai_n32_));
  OR3        m15(.A(mai_mai_n29_), .B(mai_mai_n25_), .C(mai_mai_n19_), .Y(mai01));
  AOI210     m16(.A0(mai_mai_n23_), .A1(mai_mai_n22_), .B0(mai_mai_n26_), .Y(mai_mai_n34_));
  AOI210     m17(.A0(mai_mai_n34_), .A1(i_5_), .B0(mai_mai_n26_), .Y(mai_mai_n35_));
  NO2        m18(.A(i_5_), .B(mai_mai_n26_), .Y(mai_mai_n36_));
  NO3        m19(.A(mai_mai_n36_), .B(mai_mai_n35_), .C(i_4_), .Y(mai_mai_n37_));
  NA2        m20(.A(i_0_), .B(i_6_), .Y(mai_mai_n38_));
  OAI210     m21(.A0(i_0_), .A1(i_1_), .B0(mai_mai_n38_), .Y(mai_mai_n39_));
  NO2        m22(.A(mai_mai_n38_), .B(mai_mai_n28_), .Y(mai_mai_n40_));
  NO2        m23(.A(i_6_), .B(i_5_), .Y(mai_mai_n41_));
  NO3        m24(.A(mai_mai_n41_), .B(mai_mai_n40_), .C(mai_mai_n20_), .Y(mai_mai_n42_));
  AOI210     m25(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(mai_mai_n43_));
  AO210      m26(.A0(mai_mai_n43_), .A1(mai_mai_n29_), .B0(mai_mai_n19_), .Y(mai_mai_n44_));
  INV        m27(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  OAI210     m28(.A0(mai_mai_n42_), .A1(mai_mai_n37_), .B0(mai_mai_n45_), .Y(mai02));
  NAi21      m29(.An(mai_mai_n21_), .B(mai_mai_n34_), .Y(mai_mai_n47_));
  NA3        m30(.A(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n48_));
  INV        m31(.A(mai_mai_n29_), .Y(mai_mai_n49_));
  NA2        m32(.A(mai_mai_n49_), .B(mai_mai_n47_), .Y(mai00));
  INV        m33(.A(i_5_), .Y(mai_mai_n51_));
  NO2        m34(.A(mai_mai_n51_), .B(mai_mai_n20_), .Y(mai09));
  NOi21      m35(.An(mai_mai_n32_), .B(mai_mai_n30_), .Y(mai07));
  INV        m36(.A(i_3_), .Y(mai08));
  INV        m37(.A(mai_mai_n28_), .Y(mai_mai_n55_));
  NA2        m38(.A(mai07), .B(mai_mai_n55_), .Y(mai_mai_n56_));
  XO2        m39(.A(mai_mai_n56_), .B(mai_mai_n27_), .Y(mai05));
  NO2        m40(.A(i_2_), .B(mai08), .Y(mai_mai_n58_));
  XO2        m41(.A(mai_mai_n58_), .B(i_1_), .Y(mai06));
  NA2        m42(.A(mai_mai_n18_), .B(i_0_), .Y(mai_mai_n60_));
  NO2        m43(.A(i_1_), .B(i_6_), .Y(mai_mai_n61_));
  NO3        m44(.A(mai_mai_n61_), .B(i_5_), .C(mai_mai_n32_), .Y(mai_mai_n62_));
  INV        m45(.A(mai_mai_n62_), .Y(mai_mai_n63_));
  OR2        m46(.A(mai_mai_n24_), .B(mai_mai_n18_), .Y(mai_mai_n64_));
  NO2        m47(.A(i_5_), .B(mai_mai_n39_), .Y(mai_mai_n65_));
  AOI210     m48(.A0(i_6_), .A1(i_0_), .B0(mai_mai_n65_), .Y(mai_mai_n66_));
  NA4        m49(.A(mai_mai_n66_), .B(mai_mai_n64_), .C(mai_mai_n63_), .D(mai_mai_n60_), .Y(mai03));
  NA2        m50(.A(mai_mai_n27_), .B(mai08), .Y(mai_mai_n68_));
  OAI210     m51(.A0(mai_mai_n68_), .A1(i_1_), .B0(mai_mai_n48_), .Y(mai_mai_n69_));
  OAI210     m52(.A0(mai_mai_n69_), .A1(mai_mai_n31_), .B0(i_6_), .Y(mai_mai_n70_));
  AOI210     m53(.A0(mai_mai_n30_), .A1(mai_mai_n26_), .B0(mai_mai_n28_), .Y(mai_mai_n71_));
  OR2        m54(.A(mai_mai_n71_), .B(mai_mai_n61_), .Y(mai_mai_n72_));
  NA3        m55(.A(mai_mai_n68_), .B(mai_mai_n61_), .C(i_2_), .Y(mai_mai_n73_));
  NA3        m56(.A(mai_mai_n73_), .B(mai_mai_n72_), .C(mai_mai_n70_), .Y(mai04));
  INV        u00(.A(i_5_), .Y(men_men_n18_));
  NO3        u01(.A(i_4_), .B(i_6_), .C(men_men_n18_), .Y(men_men_n19_));
  INV        u02(.A(i_4_), .Y(men_men_n20_));
  INV        u03(.A(i_5_), .Y(men_men_n21_));
  INV        u04(.A(i_1_), .Y(men_men_n22_));
  AOI210     u05(.A0(i_2_), .A1(i_3_), .B0(i_0_), .Y(men_men_n23_));
  NA2        u06(.A(men_men_n23_), .B(men_men_n22_), .Y(men_men_n24_));
  NO2        u07(.A(men_men_n24_), .B(men_men_n21_), .Y(men_men_n25_));
  INV        u08(.A(i_6_), .Y(men_men_n26_));
  NO2        u09(.A(men_men_n26_), .B(i_5_), .Y(men_men_n27_));
  INV        u10(.A(i_0_), .Y(men_men_n28_));
  NO2        u11(.A(i_2_), .B(i_1_), .Y(men_men_n29_));
  OAI210     u12(.A0(men_men_n29_), .A1(men_men_n28_), .B0(men_men_n20_), .Y(men_men_n30_));
  NO2        u13(.A(men_men_n20_), .B(i_5_), .Y(men_men_n31_));
  NO2        u14(.A(i_2_), .B(i_3_), .Y(men_men_n32_));
  NO3        u15(.A(men_men_n32_), .B(men_men_n28_), .C(men_men_n22_), .Y(men_men_n33_));
  AO220      u16(.A0(men_men_n33_), .A1(men_men_n31_), .B0(men_men_n30_), .B1(men_men_n27_), .Y(men_men_n34_));
  NA2        u17(.A(i_2_), .B(i_3_), .Y(men_men_n35_));
  NO2        u18(.A(men_men_n35_), .B(men_men_n22_), .Y(men_men_n36_));
  NO3        u19(.A(men_men_n36_), .B(men_men_n88_), .C(i_0_), .Y(men_men_n37_));
  OR4        u20(.A(men_men_n37_), .B(men_men_n34_), .C(men_men_n25_), .D(men_men_n19_), .Y(men01));
  OR2        u21(.A(i_2_), .B(i_3_), .Y(men_men_n39_));
  NA3        u22(.A(men_men_n39_), .B(i_0_), .C(i_1_), .Y(men_men_n40_));
  NA2        u23(.A(men_men_n28_), .B(men_men_n18_), .Y(men_men_n41_));
  AOI210     u24(.A0(men_men_n23_), .A1(men_men_n22_), .B0(men_men_n26_), .Y(men_men_n42_));
  AOI220     u25(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n40_), .B1(men_men_n26_), .Y(men_men_n43_));
  NA2        u26(.A(men_men_n29_), .B(men_men_n18_), .Y(men_men_n44_));
  NO2        u27(.A(men_men_n44_), .B(men_men_n26_), .Y(men_men_n45_));
  NO3        u28(.A(men_men_n45_), .B(men_men_n43_), .C(i_4_), .Y(men_men_n46_));
  NA2        u29(.A(i_0_), .B(i_6_), .Y(men_men_n47_));
  OAI210     u30(.A0(i_0_), .A1(i_1_), .B0(men_men_n47_), .Y(men_men_n48_));
  NOi31      u31(.An(men_men_n48_), .B(men_men_n23_), .C(men_men_n18_), .Y(men_men_n49_));
  NA3        u32(.A(i_1_), .B(i_6_), .C(i_5_), .Y(men_men_n50_));
  AOI210     u33(.A0(men_men_n50_), .A1(men_men_n47_), .B0(men_men_n29_), .Y(men_men_n51_));
  NO3        u34(.A(men_men_n39_), .B(i_6_), .C(i_5_), .Y(men_men_n52_));
  NO4        u35(.A(men_men_n52_), .B(men_men_n51_), .C(men_men_n49_), .D(men_men_n20_), .Y(men_men_n53_));
  NA2        u36(.A(men_men_n28_), .B(men_men_n26_), .Y(men_men_n54_));
  NO2        u37(.A(men_men_n54_), .B(men_men_n20_), .Y(men_men_n55_));
  AOI210     u38(.A0(i_0_), .A1(i_1_), .B0(i_6_), .Y(men_men_n56_));
  AO220      u39(.A0(men_men_n56_), .A1(men_men_n31_), .B0(men_men_n36_), .B1(men_men_n19_), .Y(men_men_n57_));
  AOI210     u40(.A0(men_men_n55_), .A1(men_men_n35_), .B0(men_men_n57_), .Y(men_men_n58_));
  OAI210     u41(.A0(men_men_n53_), .A1(men_men_n46_), .B0(men_men_n58_), .Y(men02));
  NA3        u42(.A(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n60_));
  AOI210     u43(.A0(men_men_n55_), .A1(men_men_n60_), .B0(men_men_n31_), .Y(men_men_n61_));
  INV        u44(.A(men_men_n61_), .Y(men00));
  OAI210     u45(.A0(men_men_n54_), .A1(men_men_n36_), .B0(i_5_), .Y(men_men_n63_));
  NO2        u46(.A(men_men_n63_), .B(men_men_n20_), .Y(men09));
  NOi21      u47(.An(men_men_n35_), .B(men_men_n32_), .Y(men07));
  INV        u48(.A(i_3_), .Y(men08));
  INV        u49(.A(men07), .Y(men_men_n67_));
  XO2        u50(.A(men_men_n67_), .B(men_men_n28_), .Y(men05));
  NAi21      u51(.An(men_men_n52_), .B(men_men_n44_), .Y(men_men_n69_));
  NA2        u52(.A(men_men_n69_), .B(i_0_), .Y(men_men_n70_));
  NO2        u53(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u54(.A(men_men_n41_), .B(men_men_n35_), .Y(men_men_n72_));
  NO2        u55(.A(men_men_n72_), .B(men_men_n37_), .Y(men_men_n73_));
  AO210      u56(.A0(men_men_n40_), .A1(men_men_n24_), .B0(men_men_n18_), .Y(men_men_n74_));
  NO2        u57(.A(men_men_n26_), .B(men_men_n18_), .Y(men_men_n75_));
  OAI210     u58(.A0(men_men_n22_), .A1(i_6_), .B0(men_men_n18_), .Y(men_men_n76_));
  NO2        u59(.A(men_men_n76_), .B(men_men_n48_), .Y(men_men_n77_));
  AOI210     u60(.A0(men_men_n75_), .A1(i_2_), .B0(men_men_n77_), .Y(men_men_n78_));
  NA4        u61(.A(men_men_n78_), .B(men_men_n74_), .C(men_men_n73_), .D(men_men_n70_), .Y(men03));
  NA2        u62(.A(men_men_n28_), .B(men08), .Y(men_men_n80_));
  OAI210     u63(.A0(men_men_n28_), .A1(men_men_n33_), .B0(i_6_), .Y(men_men_n81_));
  OR2        u64(.A(i_2_), .B(men_men_n71_), .Y(men_men_n82_));
  NA3        u65(.A(men_men_n80_), .B(men_men_n71_), .C(i_2_), .Y(men_men_n83_));
  NA3        u66(.A(men_men_n23_), .B(i_1_), .C(men_men_n26_), .Y(men_men_n84_));
  NA4        u67(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n82_), .D(men_men_n81_), .Y(men04));
  INV        u68(.A(i_5_), .Y(men_men_n88_));
  BUFFER     u69(.A(i_1_), .Y(men06));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
endmodule