// Benchmark "top" written by ABC on Thu Jun 20 14:00:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output zz01, zz02, zz00, zz07, zz05, zz06, zz03, zz04;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n136_, new_new_n137_, new_new_n138_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1044_, new_new_n1045_, new_new_n1046_, new_new_n1047_,
    new_new_n1048_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g0020(.A(new_new_n35_), .Y(zz01));
  INV        g0021(.A(i_11_), .Y(new_new_n44_));
  NO2        g0022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g0023(.A(i_2_), .Y(new_new_n46_));
  NA2        g0024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g0025(.A(i_5_), .Y(new_new_n48_));
  NO2        g0026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g0027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g0028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g0029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g0030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g0031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NA2        g0032(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n55_));
  NA3        g0033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g0034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g0035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  OAI210     g0036(.A0(new_new_n58_), .A1(new_new_n57_), .B0(new_new_n56_), .Y(new_new_n59_));
  NA2        g0037(.A(new_new_n59_), .B(i_12_), .Y(new_new_n60_));
  NAi21      g0038(.An(i_2_), .B(i_7_), .Y(new_new_n61_));
  INV        g0039(.A(i_1_), .Y(new_new_n62_));
  NA2        g0040(.A(new_new_n62_), .B(i_6_), .Y(new_new_n63_));
  NA3        g0041(.A(new_new_n63_), .B(new_new_n61_), .C(new_new_n31_), .Y(new_new_n64_));
  NA2        g0042(.A(i_1_), .B(i_10_), .Y(new_new_n65_));
  NO2        g0043(.A(new_new_n65_), .B(i_6_), .Y(new_new_n66_));
  NAi31      g0044(.An(new_new_n66_), .B(new_new_n64_), .C(new_new_n60_), .Y(new_new_n67_));
  NA2        g0045(.A(new_new_n50_), .B(i_2_), .Y(new_new_n68_));
  AOI210     g0046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n69_));
  NA2        g0047(.A(i_1_), .B(i_6_), .Y(new_new_n70_));
  NO2        g0048(.A(new_new_n70_), .B(new_new_n25_), .Y(new_new_n71_));
  INV        g0049(.A(i_0_), .Y(new_new_n72_));
  NAi21      g0050(.An(i_5_), .B(i_10_), .Y(new_new_n73_));
  NA2        g0051(.A(i_5_), .B(i_9_), .Y(new_new_n74_));
  AOI210     g0052(.A0(new_new_n74_), .A1(new_new_n73_), .B0(new_new_n72_), .Y(new_new_n75_));
  NO2        g0053(.A(new_new_n75_), .B(new_new_n71_), .Y(new_new_n76_));
  OAI210     g0054(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n76_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n77_), .A1(new_new_n67_), .B0(i_0_), .Y(new_new_n78_));
  NA2        g0056(.A(i_12_), .B(i_5_), .Y(new_new_n79_));
  NA2        g0057(.A(i_2_), .B(i_8_), .Y(new_new_n80_));
  NO2        g0058(.A(i_3_), .B(i_9_), .Y(new_new_n81_));
  NO2        g0059(.A(i_3_), .B(i_7_), .Y(new_new_n82_));
  INV        g0060(.A(i_6_), .Y(new_new_n83_));
  OR4        g0061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n84_));
  INV        g0062(.A(new_new_n84_), .Y(new_new_n85_));
  NO2        g0063(.A(i_2_), .B(i_7_), .Y(new_new_n86_));
  NAi21      g0064(.An(i_6_), .B(i_10_), .Y(new_new_n87_));
  NA2        g0065(.A(i_6_), .B(i_9_), .Y(new_new_n88_));
  AOI210     g0066(.A0(new_new_n88_), .A1(new_new_n87_), .B0(new_new_n62_), .Y(new_new_n89_));
  NA2        g0067(.A(i_2_), .B(i_6_), .Y(new_new_n90_));
  INV        g0068(.A(new_new_n89_), .Y(new_new_n91_));
  NO2        g0069(.A(new_new_n91_), .B(new_new_n79_), .Y(new_new_n92_));
  AN3        g0070(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n93_));
  NAi21      g0071(.An(i_6_), .B(i_11_), .Y(new_new_n94_));
  NO2        g0072(.A(i_5_), .B(i_8_), .Y(new_new_n95_));
  NOi21      g0073(.An(new_new_n95_), .B(new_new_n94_), .Y(new_new_n96_));
  AOI220     g0074(.A0(new_new_n96_), .A1(new_new_n61_), .B0(new_new_n93_), .B1(new_new_n32_), .Y(new_new_n97_));
  INV        g0075(.A(i_7_), .Y(new_new_n98_));
  NA2        g0076(.A(new_new_n46_), .B(new_new_n98_), .Y(new_new_n99_));
  NO2        g0077(.A(i_0_), .B(i_5_), .Y(new_new_n100_));
  NO2        g0078(.A(new_new_n100_), .B(new_new_n83_), .Y(new_new_n101_));
  NA2        g0079(.A(i_12_), .B(i_3_), .Y(new_new_n102_));
  INV        g0080(.A(new_new_n102_), .Y(new_new_n103_));
  NA3        g0081(.A(new_new_n103_), .B(new_new_n101_), .C(new_new_n99_), .Y(new_new_n104_));
  NAi21      g0082(.An(i_7_), .B(i_11_), .Y(new_new_n105_));
  NO3        g0083(.A(new_new_n105_), .B(new_new_n87_), .C(new_new_n53_), .Y(new_new_n106_));
  AN2        g0084(.A(i_2_), .B(i_10_), .Y(new_new_n107_));
  NO2        g0085(.A(new_new_n107_), .B(i_7_), .Y(new_new_n108_));
  OR2        g0086(.A(new_new_n79_), .B(new_new_n57_), .Y(new_new_n109_));
  NO2        g0087(.A(i_8_), .B(new_new_n98_), .Y(new_new_n110_));
  NO3        g0088(.A(new_new_n110_), .B(new_new_n109_), .C(new_new_n108_), .Y(new_new_n111_));
  NA2        g0089(.A(i_12_), .B(i_7_), .Y(new_new_n112_));
  NO2        g0090(.A(new_new_n62_), .B(new_new_n26_), .Y(new_new_n113_));
  NA2        g0091(.A(new_new_n113_), .B(i_0_), .Y(new_new_n114_));
  NA2        g0092(.A(i_11_), .B(i_12_), .Y(new_new_n115_));
  OAI210     g0093(.A0(new_new_n114_), .A1(new_new_n112_), .B0(new_new_n115_), .Y(new_new_n116_));
  NO2        g0094(.A(new_new_n116_), .B(new_new_n111_), .Y(new_new_n117_));
  NAi41      g0095(.An(new_new_n106_), .B(new_new_n117_), .C(new_new_n104_), .D(new_new_n97_), .Y(new_new_n118_));
  NOi21      g0096(.An(i_1_), .B(i_5_), .Y(new_new_n119_));
  NA2        g0097(.A(new_new_n119_), .B(i_11_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n98_), .B(new_new_n37_), .Y(new_new_n121_));
  NA2        g0099(.A(i_7_), .B(new_new_n25_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n122_), .B(new_new_n121_), .Y(new_new_n123_));
  NO2        g0101(.A(new_new_n123_), .B(new_new_n46_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n88_), .B(new_new_n87_), .Y(new_new_n125_));
  NAi21      g0103(.An(i_3_), .B(i_8_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(new_new_n61_), .Y(new_new_n127_));
  NOi31      g0105(.An(new_new_n127_), .B(new_new_n125_), .C(new_new_n124_), .Y(new_new_n128_));
  NO2        g0106(.A(i_1_), .B(new_new_n83_), .Y(new_new_n129_));
  NO2        g0107(.A(i_6_), .B(i_5_), .Y(new_new_n130_));
  NA2        g0108(.A(new_new_n130_), .B(i_3_), .Y(new_new_n131_));
  AO210      g0109(.A0(new_new_n131_), .A1(new_new_n47_), .B0(new_new_n129_), .Y(new_new_n132_));
  OAI220     g0110(.A0(new_new_n132_), .A1(new_new_n105_), .B0(new_new_n128_), .B1(new_new_n120_), .Y(new_new_n133_));
  NO3        g0111(.A(new_new_n133_), .B(new_new_n118_), .C(new_new_n92_), .Y(new_new_n134_));
  NA3        g0112(.A(new_new_n134_), .B(new_new_n78_), .C(new_new_n55_), .Y(zz02));
  NO2        g0113(.A(new_new_n62_), .B(new_new_n37_), .Y(new_new_n136_));
  NA2        g0114(.A(i_6_), .B(new_new_n25_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(new_new_n136_), .Y(new_new_n138_));
  NA4        g0116(.A(new_new_n138_), .B(new_new_n76_), .C(new_new_n68_), .D(new_new_n30_), .Y(zz00));
  AN2        g0117(.A(i_8_), .B(i_7_), .Y(new_new_n140_));
  NA2        g0118(.A(new_new_n140_), .B(i_6_), .Y(new_new_n141_));
  NO2        g0119(.A(i_12_), .B(i_13_), .Y(new_new_n142_));
  NAi21      g0120(.An(i_5_), .B(i_11_), .Y(new_new_n143_));
  NOi21      g0121(.An(new_new_n142_), .B(new_new_n143_), .Y(new_new_n144_));
  NO2        g0122(.A(i_0_), .B(i_1_), .Y(new_new_n145_));
  NA2        g0123(.A(i_2_), .B(i_3_), .Y(new_new_n146_));
  NO2        g0124(.A(new_new_n146_), .B(i_4_), .Y(new_new_n147_));
  NA3        g0125(.A(new_new_n147_), .B(new_new_n145_), .C(new_new_n144_), .Y(new_new_n148_));
  AN2        g0126(.A(new_new_n142_), .B(new_new_n81_), .Y(new_new_n149_));
  NO2        g0127(.A(new_new_n149_), .B(new_new_n27_), .Y(new_new_n150_));
  NA2        g0128(.A(i_1_), .B(i_5_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n72_), .B(new_new_n46_), .Y(new_new_n152_));
  NA2        g0130(.A(new_new_n152_), .B(new_new_n36_), .Y(new_new_n153_));
  NO3        g0131(.A(new_new_n153_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n154_));
  OR2        g0132(.A(i_0_), .B(i_1_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n79_), .C(i_13_), .Y(new_new_n156_));
  NAi32      g0134(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n157_));
  NAi21      g0135(.An(new_new_n157_), .B(new_new_n156_), .Y(new_new_n158_));
  NOi21      g0136(.An(i_4_), .B(i_10_), .Y(new_new_n159_));
  NA2        g0137(.A(new_new_n159_), .B(new_new_n40_), .Y(new_new_n160_));
  NO2        g0138(.A(i_3_), .B(i_5_), .Y(new_new_n161_));
  NO3        g0139(.A(new_new_n72_), .B(i_2_), .C(i_1_), .Y(new_new_n162_));
  NA2        g0140(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  OAI210     g0141(.A0(new_new_n163_), .A1(new_new_n160_), .B0(new_new_n158_), .Y(new_new_n164_));
  NO2        g0142(.A(new_new_n164_), .B(new_new_n154_), .Y(new_new_n165_));
  AOI210     g0143(.A0(new_new_n165_), .A1(new_new_n148_), .B0(new_new_n141_), .Y(new_new_n166_));
  NA2        g0144(.A(i_3_), .B(new_new_n48_), .Y(new_new_n167_));
  NOi21      g0145(.An(i_4_), .B(i_9_), .Y(new_new_n168_));
  NOi21      g0146(.An(i_11_), .B(i_13_), .Y(new_new_n169_));
  NA2        g0147(.A(new_new_n169_), .B(new_new_n168_), .Y(new_new_n170_));
  OR2        g0148(.A(new_new_n170_), .B(new_new_n167_), .Y(new_new_n171_));
  NO2        g0149(.A(i_4_), .B(i_5_), .Y(new_new_n172_));
  NAi21      g0150(.An(i_12_), .B(i_11_), .Y(new_new_n173_));
  NO2        g0151(.A(new_new_n173_), .B(i_13_), .Y(new_new_n174_));
  NA3        g0152(.A(new_new_n174_), .B(new_new_n172_), .C(new_new_n81_), .Y(new_new_n175_));
  AOI210     g0153(.A0(new_new_n175_), .A1(new_new_n171_), .B0(new_new_n1046_), .Y(new_new_n176_));
  NO2        g0154(.A(new_new_n72_), .B(new_new_n62_), .Y(new_new_n177_));
  NA2        g0155(.A(new_new_n177_), .B(new_new_n46_), .Y(new_new_n178_));
  NA2        g0156(.A(new_new_n36_), .B(i_5_), .Y(new_new_n179_));
  NAi31      g0157(.An(new_new_n179_), .B(new_new_n149_), .C(i_11_), .Y(new_new_n180_));
  NA2        g0158(.A(i_3_), .B(i_5_), .Y(new_new_n181_));
  OR2        g0159(.A(new_new_n181_), .B(new_new_n170_), .Y(new_new_n182_));
  AOI210     g0160(.A0(new_new_n182_), .A1(new_new_n180_), .B0(new_new_n178_), .Y(new_new_n183_));
  NO2        g0161(.A(new_new_n72_), .B(i_5_), .Y(new_new_n184_));
  NO2        g0162(.A(i_13_), .B(i_10_), .Y(new_new_n185_));
  NA3        g0163(.A(new_new_n185_), .B(new_new_n184_), .C(new_new_n44_), .Y(new_new_n186_));
  NO2        g0164(.A(i_2_), .B(i_1_), .Y(new_new_n187_));
  NA2        g0165(.A(new_new_n187_), .B(i_3_), .Y(new_new_n188_));
  NAi21      g0166(.An(i_4_), .B(i_12_), .Y(new_new_n189_));
  NO4        g0167(.A(new_new_n189_), .B(new_new_n188_), .C(new_new_n186_), .D(new_new_n25_), .Y(new_new_n190_));
  NO3        g0168(.A(new_new_n190_), .B(new_new_n183_), .C(new_new_n176_), .Y(new_new_n191_));
  INV        g0169(.A(i_8_), .Y(new_new_n192_));
  NO2        g0170(.A(new_new_n192_), .B(i_7_), .Y(new_new_n193_));
  NA2        g0171(.A(new_new_n193_), .B(i_6_), .Y(new_new_n194_));
  NO3        g0172(.A(i_3_), .B(new_new_n83_), .C(new_new_n48_), .Y(new_new_n195_));
  NA2        g0173(.A(new_new_n195_), .B(new_new_n110_), .Y(new_new_n196_));
  NO3        g0174(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n197_));
  NA3        g0175(.A(new_new_n197_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n198_));
  NO3        g0176(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n199_));
  OAI210     g0177(.A0(new_new_n93_), .A1(i_12_), .B0(new_new_n199_), .Y(new_new_n200_));
  AOI210     g0178(.A0(new_new_n200_), .A1(new_new_n198_), .B0(new_new_n196_), .Y(new_new_n201_));
  NO2        g0179(.A(i_3_), .B(i_8_), .Y(new_new_n202_));
  NO3        g0180(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n203_));
  NA3        g0181(.A(new_new_n203_), .B(new_new_n202_), .C(new_new_n40_), .Y(new_new_n204_));
  NO2        g0182(.A(i_13_), .B(i_9_), .Y(new_new_n205_));
  NA3        g0183(.A(new_new_n205_), .B(i_6_), .C(new_new_n192_), .Y(new_new_n206_));
  NAi21      g0184(.An(i_12_), .B(i_3_), .Y(new_new_n207_));
  NO2        g0185(.A(new_new_n44_), .B(i_5_), .Y(new_new_n208_));
  NO3        g0186(.A(i_0_), .B(i_2_), .C(new_new_n62_), .Y(new_new_n209_));
  NA3        g0187(.A(new_new_n209_), .B(new_new_n208_), .C(i_10_), .Y(new_new_n210_));
  OAI220     g0188(.A0(new_new_n210_), .A1(new_new_n206_), .B0(new_new_n57_), .B1(new_new_n204_), .Y(new_new_n211_));
  AOI210     g0189(.A0(new_new_n211_), .A1(i_7_), .B0(new_new_n201_), .Y(new_new_n212_));
  OAI220     g0190(.A0(new_new_n212_), .A1(i_4_), .B0(new_new_n194_), .B1(new_new_n191_), .Y(new_new_n213_));
  NAi21      g0191(.An(i_12_), .B(i_7_), .Y(new_new_n214_));
  NA3        g0192(.A(i_13_), .B(new_new_n192_), .C(i_10_), .Y(new_new_n215_));
  NO2        g0193(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n216_));
  NA2        g0194(.A(i_0_), .B(i_5_), .Y(new_new_n217_));
  OAI220     g0195(.A0(new_new_n83_), .A1(new_new_n188_), .B0(new_new_n178_), .B1(new_new_n131_), .Y(new_new_n218_));
  NAi31      g0196(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n219_));
  NO2        g0197(.A(new_new_n36_), .B(i_13_), .Y(new_new_n220_));
  NO2        g0198(.A(new_new_n46_), .B(new_new_n62_), .Y(new_new_n221_));
  NA3        g0199(.A(new_new_n221_), .B(i_0_), .C(new_new_n220_), .Y(new_new_n222_));
  INV        g0200(.A(i_13_), .Y(new_new_n223_));
  NO2        g0201(.A(i_12_), .B(new_new_n223_), .Y(new_new_n224_));
  NA3        g0202(.A(new_new_n224_), .B(new_new_n197_), .C(new_new_n195_), .Y(new_new_n225_));
  OAI210     g0203(.A0(new_new_n222_), .A1(new_new_n219_), .B0(new_new_n225_), .Y(new_new_n226_));
  AOI220     g0204(.A0(new_new_n226_), .A1(new_new_n140_), .B0(new_new_n218_), .B1(new_new_n216_), .Y(new_new_n227_));
  NO2        g0205(.A(i_12_), .B(new_new_n37_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n181_), .B(i_4_), .Y(new_new_n229_));
  NA2        g0207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  OR2        g0208(.A(i_8_), .B(i_7_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n231_), .B(new_new_n83_), .Y(new_new_n232_));
  NO2        g0210(.A(new_new_n53_), .B(i_1_), .Y(new_new_n233_));
  NA2        g0211(.A(new_new_n233_), .B(new_new_n232_), .Y(new_new_n234_));
  INV        g0212(.A(i_12_), .Y(new_new_n235_));
  NO3        g0213(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n236_));
  NA2        g0214(.A(i_2_), .B(i_1_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n234_), .B(new_new_n230_), .Y(new_new_n238_));
  NO3        g0216(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n239_));
  NAi21      g0217(.An(i_4_), .B(i_3_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n240_), .B(new_new_n74_), .Y(new_new_n241_));
  NO2        g0219(.A(i_0_), .B(i_6_), .Y(new_new_n242_));
  NOi41      g0220(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n243_));
  NA2        g0221(.A(new_new_n243_), .B(new_new_n242_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n237_), .B(new_new_n181_), .Y(new_new_n245_));
  NAi21      g0223(.An(new_new_n244_), .B(new_new_n245_), .Y(new_new_n246_));
  INV        g0224(.A(new_new_n246_), .Y(new_new_n247_));
  AOI220     g0225(.A0(new_new_n247_), .A1(new_new_n40_), .B0(new_new_n238_), .B1(new_new_n205_), .Y(new_new_n248_));
  NO2        g0226(.A(i_11_), .B(new_new_n223_), .Y(new_new_n249_));
  NOi21      g0227(.An(i_1_), .B(i_6_), .Y(new_new_n250_));
  NAi21      g0228(.An(i_3_), .B(i_7_), .Y(new_new_n251_));
  NO2        g0229(.A(new_new_n48_), .B(new_new_n25_), .Y(new_new_n252_));
  NO2        g0230(.A(i_12_), .B(i_3_), .Y(new_new_n253_));
  NA2        g0231(.A(new_new_n72_), .B(i_5_), .Y(new_new_n254_));
  NA3        g0232(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n255_));
  INV        g0233(.A(new_new_n141_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n235_), .B(i_13_), .Y(new_new_n257_));
  NO2        g0235(.A(new_new_n257_), .B(new_new_n74_), .Y(new_new_n258_));
  NA2        g0236(.A(new_new_n258_), .B(new_new_n256_), .Y(new_new_n259_));
  NO2        g0237(.A(new_new_n231_), .B(new_new_n37_), .Y(new_new_n260_));
  NA2        g0238(.A(i_12_), .B(i_6_), .Y(new_new_n261_));
  OR2        g0239(.A(i_13_), .B(i_9_), .Y(new_new_n262_));
  NO3        g0240(.A(new_new_n262_), .B(new_new_n261_), .C(new_new_n48_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n240_), .B(i_2_), .Y(new_new_n264_));
  NA3        g0242(.A(new_new_n264_), .B(new_new_n263_), .C(new_new_n44_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n249_), .B(i_9_), .Y(new_new_n266_));
  NA3        g0244(.A(new_new_n254_), .B(new_new_n155_), .C(new_new_n63_), .Y(new_new_n267_));
  OAI210     g0245(.A0(new_new_n267_), .A1(new_new_n266_), .B0(new_new_n265_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n152_), .B(new_new_n62_), .Y(new_new_n269_));
  NO3        g0247(.A(i_11_), .B(new_new_n223_), .C(new_new_n25_), .Y(new_new_n270_));
  NO2        g0248(.A(new_new_n251_), .B(i_8_), .Y(new_new_n271_));
  NO2        g0249(.A(i_6_), .B(new_new_n48_), .Y(new_new_n272_));
  NA3        g0250(.A(new_new_n272_), .B(new_new_n271_), .C(new_new_n270_), .Y(new_new_n273_));
  NO3        g0251(.A(new_new_n26_), .B(new_new_n83_), .C(i_5_), .Y(new_new_n274_));
  NA3        g0252(.A(new_new_n274_), .B(new_new_n260_), .C(new_new_n224_), .Y(new_new_n275_));
  AOI210     g0253(.A0(new_new_n275_), .A1(new_new_n273_), .B0(new_new_n269_), .Y(new_new_n276_));
  AOI210     g0254(.A0(new_new_n268_), .A1(new_new_n260_), .B0(new_new_n276_), .Y(new_new_n277_));
  NA4        g0255(.A(new_new_n277_), .B(new_new_n259_), .C(new_new_n248_), .D(new_new_n227_), .Y(new_new_n278_));
  NO3        g0256(.A(i_12_), .B(new_new_n223_), .C(new_new_n37_), .Y(new_new_n279_));
  INV        g0257(.A(new_new_n279_), .Y(new_new_n280_));
  NA2        g0258(.A(i_8_), .B(new_new_n98_), .Y(new_new_n281_));
  NO3        g0259(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n282_));
  AOI220     g0260(.A0(new_new_n282_), .A1(new_new_n195_), .B0(new_new_n161_), .B1(new_new_n233_), .Y(new_new_n283_));
  NO2        g0261(.A(new_new_n283_), .B(new_new_n281_), .Y(new_new_n284_));
  NO2        g0262(.A(new_new_n237_), .B(i_0_), .Y(new_new_n285_));
  AOI220     g0263(.A0(new_new_n285_), .A1(new_new_n193_), .B0(i_1_), .B1(new_new_n140_), .Y(new_new_n286_));
  NA2        g0264(.A(new_new_n272_), .B(new_new_n26_), .Y(new_new_n287_));
  NO2        g0265(.A(new_new_n287_), .B(new_new_n286_), .Y(new_new_n288_));
  NA2        g0266(.A(i_0_), .B(i_1_), .Y(new_new_n289_));
  NO2        g0267(.A(new_new_n289_), .B(i_2_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n58_), .B(i_6_), .Y(new_new_n291_));
  NA3        g0269(.A(new_new_n291_), .B(new_new_n290_), .C(new_new_n161_), .Y(new_new_n292_));
  OAI210     g0270(.A0(new_new_n163_), .A1(new_new_n141_), .B0(new_new_n292_), .Y(new_new_n293_));
  NO3        g0271(.A(new_new_n293_), .B(new_new_n288_), .C(new_new_n284_), .Y(new_new_n294_));
  NO2        g0272(.A(i_3_), .B(i_10_), .Y(new_new_n295_));
  NA3        g0273(.A(new_new_n295_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n296_));
  NO2        g0274(.A(i_2_), .B(new_new_n98_), .Y(new_new_n297_));
  NA2        g0275(.A(i_1_), .B(new_new_n36_), .Y(new_new_n298_));
  NO2        g0276(.A(new_new_n298_), .B(i_8_), .Y(new_new_n299_));
  NA3        g0277(.A(new_new_n217_), .B(new_new_n299_), .C(new_new_n297_), .Y(new_new_n300_));
  AN2        g0278(.A(i_3_), .B(i_10_), .Y(new_new_n301_));
  NA4        g0279(.A(new_new_n301_), .B(new_new_n197_), .C(new_new_n174_), .D(new_new_n172_), .Y(new_new_n302_));
  NO2        g0280(.A(i_5_), .B(new_new_n37_), .Y(new_new_n303_));
  NO2        g0281(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n304_));
  OR2        g0282(.A(new_new_n300_), .B(new_new_n296_), .Y(new_new_n305_));
  OAI220     g0283(.A0(new_new_n305_), .A1(i_6_), .B0(new_new_n294_), .B1(new_new_n280_), .Y(new_new_n306_));
  NO4        g0284(.A(new_new_n306_), .B(new_new_n278_), .C(new_new_n213_), .D(new_new_n166_), .Y(new_new_n307_));
  NO3        g0285(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n308_));
  NO2        g0286(.A(new_new_n58_), .B(new_new_n83_), .Y(new_new_n309_));
  NA2        g0287(.A(new_new_n285_), .B(new_new_n309_), .Y(new_new_n310_));
  NO3        g0288(.A(i_6_), .B(new_new_n192_), .C(i_7_), .Y(new_new_n311_));
  NA2        g0289(.A(new_new_n311_), .B(new_new_n197_), .Y(new_new_n312_));
  AOI210     g0290(.A0(new_new_n312_), .A1(new_new_n310_), .B0(new_new_n167_), .Y(new_new_n313_));
  NO2        g0291(.A(i_2_), .B(i_3_), .Y(new_new_n314_));
  OR2        g0292(.A(i_0_), .B(i_5_), .Y(new_new_n315_));
  NA2        g0293(.A(new_new_n217_), .B(new_new_n315_), .Y(new_new_n316_));
  NA4        g0294(.A(new_new_n316_), .B(new_new_n232_), .C(new_new_n314_), .D(i_1_), .Y(new_new_n317_));
  NA3        g0295(.A(new_new_n285_), .B(new_new_n161_), .C(new_new_n110_), .Y(new_new_n318_));
  NAi21      g0296(.An(i_8_), .B(i_7_), .Y(new_new_n319_));
  NO2        g0297(.A(new_new_n319_), .B(i_6_), .Y(new_new_n320_));
  NO2        g0298(.A(new_new_n155_), .B(new_new_n46_), .Y(new_new_n321_));
  NA3        g0299(.A(new_new_n321_), .B(new_new_n320_), .C(new_new_n161_), .Y(new_new_n322_));
  NA3        g0300(.A(new_new_n322_), .B(new_new_n318_), .C(new_new_n317_), .Y(new_new_n323_));
  OAI210     g0301(.A0(new_new_n323_), .A1(new_new_n313_), .B0(i_4_), .Y(new_new_n324_));
  NO2        g0302(.A(i_12_), .B(i_10_), .Y(new_new_n325_));
  NOi21      g0303(.An(i_5_), .B(i_0_), .Y(new_new_n326_));
  NO3        g0304(.A(new_new_n298_), .B(new_new_n326_), .C(new_new_n126_), .Y(new_new_n327_));
  NA4        g0305(.A(new_new_n82_), .B(new_new_n36_), .C(new_new_n83_), .D(i_8_), .Y(new_new_n328_));
  NA2        g0306(.A(new_new_n327_), .B(new_new_n325_), .Y(new_new_n329_));
  NO2        g0307(.A(i_6_), .B(i_8_), .Y(new_new_n330_));
  NOi21      g0308(.An(i_0_), .B(i_2_), .Y(new_new_n331_));
  AN2        g0309(.A(new_new_n331_), .B(new_new_n330_), .Y(new_new_n332_));
  NO2        g0310(.A(i_1_), .B(i_7_), .Y(new_new_n333_));
  AO220      g0311(.A0(new_new_n333_), .A1(new_new_n332_), .B0(new_new_n320_), .B1(new_new_n233_), .Y(new_new_n334_));
  NA3        g0312(.A(new_new_n334_), .B(i_4_), .C(i_5_), .Y(new_new_n335_));
  NA3        g0313(.A(new_new_n335_), .B(new_new_n329_), .C(new_new_n324_), .Y(new_new_n336_));
  NO3        g0314(.A(new_new_n231_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n337_));
  NO3        g0315(.A(new_new_n319_), .B(i_2_), .C(i_1_), .Y(new_new_n338_));
  OAI210     g0316(.A0(new_new_n338_), .A1(new_new_n337_), .B0(i_6_), .Y(new_new_n339_));
  NA3        g0317(.A(new_new_n250_), .B(new_new_n297_), .C(new_new_n192_), .Y(new_new_n340_));
  AOI210     g0318(.A0(new_new_n340_), .A1(new_new_n339_), .B0(new_new_n316_), .Y(new_new_n341_));
  NO2        g0319(.A(new_new_n100_), .B(new_new_n122_), .Y(new_new_n342_));
  OAI210     g0320(.A0(new_new_n342_), .A1(new_new_n341_), .B0(i_3_), .Y(new_new_n343_));
  INV        g0321(.A(new_new_n82_), .Y(new_new_n344_));
  NO2        g0322(.A(new_new_n289_), .B(new_new_n80_), .Y(new_new_n345_));
  NA2        g0323(.A(new_new_n345_), .B(new_new_n130_), .Y(new_new_n346_));
  NO2        g0324(.A(new_new_n90_), .B(new_new_n192_), .Y(new_new_n347_));
  NA3        g0325(.A(new_new_n217_), .B(new_new_n347_), .C(new_new_n62_), .Y(new_new_n348_));
  AOI210     g0326(.A0(new_new_n348_), .A1(new_new_n346_), .B0(new_new_n344_), .Y(new_new_n349_));
  NO2        g0327(.A(new_new_n192_), .B(i_9_), .Y(new_new_n350_));
  NA2        g0328(.A(new_new_n350_), .B(new_new_n155_), .Y(new_new_n351_));
  NO2        g0329(.A(new_new_n351_), .B(new_new_n46_), .Y(new_new_n352_));
  NO3        g0330(.A(new_new_n352_), .B(new_new_n349_), .C(new_new_n288_), .Y(new_new_n353_));
  AOI210     g0331(.A0(new_new_n353_), .A1(new_new_n343_), .B0(new_new_n160_), .Y(new_new_n354_));
  AOI210     g0332(.A0(new_new_n336_), .A1(new_new_n308_), .B0(new_new_n354_), .Y(new_new_n355_));
  NOi32      g0333(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n356_));
  INV        g0334(.A(new_new_n356_), .Y(new_new_n357_));
  NAi21      g0335(.An(i_0_), .B(i_6_), .Y(new_new_n358_));
  NAi21      g0336(.An(i_1_), .B(i_5_), .Y(new_new_n359_));
  NA2        g0337(.A(new_new_n359_), .B(new_new_n358_), .Y(new_new_n360_));
  NA2        g0338(.A(new_new_n360_), .B(new_new_n25_), .Y(new_new_n361_));
  OAI210     g0339(.A0(new_new_n361_), .A1(new_new_n157_), .B0(new_new_n244_), .Y(new_new_n362_));
  NAi41      g0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n363_));
  OAI220     g0341(.A0(new_new_n363_), .A1(new_new_n359_), .B0(new_new_n219_), .B1(new_new_n157_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n363_), .A1(new_new_n157_), .B0(new_new_n155_), .Y(new_new_n365_));
  NOi32      g0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n366_));
  NAi21      g0344(.An(i_6_), .B(i_1_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n366_), .C(new_new_n46_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n368_), .B(i_0_), .Y(new_new_n369_));
  OR3        g0347(.A(new_new_n369_), .B(new_new_n365_), .C(new_new_n364_), .Y(new_new_n370_));
  NO2        g0348(.A(i_1_), .B(new_new_n98_), .Y(new_new_n371_));
  NAi21      g0349(.An(i_3_), .B(i_4_), .Y(new_new_n372_));
  AN2        g0350(.A(i_6_), .B(i_7_), .Y(new_new_n373_));
  NA2        g0351(.A(i_2_), .B(i_7_), .Y(new_new_n374_));
  NO2        g0352(.A(new_new_n372_), .B(i_10_), .Y(new_new_n375_));
  AOI210     g0353(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n376_));
  OAI210     g0354(.A0(new_new_n376_), .A1(new_new_n187_), .B0(new_new_n375_), .Y(new_new_n377_));
  AOI220     g0355(.A0(new_new_n375_), .A1(new_new_n333_), .B0(new_new_n236_), .B1(new_new_n187_), .Y(new_new_n378_));
  AOI210     g0356(.A0(new_new_n378_), .A1(new_new_n377_), .B0(i_5_), .Y(new_new_n379_));
  NO3        g0357(.A(new_new_n379_), .B(new_new_n370_), .C(new_new_n362_), .Y(new_new_n380_));
  NO2        g0358(.A(new_new_n380_), .B(new_new_n357_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n382_));
  AN2        g0360(.A(i_12_), .B(i_5_), .Y(new_new_n383_));
  NO2        g0361(.A(i_4_), .B(new_new_n26_), .Y(new_new_n384_));
  NA2        g0362(.A(new_new_n384_), .B(new_new_n383_), .Y(new_new_n385_));
  NO2        g0363(.A(i_11_), .B(i_6_), .Y(new_new_n386_));
  NA3        g0364(.A(new_new_n386_), .B(new_new_n321_), .C(new_new_n223_), .Y(new_new_n387_));
  NO2        g0365(.A(new_new_n387_), .B(new_new_n385_), .Y(new_new_n388_));
  NO2        g0366(.A(new_new_n240_), .B(i_5_), .Y(new_new_n389_));
  NO2        g0367(.A(i_5_), .B(i_10_), .Y(new_new_n390_));
  AOI220     g0368(.A0(new_new_n390_), .A1(new_new_n264_), .B0(new_new_n389_), .B1(new_new_n197_), .Y(new_new_n391_));
  NA2        g0369(.A(new_new_n142_), .B(new_new_n45_), .Y(new_new_n392_));
  NO2        g0370(.A(new_new_n392_), .B(new_new_n391_), .Y(new_new_n393_));
  OAI210     g0371(.A0(new_new_n393_), .A1(new_new_n388_), .B0(new_new_n382_), .Y(new_new_n394_));
  NO2        g0372(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n395_));
  NO2        g0373(.A(new_new_n148_), .B(new_new_n83_), .Y(new_new_n396_));
  OAI210     g0374(.A0(new_new_n396_), .A1(new_new_n388_), .B0(new_new_n395_), .Y(new_new_n397_));
  NO3        g0375(.A(new_new_n83_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n398_));
  NO2        g0376(.A(i_11_), .B(i_12_), .Y(new_new_n399_));
  NA2        g0377(.A(new_new_n390_), .B(new_new_n235_), .Y(new_new_n400_));
  NA3        g0378(.A(new_new_n110_), .B(i_4_), .C(i_11_), .Y(new_new_n401_));
  OAI220     g0379(.A0(new_new_n401_), .A1(new_new_n219_), .B0(new_new_n400_), .B1(new_new_n328_), .Y(new_new_n402_));
  NAi21      g0380(.An(i_13_), .B(i_0_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n237_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n402_), .B(new_new_n404_), .Y(new_new_n405_));
  NA3        g0383(.A(new_new_n405_), .B(new_new_n397_), .C(new_new_n394_), .Y(new_new_n406_));
  NO2        g0384(.A(i_0_), .B(i_11_), .Y(new_new_n407_));
  AN2        g0385(.A(i_1_), .B(i_6_), .Y(new_new_n408_));
  NOi21      g0386(.An(i_2_), .B(i_12_), .Y(new_new_n409_));
  NA2        g0387(.A(new_new_n409_), .B(new_new_n408_), .Y(new_new_n410_));
  INV        g0388(.A(new_new_n410_), .Y(new_new_n411_));
  NA2        g0389(.A(new_new_n140_), .B(i_9_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n412_), .B(i_4_), .Y(new_new_n413_));
  NA2        g0391(.A(new_new_n411_), .B(new_new_n413_), .Y(new_new_n414_));
  OR2        g0392(.A(i_13_), .B(i_10_), .Y(new_new_n415_));
  NO2        g0393(.A(new_new_n170_), .B(new_new_n121_), .Y(new_new_n416_));
  OR2        g0394(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n98_), .B(new_new_n25_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n272_), .B(new_new_n209_), .Y(new_new_n419_));
  NO2        g0397(.A(new_new_n419_), .B(new_new_n417_), .Y(new_new_n420_));
  INV        g0398(.A(new_new_n420_), .Y(new_new_n421_));
  AOI210     g0399(.A0(new_new_n421_), .A1(new_new_n414_), .B0(new_new_n26_), .Y(new_new_n422_));
  NA2        g0400(.A(new_new_n318_), .B(new_new_n317_), .Y(new_new_n423_));
  AOI220     g0401(.A0(new_new_n291_), .A1(new_new_n282_), .B0(new_new_n285_), .B1(new_new_n309_), .Y(new_new_n424_));
  NO2        g0402(.A(new_new_n424_), .B(new_new_n167_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n181_), .B(new_new_n83_), .Y(new_new_n426_));
  AOI220     g0404(.A0(new_new_n426_), .A1(new_new_n290_), .B0(new_new_n274_), .B1(new_new_n209_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(new_new_n281_), .Y(new_new_n428_));
  NO3        g0406(.A(new_new_n428_), .B(new_new_n425_), .C(new_new_n423_), .Y(new_new_n429_));
  NA2        g0407(.A(new_new_n195_), .B(new_new_n93_), .Y(new_new_n430_));
  NA3        g0408(.A(new_new_n321_), .B(new_new_n161_), .C(new_new_n83_), .Y(new_new_n431_));
  AOI210     g0409(.A0(new_new_n431_), .A1(new_new_n430_), .B0(new_new_n319_), .Y(new_new_n432_));
  NA2        g0410(.A(new_new_n291_), .B(new_new_n233_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n433_), .B(new_new_n181_), .Y(new_new_n434_));
  NO2        g0412(.A(i_3_), .B(new_new_n48_), .Y(new_new_n435_));
  NA3        g0413(.A(new_new_n333_), .B(new_new_n332_), .C(new_new_n435_), .Y(new_new_n436_));
  NA2        g0414(.A(new_new_n311_), .B(new_new_n316_), .Y(new_new_n437_));
  OAI210     g0415(.A0(new_new_n437_), .A1(new_new_n188_), .B0(new_new_n436_), .Y(new_new_n438_));
  NO3        g0416(.A(new_new_n438_), .B(new_new_n434_), .C(new_new_n432_), .Y(new_new_n439_));
  AOI210     g0417(.A0(new_new_n439_), .A1(new_new_n429_), .B0(new_new_n266_), .Y(new_new_n440_));
  NO4        g0418(.A(new_new_n440_), .B(new_new_n422_), .C(new_new_n406_), .D(new_new_n381_), .Y(new_new_n441_));
  NO2        g0419(.A(new_new_n62_), .B(i_4_), .Y(new_new_n442_));
  NO2        g0420(.A(new_new_n72_), .B(i_13_), .Y(new_new_n443_));
  NA3        g0421(.A(new_new_n443_), .B(new_new_n442_), .C(i_2_), .Y(new_new_n444_));
  NO2        g0422(.A(i_10_), .B(i_9_), .Y(new_new_n445_));
  NAi21      g0423(.An(i_12_), .B(i_8_), .Y(new_new_n446_));
  NO2        g0424(.A(new_new_n446_), .B(i_3_), .Y(new_new_n447_));
  NA2        g0425(.A(new_new_n447_), .B(new_new_n445_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n46_), .B(i_4_), .Y(new_new_n449_));
  NA2        g0427(.A(new_new_n449_), .B(new_new_n101_), .Y(new_new_n450_));
  OAI220     g0428(.A0(new_new_n450_), .A1(new_new_n204_), .B0(new_new_n448_), .B1(new_new_n444_), .Y(new_new_n451_));
  NA2        g0429(.A(new_new_n304_), .B(i_0_), .Y(new_new_n452_));
  NO3        g0430(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n453_));
  NA2        g0431(.A(new_new_n261_), .B(new_new_n94_), .Y(new_new_n454_));
  NA2        g0432(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n455_));
  NA2        g0433(.A(i_8_), .B(i_9_), .Y(new_new_n456_));
  NO2        g0434(.A(new_new_n455_), .B(new_new_n452_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n249_), .B(new_new_n303_), .Y(new_new_n458_));
  NO3        g0436(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n459_));
  AOI210     g0437(.A0(new_new_n253_), .A1(new_new_n187_), .B0(new_new_n459_), .Y(new_new_n460_));
  NA3        g0438(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n461_));
  NA4        g0439(.A(new_new_n143_), .B(new_new_n113_), .C(new_new_n79_), .D(new_new_n23_), .Y(new_new_n462_));
  OAI220     g0440(.A0(new_new_n462_), .A1(new_new_n461_), .B0(new_new_n460_), .B1(new_new_n458_), .Y(new_new_n463_));
  NO3        g0441(.A(new_new_n463_), .B(new_new_n457_), .C(new_new_n451_), .Y(new_new_n464_));
  OR2        g0442(.A(new_new_n289_), .B(new_new_n206_), .Y(new_new_n465_));
  OA210      g0443(.A0(new_new_n351_), .A1(new_new_n98_), .B0(new_new_n292_), .Y(new_new_n466_));
  OA220      g0444(.A0(new_new_n466_), .A1(new_new_n160_), .B0(new_new_n465_), .B1(new_new_n230_), .Y(new_new_n467_));
  NA2        g0445(.A(new_new_n93_), .B(i_13_), .Y(new_new_n468_));
  NA2        g0446(.A(new_new_n426_), .B(new_new_n382_), .Y(new_new_n469_));
  NO2        g0447(.A(i_2_), .B(i_13_), .Y(new_new_n470_));
  NA3        g0448(.A(new_new_n470_), .B(new_new_n159_), .C(new_new_n96_), .Y(new_new_n471_));
  OAI220     g0449(.A0(new_new_n471_), .A1(new_new_n235_), .B0(new_new_n469_), .B1(new_new_n468_), .Y(new_new_n472_));
  NO3        g0450(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n473_));
  NO2        g0451(.A(i_6_), .B(i_7_), .Y(new_new_n474_));
  NA2        g0452(.A(new_new_n474_), .B(new_new_n473_), .Y(new_new_n475_));
  NO2        g0453(.A(i_11_), .B(i_1_), .Y(new_new_n476_));
  OR2        g0454(.A(i_11_), .B(i_8_), .Y(new_new_n477_));
  NOi21      g0455(.An(i_2_), .B(i_7_), .Y(new_new_n478_));
  NAi31      g0456(.An(new_new_n477_), .B(new_new_n478_), .C(i_0_), .Y(new_new_n479_));
  NO2        g0457(.A(new_new_n415_), .B(i_6_), .Y(new_new_n480_));
  NA3        g0458(.A(new_new_n480_), .B(new_new_n442_), .C(new_new_n74_), .Y(new_new_n481_));
  NO2        g0459(.A(new_new_n481_), .B(new_new_n479_), .Y(new_new_n482_));
  NO2        g0460(.A(i_3_), .B(new_new_n192_), .Y(new_new_n483_));
  NO2        g0461(.A(i_6_), .B(i_10_), .Y(new_new_n484_));
  NA4        g0462(.A(new_new_n484_), .B(new_new_n308_), .C(new_new_n483_), .D(new_new_n235_), .Y(new_new_n485_));
  NO2        g0463(.A(new_new_n485_), .B(new_new_n153_), .Y(new_new_n486_));
  NA2        g0464(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n487_));
  NO2        g0465(.A(new_new_n155_), .B(i_3_), .Y(new_new_n488_));
  NAi31      g0466(.An(new_new_n487_), .B(new_new_n488_), .C(new_new_n224_), .Y(new_new_n489_));
  NA3        g0467(.A(new_new_n395_), .B(new_new_n177_), .C(new_new_n147_), .Y(new_new_n490_));
  NA2        g0468(.A(new_new_n490_), .B(new_new_n489_), .Y(new_new_n491_));
  NO4        g0469(.A(new_new_n491_), .B(new_new_n486_), .C(new_new_n482_), .D(new_new_n472_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n453_), .B(new_new_n383_), .Y(new_new_n493_));
  NA2        g0471(.A(new_new_n459_), .B(new_new_n390_), .Y(new_new_n494_));
  OAI220     g0472(.A0(new_new_n494_), .A1(new_new_n222_), .B0(new_new_n493_), .B1(new_new_n56_), .Y(new_new_n495_));
  NAi21      g0473(.An(new_new_n215_), .B(new_new_n399_), .Y(new_new_n496_));
  NA2        g0474(.A(new_new_n333_), .B(new_new_n217_), .Y(new_new_n497_));
  NO2        g0475(.A(new_new_n26_), .B(i_5_), .Y(new_new_n498_));
  NO2        g0476(.A(i_0_), .B(new_new_n83_), .Y(new_new_n499_));
  NA3        g0477(.A(new_new_n499_), .B(new_new_n498_), .C(new_new_n140_), .Y(new_new_n500_));
  OR3        g0478(.A(new_new_n298_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n501_));
  OAI220     g0479(.A0(new_new_n501_), .A1(new_new_n500_), .B0(new_new_n497_), .B1(new_new_n496_), .Y(new_new_n502_));
  NA4        g0480(.A(new_new_n301_), .B(new_new_n221_), .C(new_new_n72_), .D(new_new_n235_), .Y(new_new_n503_));
  NO2        g0481(.A(new_new_n503_), .B(new_new_n475_), .Y(new_new_n504_));
  NO3        g0482(.A(new_new_n504_), .B(new_new_n502_), .C(new_new_n495_), .Y(new_new_n505_));
  NA4        g0483(.A(new_new_n505_), .B(new_new_n492_), .C(new_new_n467_), .D(new_new_n464_), .Y(new_new_n506_));
  NA2        g0484(.A(new_new_n301_), .B(new_new_n174_), .Y(new_new_n507_));
  OAI210     g0485(.A0(new_new_n296_), .A1(new_new_n179_), .B0(new_new_n507_), .Y(new_new_n508_));
  AN2        g0486(.A(new_new_n282_), .B(new_new_n232_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n509_), .B(new_new_n508_), .Y(new_new_n510_));
  NA2        g0488(.A(new_new_n120_), .B(new_new_n109_), .Y(new_new_n511_));
  AN2        g0489(.A(new_new_n511_), .B(new_new_n453_), .Y(new_new_n512_));
  NA2        g0490(.A(new_new_n308_), .B(new_new_n162_), .Y(new_new_n513_));
  OAI210     g0491(.A0(new_new_n513_), .A1(new_new_n230_), .B0(new_new_n302_), .Y(new_new_n514_));
  AOI220     g0492(.A0(new_new_n514_), .A1(new_new_n320_), .B0(new_new_n512_), .B1(new_new_n304_), .Y(new_new_n515_));
  NA4        g0493(.A(new_new_n443_), .B(new_new_n442_), .C(new_new_n202_), .D(i_2_), .Y(new_new_n516_));
  INV        g0494(.A(new_new_n516_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n356_), .B(new_new_n72_), .Y(new_new_n518_));
  NA2        g0496(.A(new_new_n373_), .B(new_new_n366_), .Y(new_new_n519_));
  NO2        g0497(.A(new_new_n36_), .B(i_8_), .Y(new_new_n520_));
  NA2        g0498(.A(new_new_n39_), .B(i_13_), .Y(new_new_n521_));
  INV        g0499(.A(new_new_n521_), .Y(new_new_n522_));
  AOI210     g0500(.A0(new_new_n517_), .A1(new_new_n203_), .B0(new_new_n522_), .Y(new_new_n523_));
  NA2        g0501(.A(new_new_n254_), .B(new_new_n63_), .Y(new_new_n524_));
  OAI210     g0502(.A0(i_8_), .A1(new_new_n524_), .B0(new_new_n132_), .Y(new_new_n525_));
  NO2        g0503(.A(i_7_), .B(new_new_n198_), .Y(new_new_n526_));
  OR2        g0504(.A(new_new_n181_), .B(i_4_), .Y(new_new_n527_));
  NO2        g0505(.A(new_new_n527_), .B(new_new_n83_), .Y(new_new_n528_));
  AOI220     g0506(.A0(new_new_n528_), .A1(new_new_n526_), .B0(new_new_n525_), .B1(new_new_n416_), .Y(new_new_n529_));
  NA4        g0507(.A(new_new_n529_), .B(new_new_n523_), .C(new_new_n515_), .D(new_new_n510_), .Y(new_new_n530_));
  NA2        g0508(.A(new_new_n389_), .B(new_new_n290_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n385_), .B(new_new_n531_), .Y(new_new_n532_));
  NA2        g0510(.A(new_new_n1047_), .B(new_new_n223_), .Y(new_new_n533_));
  NA2        g0511(.A(new_new_n484_), .B(new_new_n27_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n534_), .B(new_new_n533_), .Y(new_new_n535_));
  NOi31      g0513(.An(new_new_n311_), .B(new_new_n415_), .C(new_new_n38_), .Y(new_new_n536_));
  OAI210     g0514(.A0(new_new_n536_), .A1(new_new_n535_), .B0(new_new_n532_), .Y(new_new_n537_));
  NO2        g0515(.A(i_8_), .B(i_7_), .Y(new_new_n538_));
  OAI210     g0516(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n539_));
  NA2        g0517(.A(new_new_n539_), .B(new_new_n221_), .Y(new_new_n540_));
  OAI220     g0518(.A0(new_new_n46_), .A1(new_new_n527_), .B0(new_new_n540_), .B1(new_new_n240_), .Y(new_new_n541_));
  NA2        g0519(.A(new_new_n44_), .B(i_10_), .Y(new_new_n542_));
  NO2        g0520(.A(new_new_n542_), .B(i_6_), .Y(new_new_n543_));
  NA3        g0521(.A(new_new_n543_), .B(new_new_n541_), .C(new_new_n538_), .Y(new_new_n544_));
  AOI220     g0522(.A0(new_new_n426_), .A1(new_new_n321_), .B0(new_new_n245_), .B1(new_new_n242_), .Y(new_new_n545_));
  OAI220     g0523(.A0(new_new_n545_), .A1(new_new_n257_), .B0(new_new_n468_), .B1(new_new_n131_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n546_), .B(new_new_n260_), .Y(new_new_n547_));
  NOi31      g0525(.An(new_new_n285_), .B(new_new_n296_), .C(new_new_n179_), .Y(new_new_n548_));
  NA3        g0526(.A(new_new_n301_), .B(new_new_n172_), .C(new_new_n93_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n220_), .B(new_new_n44_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n155_), .B(i_5_), .Y(new_new_n551_));
  NA2        g0529(.A(new_new_n551_), .B(new_new_n314_), .Y(new_new_n552_));
  OAI210     g0530(.A0(new_new_n552_), .A1(new_new_n550_), .B0(new_new_n549_), .Y(new_new_n553_));
  OAI210     g0531(.A0(new_new_n553_), .A1(new_new_n548_), .B0(new_new_n459_), .Y(new_new_n554_));
  NA4        g0532(.A(new_new_n554_), .B(new_new_n547_), .C(new_new_n544_), .D(new_new_n537_), .Y(new_new_n555_));
  NA2        g0533(.A(new_new_n279_), .B(new_new_n82_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n346_), .B(new_new_n556_), .Y(new_new_n557_));
  NA2        g0535(.A(new_new_n291_), .B(new_new_n282_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n558_), .B(new_new_n171_), .Y(new_new_n559_));
  NA2        g0537(.A(i_0_), .B(new_new_n48_), .Y(new_new_n560_));
  NO2        g0538(.A(new_new_n559_), .B(new_new_n557_), .Y(new_new_n561_));
  NO4        g0539(.A(new_new_n250_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n562_));
  NO3        g0540(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n231_), .B(new_new_n36_), .Y(new_new_n564_));
  AN2        g0542(.A(new_new_n564_), .B(new_new_n563_), .Y(new_new_n565_));
  OA210      g0543(.A0(new_new_n565_), .A1(new_new_n562_), .B0(new_new_n356_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n415_), .B(i_1_), .Y(new_new_n567_));
  NOi31      g0545(.An(new_new_n567_), .B(new_new_n454_), .C(new_new_n72_), .Y(new_new_n568_));
  AN4        g0546(.A(new_new_n568_), .B(new_new_n413_), .C(new_new_n498_), .D(i_2_), .Y(new_new_n569_));
  NO2        g0547(.A(new_new_n424_), .B(new_new_n175_), .Y(new_new_n570_));
  NO3        g0548(.A(new_new_n570_), .B(new_new_n569_), .C(new_new_n566_), .Y(new_new_n571_));
  NOi21      g0549(.An(i_10_), .B(i_6_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n83_), .B(new_new_n25_), .Y(new_new_n573_));
  AOI220     g0551(.A0(new_new_n279_), .A1(new_new_n573_), .B0(new_new_n270_), .B1(new_new_n572_), .Y(new_new_n574_));
  NO2        g0552(.A(new_new_n574_), .B(new_new_n452_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n112_), .B(new_new_n23_), .Y(new_new_n576_));
  NA2        g0554(.A(new_new_n311_), .B(new_new_n162_), .Y(new_new_n577_));
  AOI220     g0555(.A0(new_new_n577_), .A1(new_new_n433_), .B0(new_new_n182_), .B1(new_new_n180_), .Y(new_new_n578_));
  NOi21      g0556(.An(new_new_n144_), .B(new_new_n328_), .Y(new_new_n579_));
  NO3        g0557(.A(new_new_n579_), .B(new_new_n578_), .C(new_new_n575_), .Y(new_new_n580_));
  NO2        g0558(.A(new_new_n518_), .B(new_new_n378_), .Y(new_new_n581_));
  INV        g0559(.A(new_new_n314_), .Y(new_new_n582_));
  NO2        g0560(.A(i_12_), .B(new_new_n83_), .Y(new_new_n583_));
  NA3        g0561(.A(new_new_n583_), .B(new_new_n270_), .C(new_new_n560_), .Y(new_new_n584_));
  NA3        g0562(.A(new_new_n386_), .B(new_new_n279_), .C(new_new_n217_), .Y(new_new_n585_));
  AOI210     g0563(.A0(new_new_n585_), .A1(new_new_n584_), .B0(new_new_n582_), .Y(new_new_n586_));
  NO3        g0564(.A(i_4_), .B(new_new_n339_), .C(new_new_n296_), .Y(new_new_n587_));
  NO3        g0565(.A(new_new_n587_), .B(new_new_n586_), .C(new_new_n581_), .Y(new_new_n588_));
  NA4        g0566(.A(new_new_n588_), .B(new_new_n580_), .C(new_new_n571_), .D(new_new_n561_), .Y(new_new_n589_));
  NO4        g0567(.A(new_new_n589_), .B(new_new_n555_), .C(new_new_n530_), .D(new_new_n506_), .Y(new_new_n590_));
  NA4        g0568(.A(new_new_n590_), .B(new_new_n441_), .C(new_new_n355_), .D(new_new_n307_), .Y(zz07));
  NO2        g0569(.A(new_new_n90_), .B(new_new_n54_), .Y(new_new_n592_));
  NO2        g0570(.A(new_new_n105_), .B(new_new_n87_), .Y(new_new_n593_));
  NA2        g0571(.A(new_new_n384_), .B(new_new_n593_), .Y(new_new_n594_));
  NA2        g0572(.A(i_11_), .B(new_new_n192_), .Y(new_new_n595_));
  INV        g0573(.A(new_new_n594_), .Y(new_new_n596_));
  NA3        g0574(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n597_));
  NO2        g0575(.A(new_new_n235_), .B(i_4_), .Y(new_new_n598_));
  NA2        g0576(.A(new_new_n598_), .B(i_8_), .Y(new_new_n599_));
  NO2        g0577(.A(new_new_n102_), .B(new_new_n597_), .Y(new_new_n600_));
  NA2        g0578(.A(i_2_), .B(new_new_n83_), .Y(new_new_n601_));
  OAI210     g0579(.A0(new_new_n86_), .A1(new_new_n202_), .B0(new_new_n203_), .Y(new_new_n602_));
  NO2        g0580(.A(i_7_), .B(new_new_n37_), .Y(new_new_n603_));
  NA2        g0581(.A(i_4_), .B(i_8_), .Y(new_new_n604_));
  AOI210     g0582(.A0(new_new_n604_), .A1(new_new_n301_), .B0(new_new_n603_), .Y(new_new_n605_));
  OAI220     g0583(.A0(new_new_n605_), .A1(new_new_n601_), .B0(new_new_n602_), .B1(i_13_), .Y(new_new_n606_));
  NO4        g0584(.A(new_new_n606_), .B(new_new_n600_), .C(new_new_n596_), .D(new_new_n592_), .Y(new_new_n607_));
  AOI210     g0585(.A0(new_new_n126_), .A1(new_new_n61_), .B0(i_10_), .Y(new_new_n608_));
  AOI210     g0586(.A0(new_new_n608_), .A1(new_new_n235_), .B0(new_new_n159_), .Y(new_new_n609_));
  OR2        g0587(.A(i_6_), .B(i_10_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n610_), .B(new_new_n23_), .Y(new_new_n611_));
  OR3        g0589(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n612_));
  NO3        g0590(.A(new_new_n612_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n613_));
  INV        g0591(.A(new_new_n199_), .Y(new_new_n614_));
  NO2        g0592(.A(new_new_n613_), .B(new_new_n611_), .Y(new_new_n615_));
  OA220      g0593(.A0(new_new_n615_), .A1(new_new_n582_), .B0(new_new_n609_), .B1(new_new_n262_), .Y(new_new_n616_));
  AOI210     g0594(.A0(new_new_n616_), .A1(new_new_n607_), .B0(new_new_n62_), .Y(new_new_n617_));
  NOi21      g0595(.An(i_11_), .B(i_7_), .Y(new_new_n618_));
  AO210      g0596(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n619_));
  NO2        g0597(.A(new_new_n619_), .B(new_new_n618_), .Y(new_new_n620_));
  NA2        g0598(.A(new_new_n620_), .B(new_new_n205_), .Y(new_new_n621_));
  NA3        g0599(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n622_));
  NAi31      g0600(.An(new_new_n622_), .B(new_new_n214_), .C(i_11_), .Y(new_new_n623_));
  AOI210     g0601(.A0(new_new_n623_), .A1(new_new_n621_), .B0(new_new_n62_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n85_), .B(new_new_n62_), .Y(new_new_n625_));
  AO210      g0603(.A0(new_new_n625_), .A1(new_new_n378_), .B0(new_new_n41_), .Y(new_new_n626_));
  NA2        g0604(.A(new_new_n224_), .B(new_new_n62_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n409_), .B(new_new_n31_), .Y(new_new_n628_));
  OR2        g0606(.A(new_new_n207_), .B(new_new_n105_), .Y(new_new_n629_));
  NA2        g0607(.A(new_new_n629_), .B(new_new_n628_), .Y(new_new_n630_));
  NO2        g0608(.A(new_new_n62_), .B(i_9_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n631_), .B(i_4_), .Y(new_new_n632_));
  NA2        g0610(.A(new_new_n632_), .B(new_new_n630_), .Y(new_new_n633_));
  NO2        g0611(.A(i_1_), .B(i_12_), .Y(new_new_n634_));
  NA3        g0612(.A(new_new_n633_), .B(new_new_n627_), .C(new_new_n626_), .Y(new_new_n635_));
  OAI210     g0613(.A0(new_new_n635_), .A1(new_new_n624_), .B0(i_6_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n235_), .B(new_new_n83_), .Y(new_new_n637_));
  NO2        g0615(.A(new_new_n637_), .B(i_11_), .Y(new_new_n638_));
  INV        g0616(.A(new_new_n455_), .Y(new_new_n639_));
  NO4        g0617(.A(new_new_n214_), .B(new_new_n126_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n640_));
  NA2        g0618(.A(new_new_n640_), .B(new_new_n631_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n235_), .B(i_6_), .Y(new_new_n642_));
  NO3        g0620(.A(new_new_n610_), .B(new_new_n231_), .C(new_new_n23_), .Y(new_new_n643_));
  INV        g0621(.A(new_new_n641_), .Y(new_new_n644_));
  NA3        g0622(.A(new_new_n538_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n645_));
  NA2        g0623(.A(new_new_n136_), .B(i_9_), .Y(new_new_n646_));
  NA3        g0624(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n46_), .B(i_1_), .Y(new_new_n648_));
  NA3        g0626(.A(new_new_n648_), .B(new_new_n261_), .C(new_new_n44_), .Y(new_new_n649_));
  OAI220     g0627(.A0(new_new_n649_), .A1(new_new_n647_), .B0(new_new_n646_), .B1(new_new_n1045_), .Y(new_new_n650_));
  NA3        g0628(.A(new_new_n631_), .B(new_new_n314_), .C(i_6_), .Y(new_new_n651_));
  NO2        g0629(.A(new_new_n651_), .B(new_new_n23_), .Y(new_new_n652_));
  AOI210     g0630(.A0(new_new_n476_), .A1(new_new_n418_), .B0(new_new_n239_), .Y(new_new_n653_));
  NO2        g0631(.A(new_new_n653_), .B(new_new_n601_), .Y(new_new_n654_));
  NAi21      g0632(.An(new_new_n645_), .B(new_new_n89_), .Y(new_new_n655_));
  NA2        g0633(.A(new_new_n648_), .B(new_new_n261_), .Y(new_new_n656_));
  NO2        g0634(.A(i_11_), .B(new_new_n37_), .Y(new_new_n657_));
  NA2        g0635(.A(new_new_n657_), .B(new_new_n24_), .Y(new_new_n658_));
  OAI210     g0636(.A0(new_new_n658_), .A1(new_new_n656_), .B0(new_new_n655_), .Y(new_new_n659_));
  OR4        g0637(.A(new_new_n659_), .B(new_new_n654_), .C(new_new_n652_), .D(new_new_n650_), .Y(new_new_n660_));
  NO3        g0638(.A(new_new_n660_), .B(new_new_n644_), .C(new_new_n639_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n235_), .B(new_new_n98_), .Y(new_new_n662_));
  NO2        g0640(.A(new_new_n662_), .B(new_new_n618_), .Y(new_new_n663_));
  NA2        g0641(.A(new_new_n663_), .B(i_1_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n664_), .B(new_new_n612_), .Y(new_new_n665_));
  NA2        g0643(.A(new_new_n665_), .B(new_new_n46_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n115_), .B(new_new_n37_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n83_), .B(i_9_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n62_), .Y(new_new_n669_));
  NA2        g0647(.A(i_1_), .B(i_3_), .Y(new_new_n670_));
  NA3        g0648(.A(new_new_n666_), .B(new_new_n661_), .C(new_new_n636_), .Y(new_new_n671_));
  NO3        g0649(.A(new_new_n477_), .B(i_3_), .C(i_7_), .Y(new_new_n672_));
  NOi21      g0650(.An(new_new_n672_), .B(i_10_), .Y(new_new_n673_));
  OA210      g0651(.A0(new_new_n673_), .A1(new_new_n243_), .B0(new_new_n83_), .Y(new_new_n674_));
  NA3        g0652(.A(new_new_n484_), .B(new_new_n520_), .C(new_new_n46_), .Y(new_new_n675_));
  NO3        g0653(.A(new_new_n478_), .B(new_new_n604_), .C(new_new_n83_), .Y(new_new_n676_));
  NA2        g0654(.A(new_new_n676_), .B(new_new_n25_), .Y(new_new_n677_));
  NA3        g0655(.A(new_new_n159_), .B(new_new_n82_), .C(new_new_n83_), .Y(new_new_n678_));
  NA3        g0656(.A(new_new_n678_), .B(new_new_n677_), .C(new_new_n675_), .Y(new_new_n679_));
  OAI210     g0657(.A0(new_new_n679_), .A1(new_new_n674_), .B0(i_1_), .Y(new_new_n680_));
  AOI210     g0658(.A0(new_new_n261_), .A1(new_new_n94_), .B0(i_1_), .Y(new_new_n681_));
  NO2        g0659(.A(new_new_n372_), .B(i_2_), .Y(new_new_n682_));
  NA2        g0660(.A(new_new_n682_), .B(new_new_n681_), .Y(new_new_n683_));
  OAI210     g0661(.A0(new_new_n651_), .A1(new_new_n446_), .B0(new_new_n683_), .Y(new_new_n684_));
  INV        g0662(.A(new_new_n684_), .Y(new_new_n685_));
  AOI210     g0663(.A0(new_new_n685_), .A1(new_new_n680_), .B0(i_13_), .Y(new_new_n686_));
  OR2        g0664(.A(i_11_), .B(i_7_), .Y(new_new_n687_));
  NA3        g0665(.A(new_new_n687_), .B(new_new_n103_), .C(new_new_n136_), .Y(new_new_n688_));
  AOI220     g0666(.A0(new_new_n470_), .A1(new_new_n159_), .B0(new_new_n449_), .B1(new_new_n136_), .Y(new_new_n689_));
  OAI210     g0667(.A0(new_new_n689_), .A1(new_new_n44_), .B0(new_new_n688_), .Y(new_new_n690_));
  AOI210     g0668(.A0(new_new_n647_), .A1(new_new_n54_), .B0(i_12_), .Y(new_new_n691_));
  NA2        g0669(.A(new_new_n243_), .B(new_new_n129_), .Y(new_new_n692_));
  OAI220     g0670(.A0(new_new_n692_), .A1(new_new_n41_), .B0(new_new_n1044_), .B1(new_new_n90_), .Y(new_new_n693_));
  AOI210     g0671(.A0(new_new_n690_), .A1(new_new_n330_), .B0(new_new_n693_), .Y(new_new_n694_));
  NA2        g0672(.A(new_new_n112_), .B(new_new_n105_), .Y(new_new_n695_));
  AOI220     g0673(.A0(new_new_n695_), .A1(new_new_n71_), .B0(new_new_n386_), .B1(new_new_n648_), .Y(new_new_n696_));
  NO2        g0674(.A(new_new_n696_), .B(new_new_n240_), .Y(new_new_n697_));
  AOI210     g0675(.A0(new_new_n446_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n125_), .B(i_13_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n647_), .B(new_new_n112_), .Y(new_new_n700_));
  INV        g0678(.A(new_new_n700_), .Y(new_new_n701_));
  OAI220     g0679(.A0(new_new_n701_), .A1(new_new_n70_), .B0(new_new_n699_), .B1(new_new_n681_), .Y(new_new_n702_));
  NO3        g0680(.A(new_new_n70_), .B(new_new_n32_), .C(new_new_n98_), .Y(new_new_n703_));
  NA2        g0681(.A(new_new_n26_), .B(new_new_n192_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n704_), .B(i_7_), .Y(new_new_n705_));
  NO3        g0683(.A(new_new_n478_), .B(new_new_n235_), .C(new_new_n83_), .Y(new_new_n706_));
  AOI210     g0684(.A0(new_new_n706_), .A1(new_new_n705_), .B0(new_new_n703_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n89_), .B(new_new_n99_), .Y(new_new_n708_));
  OAI220     g0686(.A0(new_new_n708_), .A1(new_new_n599_), .B0(new_new_n707_), .B1(new_new_n614_), .Y(new_new_n709_));
  NO3        g0687(.A(new_new_n709_), .B(new_new_n702_), .C(new_new_n697_), .Y(new_new_n710_));
  OR2        g0688(.A(i_11_), .B(i_6_), .Y(new_new_n711_));
  NA3        g0689(.A(new_new_n598_), .B(new_new_n704_), .C(i_7_), .Y(new_new_n712_));
  AOI210     g0690(.A0(new_new_n712_), .A1(new_new_n701_), .B0(new_new_n711_), .Y(new_new_n713_));
  NA3        g0691(.A(new_new_n409_), .B(new_new_n603_), .C(new_new_n94_), .Y(new_new_n714_));
  NA2        g0692(.A(new_new_n638_), .B(i_13_), .Y(new_new_n715_));
  NA2        g0693(.A(new_new_n99_), .B(new_new_n704_), .Y(new_new_n716_));
  NAi21      g0694(.An(i_11_), .B(i_12_), .Y(new_new_n717_));
  NOi41      g0695(.An(new_new_n108_), .B(new_new_n717_), .C(i_13_), .D(new_new_n83_), .Y(new_new_n718_));
  NO3        g0696(.A(new_new_n478_), .B(new_new_n583_), .C(new_new_n604_), .Y(new_new_n719_));
  AOI220     g0697(.A0(new_new_n719_), .A1(new_new_n308_), .B0(new_new_n718_), .B1(new_new_n716_), .Y(new_new_n720_));
  NA3        g0698(.A(new_new_n720_), .B(new_new_n715_), .C(new_new_n714_), .Y(new_new_n721_));
  OAI210     g0699(.A0(new_new_n721_), .A1(new_new_n713_), .B0(new_new_n62_), .Y(new_new_n722_));
  NO2        g0700(.A(i_2_), .B(i_12_), .Y(new_new_n723_));
  NA2        g0701(.A(new_new_n371_), .B(new_new_n723_), .Y(new_new_n724_));
  NA2        g0702(.A(i_8_), .B(new_new_n25_), .Y(new_new_n725_));
  NO3        g0703(.A(new_new_n725_), .B(new_new_n384_), .C(new_new_n598_), .Y(new_new_n726_));
  NA2        g0704(.A(new_new_n726_), .B(new_new_n371_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n126_), .B(i_2_), .Y(new_new_n728_));
  NA2        g0706(.A(new_new_n728_), .B(new_new_n634_), .Y(new_new_n729_));
  NA3        g0707(.A(new_new_n729_), .B(new_new_n727_), .C(new_new_n724_), .Y(new_new_n730_));
  NA3        g0708(.A(new_new_n730_), .B(new_new_n45_), .C(new_new_n223_), .Y(new_new_n731_));
  NA4        g0709(.A(new_new_n731_), .B(new_new_n722_), .C(new_new_n710_), .D(new_new_n694_), .Y(new_new_n732_));
  OR4        g0710(.A(new_new_n732_), .B(new_new_n686_), .C(new_new_n671_), .D(new_new_n617_), .Y(zz05));
  AOI210     g0711(.A0(new_new_n663_), .A1(new_new_n264_), .B0(new_new_n416_), .Y(new_new_n734_));
  AN2        g0712(.A(new_new_n24_), .B(i_10_), .Y(new_new_n735_));
  NA3        g0713(.A(new_new_n735_), .B(new_new_n723_), .C(new_new_n105_), .Y(new_new_n736_));
  NO2        g0714(.A(new_new_n599_), .B(i_11_), .Y(new_new_n737_));
  OAI210     g0715(.A0(new_new_n603_), .A1(new_new_n86_), .B0(new_new_n737_), .Y(new_new_n738_));
  NA3        g0716(.A(new_new_n738_), .B(new_new_n736_), .C(new_new_n734_), .Y(new_new_n739_));
  NO3        g0717(.A(i_11_), .B(new_new_n235_), .C(i_13_), .Y(new_new_n740_));
  NO2        g0718(.A(new_new_n122_), .B(new_new_n23_), .Y(new_new_n741_));
  NA2        g0719(.A(i_12_), .B(i_8_), .Y(new_new_n742_));
  OAI210     g0720(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n742_), .Y(new_new_n743_));
  INV        g0721(.A(new_new_n445_), .Y(new_new_n744_));
  AOI220     g0722(.A0(new_new_n314_), .A1(new_new_n576_), .B0(new_new_n743_), .B1(new_new_n741_), .Y(new_new_n745_));
  INV        g0723(.A(new_new_n745_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n746_), .B(new_new_n739_), .Y(new_new_n747_));
  INV        g0725(.A(new_new_n169_), .Y(new_new_n748_));
  INV        g0726(.A(new_new_n243_), .Y(new_new_n749_));
  OAI210     g0727(.A0(new_new_n682_), .A1(new_new_n447_), .B0(new_new_n108_), .Y(new_new_n750_));
  AOI210     g0728(.A0(new_new_n750_), .A1(new_new_n749_), .B0(new_new_n748_), .Y(new_new_n751_));
  NO2        g0729(.A(new_new_n456_), .B(new_new_n26_), .Y(new_new_n752_));
  NO2        g0730(.A(new_new_n752_), .B(new_new_n418_), .Y(new_new_n753_));
  NA2        g0731(.A(new_new_n753_), .B(i_2_), .Y(new_new_n754_));
  INV        g0732(.A(new_new_n754_), .Y(new_new_n755_));
  AOI210     g0733(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n415_), .Y(new_new_n756_));
  AOI210     g0734(.A0(new_new_n756_), .A1(new_new_n755_), .B0(new_new_n751_), .Y(new_new_n757_));
  NO2        g0735(.A(new_new_n189_), .B(new_new_n123_), .Y(new_new_n758_));
  OAI210     g0736(.A0(new_new_n758_), .A1(new_new_n741_), .B0(i_2_), .Y(new_new_n759_));
  INV        g0737(.A(new_new_n170_), .Y(new_new_n760_));
  NO3        g0738(.A(new_new_n619_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n761_));
  AOI210     g0739(.A0(new_new_n760_), .A1(new_new_n86_), .B0(new_new_n761_), .Y(new_new_n762_));
  AOI210     g0740(.A0(new_new_n762_), .A1(new_new_n759_), .B0(new_new_n192_), .Y(new_new_n763_));
  OA210      g0741(.A0(new_new_n620_), .A1(new_new_n124_), .B0(i_13_), .Y(new_new_n764_));
  NA2        g0742(.A(new_new_n199_), .B(new_new_n202_), .Y(new_new_n765_));
  NA2        g0743(.A(new_new_n149_), .B(new_new_n595_), .Y(new_new_n766_));
  AOI210     g0744(.A0(new_new_n766_), .A1(new_new_n765_), .B0(new_new_n374_), .Y(new_new_n767_));
  AOI210     g0745(.A0(new_new_n207_), .A1(new_new_n146_), .B0(new_new_n520_), .Y(new_new_n768_));
  OAI210     g0746(.A0(new_new_n768_), .A1(new_new_n224_), .B0(new_new_n418_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n99_), .B(new_new_n44_), .Y(new_new_n770_));
  INV        g0748(.A(new_new_n297_), .Y(new_new_n771_));
  NA4        g0749(.A(new_new_n771_), .B(new_new_n301_), .C(new_new_n122_), .D(new_new_n42_), .Y(new_new_n772_));
  OAI210     g0750(.A0(new_new_n772_), .A1(new_new_n770_), .B0(new_new_n769_), .Y(new_new_n773_));
  NO4        g0751(.A(new_new_n773_), .B(new_new_n767_), .C(new_new_n764_), .D(new_new_n763_), .Y(new_new_n774_));
  NA2        g0752(.A(new_new_n576_), .B(new_new_n28_), .Y(new_new_n775_));
  NA2        g0753(.A(new_new_n740_), .B(new_new_n271_), .Y(new_new_n776_));
  NA2        g0754(.A(new_new_n776_), .B(new_new_n775_), .Y(new_new_n777_));
  NO2        g0755(.A(new_new_n61_), .B(i_12_), .Y(new_new_n778_));
  NO2        g0756(.A(new_new_n778_), .B(new_new_n124_), .Y(new_new_n779_));
  NO2        g0757(.A(new_new_n779_), .B(new_new_n595_), .Y(new_new_n780_));
  AOI220     g0758(.A0(new_new_n780_), .A1(new_new_n36_), .B0(new_new_n777_), .B1(new_new_n46_), .Y(new_new_n781_));
  NA4        g0759(.A(new_new_n781_), .B(new_new_n774_), .C(new_new_n757_), .D(new_new_n747_), .Y(zz06));
  NO3        g0760(.A(new_new_n252_), .B(new_new_n303_), .C(i_1_), .Y(new_new_n783_));
  NO2        g0761(.A(new_new_n184_), .B(new_new_n137_), .Y(new_new_n784_));
  OAI210     g0762(.A0(new_new_n784_), .A1(new_new_n783_), .B0(new_new_n728_), .Y(new_new_n785_));
  NA4        g0763(.A(new_new_n390_), .B(new_new_n483_), .C(new_new_n70_), .D(new_new_n98_), .Y(new_new_n786_));
  INV        g0764(.A(new_new_n786_), .Y(new_new_n787_));
  NO2        g0765(.A(i_11_), .B(i_9_), .Y(new_new_n788_));
  NO2        g0766(.A(new_new_n787_), .B(new_new_n326_), .Y(new_new_n789_));
  AO210      g0767(.A0(new_new_n789_), .A1(new_new_n785_), .B0(i_12_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n375_), .B(new_new_n333_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n583_), .B(new_new_n62_), .Y(new_new_n792_));
  NA2        g0770(.A(new_new_n673_), .B(new_new_n70_), .Y(new_new_n793_));
  BUFFER     g0771(.A(new_new_n625_), .Y(new_new_n794_));
  NA4        g0772(.A(new_new_n794_), .B(new_new_n793_), .C(new_new_n792_), .D(new_new_n791_), .Y(new_new_n795_));
  INV        g0773(.A(new_new_n196_), .Y(new_new_n796_));
  AOI220     g0774(.A0(new_new_n796_), .A1(new_new_n788_), .B0(new_new_n795_), .B1(new_new_n72_), .Y(new_new_n797_));
  INV        g0775(.A(new_new_n325_), .Y(new_new_n798_));
  NA2        g0776(.A(new_new_n74_), .B(new_new_n129_), .Y(new_new_n799_));
  INV        g0777(.A(new_new_n122_), .Y(new_new_n800_));
  NA2        g0778(.A(new_new_n800_), .B(new_new_n46_), .Y(new_new_n801_));
  AOI210     g0779(.A0(new_new_n801_), .A1(new_new_n799_), .B0(new_new_n798_), .Y(new_new_n802_));
  NO2        g0780(.A(new_new_n250_), .B(i_9_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n803_), .B(new_new_n778_), .Y(new_new_n804_));
  AOI210     g0782(.A0(new_new_n804_), .A1(new_new_n519_), .B0(new_new_n184_), .Y(new_new_n805_));
  NO2        g0783(.A(new_new_n32_), .B(i_11_), .Y(new_new_n806_));
  NA3        g0784(.A(new_new_n806_), .B(new_new_n474_), .C(new_new_n390_), .Y(new_new_n807_));
  NAi32      g0785(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n808_));
  AOI210     g0786(.A0(new_new_n711_), .A1(new_new_n84_), .B0(new_new_n808_), .Y(new_new_n809_));
  OAI210     g0787(.A0(new_new_n672_), .A1(new_new_n564_), .B0(new_new_n563_), .Y(new_new_n810_));
  NAi31      g0788(.An(new_new_n809_), .B(new_new_n810_), .C(new_new_n807_), .Y(new_new_n811_));
  OR3        g0789(.A(new_new_n811_), .B(new_new_n805_), .C(new_new_n802_), .Y(new_new_n812_));
  NO2        g0790(.A(new_new_n687_), .B(i_2_), .Y(new_new_n813_));
  NA2        g0791(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n814_));
  OAI210     g0792(.A0(new_new_n814_), .A1(new_new_n408_), .B0(new_new_n361_), .Y(new_new_n815_));
  NA2        g0793(.A(new_new_n815_), .B(new_new_n813_), .Y(new_new_n816_));
  AO210      g0794(.A0(new_new_n360_), .A1(new_new_n350_), .B0(new_new_n398_), .Y(new_new_n817_));
  NA3        g0795(.A(new_new_n817_), .B(new_new_n253_), .C(i_7_), .Y(new_new_n818_));
  OR2        g0796(.A(new_new_n620_), .B(new_new_n447_), .Y(new_new_n819_));
  NA3        g0797(.A(new_new_n819_), .B(new_new_n145_), .C(new_new_n68_), .Y(new_new_n820_));
  AO210      g0798(.A0(new_new_n494_), .A1(new_new_n744_), .B0(new_new_n36_), .Y(new_new_n821_));
  NA4        g0799(.A(new_new_n821_), .B(new_new_n820_), .C(new_new_n818_), .D(new_new_n816_), .Y(new_new_n822_));
  OAI210     g0800(.A0(new_new_n637_), .A1(i_11_), .B0(new_new_n84_), .Y(new_new_n823_));
  NA2        g0801(.A(new_new_n823_), .B(new_new_n563_), .Y(new_new_n824_));
  OAI210     g0802(.A0(new_new_n398_), .A1(new_new_n203_), .B0(new_new_n69_), .Y(new_new_n825_));
  NA3        g0803(.A(new_new_n825_), .B(new_new_n824_), .C(new_new_n602_), .Y(new_new_n826_));
  AO210      g0804(.A0(new_new_n520_), .A1(new_new_n46_), .B0(new_new_n85_), .Y(new_new_n827_));
  NA3        g0805(.A(new_new_n827_), .B(new_new_n484_), .C(new_new_n217_), .Y(new_new_n828_));
  AOI210     g0806(.A0(new_new_n447_), .A1(new_new_n445_), .B0(new_new_n562_), .Y(new_new_n829_));
  NA2        g0807(.A(new_new_n109_), .B(new_new_n407_), .Y(new_new_n830_));
  NA2        g0808(.A(new_new_n242_), .B(new_new_n46_), .Y(new_new_n831_));
  NA3        g0809(.A(new_new_n830_), .B(new_new_n829_), .C(new_new_n828_), .Y(new_new_n832_));
  NO4        g0810(.A(new_new_n832_), .B(new_new_n826_), .C(new_new_n822_), .D(new_new_n812_), .Y(new_new_n833_));
  NA4        g0811(.A(new_new_n833_), .B(new_new_n797_), .C(new_new_n790_), .D(new_new_n380_), .Y(zz03));
  NA2        g0812(.A(i_6_), .B(i_7_), .Y(new_new_n835_));
  NO2        g0813(.A(new_new_n835_), .B(i_0_), .Y(new_new_n836_));
  NO2        g0814(.A(i_11_), .B(new_new_n235_), .Y(new_new_n837_));
  OAI210     g0815(.A0(new_new_n836_), .A1(new_new_n285_), .B0(new_new_n837_), .Y(new_new_n838_));
  NO2        g0816(.A(new_new_n838_), .B(new_new_n192_), .Y(new_new_n839_));
  NO3        g0817(.A(new_new_n452_), .B(new_new_n87_), .C(new_new_n44_), .Y(new_new_n840_));
  OA210      g0818(.A0(new_new_n840_), .A1(new_new_n839_), .B0(new_new_n172_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n409_), .B(new_new_n45_), .Y(new_new_n842_));
  NO4        g0820(.A(new_new_n376_), .B(new_new_n383_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n843_));
  NA2        g0821(.A(new_new_n184_), .B(new_new_n572_), .Y(new_new_n844_));
  NOi31      g0822(.An(new_new_n844_), .B(new_new_n843_), .C(new_new_n39_), .Y(new_new_n845_));
  NA2        g0823(.A(new_new_n698_), .B(new_new_n668_), .Y(new_new_n846_));
  NA2        g0824(.A(new_new_n331_), .B(new_new_n435_), .Y(new_new_n847_));
  OAI220     g0825(.A0(new_new_n847_), .A1(new_new_n846_), .B0(new_new_n845_), .B1(new_new_n62_), .Y(new_new_n848_));
  NOi21      g0826(.An(i_5_), .B(i_9_), .Y(new_new_n849_));
  NA2        g0827(.A(new_new_n849_), .B(new_new_n443_), .Y(new_new_n850_));
  AOI210     g0828(.A0(new_new_n261_), .A1(new_new_n476_), .B0(new_new_n676_), .Y(new_new_n851_));
  NO3        g0829(.A(new_new_n412_), .B(new_new_n261_), .C(new_new_n72_), .Y(new_new_n852_));
  NO2        g0830(.A(new_new_n173_), .B(new_new_n146_), .Y(new_new_n853_));
  AOI210     g0831(.A0(new_new_n853_), .A1(new_new_n242_), .B0(new_new_n852_), .Y(new_new_n854_));
  OAI220     g0832(.A0(new_new_n854_), .A1(new_new_n179_), .B0(new_new_n851_), .B1(new_new_n850_), .Y(new_new_n855_));
  NO3        g0833(.A(new_new_n855_), .B(new_new_n848_), .C(new_new_n841_), .Y(new_new_n856_));
  NA2        g0834(.A(new_new_n184_), .B(new_new_n24_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n667_), .B(new_new_n593_), .Y(new_new_n858_));
  NO2        g0836(.A(new_new_n858_), .B(new_new_n857_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n308_), .B(new_new_n127_), .Y(new_new_n860_));
  NAi21      g0838(.An(new_new_n160_), .B(new_new_n435_), .Y(new_new_n861_));
  OAI220     g0839(.A0(new_new_n861_), .A1(new_new_n831_), .B0(new_new_n860_), .B1(new_new_n400_), .Y(new_new_n862_));
  NO2        g0840(.A(new_new_n862_), .B(new_new_n859_), .Y(new_new_n863_));
  NO2        g0841(.A(new_new_n390_), .B(new_new_n289_), .Y(new_new_n864_));
  NA2        g0842(.A(new_new_n864_), .B(new_new_n700_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n573_), .B(i_0_), .Y(new_new_n866_));
  NO3        g0844(.A(new_new_n866_), .B(new_new_n385_), .C(new_new_n86_), .Y(new_new_n867_));
  INV        g0845(.A(new_new_n867_), .Y(new_new_n868_));
  AN2        g0846(.A(new_new_n93_), .B(new_new_n241_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n740_), .B(new_new_n326_), .Y(new_new_n870_));
  INV        g0848(.A(new_new_n57_), .Y(new_new_n871_));
  OAI220     g0849(.A0(new_new_n871_), .A1(new_new_n870_), .B0(new_new_n658_), .B1(new_new_n540_), .Y(new_new_n872_));
  NA2        g0850(.A(i_0_), .B(i_10_), .Y(new_new_n873_));
  AOI220     g0851(.A0(new_new_n331_), .A1(new_new_n95_), .B0(new_new_n184_), .B1(new_new_n82_), .Y(new_new_n874_));
  NA2        g0852(.A(new_new_n567_), .B(i_4_), .Y(new_new_n875_));
  NA2        g0853(.A(new_new_n187_), .B(new_new_n202_), .Y(new_new_n876_));
  OAI220     g0854(.A0(new_new_n876_), .A1(new_new_n870_), .B0(new_new_n875_), .B1(new_new_n874_), .Y(new_new_n877_));
  NO3        g0855(.A(new_new_n877_), .B(new_new_n872_), .C(new_new_n869_), .Y(new_new_n878_));
  NA4        g0856(.A(new_new_n878_), .B(new_new_n868_), .C(new_new_n865_), .D(new_new_n863_), .Y(new_new_n879_));
  NA2        g0857(.A(i_11_), .B(i_9_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n48_), .B(i_7_), .Y(new_new_n881_));
  NA2        g0859(.A(new_new_n395_), .B(new_new_n177_), .Y(new_new_n882_));
  NA2        g0860(.A(new_new_n882_), .B(new_new_n158_), .Y(new_new_n883_));
  NO2        g0861(.A(new_new_n880_), .B(new_new_n72_), .Y(new_new_n884_));
  NO2        g0862(.A(new_new_n173_), .B(i_0_), .Y(new_new_n885_));
  INV        g0863(.A(new_new_n885_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n474_), .B(new_new_n229_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n373_), .B(i_4_), .Y(new_new_n888_));
  OAI220     g0866(.A0(new_new_n888_), .A1(new_new_n850_), .B0(new_new_n887_), .B1(new_new_n886_), .Y(new_new_n889_));
  NO2        g0867(.A(new_new_n889_), .B(new_new_n883_), .Y(new_new_n890_));
  NA2        g0868(.A(new_new_n657_), .B(new_new_n119_), .Y(new_new_n891_));
  NO2        g0869(.A(i_6_), .B(new_new_n891_), .Y(new_new_n892_));
  AOI210     g0870(.A0(new_new_n446_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n893_));
  NA2        g0871(.A(new_new_n169_), .B(new_new_n100_), .Y(new_new_n894_));
  NOi32      g0872(.An(new_new_n893_), .Bn(new_new_n187_), .C(new_new_n894_), .Y(new_new_n895_));
  AOI210     g0873(.A0(new_new_n603_), .A1(new_new_n326_), .B0(new_new_n241_), .Y(new_new_n896_));
  NO2        g0874(.A(new_new_n896_), .B(new_new_n842_), .Y(new_new_n897_));
  NO3        g0875(.A(new_new_n897_), .B(new_new_n895_), .C(new_new_n892_), .Y(new_new_n898_));
  NOi21      g0876(.An(i_7_), .B(i_5_), .Y(new_new_n899_));
  NOi31      g0877(.An(new_new_n899_), .B(i_0_), .C(new_new_n717_), .Y(new_new_n900_));
  NA3        g0878(.A(new_new_n900_), .B(new_new_n384_), .C(i_6_), .Y(new_new_n901_));
  OA210      g0879(.A0(new_new_n894_), .A1(new_new_n519_), .B0(new_new_n901_), .Y(new_new_n902_));
  NO3        g0880(.A(new_new_n403_), .B(new_new_n363_), .C(new_new_n359_), .Y(new_new_n903_));
  NO2        g0881(.A(new_new_n255_), .B(new_new_n315_), .Y(new_new_n904_));
  INV        g0882(.A(new_new_n717_), .Y(new_new_n905_));
  AOI210     g0883(.A0(new_new_n905_), .A1(new_new_n904_), .B0(new_new_n903_), .Y(new_new_n906_));
  NA4        g0884(.A(new_new_n906_), .B(new_new_n902_), .C(new_new_n898_), .D(new_new_n890_), .Y(new_new_n907_));
  NO2        g0885(.A(new_new_n857_), .B(new_new_n237_), .Y(new_new_n908_));
  AN2        g0886(.A(new_new_n330_), .B(new_new_n326_), .Y(new_new_n909_));
  AO220      g0887(.A0(new_new_n909_), .A1(new_new_n853_), .B0(new_new_n345_), .B1(new_new_n27_), .Y(new_new_n910_));
  OAI210     g0888(.A0(new_new_n910_), .A1(new_new_n908_), .B0(i_10_), .Y(new_new_n911_));
  OA210      g0889(.A0(new_new_n474_), .A1(new_new_n221_), .B0(new_new_n473_), .Y(new_new_n912_));
  NA3        g0890(.A(new_new_n473_), .B(new_new_n409_), .C(new_new_n45_), .Y(new_new_n913_));
  OAI210     g0891(.A0(new_new_n861_), .A1(i_6_), .B0(new_new_n913_), .Y(new_new_n914_));
  NA2        g0892(.A(new_new_n884_), .B(new_new_n301_), .Y(new_new_n915_));
  NA2        g0893(.A(new_new_n186_), .B(new_new_n915_), .Y(new_new_n916_));
  AOI220     g0894(.A0(new_new_n916_), .A1(new_new_n474_), .B0(new_new_n914_), .B1(new_new_n72_), .Y(new_new_n917_));
  NA3        g0895(.A(new_new_n814_), .B(new_new_n382_), .C(new_new_n637_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n90_), .B(new_new_n44_), .Y(new_new_n919_));
  NO2        g0897(.A(new_new_n74_), .B(new_new_n742_), .Y(new_new_n920_));
  AOI220     g0898(.A0(new_new_n920_), .A1(new_new_n919_), .B0(new_new_n172_), .B1(new_new_n593_), .Y(new_new_n921_));
  AOI210     g0899(.A0(new_new_n921_), .A1(new_new_n918_), .B0(new_new_n47_), .Y(new_new_n922_));
  NO3        g0900(.A(i_5_), .B(new_new_n358_), .C(new_new_n24_), .Y(new_new_n923_));
  INV        g0901(.A(new_new_n923_), .Y(new_new_n924_));
  NAi21      g0902(.An(i_9_), .B(i_5_), .Y(new_new_n925_));
  NO2        g0903(.A(new_new_n597_), .B(new_new_n102_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n926_), .B(i_0_), .Y(new_new_n927_));
  OAI220     g0905(.A0(new_new_n927_), .A1(new_new_n83_), .B0(new_new_n924_), .B1(new_new_n170_), .Y(new_new_n928_));
  NO2        g0906(.A(new_new_n928_), .B(new_new_n922_), .Y(new_new_n929_));
  NA3        g0907(.A(new_new_n929_), .B(new_new_n917_), .C(new_new_n911_), .Y(new_new_n930_));
  NO3        g0908(.A(new_new_n930_), .B(new_new_n907_), .C(new_new_n879_), .Y(new_new_n931_));
  NO2        g0909(.A(i_0_), .B(new_new_n717_), .Y(new_new_n932_));
  NA2        g0910(.A(new_new_n72_), .B(new_new_n44_), .Y(new_new_n933_));
  NA2        g0911(.A(new_new_n873_), .B(new_new_n933_), .Y(new_new_n934_));
  NO3        g0912(.A(new_new_n102_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n935_));
  AO220      g0913(.A0(new_new_n935_), .A1(new_new_n934_), .B0(new_new_n932_), .B1(new_new_n172_), .Y(new_new_n936_));
  NO2        g0914(.A(new_new_n792_), .B(new_new_n894_), .Y(new_new_n937_));
  AOI210     g0915(.A0(new_new_n936_), .A1(new_new_n347_), .B0(new_new_n937_), .Y(new_new_n938_));
  NA2        g0916(.A(new_new_n728_), .B(new_new_n144_), .Y(new_new_n939_));
  INV        g0917(.A(new_new_n939_), .Y(new_new_n940_));
  NA3        g0918(.A(new_new_n940_), .B(new_new_n668_), .C(new_new_n72_), .Y(new_new_n941_));
  NO2        g0919(.A(new_new_n810_), .B(new_new_n403_), .Y(new_new_n942_));
  NA3        g0920(.A(new_new_n836_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n943_));
  NA2        g0921(.A(new_new_n837_), .B(i_9_), .Y(new_new_n944_));
  AOI210     g0922(.A0(new_new_n943_), .A1(new_new_n500_), .B0(new_new_n944_), .Y(new_new_n945_));
  OAI210     g0923(.A0(new_new_n242_), .A1(i_9_), .B0(new_new_n228_), .Y(new_new_n946_));
  AOI210     g0924(.A0(new_new_n946_), .A1(new_new_n866_), .B0(new_new_n151_), .Y(new_new_n947_));
  NO3        g0925(.A(new_new_n947_), .B(new_new_n945_), .C(new_new_n942_), .Y(new_new_n948_));
  NA3        g0926(.A(new_new_n948_), .B(new_new_n941_), .C(new_new_n938_), .Y(new_new_n949_));
  NA2        g0927(.A(new_new_n909_), .B(new_new_n374_), .Y(new_new_n950_));
  AOI210     g0928(.A0(new_new_n296_), .A1(new_new_n160_), .B0(new_new_n950_), .Y(new_new_n951_));
  NA3        g0929(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n44_), .Y(new_new_n952_));
  NA2        g0930(.A(new_new_n881_), .B(new_new_n488_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n952_), .A1(new_new_n160_), .B0(new_new_n953_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n954_), .B(new_new_n951_), .Y(new_new_n955_));
  NO3        g0933(.A(new_new_n873_), .B(new_new_n849_), .C(new_new_n189_), .Y(new_new_n956_));
  AOI220     g0934(.A0(new_new_n956_), .A1(i_11_), .B0(new_new_n568_), .B1(new_new_n74_), .Y(new_new_n957_));
  NO3        g0935(.A(new_new_n208_), .B(new_new_n383_), .C(i_0_), .Y(new_new_n958_));
  OAI210     g0936(.A0(new_new_n958_), .A1(new_new_n75_), .B0(i_13_), .Y(new_new_n959_));
  INV        g0937(.A(new_new_n217_), .Y(new_new_n960_));
  OAI220     g0938(.A0(new_new_n533_), .A1(new_new_n137_), .B0(new_new_n642_), .B1(new_new_n614_), .Y(new_new_n961_));
  NA3        g0939(.A(new_new_n961_), .B(i_7_), .C(new_new_n960_), .Y(new_new_n962_));
  NA4        g0940(.A(new_new_n962_), .B(new_new_n959_), .C(new_new_n957_), .D(new_new_n955_), .Y(new_new_n963_));
  NO2        g0941(.A(new_new_n240_), .B(new_new_n90_), .Y(new_new_n964_));
  AOI210     g0942(.A0(new_new_n964_), .A1(new_new_n932_), .B0(new_new_n106_), .Y(new_new_n965_));
  AOI220     g0943(.A0(new_new_n899_), .A1(new_new_n488_), .B0(new_new_n836_), .B1(new_new_n161_), .Y(new_new_n966_));
  NA2        g0944(.A(new_new_n350_), .B(new_new_n174_), .Y(new_new_n967_));
  OA220      g0945(.A0(new_new_n967_), .A1(new_new_n966_), .B0(new_new_n965_), .B1(i_5_), .Y(new_new_n968_));
  AOI210     g0946(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n173_), .Y(new_new_n969_));
  NA2        g0947(.A(new_new_n969_), .B(new_new_n912_), .Y(new_new_n970_));
  NA3        g0948(.A(new_new_n611_), .B(new_new_n184_), .C(new_new_n82_), .Y(new_new_n971_));
  NA2        g0949(.A(new_new_n971_), .B(new_new_n549_), .Y(new_new_n972_));
  NO3        g0950(.A(new_new_n842_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n493_), .B(new_new_n471_), .Y(new_new_n974_));
  NO3        g0952(.A(new_new_n974_), .B(new_new_n973_), .C(new_new_n972_), .Y(new_new_n975_));
  NA3        g0953(.A(new_new_n390_), .B(new_new_n169_), .C(new_new_n168_), .Y(new_new_n976_));
  NA3        g0954(.A(new_new_n881_), .B(new_new_n285_), .C(new_new_n228_), .Y(new_new_n977_));
  NA2        g0955(.A(new_new_n977_), .B(new_new_n976_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n390_), .B(new_new_n332_), .C(new_new_n220_), .Y(new_new_n979_));
  OAI210     g0957(.A0(new_new_n844_), .A1(new_new_n645_), .B0(new_new_n979_), .Y(new_new_n980_));
  NOi31      g0958(.An(new_new_n389_), .B(new_new_n933_), .C(new_new_n237_), .Y(new_new_n981_));
  NO3        g0959(.A(new_new_n880_), .B(new_new_n217_), .C(new_new_n189_), .Y(new_new_n982_));
  NO4        g0960(.A(new_new_n982_), .B(new_new_n981_), .C(new_new_n980_), .D(new_new_n978_), .Y(new_new_n983_));
  NA4        g0961(.A(new_new_n983_), .B(new_new_n975_), .C(new_new_n970_), .D(new_new_n968_), .Y(new_new_n984_));
  INV        g0962(.A(new_new_n613_), .Y(new_new_n985_));
  NO3        g0963(.A(new_new_n985_), .B(new_new_n560_), .C(new_new_n344_), .Y(new_new_n986_));
  INV        g0964(.A(new_new_n986_), .Y(new_new_n987_));
  NA3        g0965(.A(new_new_n301_), .B(i_5_), .C(new_new_n192_), .Y(new_new_n988_));
  NA2        g0966(.A(new_new_n988_), .B(new_new_n240_), .Y(new_new_n989_));
  NO4        g0967(.A(new_new_n237_), .B(new_new_n208_), .C(i_0_), .D(i_12_), .Y(new_new_n990_));
  AOI220     g0968(.A0(new_new_n990_), .A1(new_new_n989_), .B0(new_new_n787_), .B1(new_new_n174_), .Y(new_new_n991_));
  AN2        g0969(.A(new_new_n873_), .B(new_new_n151_), .Y(new_new_n992_));
  NO4        g0970(.A(new_new_n992_), .B(i_12_), .C(new_new_n645_), .D(new_new_n129_), .Y(new_new_n993_));
  NA2        g0971(.A(new_new_n993_), .B(new_new_n217_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n95_), .B(new_new_n572_), .C(i_11_), .Y(new_new_n995_));
  NO2        g0973(.A(new_new_n995_), .B(new_new_n153_), .Y(new_new_n996_));
  NA2        g0974(.A(new_new_n899_), .B(new_new_n470_), .Y(new_new_n997_));
  OAI220     g0975(.A0(i_7_), .A1(new_new_n988_), .B0(new_new_n997_), .B1(new_new_n669_), .Y(new_new_n998_));
  AOI210     g0976(.A0(new_new_n998_), .A1(new_new_n885_), .B0(new_new_n996_), .Y(new_new_n999_));
  NA4        g0977(.A(new_new_n999_), .B(new_new_n994_), .C(new_new_n991_), .D(new_new_n987_), .Y(new_new_n1000_));
  NO4        g0978(.A(new_new_n1000_), .B(new_new_n984_), .C(new_new_n963_), .D(new_new_n949_), .Y(new_new_n1001_));
  OAI210     g0979(.A0(new_new_n813_), .A1(new_new_n806_), .B0(new_new_n37_), .Y(new_new_n1002_));
  NA3        g0980(.A(new_new_n893_), .B(new_new_n371_), .C(i_5_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n1003_), .B(new_new_n1002_), .C(new_new_n609_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n1004_), .B(new_new_n205_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n185_), .B(new_new_n187_), .Y(new_new_n1006_));
  AO210      g0984(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1006_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n613_), .A1(new_new_n611_), .B0(new_new_n314_), .Y(new_new_n1008_));
  INV        g0986(.A(new_new_n643_), .Y(new_new_n1009_));
  NA3        g0987(.A(new_new_n1009_), .B(new_new_n1008_), .C(new_new_n1007_), .Y(new_new_n1010_));
  NO2        g0988(.A(new_new_n461_), .B(new_new_n261_), .Y(new_new_n1011_));
  NO4        g0989(.A(new_new_n231_), .B(new_new_n143_), .C(new_new_n670_), .D(new_new_n37_), .Y(new_new_n1012_));
  NO2        g0990(.A(new_new_n1012_), .B(new_new_n1011_), .Y(new_new_n1013_));
  OAI210     g0991(.A0(new_new_n995_), .A1(new_new_n146_), .B0(new_new_n1013_), .Y(new_new_n1014_));
  AOI210     g0992(.A0(new_new_n1010_), .A1(new_new_n48_), .B0(new_new_n1014_), .Y(new_new_n1015_));
  AOI210     g0993(.A0(new_new_n1015_), .A1(new_new_n1005_), .B0(new_new_n72_), .Y(new_new_n1016_));
  NO2        g0994(.A(new_new_n565_), .B(new_new_n379_), .Y(new_new_n1017_));
  NO2        g0995(.A(new_new_n1017_), .B(new_new_n748_), .Y(new_new_n1018_));
  INV        g0996(.A(new_new_n75_), .Y(new_new_n1019_));
  AOI210     g0997(.A0(new_new_n969_), .A1(new_new_n881_), .B0(new_new_n900_), .Y(new_new_n1020_));
  AOI210     g0998(.A0(new_new_n1020_), .A1(new_new_n1019_), .B0(new_new_n670_), .Y(new_new_n1021_));
  NA2        g0999(.A(new_new_n255_), .B(new_new_n56_), .Y(new_new_n1022_));
  AOI220     g1000(.A0(new_new_n1022_), .A1(new_new_n75_), .B0(new_new_n345_), .B1(new_new_n252_), .Y(new_new_n1023_));
  NO2        g1001(.A(new_new_n1023_), .B(new_new_n235_), .Y(new_new_n1024_));
  NA3        g1002(.A(new_new_n93_), .B(new_new_n303_), .C(new_new_n31_), .Y(new_new_n1025_));
  INV        g1003(.A(new_new_n1025_), .Y(new_new_n1026_));
  NO3        g1004(.A(new_new_n1026_), .B(new_new_n1024_), .C(new_new_n1021_), .Y(new_new_n1027_));
  OAI210     g1005(.A0(new_new_n263_), .A1(new_new_n156_), .B0(new_new_n86_), .Y(new_new_n1028_));
  NA3        g1006(.A(new_new_n752_), .B(new_new_n285_), .C(new_new_n79_), .Y(new_new_n1029_));
  AOI210     g1007(.A0(new_new_n1029_), .A1(new_new_n1028_), .B0(i_11_), .Y(new_new_n1030_));
  OAI210     g1008(.A0(new_new_n1048_), .A1(new_new_n893_), .B0(new_new_n205_), .Y(new_new_n1031_));
  NA2        g1009(.A(new_new_n162_), .B(i_5_), .Y(new_new_n1032_));
  AOI210     g1010(.A0(new_new_n1031_), .A1(new_new_n765_), .B0(new_new_n1032_), .Y(new_new_n1033_));
  NO4        g1011(.A(new_new_n925_), .B(new_new_n477_), .C(new_new_n251_), .D(new_new_n250_), .Y(new_new_n1034_));
  NO2        g1012(.A(new_new_n1034_), .B(new_new_n562_), .Y(new_new_n1035_));
  NO2        g1013(.A(new_new_n809_), .B(new_new_n364_), .Y(new_new_n1036_));
  AOI210     g1014(.A0(new_new_n1036_), .A1(new_new_n1035_), .B0(new_new_n41_), .Y(new_new_n1037_));
  NO3        g1015(.A(new_new_n1037_), .B(new_new_n1033_), .C(new_new_n1030_), .Y(new_new_n1038_));
  OAI210     g1016(.A0(new_new_n1027_), .A1(i_4_), .B0(new_new_n1038_), .Y(new_new_n1039_));
  NO3        g1017(.A(new_new_n1039_), .B(new_new_n1018_), .C(new_new_n1016_), .Y(new_new_n1040_));
  NA4        g1018(.A(new_new_n1040_), .B(new_new_n1001_), .C(new_new_n931_), .D(new_new_n856_), .Y(zz04));
  INV        g1019(.A(new_new_n691_), .Y(new_new_n1044_));
  INV        g1020(.A(i_2_), .Y(new_new_n1045_));
  INV        g1021(.A(i_1_), .Y(new_new_n1046_));
  INV        g1022(.A(i_12_), .Y(new_new_n1047_));
  INV        g1023(.A(i_12_), .Y(new_new_n1048_));
endmodule


