//Benchmark atmr_alu4_1266_0.0625

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n971_, mai_mai_n972_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NA2        o032(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n55_));
  NO2        o033(.A(i_1_), .B(i_6_), .Y(ori_ori_n56_));
  NA2        o034(.A(i_8_), .B(i_7_), .Y(ori_ori_n57_));
  NAi21      o035(.An(i_2_), .B(i_7_), .Y(ori_ori_n58_));
  INV        o036(.A(i_1_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(i_6_), .Y(ori_ori_n60_));
  NA3        o038(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n31_), .Y(ori_ori_n61_));
  NA2        o039(.A(i_1_), .B(i_10_), .Y(ori_ori_n62_));
  NO2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NAi21      o041(.An(ori_ori_n63_), .B(ori_ori_n61_), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n65_));
  AOI210     o043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n66_));
  NA2        o044(.A(i_1_), .B(i_6_), .Y(ori_ori_n67_));
  NO2        o045(.A(ori_ori_n67_), .B(ori_ori_n25_), .Y(ori_ori_n68_));
  INV        o046(.A(i_0_), .Y(ori_ori_n69_));
  NAi21      o047(.An(i_5_), .B(i_10_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_5_), .B(i_9_), .Y(ori_ori_n71_));
  AOI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n70_), .B0(ori_ori_n69_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n72_), .B(ori_ori_n68_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n66_), .A1(ori_ori_n65_), .B0(ori_ori_n73_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n64_), .B0(i_0_), .Y(ori_ori_n75_));
  NA2        o053(.A(i_12_), .B(i_5_), .Y(ori_ori_n76_));
  NA2        o054(.A(i_2_), .B(i_8_), .Y(ori_ori_n77_));
  NO2        o055(.A(ori_ori_n77_), .B(ori_ori_n56_), .Y(ori_ori_n78_));
  NO2        o056(.A(i_3_), .B(i_9_), .Y(ori_ori_n79_));
  NO2        o057(.A(i_3_), .B(i_7_), .Y(ori_ori_n80_));
  INV        o058(.A(i_6_), .Y(ori_ori_n81_));
  OR4        o059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n82_));
  INV        o060(.A(ori_ori_n82_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_2_), .B(i_7_), .Y(ori_ori_n84_));
  NAi21      o062(.An(i_6_), .B(i_10_), .Y(ori_ori_n85_));
  NA2        o063(.A(i_6_), .B(i_9_), .Y(ori_ori_n86_));
  AOI210     o064(.A0(ori_ori_n86_), .A1(ori_ori_n85_), .B0(ori_ori_n59_), .Y(ori_ori_n87_));
  NA2        o065(.A(i_2_), .B(i_6_), .Y(ori_ori_n88_));
  NO3        o066(.A(ori_ori_n88_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n89_), .B(ori_ori_n87_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n874_), .B0(ori_ori_n76_), .Y(ori_ori_n91_));
  AN3        o069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n92_));
  NAi21      o070(.An(i_6_), .B(i_11_), .Y(ori_ori_n93_));
  NO2        o071(.A(i_5_), .B(i_8_), .Y(ori_ori_n94_));
  NOi21      o072(.An(ori_ori_n94_), .B(ori_ori_n93_), .Y(ori_ori_n95_));
  AOI220     o073(.A0(ori_ori_n95_), .A1(ori_ori_n58_), .B0(ori_ori_n92_), .B1(ori_ori_n32_), .Y(ori_ori_n96_));
  INV        o074(.A(i_7_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n46_), .B(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o076(.A(i_0_), .B(i_5_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n81_), .Y(ori_ori_n100_));
  NA2        o078(.A(i_12_), .B(i_3_), .Y(ori_ori_n101_));
  INV        o079(.A(ori_ori_n101_), .Y(ori_ori_n102_));
  NA3        o080(.A(ori_ori_n102_), .B(ori_ori_n100_), .C(ori_ori_n98_), .Y(ori_ori_n103_));
  NAi21      o081(.An(i_7_), .B(i_11_), .Y(ori_ori_n104_));
  NO3        o082(.A(ori_ori_n104_), .B(ori_ori_n85_), .C(ori_ori_n53_), .Y(ori_ori_n105_));
  AN2        o083(.A(i_2_), .B(i_10_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(i_7_), .Y(ori_ori_n107_));
  OR2        o085(.A(ori_ori_n76_), .B(ori_ori_n56_), .Y(ori_ori_n108_));
  NO2        o086(.A(i_8_), .B(ori_ori_n97_), .Y(ori_ori_n109_));
  NO3        o087(.A(ori_ori_n109_), .B(ori_ori_n108_), .C(ori_ori_n107_), .Y(ori_ori_n110_));
  NA2        o088(.A(i_12_), .B(i_7_), .Y(ori_ori_n111_));
  NO2        o089(.A(ori_ori_n59_), .B(ori_ori_n26_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(i_0_), .Y(ori_ori_n113_));
  NA2        o091(.A(i_11_), .B(i_12_), .Y(ori_ori_n114_));
  OAI210     o092(.A0(ori_ori_n113_), .A1(ori_ori_n111_), .B0(ori_ori_n114_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n115_), .B(ori_ori_n110_), .Y(ori_ori_n116_));
  NAi41      o094(.An(ori_ori_n105_), .B(ori_ori_n116_), .C(ori_ori_n103_), .D(ori_ori_n96_), .Y(ori_ori_n117_));
  NOi21      o095(.An(i_1_), .B(i_5_), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n118_), .B(i_11_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n97_), .B(ori_ori_n37_), .Y(ori_ori_n120_));
  NA2        o098(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n121_), .B(ori_ori_n120_), .Y(ori_ori_n122_));
  NO2        o100(.A(ori_ori_n122_), .B(ori_ori_n46_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n124_));
  NAi21      o102(.An(i_3_), .B(i_8_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(ori_ori_n58_), .Y(ori_ori_n126_));
  NOi31      o104(.An(ori_ori_n126_), .B(ori_ori_n124_), .C(ori_ori_n123_), .Y(ori_ori_n127_));
  NO2        o105(.A(i_1_), .B(ori_ori_n81_), .Y(ori_ori_n128_));
  NO2        o106(.A(i_6_), .B(i_5_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(i_3_), .Y(ori_ori_n130_));
  AO210      o108(.A0(ori_ori_n130_), .A1(ori_ori_n47_), .B0(ori_ori_n128_), .Y(ori_ori_n131_));
  OAI220     o109(.A0(ori_ori_n131_), .A1(ori_ori_n104_), .B0(ori_ori_n127_), .B1(ori_ori_n119_), .Y(ori_ori_n132_));
  NO3        o110(.A(ori_ori_n132_), .B(ori_ori_n117_), .C(ori_ori_n91_), .Y(ori_ori_n133_));
  NA3        o111(.A(ori_ori_n133_), .B(ori_ori_n75_), .C(ori_ori_n55_), .Y(ori2));
  NO2        o112(.A(ori_ori_n59_), .B(ori_ori_n37_), .Y(ori_ori_n135_));
  NA2        o113(.A(i_6_), .B(ori_ori_n25_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(ori_ori_n135_), .Y(ori_ori_n137_));
  NA4        o115(.A(ori_ori_n137_), .B(ori_ori_n73_), .C(ori_ori_n65_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o116(.A(i_8_), .B(i_7_), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n139_), .B(i_6_), .Y(ori_ori_n140_));
  NO2        o118(.A(i_12_), .B(i_13_), .Y(ori_ori_n141_));
  NAi21      o119(.An(i_5_), .B(i_11_), .Y(ori_ori_n142_));
  NOi21      o120(.An(ori_ori_n141_), .B(ori_ori_n142_), .Y(ori_ori_n143_));
  NO2        o121(.A(i_0_), .B(i_1_), .Y(ori_ori_n144_));
  NA2        o122(.A(i_2_), .B(i_3_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n145_), .B(i_4_), .Y(ori_ori_n146_));
  NA3        o124(.A(ori_ori_n146_), .B(ori_ori_n144_), .C(ori_ori_n143_), .Y(ori_ori_n147_));
  AN2        o125(.A(ori_ori_n141_), .B(ori_ori_n79_), .Y(ori_ori_n148_));
  NA2        o126(.A(i_1_), .B(i_5_), .Y(ori_ori_n149_));
  OR2        o127(.A(i_0_), .B(i_1_), .Y(ori_ori_n150_));
  NO3        o128(.A(ori_ori_n150_), .B(ori_ori_n76_), .C(i_13_), .Y(ori_ori_n151_));
  NAi32      o129(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n152_));
  NAi21      o130(.An(ori_ori_n152_), .B(ori_ori_n151_), .Y(ori_ori_n153_));
  NOi21      o131(.An(i_4_), .B(i_10_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n154_), .B(ori_ori_n40_), .Y(ori_ori_n155_));
  NO2        o133(.A(i_3_), .B(i_5_), .Y(ori_ori_n156_));
  NO3        o134(.A(ori_ori_n69_), .B(i_2_), .C(i_1_), .Y(ori_ori_n157_));
  NA2        o135(.A(ori_ori_n157_), .B(ori_ori_n156_), .Y(ori_ori_n158_));
  OAI210     o136(.A0(ori_ori_n158_), .A1(ori_ori_n155_), .B0(ori_ori_n153_), .Y(ori_ori_n159_));
  INV        o137(.A(ori_ori_n159_), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n160_), .B(ori_ori_n140_), .Y(ori_ori_n161_));
  NOi21      o139(.An(i_4_), .B(i_9_), .Y(ori_ori_n162_));
  NOi21      o140(.An(i_11_), .B(i_13_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n163_), .B(ori_ori_n162_), .Y(ori_ori_n164_));
  NO2        o142(.A(i_4_), .B(i_5_), .Y(ori_ori_n165_));
  NAi21      o143(.An(i_12_), .B(i_11_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n69_), .B(ori_ori_n59_), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n167_), .B(ori_ori_n46_), .Y(ori_ori_n168_));
  NA2        o146(.A(ori_ori_n36_), .B(i_5_), .Y(ori_ori_n169_));
  NAi31      o147(.An(ori_ori_n169_), .B(ori_ori_n148_), .C(i_11_), .Y(ori_ori_n170_));
  NA2        o148(.A(i_3_), .B(i_5_), .Y(ori_ori_n171_));
  OR2        o149(.A(ori_ori_n171_), .B(ori_ori_n164_), .Y(ori_ori_n172_));
  AOI210     o150(.A0(ori_ori_n172_), .A1(ori_ori_n170_), .B0(ori_ori_n168_), .Y(ori_ori_n173_));
  NO2        o151(.A(ori_ori_n69_), .B(i_5_), .Y(ori_ori_n174_));
  NO2        o152(.A(i_13_), .B(i_10_), .Y(ori_ori_n175_));
  NA3        o153(.A(ori_ori_n175_), .B(ori_ori_n174_), .C(ori_ori_n44_), .Y(ori_ori_n176_));
  NO2        o154(.A(i_2_), .B(i_1_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n177_), .B(i_3_), .Y(ori_ori_n178_));
  NAi21      o156(.An(i_4_), .B(i_12_), .Y(ori_ori_n179_));
  INV        o157(.A(ori_ori_n173_), .Y(ori_ori_n180_));
  INV        o158(.A(i_8_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n181_), .B(i_7_), .Y(ori_ori_n182_));
  NO3        o160(.A(i_3_), .B(ori_ori_n81_), .C(ori_ori_n48_), .Y(ori_ori_n183_));
  NA2        o161(.A(ori_ori_n183_), .B(ori_ori_n109_), .Y(ori_ori_n184_));
  NO3        o162(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n185_));
  NA3        o163(.A(ori_ori_n185_), .B(ori_ori_n40_), .C(ori_ori_n44_), .Y(ori_ori_n186_));
  NO3        o164(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n186_), .B(ori_ori_n184_), .Y(ori_ori_n188_));
  NO2        o166(.A(i_3_), .B(i_8_), .Y(ori_ori_n189_));
  NO3        o167(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n190_));
  NA3        o168(.A(ori_ori_n190_), .B(ori_ori_n189_), .C(ori_ori_n40_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n99_), .B(ori_ori_n56_), .Y(ori_ori_n192_));
  INV        o170(.A(ori_ori_n192_), .Y(ori_ori_n193_));
  NO2        o171(.A(i_13_), .B(i_9_), .Y(ori_ori_n194_));
  NAi21      o172(.An(i_12_), .B(i_3_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n193_), .B(ori_ori_n191_), .Y(ori_ori_n197_));
  AOI210     o175(.A0(ori_ori_n197_), .A1(i_7_), .B0(ori_ori_n188_), .Y(ori_ori_n198_));
  OAI220     o176(.A0(ori_ori_n198_), .A1(i_4_), .B0(i_7_), .B1(ori_ori_n180_), .Y(ori_ori_n199_));
  NAi21      o177(.An(i_12_), .B(i_7_), .Y(ori_ori_n200_));
  NA3        o178(.A(i_13_), .B(ori_ori_n181_), .C(i_10_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n200_), .Y(ori_ori_n202_));
  NA2        o180(.A(i_0_), .B(i_5_), .Y(ori_ori_n203_));
  OAI220     o181(.A0(ori_ori_n81_), .A1(ori_ori_n178_), .B0(ori_ori_n168_), .B1(ori_ori_n130_), .Y(ori_ori_n204_));
  NAi31      o182(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n46_), .B(ori_ori_n59_), .Y(ori_ori_n207_));
  NA3        o185(.A(ori_ori_n207_), .B(i_0_), .C(ori_ori_n206_), .Y(ori_ori_n208_));
  INV        o186(.A(i_13_), .Y(ori_ori_n209_));
  NO2        o187(.A(i_12_), .B(ori_ori_n209_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n208_), .B(ori_ori_n205_), .Y(ori_ori_n211_));
  AOI220     o189(.A0(ori_ori_n211_), .A1(ori_ori_n139_), .B0(ori_ori_n204_), .B1(ori_ori_n202_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n213_));
  OR2        o191(.A(i_8_), .B(i_7_), .Y(ori_ori_n214_));
  NO2        o192(.A(ori_ori_n53_), .B(i_1_), .Y(ori_ori_n215_));
  INV        o193(.A(i_12_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n44_), .B(ori_ori_n216_), .Y(ori_ori_n217_));
  NO3        o195(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n218_));
  NA2        o196(.A(i_2_), .B(i_1_), .Y(ori_ori_n219_));
  NO3        o197(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n220_));
  NAi21      o198(.An(i_4_), .B(i_3_), .Y(ori_ori_n221_));
  NO2        o199(.A(i_0_), .B(i_6_), .Y(ori_ori_n222_));
  NOi41      o200(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n219_), .B(ori_ori_n171_), .Y(ori_ori_n224_));
  NO2        o202(.A(i_11_), .B(ori_ori_n209_), .Y(ori_ori_n225_));
  NOi21      o203(.An(i_1_), .B(i_6_), .Y(ori_ori_n226_));
  NAi21      o204(.An(i_3_), .B(i_7_), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n216_), .B(i_9_), .Y(ori_ori_n228_));
  OR4        o206(.A(ori_ori_n228_), .B(ori_ori_n227_), .C(ori_ori_n226_), .D(ori_ori_n174_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_12_), .B(i_3_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n69_), .B(i_5_), .Y(ori_ori_n231_));
  NA2        o209(.A(i_3_), .B(i_9_), .Y(ori_ori_n232_));
  NAi21      o210(.An(i_7_), .B(i_10_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n233_), .B(ori_ori_n232_), .Y(ori_ori_n234_));
  NA3        o212(.A(ori_ori_n234_), .B(ori_ori_n231_), .C(ori_ori_n60_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n235_), .B(ori_ori_n229_), .Y(ori_ori_n236_));
  INV        o214(.A(ori_ori_n140_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n216_), .B(i_13_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n238_), .B(ori_ori_n71_), .Y(ori_ori_n239_));
  AOI220     o217(.A0(ori_ori_n239_), .A1(ori_ori_n237_), .B0(ori_ori_n236_), .B1(ori_ori_n225_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n214_), .B(ori_ori_n37_), .Y(ori_ori_n241_));
  NA2        o219(.A(i_12_), .B(i_6_), .Y(ori_ori_n242_));
  OR2        o220(.A(i_13_), .B(i_9_), .Y(ori_ori_n243_));
  NO3        o221(.A(ori_ori_n243_), .B(ori_ori_n242_), .C(ori_ori_n48_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n221_), .B(i_2_), .Y(ori_ori_n245_));
  NA3        o223(.A(ori_ori_n245_), .B(ori_ori_n244_), .C(ori_ori_n44_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n225_), .B(i_9_), .Y(ori_ori_n247_));
  NA2        o225(.A(ori_ori_n231_), .B(ori_ori_n60_), .Y(ori_ori_n248_));
  OAI210     o226(.A0(ori_ori_n248_), .A1(ori_ori_n247_), .B0(ori_ori_n246_), .Y(ori_ori_n249_));
  NO3        o227(.A(i_11_), .B(ori_ori_n209_), .C(ori_ori_n25_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n227_), .B(i_8_), .Y(ori_ori_n251_));
  NA2        o229(.A(ori_ori_n249_), .B(ori_ori_n241_), .Y(ori_ori_n252_));
  NA3        o230(.A(ori_ori_n252_), .B(ori_ori_n240_), .C(ori_ori_n212_), .Y(ori_ori_n253_));
  NO3        o231(.A(i_12_), .B(ori_ori_n209_), .C(ori_ori_n37_), .Y(ori_ori_n254_));
  INV        o232(.A(ori_ori_n254_), .Y(ori_ori_n255_));
  NA2        o233(.A(i_8_), .B(ori_ori_n97_), .Y(ori_ori_n256_));
  AOI220     o234(.A0(i_2_), .A1(ori_ori_n183_), .B0(ori_ori_n156_), .B1(ori_ori_n215_), .Y(ori_ori_n257_));
  NO2        o235(.A(ori_ori_n257_), .B(ori_ori_n256_), .Y(ori_ori_n258_));
  NO3        o236(.A(i_0_), .B(i_2_), .C(ori_ori_n59_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n219_), .B(i_0_), .Y(ori_ori_n260_));
  AOI220     o238(.A0(ori_ori_n260_), .A1(ori_ori_n182_), .B0(ori_ori_n259_), .B1(ori_ori_n139_), .Y(ori_ori_n261_));
  NA2        o239(.A(i_5_), .B(ori_ori_n26_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n261_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n57_), .B(i_6_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n158_), .B(ori_ori_n140_), .Y(ori_ori_n265_));
  NO3        o243(.A(ori_ori_n265_), .B(ori_ori_n263_), .C(ori_ori_n258_), .Y(ori_ori_n266_));
  NO2        o244(.A(i_3_), .B(i_10_), .Y(ori_ori_n267_));
  NO2        o245(.A(i_2_), .B(ori_ori_n97_), .Y(ori_ori_n268_));
  AN2        o246(.A(i_3_), .B(i_10_), .Y(ori_ori_n269_));
  NO2        o247(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n266_), .B(ori_ori_n255_), .Y(ori_ori_n272_));
  NO4        o250(.A(ori_ori_n272_), .B(ori_ori_n253_), .C(ori_ori_n199_), .D(ori_ori_n161_), .Y(ori_ori_n273_));
  NO3        o251(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n260_), .B(i_7_), .Y(ori_ori_n275_));
  NO3        o253(.A(i_6_), .B(ori_ori_n181_), .C(i_7_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n276_), .B(ori_ori_n185_), .Y(ori_ori_n277_));
  AOI210     o255(.A0(ori_ori_n277_), .A1(ori_ori_n275_), .B0(i_5_), .Y(ori_ori_n278_));
  NO2        o256(.A(i_2_), .B(i_3_), .Y(ori_ori_n279_));
  OR2        o257(.A(i_0_), .B(i_5_), .Y(ori_ori_n280_));
  NA3        o258(.A(ori_ori_n260_), .B(ori_ori_n156_), .C(ori_ori_n109_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n150_), .B(ori_ori_n46_), .Y(ori_ori_n282_));
  INV        o260(.A(ori_ori_n281_), .Y(ori_ori_n283_));
  OAI210     o261(.A0(ori_ori_n283_), .A1(ori_ori_n278_), .B0(i_4_), .Y(ori_ori_n284_));
  NO2        o262(.A(i_12_), .B(i_10_), .Y(ori_ori_n285_));
  NOi21      o263(.An(i_5_), .B(i_0_), .Y(ori_ori_n286_));
  NO2        o264(.A(i_2_), .B(ori_ori_n97_), .Y(ori_ori_n287_));
  NO4        o265(.A(ori_ori_n287_), .B(i_4_), .C(ori_ori_n286_), .D(ori_ori_n125_), .Y(ori_ori_n288_));
  NA4        o266(.A(ori_ori_n80_), .B(ori_ori_n36_), .C(ori_ori_n81_), .D(i_8_), .Y(ori_ori_n289_));
  NA2        o267(.A(ori_ori_n288_), .B(ori_ori_n285_), .Y(ori_ori_n290_));
  NO2        o268(.A(i_6_), .B(i_8_), .Y(ori_ori_n291_));
  NOi21      o269(.An(i_0_), .B(i_2_), .Y(ori_ori_n292_));
  AN2        o270(.A(ori_ori_n292_), .B(ori_ori_n291_), .Y(ori_ori_n293_));
  NO2        o271(.A(i_1_), .B(i_7_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n290_), .B(ori_ori_n284_), .Y(ori_ori_n295_));
  NA3        o273(.A(ori_ori_n226_), .B(ori_ori_n268_), .C(ori_ori_n181_), .Y(ori_ori_n296_));
  INV        o274(.A(ori_ori_n88_), .Y(ori_ori_n297_));
  NO2        o275(.A(ori_ori_n181_), .B(i_9_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n298_), .B(ori_ori_n192_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n299_), .B(ori_ori_n46_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n300_), .B(ori_ori_n263_), .Y(ori_ori_n301_));
  AOI210     o279(.A0(ori_ori_n301_), .A1(ori_ori_n296_), .B0(ori_ori_n155_), .Y(ori_ori_n302_));
  AOI210     o280(.A0(ori_ori_n295_), .A1(ori_ori_n274_), .B0(ori_ori_n302_), .Y(ori_ori_n303_));
  NOi32      o281(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n304_));
  INV        o282(.A(ori_ori_n304_), .Y(ori_ori_n305_));
  NAi21      o283(.An(i_0_), .B(i_6_), .Y(ori_ori_n306_));
  NAi21      o284(.An(i_1_), .B(i_5_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n307_), .B(ori_ori_n306_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n308_), .B(ori_ori_n25_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n309_), .B(ori_ori_n152_), .Y(ori_ori_n310_));
  NO2        o288(.A(ori_ori_n152_), .B(ori_ori_n150_), .Y(ori_ori_n311_));
  NOi32      o289(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n312_));
  NAi21      o290(.An(i_6_), .B(i_1_), .Y(ori_ori_n313_));
  NA3        o291(.A(ori_ori_n313_), .B(ori_ori_n312_), .C(ori_ori_n46_), .Y(ori_ori_n314_));
  NO2        o292(.A(ori_ori_n314_), .B(i_0_), .Y(ori_ori_n315_));
  OR2        o293(.A(ori_ori_n315_), .B(ori_ori_n311_), .Y(ori_ori_n316_));
  NO2        o294(.A(i_1_), .B(ori_ori_n97_), .Y(ori_ori_n317_));
  NAi21      o295(.An(i_3_), .B(i_4_), .Y(ori_ori_n318_));
  NO2        o296(.A(ori_ori_n318_), .B(i_9_), .Y(ori_ori_n319_));
  AN2        o297(.A(i_6_), .B(i_7_), .Y(ori_ori_n320_));
  OAI210     o298(.A0(ori_ori_n320_), .A1(ori_ori_n317_), .B0(ori_ori_n319_), .Y(ori_ori_n321_));
  NA2        o299(.A(i_2_), .B(i_7_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n318_), .B(i_10_), .Y(ori_ori_n323_));
  NA3        o301(.A(ori_ori_n323_), .B(ori_ori_n322_), .C(ori_ori_n222_), .Y(ori_ori_n324_));
  AOI210     o302(.A0(ori_ori_n324_), .A1(ori_ori_n321_), .B0(ori_ori_n174_), .Y(ori_ori_n325_));
  AOI210     o303(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n326_));
  AOI220     o304(.A0(ori_ori_n323_), .A1(ori_ori_n294_), .B0(ori_ori_n218_), .B1(ori_ori_n177_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n327_), .B(i_5_), .Y(ori_ori_n328_));
  NO4        o306(.A(ori_ori_n328_), .B(ori_ori_n325_), .C(ori_ori_n316_), .D(ori_ori_n310_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n329_), .B(ori_ori_n305_), .Y(ori_ori_n330_));
  NO2        o308(.A(ori_ori_n57_), .B(ori_ori_n25_), .Y(ori_ori_n331_));
  AN2        o309(.A(i_12_), .B(i_5_), .Y(ori_ori_n332_));
  NO2        o310(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n333_));
  NA2        o311(.A(ori_ori_n333_), .B(ori_ori_n332_), .Y(ori_ori_n334_));
  NO2        o312(.A(i_11_), .B(i_6_), .Y(ori_ori_n335_));
  NA3        o313(.A(ori_ori_n335_), .B(ori_ori_n282_), .C(ori_ori_n209_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n336_), .B(ori_ori_n334_), .Y(ori_ori_n337_));
  NO2        o315(.A(ori_ori_n221_), .B(i_5_), .Y(ori_ori_n338_));
  NO2        o316(.A(i_5_), .B(i_10_), .Y(ori_ori_n339_));
  AOI220     o317(.A0(ori_ori_n339_), .A1(ori_ori_n245_), .B0(ori_ori_n338_), .B1(ori_ori_n185_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n141_), .B(ori_ori_n45_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n340_), .Y(ori_ori_n342_));
  OAI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n337_), .B0(ori_ori_n331_), .Y(ori_ori_n343_));
  NO2        o321(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n344_));
  NO2        o322(.A(ori_ori_n147_), .B(ori_ori_n81_), .Y(ori_ori_n345_));
  OAI210     o323(.A0(ori_ori_n345_), .A1(ori_ori_n337_), .B0(ori_ori_n344_), .Y(ori_ori_n346_));
  NO3        o324(.A(ori_ori_n81_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n347_));
  NA3        o325(.A(ori_ori_n267_), .B(ori_ori_n86_), .C(ori_ori_n71_), .Y(ori_ori_n348_));
  NO2        o326(.A(i_11_), .B(i_12_), .Y(ori_ori_n349_));
  NA2        o327(.A(ori_ori_n349_), .B(ori_ori_n36_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n348_), .B(ori_ori_n350_), .Y(ori_ori_n351_));
  NA2        o329(.A(ori_ori_n339_), .B(ori_ori_n216_), .Y(ori_ori_n352_));
  NAi21      o330(.An(i_13_), .B(i_0_), .Y(ori_ori_n353_));
  NO2        o331(.A(ori_ori_n353_), .B(ori_ori_n219_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n351_), .B(ori_ori_n354_), .Y(ori_ori_n355_));
  NA3        o333(.A(ori_ori_n355_), .B(ori_ori_n346_), .C(ori_ori_n343_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n44_), .B(ori_ori_n209_), .Y(ori_ori_n357_));
  NO2        o335(.A(i_0_), .B(i_11_), .Y(ori_ori_n358_));
  AN2        o336(.A(i_1_), .B(i_6_), .Y(ori_ori_n359_));
  NOi21      o337(.An(i_2_), .B(i_12_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n139_), .B(i_9_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n361_), .B(i_4_), .Y(ori_ori_n362_));
  OR2        o340(.A(i_13_), .B(i_10_), .Y(ori_ori_n363_));
  NO2        o341(.A(ori_ori_n164_), .B(ori_ori_n120_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n97_), .B(ori_ori_n25_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n171_), .B(ori_ori_n81_), .Y(ori_ori_n366_));
  NA2        o344(.A(ori_ori_n181_), .B(i_10_), .Y(ori_ori_n367_));
  NA3        o345(.A(ori_ori_n231_), .B(ori_ori_n60_), .C(i_2_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n264_), .B(ori_ori_n215_), .Y(ori_ori_n369_));
  OAI220     o347(.A0(ori_ori_n369_), .A1(ori_ori_n171_), .B0(ori_ori_n368_), .B1(ori_ori_n367_), .Y(ori_ori_n370_));
  INV        o348(.A(ori_ori_n370_), .Y(ori_ori_n371_));
  AOI210     o349(.A0(ori_ori_n371_), .A1(ori_ori_n281_), .B0(ori_ori_n247_), .Y(ori_ori_n372_));
  NO3        o350(.A(ori_ori_n372_), .B(ori_ori_n356_), .C(ori_ori_n330_), .Y(ori_ori_n373_));
  NO2        o351(.A(ori_ori_n69_), .B(i_13_), .Y(ori_ori_n374_));
  NO2        o352(.A(i_10_), .B(i_9_), .Y(ori_ori_n375_));
  NAi21      o353(.An(i_12_), .B(i_8_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n376_), .B(i_3_), .Y(ori_ori_n377_));
  NO2        o355(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n378_));
  NA2        o356(.A(ori_ori_n378_), .B(ori_ori_n100_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n379_), .B(ori_ori_n191_), .Y(ori_ori_n380_));
  NA2        o358(.A(ori_ori_n271_), .B(i_0_), .Y(ori_ori_n381_));
  NO3        o359(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n242_), .B(ori_ori_n93_), .Y(ori_ori_n383_));
  NA2        o361(.A(ori_ori_n383_), .B(ori_ori_n382_), .Y(ori_ori_n384_));
  NA2        o362(.A(i_8_), .B(i_9_), .Y(ori_ori_n385_));
  AOI210     o363(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n386_));
  OR2        o364(.A(ori_ori_n386_), .B(ori_ori_n385_), .Y(ori_ori_n387_));
  NA2        o365(.A(ori_ori_n254_), .B(ori_ori_n192_), .Y(ori_ori_n388_));
  OAI220     o366(.A0(ori_ori_n388_), .A1(ori_ori_n387_), .B0(ori_ori_n384_), .B1(ori_ori_n381_), .Y(ori_ori_n389_));
  NO3        o367(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n389_), .B(ori_ori_n380_), .Y(ori_ori_n391_));
  OR2        o369(.A(ori_ori_n299_), .B(ori_ori_n97_), .Y(ori_ori_n392_));
  OR2        o370(.A(ori_ori_n392_), .B(ori_ori_n155_), .Y(ori_ori_n393_));
  NA2        o371(.A(ori_ori_n92_), .B(i_13_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n366_), .B(ori_ori_n331_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n395_), .B(ori_ori_n394_), .Y(ori_ori_n396_));
  NO3        o374(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n397_));
  NO2        o375(.A(i_6_), .B(i_7_), .Y(ori_ori_n398_));
  NO2        o376(.A(i_11_), .B(i_1_), .Y(ori_ori_n399_));
  OR2        o377(.A(i_11_), .B(i_8_), .Y(ori_ori_n400_));
  NOi21      o378(.An(i_2_), .B(i_7_), .Y(ori_ori_n401_));
  NO2        o379(.A(i_6_), .B(i_10_), .Y(ori_ori_n402_));
  NA3        o380(.A(ori_ori_n223_), .B(ori_ori_n163_), .C(ori_ori_n129_), .Y(ori_ori_n403_));
  NA2        o381(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n404_));
  NA3        o382(.A(ori_ori_n344_), .B(ori_ori_n167_), .C(ori_ori_n146_), .Y(ori_ori_n405_));
  NA2        o383(.A(ori_ori_n405_), .B(ori_ori_n403_), .Y(ori_ori_n406_));
  NO2        o384(.A(ori_ori_n406_), .B(ori_ori_n396_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n382_), .B(ori_ori_n332_), .Y(ori_ori_n408_));
  NA2        o386(.A(ori_ori_n390_), .B(ori_ori_n339_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n409_), .B(ori_ori_n208_), .Y(ori_ori_n410_));
  NAi21      o388(.An(ori_ori_n201_), .B(ori_ori_n349_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n294_), .B(ori_ori_n203_), .Y(ori_ori_n412_));
  NO2        o390(.A(ori_ori_n412_), .B(ori_ori_n411_), .Y(ori_ori_n413_));
  NA2        o391(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n274_), .B(ori_ori_n218_), .Y(ori_ori_n415_));
  OAI220     o393(.A0(ori_ori_n415_), .A1(ori_ori_n368_), .B0(ori_ori_n414_), .B1(ori_ori_n394_), .Y(ori_ori_n416_));
  NO3        o394(.A(ori_ori_n416_), .B(ori_ori_n413_), .C(ori_ori_n410_), .Y(ori_ori_n417_));
  NA4        o395(.A(ori_ori_n417_), .B(ori_ori_n407_), .C(ori_ori_n393_), .D(ori_ori_n391_), .Y(ori_ori_n418_));
  NA2        o396(.A(ori_ori_n119_), .B(ori_ori_n108_), .Y(ori_ori_n419_));
  AN2        o397(.A(ori_ori_n419_), .B(ori_ori_n382_), .Y(ori_ori_n420_));
  NA2        o398(.A(ori_ori_n420_), .B(ori_ori_n271_), .Y(ori_ori_n421_));
  NA2        o399(.A(ori_ori_n304_), .B(ori_ori_n69_), .Y(ori_ori_n422_));
  NA2        o400(.A(ori_ori_n320_), .B(ori_ori_n312_), .Y(ori_ori_n423_));
  NO2        o401(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n424_));
  NA2        o402(.A(ori_ori_n39_), .B(i_13_), .Y(ori_ori_n425_));
  OAI210     o403(.A0(i_8_), .A1(ori_ori_n59_), .B0(ori_ori_n131_), .Y(ori_ori_n426_));
  NA2        o404(.A(ori_ori_n426_), .B(ori_ori_n364_), .Y(ori_ori_n427_));
  NA3        o405(.A(ori_ori_n427_), .B(ori_ori_n425_), .C(ori_ori_n421_), .Y(ori_ori_n428_));
  NO2        o406(.A(i_12_), .B(ori_ori_n181_), .Y(ori_ori_n429_));
  NO2        o407(.A(i_8_), .B(i_7_), .Y(ori_ori_n430_));
  OAI210     o408(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n431_), .B(ori_ori_n207_), .Y(ori_ori_n432_));
  NO2        o410(.A(ori_ori_n432_), .B(ori_ori_n221_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n434_));
  NO2        o412(.A(ori_ori_n434_), .B(i_6_), .Y(ori_ori_n435_));
  NA3        o413(.A(ori_ori_n435_), .B(ori_ori_n433_), .C(ori_ori_n430_), .Y(ori_ori_n436_));
  AOI220     o414(.A0(ori_ori_n366_), .A1(ori_ori_n282_), .B0(ori_ori_n224_), .B1(ori_ori_n222_), .Y(ori_ori_n437_));
  OAI220     o415(.A0(ori_ori_n437_), .A1(ori_ori_n238_), .B0(ori_ori_n394_), .B1(ori_ori_n130_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n438_), .B(ori_ori_n241_), .Y(ori_ori_n439_));
  NA3        o417(.A(ori_ori_n269_), .B(ori_ori_n165_), .C(ori_ori_n92_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n206_), .B(ori_ori_n44_), .Y(ori_ori_n441_));
  NO2        o419(.A(ori_ori_n150_), .B(i_5_), .Y(ori_ori_n442_));
  NA3        o420(.A(ori_ori_n442_), .B(ori_ori_n357_), .C(ori_ori_n279_), .Y(ori_ori_n443_));
  OAI210     o421(.A0(ori_ori_n443_), .A1(ori_ori_n441_), .B0(ori_ori_n440_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n444_), .B(ori_ori_n390_), .Y(ori_ori_n445_));
  NA3        o423(.A(ori_ori_n445_), .B(ori_ori_n439_), .C(ori_ori_n436_), .Y(ori_ori_n446_));
  AOI210     o424(.A0(ori_ori_n313_), .A1(ori_ori_n46_), .B0(ori_ori_n317_), .Y(ori_ori_n447_));
  NA2        o425(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n448_));
  NA3        o426(.A(ori_ori_n429_), .B(ori_ori_n250_), .C(ori_ori_n448_), .Y(ori_ori_n449_));
  NO2        o427(.A(ori_ori_n447_), .B(ori_ori_n449_), .Y(ori_ori_n450_));
  INV        o428(.A(ori_ori_n450_), .Y(ori_ori_n451_));
  NO4        o429(.A(ori_ori_n226_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n452_));
  NO3        o430(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n453_));
  NO2        o431(.A(ori_ori_n214_), .B(ori_ori_n36_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n363_), .B(i_1_), .Y(ori_ori_n455_));
  NOi31      o433(.An(ori_ori_n455_), .B(ori_ori_n383_), .C(ori_ori_n69_), .Y(ori_ori_n456_));
  AN4        o434(.A(ori_ori_n456_), .B(ori_ori_n362_), .C(i_3_), .D(i_2_), .Y(ori_ori_n457_));
  INV        o435(.A(ori_ori_n457_), .Y(ori_ori_n458_));
  NOi21      o436(.An(i_10_), .B(i_6_), .Y(ori_ori_n459_));
  NO2        o437(.A(ori_ori_n81_), .B(ori_ori_n25_), .Y(ori_ori_n460_));
  AOI220     o438(.A0(ori_ori_n254_), .A1(ori_ori_n460_), .B0(ori_ori_n250_), .B1(ori_ori_n459_), .Y(ori_ori_n461_));
  NO2        o439(.A(ori_ori_n461_), .B(ori_ori_n381_), .Y(ori_ori_n462_));
  NO2        o440(.A(ori_ori_n111_), .B(ori_ori_n23_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n276_), .B(ori_ori_n157_), .Y(ori_ori_n464_));
  AOI220     o442(.A0(ori_ori_n464_), .A1(ori_ori_n369_), .B0(ori_ori_n172_), .B1(ori_ori_n170_), .Y(ori_ori_n465_));
  NO2        o443(.A(ori_ori_n185_), .B(ori_ori_n37_), .Y(ori_ori_n466_));
  NOi31      o444(.An(ori_ori_n143_), .B(ori_ori_n466_), .C(ori_ori_n289_), .Y(ori_ori_n467_));
  NO3        o445(.A(ori_ori_n467_), .B(ori_ori_n465_), .C(ori_ori_n462_), .Y(ori_ori_n468_));
  NO2        o446(.A(ori_ori_n422_), .B(ori_ori_n327_), .Y(ori_ori_n469_));
  INV        o447(.A(ori_ori_n279_), .Y(ori_ori_n470_));
  NO2        o448(.A(i_12_), .B(ori_ori_n81_), .Y(ori_ori_n471_));
  NA3        o449(.A(ori_ori_n471_), .B(ori_ori_n250_), .C(ori_ori_n448_), .Y(ori_ori_n472_));
  NA3        o450(.A(ori_ori_n335_), .B(ori_ori_n254_), .C(ori_ori_n203_), .Y(ori_ori_n473_));
  AOI210     o451(.A0(ori_ori_n473_), .A1(ori_ori_n472_), .B0(ori_ori_n470_), .Y(ori_ori_n474_));
  OR2        o452(.A(i_2_), .B(i_5_), .Y(ori_ori_n475_));
  OR2        o453(.A(ori_ori_n475_), .B(ori_ori_n359_), .Y(ori_ori_n476_));
  NA2        o454(.A(ori_ori_n322_), .B(ori_ori_n222_), .Y(ori_ori_n477_));
  AOI210     o455(.A0(ori_ori_n477_), .A1(ori_ori_n476_), .B0(ori_ori_n411_), .Y(ori_ori_n478_));
  NO3        o456(.A(ori_ori_n478_), .B(ori_ori_n474_), .C(ori_ori_n469_), .Y(ori_ori_n479_));
  NA4        o457(.A(ori_ori_n479_), .B(ori_ori_n468_), .C(ori_ori_n458_), .D(ori_ori_n451_), .Y(ori_ori_n480_));
  NO4        o458(.A(ori_ori_n480_), .B(ori_ori_n446_), .C(ori_ori_n428_), .D(ori_ori_n418_), .Y(ori_ori_n481_));
  NA4        o459(.A(ori_ori_n481_), .B(ori_ori_n373_), .C(ori_ori_n303_), .D(ori_ori_n273_), .Y(ori7));
  NO2        o460(.A(ori_ori_n88_), .B(ori_ori_n54_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n104_), .B(ori_ori_n85_), .Y(ori_ori_n484_));
  NA2        o462(.A(ori_ori_n333_), .B(ori_ori_n484_), .Y(ori_ori_n485_));
  NA2        o463(.A(ori_ori_n402_), .B(ori_ori_n80_), .Y(ori_ori_n486_));
  NA2        o464(.A(i_11_), .B(ori_ori_n181_), .Y(ori_ori_n487_));
  NA2        o465(.A(ori_ori_n141_), .B(ori_ori_n487_), .Y(ori_ori_n488_));
  OAI210     o466(.A0(ori_ori_n488_), .A1(ori_ori_n486_), .B0(ori_ori_n485_), .Y(ori_ori_n489_));
  NO2        o467(.A(ori_ori_n216_), .B(i_4_), .Y(ori_ori_n490_));
  NA2        o468(.A(ori_ori_n490_), .B(i_8_), .Y(ori_ori_n491_));
  NA2        o469(.A(i_2_), .B(ori_ori_n81_), .Y(ori_ori_n492_));
  OAI210     o470(.A0(ori_ori_n84_), .A1(ori_ori_n189_), .B0(ori_ori_n190_), .Y(ori_ori_n493_));
  NO2        o471(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n494_));
  NA2        o472(.A(i_4_), .B(i_8_), .Y(ori_ori_n495_));
  AOI210     o473(.A0(ori_ori_n495_), .A1(ori_ori_n269_), .B0(ori_ori_n494_), .Y(ori_ori_n496_));
  OAI220     o474(.A0(ori_ori_n496_), .A1(ori_ori_n492_), .B0(ori_ori_n493_), .B1(i_13_), .Y(ori_ori_n497_));
  NO3        o475(.A(ori_ori_n497_), .B(ori_ori_n489_), .C(ori_ori_n483_), .Y(ori_ori_n498_));
  AOI210     o476(.A0(ori_ori_n125_), .A1(ori_ori_n58_), .B0(i_10_), .Y(ori_ori_n499_));
  AOI210     o477(.A0(ori_ori_n499_), .A1(ori_ori_n216_), .B0(ori_ori_n154_), .Y(ori_ori_n500_));
  OR2        o478(.A(i_6_), .B(i_10_), .Y(ori_ori_n501_));
  OR3        o479(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n502_));
  INV        o480(.A(ori_ori_n187_), .Y(ori_ori_n503_));
  OR2        o481(.A(ori_ori_n500_), .B(ori_ori_n243_), .Y(ori_ori_n504_));
  AOI210     o482(.A0(ori_ori_n504_), .A1(ori_ori_n498_), .B0(ori_ori_n59_), .Y(ori_ori_n505_));
  NOi21      o483(.An(i_11_), .B(i_7_), .Y(ori_ori_n506_));
  AO210      o484(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n507_));
  NO2        o485(.A(ori_ori_n507_), .B(ori_ori_n506_), .Y(ori_ori_n508_));
  NA2        o486(.A(ori_ori_n508_), .B(ori_ori_n194_), .Y(ori_ori_n509_));
  NA3        o487(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n510_));
  NAi31      o488(.An(ori_ori_n510_), .B(ori_ori_n200_), .C(i_11_), .Y(ori_ori_n511_));
  AOI210     o489(.A0(ori_ori_n511_), .A1(ori_ori_n509_), .B0(ori_ori_n59_), .Y(ori_ori_n512_));
  NA2        o490(.A(ori_ori_n83_), .B(ori_ori_n59_), .Y(ori_ori_n513_));
  AO210      o491(.A0(ori_ori_n513_), .A1(ori_ori_n327_), .B0(ori_ori_n41_), .Y(ori_ori_n514_));
  NO3        o492(.A(ori_ori_n233_), .B(ori_ori_n195_), .C(ori_ori_n487_), .Y(ori_ori_n515_));
  OAI210     o493(.A0(ori_ori_n515_), .A1(ori_ori_n210_), .B0(ori_ori_n59_), .Y(ori_ori_n516_));
  NA2        o494(.A(ori_ori_n360_), .B(ori_ori_n31_), .Y(ori_ori_n517_));
  OR2        o495(.A(ori_ori_n195_), .B(ori_ori_n104_), .Y(ori_ori_n518_));
  NA2        o496(.A(ori_ori_n518_), .B(ori_ori_n517_), .Y(ori_ori_n519_));
  NO2        o497(.A(i_1_), .B(i_4_), .Y(ori_ori_n520_));
  NA2        o498(.A(ori_ori_n520_), .B(ori_ori_n519_), .Y(ori_ori_n521_));
  NO2        o499(.A(i_1_), .B(i_12_), .Y(ori_ori_n522_));
  NA3        o500(.A(ori_ori_n521_), .B(ori_ori_n516_), .C(ori_ori_n514_), .Y(ori_ori_n523_));
  OAI210     o501(.A0(ori_ori_n523_), .A1(ori_ori_n512_), .B0(i_6_), .Y(ori_ori_n524_));
  NO2        o502(.A(ori_ori_n510_), .B(ori_ori_n104_), .Y(ori_ori_n525_));
  NA2        o503(.A(ori_ori_n525_), .B(ori_ori_n471_), .Y(ori_ori_n526_));
  NO2        o504(.A(i_6_), .B(i_11_), .Y(ori_ori_n527_));
  NA2        o505(.A(ori_ori_n526_), .B(ori_ori_n384_), .Y(ori_ori_n528_));
  NO3        o506(.A(ori_ori_n501_), .B(ori_ori_n214_), .C(ori_ori_n23_), .Y(ori_ori_n529_));
  AOI210     o507(.A0(i_1_), .A1(ori_ori_n234_), .B0(ori_ori_n529_), .Y(ori_ori_n530_));
  NO2        o508(.A(ori_ori_n530_), .B(ori_ori_n44_), .Y(ori_ori_n531_));
  NA3        o509(.A(ori_ori_n430_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n532_));
  INV        o510(.A(i_2_), .Y(ori_ori_n533_));
  NA2        o511(.A(ori_ori_n135_), .B(i_9_), .Y(ori_ori_n534_));
  NO2        o512(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n535_));
  NO2        o513(.A(ori_ori_n534_), .B(ori_ori_n533_), .Y(ori_ori_n536_));
  AOI210     o514(.A0(ori_ori_n399_), .A1(ori_ori_n365_), .B0(ori_ori_n220_), .Y(ori_ori_n537_));
  NO2        o515(.A(ori_ori_n537_), .B(ori_ori_n492_), .Y(ori_ori_n538_));
  NAi21      o516(.An(ori_ori_n532_), .B(ori_ori_n87_), .Y(ori_ori_n539_));
  NA2        o517(.A(ori_ori_n535_), .B(ori_ori_n242_), .Y(ori_ori_n540_));
  NO2        o518(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n541_));
  NA2        o519(.A(ori_ori_n541_), .B(ori_ori_n24_), .Y(ori_ori_n542_));
  OAI210     o520(.A0(ori_ori_n542_), .A1(ori_ori_n540_), .B0(ori_ori_n539_), .Y(ori_ori_n543_));
  OR3        o521(.A(ori_ori_n543_), .B(ori_ori_n538_), .C(ori_ori_n536_), .Y(ori_ori_n544_));
  NO3        o522(.A(ori_ori_n544_), .B(ori_ori_n531_), .C(ori_ori_n528_), .Y(ori_ori_n545_));
  NO2        o523(.A(ori_ori_n216_), .B(ori_ori_n97_), .Y(ori_ori_n546_));
  NO2        o524(.A(ori_ori_n546_), .B(ori_ori_n506_), .Y(ori_ori_n547_));
  NA2        o525(.A(ori_ori_n547_), .B(i_1_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n548_), .B(ori_ori_n502_), .Y(ori_ori_n549_));
  NA2        o527(.A(ori_ori_n549_), .B(ori_ori_n46_), .Y(ori_ori_n550_));
  NA2        o528(.A(i_3_), .B(ori_ori_n181_), .Y(ori_ori_n551_));
  NO2        o529(.A(ori_ori_n551_), .B(ori_ori_n111_), .Y(ori_ori_n552_));
  AN2        o530(.A(ori_ori_n552_), .B(ori_ori_n435_), .Y(ori_ori_n553_));
  NO2        o531(.A(ori_ori_n214_), .B(ori_ori_n44_), .Y(ori_ori_n554_));
  NO3        o532(.A(ori_ori_n554_), .B(ori_ori_n271_), .C(ori_ori_n217_), .Y(ori_ori_n555_));
  NO2        o533(.A(ori_ori_n114_), .B(ori_ori_n37_), .Y(ori_ori_n556_));
  NO2        o534(.A(ori_ori_n556_), .B(i_6_), .Y(ori_ori_n557_));
  NO2        o535(.A(ori_ori_n81_), .B(i_9_), .Y(ori_ori_n558_));
  NO2        o536(.A(ori_ori_n558_), .B(ori_ori_n59_), .Y(ori_ori_n559_));
  NO2        o537(.A(ori_ori_n559_), .B(ori_ori_n522_), .Y(ori_ori_n560_));
  NO4        o538(.A(ori_ori_n560_), .B(ori_ori_n557_), .C(ori_ori_n555_), .D(i_4_), .Y(ori_ori_n561_));
  NA2        o539(.A(i_1_), .B(i_3_), .Y(ori_ori_n562_));
  NO2        o540(.A(ori_ori_n385_), .B(ori_ori_n88_), .Y(ori_ori_n563_));
  AOI210     o541(.A0(ori_ori_n554_), .A1(ori_ori_n459_), .B0(ori_ori_n563_), .Y(ori_ori_n564_));
  NO2        o542(.A(ori_ori_n564_), .B(ori_ori_n562_), .Y(ori_ori_n565_));
  NO3        o543(.A(ori_ori_n565_), .B(ori_ori_n561_), .C(ori_ori_n553_), .Y(ori_ori_n566_));
  NA4        o544(.A(ori_ori_n566_), .B(ori_ori_n550_), .C(ori_ori_n545_), .D(ori_ori_n524_), .Y(ori_ori_n567_));
  NO3        o545(.A(ori_ori_n400_), .B(i_3_), .C(i_7_), .Y(ori_ori_n568_));
  NOi21      o546(.An(ori_ori_n568_), .B(i_10_), .Y(ori_ori_n569_));
  OA210      o547(.A0(ori_ori_n569_), .A1(ori_ori_n223_), .B0(ori_ori_n81_), .Y(ori_ori_n570_));
  NA3        o548(.A(ori_ori_n402_), .B(ori_ori_n424_), .C(ori_ori_n46_), .Y(ori_ori_n571_));
  NO3        o549(.A(ori_ori_n401_), .B(ori_ori_n495_), .C(ori_ori_n81_), .Y(ori_ori_n572_));
  NA2        o550(.A(ori_ori_n572_), .B(ori_ori_n25_), .Y(ori_ori_n573_));
  NA2        o551(.A(ori_ori_n573_), .B(ori_ori_n571_), .Y(ori_ori_n574_));
  OAI210     o552(.A0(ori_ori_n574_), .A1(ori_ori_n570_), .B0(i_1_), .Y(ori_ori_n575_));
  AOI210     o553(.A0(ori_ori_n242_), .A1(ori_ori_n93_), .B0(i_1_), .Y(ori_ori_n576_));
  NO2        o554(.A(ori_ori_n318_), .B(i_2_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n577_), .B(ori_ori_n576_), .Y(ori_ori_n578_));
  AOI210     o556(.A0(ori_ori_n578_), .A1(ori_ori_n575_), .B0(i_13_), .Y(ori_ori_n579_));
  NO2        o557(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n401_), .B(ori_ori_n24_), .Y(ori_ori_n581_));
  NO2        o559(.A(ori_ori_n873_), .B(ori_ori_n88_), .Y(ori_ori_n582_));
  INV        o560(.A(ori_ori_n582_), .Y(ori_ori_n583_));
  INV        o561(.A(ori_ori_n111_), .Y(ori_ori_n584_));
  AOI220     o562(.A0(ori_ori_n584_), .A1(ori_ori_n68_), .B0(ori_ori_n335_), .B1(ori_ori_n535_), .Y(ori_ori_n585_));
  NO2        o563(.A(ori_ori_n585_), .B(ori_ori_n221_), .Y(ori_ori_n586_));
  AOI210     o564(.A0(ori_ori_n376_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n587_));
  NOi31      o565(.An(ori_ori_n587_), .B(ori_ori_n486_), .C(ori_ori_n44_), .Y(ori_ori_n588_));
  NA2        o566(.A(ori_ori_n124_), .B(i_13_), .Y(ori_ori_n589_));
  NO2        o567(.A(ori_ori_n589_), .B(ori_ori_n576_), .Y(ori_ori_n590_));
  NO3        o568(.A(ori_ori_n67_), .B(ori_ori_n32_), .C(ori_ori_n97_), .Y(ori_ori_n591_));
  NA2        o569(.A(ori_ori_n26_), .B(ori_ori_n181_), .Y(ori_ori_n592_));
  NA2        o570(.A(ori_ori_n592_), .B(i_7_), .Y(ori_ori_n593_));
  NO3        o571(.A(ori_ori_n401_), .B(ori_ori_n216_), .C(ori_ori_n81_), .Y(ori_ori_n594_));
  AOI210     o572(.A0(ori_ori_n594_), .A1(ori_ori_n593_), .B0(ori_ori_n591_), .Y(ori_ori_n595_));
  AOI220     o573(.A0(ori_ori_n335_), .A1(ori_ori_n535_), .B0(ori_ori_n87_), .B1(ori_ori_n98_), .Y(ori_ori_n596_));
  OAI220     o574(.A0(ori_ori_n596_), .A1(ori_ori_n491_), .B0(ori_ori_n595_), .B1(ori_ori_n503_), .Y(ori_ori_n597_));
  NO4        o575(.A(ori_ori_n597_), .B(ori_ori_n590_), .C(ori_ori_n588_), .D(ori_ori_n586_), .Y(ori_ori_n598_));
  OR2        o576(.A(i_11_), .B(i_6_), .Y(ori_ori_n599_));
  NA3        o577(.A(ori_ori_n490_), .B(ori_ori_n592_), .C(i_7_), .Y(ori_ori_n600_));
  NO2        o578(.A(ori_ori_n600_), .B(ori_ori_n599_), .Y(ori_ori_n601_));
  NA3        o579(.A(ori_ori_n360_), .B(ori_ori_n494_), .C(ori_ori_n93_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n527_), .B(i_13_), .Y(ori_ori_n603_));
  NAi21      o581(.An(i_11_), .B(i_12_), .Y(ori_ori_n604_));
  NO3        o582(.A(ori_ori_n401_), .B(ori_ori_n471_), .C(ori_ori_n495_), .Y(ori_ori_n605_));
  NA2        o583(.A(ori_ori_n605_), .B(ori_ori_n274_), .Y(ori_ori_n606_));
  NA3        o584(.A(ori_ori_n606_), .B(ori_ori_n603_), .C(ori_ori_n602_), .Y(ori_ori_n607_));
  OAI210     o585(.A0(ori_ori_n607_), .A1(ori_ori_n601_), .B0(ori_ori_n59_), .Y(ori_ori_n608_));
  NO2        o586(.A(i_2_), .B(i_12_), .Y(ori_ori_n609_));
  NA2        o587(.A(ori_ori_n317_), .B(ori_ori_n609_), .Y(ori_ori_n610_));
  NO2        o588(.A(ori_ori_n125_), .B(i_2_), .Y(ori_ori_n611_));
  NA2        o589(.A(ori_ori_n611_), .B(ori_ori_n522_), .Y(ori_ori_n612_));
  NA2        o590(.A(ori_ori_n612_), .B(ori_ori_n610_), .Y(ori_ori_n613_));
  NA3        o591(.A(ori_ori_n613_), .B(ori_ori_n45_), .C(ori_ori_n209_), .Y(ori_ori_n614_));
  NA4        o592(.A(ori_ori_n614_), .B(ori_ori_n608_), .C(ori_ori_n598_), .D(ori_ori_n583_), .Y(ori_ori_n615_));
  OR4        o593(.A(ori_ori_n615_), .B(ori_ori_n579_), .C(ori_ori_n567_), .D(ori_ori_n505_), .Y(ori5));
  NA2        o594(.A(ori_ori_n547_), .B(ori_ori_n245_), .Y(ori_ori_n617_));
  AN2        o595(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n618_));
  NA3        o596(.A(ori_ori_n618_), .B(ori_ori_n609_), .C(ori_ori_n104_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n491_), .B(i_11_), .Y(ori_ori_n620_));
  NA2        o598(.A(ori_ori_n84_), .B(ori_ori_n620_), .Y(ori_ori_n621_));
  NA3        o599(.A(ori_ori_n621_), .B(ori_ori_n619_), .C(ori_ori_n617_), .Y(ori_ori_n622_));
  NO3        o600(.A(i_11_), .B(ori_ori_n216_), .C(i_13_), .Y(ori_ori_n623_));
  NO2        o601(.A(ori_ori_n121_), .B(ori_ori_n23_), .Y(ori_ori_n624_));
  NA2        o602(.A(i_12_), .B(i_8_), .Y(ori_ori_n625_));
  OAI210     o603(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n625_), .Y(ori_ori_n626_));
  INV        o604(.A(ori_ori_n375_), .Y(ori_ori_n627_));
  AOI220     o605(.A0(ori_ori_n279_), .A1(ori_ori_n463_), .B0(ori_ori_n626_), .B1(ori_ori_n624_), .Y(ori_ori_n628_));
  INV        o606(.A(ori_ori_n628_), .Y(ori_ori_n629_));
  NO2        o607(.A(ori_ori_n629_), .B(ori_ori_n622_), .Y(ori_ori_n630_));
  INV        o608(.A(ori_ori_n163_), .Y(ori_ori_n631_));
  INV        o609(.A(ori_ori_n223_), .Y(ori_ori_n632_));
  OAI210     o610(.A0(ori_ori_n577_), .A1(ori_ori_n377_), .B0(ori_ori_n107_), .Y(ori_ori_n633_));
  AOI210     o611(.A0(ori_ori_n633_), .A1(ori_ori_n632_), .B0(ori_ori_n631_), .Y(ori_ori_n634_));
  NO2        o612(.A(ori_ori_n385_), .B(ori_ori_n26_), .Y(ori_ori_n635_));
  NO2        o613(.A(ori_ori_n635_), .B(ori_ori_n365_), .Y(ori_ori_n636_));
  NA2        o614(.A(ori_ori_n636_), .B(i_2_), .Y(ori_ori_n637_));
  INV        o615(.A(ori_ori_n637_), .Y(ori_ori_n638_));
  AOI210     o616(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n363_), .Y(ori_ori_n639_));
  AOI210     o617(.A0(ori_ori_n639_), .A1(ori_ori_n638_), .B0(ori_ori_n634_), .Y(ori_ori_n640_));
  NO2        o618(.A(ori_ori_n179_), .B(ori_ori_n122_), .Y(ori_ori_n641_));
  OAI210     o619(.A0(ori_ori_n641_), .A1(ori_ori_n624_), .B0(i_2_), .Y(ori_ori_n642_));
  INV        o620(.A(ori_ori_n164_), .Y(ori_ori_n643_));
  NA2        o621(.A(ori_ori_n643_), .B(ori_ori_n84_), .Y(ori_ori_n644_));
  AOI210     o622(.A0(ori_ori_n644_), .A1(ori_ori_n642_), .B0(ori_ori_n181_), .Y(ori_ori_n645_));
  OA210      o623(.A0(ori_ori_n508_), .A1(ori_ori_n123_), .B0(i_13_), .Y(ori_ori_n646_));
  NA2        o624(.A(ori_ori_n187_), .B(ori_ori_n189_), .Y(ori_ori_n647_));
  NA2        o625(.A(ori_ori_n148_), .B(ori_ori_n487_), .Y(ori_ori_n648_));
  AOI210     o626(.A0(ori_ori_n648_), .A1(ori_ori_n647_), .B0(ori_ori_n322_), .Y(ori_ori_n649_));
  AOI210     o627(.A0(ori_ori_n195_), .A1(ori_ori_n145_), .B0(ori_ori_n424_), .Y(ori_ori_n650_));
  NA2        o628(.A(ori_ori_n650_), .B(ori_ori_n365_), .Y(ori_ori_n651_));
  NO2        o629(.A(ori_ori_n98_), .B(ori_ori_n44_), .Y(ori_ori_n652_));
  INV        o630(.A(ori_ori_n268_), .Y(ori_ori_n653_));
  NA4        o631(.A(ori_ori_n653_), .B(ori_ori_n269_), .C(ori_ori_n121_), .D(ori_ori_n42_), .Y(ori_ori_n654_));
  OAI210     o632(.A0(ori_ori_n654_), .A1(ori_ori_n652_), .B0(ori_ori_n651_), .Y(ori_ori_n655_));
  NO4        o633(.A(ori_ori_n655_), .B(ori_ori_n649_), .C(ori_ori_n646_), .D(ori_ori_n645_), .Y(ori_ori_n656_));
  NA2        o634(.A(ori_ori_n463_), .B(ori_ori_n28_), .Y(ori_ori_n657_));
  NA2        o635(.A(ori_ori_n623_), .B(ori_ori_n251_), .Y(ori_ori_n658_));
  NA2        o636(.A(ori_ori_n658_), .B(ori_ori_n657_), .Y(ori_ori_n659_));
  NO2        o637(.A(ori_ori_n58_), .B(i_12_), .Y(ori_ori_n660_));
  NO2        o638(.A(ori_ori_n660_), .B(ori_ori_n123_), .Y(ori_ori_n661_));
  NO2        o639(.A(ori_ori_n661_), .B(ori_ori_n487_), .Y(ori_ori_n662_));
  AOI220     o640(.A0(ori_ori_n662_), .A1(ori_ori_n36_), .B0(ori_ori_n659_), .B1(ori_ori_n46_), .Y(ori_ori_n663_));
  NA4        o641(.A(ori_ori_n663_), .B(ori_ori_n656_), .C(ori_ori_n640_), .D(ori_ori_n630_), .Y(ori6));
  NO3        o642(.A(i_9_), .B(ori_ori_n270_), .C(i_1_), .Y(ori_ori_n665_));
  NO2        o643(.A(ori_ori_n174_), .B(ori_ori_n136_), .Y(ori_ori_n666_));
  OAI210     o644(.A0(ori_ori_n666_), .A1(ori_ori_n665_), .B0(ori_ori_n611_), .Y(ori_ori_n667_));
  NO2        o645(.A(ori_ori_n205_), .B(ori_ori_n404_), .Y(ori_ori_n668_));
  INV        o646(.A(ori_ori_n286_), .Y(ori_ori_n669_));
  AO210      o647(.A0(ori_ori_n669_), .A1(ori_ori_n667_), .B0(i_12_), .Y(ori_ori_n670_));
  NA2        o648(.A(ori_ori_n471_), .B(ori_ori_n59_), .Y(ori_ori_n671_));
  NA2        o649(.A(ori_ori_n569_), .B(ori_ori_n67_), .Y(ori_ori_n672_));
  BUFFER     o650(.A(ori_ori_n513_), .Y(ori_ori_n673_));
  NA3        o651(.A(ori_ori_n673_), .B(ori_ori_n672_), .C(ori_ori_n671_), .Y(ori_ori_n674_));
  NA2        o652(.A(ori_ori_n674_), .B(ori_ori_n69_), .Y(ori_ori_n675_));
  INV        o653(.A(ori_ori_n285_), .Y(ori_ori_n676_));
  NA2        o654(.A(ori_ori_n71_), .B(ori_ori_n128_), .Y(ori_ori_n677_));
  NO2        o655(.A(ori_ori_n677_), .B(ori_ori_n676_), .Y(ori_ori_n678_));
  NO2        o656(.A(ori_ori_n226_), .B(i_9_), .Y(ori_ori_n679_));
  NA2        o657(.A(ori_ori_n679_), .B(ori_ori_n660_), .Y(ori_ori_n680_));
  AOI210     o658(.A0(ori_ori_n680_), .A1(ori_ori_n423_), .B0(ori_ori_n174_), .Y(ori_ori_n681_));
  NO2        o659(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n682_));
  NA3        o660(.A(ori_ori_n682_), .B(ori_ori_n398_), .C(ori_ori_n339_), .Y(ori_ori_n683_));
  NAi32      o661(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n684_));
  NO2        o662(.A(ori_ori_n599_), .B(ori_ori_n684_), .Y(ori_ori_n685_));
  OAI210     o663(.A0(ori_ori_n568_), .A1(ori_ori_n454_), .B0(ori_ori_n453_), .Y(ori_ori_n686_));
  NAi31      o664(.An(ori_ori_n685_), .B(ori_ori_n686_), .C(ori_ori_n683_), .Y(ori_ori_n687_));
  OR3        o665(.A(ori_ori_n687_), .B(ori_ori_n681_), .C(ori_ori_n678_), .Y(ori_ori_n688_));
  AO220      o666(.A0(ori_ori_n308_), .A1(ori_ori_n298_), .B0(ori_ori_n347_), .B1(ori_ori_n487_), .Y(ori_ori_n689_));
  NA3        o667(.A(ori_ori_n689_), .B(ori_ori_n230_), .C(i_7_), .Y(ori_ori_n690_));
  NA3        o668(.A(ori_ori_n377_), .B(ori_ori_n144_), .C(ori_ori_n65_), .Y(ori_ori_n691_));
  AO210      o669(.A0(ori_ori_n409_), .A1(ori_ori_n627_), .B0(ori_ori_n36_), .Y(ori_ori_n692_));
  NA3        o670(.A(ori_ori_n692_), .B(ori_ori_n691_), .C(ori_ori_n690_), .Y(ori_ori_n693_));
  OAI210     o671(.A0(i_6_), .A1(i_11_), .B0(ori_ori_n82_), .Y(ori_ori_n694_));
  AOI220     o672(.A0(ori_ori_n694_), .A1(ori_ori_n453_), .B0(ori_ori_n668_), .B1(ori_ori_n593_), .Y(ori_ori_n695_));
  NA3        o673(.A(ori_ori_n322_), .B(ori_ori_n218_), .C(ori_ori_n144_), .Y(ori_ori_n696_));
  NA2        o674(.A(ori_ori_n347_), .B(ori_ori_n66_), .Y(ori_ori_n697_));
  NA4        o675(.A(ori_ori_n697_), .B(ori_ori_n696_), .C(ori_ori_n695_), .D(ori_ori_n493_), .Y(ori_ori_n698_));
  AO210      o676(.A0(ori_ori_n424_), .A1(ori_ori_n46_), .B0(ori_ori_n83_), .Y(ori_ori_n699_));
  NA3        o677(.A(ori_ori_n699_), .B(ori_ori_n402_), .C(ori_ori_n203_), .Y(ori_ori_n700_));
  AOI210     o678(.A0(ori_ori_n377_), .A1(ori_ori_n375_), .B0(ori_ori_n452_), .Y(ori_ori_n701_));
  NO2        o679(.A(ori_ori_n501_), .B(ori_ori_n98_), .Y(ori_ori_n702_));
  OAI210     o680(.A0(ori_ori_n702_), .A1(ori_ori_n108_), .B0(ori_ori_n358_), .Y(ori_ori_n703_));
  NA2        o681(.A(ori_ori_n222_), .B(ori_ori_n46_), .Y(ori_ori_n704_));
  INV        o682(.A(ori_ori_n476_), .Y(ori_ori_n705_));
  NA3        o683(.A(ori_ori_n705_), .B(ori_ori_n285_), .C(i_7_), .Y(ori_ori_n706_));
  NA4        o684(.A(ori_ori_n706_), .B(ori_ori_n703_), .C(ori_ori_n701_), .D(ori_ori_n700_), .Y(ori_ori_n707_));
  NO4        o685(.A(ori_ori_n707_), .B(ori_ori_n698_), .C(ori_ori_n693_), .D(ori_ori_n688_), .Y(ori_ori_n708_));
  NA4        o686(.A(ori_ori_n708_), .B(ori_ori_n675_), .C(ori_ori_n670_), .D(ori_ori_n329_), .Y(ori3));
  NA2        o687(.A(i_12_), .B(i_10_), .Y(ori_ori_n710_));
  NO2        o688(.A(i_11_), .B(ori_ori_n216_), .Y(ori_ori_n711_));
  NA2        o689(.A(ori_ori_n696_), .B(ori_ori_n493_), .Y(ori_ori_n712_));
  NA2        o690(.A(ori_ori_n712_), .B(ori_ori_n40_), .Y(ori_ori_n713_));
  NO3        o691(.A(ori_ori_n518_), .B(ori_ori_n385_), .C(ori_ori_n128_), .Y(ori_ori_n714_));
  NA2        o692(.A(ori_ori_n360_), .B(ori_ori_n45_), .Y(ori_ori_n715_));
  INV        o693(.A(ori_ori_n714_), .Y(ori_ori_n716_));
  AOI210     o694(.A0(ori_ori_n716_), .A1(ori_ori_n713_), .B0(ori_ori_n48_), .Y(ori_ori_n717_));
  NO4        o695(.A(ori_ori_n326_), .B(ori_ori_n332_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n718_));
  NA2        o696(.A(ori_ori_n587_), .B(ori_ori_n558_), .Y(ori_ori_n719_));
  NA2        o697(.A(ori_ori_n292_), .B(i_5_), .Y(ori_ori_n720_));
  OAI220     o698(.A0(ori_ori_n720_), .A1(ori_ori_n719_), .B0(ori_ori_n875_), .B1(ori_ori_n59_), .Y(ori_ori_n721_));
  NOi21      o699(.An(i_5_), .B(i_9_), .Y(ori_ori_n722_));
  NA2        o700(.A(ori_ori_n722_), .B(ori_ori_n374_), .Y(ori_ori_n723_));
  BUFFER     o701(.A(ori_ori_n242_), .Y(ori_ori_n724_));
  AOI210     o702(.A0(ori_ori_n724_), .A1(ori_ori_n399_), .B0(ori_ori_n572_), .Y(ori_ori_n725_));
  NO3        o703(.A(ori_ori_n361_), .B(ori_ori_n242_), .C(ori_ori_n69_), .Y(ori_ori_n726_));
  NO2        o704(.A(ori_ori_n166_), .B(ori_ori_n145_), .Y(ori_ori_n727_));
  AOI210     o705(.A0(ori_ori_n727_), .A1(ori_ori_n222_), .B0(ori_ori_n726_), .Y(ori_ori_n728_));
  OAI220     o706(.A0(ori_ori_n728_), .A1(ori_ori_n169_), .B0(ori_ori_n725_), .B1(ori_ori_n723_), .Y(ori_ori_n729_));
  NO3        o707(.A(ori_ori_n729_), .B(ori_ori_n721_), .C(ori_ori_n717_), .Y(ori_ori_n730_));
  NA2        o708(.A(ori_ori_n174_), .B(ori_ori_n24_), .Y(ori_ori_n731_));
  NO2        o709(.A(ori_ori_n556_), .B(ori_ori_n484_), .Y(ori_ori_n732_));
  NO2        o710(.A(ori_ori_n732_), .B(ori_ori_n731_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n274_), .B(ori_ori_n126_), .Y(ori_ori_n734_));
  NAi21      o712(.An(ori_ori_n155_), .B(i_5_), .Y(ori_ori_n735_));
  OAI220     o713(.A0(ori_ori_n735_), .A1(ori_ori_n704_), .B0(ori_ori_n734_), .B1(ori_ori_n352_), .Y(ori_ori_n736_));
  NO2        o714(.A(ori_ori_n736_), .B(ori_ori_n733_), .Y(ori_ori_n737_));
  NA2        o715(.A(ori_ori_n460_), .B(i_0_), .Y(ori_ori_n738_));
  NO3        o716(.A(ori_ori_n738_), .B(ori_ori_n334_), .C(ori_ori_n84_), .Y(ori_ori_n739_));
  NO4        o717(.A(ori_ori_n475_), .B(ori_ori_n200_), .C(ori_ori_n363_), .D(ori_ori_n359_), .Y(ori_ori_n740_));
  AOI210     o718(.A0(ori_ori_n740_), .A1(i_11_), .B0(ori_ori_n739_), .Y(ori_ori_n741_));
  INV        o719(.A(ori_ori_n398_), .Y(ori_ori_n742_));
  NA2        o720(.A(ori_ori_n623_), .B(ori_ori_n286_), .Y(ori_ori_n743_));
  AOI210     o721(.A0(ori_ori_n402_), .A1(ori_ori_n84_), .B0(ori_ori_n56_), .Y(ori_ori_n744_));
  OAI220     o722(.A0(ori_ori_n744_), .A1(ori_ori_n743_), .B0(ori_ori_n542_), .B1(ori_ori_n432_), .Y(ori_ori_n745_));
  NO2        o723(.A(ori_ori_n228_), .B(ori_ori_n149_), .Y(ori_ori_n746_));
  NA2        o724(.A(i_0_), .B(i_10_), .Y(ori_ori_n747_));
  INV        o725(.A(ori_ori_n434_), .Y(ori_ori_n748_));
  NO4        o726(.A(ori_ori_n111_), .B(ori_ori_n56_), .C(ori_ori_n551_), .D(i_5_), .Y(ori_ori_n749_));
  AO220      o727(.A0(ori_ori_n749_), .A1(ori_ori_n748_), .B0(ori_ori_n746_), .B1(i_6_), .Y(ori_ori_n750_));
  NA2        o728(.A(ori_ori_n177_), .B(ori_ori_n189_), .Y(ori_ori_n751_));
  NO2        o729(.A(ori_ori_n751_), .B(ori_ori_n743_), .Y(ori_ori_n752_));
  NO3        o730(.A(ori_ori_n752_), .B(ori_ori_n750_), .C(ori_ori_n745_), .Y(ori_ori_n753_));
  NA3        o731(.A(ori_ori_n753_), .B(ori_ori_n741_), .C(ori_ori_n737_), .Y(ori_ori_n754_));
  NA2        o732(.A(i_11_), .B(i_9_), .Y(ori_ori_n755_));
  NA2        o733(.A(ori_ori_n344_), .B(ori_ori_n167_), .Y(ori_ori_n756_));
  NA2        o734(.A(ori_ori_n756_), .B(ori_ori_n153_), .Y(ori_ori_n757_));
  NO2        o735(.A(ori_ori_n755_), .B(ori_ori_n69_), .Y(ori_ori_n758_));
  NO2        o736(.A(ori_ori_n166_), .B(i_0_), .Y(ori_ori_n759_));
  INV        o737(.A(ori_ori_n757_), .Y(ori_ori_n760_));
  NA2        o738(.A(ori_ori_n541_), .B(ori_ori_n118_), .Y(ori_ori_n761_));
  NO2        o739(.A(i_6_), .B(ori_ori_n761_), .Y(ori_ori_n762_));
  AOI210     o740(.A0(ori_ori_n376_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n763_));
  NA2        o741(.A(ori_ori_n163_), .B(ori_ori_n99_), .Y(ori_ori_n764_));
  NOi32      o742(.An(ori_ori_n763_), .Bn(ori_ori_n177_), .C(ori_ori_n764_), .Y(ori_ori_n765_));
  NA2        o743(.A(ori_ori_n494_), .B(ori_ori_n286_), .Y(ori_ori_n766_));
  NO2        o744(.A(ori_ori_n766_), .B(ori_ori_n715_), .Y(ori_ori_n767_));
  NO3        o745(.A(ori_ori_n767_), .B(ori_ori_n765_), .C(ori_ori_n762_), .Y(ori_ori_n768_));
  NOi21      o746(.An(i_7_), .B(i_5_), .Y(ori_ori_n769_));
  NOi31      o747(.An(ori_ori_n769_), .B(i_0_), .C(ori_ori_n604_), .Y(ori_ori_n770_));
  NA3        o748(.A(ori_ori_n770_), .B(ori_ori_n333_), .C(i_6_), .Y(ori_ori_n771_));
  OA210      o749(.A0(ori_ori_n764_), .A1(ori_ori_n423_), .B0(ori_ori_n771_), .Y(ori_ori_n772_));
  INV        o750(.A(ori_ori_n280_), .Y(ori_ori_n773_));
  NA3        o751(.A(ori_ori_n772_), .B(ori_ori_n768_), .C(ori_ori_n760_), .Y(ori_ori_n774_));
  NO2        o752(.A(ori_ori_n710_), .B(ori_ori_n279_), .Y(ori_ori_n775_));
  NA2        o753(.A(ori_ori_n775_), .B(ori_ori_n758_), .Y(ori_ori_n776_));
  NA3        o754(.A(ori_ori_n397_), .B(ori_ori_n360_), .C(ori_ori_n45_), .Y(ori_ori_n777_));
  OAI210     o755(.A0(ori_ori_n735_), .A1(ori_ori_n742_), .B0(ori_ori_n777_), .Y(ori_ori_n778_));
  NO2        o756(.A(ori_ori_n230_), .B(ori_ori_n46_), .Y(ori_ori_n779_));
  NA2        o757(.A(ori_ori_n758_), .B(ori_ori_n269_), .Y(ori_ori_n780_));
  OAI210     o758(.A0(ori_ori_n779_), .A1(ori_ori_n176_), .B0(ori_ori_n780_), .Y(ori_ori_n781_));
  AOI220     o759(.A0(ori_ori_n781_), .A1(ori_ori_n398_), .B0(ori_ori_n778_), .B1(ori_ori_n69_), .Y(ori_ori_n782_));
  NO2        o760(.A(ori_ori_n71_), .B(ori_ori_n625_), .Y(ori_ori_n783_));
  AOI210     o761(.A0(ori_ori_n165_), .A1(ori_ori_n484_), .B0(ori_ori_n783_), .Y(ori_ori_n784_));
  NO2        o762(.A(ori_ori_n784_), .B(ori_ori_n47_), .Y(ori_ori_n785_));
  NO3        o763(.A(ori_ori_n475_), .B(ori_ori_n306_), .C(ori_ori_n24_), .Y(ori_ori_n786_));
  AOI210     o764(.A0(ori_ori_n581_), .A1(ori_ori_n442_), .B0(ori_ori_n786_), .Y(ori_ori_n787_));
  NAi21      o765(.An(i_9_), .B(i_5_), .Y(ori_ori_n788_));
  NO2        o766(.A(ori_ori_n787_), .B(ori_ori_n164_), .Y(ori_ori_n789_));
  NO2        o767(.A(ori_ori_n789_), .B(ori_ori_n785_), .Y(ori_ori_n790_));
  NA3        o768(.A(ori_ori_n790_), .B(ori_ori_n782_), .C(ori_ori_n776_), .Y(ori_ori_n791_));
  NO3        o769(.A(ori_ori_n791_), .B(ori_ori_n774_), .C(ori_ori_n754_), .Y(ori_ori_n792_));
  NO2        o770(.A(i_0_), .B(ori_ori_n604_), .Y(ori_ori_n793_));
  NA2        o771(.A(ori_ori_n69_), .B(ori_ori_n44_), .Y(ori_ori_n794_));
  AN2        o772(.A(ori_ori_n793_), .B(ori_ori_n165_), .Y(ori_ori_n795_));
  NO2        o773(.A(ori_ori_n671_), .B(ori_ori_n764_), .Y(ori_ori_n796_));
  AOI210     o774(.A0(ori_ori_n795_), .A1(ori_ori_n297_), .B0(ori_ori_n796_), .Y(ori_ori_n797_));
  NO2        o775(.A(ori_ori_n686_), .B(ori_ori_n353_), .Y(ori_ori_n798_));
  NA2        o776(.A(ori_ori_n222_), .B(ori_ori_n213_), .Y(ori_ori_n799_));
  AOI210     o777(.A0(ori_ori_n799_), .A1(ori_ori_n738_), .B0(ori_ori_n149_), .Y(ori_ori_n800_));
  NO2        o778(.A(ori_ori_n800_), .B(ori_ori_n798_), .Y(ori_ori_n801_));
  NA2        o779(.A(ori_ori_n801_), .B(ori_ori_n797_), .Y(ori_ori_n802_));
  NO3        o780(.A(ori_ori_n747_), .B(ori_ori_n722_), .C(ori_ori_n179_), .Y(ori_ori_n803_));
  AOI220     o781(.A0(ori_ori_n803_), .A1(i_11_), .B0(ori_ori_n456_), .B1(ori_ori_n71_), .Y(ori_ori_n804_));
  NO3        o782(.A(ori_ori_n196_), .B(ori_ori_n332_), .C(i_0_), .Y(ori_ori_n805_));
  OAI210     o783(.A0(ori_ori_n805_), .A1(ori_ori_n72_), .B0(i_13_), .Y(ori_ori_n806_));
  NA2        o784(.A(ori_ori_n806_), .B(ori_ori_n804_), .Y(ori_ori_n807_));
  INV        o785(.A(ori_ori_n105_), .Y(ori_ori_n808_));
  OR2        o786(.A(ori_ori_n808_), .B(i_5_), .Y(ori_ori_n809_));
  NO3        o787(.A(ori_ori_n715_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n810_));
  NA2        o788(.A(ori_ori_n408_), .B(ori_ori_n403_), .Y(ori_ori_n811_));
  NO2        o789(.A(ori_ori_n811_), .B(ori_ori_n810_), .Y(ori_ori_n812_));
  NA3        o790(.A(ori_ori_n339_), .B(ori_ori_n163_), .C(ori_ori_n162_), .Y(ori_ori_n813_));
  INV        o791(.A(ori_ori_n813_), .Y(ori_ori_n814_));
  NA3        o792(.A(ori_ori_n339_), .B(ori_ori_n293_), .C(ori_ori_n206_), .Y(ori_ori_n815_));
  INV        o793(.A(ori_ori_n815_), .Y(ori_ori_n816_));
  NOi31      o794(.An(ori_ori_n338_), .B(ori_ori_n794_), .C(ori_ori_n219_), .Y(ori_ori_n817_));
  NO3        o795(.A(ori_ori_n755_), .B(ori_ori_n203_), .C(ori_ori_n179_), .Y(ori_ori_n818_));
  NO4        o796(.A(ori_ori_n818_), .B(ori_ori_n817_), .C(ori_ori_n816_), .D(ori_ori_n814_), .Y(ori_ori_n819_));
  NA3        o797(.A(ori_ori_n819_), .B(ori_ori_n812_), .C(ori_ori_n809_), .Y(ori_ori_n820_));
  NO2        o798(.A(ori_ori_n81_), .B(i_5_), .Y(ori_ori_n821_));
  NA3        o799(.A(ori_ori_n711_), .B(ori_ori_n106_), .C(ori_ori_n121_), .Y(ori_ori_n822_));
  INV        o800(.A(ori_ori_n822_), .Y(ori_ori_n823_));
  NA2        o801(.A(ori_ori_n823_), .B(ori_ori_n821_), .Y(ori_ori_n824_));
  NA3        o802(.A(ori_ori_n269_), .B(i_5_), .C(ori_ori_n181_), .Y(ori_ori_n825_));
  NAi31      o803(.An(ori_ori_n220_), .B(ori_ori_n825_), .C(ori_ori_n221_), .Y(ori_ori_n826_));
  NO4        o804(.A(ori_ori_n219_), .B(ori_ori_n196_), .C(i_0_), .D(i_12_), .Y(ori_ori_n827_));
  NA2        o805(.A(ori_ori_n827_), .B(ori_ori_n826_), .Y(ori_ori_n828_));
  AN2        o806(.A(ori_ori_n747_), .B(ori_ori_n149_), .Y(ori_ori_n829_));
  NO4        o807(.A(ori_ori_n829_), .B(i_12_), .C(ori_ori_n532_), .D(ori_ori_n128_), .Y(ori_ori_n830_));
  NA2        o808(.A(ori_ori_n830_), .B(ori_ori_n203_), .Y(ori_ori_n831_));
  NA3        o809(.A(ori_ori_n94_), .B(ori_ori_n459_), .C(i_11_), .Y(ori_ori_n832_));
  NO2        o810(.A(ori_ori_n832_), .B(ori_ori_n69_), .Y(ori_ori_n833_));
  NA2        o811(.A(ori_ori_n60_), .B(ori_ori_n97_), .Y(ori_ori_n834_));
  NO2        o812(.A(ori_ori_n834_), .B(ori_ori_n825_), .Y(ori_ori_n835_));
  AOI210     o813(.A0(ori_ori_n835_), .A1(ori_ori_n759_), .B0(ori_ori_n833_), .Y(ori_ori_n836_));
  NA4        o814(.A(ori_ori_n836_), .B(ori_ori_n831_), .C(ori_ori_n828_), .D(ori_ori_n824_), .Y(ori_ori_n837_));
  NO4        o815(.A(ori_ori_n837_), .B(ori_ori_n820_), .C(ori_ori_n807_), .D(ori_ori_n802_), .Y(ori_ori_n838_));
  NA2        o816(.A(ori_ori_n682_), .B(ori_ori_n37_), .Y(ori_ori_n839_));
  NA3        o817(.A(ori_ori_n763_), .B(ori_ori_n317_), .C(i_5_), .Y(ori_ori_n840_));
  NA3        o818(.A(ori_ori_n840_), .B(ori_ori_n839_), .C(ori_ori_n500_), .Y(ori_ori_n841_));
  NA2        o819(.A(ori_ori_n841_), .B(ori_ori_n194_), .Y(ori_ori_n842_));
  BUFFER     o820(.A(ori_ori_n318_), .Y(ori_ori_n843_));
  NA2        o821(.A(ori_ori_n175_), .B(ori_ori_n177_), .Y(ori_ori_n844_));
  AO210      o822(.A0(ori_ori_n843_), .A1(ori_ori_n33_), .B0(ori_ori_n844_), .Y(ori_ori_n845_));
  INV        o823(.A(ori_ori_n529_), .Y(ori_ori_n846_));
  NA2        o824(.A(ori_ori_n846_), .B(ori_ori_n845_), .Y(ori_ori_n847_));
  AOI210     o825(.A0(ori_ori_n847_), .A1(ori_ori_n48_), .B0(ori_ori_n740_), .Y(ori_ori_n848_));
  AOI210     o826(.A0(ori_ori_n848_), .A1(ori_ori_n842_), .B0(ori_ori_n69_), .Y(ori_ori_n849_));
  INV        o827(.A(ori_ori_n72_), .Y(ori_ori_n850_));
  INV        o828(.A(ori_ori_n770_), .Y(ori_ori_n851_));
  AOI210     o829(.A0(ori_ori_n851_), .A1(ori_ori_n850_), .B0(ori_ori_n562_), .Y(ori_ori_n852_));
  INV        o830(.A(ori_ori_n852_), .Y(ori_ori_n853_));
  OAI210     o831(.A0(ori_ori_n244_), .A1(ori_ori_n151_), .B0(ori_ori_n84_), .Y(ori_ori_n854_));
  NA3        o832(.A(ori_ori_n635_), .B(ori_ori_n260_), .C(ori_ori_n76_), .Y(ori_ori_n855_));
  AOI210     o833(.A0(ori_ori_n855_), .A1(ori_ori_n854_), .B0(i_11_), .Y(ori_ori_n856_));
  NA2        o834(.A(ori_ori_n495_), .B(ori_ori_n200_), .Y(ori_ori_n857_));
  OAI210     o835(.A0(ori_ori_n857_), .A1(ori_ori_n763_), .B0(ori_ori_n194_), .Y(ori_ori_n858_));
  NA2        o836(.A(ori_ori_n157_), .B(i_5_), .Y(ori_ori_n859_));
  NO2        o837(.A(ori_ori_n858_), .B(ori_ori_n859_), .Y(ori_ori_n860_));
  NO3        o838(.A(ori_ori_n57_), .B(ori_ori_n56_), .C(i_4_), .Y(ori_ori_n861_));
  OAI210     o839(.A0(ori_ori_n773_), .A1(ori_ori_n270_), .B0(ori_ori_n861_), .Y(ori_ori_n862_));
  NO2        o840(.A(ori_ori_n862_), .B(ori_ori_n604_), .Y(ori_ori_n863_));
  NO4        o841(.A(ori_ori_n788_), .B(ori_ori_n400_), .C(ori_ori_n227_), .D(ori_ori_n226_), .Y(ori_ori_n864_));
  NO2        o842(.A(ori_ori_n864_), .B(ori_ori_n452_), .Y(ori_ori_n865_));
  NO2        o843(.A(ori_ori_n865_), .B(ori_ori_n41_), .Y(ori_ori_n866_));
  NO4        o844(.A(ori_ori_n866_), .B(ori_ori_n863_), .C(ori_ori_n860_), .D(ori_ori_n856_), .Y(ori_ori_n867_));
  OAI210     o845(.A0(ori_ori_n853_), .A1(i_4_), .B0(ori_ori_n867_), .Y(ori_ori_n868_));
  NO2        o846(.A(ori_ori_n868_), .B(ori_ori_n849_), .Y(ori_ori_n869_));
  NA4        o847(.A(ori_ori_n869_), .B(ori_ori_n838_), .C(ori_ori_n792_), .D(ori_ori_n730_), .Y(ori4));
  INV        o848(.A(ori_ori_n580_), .Y(ori_ori_n873_));
  INV        o849(.A(ori_ori_n78_), .Y(ori_ori_n874_));
  INV        o850(.A(ori_ori_n718_), .Y(ori_ori_n875_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m021(.A(mai_mai_n35_), .Y(mai1));
  INV        m022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m064(.A(i_6_), .Y(mai_mai_n87_));
  NO2        m065(.A(i_2_), .B(i_7_), .Y(mai_mai_n88_));
  INV        m066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  OAI210     m067(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NAi21      m068(.An(i_6_), .B(i_10_), .Y(mai_mai_n91_));
  NA2        m069(.A(i_6_), .B(i_9_), .Y(mai_mai_n92_));
  AOI210     m070(.A0(mai_mai_n92_), .A1(mai_mai_n91_), .B0(mai_mai_n64_), .Y(mai_mai_n93_));
  NA2        m071(.A(i_2_), .B(i_6_), .Y(mai_mai_n94_));
  NO3        m072(.A(mai_mai_n94_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n95_));
  NO2        m073(.A(mai_mai_n95_), .B(mai_mai_n93_), .Y(mai_mai_n96_));
  AOI210     m074(.A0(mai_mai_n96_), .A1(mai_mai_n90_), .B0(mai_mai_n81_), .Y(mai_mai_n97_));
  AN3        m075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n98_));
  NAi21      m076(.An(i_6_), .B(i_11_), .Y(mai_mai_n99_));
  NO2        m077(.A(i_5_), .B(i_8_), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n98_), .B(mai_mai_n32_), .Y(mai_mai_n101_));
  INV        m079(.A(i_7_), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n47_), .B(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m081(.A(i_0_), .B(i_5_), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n104_), .B(mai_mai_n87_), .Y(mai_mai_n105_));
  NA2        m083(.A(i_12_), .B(i_3_), .Y(mai_mai_n106_));
  INV        m084(.A(mai_mai_n106_), .Y(mai_mai_n107_));
  NA3        m085(.A(mai_mai_n107_), .B(mai_mai_n105_), .C(mai_mai_n103_), .Y(mai_mai_n108_));
  NAi21      m086(.An(i_7_), .B(i_11_), .Y(mai_mai_n109_));
  NO3        m087(.A(mai_mai_n109_), .B(mai_mai_n91_), .C(mai_mai_n54_), .Y(mai_mai_n110_));
  AN2        m088(.A(i_2_), .B(i_10_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n111_), .B(i_7_), .Y(mai_mai_n112_));
  OR2        m090(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n113_));
  NO2        m091(.A(i_8_), .B(mai_mai_n102_), .Y(mai_mai_n114_));
  NA2        m092(.A(i_12_), .B(i_7_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n116_));
  NA2        m094(.A(i_11_), .B(i_12_), .Y(mai_mai_n117_));
  NAi41      m095(.An(mai_mai_n110_), .B(mai_mai_n117_), .C(mai_mai_n108_), .D(mai_mai_n101_), .Y(mai_mai_n118_));
  NOi21      m096(.An(i_1_), .B(i_5_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(i_11_), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n102_), .B(mai_mai_n37_), .Y(mai_mai_n121_));
  NA2        m099(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n122_));
  NA2        m100(.A(mai_mai_n122_), .B(mai_mai_n121_), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n123_), .B(mai_mai_n47_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n92_), .B(mai_mai_n91_), .Y(mai_mai_n125_));
  NAi21      m103(.An(i_3_), .B(i_8_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n126_), .B(mai_mai_n63_), .Y(mai_mai_n127_));
  NOi31      m105(.An(mai_mai_n127_), .B(mai_mai_n125_), .C(mai_mai_n124_), .Y(mai_mai_n128_));
  NO2        m106(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n129_));
  NO2        m107(.A(i_6_), .B(i_5_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(i_3_), .Y(mai_mai_n131_));
  AO210      m109(.A0(mai_mai_n131_), .A1(mai_mai_n48_), .B0(mai_mai_n129_), .Y(mai_mai_n132_));
  OAI220     m110(.A0(mai_mai_n132_), .A1(mai_mai_n109_), .B0(mai_mai_n128_), .B1(mai_mai_n120_), .Y(mai_mai_n133_));
  NO3        m111(.A(mai_mai_n133_), .B(mai_mai_n118_), .C(mai_mai_n97_), .Y(mai_mai_n134_));
  NA3        m112(.A(mai_mai_n134_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m113(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n136_));
  NA2        m114(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n138_));
  NA4        m116(.A(mai_mai_n138_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m117(.A(i_8_), .B(i_7_), .Y(mai_mai_n140_));
  NA2        m118(.A(mai_mai_n140_), .B(i_6_), .Y(mai_mai_n141_));
  NO2        m119(.A(i_12_), .B(i_13_), .Y(mai_mai_n142_));
  NAi21      m120(.An(i_5_), .B(i_11_), .Y(mai_mai_n143_));
  NOi21      m121(.An(mai_mai_n142_), .B(mai_mai_n143_), .Y(mai_mai_n144_));
  NO2        m122(.A(i_0_), .B(i_1_), .Y(mai_mai_n145_));
  NA2        m123(.A(i_2_), .B(i_3_), .Y(mai_mai_n146_));
  NO2        m124(.A(mai_mai_n146_), .B(i_4_), .Y(mai_mai_n147_));
  NA3        m125(.A(mai_mai_n147_), .B(mai_mai_n145_), .C(mai_mai_n144_), .Y(mai_mai_n148_));
  OR2        m126(.A(mai_mai_n148_), .B(mai_mai_n25_), .Y(mai_mai_n149_));
  AN2        m127(.A(mai_mai_n142_), .B(mai_mai_n84_), .Y(mai_mai_n150_));
  NO2        m128(.A(mai_mai_n150_), .B(mai_mai_n27_), .Y(mai_mai_n151_));
  NA2        m129(.A(i_1_), .B(i_5_), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n74_), .B(mai_mai_n47_), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n153_), .B(mai_mai_n36_), .Y(mai_mai_n154_));
  NO3        m132(.A(mai_mai_n154_), .B(mai_mai_n152_), .C(mai_mai_n151_), .Y(mai_mai_n155_));
  OR2        m133(.A(i_0_), .B(i_1_), .Y(mai_mai_n156_));
  NO3        m134(.A(mai_mai_n156_), .B(mai_mai_n81_), .C(i_13_), .Y(mai_mai_n157_));
  NAi32      m135(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n158_));
  NOi21      m136(.An(i_4_), .B(i_10_), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n159_), .B(mai_mai_n40_), .Y(mai_mai_n160_));
  NO2        m138(.A(i_3_), .B(i_5_), .Y(mai_mai_n161_));
  INV        m139(.A(mai_mai_n155_), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n162_), .A1(mai_mai_n149_), .B0(mai_mai_n141_), .Y(mai_mai_n163_));
  NA3        m141(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_4_), .B(i_9_), .Y(mai_mai_n165_));
  NOi21      m143(.An(i_11_), .B(i_13_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  BUFFER     m145(.A(mai_mai_n167_), .Y(mai_mai_n168_));
  NO2        m146(.A(i_4_), .B(i_5_), .Y(mai_mai_n169_));
  NAi21      m147(.An(i_12_), .B(i_11_), .Y(mai_mai_n170_));
  NO2        m148(.A(mai_mai_n170_), .B(i_13_), .Y(mai_mai_n171_));
  NA3        m149(.A(mai_mai_n171_), .B(mai_mai_n169_), .C(mai_mai_n84_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(mai_mai_n172_), .A1(mai_mai_n168_), .B0(mai_mai_n164_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n175_));
  NA2        m153(.A(i_3_), .B(i_5_), .Y(mai_mai_n176_));
  NO2        m154(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n177_));
  NO2        m155(.A(i_13_), .B(i_10_), .Y(mai_mai_n178_));
  NA3        m156(.A(mai_mai_n178_), .B(mai_mai_n177_), .C(mai_mai_n45_), .Y(mai_mai_n179_));
  NO2        m157(.A(i_2_), .B(i_1_), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n180_), .B(i_3_), .Y(mai_mai_n181_));
  NAi21      m159(.An(i_4_), .B(i_12_), .Y(mai_mai_n182_));
  NO4        m160(.A(mai_mai_n182_), .B(mai_mai_n181_), .C(mai_mai_n179_), .D(mai_mai_n25_), .Y(mai_mai_n183_));
  NO2        m161(.A(mai_mai_n183_), .B(mai_mai_n173_), .Y(mai_mai_n184_));
  INV        m162(.A(i_8_), .Y(mai_mai_n185_));
  NO2        m163(.A(mai_mai_n185_), .B(i_7_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n186_), .B(i_6_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(mai_mai_n114_), .Y(mai_mai_n189_));
  NO3        m167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n190_));
  NA3        m168(.A(mai_mai_n190_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n191_));
  NO3        m169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n192_));
  OAI210     m170(.A0(mai_mai_n98_), .A1(i_12_), .B0(mai_mai_n192_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n193_), .B(mai_mai_n189_), .Y(mai_mai_n194_));
  NO2        m172(.A(i_3_), .B(i_8_), .Y(mai_mai_n195_));
  NO3        m173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n104_), .B(mai_mai_n59_), .Y(mai_mai_n197_));
  NO2        m175(.A(i_13_), .B(i_9_), .Y(mai_mai_n198_));
  NA3        m176(.A(mai_mai_n198_), .B(i_6_), .C(mai_mai_n185_), .Y(mai_mai_n199_));
  NAi21      m177(.An(i_12_), .B(i_3_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n201_));
  NO3        m179(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n202_));
  NA3        m180(.A(mai_mai_n202_), .B(mai_mai_n201_), .C(i_10_), .Y(mai_mai_n203_));
  NO2        m181(.A(mai_mai_n203_), .B(mai_mai_n199_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(mai_mai_n194_), .Y(mai_mai_n205_));
  OAI220     m183(.A0(mai_mai_n205_), .A1(i_4_), .B0(mai_mai_n187_), .B1(mai_mai_n184_), .Y(mai_mai_n206_));
  NAi21      m184(.An(i_12_), .B(i_7_), .Y(mai_mai_n207_));
  NA3        m185(.A(i_13_), .B(mai_mai_n185_), .C(i_10_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n209_));
  NA2        m187(.A(i_0_), .B(i_5_), .Y(mai_mai_n210_));
  NA2        m188(.A(mai_mai_n210_), .B(mai_mai_n105_), .Y(mai_mai_n211_));
  OAI220     m189(.A0(mai_mai_n211_), .A1(mai_mai_n181_), .B0(i_2_), .B1(mai_mai_n131_), .Y(mai_mai_n212_));
  NAi31      m190(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n216_));
  INV        m194(.A(i_13_), .Y(mai_mai_n217_));
  NO2        m195(.A(i_12_), .B(mai_mai_n217_), .Y(mai_mai_n218_));
  NA3        m196(.A(mai_mai_n218_), .B(mai_mai_n190_), .C(mai_mai_n188_), .Y(mai_mai_n219_));
  INV        m197(.A(mai_mai_n219_), .Y(mai_mai_n220_));
  AOI220     m198(.A0(mai_mai_n220_), .A1(mai_mai_n140_), .B0(mai_mai_n212_), .B1(mai_mai_n209_), .Y(mai_mai_n221_));
  NO2        m199(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n176_), .B(i_4_), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n223_), .B(mai_mai_n222_), .Y(mai_mai_n224_));
  OR2        m202(.A(i_8_), .B(i_7_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n225_), .B(mai_mai_n87_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n227_));
  NA2        m205(.A(mai_mai_n227_), .B(mai_mai_n226_), .Y(mai_mai_n228_));
  INV        m206(.A(i_12_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n45_), .B(mai_mai_n229_), .Y(mai_mai_n230_));
  NO3        m208(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n231_));
  NA2        m209(.A(i_2_), .B(i_1_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n228_), .B(mai_mai_n224_), .Y(mai_mai_n233_));
  NO3        m211(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n234_));
  NAi21      m212(.An(i_4_), .B(i_3_), .Y(mai_mai_n235_));
  NO2        m213(.A(i_0_), .B(i_6_), .Y(mai_mai_n236_));
  NOi41      m214(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n237_), .B(mai_mai_n236_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n232_), .B(mai_mai_n176_), .Y(mai_mai_n239_));
  NAi21      m217(.An(mai_mai_n238_), .B(mai_mai_n239_), .Y(mai_mai_n240_));
  INV        m218(.A(mai_mai_n240_), .Y(mai_mai_n241_));
  AOI220     m219(.A0(mai_mai_n241_), .A1(mai_mai_n40_), .B0(mai_mai_n233_), .B1(mai_mai_n198_), .Y(mai_mai_n242_));
  NO2        m220(.A(i_11_), .B(mai_mai_n217_), .Y(mai_mai_n243_));
  NOi21      m221(.An(i_1_), .B(i_6_), .Y(mai_mai_n244_));
  NAi21      m222(.An(i_3_), .B(i_7_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n246_));
  NO2        m224(.A(i_12_), .B(i_3_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n248_));
  NA3        m226(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n225_), .B(mai_mai_n37_), .Y(mai_mai_n250_));
  NA2        m228(.A(i_12_), .B(i_6_), .Y(mai_mai_n251_));
  OR2        m229(.A(i_13_), .B(i_9_), .Y(mai_mai_n252_));
  NO3        m230(.A(mai_mai_n252_), .B(mai_mai_n251_), .C(mai_mai_n49_), .Y(mai_mai_n253_));
  NO2        m231(.A(mai_mai_n235_), .B(i_2_), .Y(mai_mai_n254_));
  NA3        m232(.A(mai_mai_n254_), .B(mai_mai_n253_), .C(mai_mai_n45_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n243_), .B(i_9_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n248_), .B(mai_mai_n65_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n257_), .A1(mai_mai_n256_), .B0(mai_mai_n255_), .Y(mai_mai_n258_));
  NA2        m236(.A(mai_mai_n153_), .B(mai_mai_n64_), .Y(mai_mai_n259_));
  NO3        m237(.A(i_11_), .B(mai_mai_n217_), .C(mai_mai_n25_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n245_), .B(i_8_), .Y(mai_mai_n261_));
  NA3        m239(.A(i_5_), .B(mai_mai_n261_), .C(mai_mai_n260_), .Y(mai_mai_n262_));
  NO3        m240(.A(mai_mai_n26_), .B(mai_mai_n87_), .C(i_5_), .Y(mai_mai_n263_));
  NA3        m241(.A(mai_mai_n263_), .B(mai_mai_n250_), .C(mai_mai_n218_), .Y(mai_mai_n264_));
  AOI210     m242(.A0(mai_mai_n264_), .A1(mai_mai_n262_), .B0(mai_mai_n259_), .Y(mai_mai_n265_));
  AOI210     m243(.A0(mai_mai_n258_), .A1(mai_mai_n250_), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  NA3        m244(.A(mai_mai_n266_), .B(mai_mai_n242_), .C(mai_mai_n221_), .Y(mai_mai_n267_));
  NO3        m245(.A(i_12_), .B(mai_mai_n217_), .C(mai_mai_n37_), .Y(mai_mai_n268_));
  INV        m246(.A(mai_mai_n268_), .Y(mai_mai_n269_));
  NA2        m247(.A(i_8_), .B(mai_mai_n102_), .Y(mai_mai_n270_));
  NO3        m248(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n232_), .B(i_0_), .Y(mai_mai_n272_));
  NA2        m250(.A(i_0_), .B(i_1_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n273_), .B(i_2_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n275_));
  NA3        m253(.A(mai_mai_n275_), .B(mai_mai_n274_), .C(mai_mai_n161_), .Y(mai_mai_n276_));
  NO2        m254(.A(i_3_), .B(i_10_), .Y(mai_mai_n277_));
  NA3        m255(.A(mai_mai_n277_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n278_));
  NO2        m256(.A(i_2_), .B(mai_mai_n102_), .Y(mai_mai_n279_));
  NO2        m257(.A(i_4_), .B(i_8_), .Y(mai_mai_n280_));
  NOi21      m258(.An(mai_mai_n210_), .B(mai_mai_n104_), .Y(mai_mai_n281_));
  NA3        m259(.A(mai_mai_n281_), .B(mai_mai_n280_), .C(mai_mai_n279_), .Y(mai_mai_n282_));
  AN2        m260(.A(i_3_), .B(i_10_), .Y(mai_mai_n283_));
  NA4        m261(.A(mai_mai_n283_), .B(mai_mai_n190_), .C(mai_mai_n171_), .D(mai_mai_n169_), .Y(mai_mai_n284_));
  NO2        m262(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n286_));
  OR2        m264(.A(mai_mai_n282_), .B(mai_mai_n278_), .Y(mai_mai_n287_));
  OAI220     m265(.A0(mai_mai_n287_), .A1(i_6_), .B0(mai_mai_n276_), .B1(mai_mai_n269_), .Y(mai_mai_n288_));
  NO4        m266(.A(mai_mai_n288_), .B(mai_mai_n267_), .C(mai_mai_n206_), .D(mai_mai_n163_), .Y(mai_mai_n289_));
  NO3        m267(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n290_));
  NO2        m268(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n291_));
  NO3        m269(.A(i_6_), .B(mai_mai_n185_), .C(i_7_), .Y(mai_mai_n292_));
  NO2        m270(.A(i_2_), .B(i_3_), .Y(mai_mai_n293_));
  OR2        m271(.A(i_0_), .B(i_5_), .Y(mai_mai_n294_));
  NA2        m272(.A(mai_mai_n210_), .B(mai_mai_n294_), .Y(mai_mai_n295_));
  NA4        m273(.A(mai_mai_n295_), .B(mai_mai_n226_), .C(mai_mai_n293_), .D(i_1_), .Y(mai_mai_n296_));
  NAi21      m274(.An(i_8_), .B(i_7_), .Y(mai_mai_n297_));
  NO2        m275(.A(mai_mai_n297_), .B(i_6_), .Y(mai_mai_n298_));
  NO2        m276(.A(mai_mai_n156_), .B(mai_mai_n47_), .Y(mai_mai_n299_));
  NA3        m277(.A(mai_mai_n299_), .B(mai_mai_n298_), .C(mai_mai_n161_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n300_), .B(mai_mai_n296_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n301_), .B(i_4_), .Y(mai_mai_n302_));
  NO2        m280(.A(i_12_), .B(i_10_), .Y(mai_mai_n303_));
  NOi21      m281(.An(i_5_), .B(i_0_), .Y(mai_mai_n304_));
  NO2        m282(.A(i_6_), .B(i_8_), .Y(mai_mai_n305_));
  NOi21      m283(.An(i_0_), .B(i_2_), .Y(mai_mai_n306_));
  AN2        m284(.A(mai_mai_n306_), .B(mai_mai_n305_), .Y(mai_mai_n307_));
  NO2        m285(.A(i_1_), .B(i_7_), .Y(mai_mai_n308_));
  AO220      m286(.A0(mai_mai_n308_), .A1(mai_mai_n307_), .B0(mai_mai_n298_), .B1(mai_mai_n227_), .Y(mai_mai_n309_));
  NA2        m287(.A(mai_mai_n309_), .B(mai_mai_n42_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n310_), .B(mai_mai_n302_), .Y(mai_mai_n311_));
  NO3        m289(.A(mai_mai_n225_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n312_));
  NO3        m290(.A(mai_mai_n297_), .B(i_2_), .C(i_1_), .Y(mai_mai_n313_));
  OAI210     m291(.A0(mai_mai_n313_), .A1(mai_mai_n312_), .B0(i_6_), .Y(mai_mai_n314_));
  INV        m292(.A(mai_mai_n314_), .Y(mai_mai_n315_));
  NOi21      m293(.An(mai_mai_n152_), .B(mai_mai_n105_), .Y(mai_mai_n316_));
  NO2        m294(.A(mai_mai_n316_), .B(mai_mai_n122_), .Y(mai_mai_n317_));
  OAI210     m295(.A0(mai_mai_n317_), .A1(mai_mai_n315_), .B0(i_3_), .Y(mai_mai_n318_));
  NO2        m296(.A(mai_mai_n273_), .B(mai_mai_n82_), .Y(mai_mai_n319_));
  NA2        m297(.A(mai_mai_n319_), .B(mai_mai_n130_), .Y(mai_mai_n320_));
  NO2        m298(.A(mai_mai_n94_), .B(mai_mai_n185_), .Y(mai_mai_n321_));
  NA3        m299(.A(mai_mai_n281_), .B(mai_mai_n321_), .C(mai_mai_n64_), .Y(mai_mai_n322_));
  AOI210     m300(.A0(mai_mai_n322_), .A1(mai_mai_n320_), .B0(i_7_), .Y(mai_mai_n323_));
  NO2        m301(.A(mai_mai_n185_), .B(i_9_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n324_), .B(mai_mai_n197_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n325_), .B(mai_mai_n47_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n326_), .B(mai_mai_n323_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n327_), .A1(mai_mai_n318_), .B0(mai_mai_n160_), .Y(mai_mai_n328_));
  AOI210     m306(.A0(mai_mai_n311_), .A1(mai_mai_n290_), .B0(mai_mai_n328_), .Y(mai_mai_n329_));
  NOi32      m307(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n330_));
  INV        m308(.A(mai_mai_n330_), .Y(mai_mai_n331_));
  NAi21      m309(.An(i_0_), .B(i_6_), .Y(mai_mai_n332_));
  NAi21      m310(.An(i_1_), .B(i_5_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n333_), .B(mai_mai_n332_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n334_), .B(mai_mai_n25_), .Y(mai_mai_n335_));
  OAI210     m313(.A0(mai_mai_n335_), .A1(mai_mai_n158_), .B0(mai_mai_n238_), .Y(mai_mai_n336_));
  NAi41      m314(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n337_));
  OAI220     m315(.A0(mai_mai_n337_), .A1(mai_mai_n333_), .B0(mai_mai_n213_), .B1(mai_mai_n158_), .Y(mai_mai_n338_));
  AOI210     m316(.A0(mai_mai_n337_), .A1(mai_mai_n158_), .B0(mai_mai_n156_), .Y(mai_mai_n339_));
  NOi32      m317(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n340_));
  NAi21      m318(.An(i_6_), .B(i_1_), .Y(mai_mai_n341_));
  NA3        m319(.A(mai_mai_n341_), .B(mai_mai_n340_), .C(mai_mai_n47_), .Y(mai_mai_n342_));
  NO2        m320(.A(mai_mai_n342_), .B(i_0_), .Y(mai_mai_n343_));
  OR3        m321(.A(mai_mai_n343_), .B(mai_mai_n339_), .C(mai_mai_n338_), .Y(mai_mai_n344_));
  NO2        m322(.A(i_1_), .B(mai_mai_n102_), .Y(mai_mai_n345_));
  NAi21      m323(.An(i_3_), .B(i_4_), .Y(mai_mai_n346_));
  NO2        m324(.A(mai_mai_n346_), .B(i_9_), .Y(mai_mai_n347_));
  AN2        m325(.A(i_6_), .B(i_7_), .Y(mai_mai_n348_));
  OAI210     m326(.A0(mai_mai_n348_), .A1(mai_mai_n345_), .B0(mai_mai_n347_), .Y(mai_mai_n349_));
  NA2        m327(.A(i_2_), .B(i_7_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n346_), .B(i_10_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n349_), .B(mai_mai_n177_), .Y(mai_mai_n352_));
  AOI210     m330(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n180_), .B0(mai_mai_n351_), .Y(mai_mai_n354_));
  AOI220     m332(.A0(mai_mai_n351_), .A1(mai_mai_n308_), .B0(mai_mai_n231_), .B1(mai_mai_n180_), .Y(mai_mai_n355_));
  AOI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n354_), .B0(i_5_), .Y(mai_mai_n356_));
  NO4        m334(.A(mai_mai_n356_), .B(mai_mai_n352_), .C(mai_mai_n344_), .D(mai_mai_n336_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n357_), .B(mai_mai_n331_), .Y(mai_mai_n358_));
  AN2        m336(.A(i_12_), .B(i_5_), .Y(mai_mai_n359_));
  NO2        m337(.A(i_11_), .B(i_6_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n235_), .B(i_5_), .Y(mai_mai_n361_));
  NO2        m339(.A(i_5_), .B(i_10_), .Y(mai_mai_n362_));
  NO2        m340(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n363_));
  NO3        m341(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n364_));
  NO2        m342(.A(i_11_), .B(i_12_), .Y(mai_mai_n365_));
  NA3        m343(.A(mai_mai_n114_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n366_));
  NO2        m344(.A(mai_mai_n366_), .B(mai_mai_n213_), .Y(mai_mai_n367_));
  NAi21      m345(.An(i_13_), .B(i_0_), .Y(mai_mai_n368_));
  INV        m346(.A(mai_mai_n368_), .Y(mai_mai_n369_));
  NA2        m347(.A(mai_mai_n367_), .B(mai_mai_n369_), .Y(mai_mai_n370_));
  INV        m348(.A(mai_mai_n370_), .Y(mai_mai_n371_));
  NO3        m349(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n372_));
  NO2        m350(.A(i_0_), .B(i_11_), .Y(mai_mai_n373_));
  INV        m351(.A(i_5_), .Y(mai_mai_n374_));
  AN2        m352(.A(i_1_), .B(i_6_), .Y(mai_mai_n375_));
  NOi21      m353(.An(i_2_), .B(i_12_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n376_), .B(mai_mai_n375_), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n377_), .B(mai_mai_n374_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n140_), .B(i_9_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(i_4_), .Y(mai_mai_n380_));
  NA2        m358(.A(mai_mai_n378_), .B(mai_mai_n380_), .Y(mai_mai_n381_));
  NAi21      m359(.An(i_9_), .B(i_4_), .Y(mai_mai_n382_));
  OR2        m360(.A(i_13_), .B(i_10_), .Y(mai_mai_n383_));
  NO3        m361(.A(mai_mai_n383_), .B(mai_mai_n117_), .C(mai_mai_n382_), .Y(mai_mai_n384_));
  NO2        m362(.A(mai_mai_n167_), .B(mai_mai_n121_), .Y(mai_mai_n385_));
  OR2        m363(.A(mai_mai_n208_), .B(mai_mai_n207_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n102_), .B(mai_mai_n25_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n268_), .B(mai_mai_n387_), .Y(mai_mai_n388_));
  NA2        m366(.A(i_5_), .B(mai_mai_n202_), .Y(mai_mai_n389_));
  OAI220     m367(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n388_), .B1(mai_mai_n316_), .Y(mai_mai_n390_));
  INV        m368(.A(mai_mai_n390_), .Y(mai_mai_n391_));
  AOI210     m369(.A0(mai_mai_n391_), .A1(mai_mai_n381_), .B0(mai_mai_n26_), .Y(mai_mai_n392_));
  INV        m370(.A(mai_mai_n296_), .Y(mai_mai_n393_));
  AOI220     m371(.A0(mai_mai_n275_), .A1(mai_mai_n271_), .B0(mai_mai_n272_), .B1(mai_mai_n291_), .Y(mai_mai_n394_));
  NO2        m372(.A(mai_mai_n394_), .B(i_5_), .Y(mai_mai_n395_));
  AOI220     m373(.A0(i_3_), .A1(mai_mai_n274_), .B0(mai_mai_n263_), .B1(mai_mai_n202_), .Y(mai_mai_n396_));
  NO2        m374(.A(mai_mai_n396_), .B(mai_mai_n270_), .Y(mai_mai_n397_));
  NO3        m375(.A(mai_mai_n397_), .B(mai_mai_n395_), .C(mai_mai_n393_), .Y(mai_mai_n398_));
  NA2        m376(.A(mai_mai_n188_), .B(mai_mai_n98_), .Y(mai_mai_n399_));
  NA3        m377(.A(mai_mai_n299_), .B(mai_mai_n161_), .C(mai_mai_n87_), .Y(mai_mai_n400_));
  AOI210     m378(.A0(mai_mai_n400_), .A1(mai_mai_n399_), .B0(mai_mai_n297_), .Y(mai_mai_n401_));
  NA3        m379(.A(mai_mai_n308_), .B(mai_mai_n307_), .C(i_5_), .Y(mai_mai_n402_));
  INV        m380(.A(mai_mai_n292_), .Y(mai_mai_n403_));
  OAI210     m381(.A0(mai_mai_n403_), .A1(mai_mai_n181_), .B0(mai_mai_n402_), .Y(mai_mai_n404_));
  NO2        m382(.A(mai_mai_n404_), .B(mai_mai_n401_), .Y(mai_mai_n405_));
  AOI210     m383(.A0(mai_mai_n405_), .A1(mai_mai_n398_), .B0(mai_mai_n256_), .Y(mai_mai_n406_));
  NO4        m384(.A(mai_mai_n406_), .B(mai_mai_n392_), .C(mai_mai_n371_), .D(mai_mai_n358_), .Y(mai_mai_n407_));
  NO2        m385(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n408_));
  NO2        m386(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n409_));
  NO2        m387(.A(i_10_), .B(i_9_), .Y(mai_mai_n410_));
  NAi21      m388(.An(i_12_), .B(i_8_), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n411_), .B(i_3_), .Y(mai_mai_n412_));
  NA2        m390(.A(mai_mai_n286_), .B(i_0_), .Y(mai_mai_n413_));
  NO3        m391(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n414_));
  NA2        m392(.A(mai_mai_n251_), .B(mai_mai_n99_), .Y(mai_mai_n415_));
  NA2        m393(.A(mai_mai_n415_), .B(mai_mai_n414_), .Y(mai_mai_n416_));
  NA2        m394(.A(i_8_), .B(i_9_), .Y(mai_mai_n417_));
  NA2        m395(.A(mai_mai_n268_), .B(mai_mai_n197_), .Y(mai_mai_n418_));
  OAI220     m396(.A0(mai_mai_n418_), .A1(mai_mai_n417_), .B0(mai_mai_n416_), .B1(mai_mai_n413_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n243_), .B(mai_mai_n285_), .Y(mai_mai_n420_));
  NO3        m398(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n421_));
  INV        m399(.A(mai_mai_n421_), .Y(mai_mai_n422_));
  NA3        m400(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n423_));
  NA4        m401(.A(mai_mai_n143_), .B(mai_mai_n116_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n424_));
  OAI220     m402(.A0(mai_mai_n424_), .A1(mai_mai_n423_), .B0(mai_mai_n422_), .B1(mai_mai_n420_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n425_), .B(mai_mai_n419_), .Y(mai_mai_n426_));
  OR2        m404(.A(mai_mai_n273_), .B(mai_mai_n199_), .Y(mai_mai_n427_));
  OA210      m405(.A0(mai_mai_n325_), .A1(mai_mai_n102_), .B0(mai_mai_n276_), .Y(mai_mai_n428_));
  OA220      m406(.A0(mai_mai_n428_), .A1(mai_mai_n160_), .B0(mai_mai_n427_), .B1(mai_mai_n224_), .Y(mai_mai_n429_));
  NO2        m407(.A(i_2_), .B(i_13_), .Y(mai_mai_n430_));
  NO3        m408(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n431_));
  NO2        m409(.A(i_6_), .B(i_7_), .Y(mai_mai_n432_));
  NA2        m410(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  NO2        m411(.A(i_11_), .B(i_1_), .Y(mai_mai_n434_));
  OR2        m412(.A(i_11_), .B(i_8_), .Y(mai_mai_n435_));
  NOi21      m413(.An(i_2_), .B(i_7_), .Y(mai_mai_n436_));
  NAi31      m414(.An(mai_mai_n435_), .B(mai_mai_n436_), .C(i_0_), .Y(mai_mai_n437_));
  INV        m415(.A(mai_mai_n383_), .Y(mai_mai_n438_));
  NA3        m416(.A(mai_mai_n438_), .B(mai_mai_n408_), .C(mai_mai_n76_), .Y(mai_mai_n439_));
  NO2        m417(.A(mai_mai_n439_), .B(mai_mai_n437_), .Y(mai_mai_n440_));
  NO2        m418(.A(i_3_), .B(mai_mai_n185_), .Y(mai_mai_n441_));
  NO2        m419(.A(i_6_), .B(i_10_), .Y(mai_mai_n442_));
  NA4        m420(.A(mai_mai_n442_), .B(mai_mai_n290_), .C(mai_mai_n441_), .D(mai_mai_n229_), .Y(mai_mai_n443_));
  NO2        m421(.A(mai_mai_n443_), .B(mai_mai_n154_), .Y(mai_mai_n444_));
  NA3        m422(.A(mai_mai_n237_), .B(mai_mai_n166_), .C(mai_mai_n130_), .Y(mai_mai_n445_));
  NA2        m423(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n446_));
  NO2        m424(.A(mai_mai_n156_), .B(i_3_), .Y(mai_mai_n447_));
  NAi31      m425(.An(mai_mai_n446_), .B(mai_mai_n447_), .C(mai_mai_n218_), .Y(mai_mai_n448_));
  NA3        m426(.A(mai_mai_n363_), .B(mai_mai_n174_), .C(mai_mai_n147_), .Y(mai_mai_n449_));
  NA3        m427(.A(mai_mai_n449_), .B(mai_mai_n448_), .C(mai_mai_n445_), .Y(mai_mai_n450_));
  NO3        m428(.A(mai_mai_n450_), .B(mai_mai_n444_), .C(mai_mai_n440_), .Y(mai_mai_n451_));
  NA2        m429(.A(mai_mai_n414_), .B(mai_mai_n359_), .Y(mai_mai_n452_));
  NAi21      m430(.An(mai_mai_n208_), .B(mai_mai_n365_), .Y(mai_mai_n453_));
  NA2        m431(.A(mai_mai_n308_), .B(mai_mai_n210_), .Y(mai_mai_n454_));
  NO2        m432(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n455_));
  NO2        m433(.A(i_0_), .B(mai_mai_n87_), .Y(mai_mai_n456_));
  NA3        m434(.A(mai_mai_n456_), .B(mai_mai_n455_), .C(mai_mai_n140_), .Y(mai_mai_n457_));
  OR3        m435(.A(i_4_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n458_));
  OAI220     m436(.A0(mai_mai_n458_), .A1(mai_mai_n457_), .B0(mai_mai_n454_), .B1(mai_mai_n453_), .Y(mai_mai_n459_));
  NA4        m437(.A(mai_mai_n283_), .B(mai_mai_n216_), .C(mai_mai_n74_), .D(mai_mai_n229_), .Y(mai_mai_n460_));
  NO2        m438(.A(mai_mai_n460_), .B(mai_mai_n433_), .Y(mai_mai_n461_));
  NO2        m439(.A(mai_mai_n461_), .B(mai_mai_n459_), .Y(mai_mai_n462_));
  NA4        m440(.A(mai_mai_n462_), .B(mai_mai_n451_), .C(mai_mai_n429_), .D(mai_mai_n426_), .Y(mai_mai_n463_));
  NA3        m441(.A(mai_mai_n283_), .B(mai_mai_n171_), .C(mai_mai_n169_), .Y(mai_mai_n464_));
  INV        m442(.A(mai_mai_n464_), .Y(mai_mai_n465_));
  BUFFER     m443(.A(mai_mai_n226_), .Y(mai_mai_n466_));
  NA2        m444(.A(mai_mai_n466_), .B(mai_mai_n465_), .Y(mai_mai_n467_));
  NA2        m445(.A(mai_mai_n290_), .B(i_0_), .Y(mai_mai_n468_));
  OAI210     m446(.A0(mai_mai_n468_), .A1(mai_mai_n224_), .B0(mai_mai_n284_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n469_), .B(mai_mai_n298_), .Y(mai_mai_n470_));
  NA2        m448(.A(mai_mai_n359_), .B(mai_mai_n217_), .Y(mai_mai_n471_));
  NA2        m449(.A(mai_mai_n330_), .B(mai_mai_n74_), .Y(mai_mai_n472_));
  NA2        m450(.A(mai_mai_n348_), .B(mai_mai_n340_), .Y(mai_mai_n473_));
  OR2        m451(.A(mai_mai_n471_), .B(mai_mai_n473_), .Y(mai_mai_n474_));
  NO2        m452(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n475_));
  NAi41      m453(.An(mai_mai_n472_), .B(mai_mai_n442_), .C(mai_mai_n475_), .D(mai_mai_n47_), .Y(mai_mai_n476_));
  AOI210     m454(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n384_), .Y(mai_mai_n477_));
  NA3        m455(.A(mai_mai_n477_), .B(mai_mai_n476_), .C(mai_mai_n474_), .Y(mai_mai_n478_));
  INV        m456(.A(mai_mai_n478_), .Y(mai_mai_n479_));
  NA2        m457(.A(mai_mai_n248_), .B(mai_mai_n65_), .Y(mai_mai_n480_));
  OAI210     m458(.A0(i_8_), .A1(mai_mai_n480_), .B0(mai_mai_n132_), .Y(mai_mai_n481_));
  AOI210     m459(.A0(mai_mai_n186_), .A1(i_9_), .B0(mai_mai_n250_), .Y(mai_mai_n482_));
  NO2        m460(.A(mai_mai_n482_), .B(mai_mai_n191_), .Y(mai_mai_n483_));
  OR2        m461(.A(mai_mai_n176_), .B(i_4_), .Y(mai_mai_n484_));
  INV        m462(.A(mai_mai_n484_), .Y(mai_mai_n485_));
  AOI220     m463(.A0(mai_mai_n485_), .A1(mai_mai_n483_), .B0(mai_mai_n481_), .B1(mai_mai_n385_), .Y(mai_mai_n486_));
  NA4        m464(.A(mai_mai_n486_), .B(mai_mai_n479_), .C(mai_mai_n470_), .D(mai_mai_n467_), .Y(mai_mai_n487_));
  NA2        m465(.A(mai_mai_n361_), .B(mai_mai_n274_), .Y(mai_mai_n488_));
  OAI210     m466(.A0(mai_mai_n972_), .A1(mai_mai_n164_), .B0(mai_mai_n488_), .Y(mai_mai_n489_));
  NO2        m467(.A(i_12_), .B(mai_mai_n185_), .Y(mai_mai_n490_));
  NA2        m468(.A(mai_mai_n490_), .B(mai_mai_n217_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n442_), .B(mai_mai_n27_), .Y(mai_mai_n492_));
  NO2        m470(.A(mai_mai_n492_), .B(mai_mai_n491_), .Y(mai_mai_n493_));
  NOi31      m471(.An(mai_mai_n292_), .B(mai_mai_n383_), .C(mai_mai_n38_), .Y(mai_mai_n494_));
  OAI210     m472(.A0(mai_mai_n494_), .A1(mai_mai_n493_), .B0(mai_mai_n489_), .Y(mai_mai_n495_));
  AOI220     m473(.A0(mai_mai_n299_), .A1(mai_mai_n40_), .B0(mai_mai_n227_), .B1(mai_mai_n198_), .Y(mai_mai_n496_));
  NO2        m474(.A(mai_mai_n496_), .B(mai_mai_n484_), .Y(mai_mai_n497_));
  NA2        m475(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n498_));
  NO2        m476(.A(mai_mai_n498_), .B(i_6_), .Y(mai_mai_n499_));
  NA2        m477(.A(mai_mai_n499_), .B(mai_mai_n497_), .Y(mai_mai_n500_));
  NOi31      m478(.An(mai_mai_n272_), .B(mai_mai_n278_), .C(mai_mai_n175_), .Y(mai_mai_n501_));
  NA3        m479(.A(mai_mai_n283_), .B(mai_mai_n169_), .C(mai_mai_n98_), .Y(mai_mai_n502_));
  NO2        m480(.A(mai_mai_n156_), .B(i_5_), .Y(mai_mai_n503_));
  NA2        m481(.A(mai_mai_n503_), .B(mai_mai_n293_), .Y(mai_mai_n504_));
  NA2        m482(.A(mai_mai_n504_), .B(mai_mai_n502_), .Y(mai_mai_n505_));
  OAI210     m483(.A0(mai_mai_n505_), .A1(mai_mai_n501_), .B0(mai_mai_n421_), .Y(mai_mai_n506_));
  NA3        m484(.A(mai_mai_n506_), .B(mai_mai_n500_), .C(mai_mai_n495_), .Y(mai_mai_n507_));
  NA3        m485(.A(mai_mai_n210_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n508_));
  NA2        m486(.A(mai_mai_n268_), .B(mai_mai_n85_), .Y(mai_mai_n509_));
  AOI210     m487(.A0(mai_mai_n508_), .A1(mai_mai_n320_), .B0(mai_mai_n509_), .Y(mai_mai_n510_));
  NA2        m488(.A(mai_mai_n275_), .B(mai_mai_n271_), .Y(mai_mai_n511_));
  NO2        m489(.A(mai_mai_n511_), .B(mai_mai_n168_), .Y(mai_mai_n512_));
  NA2        m490(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n513_));
  NA2        m491(.A(mai_mai_n410_), .B(mai_mai_n214_), .Y(mai_mai_n514_));
  NO2        m492(.A(mai_mai_n513_), .B(mai_mai_n514_), .Y(mai_mai_n515_));
  AOI210     m493(.A0(mai_mai_n341_), .A1(mai_mai_n47_), .B0(mai_mai_n345_), .Y(mai_mai_n516_));
  NA2        m494(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n517_));
  NA3        m495(.A(mai_mai_n490_), .B(mai_mai_n260_), .C(mai_mai_n517_), .Y(mai_mai_n518_));
  NO2        m496(.A(mai_mai_n516_), .B(mai_mai_n518_), .Y(mai_mai_n519_));
  NO4        m497(.A(mai_mai_n519_), .B(mai_mai_n515_), .C(mai_mai_n512_), .D(mai_mai_n510_), .Y(mai_mai_n520_));
  NO4        m498(.A(mai_mai_n244_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n521_));
  NO3        m499(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n522_));
  NO2        m500(.A(mai_mai_n225_), .B(mai_mai_n36_), .Y(mai_mai_n523_));
  AN2        m501(.A(mai_mai_n523_), .B(mai_mai_n522_), .Y(mai_mai_n524_));
  OA210      m502(.A0(mai_mai_n524_), .A1(mai_mai_n521_), .B0(mai_mai_n330_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n383_), .B(i_1_), .Y(mai_mai_n526_));
  NOi31      m504(.An(mai_mai_n526_), .B(mai_mai_n415_), .C(mai_mai_n74_), .Y(mai_mai_n527_));
  AN4        m505(.A(mai_mai_n527_), .B(mai_mai_n380_), .C(mai_mai_n455_), .D(i_2_), .Y(mai_mai_n528_));
  NO2        m506(.A(mai_mai_n394_), .B(mai_mai_n172_), .Y(mai_mai_n529_));
  NO3        m507(.A(mai_mai_n529_), .B(mai_mai_n528_), .C(mai_mai_n525_), .Y(mai_mai_n530_));
  NOi21      m508(.An(i_10_), .B(i_6_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n532_));
  AOI220     m510(.A0(mai_mai_n268_), .A1(mai_mai_n532_), .B0(mai_mai_n260_), .B1(mai_mai_n531_), .Y(mai_mai_n533_));
  NO2        m511(.A(mai_mai_n533_), .B(mai_mai_n413_), .Y(mai_mai_n534_));
  NO2        m512(.A(mai_mai_n115_), .B(mai_mai_n23_), .Y(mai_mai_n535_));
  INV        m513(.A(mai_mai_n534_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n472_), .B(mai_mai_n355_), .Y(mai_mai_n537_));
  INV        m515(.A(mai_mai_n293_), .Y(mai_mai_n538_));
  NO2        m516(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n539_));
  NA3        m517(.A(mai_mai_n539_), .B(mai_mai_n260_), .C(mai_mai_n517_), .Y(mai_mai_n540_));
  NA3        m518(.A(mai_mai_n360_), .B(mai_mai_n268_), .C(mai_mai_n210_), .Y(mai_mai_n541_));
  AOI210     m519(.A0(mai_mai_n541_), .A1(mai_mai_n540_), .B0(mai_mai_n538_), .Y(mai_mai_n542_));
  NO3        m520(.A(i_4_), .B(mai_mai_n314_), .C(mai_mai_n278_), .Y(mai_mai_n543_));
  OR2        m521(.A(i_2_), .B(i_5_), .Y(mai_mai_n544_));
  OR2        m522(.A(mai_mai_n544_), .B(mai_mai_n375_), .Y(mai_mai_n545_));
  NO2        m523(.A(mai_mai_n545_), .B(mai_mai_n453_), .Y(mai_mai_n546_));
  NO4        m524(.A(mai_mai_n546_), .B(mai_mai_n543_), .C(mai_mai_n542_), .D(mai_mai_n537_), .Y(mai_mai_n547_));
  NA4        m525(.A(mai_mai_n547_), .B(mai_mai_n536_), .C(mai_mai_n530_), .D(mai_mai_n520_), .Y(mai_mai_n548_));
  NO4        m526(.A(mai_mai_n548_), .B(mai_mai_n507_), .C(mai_mai_n487_), .D(mai_mai_n463_), .Y(mai_mai_n549_));
  NA4        m527(.A(mai_mai_n549_), .B(mai_mai_n407_), .C(mai_mai_n329_), .D(mai_mai_n289_), .Y(mai7));
  NO2        m528(.A(mai_mai_n94_), .B(mai_mai_n55_), .Y(mai_mai_n551_));
  NA2        m529(.A(i_11_), .B(mai_mai_n185_), .Y(mai_mai_n552_));
  NA3        m530(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n553_));
  NO2        m531(.A(mai_mai_n229_), .B(i_4_), .Y(mai_mai_n554_));
  NA2        m532(.A(mai_mai_n554_), .B(i_8_), .Y(mai_mai_n555_));
  NO2        m533(.A(mai_mai_n106_), .B(mai_mai_n553_), .Y(mai_mai_n556_));
  NA2        m534(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n557_));
  OAI210     m535(.A0(mai_mai_n88_), .A1(mai_mai_n195_), .B0(mai_mai_n196_), .Y(mai_mai_n558_));
  NO2        m536(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n559_));
  NA2        m537(.A(i_4_), .B(i_8_), .Y(mai_mai_n560_));
  AOI210     m538(.A0(mai_mai_n560_), .A1(mai_mai_n283_), .B0(mai_mai_n559_), .Y(mai_mai_n561_));
  OAI220     m539(.A0(mai_mai_n561_), .A1(mai_mai_n557_), .B0(mai_mai_n558_), .B1(i_13_), .Y(mai_mai_n562_));
  NO3        m540(.A(mai_mai_n562_), .B(mai_mai_n556_), .C(mai_mai_n551_), .Y(mai_mai_n563_));
  INV        m541(.A(mai_mai_n159_), .Y(mai_mai_n564_));
  OR2        m542(.A(i_6_), .B(i_10_), .Y(mai_mai_n565_));
  NO2        m543(.A(mai_mai_n565_), .B(mai_mai_n23_), .Y(mai_mai_n566_));
  OR3        m544(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n567_));
  NO3        m545(.A(mai_mai_n567_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n568_));
  INV        m546(.A(mai_mai_n192_), .Y(mai_mai_n569_));
  NO2        m547(.A(mai_mai_n568_), .B(mai_mai_n566_), .Y(mai_mai_n570_));
  OA220      m548(.A0(mai_mai_n570_), .A1(mai_mai_n538_), .B0(mai_mai_n564_), .B1(mai_mai_n252_), .Y(mai_mai_n571_));
  AOI210     m549(.A0(mai_mai_n571_), .A1(mai_mai_n563_), .B0(mai_mai_n64_), .Y(mai_mai_n572_));
  NOi21      m550(.An(i_11_), .B(i_7_), .Y(mai_mai_n573_));
  AO210      m551(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n574_));
  NO2        m552(.A(mai_mai_n574_), .B(mai_mai_n573_), .Y(mai_mai_n575_));
  NA2        m553(.A(mai_mai_n575_), .B(mai_mai_n198_), .Y(mai_mai_n576_));
  NA3        m554(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n577_));
  NAi31      m555(.An(mai_mai_n577_), .B(mai_mai_n207_), .C(i_11_), .Y(mai_mai_n578_));
  AOI210     m556(.A0(mai_mai_n578_), .A1(mai_mai_n576_), .B0(mai_mai_n64_), .Y(mai_mai_n579_));
  NO3        m557(.A(i_7_), .B(mai_mai_n200_), .C(mai_mai_n552_), .Y(mai_mai_n580_));
  OAI210     m558(.A0(mai_mai_n580_), .A1(mai_mai_n218_), .B0(mai_mai_n64_), .Y(mai_mai_n581_));
  NO2        m559(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n582_));
  NO2        m560(.A(i_1_), .B(i_12_), .Y(mai_mai_n583_));
  NA3        m561(.A(mai_mai_n583_), .B(mai_mai_n111_), .C(mai_mai_n24_), .Y(mai_mai_n584_));
  BUFFER     m562(.A(mai_mai_n584_), .Y(mai_mai_n585_));
  NA2        m563(.A(mai_mai_n585_), .B(mai_mai_n581_), .Y(mai_mai_n586_));
  OAI210     m564(.A0(mai_mai_n586_), .A1(mai_mai_n579_), .B0(i_6_), .Y(mai_mai_n587_));
  NO2        m565(.A(mai_mai_n577_), .B(mai_mai_n109_), .Y(mai_mai_n588_));
  NA2        m566(.A(mai_mai_n588_), .B(mai_mai_n539_), .Y(mai_mai_n589_));
  NO2        m567(.A(i_6_), .B(i_11_), .Y(mai_mai_n590_));
  NA2        m568(.A(mai_mai_n589_), .B(mai_mai_n416_), .Y(mai_mai_n591_));
  NO4        m569(.A(mai_mai_n207_), .B(mai_mai_n126_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n592_));
  NA2        m570(.A(mai_mai_n592_), .B(mai_mai_n582_), .Y(mai_mai_n593_));
  NA2        m571(.A(mai_mai_n229_), .B(i_6_), .Y(mai_mai_n594_));
  INV        m572(.A(mai_mai_n593_), .Y(mai_mai_n595_));
  INV        m573(.A(i_2_), .Y(mai_mai_n596_));
  NA2        m574(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n597_));
  NA3        m575(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n598_));
  NO2        m576(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n599_));
  NA3        m577(.A(mai_mai_n599_), .B(mai_mai_n251_), .C(mai_mai_n45_), .Y(mai_mai_n600_));
  OAI220     m578(.A0(mai_mai_n600_), .A1(mai_mai_n598_), .B0(mai_mai_n597_), .B1(mai_mai_n596_), .Y(mai_mai_n601_));
  NA3        m579(.A(mai_mai_n582_), .B(mai_mai_n293_), .C(i_6_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n602_), .B(mai_mai_n23_), .Y(mai_mai_n603_));
  AOI210     m581(.A0(mai_mai_n434_), .A1(mai_mai_n387_), .B0(mai_mai_n234_), .Y(mai_mai_n604_));
  NO2        m582(.A(mai_mai_n604_), .B(mai_mai_n557_), .Y(mai_mai_n605_));
  NO2        m583(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n606_));
  OR3        m584(.A(mai_mai_n605_), .B(mai_mai_n603_), .C(mai_mai_n601_), .Y(mai_mai_n607_));
  NO3        m585(.A(mai_mai_n607_), .B(mai_mai_n595_), .C(mai_mai_n591_), .Y(mai_mai_n608_));
  NO2        m586(.A(mai_mai_n229_), .B(mai_mai_n102_), .Y(mai_mai_n609_));
  NO2        m587(.A(mai_mai_n609_), .B(mai_mai_n573_), .Y(mai_mai_n610_));
  NA2        m588(.A(mai_mai_n610_), .B(i_1_), .Y(mai_mai_n611_));
  NO2        m589(.A(mai_mai_n611_), .B(mai_mai_n567_), .Y(mai_mai_n612_));
  NO2        m590(.A(mai_mai_n382_), .B(mai_mai_n87_), .Y(mai_mai_n613_));
  NA2        m591(.A(mai_mai_n612_), .B(mai_mai_n47_), .Y(mai_mai_n614_));
  NA2        m592(.A(i_3_), .B(mai_mai_n185_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n615_), .B(mai_mai_n115_), .Y(mai_mai_n616_));
  AN2        m594(.A(mai_mai_n616_), .B(mai_mai_n499_), .Y(mai_mai_n617_));
  NO2        m595(.A(mai_mai_n225_), .B(mai_mai_n45_), .Y(mai_mai_n618_));
  NO3        m596(.A(mai_mai_n618_), .B(mai_mai_n286_), .C(mai_mai_n230_), .Y(mai_mai_n619_));
  NO2        m597(.A(mai_mai_n117_), .B(mai_mai_n37_), .Y(mai_mai_n620_));
  NO2        m598(.A(mai_mai_n620_), .B(i_6_), .Y(mai_mai_n621_));
  NO2        m599(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n622_));
  NO2        m600(.A(mai_mai_n622_), .B(mai_mai_n64_), .Y(mai_mai_n623_));
  NO2        m601(.A(mai_mai_n623_), .B(mai_mai_n583_), .Y(mai_mai_n624_));
  NO4        m602(.A(mai_mai_n624_), .B(mai_mai_n621_), .C(mai_mai_n619_), .D(i_4_), .Y(mai_mai_n625_));
  NA2        m603(.A(i_1_), .B(i_3_), .Y(mai_mai_n626_));
  NO2        m604(.A(mai_mai_n417_), .B(mai_mai_n94_), .Y(mai_mai_n627_));
  AOI210     m605(.A0(mai_mai_n618_), .A1(mai_mai_n531_), .B0(mai_mai_n627_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n628_), .B(mai_mai_n626_), .Y(mai_mai_n629_));
  NO3        m607(.A(mai_mai_n629_), .B(mai_mai_n625_), .C(mai_mai_n617_), .Y(mai_mai_n630_));
  NA4        m608(.A(mai_mai_n630_), .B(mai_mai_n614_), .C(mai_mai_n608_), .D(mai_mai_n587_), .Y(mai_mai_n631_));
  NO3        m609(.A(mai_mai_n435_), .B(i_3_), .C(i_7_), .Y(mai_mai_n632_));
  NOi21      m610(.An(mai_mai_n632_), .B(i_10_), .Y(mai_mai_n633_));
  OA210      m611(.A0(mai_mai_n633_), .A1(mai_mai_n237_), .B0(mai_mai_n87_), .Y(mai_mai_n634_));
  NA2        m612(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n635_));
  NA3        m613(.A(mai_mai_n159_), .B(mai_mai_n85_), .C(mai_mai_n87_), .Y(mai_mai_n636_));
  NA2        m614(.A(mai_mai_n636_), .B(mai_mai_n635_), .Y(mai_mai_n637_));
  OAI210     m615(.A0(mai_mai_n637_), .A1(mai_mai_n634_), .B0(i_1_), .Y(mai_mai_n638_));
  AOI210     m616(.A0(mai_mai_n251_), .A1(mai_mai_n99_), .B0(i_1_), .Y(mai_mai_n639_));
  NO2        m617(.A(mai_mai_n346_), .B(i_2_), .Y(mai_mai_n640_));
  NA2        m618(.A(mai_mai_n640_), .B(mai_mai_n639_), .Y(mai_mai_n641_));
  OAI210     m619(.A0(mai_mai_n602_), .A1(mai_mai_n411_), .B0(mai_mai_n641_), .Y(mai_mai_n642_));
  INV        m620(.A(mai_mai_n642_), .Y(mai_mai_n643_));
  AOI210     m621(.A0(mai_mai_n643_), .A1(mai_mai_n638_), .B0(i_13_), .Y(mai_mai_n644_));
  OR2        m622(.A(i_11_), .B(i_7_), .Y(mai_mai_n645_));
  NA3        m623(.A(mai_mai_n645_), .B(mai_mai_n107_), .C(mai_mai_n136_), .Y(mai_mai_n646_));
  AOI220     m624(.A0(mai_mai_n430_), .A1(mai_mai_n159_), .B0(i_2_), .B1(mai_mai_n136_), .Y(mai_mai_n647_));
  OAI210     m625(.A0(mai_mai_n647_), .A1(mai_mai_n45_), .B0(mai_mai_n646_), .Y(mai_mai_n648_));
  NO2        m626(.A(mai_mai_n55_), .B(i_12_), .Y(mai_mai_n649_));
  NO2        m627(.A(mai_mai_n436_), .B(mai_mai_n24_), .Y(mai_mai_n650_));
  AOI220     m628(.A0(mai_mai_n650_), .A1(mai_mai_n613_), .B0(mai_mai_n237_), .B1(mai_mai_n129_), .Y(mai_mai_n651_));
  OAI220     m629(.A0(mai_mai_n651_), .A1(mai_mai_n41_), .B0(mai_mai_n971_), .B1(mai_mai_n94_), .Y(mai_mai_n652_));
  AOI210     m630(.A0(mai_mai_n648_), .A1(mai_mai_n305_), .B0(mai_mai_n652_), .Y(mai_mai_n653_));
  INV        m631(.A(mai_mai_n115_), .Y(mai_mai_n654_));
  AOI220     m632(.A0(mai_mai_n654_), .A1(mai_mai_n73_), .B0(mai_mai_n360_), .B1(mai_mai_n599_), .Y(mai_mai_n655_));
  NO2        m633(.A(mai_mai_n655_), .B(mai_mai_n235_), .Y(mai_mai_n656_));
  NA2        m634(.A(mai_mai_n125_), .B(i_13_), .Y(mai_mai_n657_));
  NO2        m635(.A(mai_mai_n598_), .B(mai_mai_n115_), .Y(mai_mai_n658_));
  INV        m636(.A(mai_mai_n658_), .Y(mai_mai_n659_));
  OAI220     m637(.A0(mai_mai_n659_), .A1(mai_mai_n72_), .B0(mai_mai_n657_), .B1(mai_mai_n639_), .Y(mai_mai_n660_));
  NA2        m638(.A(mai_mai_n26_), .B(mai_mai_n185_), .Y(mai_mai_n661_));
  NA2        m639(.A(mai_mai_n661_), .B(i_7_), .Y(mai_mai_n662_));
  NO3        m640(.A(mai_mai_n436_), .B(mai_mai_n229_), .C(mai_mai_n87_), .Y(mai_mai_n663_));
  NA2        m641(.A(mai_mai_n663_), .B(mai_mai_n662_), .Y(mai_mai_n664_));
  NA2        m642(.A(mai_mai_n93_), .B(mai_mai_n103_), .Y(mai_mai_n665_));
  OAI220     m643(.A0(mai_mai_n665_), .A1(mai_mai_n555_), .B0(mai_mai_n664_), .B1(mai_mai_n569_), .Y(mai_mai_n666_));
  NO3        m644(.A(mai_mai_n666_), .B(mai_mai_n660_), .C(mai_mai_n656_), .Y(mai_mai_n667_));
  OR2        m645(.A(i_11_), .B(i_6_), .Y(mai_mai_n668_));
  NA3        m646(.A(mai_mai_n554_), .B(mai_mai_n661_), .C(i_7_), .Y(mai_mai_n669_));
  AOI210     m647(.A0(mai_mai_n669_), .A1(mai_mai_n659_), .B0(mai_mai_n668_), .Y(mai_mai_n670_));
  NA3        m648(.A(mai_mai_n376_), .B(mai_mai_n559_), .C(mai_mai_n99_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n590_), .B(i_13_), .Y(mai_mai_n672_));
  NAi21      m650(.An(i_11_), .B(i_12_), .Y(mai_mai_n673_));
  NOi41      m651(.An(mai_mai_n112_), .B(mai_mai_n673_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n674_));
  NO3        m652(.A(mai_mai_n436_), .B(mai_mai_n539_), .C(mai_mai_n560_), .Y(mai_mai_n675_));
  AOI210     m653(.A0(mai_mai_n675_), .A1(mai_mai_n290_), .B0(mai_mai_n674_), .Y(mai_mai_n676_));
  NA3        m654(.A(mai_mai_n676_), .B(mai_mai_n672_), .C(mai_mai_n671_), .Y(mai_mai_n677_));
  OAI210     m655(.A0(mai_mai_n677_), .A1(mai_mai_n670_), .B0(mai_mai_n64_), .Y(mai_mai_n678_));
  NO2        m656(.A(i_2_), .B(i_12_), .Y(mai_mai_n679_));
  NA2        m657(.A(mai_mai_n345_), .B(mai_mai_n679_), .Y(mai_mai_n680_));
  NO3        m658(.A(i_9_), .B(i_3_), .C(mai_mai_n554_), .Y(mai_mai_n681_));
  NA2        m659(.A(mai_mai_n681_), .B(mai_mai_n345_), .Y(mai_mai_n682_));
  NA2        m660(.A(mai_mai_n682_), .B(mai_mai_n680_), .Y(mai_mai_n683_));
  NA3        m661(.A(mai_mai_n683_), .B(mai_mai_n46_), .C(mai_mai_n217_), .Y(mai_mai_n684_));
  NA4        m662(.A(mai_mai_n684_), .B(mai_mai_n678_), .C(mai_mai_n667_), .D(mai_mai_n653_), .Y(mai_mai_n685_));
  OR4        m663(.A(mai_mai_n685_), .B(mai_mai_n644_), .C(mai_mai_n631_), .D(mai_mai_n572_), .Y(mai5));
  NA2        m664(.A(mai_mai_n610_), .B(mai_mai_n254_), .Y(mai_mai_n687_));
  AN2        m665(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n688_));
  NA3        m666(.A(mai_mai_n688_), .B(mai_mai_n679_), .C(mai_mai_n109_), .Y(mai_mai_n689_));
  NO2        m667(.A(mai_mai_n555_), .B(i_11_), .Y(mai_mai_n690_));
  NA2        m668(.A(mai_mai_n88_), .B(mai_mai_n690_), .Y(mai_mai_n691_));
  NA3        m669(.A(mai_mai_n691_), .B(mai_mai_n689_), .C(mai_mai_n687_), .Y(mai_mai_n692_));
  NO3        m670(.A(i_11_), .B(mai_mai_n229_), .C(i_13_), .Y(mai_mai_n693_));
  NO2        m671(.A(mai_mai_n122_), .B(mai_mai_n23_), .Y(mai_mai_n694_));
  NA2        m672(.A(i_12_), .B(i_8_), .Y(mai_mai_n695_));
  OAI210     m673(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n695_), .Y(mai_mai_n696_));
  INV        m674(.A(mai_mai_n410_), .Y(mai_mai_n697_));
  AOI220     m675(.A0(mai_mai_n293_), .A1(mai_mai_n535_), .B0(mai_mai_n696_), .B1(mai_mai_n694_), .Y(mai_mai_n698_));
  INV        m676(.A(mai_mai_n698_), .Y(mai_mai_n699_));
  NO2        m677(.A(mai_mai_n699_), .B(mai_mai_n692_), .Y(mai_mai_n700_));
  INV        m678(.A(mai_mai_n166_), .Y(mai_mai_n701_));
  INV        m679(.A(mai_mai_n237_), .Y(mai_mai_n702_));
  OAI210     m680(.A0(mai_mai_n640_), .A1(mai_mai_n412_), .B0(mai_mai_n112_), .Y(mai_mai_n703_));
  AOI210     m681(.A0(mai_mai_n703_), .A1(mai_mai_n702_), .B0(mai_mai_n701_), .Y(mai_mai_n704_));
  NO2        m682(.A(mai_mai_n417_), .B(mai_mai_n26_), .Y(mai_mai_n705_));
  NO2        m683(.A(mai_mai_n705_), .B(mai_mai_n387_), .Y(mai_mai_n706_));
  NA2        m684(.A(mai_mai_n706_), .B(i_2_), .Y(mai_mai_n707_));
  INV        m685(.A(mai_mai_n707_), .Y(mai_mai_n708_));
  AOI210     m686(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n383_), .Y(mai_mai_n709_));
  AOI210     m687(.A0(mai_mai_n709_), .A1(mai_mai_n708_), .B0(mai_mai_n704_), .Y(mai_mai_n710_));
  NO2        m688(.A(mai_mai_n182_), .B(mai_mai_n123_), .Y(mai_mai_n711_));
  OAI210     m689(.A0(mai_mai_n711_), .A1(mai_mai_n694_), .B0(i_2_), .Y(mai_mai_n712_));
  INV        m690(.A(mai_mai_n167_), .Y(mai_mai_n713_));
  NO3        m691(.A(mai_mai_n574_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n714_));
  AOI210     m692(.A0(mai_mai_n713_), .A1(mai_mai_n88_), .B0(mai_mai_n714_), .Y(mai_mai_n715_));
  AOI210     m693(.A0(mai_mai_n715_), .A1(mai_mai_n712_), .B0(mai_mai_n185_), .Y(mai_mai_n716_));
  OA210      m694(.A0(mai_mai_n575_), .A1(mai_mai_n124_), .B0(i_13_), .Y(mai_mai_n717_));
  NA2        m695(.A(mai_mai_n192_), .B(mai_mai_n195_), .Y(mai_mai_n718_));
  NA2        m696(.A(mai_mai_n150_), .B(mai_mai_n552_), .Y(mai_mai_n719_));
  AOI210     m697(.A0(mai_mai_n719_), .A1(mai_mai_n718_), .B0(mai_mai_n350_), .Y(mai_mai_n720_));
  AOI210     m698(.A0(mai_mai_n200_), .A1(mai_mai_n146_), .B0(mai_mai_n475_), .Y(mai_mai_n721_));
  NA2        m699(.A(mai_mai_n721_), .B(mai_mai_n387_), .Y(mai_mai_n722_));
  NO2        m700(.A(mai_mai_n103_), .B(mai_mai_n45_), .Y(mai_mai_n723_));
  INV        m701(.A(mai_mai_n279_), .Y(mai_mai_n724_));
  NA4        m702(.A(mai_mai_n724_), .B(mai_mai_n283_), .C(mai_mai_n122_), .D(mai_mai_n43_), .Y(mai_mai_n725_));
  OAI210     m703(.A0(mai_mai_n725_), .A1(mai_mai_n723_), .B0(mai_mai_n722_), .Y(mai_mai_n726_));
  NO4        m704(.A(mai_mai_n726_), .B(mai_mai_n720_), .C(mai_mai_n717_), .D(mai_mai_n716_), .Y(mai_mai_n727_));
  NA2        m705(.A(mai_mai_n535_), .B(mai_mai_n28_), .Y(mai_mai_n728_));
  NA2        m706(.A(mai_mai_n693_), .B(mai_mai_n261_), .Y(mai_mai_n729_));
  NA2        m707(.A(mai_mai_n729_), .B(mai_mai_n728_), .Y(mai_mai_n730_));
  NO2        m708(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n731_));
  NO2        m709(.A(mai_mai_n731_), .B(mai_mai_n124_), .Y(mai_mai_n732_));
  NO2        m710(.A(mai_mai_n732_), .B(mai_mai_n552_), .Y(mai_mai_n733_));
  AOI220     m711(.A0(mai_mai_n733_), .A1(mai_mai_n36_), .B0(mai_mai_n730_), .B1(mai_mai_n47_), .Y(mai_mai_n734_));
  NA4        m712(.A(mai_mai_n734_), .B(mai_mai_n727_), .C(mai_mai_n710_), .D(mai_mai_n700_), .Y(mai6));
  NA4        m713(.A(mai_mai_n362_), .B(mai_mai_n441_), .C(mai_mai_n72_), .D(mai_mai_n102_), .Y(mai_mai_n736_));
  INV        m714(.A(mai_mai_n736_), .Y(mai_mai_n737_));
  NO2        m715(.A(mai_mai_n213_), .B(mai_mai_n446_), .Y(mai_mai_n738_));
  NO2        m716(.A(i_11_), .B(i_9_), .Y(mai_mai_n739_));
  NO2        m717(.A(mai_mai_n737_), .B(mai_mai_n304_), .Y(mai_mai_n740_));
  OR2        m718(.A(mai_mai_n740_), .B(i_12_), .Y(mai_mai_n741_));
  NA2        m719(.A(mai_mai_n351_), .B(mai_mai_n308_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n539_), .B(mai_mai_n64_), .Y(mai_mai_n743_));
  NA2        m721(.A(mai_mai_n633_), .B(mai_mai_n72_), .Y(mai_mai_n744_));
  NA3        m722(.A(mai_mai_n744_), .B(mai_mai_n743_), .C(mai_mai_n742_), .Y(mai_mai_n745_));
  INV        m723(.A(mai_mai_n189_), .Y(mai_mai_n746_));
  AOI220     m724(.A0(mai_mai_n746_), .A1(mai_mai_n739_), .B0(mai_mai_n745_), .B1(mai_mai_n74_), .Y(mai_mai_n747_));
  INV        m725(.A(mai_mai_n303_), .Y(mai_mai_n748_));
  NA2        m726(.A(mai_mai_n76_), .B(mai_mai_n129_), .Y(mai_mai_n749_));
  INV        m727(.A(mai_mai_n122_), .Y(mai_mai_n750_));
  NA2        m728(.A(mai_mai_n750_), .B(mai_mai_n47_), .Y(mai_mai_n751_));
  AOI210     m729(.A0(mai_mai_n751_), .A1(mai_mai_n749_), .B0(mai_mai_n748_), .Y(mai_mai_n752_));
  NO2        m730(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n753_));
  NA3        m731(.A(mai_mai_n753_), .B(mai_mai_n432_), .C(mai_mai_n362_), .Y(mai_mai_n754_));
  NAi32      m732(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n755_));
  NO2        m733(.A(mai_mai_n668_), .B(mai_mai_n755_), .Y(mai_mai_n756_));
  OAI210     m734(.A0(mai_mai_n632_), .A1(mai_mai_n523_), .B0(mai_mai_n522_), .Y(mai_mai_n757_));
  NAi31      m735(.An(mai_mai_n756_), .B(mai_mai_n757_), .C(mai_mai_n754_), .Y(mai_mai_n758_));
  OR2        m736(.A(mai_mai_n758_), .B(mai_mai_n752_), .Y(mai_mai_n759_));
  NO2        m737(.A(mai_mai_n645_), .B(i_2_), .Y(mai_mai_n760_));
  NA2        m738(.A(mai_mai_n49_), .B(mai_mai_n37_), .Y(mai_mai_n761_));
  NO2        m739(.A(mai_mai_n761_), .B(mai_mai_n375_), .Y(mai_mai_n762_));
  NA2        m740(.A(mai_mai_n762_), .B(mai_mai_n760_), .Y(mai_mai_n763_));
  AO210      m741(.A0(mai_mai_n334_), .A1(mai_mai_n324_), .B0(mai_mai_n364_), .Y(mai_mai_n764_));
  NA3        m742(.A(mai_mai_n764_), .B(mai_mai_n247_), .C(i_7_), .Y(mai_mai_n765_));
  BUFFER     m743(.A(mai_mai_n575_), .Y(mai_mai_n766_));
  NA3        m744(.A(mai_mai_n766_), .B(mai_mai_n145_), .C(mai_mai_n70_), .Y(mai_mai_n767_));
  OR2        m745(.A(mai_mai_n697_), .B(mai_mai_n36_), .Y(mai_mai_n768_));
  NA4        m746(.A(mai_mai_n768_), .B(mai_mai_n767_), .C(mai_mai_n765_), .D(mai_mai_n763_), .Y(mai_mai_n769_));
  NO2        m747(.A(i_6_), .B(i_11_), .Y(mai_mai_n770_));
  AOI220     m748(.A0(mai_mai_n770_), .A1(mai_mai_n522_), .B0(mai_mai_n738_), .B1(mai_mai_n662_), .Y(mai_mai_n771_));
  NA3        m749(.A(mai_mai_n350_), .B(mai_mai_n231_), .C(mai_mai_n145_), .Y(mai_mai_n772_));
  NA2        m750(.A(mai_mai_n364_), .B(mai_mai_n71_), .Y(mai_mai_n773_));
  NA4        m751(.A(mai_mai_n773_), .B(mai_mai_n772_), .C(mai_mai_n771_), .D(mai_mai_n558_), .Y(mai_mai_n774_));
  AOI210     m752(.A0(mai_mai_n412_), .A1(mai_mai_n410_), .B0(mai_mai_n521_), .Y(mai_mai_n775_));
  NO2        m753(.A(mai_mai_n565_), .B(mai_mai_n103_), .Y(mai_mai_n776_));
  OAI210     m754(.A0(mai_mai_n776_), .A1(mai_mai_n113_), .B0(mai_mai_n373_), .Y(mai_mai_n777_));
  INV        m755(.A(mai_mai_n545_), .Y(mai_mai_n778_));
  NA3        m756(.A(mai_mai_n778_), .B(mai_mai_n303_), .C(i_7_), .Y(mai_mai_n779_));
  NA3        m757(.A(mai_mai_n779_), .B(mai_mai_n777_), .C(mai_mai_n775_), .Y(mai_mai_n780_));
  NO4        m758(.A(mai_mai_n780_), .B(mai_mai_n774_), .C(mai_mai_n769_), .D(mai_mai_n759_), .Y(mai_mai_n781_));
  NA4        m759(.A(mai_mai_n781_), .B(mai_mai_n747_), .C(mai_mai_n741_), .D(mai_mai_n357_), .Y(mai3));
  NA2        m760(.A(i_12_), .B(i_10_), .Y(mai_mai_n783_));
  NA2        m761(.A(i_6_), .B(i_7_), .Y(mai_mai_n784_));
  NO2        m762(.A(mai_mai_n784_), .B(i_0_), .Y(mai_mai_n785_));
  NO2        m763(.A(i_11_), .B(mai_mai_n229_), .Y(mai_mai_n786_));
  NA2        m764(.A(mai_mai_n272_), .B(mai_mai_n786_), .Y(mai_mai_n787_));
  NO2        m765(.A(mai_mai_n787_), .B(mai_mai_n185_), .Y(mai_mai_n788_));
  NO3        m766(.A(mai_mai_n413_), .B(mai_mai_n91_), .C(mai_mai_n45_), .Y(mai_mai_n789_));
  OA210      m767(.A0(mai_mai_n789_), .A1(mai_mai_n788_), .B0(mai_mai_n169_), .Y(mai_mai_n790_));
  NA2        m768(.A(mai_mai_n772_), .B(mai_mai_n349_), .Y(mai_mai_n791_));
  NA2        m769(.A(mai_mai_n791_), .B(mai_mai_n40_), .Y(mai_mai_n792_));
  NOi21      m770(.An(mai_mai_n98_), .B(mai_mai_n706_), .Y(mai_mai_n793_));
  NA2        m771(.A(mai_mai_n376_), .B(mai_mai_n46_), .Y(mai_mai_n794_));
  AN2        m772(.A(mai_mai_n415_), .B(mai_mai_n56_), .Y(mai_mai_n795_));
  NO2        m773(.A(mai_mai_n795_), .B(mai_mai_n793_), .Y(mai_mai_n796_));
  AOI210     m774(.A0(mai_mai_n796_), .A1(mai_mai_n792_), .B0(mai_mai_n49_), .Y(mai_mai_n797_));
  NO4        m775(.A(mai_mai_n353_), .B(mai_mai_n359_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n798_));
  NA2        m776(.A(mai_mai_n177_), .B(mai_mai_n531_), .Y(mai_mai_n799_));
  NOi21      m777(.An(mai_mai_n799_), .B(mai_mai_n798_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n800_), .B(mai_mai_n64_), .Y(mai_mai_n801_));
  NOi21      m779(.An(i_5_), .B(i_9_), .Y(mai_mai_n802_));
  NA2        m780(.A(mai_mai_n802_), .B(mai_mai_n409_), .Y(mai_mai_n803_));
  BUFFER     m781(.A(mai_mai_n251_), .Y(mai_mai_n804_));
  NA2        m782(.A(mai_mai_n804_), .B(mai_mai_n434_), .Y(mai_mai_n805_));
  NO3        m783(.A(mai_mai_n379_), .B(mai_mai_n251_), .C(mai_mai_n74_), .Y(mai_mai_n806_));
  NO2        m784(.A(mai_mai_n170_), .B(mai_mai_n146_), .Y(mai_mai_n807_));
  AOI210     m785(.A0(mai_mai_n807_), .A1(mai_mai_n236_), .B0(mai_mai_n806_), .Y(mai_mai_n808_));
  OAI220     m786(.A0(mai_mai_n808_), .A1(mai_mai_n175_), .B0(mai_mai_n805_), .B1(mai_mai_n803_), .Y(mai_mai_n809_));
  NO4        m787(.A(mai_mai_n809_), .B(mai_mai_n801_), .C(mai_mai_n797_), .D(mai_mai_n790_), .Y(mai_mai_n810_));
  NA2        m788(.A(mai_mai_n177_), .B(mai_mai_n24_), .Y(mai_mai_n811_));
  NO2        m789(.A(mai_mai_n362_), .B(mai_mai_n273_), .Y(mai_mai_n812_));
  NA2        m790(.A(mai_mai_n812_), .B(mai_mai_n658_), .Y(mai_mai_n813_));
  NA2        m791(.A(mai_mai_n532_), .B(i_0_), .Y(mai_mai_n814_));
  NO4        m792(.A(mai_mai_n544_), .B(mai_mai_n207_), .C(mai_mai_n383_), .D(mai_mai_n375_), .Y(mai_mai_n815_));
  NA2        m793(.A(mai_mai_n815_), .B(i_11_), .Y(mai_mai_n816_));
  NA2        m794(.A(mai_mai_n693_), .B(mai_mai_n304_), .Y(mai_mai_n817_));
  AOI210     m795(.A0(mai_mai_n442_), .A1(mai_mai_n88_), .B0(mai_mai_n59_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n818_), .B(mai_mai_n817_), .Y(mai_mai_n819_));
  INV        m797(.A(mai_mai_n498_), .Y(mai_mai_n820_));
  NO4        m798(.A(mai_mai_n115_), .B(mai_mai_n59_), .C(mai_mai_n615_), .D(i_5_), .Y(mai_mai_n821_));
  AN2        m799(.A(mai_mai_n821_), .B(mai_mai_n820_), .Y(mai_mai_n822_));
  AOI220     m800(.A0(mai_mai_n306_), .A1(mai_mai_n100_), .B0(mai_mai_n177_), .B1(mai_mai_n85_), .Y(mai_mai_n823_));
  NA2        m801(.A(mai_mai_n526_), .B(i_4_), .Y(mai_mai_n824_));
  NO2        m802(.A(mai_mai_n824_), .B(mai_mai_n823_), .Y(mai_mai_n825_));
  NO3        m803(.A(mai_mai_n825_), .B(mai_mai_n822_), .C(mai_mai_n819_), .Y(mai_mai_n826_));
  NA3        m804(.A(mai_mai_n826_), .B(mai_mai_n816_), .C(mai_mai_n813_), .Y(mai_mai_n827_));
  NO2        m805(.A(mai_mai_n104_), .B(mai_mai_n37_), .Y(mai_mai_n828_));
  NA2        m806(.A(i_11_), .B(i_9_), .Y(mai_mai_n829_));
  NO3        m807(.A(i_12_), .B(mai_mai_n829_), .C(mai_mai_n557_), .Y(mai_mai_n830_));
  AN2        m808(.A(mai_mai_n830_), .B(mai_mai_n828_), .Y(mai_mai_n831_));
  NO2        m809(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n832_));
  NA2        m810(.A(mai_mai_n363_), .B(mai_mai_n174_), .Y(mai_mai_n833_));
  INV        m811(.A(mai_mai_n833_), .Y(mai_mai_n834_));
  NO2        m812(.A(mai_mai_n829_), .B(mai_mai_n74_), .Y(mai_mai_n835_));
  NO2        m813(.A(mai_mai_n170_), .B(i_0_), .Y(mai_mai_n836_));
  INV        m814(.A(mai_mai_n836_), .Y(mai_mai_n837_));
  NA2        m815(.A(mai_mai_n432_), .B(mai_mai_n223_), .Y(mai_mai_n838_));
  AOI210     m816(.A0(mai_mai_n348_), .A1(mai_mai_n42_), .B0(mai_mai_n372_), .Y(mai_mai_n839_));
  OAI220     m817(.A0(mai_mai_n839_), .A1(mai_mai_n803_), .B0(mai_mai_n838_), .B1(mai_mai_n837_), .Y(mai_mai_n840_));
  NO3        m818(.A(mai_mai_n840_), .B(mai_mai_n834_), .C(mai_mai_n831_), .Y(mai_mai_n841_));
  NA2        m819(.A(mai_mai_n606_), .B(mai_mai_n119_), .Y(mai_mai_n842_));
  NO2        m820(.A(i_6_), .B(mai_mai_n842_), .Y(mai_mai_n843_));
  NA2        m821(.A(mai_mai_n166_), .B(mai_mai_n104_), .Y(mai_mai_n844_));
  NA2        m822(.A(mai_mai_n559_), .B(mai_mai_n304_), .Y(mai_mai_n845_));
  NO2        m823(.A(mai_mai_n845_), .B(mai_mai_n794_), .Y(mai_mai_n846_));
  NO2        m824(.A(mai_mai_n846_), .B(mai_mai_n843_), .Y(mai_mai_n847_));
  NOi21      m825(.An(i_7_), .B(i_5_), .Y(mai_mai_n848_));
  NO3        m826(.A(mai_mai_n368_), .B(mai_mai_n337_), .C(mai_mai_n333_), .Y(mai_mai_n849_));
  NO2        m827(.A(mai_mai_n249_), .B(mai_mai_n294_), .Y(mai_mai_n850_));
  INV        m828(.A(mai_mai_n673_), .Y(mai_mai_n851_));
  AOI210     m829(.A0(mai_mai_n851_), .A1(mai_mai_n850_), .B0(mai_mai_n849_), .Y(mai_mai_n852_));
  NA3        m830(.A(mai_mai_n852_), .B(mai_mai_n847_), .C(mai_mai_n841_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n811_), .B(mai_mai_n232_), .Y(mai_mai_n854_));
  AN2        m832(.A(mai_mai_n305_), .B(mai_mai_n304_), .Y(mai_mai_n855_));
  AN2        m833(.A(mai_mai_n855_), .B(mai_mai_n807_), .Y(mai_mai_n856_));
  OAI210     m834(.A0(mai_mai_n856_), .A1(mai_mai_n854_), .B0(i_10_), .Y(mai_mai_n857_));
  NO2        m835(.A(mai_mai_n783_), .B(mai_mai_n293_), .Y(mai_mai_n858_));
  OA210      m836(.A0(mai_mai_n432_), .A1(mai_mai_n216_), .B0(mai_mai_n431_), .Y(mai_mai_n859_));
  NA2        m837(.A(mai_mai_n858_), .B(mai_mai_n835_), .Y(mai_mai_n860_));
  NA2        m838(.A(mai_mai_n835_), .B(mai_mai_n283_), .Y(mai_mai_n861_));
  OAI210     m839(.A0(i_2_), .A1(mai_mai_n179_), .B0(mai_mai_n861_), .Y(mai_mai_n862_));
  NA2        m840(.A(mai_mai_n862_), .B(mai_mai_n432_), .Y(mai_mai_n863_));
  NO3        m841(.A(mai_mai_n544_), .B(mai_mai_n332_), .C(mai_mai_n24_), .Y(mai_mai_n864_));
  AOI210     m842(.A0(mai_mai_n650_), .A1(mai_mai_n503_), .B0(mai_mai_n864_), .Y(mai_mai_n865_));
  NAi21      m843(.An(i_9_), .B(i_5_), .Y(mai_mai_n866_));
  NO2        m844(.A(mai_mai_n866_), .B(mai_mai_n368_), .Y(mai_mai_n867_));
  NO2        m845(.A(mai_mai_n553_), .B(mai_mai_n106_), .Y(mai_mai_n868_));
  AOI220     m846(.A0(mai_mai_n868_), .A1(i_0_), .B0(mai_mai_n867_), .B1(mai_mai_n575_), .Y(mai_mai_n869_));
  OAI220     m847(.A0(mai_mai_n869_), .A1(mai_mai_n87_), .B0(mai_mai_n865_), .B1(mai_mai_n167_), .Y(mai_mai_n870_));
  NO2        m848(.A(mai_mai_n870_), .B(mai_mai_n478_), .Y(mai_mai_n871_));
  NA4        m849(.A(mai_mai_n871_), .B(mai_mai_n863_), .C(mai_mai_n860_), .D(mai_mai_n857_), .Y(mai_mai_n872_));
  NO3        m850(.A(mai_mai_n872_), .B(mai_mai_n853_), .C(mai_mai_n827_), .Y(mai_mai_n873_));
  NO2        m851(.A(i_0_), .B(mai_mai_n673_), .Y(mai_mai_n874_));
  NO3        m852(.A(mai_mai_n106_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n875_));
  AO220      m853(.A0(mai_mai_n875_), .A1(mai_mai_n45_), .B0(mai_mai_n874_), .B1(mai_mai_n169_), .Y(mai_mai_n876_));
  AOI210     m854(.A0(mai_mai_n743_), .A1(mai_mai_n635_), .B0(mai_mai_n844_), .Y(mai_mai_n877_));
  AOI210     m855(.A0(mai_mai_n876_), .A1(mai_mai_n321_), .B0(mai_mai_n877_), .Y(mai_mai_n878_));
  NA2        m856(.A(i_8_), .B(mai_mai_n144_), .Y(mai_mai_n879_));
  INV        m857(.A(mai_mai_n879_), .Y(mai_mai_n880_));
  NA3        m858(.A(mai_mai_n880_), .B(mai_mai_n622_), .C(mai_mai_n74_), .Y(mai_mai_n881_));
  NO2        m859(.A(mai_mai_n757_), .B(mai_mai_n368_), .Y(mai_mai_n882_));
  NA3        m860(.A(mai_mai_n785_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n883_));
  NA2        m861(.A(mai_mai_n786_), .B(i_9_), .Y(mai_mai_n884_));
  AOI210     m862(.A0(mai_mai_n883_), .A1(mai_mai_n457_), .B0(mai_mai_n884_), .Y(mai_mai_n885_));
  OAI210     m863(.A0(mai_mai_n236_), .A1(i_9_), .B0(mai_mai_n222_), .Y(mai_mai_n886_));
  AOI210     m864(.A0(mai_mai_n886_), .A1(mai_mai_n814_), .B0(mai_mai_n152_), .Y(mai_mai_n887_));
  NO3        m865(.A(mai_mai_n887_), .B(mai_mai_n885_), .C(mai_mai_n882_), .Y(mai_mai_n888_));
  NA3        m866(.A(mai_mai_n888_), .B(mai_mai_n881_), .C(mai_mai_n878_), .Y(mai_mai_n889_));
  NA2        m867(.A(mai_mai_n855_), .B(mai_mai_n350_), .Y(mai_mai_n890_));
  AOI210     m868(.A0(mai_mai_n278_), .A1(mai_mai_n160_), .B0(mai_mai_n890_), .Y(mai_mai_n891_));
  NA3        m869(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n892_));
  NA2        m870(.A(mai_mai_n832_), .B(mai_mai_n447_), .Y(mai_mai_n893_));
  AOI210     m871(.A0(mai_mai_n892_), .A1(mai_mai_n160_), .B0(mai_mai_n893_), .Y(mai_mai_n894_));
  NO2        m872(.A(mai_mai_n894_), .B(mai_mai_n891_), .Y(mai_mai_n895_));
  NA2        m873(.A(mai_mai_n527_), .B(mai_mai_n76_), .Y(mai_mai_n896_));
  NO3        m874(.A(mai_mai_n201_), .B(mai_mai_n359_), .C(i_0_), .Y(mai_mai_n897_));
  OAI210     m875(.A0(mai_mai_n897_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n898_));
  INV        m876(.A(mai_mai_n210_), .Y(mai_mai_n899_));
  OAI220     m877(.A0(mai_mai_n491_), .A1(mai_mai_n137_), .B0(mai_mai_n594_), .B1(mai_mai_n569_), .Y(mai_mai_n900_));
  NA3        m878(.A(mai_mai_n900_), .B(i_7_), .C(mai_mai_n899_), .Y(mai_mai_n901_));
  NA4        m879(.A(mai_mai_n901_), .B(mai_mai_n898_), .C(mai_mai_n896_), .D(mai_mai_n895_), .Y(mai_mai_n902_));
  NO2        m880(.A(mai_mai_n235_), .B(mai_mai_n94_), .Y(mai_mai_n903_));
  AOI210     m881(.A0(mai_mai_n903_), .A1(mai_mai_n874_), .B0(mai_mai_n110_), .Y(mai_mai_n904_));
  NA2        m882(.A(mai_mai_n848_), .B(mai_mai_n447_), .Y(mai_mai_n905_));
  NA2        m883(.A(mai_mai_n324_), .B(mai_mai_n171_), .Y(mai_mai_n906_));
  OA220      m884(.A0(mai_mai_n906_), .A1(mai_mai_n905_), .B0(mai_mai_n904_), .B1(i_5_), .Y(mai_mai_n907_));
  AOI210     m885(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n170_), .Y(mai_mai_n908_));
  NA2        m886(.A(mai_mai_n908_), .B(mai_mai_n859_), .Y(mai_mai_n909_));
  NA3        m887(.A(mai_mai_n566_), .B(mai_mai_n177_), .C(mai_mai_n85_), .Y(mai_mai_n910_));
  NA2        m888(.A(mai_mai_n910_), .B(mai_mai_n502_), .Y(mai_mai_n911_));
  NO3        m889(.A(mai_mai_n794_), .B(mai_mai_n55_), .C(mai_mai_n49_), .Y(mai_mai_n912_));
  NA2        m890(.A(mai_mai_n452_), .B(mai_mai_n445_), .Y(mai_mai_n913_));
  NO3        m891(.A(mai_mai_n913_), .B(mai_mai_n912_), .C(mai_mai_n911_), .Y(mai_mai_n914_));
  NA3        m892(.A(mai_mai_n832_), .B(mai_mai_n272_), .C(mai_mai_n222_), .Y(mai_mai_n915_));
  INV        m893(.A(mai_mai_n915_), .Y(mai_mai_n916_));
  NO3        m894(.A(mai_mai_n829_), .B(mai_mai_n210_), .C(mai_mai_n182_), .Y(mai_mai_n917_));
  NO2        m895(.A(mai_mai_n917_), .B(mai_mai_n916_), .Y(mai_mai_n918_));
  NA4        m896(.A(mai_mai_n918_), .B(mai_mai_n914_), .C(mai_mai_n909_), .D(mai_mai_n907_), .Y(mai_mai_n919_));
  INV        m897(.A(mai_mai_n568_), .Y(mai_mai_n920_));
  NO3        m898(.A(mai_mai_n920_), .B(mai_mai_n517_), .C(i_7_), .Y(mai_mai_n921_));
  INV        m899(.A(mai_mai_n921_), .Y(mai_mai_n922_));
  NA3        m900(.A(mai_mai_n283_), .B(i_5_), .C(mai_mai_n185_), .Y(mai_mai_n923_));
  NAi31      m901(.An(mai_mai_n234_), .B(mai_mai_n923_), .C(mai_mai_n235_), .Y(mai_mai_n924_));
  NO4        m902(.A(mai_mai_n232_), .B(mai_mai_n201_), .C(i_0_), .D(i_12_), .Y(mai_mai_n925_));
  AOI220     m903(.A0(mai_mai_n925_), .A1(mai_mai_n924_), .B0(mai_mai_n737_), .B1(mai_mai_n171_), .Y(mai_mai_n926_));
  NA2        m904(.A(mai_mai_n848_), .B(mai_mai_n430_), .Y(mai_mai_n927_));
  OAI220     m905(.A0(i_7_), .A1(mai_mai_n923_), .B0(mai_mai_n927_), .B1(mai_mai_n623_), .Y(mai_mai_n928_));
  NA2        m906(.A(mai_mai_n928_), .B(mai_mai_n836_), .Y(mai_mai_n929_));
  NA3        m907(.A(mai_mai_n929_), .B(mai_mai_n926_), .C(mai_mai_n922_), .Y(mai_mai_n930_));
  NO4        m908(.A(mai_mai_n930_), .B(mai_mai_n919_), .C(mai_mai_n902_), .D(mai_mai_n889_), .Y(mai_mai_n931_));
  OAI210     m909(.A0(mai_mai_n760_), .A1(mai_mai_n753_), .B0(mai_mai_n37_), .Y(mai_mai_n932_));
  NA2        m910(.A(mai_mai_n932_), .B(mai_mai_n564_), .Y(mai_mai_n933_));
  NA2        m911(.A(mai_mai_n933_), .B(mai_mai_n198_), .Y(mai_mai_n934_));
  NA2        m912(.A(mai_mai_n178_), .B(mai_mai_n180_), .Y(mai_mai_n935_));
  AO210      m913(.A0(mai_mai_n645_), .A1(mai_mai_n33_), .B0(mai_mai_n935_), .Y(mai_mai_n936_));
  OAI210     m914(.A0(mai_mai_n568_), .A1(mai_mai_n566_), .B0(mai_mai_n293_), .Y(mai_mai_n937_));
  NAi31      m915(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n938_));
  NO2        m916(.A(mai_mai_n71_), .B(mai_mai_n938_), .Y(mai_mai_n939_));
  INV        m917(.A(mai_mai_n939_), .Y(mai_mai_n940_));
  NA3        m918(.A(mai_mai_n940_), .B(mai_mai_n937_), .C(mai_mai_n936_), .Y(mai_mai_n941_));
  NO2        m919(.A(mai_mai_n423_), .B(mai_mai_n251_), .Y(mai_mai_n942_));
  NO4        m920(.A(mai_mai_n225_), .B(mai_mai_n143_), .C(mai_mai_n626_), .D(mai_mai_n37_), .Y(mai_mai_n943_));
  NO3        m921(.A(mai_mai_n943_), .B(mai_mai_n942_), .C(mai_mai_n815_), .Y(mai_mai_n944_));
  INV        m922(.A(mai_mai_n944_), .Y(mai_mai_n945_));
  AOI210     m923(.A0(mai_mai_n941_), .A1(mai_mai_n49_), .B0(mai_mai_n945_), .Y(mai_mai_n946_));
  AOI210     m924(.A0(mai_mai_n946_), .A1(mai_mai_n934_), .B0(mai_mai_n74_), .Y(mai_mai_n947_));
  NO2        m925(.A(mai_mai_n524_), .B(mai_mai_n356_), .Y(mai_mai_n948_));
  NO2        m926(.A(mai_mai_n948_), .B(mai_mai_n701_), .Y(mai_mai_n949_));
  NA2        m927(.A(mai_mai_n908_), .B(mai_mai_n832_), .Y(mai_mai_n950_));
  NO2        m928(.A(mai_mai_n950_), .B(mai_mai_n626_), .Y(mai_mai_n951_));
  NA2        m929(.A(mai_mai_n249_), .B(mai_mai_n58_), .Y(mai_mai_n952_));
  AOI220     m930(.A0(mai_mai_n952_), .A1(mai_mai_n77_), .B0(mai_mai_n319_), .B1(mai_mai_n246_), .Y(mai_mai_n953_));
  NO2        m931(.A(mai_mai_n953_), .B(mai_mai_n229_), .Y(mai_mai_n954_));
  NA3        m932(.A(mai_mai_n98_), .B(mai_mai_n285_), .C(mai_mai_n31_), .Y(mai_mai_n955_));
  INV        m933(.A(mai_mai_n955_), .Y(mai_mai_n956_));
  NO3        m934(.A(mai_mai_n956_), .B(mai_mai_n954_), .C(mai_mai_n951_), .Y(mai_mai_n957_));
  OAI210     m935(.A0(mai_mai_n253_), .A1(mai_mai_n157_), .B0(mai_mai_n88_), .Y(mai_mai_n958_));
  NA3        m936(.A(mai_mai_n705_), .B(mai_mai_n272_), .C(mai_mai_n81_), .Y(mai_mai_n959_));
  AOI210     m937(.A0(mai_mai_n959_), .A1(mai_mai_n958_), .B0(i_11_), .Y(mai_mai_n960_));
  NO4        m938(.A(mai_mai_n866_), .B(mai_mai_n435_), .C(mai_mai_n245_), .D(mai_mai_n244_), .Y(mai_mai_n961_));
  NO2        m939(.A(mai_mai_n961_), .B(mai_mai_n521_), .Y(mai_mai_n962_));
  INV        m940(.A(mai_mai_n338_), .Y(mai_mai_n963_));
  AOI210     m941(.A0(mai_mai_n963_), .A1(mai_mai_n962_), .B0(mai_mai_n41_), .Y(mai_mai_n964_));
  NO2        m942(.A(mai_mai_n964_), .B(mai_mai_n960_), .Y(mai_mai_n965_));
  OAI210     m943(.A0(mai_mai_n957_), .A1(i_4_), .B0(mai_mai_n965_), .Y(mai_mai_n966_));
  NO3        m944(.A(mai_mai_n966_), .B(mai_mai_n949_), .C(mai_mai_n947_), .Y(mai_mai_n967_));
  NA4        m945(.A(mai_mai_n967_), .B(mai_mai_n931_), .C(mai_mai_n873_), .D(mai_mai_n810_), .Y(mai4));
  INV        m946(.A(mai_mai_n649_), .Y(mai_mai_n971_));
  INV        m947(.A(i_12_), .Y(mai_mai_n972_));
  NAi21      u000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u002(.A(i_9_), .Y(men_men_n25_));
  INV        u003(.A(i_3_), .Y(men_men_n26_));
  NO2        u004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u013(.A(i_4_), .Y(men_men_n36_));
  INV        u014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u018(.A(men_men_n40_), .Y(men_men_n41_));
  NAi31      u019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u020(.A(men_men_n35_), .Y(men1));
  INV        u021(.A(i_11_), .Y(men_men_n44_));
  NO2        u022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u023(.A(i_2_), .Y(men_men_n46_));
  NA2        u024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u025(.A(i_5_), .Y(men_men_n48_));
  NO2        u026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  NA2        u028(.A(i_0_), .B(i_2_), .Y(men_men_n51_));
  NA2        u029(.A(i_7_), .B(i_9_), .Y(men_men_n52_));
  NO2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NA3        u031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n54_));
  NO2        u032(.A(i_1_), .B(i_6_), .Y(men_men_n55_));
  NA2        u033(.A(i_8_), .B(i_7_), .Y(men_men_n56_));
  OAI210     u034(.A0(men_men_n56_), .A1(men_men_n55_), .B0(men_men_n54_), .Y(men_men_n57_));
  NA2        u035(.A(men_men_n57_), .B(i_12_), .Y(men_men_n58_));
  NAi21      u036(.An(i_2_), .B(i_7_), .Y(men_men_n59_));
  INV        u037(.A(i_1_), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n60_), .B(i_6_), .Y(men_men_n61_));
  NA3        u039(.A(men_men_n61_), .B(men_men_n59_), .C(men_men_n31_), .Y(men_men_n62_));
  NA2        u040(.A(i_1_), .B(i_10_), .Y(men_men_n63_));
  NO2        u041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NAi31      u042(.An(men_men_n64_), .B(men_men_n62_), .C(men_men_n58_), .Y(men_men_n65_));
  NA2        u043(.A(men_men_n50_), .B(i_2_), .Y(men_men_n66_));
  AOI210     u044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n67_));
  NA2        u045(.A(i_1_), .B(i_6_), .Y(men_men_n68_));
  NO2        u046(.A(men_men_n68_), .B(men_men_n25_), .Y(men_men_n69_));
  INV        u047(.A(i_0_), .Y(men_men_n70_));
  NAi21      u048(.An(i_5_), .B(i_10_), .Y(men_men_n71_));
  NA2        u049(.A(i_5_), .B(i_9_), .Y(men_men_n72_));
  AOI210     u050(.A0(men_men_n72_), .A1(men_men_n71_), .B0(men_men_n70_), .Y(men_men_n73_));
  NO2        u051(.A(men_men_n73_), .B(men_men_n69_), .Y(men_men_n74_));
  OAI210     u052(.A0(men_men_n67_), .A1(men_men_n66_), .B0(men_men_n74_), .Y(men_men_n75_));
  OAI210     u053(.A0(men_men_n75_), .A1(men_men_n65_), .B0(i_0_), .Y(men_men_n76_));
  NA2        u054(.A(i_12_), .B(i_5_), .Y(men_men_n77_));
  NA2        u055(.A(i_2_), .B(i_8_), .Y(men_men_n78_));
  NO2        u056(.A(i_3_), .B(i_9_), .Y(men_men_n79_));
  NO2        u057(.A(i_3_), .B(i_7_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n79_), .B(men_men_n60_), .Y(men_men_n81_));
  INV        u059(.A(i_6_), .Y(men_men_n82_));
  OR4        u060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n83_));
  INV        u061(.A(men_men_n83_), .Y(men_men_n84_));
  NO2        u062(.A(i_2_), .B(i_7_), .Y(men_men_n85_));
  NO2        u063(.A(men_men_n84_), .B(men_men_n85_), .Y(men_men_n86_));
  NA2        u064(.A(men_men_n81_), .B(men_men_n86_), .Y(men_men_n87_));
  NAi21      u065(.An(i_6_), .B(i_10_), .Y(men_men_n88_));
  NA2        u066(.A(i_6_), .B(i_9_), .Y(men_men_n89_));
  AOI210     u067(.A0(men_men_n89_), .A1(men_men_n88_), .B0(men_men_n60_), .Y(men_men_n90_));
  NA2        u068(.A(i_2_), .B(i_6_), .Y(men_men_n91_));
  INV        u069(.A(men_men_n90_), .Y(men_men_n92_));
  AOI210     u070(.A0(men_men_n92_), .A1(men_men_n87_), .B0(men_men_n77_), .Y(men_men_n93_));
  AN3        u071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n94_));
  NAi21      u072(.An(i_6_), .B(i_11_), .Y(men_men_n95_));
  NO2        u073(.A(i_5_), .B(i_8_), .Y(men_men_n96_));
  NOi21      u074(.An(men_men_n96_), .B(men_men_n95_), .Y(men_men_n97_));
  AOI220     u075(.A0(men_men_n97_), .A1(men_men_n59_), .B0(men_men_n94_), .B1(men_men_n32_), .Y(men_men_n98_));
  INV        u076(.A(i_7_), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n46_), .B(men_men_n99_), .Y(men_men_n100_));
  NO2        u078(.A(i_0_), .B(i_5_), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n101_), .B(men_men_n82_), .Y(men_men_n102_));
  NA2        u080(.A(i_12_), .B(i_3_), .Y(men_men_n103_));
  INV        u081(.A(men_men_n103_), .Y(men_men_n104_));
  NA3        u082(.A(men_men_n104_), .B(men_men_n102_), .C(men_men_n100_), .Y(men_men_n105_));
  NAi21      u083(.An(i_7_), .B(i_11_), .Y(men_men_n106_));
  AN2        u084(.A(i_2_), .B(i_10_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(i_7_), .Y(men_men_n108_));
  OR2        u086(.A(men_men_n77_), .B(men_men_n55_), .Y(men_men_n109_));
  NO2        u087(.A(i_8_), .B(men_men_n99_), .Y(men_men_n110_));
  NO3        u088(.A(men_men_n110_), .B(men_men_n109_), .C(men_men_n108_), .Y(men_men_n111_));
  NA2        u089(.A(i_12_), .B(i_7_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n60_), .B(men_men_n26_), .Y(men_men_n113_));
  NA2        u091(.A(men_men_n113_), .B(i_0_), .Y(men_men_n114_));
  NA2        u092(.A(i_11_), .B(i_12_), .Y(men_men_n115_));
  OAI210     u093(.A0(men_men_n114_), .A1(men_men_n112_), .B0(men_men_n115_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n116_), .B(men_men_n111_), .Y(men_men_n117_));
  NA3        u095(.A(men_men_n117_), .B(men_men_n105_), .C(men_men_n98_), .Y(men_men_n118_));
  NOi21      u096(.An(i_1_), .B(i_5_), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n119_), .B(i_11_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n99_), .B(men_men_n37_), .Y(men_men_n121_));
  NA2        u099(.A(i_7_), .B(men_men_n25_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n123_), .B(men_men_n46_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n89_), .B(men_men_n88_), .Y(men_men_n125_));
  NAi21      u103(.An(i_3_), .B(i_8_), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n126_), .B(men_men_n59_), .Y(men_men_n127_));
  NOi31      u105(.An(men_men_n127_), .B(men_men_n125_), .C(men_men_n124_), .Y(men_men_n128_));
  NO2        u106(.A(i_1_), .B(men_men_n82_), .Y(men_men_n129_));
  NO2        u107(.A(i_6_), .B(i_5_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n130_), .B(i_3_), .Y(men_men_n131_));
  OAI220     u109(.A0(men_men_n131_), .A1(men_men_n106_), .B0(men_men_n128_), .B1(men_men_n120_), .Y(men_men_n132_));
  NO3        u110(.A(men_men_n132_), .B(men_men_n118_), .C(men_men_n93_), .Y(men_men_n133_));
  NA2        u111(.A(men_men_n133_), .B(men_men_n76_), .Y(men2));
  NO2        u112(.A(men_men_n60_), .B(men_men_n37_), .Y(men_men_n135_));
  NA2        u113(.A(i_6_), .B(men_men_n25_), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n136_), .B(men_men_n135_), .Y(men_men_n137_));
  NA4        u115(.A(men_men_n137_), .B(men_men_n74_), .C(men_men_n66_), .D(men_men_n30_), .Y(men0));
  AN2        u116(.A(i_8_), .B(i_7_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n139_), .B(i_6_), .Y(men_men_n140_));
  NO2        u118(.A(i_12_), .B(i_13_), .Y(men_men_n141_));
  NAi21      u119(.An(i_5_), .B(i_11_), .Y(men_men_n142_));
  NOi21      u120(.An(men_men_n141_), .B(men_men_n142_), .Y(men_men_n143_));
  NO2        u121(.A(i_0_), .B(i_1_), .Y(men_men_n144_));
  NA2        u122(.A(i_2_), .B(i_3_), .Y(men_men_n145_));
  NO2        u123(.A(men_men_n145_), .B(i_4_), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n146_), .B(men_men_n143_), .Y(men_men_n147_));
  AN2        u125(.A(men_men_n141_), .B(men_men_n79_), .Y(men_men_n148_));
  NO2        u126(.A(men_men_n148_), .B(men_men_n27_), .Y(men_men_n149_));
  NA2        u127(.A(i_1_), .B(i_5_), .Y(men_men_n150_));
  NO2        u128(.A(men_men_n70_), .B(men_men_n46_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n151_), .B(men_men_n36_), .Y(men_men_n152_));
  NO3        u130(.A(men_men_n152_), .B(men_men_n150_), .C(men_men_n149_), .Y(men_men_n153_));
  OR2        u131(.A(i_0_), .B(i_1_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n154_), .B(men_men_n77_), .C(i_13_), .Y(men_men_n155_));
  NAi32      u133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n156_));
  NAi21      u134(.An(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  NOi21      u135(.An(i_4_), .B(i_10_), .Y(men_men_n158_));
  NA2        u136(.A(men_men_n158_), .B(men_men_n40_), .Y(men_men_n159_));
  NO2        u137(.A(i_3_), .B(i_5_), .Y(men_men_n160_));
  NO3        u138(.A(men_men_n70_), .B(i_2_), .C(i_1_), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n161_), .B(men_men_n160_), .Y(men_men_n162_));
  OAI210     u140(.A0(men_men_n162_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n163_));
  NO2        u141(.A(men_men_n163_), .B(men_men_n153_), .Y(men_men_n164_));
  AOI210     u142(.A0(men_men_n164_), .A1(men_men_n147_), .B0(men_men_n140_), .Y(men_men_n165_));
  NA2        u143(.A(men_men_n70_), .B(i_1_), .Y(men_men_n166_));
  NA2        u144(.A(i_3_), .B(men_men_n48_), .Y(men_men_n167_));
  NOi21      u145(.An(i_4_), .B(i_9_), .Y(men_men_n168_));
  NOi21      u146(.An(i_11_), .B(i_13_), .Y(men_men_n169_));
  NA2        u147(.A(men_men_n169_), .B(men_men_n168_), .Y(men_men_n170_));
  OR2        u148(.A(men_men_n170_), .B(men_men_n167_), .Y(men_men_n171_));
  NO2        u149(.A(i_4_), .B(i_5_), .Y(men_men_n172_));
  NAi21      u150(.An(i_12_), .B(i_11_), .Y(men_men_n173_));
  NO2        u151(.A(men_men_n173_), .B(i_13_), .Y(men_men_n174_));
  NA3        u152(.A(men_men_n174_), .B(men_men_n172_), .C(men_men_n79_), .Y(men_men_n175_));
  AOI210     u153(.A0(men_men_n175_), .A1(men_men_n171_), .B0(men_men_n166_), .Y(men_men_n176_));
  NO2        u154(.A(men_men_n70_), .B(men_men_n60_), .Y(men_men_n177_));
  INV        u155(.A(men_men_n177_), .Y(men_men_n178_));
  NA2        u156(.A(men_men_n36_), .B(i_5_), .Y(men_men_n179_));
  NAi31      u157(.An(men_men_n179_), .B(men_men_n148_), .C(i_11_), .Y(men_men_n180_));
  NA2        u158(.A(i_3_), .B(i_5_), .Y(men_men_n181_));
  OR2        u159(.A(men_men_n181_), .B(men_men_n170_), .Y(men_men_n182_));
  AOI210     u160(.A0(men_men_n182_), .A1(men_men_n180_), .B0(men_men_n178_), .Y(men_men_n183_));
  NO2        u161(.A(men_men_n70_), .B(i_5_), .Y(men_men_n184_));
  NO2        u162(.A(i_13_), .B(i_10_), .Y(men_men_n185_));
  NA3        u163(.A(men_men_n185_), .B(men_men_n184_), .C(men_men_n44_), .Y(men_men_n186_));
  NO2        u164(.A(i_2_), .B(i_1_), .Y(men_men_n187_));
  NA2        u165(.A(men_men_n187_), .B(i_3_), .Y(men_men_n188_));
  NAi21      u166(.An(i_4_), .B(i_12_), .Y(men_men_n189_));
  NO4        u167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n186_), .D(men_men_n25_), .Y(men_men_n190_));
  NO3        u168(.A(men_men_n190_), .B(men_men_n183_), .C(men_men_n176_), .Y(men_men_n191_));
  INV        u169(.A(i_8_), .Y(men_men_n192_));
  NA2        u170(.A(i_8_), .B(i_6_), .Y(men_men_n193_));
  NO3        u171(.A(i_3_), .B(men_men_n82_), .C(men_men_n48_), .Y(men_men_n194_));
  NA2        u172(.A(men_men_n194_), .B(men_men_n110_), .Y(men_men_n195_));
  NO3        u173(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n196_));
  NA3        u174(.A(men_men_n196_), .B(men_men_n40_), .C(men_men_n44_), .Y(men_men_n197_));
  NO3        u175(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n198_));
  OAI210     u176(.A0(men_men_n94_), .A1(i_12_), .B0(men_men_n198_), .Y(men_men_n199_));
  AOI210     u177(.A0(men_men_n199_), .A1(men_men_n197_), .B0(men_men_n195_), .Y(men_men_n200_));
  NO2        u178(.A(i_3_), .B(i_8_), .Y(men_men_n201_));
  NO3        u179(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n202_));
  NA3        u180(.A(men_men_n202_), .B(men_men_n201_), .C(men_men_n40_), .Y(men_men_n203_));
  INV        u181(.A(i_1_), .Y(men_men_n204_));
  NO2        u182(.A(i_13_), .B(i_9_), .Y(men_men_n205_));
  NA3        u183(.A(men_men_n205_), .B(i_6_), .C(men_men_n192_), .Y(men_men_n206_));
  NAi21      u184(.An(i_12_), .B(i_3_), .Y(men_men_n207_));
  OR2        u185(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n44_), .B(i_5_), .Y(men_men_n209_));
  NO3        u187(.A(i_0_), .B(i_2_), .C(men_men_n60_), .Y(men_men_n210_));
  INV        u188(.A(men_men_n210_), .Y(men_men_n211_));
  OAI220     u189(.A0(men_men_n211_), .A1(men_men_n208_), .B0(men_men_n204_), .B1(men_men_n203_), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n212_), .A1(i_7_), .B0(men_men_n200_), .Y(men_men_n213_));
  OAI220     u191(.A0(men_men_n213_), .A1(i_4_), .B0(men_men_n193_), .B1(men_men_n191_), .Y(men_men_n214_));
  NA3        u192(.A(i_13_), .B(men_men_n192_), .C(i_10_), .Y(men_men_n215_));
  NA2        u193(.A(i_0_), .B(i_5_), .Y(men_men_n216_));
  NAi31      u194(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n36_), .B(i_13_), .Y(men_men_n218_));
  NO2        u196(.A(men_men_n70_), .B(men_men_n26_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n46_), .B(men_men_n60_), .Y(men_men_n220_));
  NA3        u198(.A(men_men_n220_), .B(men_men_n219_), .C(men_men_n218_), .Y(men_men_n221_));
  INV        u199(.A(i_13_), .Y(men_men_n222_));
  NO2        u200(.A(i_12_), .B(men_men_n222_), .Y(men_men_n223_));
  NA3        u201(.A(men_men_n223_), .B(men_men_n196_), .C(men_men_n194_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n221_), .A1(men_men_n217_), .B0(men_men_n224_), .Y(men_men_n225_));
  NA2        u203(.A(men_men_n225_), .B(men_men_n139_), .Y(men_men_n226_));
  NO2        u204(.A(i_12_), .B(men_men_n37_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n181_), .B(i_4_), .Y(men_men_n228_));
  NA2        u206(.A(men_men_n228_), .B(men_men_n227_), .Y(men_men_n229_));
  OR2        u207(.A(i_8_), .B(i_7_), .Y(men_men_n230_));
  NO2        u208(.A(men_men_n230_), .B(men_men_n82_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n51_), .B(i_1_), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n232_), .B(men_men_n231_), .Y(men_men_n233_));
  INV        u211(.A(i_12_), .Y(men_men_n234_));
  NO3        u212(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n235_));
  NA2        u213(.A(i_2_), .B(i_1_), .Y(men_men_n236_));
  NO2        u214(.A(men_men_n233_), .B(men_men_n229_), .Y(men_men_n237_));
  NO3        u215(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n238_));
  NAi21      u216(.An(i_4_), .B(i_3_), .Y(men_men_n239_));
  INV        u217(.A(men_men_n72_), .Y(men_men_n240_));
  NO2        u218(.A(i_0_), .B(i_6_), .Y(men_men_n241_));
  NOi41      u219(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n242_));
  NA2        u220(.A(men_men_n242_), .B(men_men_n241_), .Y(men_men_n243_));
  NO2        u221(.A(men_men_n236_), .B(men_men_n181_), .Y(men_men_n244_));
  NAi21      u222(.An(men_men_n243_), .B(men_men_n244_), .Y(men_men_n245_));
  INV        u223(.A(men_men_n245_), .Y(men_men_n246_));
  AOI210     u224(.A0(men_men_n246_), .A1(men_men_n40_), .B0(men_men_n237_), .Y(men_men_n247_));
  NO2        u225(.A(i_11_), .B(men_men_n222_), .Y(men_men_n248_));
  NOi21      u226(.An(i_1_), .B(i_6_), .Y(men_men_n249_));
  NAi21      u227(.An(i_3_), .B(i_7_), .Y(men_men_n250_));
  NA2        u228(.A(men_men_n234_), .B(i_9_), .Y(men_men_n251_));
  OR4        u229(.A(men_men_n251_), .B(men_men_n250_), .C(men_men_n249_), .D(men_men_n184_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n48_), .B(men_men_n25_), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n70_), .B(i_5_), .Y(men_men_n254_));
  NA2        u232(.A(i_3_), .B(i_9_), .Y(men_men_n255_));
  NAi21      u233(.An(i_7_), .B(i_10_), .Y(men_men_n256_));
  NO2        u234(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  NA3        u235(.A(men_men_n257_), .B(men_men_n254_), .C(men_men_n61_), .Y(men_men_n258_));
  NA2        u236(.A(men_men_n258_), .B(men_men_n252_), .Y(men_men_n259_));
  NA3        u237(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n260_));
  INV        u238(.A(men_men_n140_), .Y(men_men_n261_));
  NA2        u239(.A(men_men_n234_), .B(i_13_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n262_), .B(men_men_n72_), .Y(men_men_n263_));
  AOI220     u241(.A0(men_men_n263_), .A1(men_men_n261_), .B0(men_men_n259_), .B1(men_men_n248_), .Y(men_men_n264_));
  NO2        u242(.A(men_men_n230_), .B(men_men_n37_), .Y(men_men_n265_));
  NA2        u243(.A(i_12_), .B(i_6_), .Y(men_men_n266_));
  OR2        u244(.A(i_13_), .B(i_9_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n239_), .B(i_2_), .Y(men_men_n268_));
  NA2        u246(.A(men_men_n248_), .B(i_9_), .Y(men_men_n269_));
  NA2        u247(.A(men_men_n151_), .B(men_men_n60_), .Y(men_men_n270_));
  NO3        u248(.A(i_11_), .B(men_men_n222_), .C(men_men_n25_), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n250_), .B(i_8_), .Y(men_men_n272_));
  NO2        u250(.A(i_6_), .B(men_men_n48_), .Y(men_men_n273_));
  NA3        u251(.A(men_men_n273_), .B(men_men_n272_), .C(men_men_n271_), .Y(men_men_n274_));
  NA3        u252(.A(i_6_), .B(men_men_n265_), .C(men_men_n223_), .Y(men_men_n275_));
  AOI210     u253(.A0(men_men_n275_), .A1(men_men_n274_), .B0(men_men_n270_), .Y(men_men_n276_));
  INV        u254(.A(men_men_n276_), .Y(men_men_n277_));
  NA4        u255(.A(men_men_n277_), .B(men_men_n264_), .C(men_men_n247_), .D(men_men_n226_), .Y(men_men_n278_));
  NO3        u256(.A(i_12_), .B(men_men_n222_), .C(men_men_n37_), .Y(men_men_n279_));
  INV        u257(.A(men_men_n279_), .Y(men_men_n280_));
  NA2        u258(.A(i_8_), .B(men_men_n99_), .Y(men_men_n281_));
  NOi21      u259(.An(men_men_n160_), .B(men_men_n82_), .Y(men_men_n282_));
  NO3        u260(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n283_));
  AOI220     u261(.A0(men_men_n283_), .A1(men_men_n194_), .B0(men_men_n282_), .B1(men_men_n232_), .Y(men_men_n284_));
  NO2        u262(.A(men_men_n284_), .B(men_men_n281_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n236_), .B(i_0_), .Y(men_men_n286_));
  AOI220     u264(.A0(men_men_n286_), .A1(i_8_), .B0(i_1_), .B1(men_men_n139_), .Y(men_men_n287_));
  NA2        u265(.A(men_men_n273_), .B(men_men_n26_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n288_), .B(men_men_n287_), .Y(men_men_n289_));
  NA2        u267(.A(i_0_), .B(i_1_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n290_), .B(i_2_), .Y(men_men_n291_));
  NO2        u269(.A(men_men_n56_), .B(i_6_), .Y(men_men_n292_));
  NA3        u270(.A(men_men_n292_), .B(men_men_n291_), .C(men_men_n160_), .Y(men_men_n293_));
  OAI210     u271(.A0(men_men_n162_), .A1(men_men_n140_), .B0(men_men_n293_), .Y(men_men_n294_));
  NO3        u272(.A(men_men_n294_), .B(men_men_n289_), .C(men_men_n285_), .Y(men_men_n295_));
  NO2        u273(.A(i_3_), .B(i_10_), .Y(men_men_n296_));
  NA3        u274(.A(men_men_n296_), .B(men_men_n40_), .C(men_men_n44_), .Y(men_men_n297_));
  NO2        u275(.A(i_2_), .B(men_men_n99_), .Y(men_men_n298_));
  NA2        u276(.A(i_1_), .B(men_men_n36_), .Y(men_men_n299_));
  NO2        u277(.A(men_men_n299_), .B(i_8_), .Y(men_men_n300_));
  NA2        u278(.A(men_men_n300_), .B(men_men_n298_), .Y(men_men_n301_));
  AN2        u279(.A(i_3_), .B(i_10_), .Y(men_men_n302_));
  NA4        u280(.A(men_men_n302_), .B(men_men_n196_), .C(men_men_n174_), .D(men_men_n172_), .Y(men_men_n303_));
  NO2        u281(.A(i_5_), .B(men_men_n37_), .Y(men_men_n304_));
  NO2        u282(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n305_));
  OR2        u283(.A(men_men_n301_), .B(men_men_n297_), .Y(men_men_n306_));
  OAI220     u284(.A0(men_men_n306_), .A1(i_6_), .B0(men_men_n295_), .B1(men_men_n280_), .Y(men_men_n307_));
  NO4        u285(.A(men_men_n307_), .B(men_men_n278_), .C(men_men_n214_), .D(men_men_n165_), .Y(men_men_n308_));
  NO3        u286(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n309_));
  NO2        u287(.A(men_men_n56_), .B(men_men_n82_), .Y(men_men_n310_));
  NO3        u288(.A(i_6_), .B(men_men_n192_), .C(i_7_), .Y(men_men_n311_));
  INV        u289(.A(men_men_n311_), .Y(men_men_n312_));
  NO2        u290(.A(men_men_n312_), .B(men_men_n167_), .Y(men_men_n313_));
  NO2        u291(.A(i_2_), .B(i_3_), .Y(men_men_n314_));
  OR2        u292(.A(i_0_), .B(i_5_), .Y(men_men_n315_));
  NA2        u293(.A(men_men_n216_), .B(men_men_n315_), .Y(men_men_n316_));
  NA4        u294(.A(men_men_n316_), .B(men_men_n231_), .C(men_men_n314_), .D(i_1_), .Y(men_men_n317_));
  NA3        u295(.A(men_men_n286_), .B(men_men_n282_), .C(men_men_n110_), .Y(men_men_n318_));
  NAi21      u296(.An(i_8_), .B(i_7_), .Y(men_men_n319_));
  NO2        u297(.A(men_men_n319_), .B(i_6_), .Y(men_men_n320_));
  NO2        u298(.A(men_men_n154_), .B(men_men_n46_), .Y(men_men_n321_));
  NA3        u299(.A(men_men_n321_), .B(men_men_n320_), .C(men_men_n160_), .Y(men_men_n322_));
  NA3        u300(.A(men_men_n322_), .B(men_men_n318_), .C(men_men_n317_), .Y(men_men_n323_));
  OAI210     u301(.A0(men_men_n323_), .A1(men_men_n313_), .B0(i_4_), .Y(men_men_n324_));
  NO2        u302(.A(i_12_), .B(i_10_), .Y(men_men_n325_));
  NOi21      u303(.An(i_5_), .B(i_0_), .Y(men_men_n326_));
  NO3        u304(.A(men_men_n299_), .B(men_men_n326_), .C(men_men_n126_), .Y(men_men_n327_));
  NA4        u305(.A(men_men_n80_), .B(men_men_n36_), .C(men_men_n82_), .D(i_8_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n327_), .B(men_men_n325_), .Y(men_men_n329_));
  NO2        u307(.A(i_6_), .B(i_8_), .Y(men_men_n330_));
  NOi21      u308(.An(i_0_), .B(i_2_), .Y(men_men_n331_));
  AN2        u309(.A(men_men_n331_), .B(men_men_n330_), .Y(men_men_n332_));
  NO2        u310(.A(i_1_), .B(i_7_), .Y(men_men_n333_));
  AO220      u311(.A0(men_men_n333_), .A1(men_men_n332_), .B0(men_men_n320_), .B1(men_men_n232_), .Y(men_men_n334_));
  NA3        u312(.A(men_men_n334_), .B(i_4_), .C(i_5_), .Y(men_men_n335_));
  NA3        u313(.A(men_men_n335_), .B(men_men_n329_), .C(men_men_n324_), .Y(men_men_n336_));
  NO3        u314(.A(men_men_n230_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n337_));
  NO3        u315(.A(men_men_n319_), .B(i_2_), .C(i_1_), .Y(men_men_n338_));
  OAI210     u316(.A0(men_men_n338_), .A1(men_men_n337_), .B0(i_6_), .Y(men_men_n339_));
  NA3        u317(.A(men_men_n249_), .B(men_men_n298_), .C(men_men_n192_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n340_), .A1(men_men_n339_), .B0(men_men_n316_), .Y(men_men_n341_));
  NOi21      u319(.An(men_men_n150_), .B(men_men_n102_), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n122_), .Y(men_men_n343_));
  OAI210     u321(.A0(men_men_n343_), .A1(men_men_n341_), .B0(i_3_), .Y(men_men_n344_));
  INV        u322(.A(men_men_n80_), .Y(men_men_n345_));
  NO2        u323(.A(men_men_n290_), .B(men_men_n78_), .Y(men_men_n346_));
  NA2        u324(.A(men_men_n346_), .B(men_men_n130_), .Y(men_men_n347_));
  NO2        u325(.A(men_men_n91_), .B(men_men_n192_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n348_), .B(men_men_n60_), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n349_), .A1(men_men_n347_), .B0(men_men_n345_), .Y(men_men_n350_));
  INV        u328(.A(i_9_), .Y(men_men_n351_));
  NO2        u329(.A(men_men_n350_), .B(men_men_n289_), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n352_), .A1(men_men_n344_), .B0(men_men_n159_), .Y(men_men_n353_));
  AOI210     u331(.A0(men_men_n336_), .A1(men_men_n309_), .B0(men_men_n353_), .Y(men_men_n354_));
  NOi32      u332(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n355_));
  INV        u333(.A(men_men_n355_), .Y(men_men_n356_));
  NAi21      u334(.An(i_1_), .B(i_5_), .Y(men_men_n357_));
  INV        u335(.A(men_men_n243_), .Y(men_men_n358_));
  NAi41      u336(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n359_));
  OAI220     u337(.A0(men_men_n359_), .A1(men_men_n357_), .B0(men_men_n217_), .B1(men_men_n156_), .Y(men_men_n360_));
  AOI210     u338(.A0(men_men_n359_), .A1(men_men_n156_), .B0(men_men_n154_), .Y(men_men_n361_));
  NOi32      u339(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n362_));
  OR2        u340(.A(men_men_n361_), .B(men_men_n360_), .Y(men_men_n363_));
  NO2        u341(.A(i_1_), .B(men_men_n99_), .Y(men_men_n364_));
  NAi21      u342(.An(i_3_), .B(i_4_), .Y(men_men_n365_));
  NO2        u343(.A(men_men_n365_), .B(i_9_), .Y(men_men_n366_));
  AN2        u344(.A(i_6_), .B(i_7_), .Y(men_men_n367_));
  OAI210     u345(.A0(men_men_n367_), .A1(men_men_n364_), .B0(men_men_n366_), .Y(men_men_n368_));
  NA2        u346(.A(i_2_), .B(i_7_), .Y(men_men_n369_));
  NO2        u347(.A(men_men_n365_), .B(i_10_), .Y(men_men_n370_));
  NA3        u348(.A(men_men_n370_), .B(men_men_n369_), .C(men_men_n241_), .Y(men_men_n371_));
  AOI210     u349(.A0(men_men_n371_), .A1(men_men_n368_), .B0(men_men_n184_), .Y(men_men_n372_));
  AOI210     u350(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n187_), .B0(men_men_n370_), .Y(men_men_n374_));
  AOI220     u352(.A0(men_men_n370_), .A1(men_men_n333_), .B0(men_men_n235_), .B1(men_men_n187_), .Y(men_men_n375_));
  AOI210     u353(.A0(men_men_n375_), .A1(men_men_n374_), .B0(i_5_), .Y(men_men_n376_));
  NO4        u354(.A(men_men_n376_), .B(men_men_n372_), .C(men_men_n363_), .D(men_men_n358_), .Y(men_men_n377_));
  NO2        u355(.A(men_men_n377_), .B(men_men_n356_), .Y(men_men_n378_));
  NO2        u356(.A(men_men_n56_), .B(men_men_n25_), .Y(men_men_n379_));
  AN2        u357(.A(i_12_), .B(i_5_), .Y(men_men_n380_));
  NO2        u358(.A(i_4_), .B(men_men_n26_), .Y(men_men_n381_));
  NA2        u359(.A(men_men_n381_), .B(men_men_n380_), .Y(men_men_n382_));
  NO2        u360(.A(i_11_), .B(i_6_), .Y(men_men_n383_));
  NA3        u361(.A(men_men_n383_), .B(men_men_n321_), .C(men_men_n222_), .Y(men_men_n384_));
  NO2        u362(.A(men_men_n384_), .B(men_men_n382_), .Y(men_men_n385_));
  NO2        u363(.A(men_men_n239_), .B(i_5_), .Y(men_men_n386_));
  NO2        u364(.A(i_5_), .B(i_10_), .Y(men_men_n387_));
  NA2        u365(.A(men_men_n141_), .B(men_men_n45_), .Y(men_men_n388_));
  NO2        u366(.A(men_men_n388_), .B(men_men_n239_), .Y(men_men_n389_));
  OAI210     u367(.A0(men_men_n389_), .A1(men_men_n385_), .B0(men_men_n379_), .Y(men_men_n390_));
  NO2        u368(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n391_));
  NA2        u369(.A(men_men_n385_), .B(men_men_n391_), .Y(men_men_n392_));
  NO3        u370(.A(men_men_n82_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n393_));
  NA3        u371(.A(men_men_n296_), .B(men_men_n89_), .C(men_men_n52_), .Y(men_men_n394_));
  NO2        u372(.A(i_11_), .B(i_12_), .Y(men_men_n395_));
  NA2        u373(.A(men_men_n395_), .B(men_men_n36_), .Y(men_men_n396_));
  NO2        u374(.A(men_men_n394_), .B(men_men_n396_), .Y(men_men_n397_));
  NA2        u375(.A(men_men_n387_), .B(men_men_n234_), .Y(men_men_n398_));
  NA3        u376(.A(men_men_n110_), .B(i_4_), .C(i_11_), .Y(men_men_n399_));
  NO2        u377(.A(men_men_n399_), .B(men_men_n217_), .Y(men_men_n400_));
  NAi21      u378(.An(i_13_), .B(i_0_), .Y(men_men_n401_));
  NO2        u379(.A(men_men_n401_), .B(men_men_n236_), .Y(men_men_n402_));
  OAI210     u380(.A0(men_men_n400_), .A1(men_men_n397_), .B0(men_men_n402_), .Y(men_men_n403_));
  NA3        u381(.A(men_men_n403_), .B(men_men_n392_), .C(men_men_n390_), .Y(men_men_n404_));
  NO3        u382(.A(i_1_), .B(i_12_), .C(men_men_n82_), .Y(men_men_n405_));
  NO2        u383(.A(i_0_), .B(i_11_), .Y(men_men_n406_));
  AN2        u384(.A(i_1_), .B(i_6_), .Y(men_men_n407_));
  NOi21      u385(.An(i_2_), .B(i_12_), .Y(men_men_n408_));
  NA2        u386(.A(men_men_n408_), .B(men_men_n407_), .Y(men_men_n409_));
  INV        u387(.A(men_men_n409_), .Y(men_men_n410_));
  NA2        u388(.A(men_men_n139_), .B(i_9_), .Y(men_men_n411_));
  NO2        u389(.A(men_men_n411_), .B(i_4_), .Y(men_men_n412_));
  NA2        u390(.A(men_men_n410_), .B(men_men_n412_), .Y(men_men_n413_));
  NAi21      u391(.An(i_9_), .B(i_4_), .Y(men_men_n414_));
  OR2        u392(.A(i_13_), .B(i_10_), .Y(men_men_n415_));
  NO3        u393(.A(men_men_n415_), .B(men_men_n115_), .C(men_men_n414_), .Y(men_men_n416_));
  NO2        u394(.A(men_men_n99_), .B(men_men_n25_), .Y(men_men_n417_));
  NA2        u395(.A(men_men_n279_), .B(men_men_n417_), .Y(men_men_n418_));
  NA2        u396(.A(men_men_n273_), .B(men_men_n210_), .Y(men_men_n419_));
  OAI220     u397(.A0(men_men_n419_), .A1(men_men_n215_), .B0(men_men_n418_), .B1(men_men_n342_), .Y(men_men_n420_));
  INV        u398(.A(men_men_n420_), .Y(men_men_n421_));
  AOI210     u399(.A0(men_men_n421_), .A1(men_men_n413_), .B0(men_men_n26_), .Y(men_men_n422_));
  NA2        u400(.A(men_men_n318_), .B(men_men_n317_), .Y(men_men_n423_));
  AOI220     u401(.A0(men_men_n292_), .A1(men_men_n283_), .B0(men_men_n286_), .B1(men_men_n310_), .Y(men_men_n424_));
  NO2        u402(.A(men_men_n424_), .B(men_men_n167_), .Y(men_men_n425_));
  NO2        u403(.A(men_men_n181_), .B(men_men_n82_), .Y(men_men_n426_));
  AOI220     u404(.A0(men_men_n426_), .A1(men_men_n291_), .B0(i_6_), .B1(men_men_n210_), .Y(men_men_n427_));
  NO2        u405(.A(men_men_n427_), .B(men_men_n281_), .Y(men_men_n428_));
  NO3        u406(.A(men_men_n428_), .B(men_men_n425_), .C(men_men_n423_), .Y(men_men_n429_));
  NA2        u407(.A(men_men_n194_), .B(men_men_n94_), .Y(men_men_n430_));
  NA3        u408(.A(men_men_n321_), .B(men_men_n160_), .C(men_men_n82_), .Y(men_men_n431_));
  AOI210     u409(.A0(men_men_n431_), .A1(men_men_n430_), .B0(men_men_n319_), .Y(men_men_n432_));
  NA2        u410(.A(men_men_n192_), .B(i_10_), .Y(men_men_n433_));
  NA3        u411(.A(men_men_n254_), .B(men_men_n61_), .C(i_2_), .Y(men_men_n434_));
  NA2        u412(.A(men_men_n292_), .B(men_men_n232_), .Y(men_men_n435_));
  OAI220     u413(.A0(men_men_n435_), .A1(men_men_n181_), .B0(men_men_n434_), .B1(men_men_n433_), .Y(men_men_n436_));
  NO2        u414(.A(i_3_), .B(men_men_n48_), .Y(men_men_n437_));
  NA3        u415(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n437_), .Y(men_men_n438_));
  NA2        u416(.A(men_men_n311_), .B(men_men_n316_), .Y(men_men_n439_));
  OAI210     u417(.A0(men_men_n439_), .A1(men_men_n188_), .B0(men_men_n438_), .Y(men_men_n440_));
  NO3        u418(.A(men_men_n440_), .B(men_men_n436_), .C(men_men_n432_), .Y(men_men_n441_));
  AOI210     u419(.A0(men_men_n441_), .A1(men_men_n429_), .B0(men_men_n269_), .Y(men_men_n442_));
  NO4        u420(.A(men_men_n442_), .B(men_men_n422_), .C(men_men_n404_), .D(men_men_n378_), .Y(men_men_n443_));
  NO2        u421(.A(men_men_n60_), .B(i_4_), .Y(men_men_n444_));
  NO2        u422(.A(men_men_n70_), .B(i_13_), .Y(men_men_n445_));
  NO2        u423(.A(i_10_), .B(i_9_), .Y(men_men_n446_));
  NAi21      u424(.An(i_12_), .B(i_8_), .Y(men_men_n447_));
  NO2        u425(.A(men_men_n447_), .B(i_3_), .Y(men_men_n448_));
  NO2        u426(.A(men_men_n46_), .B(i_4_), .Y(men_men_n449_));
  NA2        u427(.A(men_men_n449_), .B(men_men_n102_), .Y(men_men_n450_));
  NO2        u428(.A(men_men_n450_), .B(men_men_n203_), .Y(men_men_n451_));
  NA2        u429(.A(men_men_n305_), .B(i_0_), .Y(men_men_n452_));
  NO3        u430(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n453_));
  NA2        u431(.A(men_men_n266_), .B(men_men_n95_), .Y(men_men_n454_));
  NA2        u432(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  NA2        u433(.A(i_8_), .B(i_9_), .Y(men_men_n456_));
  NA2        u434(.A(men_men_n248_), .B(men_men_n304_), .Y(men_men_n457_));
  NO3        u435(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n458_));
  INV        u436(.A(men_men_n458_), .Y(men_men_n459_));
  NA3        u437(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n460_));
  NA4        u438(.A(men_men_n142_), .B(men_men_n113_), .C(men_men_n77_), .D(men_men_n23_), .Y(men_men_n461_));
  OAI220     u439(.A0(men_men_n461_), .A1(men_men_n460_), .B0(men_men_n459_), .B1(men_men_n457_), .Y(men_men_n462_));
  NO2        u440(.A(men_men_n462_), .B(men_men_n451_), .Y(men_men_n463_));
  NA2        u441(.A(men_men_n291_), .B(men_men_n106_), .Y(men_men_n464_));
  OR2        u442(.A(men_men_n464_), .B(men_men_n206_), .Y(men_men_n465_));
  BUFFER     u443(.A(men_men_n293_), .Y(men_men_n466_));
  OA220      u444(.A0(men_men_n466_), .A1(men_men_n159_), .B0(men_men_n465_), .B1(men_men_n229_), .Y(men_men_n467_));
  NA2        u445(.A(men_men_n94_), .B(i_13_), .Y(men_men_n468_));
  NA2        u446(.A(men_men_n426_), .B(men_men_n379_), .Y(men_men_n469_));
  NO2        u447(.A(i_2_), .B(i_13_), .Y(men_men_n470_));
  NO2        u448(.A(men_men_n469_), .B(men_men_n468_), .Y(men_men_n471_));
  NO3        u449(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n472_));
  NO2        u450(.A(i_6_), .B(i_7_), .Y(men_men_n473_));
  NA2        u451(.A(men_men_n473_), .B(men_men_n472_), .Y(men_men_n474_));
  NO2        u452(.A(i_11_), .B(i_1_), .Y(men_men_n475_));
  NO2        u453(.A(men_men_n70_), .B(i_3_), .Y(men_men_n476_));
  NOi21      u454(.An(i_2_), .B(i_7_), .Y(men_men_n477_));
  NAi31      u455(.An(i_11_), .B(men_men_n477_), .C(men_men_n476_), .Y(men_men_n478_));
  NO2        u456(.A(men_men_n415_), .B(i_6_), .Y(men_men_n479_));
  NA2        u457(.A(men_men_n479_), .B(men_men_n444_), .Y(men_men_n480_));
  NO2        u458(.A(men_men_n480_), .B(men_men_n478_), .Y(men_men_n481_));
  NO2        u459(.A(i_3_), .B(men_men_n192_), .Y(men_men_n482_));
  NO2        u460(.A(i_6_), .B(i_10_), .Y(men_men_n483_));
  NA4        u461(.A(men_men_n483_), .B(men_men_n309_), .C(men_men_n482_), .D(men_men_n234_), .Y(men_men_n484_));
  NO2        u462(.A(men_men_n484_), .B(men_men_n152_), .Y(men_men_n485_));
  NA2        u463(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n486_));
  NO2        u464(.A(men_men_n154_), .B(i_3_), .Y(men_men_n487_));
  NAi31      u465(.An(men_men_n486_), .B(men_men_n487_), .C(men_men_n223_), .Y(men_men_n488_));
  NA3        u466(.A(men_men_n391_), .B(men_men_n177_), .C(men_men_n146_), .Y(men_men_n489_));
  NA2        u467(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n490_));
  NO4        u468(.A(men_men_n490_), .B(men_men_n485_), .C(men_men_n481_), .D(men_men_n471_), .Y(men_men_n491_));
  NA2        u469(.A(men_men_n458_), .B(men_men_n387_), .Y(men_men_n492_));
  NO2        u470(.A(men_men_n492_), .B(men_men_n221_), .Y(men_men_n493_));
  NAi21      u471(.An(men_men_n215_), .B(men_men_n395_), .Y(men_men_n494_));
  NO2        u472(.A(men_men_n26_), .B(i_5_), .Y(men_men_n495_));
  NO2        u473(.A(i_0_), .B(men_men_n82_), .Y(men_men_n496_));
  NA3        u474(.A(men_men_n496_), .B(men_men_n495_), .C(men_men_n139_), .Y(men_men_n497_));
  OR3        u475(.A(men_men_n299_), .B(men_men_n38_), .C(men_men_n46_), .Y(men_men_n498_));
  NO2        u476(.A(men_men_n498_), .B(men_men_n497_), .Y(men_men_n499_));
  NA2        u477(.A(men_men_n27_), .B(i_10_), .Y(men_men_n500_));
  NA2        u478(.A(men_men_n309_), .B(men_men_n235_), .Y(men_men_n501_));
  OAI220     u479(.A0(men_men_n501_), .A1(men_men_n434_), .B0(men_men_n500_), .B1(men_men_n468_), .Y(men_men_n502_));
  NA4        u480(.A(men_men_n302_), .B(men_men_n220_), .C(men_men_n70_), .D(men_men_n234_), .Y(men_men_n503_));
  NO2        u481(.A(men_men_n503_), .B(men_men_n474_), .Y(men_men_n504_));
  NO4        u482(.A(men_men_n504_), .B(men_men_n502_), .C(men_men_n499_), .D(men_men_n493_), .Y(men_men_n505_));
  NA4        u483(.A(men_men_n505_), .B(men_men_n491_), .C(men_men_n467_), .D(men_men_n463_), .Y(men_men_n506_));
  NA3        u484(.A(men_men_n302_), .B(men_men_n174_), .C(men_men_n172_), .Y(men_men_n507_));
  OAI210     u485(.A0(men_men_n297_), .A1(men_men_n179_), .B0(men_men_n507_), .Y(men_men_n508_));
  BUFFER     u486(.A(men_men_n283_), .Y(men_men_n509_));
  NA2        u487(.A(men_men_n509_), .B(men_men_n508_), .Y(men_men_n510_));
  NA2        u488(.A(men_men_n120_), .B(men_men_n109_), .Y(men_men_n511_));
  AN2        u489(.A(men_men_n511_), .B(men_men_n453_), .Y(men_men_n512_));
  NA2        u490(.A(men_men_n309_), .B(men_men_n161_), .Y(men_men_n513_));
  OAI210     u491(.A0(men_men_n513_), .A1(men_men_n229_), .B0(men_men_n303_), .Y(men_men_n514_));
  AOI220     u492(.A0(men_men_n514_), .A1(men_men_n320_), .B0(men_men_n512_), .B1(men_men_n305_), .Y(men_men_n515_));
  NA2        u493(.A(men_men_n380_), .B(men_men_n222_), .Y(men_men_n516_));
  NA2        u494(.A(men_men_n355_), .B(men_men_n70_), .Y(men_men_n517_));
  NA2        u495(.A(men_men_n367_), .B(men_men_n362_), .Y(men_men_n518_));
  AO210      u496(.A0(men_men_n517_), .A1(men_men_n516_), .B0(men_men_n518_), .Y(men_men_n519_));
  NO2        u497(.A(men_men_n36_), .B(i_8_), .Y(men_men_n520_));
  NAi41      u498(.An(men_men_n517_), .B(men_men_n483_), .C(men_men_n520_), .D(men_men_n46_), .Y(men_men_n521_));
  AOI210     u499(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n416_), .Y(men_men_n522_));
  NA3        u500(.A(men_men_n522_), .B(men_men_n521_), .C(men_men_n519_), .Y(men_men_n523_));
  INV        u501(.A(men_men_n523_), .Y(men_men_n524_));
  NO2        u502(.A(i_7_), .B(men_men_n197_), .Y(men_men_n525_));
  NO2        u503(.A(men_men_n181_), .B(men_men_n82_), .Y(men_men_n526_));
  NA2        u504(.A(men_men_n526_), .B(men_men_n525_), .Y(men_men_n527_));
  NA4        u505(.A(men_men_n527_), .B(men_men_n524_), .C(men_men_n515_), .D(men_men_n510_), .Y(men_men_n528_));
  NA2        u506(.A(men_men_n386_), .B(men_men_n291_), .Y(men_men_n529_));
  OAI210     u507(.A0(men_men_n382_), .A1(men_men_n166_), .B0(men_men_n529_), .Y(men_men_n530_));
  NA2        u508(.A(men_men_n1016_), .B(men_men_n222_), .Y(men_men_n531_));
  NO3        u509(.A(men_men_n1014_), .B(men_men_n531_), .C(men_men_n464_), .Y(men_men_n532_));
  NOi31      u510(.An(men_men_n311_), .B(men_men_n415_), .C(men_men_n38_), .Y(men_men_n533_));
  OAI210     u511(.A0(men_men_n533_), .A1(men_men_n532_), .B0(men_men_n530_), .Y(men_men_n534_));
  NO2        u512(.A(i_8_), .B(i_7_), .Y(men_men_n535_));
  INV        u513(.A(i_5_), .Y(men_men_n536_));
  NA2        u514(.A(men_men_n536_), .B(men_men_n220_), .Y(men_men_n537_));
  AOI220     u515(.A0(men_men_n321_), .A1(men_men_n40_), .B0(men_men_n232_), .B1(men_men_n205_), .Y(men_men_n538_));
  OAI220     u516(.A0(men_men_n538_), .A1(men_men_n181_), .B0(men_men_n537_), .B1(men_men_n239_), .Y(men_men_n539_));
  NA2        u517(.A(men_men_n44_), .B(i_10_), .Y(men_men_n540_));
  NO2        u518(.A(men_men_n540_), .B(i_6_), .Y(men_men_n541_));
  NA3        u519(.A(men_men_n541_), .B(men_men_n539_), .C(men_men_n535_), .Y(men_men_n542_));
  AOI220     u520(.A0(men_men_n426_), .A1(men_men_n321_), .B0(men_men_n244_), .B1(men_men_n241_), .Y(men_men_n543_));
  OAI220     u521(.A0(men_men_n543_), .A1(men_men_n262_), .B0(men_men_n468_), .B1(men_men_n131_), .Y(men_men_n544_));
  NA2        u522(.A(men_men_n544_), .B(men_men_n265_), .Y(men_men_n545_));
  NOi21      u523(.An(men_men_n286_), .B(men_men_n297_), .Y(men_men_n546_));
  NA2        u524(.A(men_men_n546_), .B(men_men_n458_), .Y(men_men_n547_));
  NA4        u525(.A(men_men_n547_), .B(men_men_n545_), .C(men_men_n542_), .D(men_men_n534_), .Y(men_men_n548_));
  NA3        u526(.A(men_men_n216_), .B(men_men_n68_), .C(men_men_n44_), .Y(men_men_n549_));
  NA2        u527(.A(men_men_n279_), .B(men_men_n80_), .Y(men_men_n550_));
  AOI210     u528(.A0(men_men_n549_), .A1(men_men_n347_), .B0(men_men_n550_), .Y(men_men_n551_));
  NA2        u529(.A(men_men_n292_), .B(men_men_n283_), .Y(men_men_n552_));
  NO2        u530(.A(men_men_n552_), .B(men_men_n171_), .Y(men_men_n553_));
  NA2        u531(.A(men_men_n220_), .B(men_men_n219_), .Y(men_men_n554_));
  NA2        u532(.A(men_men_n446_), .B(men_men_n218_), .Y(men_men_n555_));
  NO2        u533(.A(men_men_n554_), .B(men_men_n555_), .Y(men_men_n556_));
  NO3        u534(.A(men_men_n556_), .B(men_men_n553_), .C(men_men_n551_), .Y(men_men_n557_));
  NO4        u535(.A(men_men_n249_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n558_));
  NO3        u536(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n559_));
  NO2        u537(.A(men_men_n230_), .B(men_men_n36_), .Y(men_men_n560_));
  AN2        u538(.A(men_men_n560_), .B(men_men_n559_), .Y(men_men_n561_));
  OA210      u539(.A0(men_men_n561_), .A1(men_men_n558_), .B0(men_men_n355_), .Y(men_men_n562_));
  NO2        u540(.A(men_men_n415_), .B(i_1_), .Y(men_men_n563_));
  NOi31      u541(.An(men_men_n563_), .B(men_men_n454_), .C(men_men_n70_), .Y(men_men_n564_));
  NO2        u542(.A(men_men_n424_), .B(men_men_n175_), .Y(men_men_n565_));
  NO2        u543(.A(men_men_n565_), .B(men_men_n562_), .Y(men_men_n566_));
  NOi21      u544(.An(i_10_), .B(i_6_), .Y(men_men_n567_));
  NO2        u545(.A(men_men_n82_), .B(men_men_n25_), .Y(men_men_n568_));
  NO2        u546(.A(men_men_n112_), .B(men_men_n23_), .Y(men_men_n569_));
  NA2        u547(.A(men_men_n311_), .B(men_men_n161_), .Y(men_men_n570_));
  AOI220     u548(.A0(men_men_n570_), .A1(men_men_n435_), .B0(men_men_n182_), .B1(men_men_n180_), .Y(men_men_n571_));
  NOi21      u549(.An(men_men_n143_), .B(men_men_n328_), .Y(men_men_n572_));
  NO2        u550(.A(men_men_n572_), .B(men_men_n571_), .Y(men_men_n573_));
  NO2        u551(.A(i_12_), .B(men_men_n82_), .Y(men_men_n574_));
  NA2        u552(.A(men_men_n172_), .B(i_0_), .Y(men_men_n575_));
  NO3        u553(.A(men_men_n575_), .B(men_men_n339_), .C(men_men_n297_), .Y(men_men_n576_));
  INV        u554(.A(men_men_n196_), .Y(men_men_n577_));
  NO2        u555(.A(men_men_n577_), .B(men_men_n494_), .Y(men_men_n578_));
  NO2        u556(.A(men_men_n578_), .B(men_men_n576_), .Y(men_men_n579_));
  NA4        u557(.A(men_men_n579_), .B(men_men_n573_), .C(men_men_n566_), .D(men_men_n557_), .Y(men_men_n580_));
  NO4        u558(.A(men_men_n580_), .B(men_men_n548_), .C(men_men_n528_), .D(men_men_n506_), .Y(men_men_n581_));
  NA4        u559(.A(men_men_n581_), .B(men_men_n443_), .C(men_men_n354_), .D(men_men_n308_), .Y(men7));
  NO2        u560(.A(men_men_n91_), .B(men_men_n52_), .Y(men_men_n583_));
  NO2        u561(.A(men_men_n106_), .B(men_men_n88_), .Y(men_men_n584_));
  NA2        u562(.A(men_men_n381_), .B(men_men_n584_), .Y(men_men_n585_));
  NA2        u563(.A(men_men_n483_), .B(men_men_n80_), .Y(men_men_n586_));
  NA2        u564(.A(i_11_), .B(men_men_n192_), .Y(men_men_n587_));
  NA2        u565(.A(men_men_n141_), .B(men_men_n587_), .Y(men_men_n588_));
  OAI210     u566(.A0(men_men_n588_), .A1(men_men_n586_), .B0(men_men_n585_), .Y(men_men_n589_));
  NA3        u567(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n590_));
  NO2        u568(.A(men_men_n234_), .B(i_4_), .Y(men_men_n591_));
  NA2        u569(.A(men_men_n591_), .B(i_8_), .Y(men_men_n592_));
  NO2        u570(.A(men_men_n103_), .B(men_men_n590_), .Y(men_men_n593_));
  NA2        u571(.A(i_2_), .B(men_men_n82_), .Y(men_men_n594_));
  OAI210     u572(.A0(men_men_n85_), .A1(men_men_n201_), .B0(men_men_n202_), .Y(men_men_n595_));
  NO2        u573(.A(i_7_), .B(men_men_n37_), .Y(men_men_n596_));
  NA2        u574(.A(i_4_), .B(i_8_), .Y(men_men_n597_));
  AOI210     u575(.A0(men_men_n597_), .A1(men_men_n302_), .B0(men_men_n596_), .Y(men_men_n598_));
  OAI220     u576(.A0(men_men_n598_), .A1(men_men_n594_), .B0(men_men_n595_), .B1(i_13_), .Y(men_men_n599_));
  NO4        u577(.A(men_men_n599_), .B(men_men_n593_), .C(men_men_n589_), .D(men_men_n583_), .Y(men_men_n600_));
  AOI210     u578(.A0(men_men_n126_), .A1(men_men_n59_), .B0(i_10_), .Y(men_men_n601_));
  AOI210     u579(.A0(men_men_n601_), .A1(men_men_n234_), .B0(men_men_n158_), .Y(men_men_n602_));
  OR2        u580(.A(i_6_), .B(i_10_), .Y(men_men_n603_));
  NO2        u581(.A(men_men_n603_), .B(men_men_n23_), .Y(men_men_n604_));
  OR3        u582(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n605_));
  NO3        u583(.A(men_men_n605_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n606_));
  INV        u584(.A(men_men_n198_), .Y(men_men_n607_));
  NO2        u585(.A(men_men_n606_), .B(men_men_n604_), .Y(men_men_n608_));
  OA220      u586(.A0(men_men_n608_), .A1(i_2_), .B0(men_men_n602_), .B1(men_men_n267_), .Y(men_men_n609_));
  AOI210     u587(.A0(men_men_n609_), .A1(men_men_n600_), .B0(men_men_n60_), .Y(men_men_n610_));
  NOi21      u588(.An(i_11_), .B(i_7_), .Y(men_men_n611_));
  AO210      u589(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n612_));
  NO2        u590(.A(men_men_n612_), .B(men_men_n611_), .Y(men_men_n613_));
  NA2        u591(.A(men_men_n613_), .B(men_men_n205_), .Y(men_men_n614_));
  NO2        u592(.A(men_men_n614_), .B(men_men_n60_), .Y(men_men_n615_));
  NA2        u593(.A(men_men_n84_), .B(men_men_n60_), .Y(men_men_n616_));
  AO210      u594(.A0(men_men_n616_), .A1(men_men_n375_), .B0(men_men_n41_), .Y(men_men_n617_));
  NA2        u595(.A(men_men_n223_), .B(men_men_n60_), .Y(men_men_n618_));
  NA2        u596(.A(men_men_n408_), .B(men_men_n31_), .Y(men_men_n619_));
  OR2        u597(.A(men_men_n207_), .B(men_men_n106_), .Y(men_men_n620_));
  NA2        u598(.A(men_men_n620_), .B(men_men_n619_), .Y(men_men_n621_));
  NO2        u599(.A(men_men_n60_), .B(i_9_), .Y(men_men_n622_));
  NO2        u600(.A(men_men_n622_), .B(i_4_), .Y(men_men_n623_));
  NA2        u601(.A(men_men_n623_), .B(men_men_n621_), .Y(men_men_n624_));
  NO2        u602(.A(i_1_), .B(i_12_), .Y(men_men_n625_));
  NA3        u603(.A(men_men_n625_), .B(men_men_n107_), .C(men_men_n24_), .Y(men_men_n626_));
  NA4        u604(.A(men_men_n626_), .B(men_men_n624_), .C(men_men_n618_), .D(men_men_n617_), .Y(men_men_n627_));
  OAI210     u605(.A0(men_men_n627_), .A1(men_men_n615_), .B0(i_6_), .Y(men_men_n628_));
  NO2        u606(.A(men_men_n234_), .B(men_men_n82_), .Y(men_men_n629_));
  NO2        u607(.A(men_men_n629_), .B(i_11_), .Y(men_men_n630_));
  INV        u608(.A(men_men_n455_), .Y(men_men_n631_));
  NO4        u609(.A(i_12_), .B(men_men_n126_), .C(i_13_), .D(men_men_n82_), .Y(men_men_n632_));
  NA2        u610(.A(men_men_n632_), .B(men_men_n622_), .Y(men_men_n633_));
  NO3        u611(.A(men_men_n603_), .B(men_men_n230_), .C(men_men_n23_), .Y(men_men_n634_));
  AOI210     u612(.A0(i_1_), .A1(men_men_n257_), .B0(men_men_n634_), .Y(men_men_n635_));
  OAI210     u613(.A0(men_men_n635_), .A1(men_men_n44_), .B0(men_men_n633_), .Y(men_men_n636_));
  NA3        u614(.A(men_men_n535_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n637_));
  NA2        u615(.A(men_men_n135_), .B(i_9_), .Y(men_men_n638_));
  NA3        u616(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n639_));
  NO2        u617(.A(men_men_n46_), .B(i_1_), .Y(men_men_n640_));
  NA3        u618(.A(men_men_n640_), .B(men_men_n266_), .C(men_men_n44_), .Y(men_men_n641_));
  OAI220     u619(.A0(men_men_n641_), .A1(men_men_n639_), .B0(men_men_n638_), .B1(men_men_n1013_), .Y(men_men_n642_));
  NA3        u620(.A(men_men_n622_), .B(men_men_n314_), .C(i_6_), .Y(men_men_n643_));
  NO2        u621(.A(men_men_n643_), .B(men_men_n23_), .Y(men_men_n644_));
  AOI210     u622(.A0(men_men_n475_), .A1(men_men_n417_), .B0(men_men_n238_), .Y(men_men_n645_));
  NO2        u623(.A(men_men_n645_), .B(men_men_n594_), .Y(men_men_n646_));
  NAi21      u624(.An(men_men_n637_), .B(men_men_n90_), .Y(men_men_n647_));
  NA2        u625(.A(men_men_n640_), .B(men_men_n266_), .Y(men_men_n648_));
  NO2        u626(.A(i_11_), .B(men_men_n37_), .Y(men_men_n649_));
  NA2        u627(.A(men_men_n649_), .B(men_men_n24_), .Y(men_men_n650_));
  OAI210     u628(.A0(men_men_n650_), .A1(men_men_n648_), .B0(men_men_n647_), .Y(men_men_n651_));
  OR4        u629(.A(men_men_n651_), .B(men_men_n646_), .C(men_men_n644_), .D(men_men_n642_), .Y(men_men_n652_));
  NO3        u630(.A(men_men_n652_), .B(men_men_n636_), .C(men_men_n631_), .Y(men_men_n653_));
  NO2        u631(.A(men_men_n234_), .B(men_men_n99_), .Y(men_men_n654_));
  NO2        u632(.A(men_men_n654_), .B(men_men_n611_), .Y(men_men_n655_));
  NO2        u633(.A(men_men_n414_), .B(men_men_n82_), .Y(men_men_n656_));
  NO2        u634(.A(men_men_n115_), .B(men_men_n37_), .Y(men_men_n657_));
  NO2        u635(.A(men_men_n82_), .B(i_9_), .Y(men_men_n658_));
  NO2        u636(.A(men_men_n658_), .B(men_men_n60_), .Y(men_men_n659_));
  NA2        u637(.A(i_1_), .B(i_3_), .Y(men_men_n660_));
  NA2        u638(.A(men_men_n653_), .B(men_men_n628_), .Y(men_men_n661_));
  NA2        u639(.A(men_men_n367_), .B(men_men_n366_), .Y(men_men_n662_));
  NO3        u640(.A(men_men_n477_), .B(men_men_n597_), .C(men_men_n82_), .Y(men_men_n663_));
  NA2        u641(.A(men_men_n663_), .B(men_men_n25_), .Y(men_men_n664_));
  NA3        u642(.A(men_men_n158_), .B(men_men_n80_), .C(men_men_n82_), .Y(men_men_n665_));
  NA3        u643(.A(men_men_n665_), .B(men_men_n664_), .C(men_men_n662_), .Y(men_men_n666_));
  NA2        u644(.A(men_men_n666_), .B(i_1_), .Y(men_men_n667_));
  AOI210     u645(.A0(men_men_n266_), .A1(men_men_n95_), .B0(i_1_), .Y(men_men_n668_));
  NO2        u646(.A(men_men_n365_), .B(i_2_), .Y(men_men_n669_));
  NA2        u647(.A(men_men_n669_), .B(men_men_n668_), .Y(men_men_n670_));
  AOI210     u648(.A0(men_men_n670_), .A1(men_men_n667_), .B0(i_13_), .Y(men_men_n671_));
  OR2        u649(.A(i_11_), .B(i_7_), .Y(men_men_n672_));
  NA3        u650(.A(men_men_n672_), .B(men_men_n104_), .C(men_men_n135_), .Y(men_men_n673_));
  AOI220     u651(.A0(men_men_n470_), .A1(men_men_n158_), .B0(men_men_n449_), .B1(men_men_n135_), .Y(men_men_n674_));
  OAI210     u652(.A0(men_men_n674_), .A1(men_men_n44_), .B0(men_men_n673_), .Y(men_men_n675_));
  NO2        u653(.A(men_men_n52_), .B(i_12_), .Y(men_men_n676_));
  NO2        u654(.A(men_men_n477_), .B(men_men_n24_), .Y(men_men_n677_));
  AOI220     u655(.A0(men_men_n677_), .A1(men_men_n656_), .B0(men_men_n242_), .B1(men_men_n129_), .Y(men_men_n678_));
  OAI220     u656(.A0(men_men_n678_), .A1(men_men_n41_), .B0(men_men_n1012_), .B1(men_men_n91_), .Y(men_men_n679_));
  AOI210     u657(.A0(men_men_n675_), .A1(men_men_n330_), .B0(men_men_n679_), .Y(men_men_n680_));
  NA2        u658(.A(men_men_n383_), .B(men_men_n640_), .Y(men_men_n681_));
  NO2        u659(.A(men_men_n681_), .B(men_men_n239_), .Y(men_men_n682_));
  AOI210     u660(.A0(men_men_n447_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n683_));
  NOi31      u661(.An(men_men_n683_), .B(men_men_n586_), .C(men_men_n44_), .Y(men_men_n684_));
  NA2        u662(.A(men_men_n125_), .B(i_13_), .Y(men_men_n685_));
  NO2        u663(.A(men_men_n639_), .B(men_men_n112_), .Y(men_men_n686_));
  INV        u664(.A(men_men_n686_), .Y(men_men_n687_));
  OAI220     u665(.A0(men_men_n687_), .A1(men_men_n68_), .B0(men_men_n685_), .B1(men_men_n668_), .Y(men_men_n688_));
  NO3        u666(.A(men_men_n68_), .B(men_men_n32_), .C(men_men_n99_), .Y(men_men_n689_));
  NA2        u667(.A(men_men_n26_), .B(men_men_n192_), .Y(men_men_n690_));
  INV        u668(.A(i_7_), .Y(men_men_n691_));
  INV        u669(.A(men_men_n689_), .Y(men_men_n692_));
  AOI220     u670(.A0(men_men_n383_), .A1(men_men_n640_), .B0(men_men_n90_), .B1(men_men_n100_), .Y(men_men_n693_));
  OAI220     u671(.A0(men_men_n693_), .A1(men_men_n592_), .B0(men_men_n692_), .B1(men_men_n607_), .Y(men_men_n694_));
  NO4        u672(.A(men_men_n694_), .B(men_men_n688_), .C(men_men_n684_), .D(men_men_n682_), .Y(men_men_n695_));
  OR2        u673(.A(i_11_), .B(i_6_), .Y(men_men_n696_));
  NA3        u674(.A(men_men_n591_), .B(men_men_n690_), .C(i_7_), .Y(men_men_n697_));
  AOI210     u675(.A0(men_men_n697_), .A1(men_men_n687_), .B0(men_men_n696_), .Y(men_men_n698_));
  NA3        u676(.A(men_men_n408_), .B(men_men_n596_), .C(men_men_n95_), .Y(men_men_n699_));
  NA2        u677(.A(men_men_n630_), .B(i_13_), .Y(men_men_n700_));
  NA2        u678(.A(men_men_n100_), .B(men_men_n690_), .Y(men_men_n701_));
  NAi21      u679(.An(i_11_), .B(i_12_), .Y(men_men_n702_));
  NOi41      u680(.An(men_men_n108_), .B(men_men_n702_), .C(i_13_), .D(men_men_n82_), .Y(men_men_n703_));
  NA2        u681(.A(men_men_n703_), .B(men_men_n701_), .Y(men_men_n704_));
  NA3        u682(.A(men_men_n704_), .B(men_men_n700_), .C(men_men_n699_), .Y(men_men_n705_));
  OAI210     u683(.A0(men_men_n705_), .A1(men_men_n698_), .B0(men_men_n60_), .Y(men_men_n706_));
  NO2        u684(.A(i_2_), .B(i_12_), .Y(men_men_n707_));
  NA2        u685(.A(men_men_n364_), .B(men_men_n707_), .Y(men_men_n708_));
  NA2        u686(.A(i_8_), .B(men_men_n25_), .Y(men_men_n709_));
  NO3        u687(.A(men_men_n709_), .B(men_men_n381_), .C(men_men_n591_), .Y(men_men_n710_));
  OAI210     u688(.A0(men_men_n710_), .A1(men_men_n366_), .B0(men_men_n364_), .Y(men_men_n711_));
  NO2        u689(.A(men_men_n126_), .B(i_2_), .Y(men_men_n712_));
  NA2        u690(.A(men_men_n712_), .B(men_men_n625_), .Y(men_men_n713_));
  NA3        u691(.A(men_men_n713_), .B(men_men_n711_), .C(men_men_n708_), .Y(men_men_n714_));
  NA3        u692(.A(men_men_n714_), .B(men_men_n45_), .C(men_men_n222_), .Y(men_men_n715_));
  NA4        u693(.A(men_men_n715_), .B(men_men_n706_), .C(men_men_n695_), .D(men_men_n680_), .Y(men_men_n716_));
  OR4        u694(.A(men_men_n716_), .B(men_men_n671_), .C(men_men_n661_), .D(men_men_n610_), .Y(men5));
  NA2        u695(.A(men_men_n655_), .B(men_men_n268_), .Y(men_men_n718_));
  AN2        u696(.A(men_men_n24_), .B(i_10_), .Y(men_men_n719_));
  NA3        u697(.A(men_men_n719_), .B(men_men_n707_), .C(men_men_n106_), .Y(men_men_n720_));
  NO2        u698(.A(men_men_n592_), .B(i_11_), .Y(men_men_n721_));
  NA2        u699(.A(men_men_n85_), .B(men_men_n721_), .Y(men_men_n722_));
  NA3        u700(.A(men_men_n722_), .B(men_men_n720_), .C(men_men_n718_), .Y(men_men_n723_));
  NO3        u701(.A(i_11_), .B(men_men_n234_), .C(i_13_), .Y(men_men_n724_));
  NO2        u702(.A(men_men_n122_), .B(men_men_n23_), .Y(men_men_n725_));
  NA2        u703(.A(i_12_), .B(i_8_), .Y(men_men_n726_));
  OAI210     u704(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n726_), .Y(men_men_n727_));
  INV        u705(.A(men_men_n446_), .Y(men_men_n728_));
  AOI220     u706(.A0(men_men_n314_), .A1(men_men_n569_), .B0(men_men_n727_), .B1(men_men_n725_), .Y(men_men_n729_));
  INV        u707(.A(men_men_n729_), .Y(men_men_n730_));
  NO2        u708(.A(men_men_n730_), .B(men_men_n723_), .Y(men_men_n731_));
  INV        u709(.A(men_men_n169_), .Y(men_men_n732_));
  INV        u710(.A(men_men_n242_), .Y(men_men_n733_));
  OAI210     u711(.A0(men_men_n669_), .A1(men_men_n448_), .B0(men_men_n108_), .Y(men_men_n734_));
  AOI210     u712(.A0(men_men_n734_), .A1(men_men_n733_), .B0(men_men_n732_), .Y(men_men_n735_));
  NO2        u713(.A(men_men_n456_), .B(men_men_n26_), .Y(men_men_n736_));
  NO2        u714(.A(men_men_n736_), .B(men_men_n417_), .Y(men_men_n737_));
  NA2        u715(.A(men_men_n737_), .B(i_2_), .Y(men_men_n738_));
  INV        u716(.A(men_men_n738_), .Y(men_men_n739_));
  AOI210     u717(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n415_), .Y(men_men_n740_));
  AOI210     u718(.A0(men_men_n740_), .A1(men_men_n739_), .B0(men_men_n735_), .Y(men_men_n741_));
  NO2        u719(.A(men_men_n189_), .B(men_men_n123_), .Y(men_men_n742_));
  OAI210     u720(.A0(men_men_n742_), .A1(men_men_n725_), .B0(i_2_), .Y(men_men_n743_));
  INV        u721(.A(men_men_n170_), .Y(men_men_n744_));
  NO3        u722(.A(men_men_n612_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n745_));
  AOI210     u723(.A0(men_men_n744_), .A1(men_men_n85_), .B0(men_men_n745_), .Y(men_men_n746_));
  AOI210     u724(.A0(men_men_n746_), .A1(men_men_n743_), .B0(men_men_n192_), .Y(men_men_n747_));
  OA210      u725(.A0(men_men_n613_), .A1(men_men_n124_), .B0(i_13_), .Y(men_men_n748_));
  NA2        u726(.A(men_men_n148_), .B(men_men_n587_), .Y(men_men_n749_));
  NO2        u727(.A(men_men_n749_), .B(men_men_n369_), .Y(men_men_n750_));
  AOI210     u728(.A0(men_men_n207_), .A1(men_men_n145_), .B0(men_men_n520_), .Y(men_men_n751_));
  NA2        u729(.A(men_men_n751_), .B(men_men_n417_), .Y(men_men_n752_));
  NO2        u730(.A(men_men_n100_), .B(men_men_n44_), .Y(men_men_n753_));
  INV        u731(.A(men_men_n298_), .Y(men_men_n754_));
  NA4        u732(.A(men_men_n754_), .B(men_men_n302_), .C(men_men_n122_), .D(men_men_n42_), .Y(men_men_n755_));
  OAI210     u733(.A0(men_men_n755_), .A1(men_men_n753_), .B0(men_men_n752_), .Y(men_men_n756_));
  NO4        u734(.A(men_men_n756_), .B(men_men_n750_), .C(men_men_n748_), .D(men_men_n747_), .Y(men_men_n757_));
  NA2        u735(.A(men_men_n569_), .B(men_men_n28_), .Y(men_men_n758_));
  NA2        u736(.A(men_men_n724_), .B(men_men_n272_), .Y(men_men_n759_));
  NA2        u737(.A(men_men_n759_), .B(men_men_n758_), .Y(men_men_n760_));
  NO2        u738(.A(men_men_n59_), .B(i_12_), .Y(men_men_n761_));
  NO2        u739(.A(men_men_n761_), .B(men_men_n124_), .Y(men_men_n762_));
  NO2        u740(.A(men_men_n762_), .B(men_men_n587_), .Y(men_men_n763_));
  AOI220     u741(.A0(men_men_n763_), .A1(men_men_n36_), .B0(men_men_n760_), .B1(men_men_n46_), .Y(men_men_n764_));
  NA4        u742(.A(men_men_n764_), .B(men_men_n757_), .C(men_men_n741_), .D(men_men_n731_), .Y(men6));
  NO3        u743(.A(men_men_n253_), .B(men_men_n304_), .C(i_1_), .Y(men_men_n766_));
  NO2        u744(.A(men_men_n184_), .B(men_men_n136_), .Y(men_men_n767_));
  OAI210     u745(.A0(men_men_n767_), .A1(men_men_n766_), .B0(men_men_n712_), .Y(men_men_n768_));
  NA4        u746(.A(men_men_n387_), .B(men_men_n482_), .C(men_men_n68_), .D(men_men_n99_), .Y(men_men_n769_));
  INV        u747(.A(men_men_n769_), .Y(men_men_n770_));
  NO2        u748(.A(men_men_n217_), .B(men_men_n486_), .Y(men_men_n771_));
  NO2        u749(.A(i_11_), .B(i_9_), .Y(men_men_n772_));
  NO2        u750(.A(men_men_n770_), .B(men_men_n326_), .Y(men_men_n773_));
  AO210      u751(.A0(men_men_n773_), .A1(men_men_n768_), .B0(i_12_), .Y(men_men_n774_));
  NA2        u752(.A(men_men_n370_), .B(men_men_n333_), .Y(men_men_n775_));
  NA2        u753(.A(men_men_n574_), .B(men_men_n60_), .Y(men_men_n776_));
  BUFFER     u754(.A(men_men_n616_), .Y(men_men_n777_));
  NA3        u755(.A(men_men_n777_), .B(men_men_n776_), .C(men_men_n775_), .Y(men_men_n778_));
  INV        u756(.A(men_men_n195_), .Y(men_men_n779_));
  AOI220     u757(.A0(men_men_n779_), .A1(men_men_n772_), .B0(men_men_n778_), .B1(men_men_n70_), .Y(men_men_n780_));
  INV        u758(.A(men_men_n325_), .Y(men_men_n781_));
  NA2        u759(.A(men_men_n72_), .B(men_men_n129_), .Y(men_men_n782_));
  INV        u760(.A(men_men_n122_), .Y(men_men_n783_));
  NA2        u761(.A(men_men_n783_), .B(men_men_n46_), .Y(men_men_n784_));
  AOI210     u762(.A0(men_men_n784_), .A1(men_men_n782_), .B0(men_men_n781_), .Y(men_men_n785_));
  NO2        u763(.A(men_men_n249_), .B(i_9_), .Y(men_men_n786_));
  NA2        u764(.A(men_men_n786_), .B(men_men_n761_), .Y(men_men_n787_));
  AOI210     u765(.A0(men_men_n787_), .A1(men_men_n518_), .B0(men_men_n184_), .Y(men_men_n788_));
  NAi32      u766(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n789_));
  NO2        u767(.A(men_men_n696_), .B(men_men_n789_), .Y(men_men_n790_));
  OR3        u768(.A(men_men_n790_), .B(men_men_n788_), .C(men_men_n785_), .Y(men_men_n791_));
  NO2        u769(.A(men_men_n672_), .B(i_2_), .Y(men_men_n792_));
  NA2        u770(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n793_));
  NO2        u771(.A(men_men_n793_), .B(men_men_n407_), .Y(men_men_n794_));
  NA2        u772(.A(men_men_n794_), .B(men_men_n792_), .Y(men_men_n795_));
  OR2        u773(.A(men_men_n613_), .B(men_men_n448_), .Y(men_men_n796_));
  NA3        u774(.A(men_men_n796_), .B(men_men_n144_), .C(men_men_n66_), .Y(men_men_n797_));
  AO210      u775(.A0(men_men_n492_), .A1(men_men_n728_), .B0(men_men_n36_), .Y(men_men_n798_));
  NA3        u776(.A(men_men_n798_), .B(men_men_n797_), .C(men_men_n795_), .Y(men_men_n799_));
  OAI210     u777(.A0(men_men_n629_), .A1(i_11_), .B0(men_men_n83_), .Y(men_men_n800_));
  AOI220     u778(.A0(men_men_n800_), .A1(men_men_n559_), .B0(men_men_n771_), .B1(men_men_n691_), .Y(men_men_n801_));
  NA2        u779(.A(men_men_n393_), .B(men_men_n67_), .Y(men_men_n802_));
  NA3        u780(.A(men_men_n802_), .B(men_men_n801_), .C(men_men_n595_), .Y(men_men_n803_));
  AO210      u781(.A0(men_men_n520_), .A1(men_men_n46_), .B0(men_men_n84_), .Y(men_men_n804_));
  NA3        u782(.A(men_men_n804_), .B(men_men_n483_), .C(men_men_n216_), .Y(men_men_n805_));
  AOI210     u783(.A0(men_men_n448_), .A1(men_men_n446_), .B0(men_men_n558_), .Y(men_men_n806_));
  NA2        u784(.A(men_men_n109_), .B(men_men_n406_), .Y(men_men_n807_));
  INV        u785(.A(men_men_n241_), .Y(men_men_n808_));
  NA3        u786(.A(men_men_n807_), .B(men_men_n806_), .C(men_men_n805_), .Y(men_men_n809_));
  NO4        u787(.A(men_men_n809_), .B(men_men_n803_), .C(men_men_n799_), .D(men_men_n791_), .Y(men_men_n810_));
  NA4        u788(.A(men_men_n810_), .B(men_men_n780_), .C(men_men_n774_), .D(men_men_n377_), .Y(men3));
  NA2        u789(.A(i_6_), .B(i_7_), .Y(men_men_n812_));
  NO2        u790(.A(men_men_n812_), .B(i_0_), .Y(men_men_n813_));
  NO2        u791(.A(i_11_), .B(men_men_n234_), .Y(men_men_n814_));
  OAI210     u792(.A0(men_men_n813_), .A1(men_men_n286_), .B0(men_men_n814_), .Y(men_men_n815_));
  NO2        u793(.A(men_men_n815_), .B(men_men_n192_), .Y(men_men_n816_));
  NO3        u794(.A(men_men_n452_), .B(men_men_n88_), .C(men_men_n44_), .Y(men_men_n817_));
  OA210      u795(.A0(men_men_n817_), .A1(men_men_n816_), .B0(men_men_n172_), .Y(men_men_n818_));
  NA2        u796(.A(men_men_n595_), .B(men_men_n368_), .Y(men_men_n819_));
  NA2        u797(.A(men_men_n819_), .B(men_men_n40_), .Y(men_men_n820_));
  NO3        u798(.A(men_men_n620_), .B(men_men_n456_), .C(men_men_n129_), .Y(men_men_n821_));
  AN2        u799(.A(men_men_n454_), .B(men_men_n53_), .Y(men_men_n822_));
  NO2        u800(.A(men_men_n822_), .B(men_men_n821_), .Y(men_men_n823_));
  AOI210     u801(.A0(men_men_n823_), .A1(men_men_n820_), .B0(men_men_n48_), .Y(men_men_n824_));
  NO4        u802(.A(men_men_n373_), .B(men_men_n380_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n825_));
  NA2        u803(.A(men_men_n184_), .B(men_men_n567_), .Y(men_men_n826_));
  NOi21      u804(.An(men_men_n826_), .B(men_men_n825_), .Y(men_men_n827_));
  NO2        u805(.A(men_men_n827_), .B(men_men_n60_), .Y(men_men_n828_));
  NOi21      u806(.An(i_5_), .B(i_9_), .Y(men_men_n829_));
  NA2        u807(.A(men_men_n829_), .B(men_men_n445_), .Y(men_men_n830_));
  BUFFER     u808(.A(men_men_n266_), .Y(men_men_n831_));
  AOI210     u809(.A0(men_men_n831_), .A1(men_men_n475_), .B0(men_men_n663_), .Y(men_men_n832_));
  NO2        u810(.A(men_men_n173_), .B(men_men_n145_), .Y(men_men_n833_));
  NO2        u811(.A(men_men_n832_), .B(men_men_n830_), .Y(men_men_n834_));
  NO4        u812(.A(men_men_n834_), .B(men_men_n828_), .C(men_men_n824_), .D(men_men_n818_), .Y(men_men_n835_));
  NA2        u813(.A(men_men_n184_), .B(men_men_n24_), .Y(men_men_n836_));
  NO2        u814(.A(men_men_n657_), .B(men_men_n584_), .Y(men_men_n837_));
  NO2        u815(.A(men_men_n837_), .B(men_men_n836_), .Y(men_men_n838_));
  NA2        u816(.A(men_men_n309_), .B(men_men_n127_), .Y(men_men_n839_));
  NAi21      u817(.An(men_men_n159_), .B(men_men_n437_), .Y(men_men_n840_));
  OAI220     u818(.A0(men_men_n840_), .A1(men_men_n808_), .B0(men_men_n839_), .B1(men_men_n398_), .Y(men_men_n841_));
  NO2        u819(.A(men_men_n841_), .B(men_men_n838_), .Y(men_men_n842_));
  NO2        u820(.A(men_men_n387_), .B(men_men_n290_), .Y(men_men_n843_));
  NA2        u821(.A(men_men_n843_), .B(men_men_n686_), .Y(men_men_n844_));
  NA2        u822(.A(men_men_n568_), .B(i_0_), .Y(men_men_n845_));
  NO3        u823(.A(men_men_n845_), .B(men_men_n382_), .C(men_men_n85_), .Y(men_men_n846_));
  INV        u824(.A(men_men_n846_), .Y(men_men_n847_));
  AN2        u825(.A(men_men_n94_), .B(men_men_n240_), .Y(men_men_n848_));
  NA2        u826(.A(men_men_n724_), .B(men_men_n326_), .Y(men_men_n849_));
  INV        u827(.A(men_men_n55_), .Y(men_men_n850_));
  OAI220     u828(.A0(men_men_n850_), .A1(men_men_n849_), .B0(men_men_n650_), .B1(men_men_n537_), .Y(men_men_n851_));
  NO2        u829(.A(men_men_n251_), .B(men_men_n150_), .Y(men_men_n852_));
  NA2        u830(.A(i_0_), .B(i_10_), .Y(men_men_n853_));
  AN2        u831(.A(men_men_n852_), .B(i_6_), .Y(men_men_n854_));
  AOI220     u832(.A0(men_men_n331_), .A1(men_men_n96_), .B0(men_men_n184_), .B1(men_men_n80_), .Y(men_men_n855_));
  NA2        u833(.A(men_men_n563_), .B(i_4_), .Y(men_men_n856_));
  NA2        u834(.A(men_men_n187_), .B(men_men_n201_), .Y(men_men_n857_));
  OAI220     u835(.A0(men_men_n857_), .A1(men_men_n849_), .B0(men_men_n856_), .B1(men_men_n855_), .Y(men_men_n858_));
  NO4        u836(.A(men_men_n858_), .B(men_men_n854_), .C(men_men_n851_), .D(men_men_n848_), .Y(men_men_n859_));
  NA4        u837(.A(men_men_n859_), .B(men_men_n847_), .C(men_men_n844_), .D(men_men_n842_), .Y(men_men_n860_));
  NO2        u838(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n861_));
  NA2        u839(.A(i_11_), .B(i_9_), .Y(men_men_n862_));
  NO3        u840(.A(i_12_), .B(men_men_n862_), .C(men_men_n594_), .Y(men_men_n863_));
  AN2        u841(.A(men_men_n863_), .B(men_men_n861_), .Y(men_men_n864_));
  NO2        u842(.A(men_men_n48_), .B(i_7_), .Y(men_men_n865_));
  NA2        u843(.A(men_men_n391_), .B(men_men_n177_), .Y(men_men_n866_));
  NA2        u844(.A(men_men_n866_), .B(men_men_n157_), .Y(men_men_n867_));
  NO2        u845(.A(men_men_n173_), .B(i_0_), .Y(men_men_n868_));
  INV        u846(.A(men_men_n868_), .Y(men_men_n869_));
  NA2        u847(.A(men_men_n473_), .B(men_men_n228_), .Y(men_men_n870_));
  INV        u848(.A(men_men_n405_), .Y(men_men_n871_));
  OAI220     u849(.A0(men_men_n871_), .A1(men_men_n830_), .B0(men_men_n870_), .B1(men_men_n869_), .Y(men_men_n872_));
  NO3        u850(.A(men_men_n872_), .B(men_men_n867_), .C(men_men_n864_), .Y(men_men_n873_));
  NA2        u851(.A(men_men_n649_), .B(men_men_n119_), .Y(men_men_n874_));
  NO2        u852(.A(i_6_), .B(men_men_n874_), .Y(men_men_n875_));
  AOI210     u853(.A0(men_men_n447_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n876_));
  NA2        u854(.A(men_men_n169_), .B(men_men_n101_), .Y(men_men_n877_));
  NOi32      u855(.An(men_men_n876_), .Bn(men_men_n187_), .C(men_men_n877_), .Y(men_men_n878_));
  NO2        u856(.A(men_men_n878_), .B(men_men_n875_), .Y(men_men_n879_));
  NOi21      u857(.An(i_7_), .B(i_5_), .Y(men_men_n880_));
  NOi31      u858(.An(men_men_n880_), .B(i_0_), .C(men_men_n702_), .Y(men_men_n881_));
  NA3        u859(.A(men_men_n881_), .B(men_men_n381_), .C(i_6_), .Y(men_men_n882_));
  OA210      u860(.A0(men_men_n877_), .A1(men_men_n518_), .B0(men_men_n882_), .Y(men_men_n883_));
  NO3        u861(.A(men_men_n401_), .B(men_men_n359_), .C(men_men_n357_), .Y(men_men_n884_));
  NO2        u862(.A(men_men_n260_), .B(men_men_n315_), .Y(men_men_n885_));
  NO2        u863(.A(men_men_n702_), .B(men_men_n255_), .Y(men_men_n886_));
  AOI210     u864(.A0(men_men_n886_), .A1(men_men_n885_), .B0(men_men_n884_), .Y(men_men_n887_));
  NA4        u865(.A(men_men_n887_), .B(men_men_n883_), .C(men_men_n879_), .D(men_men_n873_), .Y(men_men_n888_));
  NO2        u866(.A(men_men_n836_), .B(men_men_n236_), .Y(men_men_n889_));
  AN2        u867(.A(men_men_n330_), .B(men_men_n326_), .Y(men_men_n890_));
  AN2        u868(.A(men_men_n890_), .B(men_men_n833_), .Y(men_men_n891_));
  OAI210     u869(.A0(men_men_n891_), .A1(men_men_n889_), .B0(i_10_), .Y(men_men_n892_));
  OA210      u870(.A0(men_men_n473_), .A1(men_men_n220_), .B0(men_men_n472_), .Y(men_men_n893_));
  NA3        u871(.A(men_men_n472_), .B(men_men_n408_), .C(men_men_n45_), .Y(men_men_n894_));
  INV        u872(.A(men_men_n894_), .Y(men_men_n895_));
  NO2        u873(.A(i_3_), .B(men_men_n186_), .Y(men_men_n896_));
  AOI220     u874(.A0(men_men_n896_), .A1(men_men_n473_), .B0(men_men_n895_), .B1(men_men_n70_), .Y(men_men_n897_));
  NA3        u875(.A(men_men_n793_), .B(men_men_n379_), .C(men_men_n629_), .Y(men_men_n898_));
  NA2        u876(.A(men_men_n91_), .B(men_men_n44_), .Y(men_men_n899_));
  NO2        u877(.A(men_men_n72_), .B(men_men_n726_), .Y(men_men_n900_));
  AOI220     u878(.A0(men_men_n900_), .A1(men_men_n899_), .B0(men_men_n172_), .B1(men_men_n584_), .Y(men_men_n901_));
  AOI210     u879(.A0(men_men_n901_), .A1(men_men_n898_), .B0(men_men_n47_), .Y(men_men_n902_));
  NAi21      u880(.An(i_9_), .B(i_5_), .Y(men_men_n903_));
  NO2        u881(.A(men_men_n903_), .B(men_men_n401_), .Y(men_men_n904_));
  NO2        u882(.A(men_men_n590_), .B(men_men_n103_), .Y(men_men_n905_));
  AOI220     u883(.A0(men_men_n905_), .A1(i_0_), .B0(men_men_n904_), .B1(men_men_n613_), .Y(men_men_n906_));
  NO2        u884(.A(men_men_n906_), .B(men_men_n82_), .Y(men_men_n907_));
  NO3        u885(.A(men_men_n907_), .B(men_men_n902_), .C(men_men_n523_), .Y(men_men_n908_));
  NA3        u886(.A(men_men_n908_), .B(men_men_n897_), .C(men_men_n892_), .Y(men_men_n909_));
  NO3        u887(.A(men_men_n909_), .B(men_men_n888_), .C(men_men_n860_), .Y(men_men_n910_));
  NA2        u888(.A(men_men_n70_), .B(men_men_n44_), .Y(men_men_n911_));
  NA2        u889(.A(men_men_n853_), .B(men_men_n911_), .Y(men_men_n912_));
  NO3        u890(.A(men_men_n103_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n913_));
  AN2        u891(.A(men_men_n913_), .B(men_men_n912_), .Y(men_men_n914_));
  AOI210     u892(.A0(men_men_n776_), .A1(men_men_n662_), .B0(men_men_n877_), .Y(men_men_n915_));
  AOI210     u893(.A0(men_men_n914_), .A1(men_men_n348_), .B0(men_men_n915_), .Y(men_men_n916_));
  NA2        u894(.A(men_men_n712_), .B(men_men_n143_), .Y(men_men_n917_));
  INV        u895(.A(men_men_n917_), .Y(men_men_n918_));
  NA3        u896(.A(men_men_n918_), .B(men_men_n658_), .C(men_men_n70_), .Y(men_men_n919_));
  NA3        u897(.A(men_men_n813_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n920_));
  NA2        u898(.A(men_men_n814_), .B(i_9_), .Y(men_men_n921_));
  AOI210     u899(.A0(men_men_n920_), .A1(men_men_n497_), .B0(men_men_n921_), .Y(men_men_n922_));
  NA2        u900(.A(men_men_n241_), .B(men_men_n227_), .Y(men_men_n923_));
  AOI210     u901(.A0(men_men_n923_), .A1(men_men_n845_), .B0(men_men_n150_), .Y(men_men_n924_));
  NO2        u902(.A(men_men_n924_), .B(men_men_n922_), .Y(men_men_n925_));
  NA3        u903(.A(men_men_n925_), .B(men_men_n919_), .C(men_men_n916_), .Y(men_men_n926_));
  NA2        u904(.A(men_men_n890_), .B(men_men_n369_), .Y(men_men_n927_));
  AOI210     u905(.A0(men_men_n297_), .A1(men_men_n159_), .B0(men_men_n927_), .Y(men_men_n928_));
  NA2        u906(.A(men_men_n40_), .B(men_men_n44_), .Y(men_men_n929_));
  NA2        u907(.A(men_men_n865_), .B(men_men_n487_), .Y(men_men_n930_));
  AOI210     u908(.A0(men_men_n929_), .A1(men_men_n159_), .B0(men_men_n930_), .Y(men_men_n931_));
  NO2        u909(.A(men_men_n931_), .B(men_men_n928_), .Y(men_men_n932_));
  NO3        u910(.A(men_men_n853_), .B(men_men_n829_), .C(men_men_n189_), .Y(men_men_n933_));
  AOI220     u911(.A0(men_men_n933_), .A1(i_11_), .B0(men_men_n564_), .B1(men_men_n72_), .Y(men_men_n934_));
  NO3        u912(.A(men_men_n209_), .B(men_men_n380_), .C(i_0_), .Y(men_men_n935_));
  OAI210     u913(.A0(men_men_n935_), .A1(men_men_n73_), .B0(i_13_), .Y(men_men_n936_));
  INV        u914(.A(men_men_n216_), .Y(men_men_n937_));
  NO2        u915(.A(men_men_n531_), .B(men_men_n136_), .Y(men_men_n938_));
  NA3        u916(.A(men_men_n938_), .B(men_men_n1017_), .C(men_men_n937_), .Y(men_men_n939_));
  NA4        u917(.A(men_men_n939_), .B(men_men_n936_), .C(men_men_n934_), .D(men_men_n932_), .Y(men_men_n940_));
  AOI220     u918(.A0(men_men_n880_), .A1(men_men_n487_), .B0(men_men_n813_), .B1(men_men_n160_), .Y(men_men_n941_));
  NA2        u919(.A(men_men_n351_), .B(men_men_n174_), .Y(men_men_n942_));
  OR2        u920(.A(men_men_n942_), .B(men_men_n941_), .Y(men_men_n943_));
  AOI210     u921(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n173_), .Y(men_men_n944_));
  NA2        u922(.A(men_men_n944_), .B(men_men_n893_), .Y(men_men_n945_));
  NA3        u923(.A(men_men_n387_), .B(men_men_n169_), .C(men_men_n168_), .Y(men_men_n946_));
  NA3        u924(.A(men_men_n865_), .B(men_men_n286_), .C(men_men_n227_), .Y(men_men_n947_));
  NA2        u925(.A(men_men_n947_), .B(men_men_n946_), .Y(men_men_n948_));
  NA3        u926(.A(men_men_n387_), .B(men_men_n332_), .C(men_men_n218_), .Y(men_men_n949_));
  INV        u927(.A(men_men_n949_), .Y(men_men_n950_));
  NOi31      u928(.An(men_men_n386_), .B(men_men_n911_), .C(men_men_n236_), .Y(men_men_n951_));
  NO3        u929(.A(men_men_n951_), .B(men_men_n950_), .C(men_men_n948_), .Y(men_men_n952_));
  NA3        u930(.A(men_men_n952_), .B(men_men_n945_), .C(men_men_n943_), .Y(men_men_n953_));
  NO2        u931(.A(men_men_n82_), .B(i_5_), .Y(men_men_n954_));
  NA3        u932(.A(men_men_n814_), .B(men_men_n107_), .C(men_men_n122_), .Y(men_men_n955_));
  INV        u933(.A(men_men_n955_), .Y(men_men_n956_));
  NA2        u934(.A(men_men_n956_), .B(men_men_n954_), .Y(men_men_n957_));
  NA2        u935(.A(men_men_n770_), .B(men_men_n174_), .Y(men_men_n958_));
  AN2        u936(.A(men_men_n853_), .B(men_men_n150_), .Y(men_men_n959_));
  NO4        u937(.A(men_men_n959_), .B(i_12_), .C(men_men_n637_), .D(men_men_n129_), .Y(men_men_n960_));
  NA2        u938(.A(men_men_n960_), .B(men_men_n216_), .Y(men_men_n961_));
  NA3        u939(.A(men_men_n96_), .B(men_men_n567_), .C(i_11_), .Y(men_men_n962_));
  NO2        u940(.A(men_men_n962_), .B(men_men_n152_), .Y(men_men_n963_));
  NA2        u941(.A(men_men_n880_), .B(men_men_n470_), .Y(men_men_n964_));
  NO2        u942(.A(men_men_n964_), .B(men_men_n659_), .Y(men_men_n965_));
  AOI210     u943(.A0(men_men_n965_), .A1(men_men_n868_), .B0(men_men_n963_), .Y(men_men_n966_));
  NA4        u944(.A(men_men_n966_), .B(men_men_n961_), .C(men_men_n958_), .D(men_men_n957_), .Y(men_men_n967_));
  NO4        u945(.A(men_men_n967_), .B(men_men_n953_), .C(men_men_n940_), .D(men_men_n926_), .Y(men_men_n968_));
  NA2        u946(.A(men_men_n792_), .B(men_men_n37_), .Y(men_men_n969_));
  NA3        u947(.A(men_men_n876_), .B(men_men_n364_), .C(i_5_), .Y(men_men_n970_));
  NA3        u948(.A(men_men_n970_), .B(men_men_n969_), .C(men_men_n602_), .Y(men_men_n971_));
  NA2        u949(.A(men_men_n971_), .B(men_men_n205_), .Y(men_men_n972_));
  NA2        u950(.A(men_men_n185_), .B(men_men_n187_), .Y(men_men_n973_));
  AO210      u951(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n973_), .Y(men_men_n974_));
  OAI210     u952(.A0(men_men_n606_), .A1(men_men_n604_), .B0(men_men_n314_), .Y(men_men_n975_));
  NAi31      u953(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n976_));
  AOI210     u954(.A0(men_men_n115_), .A1(men_men_n67_), .B0(men_men_n976_), .Y(men_men_n977_));
  NO2        u955(.A(men_men_n977_), .B(men_men_n634_), .Y(men_men_n978_));
  NA3        u956(.A(men_men_n978_), .B(men_men_n975_), .C(men_men_n974_), .Y(men_men_n979_));
  NO2        u957(.A(men_men_n460_), .B(men_men_n266_), .Y(men_men_n980_));
  NO4        u958(.A(men_men_n230_), .B(men_men_n142_), .C(men_men_n660_), .D(men_men_n37_), .Y(men_men_n981_));
  NO2        u959(.A(men_men_n981_), .B(men_men_n980_), .Y(men_men_n982_));
  OAI210     u960(.A0(men_men_n962_), .A1(men_men_n145_), .B0(men_men_n982_), .Y(men_men_n983_));
  AOI210     u961(.A0(men_men_n979_), .A1(men_men_n48_), .B0(men_men_n983_), .Y(men_men_n984_));
  AOI210     u962(.A0(men_men_n984_), .A1(men_men_n972_), .B0(men_men_n70_), .Y(men_men_n985_));
  NO2        u963(.A(men_men_n561_), .B(men_men_n376_), .Y(men_men_n986_));
  NO2        u964(.A(men_men_n986_), .B(men_men_n732_), .Y(men_men_n987_));
  OAI210     u965(.A0(men_men_n77_), .A1(men_men_n52_), .B0(men_men_n106_), .Y(men_men_n988_));
  NA2        u966(.A(men_men_n988_), .B(men_men_n73_), .Y(men_men_n989_));
  AOI210     u967(.A0(men_men_n944_), .A1(men_men_n865_), .B0(men_men_n881_), .Y(men_men_n990_));
  AOI210     u968(.A0(men_men_n990_), .A1(men_men_n989_), .B0(men_men_n660_), .Y(men_men_n991_));
  NA2        u969(.A(men_men_n260_), .B(men_men_n54_), .Y(men_men_n992_));
  AOI220     u970(.A0(men_men_n992_), .A1(men_men_n73_), .B0(men_men_n346_), .B1(men_men_n253_), .Y(men_men_n993_));
  NO2        u971(.A(men_men_n993_), .B(men_men_n234_), .Y(men_men_n994_));
  NA3        u972(.A(men_men_n94_), .B(men_men_n304_), .C(men_men_n31_), .Y(men_men_n995_));
  INV        u973(.A(men_men_n995_), .Y(men_men_n996_));
  NO3        u974(.A(men_men_n996_), .B(men_men_n994_), .C(men_men_n991_), .Y(men_men_n997_));
  OAI210     u975(.A0(men_men_n1015_), .A1(men_men_n876_), .B0(men_men_n205_), .Y(men_men_n998_));
  NA2        u976(.A(men_men_n161_), .B(i_5_), .Y(men_men_n999_));
  NO2        u977(.A(men_men_n998_), .B(men_men_n999_), .Y(men_men_n1000_));
  NO3        u978(.A(men_men_n56_), .B(men_men_n55_), .C(i_4_), .Y(men_men_n1001_));
  OAI210     u979(.A0(men_men_n885_), .A1(men_men_n304_), .B0(men_men_n1001_), .Y(men_men_n1002_));
  NO2        u980(.A(men_men_n1002_), .B(men_men_n702_), .Y(men_men_n1003_));
  INV        u981(.A(men_men_n360_), .Y(men_men_n1004_));
  NO2        u982(.A(men_men_n1004_), .B(men_men_n41_), .Y(men_men_n1005_));
  NO3        u983(.A(men_men_n1005_), .B(men_men_n1003_), .C(men_men_n1000_), .Y(men_men_n1006_));
  OAI210     u984(.A0(men_men_n997_), .A1(i_4_), .B0(men_men_n1006_), .Y(men_men_n1007_));
  NO3        u985(.A(men_men_n1007_), .B(men_men_n987_), .C(men_men_n985_), .Y(men_men_n1008_));
  NA4        u986(.A(men_men_n1008_), .B(men_men_n968_), .C(men_men_n910_), .D(men_men_n835_), .Y(men4));
  INV        u987(.A(men_men_n676_), .Y(men_men_n1012_));
  INV        u988(.A(i_2_), .Y(men_men_n1013_));
  INV        u989(.A(men_men_n483_), .Y(men_men_n1014_));
  INV        u990(.A(i_12_), .Y(men_men_n1015_));
  INV        u991(.A(i_12_), .Y(men_men_n1016_));
  INV        u992(.A(i_3_), .Y(men_men_n1017_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule