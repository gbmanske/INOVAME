// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n128_, new_new_n129_, new_new_n130_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n665_, new_new_n666_,
    new_new_n667_, new_new_n668_, new_new_n669_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n674_,
    new_new_n675_, new_new_n676_, new_new_n677_, new_new_n678_,
    new_new_n679_, new_new_n680_, new_new_n681_, new_new_n682_,
    new_new_n683_, new_new_n684_, new_new_n685_, new_new_n686_,
    new_new_n687_, new_new_n688_, new_new_n689_, new_new_n690_,
    new_new_n691_, new_new_n692_, new_new_n693_, new_new_n694_,
    new_new_n695_, new_new_n696_, new_new_n697_, new_new_n698_,
    new_new_n699_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n712_, new_new_n713_, new_new_n714_, new_new_n715_,
    new_new_n716_, new_new_n717_, new_new_n718_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n722_, new_new_n723_,
    new_new_n724_, new_new_n725_, new_new_n726_, new_new_n727_,
    new_new_n728_, new_new_n729_, new_new_n730_, new_new_n731_,
    new_new_n732_, new_new_n733_, new_new_n734_, new_new_n735_,
    new_new_n736_, new_new_n737_, new_new_n738_, new_new_n739_,
    new_new_n740_, new_new_n741_, new_new_n742_, new_new_n743_,
    new_new_n744_, new_new_n745_, new_new_n746_, new_new_n747_,
    new_new_n748_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n944_, new_new_n945_, new_new_n946_, new_new_n947_,
    new_new_n948_, new_new_n949_, new_new_n950_, new_new_n951_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(mai1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  NAi21      g035(.An(i_2_), .B(i_7_), .Y(new_new_n58_));
  INV        g036(.A(i_1_), .Y(new_new_n59_));
  NA2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NA2        g038(.A(i_1_), .B(i_10_), .Y(new_new_n61_));
  NO2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n50_), .B(i_2_), .Y(new_new_n63_));
  AOI210     g041(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_6_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(new_new_n25_), .Y(new_new_n66_));
  INV        g044(.A(i_0_), .Y(new_new_n67_));
  NAi21      g045(.An(i_5_), .B(i_10_), .Y(new_new_n68_));
  NA2        g046(.A(i_5_), .B(i_9_), .Y(new_new_n69_));
  AOI210     g047(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n67_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n66_), .Y(new_new_n71_));
  OAI210     g049(.A0(new_new_n64_), .A1(new_new_n63_), .B0(new_new_n71_), .Y(new_new_n72_));
  OAI210     g050(.A0(new_new_n72_), .A1(new_new_n62_), .B0(i_0_), .Y(new_new_n73_));
  NA2        g051(.A(i_12_), .B(i_5_), .Y(new_new_n74_));
  NA2        g052(.A(i_2_), .B(i_8_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_9_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_7_), .Y(new_new_n77_));
  NO3        g055(.A(new_new_n77_), .B(new_new_n76_), .C(new_new_n59_), .Y(new_new_n78_));
  INV        g056(.A(i_6_), .Y(new_new_n79_));
  OR4        g057(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n80_), .Y(new_new_n81_));
  NO2        g059(.A(i_2_), .B(i_7_), .Y(new_new_n82_));
  NA2        g060(.A(new_new_n78_), .B(new_new_n80_), .Y(new_new_n83_));
  NAi21      g061(.An(i_6_), .B(i_10_), .Y(new_new_n84_));
  NA2        g062(.A(i_6_), .B(i_9_), .Y(new_new_n85_));
  AOI210     g063(.A0(new_new_n85_), .A1(new_new_n84_), .B0(new_new_n59_), .Y(new_new_n86_));
  NA2        g064(.A(i_2_), .B(i_6_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n83_), .B(new_new_n74_), .Y(new_new_n88_));
  AN3        g066(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n89_));
  NAi21      g067(.An(i_6_), .B(i_11_), .Y(new_new_n90_));
  NO2        g068(.A(i_5_), .B(i_8_), .Y(new_new_n91_));
  NOi21      g069(.An(new_new_n91_), .B(new_new_n90_), .Y(new_new_n92_));
  AOI220     g070(.A0(new_new_n92_), .A1(new_new_n58_), .B0(new_new_n89_), .B1(new_new_n32_), .Y(new_new_n93_));
  INV        g071(.A(i_7_), .Y(new_new_n94_));
  NA2        g072(.A(new_new_n46_), .B(new_new_n94_), .Y(new_new_n95_));
  NO2        g073(.A(i_0_), .B(i_5_), .Y(new_new_n96_));
  NO2        g074(.A(new_new_n96_), .B(new_new_n79_), .Y(new_new_n97_));
  NA2        g075(.A(i_12_), .B(i_3_), .Y(new_new_n98_));
  INV        g076(.A(new_new_n98_), .Y(new_new_n99_));
  NA2        g077(.A(new_new_n99_), .B(new_new_n97_), .Y(new_new_n100_));
  NAi21      g078(.An(i_7_), .B(i_11_), .Y(new_new_n101_));
  AN2        g079(.A(i_2_), .B(i_10_), .Y(new_new_n102_));
  NO2        g080(.A(new_new_n102_), .B(i_7_), .Y(new_new_n103_));
  OR2        g081(.A(new_new_n74_), .B(new_new_n56_), .Y(new_new_n104_));
  NO2        g082(.A(i_8_), .B(new_new_n94_), .Y(new_new_n105_));
  NO3        g083(.A(new_new_n105_), .B(new_new_n104_), .C(new_new_n103_), .Y(new_new_n106_));
  NA2        g084(.A(i_12_), .B(i_7_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n59_), .B(new_new_n26_), .Y(new_new_n108_));
  NA2        g086(.A(new_new_n108_), .B(i_0_), .Y(new_new_n109_));
  NA2        g087(.A(i_11_), .B(i_12_), .Y(new_new_n110_));
  OAI210     g088(.A0(new_new_n109_), .A1(new_new_n107_), .B0(new_new_n110_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(new_new_n106_), .Y(new_new_n112_));
  NA3        g090(.A(new_new_n112_), .B(new_new_n100_), .C(new_new_n93_), .Y(new_new_n113_));
  NOi21      g091(.An(i_1_), .B(i_5_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(i_11_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n94_), .B(new_new_n37_), .Y(new_new_n116_));
  NA2        g094(.A(i_7_), .B(new_new_n25_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(new_new_n116_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n118_), .B(new_new_n46_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n85_), .B(new_new_n84_), .Y(new_new_n120_));
  NAi21      g098(.An(i_3_), .B(i_8_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(new_new_n58_), .Y(new_new_n122_));
  NO2        g100(.A(i_6_), .B(i_5_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(i_3_), .Y(new_new_n124_));
  NO2        g102(.A(new_new_n122_), .B(new_new_n115_), .Y(new_new_n125_));
  NO3        g103(.A(new_new_n125_), .B(new_new_n113_), .C(new_new_n88_), .Y(new_new_n126_));
  NA3        g104(.A(new_new_n126_), .B(new_new_n73_), .C(new_new_n55_), .Y(mai2));
  NO2        g105(.A(new_new_n59_), .B(new_new_n37_), .Y(new_new_n128_));
  NA2        g106(.A(i_6_), .B(new_new_n25_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n129_), .B(new_new_n128_), .Y(new_new_n130_));
  NA4        g108(.A(new_new_n130_), .B(new_new_n71_), .C(new_new_n63_), .D(new_new_n30_), .Y(mai0));
  AN2        g109(.A(i_8_), .B(i_7_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n132_), .B(i_6_), .Y(new_new_n133_));
  NO2        g111(.A(i_12_), .B(i_13_), .Y(new_new_n134_));
  NAi21      g112(.An(i_5_), .B(i_11_), .Y(new_new_n135_));
  NOi21      g113(.An(new_new_n134_), .B(new_new_n135_), .Y(new_new_n136_));
  NO2        g114(.A(i_0_), .B(i_1_), .Y(new_new_n137_));
  NA2        g115(.A(i_2_), .B(i_3_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n138_), .B(i_4_), .Y(new_new_n139_));
  NA3        g117(.A(new_new_n139_), .B(new_new_n137_), .C(new_new_n136_), .Y(new_new_n140_));
  AN2        g118(.A(new_new_n134_), .B(new_new_n76_), .Y(new_new_n141_));
  NA2        g119(.A(i_1_), .B(i_5_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n67_), .B(new_new_n46_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n36_), .Y(new_new_n144_));
  NO3        g122(.A(new_new_n144_), .B(new_new_n142_), .C(i_13_), .Y(new_new_n145_));
  OR2        g123(.A(i_0_), .B(i_1_), .Y(new_new_n146_));
  NO3        g124(.A(new_new_n146_), .B(new_new_n74_), .C(i_13_), .Y(new_new_n147_));
  NAi32      g125(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n148_));
  NAi21      g126(.An(new_new_n148_), .B(new_new_n147_), .Y(new_new_n149_));
  NOi21      g127(.An(i_4_), .B(i_10_), .Y(new_new_n150_));
  NA2        g128(.A(new_new_n150_), .B(new_new_n40_), .Y(new_new_n151_));
  NO2        g129(.A(i_3_), .B(i_5_), .Y(new_new_n152_));
  NO3        g130(.A(new_new_n67_), .B(i_2_), .C(i_1_), .Y(new_new_n153_));
  NA2        g131(.A(new_new_n153_), .B(new_new_n152_), .Y(new_new_n154_));
  OAI210     g132(.A0(new_new_n154_), .A1(new_new_n151_), .B0(new_new_n149_), .Y(new_new_n155_));
  NO2        g133(.A(new_new_n155_), .B(new_new_n145_), .Y(new_new_n156_));
  AOI210     g134(.A0(new_new_n156_), .A1(new_new_n140_), .B0(new_new_n133_), .Y(new_new_n157_));
  NA2        g135(.A(i_3_), .B(new_new_n48_), .Y(new_new_n158_));
  NOi21      g136(.An(i_4_), .B(i_9_), .Y(new_new_n159_));
  NOi21      g137(.An(i_11_), .B(i_13_), .Y(new_new_n160_));
  NA2        g138(.A(new_new_n160_), .B(new_new_n159_), .Y(new_new_n161_));
  OR2        g139(.A(new_new_n161_), .B(new_new_n158_), .Y(new_new_n162_));
  NO2        g140(.A(i_4_), .B(i_5_), .Y(new_new_n163_));
  NAi21      g141(.An(i_12_), .B(i_11_), .Y(new_new_n164_));
  NO2        g142(.A(new_new_n164_), .B(i_13_), .Y(new_new_n165_));
  NA3        g143(.A(new_new_n165_), .B(new_new_n163_), .C(new_new_n76_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(new_new_n162_), .Y(new_new_n167_));
  NO2        g145(.A(new_new_n67_), .B(new_new_n59_), .Y(new_new_n168_));
  NA2        g146(.A(new_new_n168_), .B(new_new_n46_), .Y(new_new_n169_));
  NA2        g147(.A(new_new_n36_), .B(i_5_), .Y(new_new_n170_));
  NAi31      g148(.An(new_new_n170_), .B(new_new_n141_), .C(i_11_), .Y(new_new_n171_));
  NA2        g149(.A(i_3_), .B(i_5_), .Y(new_new_n172_));
  AOI210     g150(.A0(new_new_n161_), .A1(new_new_n171_), .B0(new_new_n169_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n67_), .B(i_5_), .Y(new_new_n174_));
  NO2        g152(.A(i_13_), .B(i_10_), .Y(new_new_n175_));
  NA3        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n44_), .Y(new_new_n176_));
  NO2        g154(.A(i_2_), .B(i_1_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n177_), .B(i_3_), .Y(new_new_n178_));
  NAi21      g156(.An(i_4_), .B(i_12_), .Y(new_new_n179_));
  NO3        g157(.A(new_new_n179_), .B(new_new_n178_), .C(new_new_n176_), .Y(new_new_n180_));
  NO3        g158(.A(new_new_n180_), .B(new_new_n173_), .C(new_new_n167_), .Y(new_new_n181_));
  INV        g159(.A(i_8_), .Y(new_new_n182_));
  INV        g160(.A(i_6_), .Y(new_new_n183_));
  NO3        g161(.A(i_3_), .B(new_new_n79_), .C(new_new_n48_), .Y(new_new_n184_));
  NA2        g162(.A(new_new_n184_), .B(new_new_n105_), .Y(new_new_n185_));
  NO3        g163(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n186_));
  NA3        g164(.A(new_new_n186_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n187_));
  NO3        g165(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n188_));
  INV        g166(.A(new_new_n188_), .Y(new_new_n189_));
  AOI210     g167(.A0(new_new_n189_), .A1(new_new_n187_), .B0(new_new_n185_), .Y(new_new_n190_));
  NO2        g168(.A(i_3_), .B(i_8_), .Y(new_new_n191_));
  NO3        g169(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n192_));
  NA3        g170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n40_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n96_), .B(new_new_n56_), .Y(new_new_n194_));
  NO2        g172(.A(i_13_), .B(i_9_), .Y(new_new_n195_));
  NA3        g173(.A(new_new_n195_), .B(i_6_), .C(new_new_n182_), .Y(new_new_n196_));
  BUFFER     g174(.A(new_new_n196_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n44_), .B(i_5_), .Y(new_new_n198_));
  NO3        g176(.A(i_0_), .B(i_2_), .C(new_new_n59_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(new_new_n198_), .C(i_10_), .Y(new_new_n200_));
  OAI210     g178(.A0(new_new_n200_), .A1(new_new_n197_), .B0(new_new_n193_), .Y(new_new_n201_));
  AOI210     g179(.A0(new_new_n201_), .A1(i_7_), .B0(new_new_n190_), .Y(new_new_n202_));
  OAI220     g180(.A0(new_new_n202_), .A1(i_4_), .B0(new_new_n183_), .B1(new_new_n181_), .Y(new_new_n203_));
  NA3        g181(.A(i_13_), .B(new_new_n182_), .C(i_10_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n204_), .B(i_12_), .Y(new_new_n205_));
  NA2        g183(.A(i_0_), .B(i_5_), .Y(new_new_n206_));
  OAI220     g184(.A0(new_new_n79_), .A1(new_new_n178_), .B0(new_new_n169_), .B1(new_new_n124_), .Y(new_new_n207_));
  NAi31      g185(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n36_), .B(i_13_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n46_), .B(new_new_n59_), .Y(new_new_n210_));
  NA3        g188(.A(new_new_n210_), .B(i_3_), .C(new_new_n209_), .Y(new_new_n211_));
  INV        g189(.A(i_13_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(new_new_n212_), .Y(new_new_n213_));
  NA3        g191(.A(new_new_n213_), .B(new_new_n186_), .C(new_new_n184_), .Y(new_new_n214_));
  OAI210     g192(.A0(new_new_n211_), .A1(new_new_n208_), .B0(new_new_n214_), .Y(new_new_n215_));
  AOI220     g193(.A0(new_new_n215_), .A1(new_new_n132_), .B0(new_new_n207_), .B1(new_new_n205_), .Y(new_new_n216_));
  NO2        g194(.A(i_12_), .B(new_new_n37_), .Y(new_new_n217_));
  NO2        g195(.A(new_new_n172_), .B(i_4_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  OR2        g197(.A(i_8_), .B(i_7_), .Y(new_new_n220_));
  NO2        g198(.A(new_new_n220_), .B(new_new_n79_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n53_), .B(i_1_), .Y(new_new_n222_));
  NA2        g200(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n223_));
  INV        g201(.A(i_12_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n44_), .B(new_new_n224_), .Y(new_new_n225_));
  NO3        g203(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n226_));
  NA2        g204(.A(i_2_), .B(i_1_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n223_), .B(new_new_n219_), .Y(new_new_n228_));
  NAi21      g206(.An(i_4_), .B(i_3_), .Y(new_new_n229_));
  INV        g207(.A(new_new_n69_), .Y(new_new_n230_));
  NO2        g208(.A(i_0_), .B(i_6_), .Y(new_new_n231_));
  NOi41      g209(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n227_), .B(new_new_n172_), .Y(new_new_n234_));
  NAi21      g212(.An(new_new_n233_), .B(new_new_n234_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n235_), .Y(new_new_n236_));
  AOI210     g214(.A0(new_new_n236_), .A1(new_new_n40_), .B0(new_new_n228_), .Y(new_new_n237_));
  NO2        g215(.A(i_11_), .B(new_new_n212_), .Y(new_new_n238_));
  NOi21      g216(.An(i_1_), .B(i_6_), .Y(new_new_n239_));
  NAi21      g217(.An(i_3_), .B(i_7_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n224_), .B(i_9_), .Y(new_new_n241_));
  NO2        g219(.A(i_12_), .B(i_3_), .Y(new_new_n242_));
  NA3        g220(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n243_));
  INV        g221(.A(new_new_n133_), .Y(new_new_n244_));
  NA2        g222(.A(new_new_n224_), .B(i_13_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n245_), .B(new_new_n69_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n246_), .B(new_new_n244_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n220_), .B(new_new_n37_), .Y(new_new_n248_));
  NA2        g226(.A(i_12_), .B(i_6_), .Y(new_new_n249_));
  OR2        g227(.A(i_13_), .B(i_9_), .Y(new_new_n250_));
  NO3        g228(.A(new_new_n250_), .B(new_new_n249_), .C(new_new_n48_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n229_), .B(i_2_), .Y(new_new_n252_));
  NA3        g230(.A(new_new_n252_), .B(new_new_n251_), .C(new_new_n44_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n238_), .B(i_9_), .Y(new_new_n254_));
  OAI210     g232(.A0(new_new_n59_), .A1(new_new_n254_), .B0(new_new_n253_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n143_), .B(new_new_n59_), .Y(new_new_n256_));
  NO3        g234(.A(i_11_), .B(new_new_n212_), .C(new_new_n25_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n240_), .B(i_8_), .Y(new_new_n258_));
  NO2        g236(.A(i_6_), .B(new_new_n48_), .Y(new_new_n259_));
  NA3        g237(.A(new_new_n259_), .B(new_new_n258_), .C(new_new_n257_), .Y(new_new_n260_));
  NA3        g238(.A(i_3_), .B(new_new_n248_), .C(new_new_n213_), .Y(new_new_n261_));
  AOI210     g239(.A0(new_new_n261_), .A1(new_new_n260_), .B0(new_new_n256_), .Y(new_new_n262_));
  AOI210     g240(.A0(new_new_n255_), .A1(new_new_n248_), .B0(new_new_n262_), .Y(new_new_n263_));
  NA4        g241(.A(new_new_n263_), .B(new_new_n247_), .C(new_new_n237_), .D(new_new_n216_), .Y(new_new_n264_));
  NO3        g242(.A(i_12_), .B(new_new_n212_), .C(new_new_n37_), .Y(new_new_n265_));
  INV        g243(.A(new_new_n265_), .Y(new_new_n266_));
  NA2        g244(.A(i_8_), .B(new_new_n94_), .Y(new_new_n267_));
  NO3        g245(.A(i_0_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n268_));
  AOI220     g246(.A0(new_new_n268_), .A1(new_new_n184_), .B0(new_new_n152_), .B1(new_new_n222_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n269_), .B(new_new_n267_), .Y(new_new_n270_));
  NO3        g248(.A(i_0_), .B(i_2_), .C(new_new_n59_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n227_), .B(i_0_), .Y(new_new_n272_));
  AOI220     g250(.A0(new_new_n272_), .A1(new_new_n946_), .B0(new_new_n271_), .B1(new_new_n132_), .Y(new_new_n273_));
  NA2        g251(.A(new_new_n259_), .B(new_new_n26_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n274_), .B(new_new_n273_), .Y(new_new_n275_));
  NA2        g253(.A(i_0_), .B(i_1_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(i_2_), .Y(new_new_n277_));
  NO2        g255(.A(new_new_n57_), .B(i_6_), .Y(new_new_n278_));
  NA3        g256(.A(new_new_n278_), .B(new_new_n277_), .C(new_new_n152_), .Y(new_new_n279_));
  OAI210     g257(.A0(new_new_n154_), .A1(new_new_n133_), .B0(new_new_n279_), .Y(new_new_n280_));
  NO3        g258(.A(new_new_n280_), .B(new_new_n275_), .C(new_new_n270_), .Y(new_new_n281_));
  NO2        g259(.A(i_3_), .B(i_10_), .Y(new_new_n282_));
  NA3        g260(.A(new_new_n282_), .B(new_new_n40_), .C(new_new_n44_), .Y(new_new_n283_));
  NO2        g261(.A(i_2_), .B(new_new_n94_), .Y(new_new_n284_));
  NA2        g262(.A(i_1_), .B(new_new_n36_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n285_), .B(i_8_), .Y(new_new_n286_));
  INV        g264(.A(new_new_n286_), .Y(new_new_n287_));
  AN2        g265(.A(i_3_), .B(i_10_), .Y(new_new_n288_));
  NA3        g266(.A(new_new_n186_), .B(new_new_n165_), .C(new_new_n163_), .Y(new_new_n289_));
  NO2        g267(.A(i_5_), .B(new_new_n37_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n291_));
  OR2        g269(.A(new_new_n287_), .B(new_new_n283_), .Y(new_new_n292_));
  OAI220     g270(.A0(new_new_n292_), .A1(i_6_), .B0(new_new_n281_), .B1(new_new_n266_), .Y(new_new_n293_));
  NO4        g271(.A(new_new_n293_), .B(new_new_n264_), .C(new_new_n203_), .D(new_new_n157_), .Y(new_new_n294_));
  NO3        g272(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n295_));
  NO3        g273(.A(i_6_), .B(new_new_n182_), .C(i_7_), .Y(new_new_n296_));
  AOI210     g274(.A0(i_1_), .A1(new_new_n227_), .B0(new_new_n158_), .Y(new_new_n297_));
  NO2        g275(.A(i_2_), .B(i_3_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n206_), .B(i_5_), .Y(new_new_n299_));
  NA4        g277(.A(new_new_n299_), .B(new_new_n221_), .C(new_new_n298_), .D(i_1_), .Y(new_new_n300_));
  NA3        g278(.A(new_new_n272_), .B(new_new_n152_), .C(new_new_n105_), .Y(new_new_n301_));
  NAi21      g279(.An(i_8_), .B(i_7_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n302_), .B(i_6_), .Y(new_new_n303_));
  NA3        g281(.A(i_2_), .B(new_new_n303_), .C(new_new_n152_), .Y(new_new_n304_));
  NA3        g282(.A(new_new_n304_), .B(new_new_n301_), .C(new_new_n300_), .Y(new_new_n305_));
  OAI210     g283(.A0(new_new_n305_), .A1(new_new_n297_), .B0(i_4_), .Y(new_new_n306_));
  NO2        g284(.A(i_12_), .B(i_10_), .Y(new_new_n307_));
  NOi21      g285(.An(i_5_), .B(i_0_), .Y(new_new_n308_));
  NO3        g286(.A(new_new_n285_), .B(new_new_n308_), .C(new_new_n121_), .Y(new_new_n309_));
  NA4        g287(.A(new_new_n77_), .B(new_new_n36_), .C(new_new_n79_), .D(i_8_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n309_), .B(new_new_n307_), .Y(new_new_n311_));
  NO2        g289(.A(i_6_), .B(i_8_), .Y(new_new_n312_));
  NOi21      g290(.An(i_0_), .B(i_2_), .Y(new_new_n313_));
  AN2        g291(.A(new_new_n313_), .B(new_new_n312_), .Y(new_new_n314_));
  NO2        g292(.A(i_1_), .B(i_7_), .Y(new_new_n315_));
  AO220      g293(.A0(new_new_n315_), .A1(new_new_n314_), .B0(new_new_n303_), .B1(new_new_n222_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(i_4_), .Y(new_new_n317_));
  NA3        g295(.A(new_new_n317_), .B(new_new_n311_), .C(new_new_n306_), .Y(new_new_n318_));
  NO3        g296(.A(new_new_n220_), .B(new_new_n46_), .C(i_1_), .Y(new_new_n319_));
  NO3        g297(.A(new_new_n302_), .B(i_2_), .C(i_1_), .Y(new_new_n320_));
  OAI210     g298(.A0(new_new_n320_), .A1(new_new_n319_), .B0(i_6_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n239_), .B(new_new_n284_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n322_), .B(new_new_n321_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n323_), .B(i_3_), .Y(new_new_n324_));
  NO2        g302(.A(new_new_n276_), .B(new_new_n75_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n325_), .B(new_new_n123_), .Y(new_new_n326_));
  NO2        g304(.A(new_new_n87_), .B(new_new_n182_), .Y(new_new_n327_));
  AOI210     g305(.A0(new_new_n87_), .A1(new_new_n326_), .B0(i_3_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n182_), .B(i_9_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n329_), .B(new_new_n194_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n328_), .B(new_new_n275_), .Y(new_new_n331_));
  AOI210     g309(.A0(new_new_n331_), .A1(new_new_n324_), .B0(new_new_n151_), .Y(new_new_n332_));
  AOI210     g310(.A0(new_new_n318_), .A1(new_new_n295_), .B0(new_new_n332_), .Y(new_new_n333_));
  NOi32      g311(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n334_));
  INV        g312(.A(new_new_n334_), .Y(new_new_n335_));
  NAi21      g313(.An(i_0_), .B(i_6_), .Y(new_new_n336_));
  NAi21      g314(.An(i_1_), .B(i_5_), .Y(new_new_n337_));
  NA2        g315(.A(new_new_n337_), .B(new_new_n336_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n338_), .B(new_new_n25_), .Y(new_new_n339_));
  OAI210     g317(.A0(new_new_n339_), .A1(new_new_n148_), .B0(new_new_n233_), .Y(new_new_n340_));
  NAi41      g318(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n341_));
  OAI220     g319(.A0(new_new_n341_), .A1(new_new_n337_), .B0(new_new_n208_), .B1(new_new_n148_), .Y(new_new_n342_));
  AOI210     g320(.A0(new_new_n341_), .A1(new_new_n148_), .B0(new_new_n146_), .Y(new_new_n343_));
  OR2        g321(.A(new_new_n343_), .B(new_new_n342_), .Y(new_new_n344_));
  NO2        g322(.A(i_1_), .B(new_new_n94_), .Y(new_new_n345_));
  NAi21      g323(.An(i_3_), .B(i_4_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n346_), .B(i_9_), .Y(new_new_n347_));
  OAI210     g325(.A0(i_6_), .A1(new_new_n345_), .B0(new_new_n347_), .Y(new_new_n348_));
  NA2        g326(.A(i_2_), .B(i_7_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n346_), .B(i_10_), .Y(new_new_n350_));
  NA3        g328(.A(new_new_n350_), .B(new_new_n349_), .C(new_new_n231_), .Y(new_new_n351_));
  AOI210     g329(.A0(new_new_n351_), .A1(new_new_n348_), .B0(new_new_n174_), .Y(new_new_n352_));
  AOI210     g330(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n353_));
  OAI210     g331(.A0(new_new_n353_), .A1(new_new_n177_), .B0(new_new_n350_), .Y(new_new_n354_));
  AOI220     g332(.A0(new_new_n350_), .A1(new_new_n315_), .B0(new_new_n226_), .B1(new_new_n177_), .Y(new_new_n355_));
  AOI210     g333(.A0(new_new_n355_), .A1(new_new_n354_), .B0(i_5_), .Y(new_new_n356_));
  NO4        g334(.A(new_new_n356_), .B(new_new_n352_), .C(new_new_n344_), .D(new_new_n340_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(new_new_n335_), .Y(new_new_n358_));
  NO2        g336(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n359_));
  AN2        g337(.A(i_12_), .B(i_5_), .Y(new_new_n360_));
  NO2        g338(.A(i_4_), .B(new_new_n26_), .Y(new_new_n361_));
  NA2        g339(.A(new_new_n361_), .B(new_new_n360_), .Y(new_new_n362_));
  NO2        g340(.A(i_11_), .B(i_6_), .Y(new_new_n363_));
  NA3        g341(.A(new_new_n363_), .B(i_2_), .C(new_new_n212_), .Y(new_new_n364_));
  NO2        g342(.A(new_new_n364_), .B(new_new_n362_), .Y(new_new_n365_));
  INV        g343(.A(i_5_), .Y(new_new_n366_));
  NO2        g344(.A(i_5_), .B(i_10_), .Y(new_new_n367_));
  AOI220     g345(.A0(new_new_n367_), .A1(new_new_n252_), .B0(new_new_n366_), .B1(new_new_n186_), .Y(new_new_n368_));
  NA2        g346(.A(new_new_n134_), .B(new_new_n45_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(new_new_n368_), .Y(new_new_n370_));
  OAI210     g348(.A0(new_new_n370_), .A1(new_new_n365_), .B0(new_new_n359_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n372_));
  NO2        g350(.A(new_new_n140_), .B(new_new_n79_), .Y(new_new_n373_));
  OAI210     g351(.A0(new_new_n373_), .A1(new_new_n365_), .B0(new_new_n372_), .Y(new_new_n374_));
  NO3        g352(.A(new_new_n79_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n375_));
  NA2        g353(.A(new_new_n367_), .B(new_new_n224_), .Y(new_new_n376_));
  OAI210     g354(.A0(new_new_n376_), .A1(new_new_n310_), .B0(new_new_n208_), .Y(new_new_n377_));
  NAi21      g355(.An(i_13_), .B(i_0_), .Y(new_new_n378_));
  NO2        g356(.A(new_new_n378_), .B(new_new_n227_), .Y(new_new_n379_));
  NA2        g357(.A(new_new_n377_), .B(new_new_n379_), .Y(new_new_n380_));
  NA3        g358(.A(new_new_n380_), .B(new_new_n374_), .C(new_new_n371_), .Y(new_new_n381_));
  NA2        g359(.A(new_new_n44_), .B(new_new_n212_), .Y(new_new_n382_));
  NO2        g360(.A(i_0_), .B(i_11_), .Y(new_new_n383_));
  INV        g361(.A(i_5_), .Y(new_new_n384_));
  AN2        g362(.A(i_1_), .B(i_6_), .Y(new_new_n385_));
  NOi21      g363(.An(i_2_), .B(i_12_), .Y(new_new_n386_));
  NA2        g364(.A(new_new_n386_), .B(new_new_n385_), .Y(new_new_n387_));
  NO2        g365(.A(new_new_n387_), .B(new_new_n384_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n132_), .B(i_9_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(i_4_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n388_), .B(new_new_n390_), .Y(new_new_n391_));
  NAi21      g369(.An(i_9_), .B(i_4_), .Y(new_new_n392_));
  OR2        g370(.A(i_13_), .B(i_10_), .Y(new_new_n393_));
  NO3        g371(.A(new_new_n393_), .B(new_new_n110_), .C(new_new_n392_), .Y(new_new_n394_));
  BUFFER     g372(.A(new_new_n204_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n94_), .B(new_new_n25_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n259_), .B(new_new_n199_), .Y(new_new_n397_));
  NO2        g375(.A(new_new_n397_), .B(new_new_n395_), .Y(new_new_n398_));
  INV        g376(.A(new_new_n398_), .Y(new_new_n399_));
  AOI210     g377(.A0(new_new_n399_), .A1(new_new_n391_), .B0(new_new_n26_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n301_), .B(new_new_n300_), .Y(new_new_n401_));
  AOI220     g379(.A0(new_new_n278_), .A1(new_new_n268_), .B0(new_new_n272_), .B1(i_6_), .Y(new_new_n402_));
  NO2        g380(.A(new_new_n402_), .B(new_new_n158_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n172_), .B(new_new_n79_), .Y(new_new_n404_));
  AOI220     g382(.A0(new_new_n404_), .A1(new_new_n277_), .B0(i_3_), .B1(new_new_n199_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n405_), .B(new_new_n267_), .Y(new_new_n406_));
  NO3        g384(.A(new_new_n406_), .B(new_new_n403_), .C(new_new_n401_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n184_), .B(new_new_n89_), .Y(new_new_n408_));
  NA3        g386(.A(i_2_), .B(new_new_n152_), .C(new_new_n79_), .Y(new_new_n409_));
  AOI210     g387(.A0(new_new_n409_), .A1(new_new_n408_), .B0(new_new_n302_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n278_), .B(new_new_n222_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n411_), .B(new_new_n172_), .Y(new_new_n412_));
  NA3        g390(.A(new_new_n315_), .B(new_new_n314_), .C(i_5_), .Y(new_new_n413_));
  INV        g391(.A(new_new_n296_), .Y(new_new_n414_));
  OAI210     g392(.A0(new_new_n414_), .A1(new_new_n178_), .B0(new_new_n413_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n412_), .C(new_new_n410_), .Y(new_new_n416_));
  AOI210     g394(.A0(new_new_n416_), .A1(new_new_n407_), .B0(new_new_n254_), .Y(new_new_n417_));
  NO4        g395(.A(new_new_n417_), .B(new_new_n400_), .C(new_new_n381_), .D(new_new_n358_), .Y(new_new_n418_));
  NO2        g396(.A(new_new_n67_), .B(i_13_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n419_), .B(i_2_), .Y(new_new_n420_));
  NO2        g398(.A(i_10_), .B(i_9_), .Y(new_new_n421_));
  NAi21      g399(.An(i_12_), .B(i_8_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n422_), .B(i_3_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n423_), .B(new_new_n421_), .Y(new_new_n424_));
  NA2        g402(.A(i_2_), .B(new_new_n97_), .Y(new_new_n425_));
  OAI220     g403(.A0(new_new_n425_), .A1(new_new_n193_), .B0(new_new_n424_), .B1(new_new_n420_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n291_), .B(i_0_), .Y(new_new_n427_));
  NO3        g405(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n249_), .B(new_new_n90_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NA2        g408(.A(i_8_), .B(i_9_), .Y(new_new_n431_));
  NO2        g409(.A(i_7_), .B(i_2_), .Y(new_new_n432_));
  OR2        g410(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n265_), .B(new_new_n194_), .Y(new_new_n434_));
  NO2        g412(.A(new_new_n434_), .B(new_new_n433_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n238_), .B(new_new_n290_), .Y(new_new_n436_));
  NO3        g414(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n437_));
  INV        g415(.A(new_new_n437_), .Y(new_new_n438_));
  NA3        g416(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n439_));
  NA3        g417(.A(new_new_n135_), .B(new_new_n108_), .C(new_new_n23_), .Y(new_new_n440_));
  OAI220     g418(.A0(new_new_n440_), .A1(new_new_n439_), .B0(new_new_n438_), .B1(new_new_n436_), .Y(new_new_n441_));
  NO3        g419(.A(new_new_n441_), .B(new_new_n435_), .C(new_new_n426_), .Y(new_new_n442_));
  OR2        g420(.A(new_new_n276_), .B(new_new_n196_), .Y(new_new_n443_));
  OA210      g421(.A0(new_new_n330_), .A1(new_new_n94_), .B0(new_new_n279_), .Y(new_new_n444_));
  OA220      g422(.A0(new_new_n444_), .A1(new_new_n151_), .B0(new_new_n443_), .B1(new_new_n219_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n89_), .B(i_13_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n404_), .B(new_new_n359_), .Y(new_new_n447_));
  NO2        g425(.A(i_2_), .B(i_13_), .Y(new_new_n448_));
  NA3        g426(.A(new_new_n448_), .B(new_new_n150_), .C(new_new_n92_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n447_), .B(new_new_n446_), .Y(new_new_n450_));
  NO3        g428(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n451_));
  NO2        g429(.A(i_6_), .B(i_7_), .Y(new_new_n452_));
  OR2        g430(.A(i_11_), .B(i_8_), .Y(new_new_n453_));
  NOi21      g431(.An(i_2_), .B(i_7_), .Y(new_new_n454_));
  NAi31      g432(.An(new_new_n453_), .B(new_new_n454_), .C(new_new_n945_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n393_), .B(i_6_), .Y(new_new_n456_));
  NA2        g434(.A(new_new_n456_), .B(new_new_n950_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n457_), .B(new_new_n455_), .Y(new_new_n458_));
  NO2        g436(.A(i_3_), .B(new_new_n182_), .Y(new_new_n459_));
  NO2        g437(.A(i_6_), .B(i_10_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n461_));
  NO2        g439(.A(new_new_n146_), .B(i_3_), .Y(new_new_n462_));
  NAi31      g440(.An(new_new_n461_), .B(new_new_n462_), .C(new_new_n213_), .Y(new_new_n463_));
  NA3        g441(.A(new_new_n372_), .B(new_new_n168_), .C(new_new_n139_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n464_), .B(new_new_n463_), .Y(new_new_n465_));
  NO3        g443(.A(new_new_n465_), .B(new_new_n458_), .C(new_new_n450_), .Y(new_new_n466_));
  NA2        g444(.A(new_new_n428_), .B(new_new_n360_), .Y(new_new_n467_));
  NA2        g445(.A(new_new_n437_), .B(new_new_n367_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n468_), .B(new_new_n211_), .Y(new_new_n469_));
  NO2        g447(.A(i_0_), .B(new_new_n79_), .Y(new_new_n470_));
  NA3        g448(.A(new_new_n470_), .B(i_3_), .C(new_new_n132_), .Y(new_new_n471_));
  OR3        g449(.A(new_new_n285_), .B(new_new_n38_), .C(new_new_n46_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n472_), .B(new_new_n471_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n27_), .B(i_10_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n446_), .Y(new_new_n475_));
  NO3        g453(.A(new_new_n475_), .B(new_new_n473_), .C(new_new_n469_), .Y(new_new_n476_));
  NA4        g454(.A(new_new_n476_), .B(new_new_n466_), .C(new_new_n445_), .D(new_new_n442_), .Y(new_new_n477_));
  NA3        g455(.A(new_new_n288_), .B(new_new_n165_), .C(new_new_n163_), .Y(new_new_n478_));
  INV        g456(.A(new_new_n478_), .Y(new_new_n479_));
  BUFFER     g457(.A(new_new_n221_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n480_), .B(new_new_n479_), .Y(new_new_n481_));
  NA2        g459(.A(new_new_n115_), .B(new_new_n104_), .Y(new_new_n482_));
  AN2        g460(.A(new_new_n482_), .B(new_new_n428_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n295_), .B(new_new_n153_), .Y(new_new_n484_));
  OAI210     g462(.A0(new_new_n484_), .A1(new_new_n219_), .B0(new_new_n289_), .Y(new_new_n485_));
  AOI220     g463(.A0(new_new_n485_), .A1(new_new_n303_), .B0(new_new_n483_), .B1(new_new_n291_), .Y(new_new_n486_));
  NA4        g464(.A(new_new_n419_), .B(new_new_n950_), .C(new_new_n191_), .D(i_2_), .Y(new_new_n487_));
  INV        g465(.A(new_new_n487_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n334_), .B(new_new_n67_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n36_), .B(i_8_), .Y(new_new_n490_));
  AOI210     g468(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n394_), .Y(new_new_n491_));
  INV        g469(.A(new_new_n491_), .Y(new_new_n492_));
  AOI210     g470(.A0(new_new_n488_), .A1(new_new_n192_), .B0(new_new_n492_), .Y(new_new_n493_));
  NO2        g471(.A(i_7_), .B(new_new_n187_), .Y(new_new_n494_));
  OR2        g472(.A(new_new_n172_), .B(i_4_), .Y(new_new_n495_));
  INV        g473(.A(new_new_n495_), .Y(new_new_n496_));
  NA2        g474(.A(new_new_n496_), .B(new_new_n494_), .Y(new_new_n497_));
  NA4        g475(.A(new_new_n497_), .B(new_new_n493_), .C(new_new_n486_), .D(new_new_n481_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n366_), .B(new_new_n277_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n362_), .B(new_new_n499_), .Y(new_new_n500_));
  NO2        g478(.A(i_12_), .B(new_new_n182_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n501_), .B(new_new_n212_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n460_), .B(new_new_n27_), .Y(new_new_n503_));
  NO2        g481(.A(new_new_n503_), .B(new_new_n502_), .Y(new_new_n504_));
  NOi21      g482(.An(new_new_n296_), .B(new_new_n38_), .Y(new_new_n505_));
  OAI210     g483(.A0(new_new_n505_), .A1(new_new_n504_), .B0(new_new_n500_), .Y(new_new_n506_));
  NO2        g484(.A(i_8_), .B(i_7_), .Y(new_new_n507_));
  INV        g485(.A(new_new_n210_), .Y(new_new_n508_));
  OAI220     g486(.A0(new_new_n46_), .A1(new_new_n495_), .B0(new_new_n508_), .B1(new_new_n229_), .Y(new_new_n509_));
  NO2        g487(.A(new_new_n949_), .B(i_6_), .Y(new_new_n510_));
  NA3        g488(.A(new_new_n510_), .B(new_new_n509_), .C(new_new_n507_), .Y(new_new_n511_));
  AOI220     g489(.A0(new_new_n404_), .A1(i_2_), .B0(new_new_n234_), .B1(new_new_n231_), .Y(new_new_n512_));
  OAI220     g490(.A0(new_new_n512_), .A1(new_new_n245_), .B0(new_new_n446_), .B1(new_new_n124_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n513_), .B(new_new_n248_), .Y(new_new_n514_));
  NA3        g492(.A(new_new_n288_), .B(new_new_n163_), .C(new_new_n89_), .Y(new_new_n515_));
  NO2        g493(.A(new_new_n209_), .B(new_new_n44_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n146_), .B(i_5_), .Y(new_new_n517_));
  NA2        g495(.A(new_new_n517_), .B(new_new_n382_), .Y(new_new_n518_));
  NO2        g496(.A(new_new_n518_), .B(new_new_n516_), .Y(new_new_n519_));
  NA2        g497(.A(new_new_n519_), .B(new_new_n437_), .Y(new_new_n520_));
  NA4        g498(.A(new_new_n520_), .B(new_new_n514_), .C(new_new_n511_), .D(new_new_n506_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n206_), .B(new_new_n65_), .C(new_new_n44_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n265_), .B(new_new_n77_), .Y(new_new_n523_));
  AOI210     g501(.A0(new_new_n522_), .A1(new_new_n326_), .B0(new_new_n523_), .Y(new_new_n524_));
  AOI210     g502(.A0(i_6_), .A1(new_new_n46_), .B0(new_new_n345_), .Y(new_new_n525_));
  NA2        g503(.A(new_new_n501_), .B(new_new_n257_), .Y(new_new_n526_));
  NO2        g504(.A(new_new_n525_), .B(new_new_n526_), .Y(new_new_n527_));
  NO2        g505(.A(new_new_n527_), .B(new_new_n524_), .Y(new_new_n528_));
  NO4        g506(.A(new_new_n239_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n529_));
  NO3        g507(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n530_));
  NO2        g508(.A(new_new_n220_), .B(new_new_n36_), .Y(new_new_n531_));
  AN2        g509(.A(new_new_n531_), .B(new_new_n530_), .Y(new_new_n532_));
  OA210      g510(.A0(new_new_n532_), .A1(new_new_n529_), .B0(new_new_n334_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n393_), .B(i_1_), .Y(new_new_n534_));
  NOi31      g512(.An(new_new_n534_), .B(new_new_n429_), .C(new_new_n67_), .Y(new_new_n535_));
  AN3        g513(.A(new_new_n535_), .B(new_new_n390_), .C(i_2_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n402_), .B(new_new_n166_), .Y(new_new_n537_));
  NO3        g515(.A(new_new_n537_), .B(new_new_n536_), .C(new_new_n533_), .Y(new_new_n538_));
  NOi21      g516(.An(i_10_), .B(i_6_), .Y(new_new_n539_));
  NA2        g517(.A(new_new_n257_), .B(new_new_n539_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n540_), .B(new_new_n427_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n107_), .B(new_new_n23_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n296_), .B(new_new_n153_), .Y(new_new_n543_));
  AOI220     g521(.A0(new_new_n543_), .A1(new_new_n411_), .B0(new_new_n161_), .B1(new_new_n171_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n186_), .B(new_new_n37_), .Y(new_new_n545_));
  NOi31      g523(.An(new_new_n136_), .B(new_new_n545_), .C(new_new_n310_), .Y(new_new_n546_));
  NO3        g524(.A(new_new_n546_), .B(new_new_n544_), .C(new_new_n541_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n489_), .B(new_new_n355_), .Y(new_new_n548_));
  NO2        g526(.A(i_12_), .B(new_new_n79_), .Y(new_new_n549_));
  NO3        g527(.A(i_4_), .B(new_new_n321_), .C(new_new_n283_), .Y(new_new_n550_));
  BUFFER     g528(.A(i_5_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n550_), .B(new_new_n548_), .Y(new_new_n552_));
  NA4        g530(.A(new_new_n552_), .B(new_new_n547_), .C(new_new_n538_), .D(new_new_n528_), .Y(new_new_n553_));
  NO4        g531(.A(new_new_n553_), .B(new_new_n521_), .C(new_new_n498_), .D(new_new_n477_), .Y(new_new_n554_));
  NA4        g532(.A(new_new_n554_), .B(new_new_n418_), .C(new_new_n333_), .D(new_new_n294_), .Y(mai7));
  NO2        g533(.A(new_new_n101_), .B(new_new_n84_), .Y(new_new_n556_));
  NA2        g534(.A(new_new_n460_), .B(new_new_n77_), .Y(new_new_n557_));
  NA3        g535(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n224_), .B(i_4_), .Y(new_new_n559_));
  NA2        g537(.A(new_new_n559_), .B(i_8_), .Y(new_new_n560_));
  NO2        g538(.A(new_new_n98_), .B(new_new_n558_), .Y(new_new_n561_));
  OAI210     g539(.A0(new_new_n82_), .A1(new_new_n191_), .B0(new_new_n192_), .Y(new_new_n562_));
  NO2        g540(.A(i_7_), .B(new_new_n37_), .Y(new_new_n563_));
  NO2        g541(.A(new_new_n562_), .B(i_13_), .Y(new_new_n564_));
  NO3        g542(.A(new_new_n564_), .B(new_new_n561_), .C(new_new_n556_), .Y(new_new_n565_));
  AOI210     g543(.A0(new_new_n121_), .A1(new_new_n58_), .B0(i_10_), .Y(new_new_n566_));
  AOI210     g544(.A0(new_new_n566_), .A1(new_new_n224_), .B0(new_new_n150_), .Y(new_new_n567_));
  NO2        g545(.A(i_10_), .B(new_new_n23_), .Y(new_new_n568_));
  OR3        g546(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n569_));
  NO3        g547(.A(new_new_n569_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n570_));
  INV        g548(.A(new_new_n188_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n570_), .B(new_new_n568_), .Y(new_new_n572_));
  OA220      g550(.A0(new_new_n572_), .A1(i_2_), .B0(new_new_n567_), .B1(new_new_n250_), .Y(new_new_n573_));
  AOI210     g551(.A0(new_new_n573_), .A1(new_new_n565_), .B0(new_new_n59_), .Y(new_new_n574_));
  NOi21      g552(.An(i_11_), .B(i_7_), .Y(new_new_n575_));
  AO210      g553(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n576_));
  NO2        g554(.A(new_new_n576_), .B(new_new_n575_), .Y(new_new_n577_));
  NA2        g555(.A(new_new_n577_), .B(new_new_n195_), .Y(new_new_n578_));
  NA3        g556(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n578_), .B(new_new_n59_), .Y(new_new_n580_));
  AO210      g558(.A0(new_new_n80_), .A1(new_new_n355_), .B0(new_new_n41_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n213_), .B(new_new_n59_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n59_), .B(i_9_), .Y(new_new_n583_));
  NO2        g561(.A(i_1_), .B(i_12_), .Y(new_new_n584_));
  NA2        g562(.A(new_new_n582_), .B(new_new_n581_), .Y(new_new_n585_));
  OAI210     g563(.A0(new_new_n585_), .A1(new_new_n580_), .B0(i_6_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n579_), .B(new_new_n101_), .Y(new_new_n587_));
  NA2        g565(.A(new_new_n587_), .B(new_new_n549_), .Y(new_new_n588_));
  NO2        g566(.A(i_6_), .B(i_11_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n588_), .B(new_new_n430_), .Y(new_new_n590_));
  NO4        g568(.A(i_12_), .B(new_new_n121_), .C(i_13_), .D(new_new_n79_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n583_), .Y(new_new_n592_));
  NO3        g570(.A(i_10_), .B(new_new_n220_), .C(new_new_n23_), .Y(new_new_n593_));
  INV        g571(.A(new_new_n592_), .Y(new_new_n594_));
  NA3        g572(.A(new_new_n507_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n128_), .B(i_9_), .Y(new_new_n596_));
  NA2        g574(.A(i_3_), .B(i_9_), .Y(new_new_n597_));
  NO2        g575(.A(new_new_n596_), .B(new_new_n944_), .Y(new_new_n598_));
  NA3        g576(.A(new_new_n583_), .B(new_new_n298_), .C(i_6_), .Y(new_new_n599_));
  NO2        g577(.A(new_new_n599_), .B(new_new_n23_), .Y(new_new_n600_));
  NO2        g578(.A(i_11_), .B(new_new_n37_), .Y(new_new_n601_));
  NA2        g579(.A(new_new_n601_), .B(new_new_n24_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n602_), .B(i_6_), .Y(new_new_n603_));
  OR3        g581(.A(new_new_n603_), .B(new_new_n600_), .C(new_new_n598_), .Y(new_new_n604_));
  NO3        g582(.A(new_new_n604_), .B(new_new_n594_), .C(new_new_n590_), .Y(new_new_n605_));
  NO2        g583(.A(new_new_n392_), .B(new_new_n79_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n220_), .B(new_new_n44_), .Y(new_new_n607_));
  NO3        g585(.A(new_new_n607_), .B(new_new_n291_), .C(new_new_n225_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n110_), .B(new_new_n37_), .Y(new_new_n609_));
  NO2        g587(.A(new_new_n609_), .B(i_6_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n79_), .B(i_9_), .Y(new_new_n611_));
  NO2        g589(.A(new_new_n611_), .B(new_new_n59_), .Y(new_new_n612_));
  NO2        g590(.A(new_new_n612_), .B(new_new_n584_), .Y(new_new_n613_));
  NO4        g591(.A(new_new_n613_), .B(new_new_n610_), .C(new_new_n608_), .D(i_4_), .Y(new_new_n614_));
  NA2        g592(.A(i_1_), .B(i_3_), .Y(new_new_n615_));
  INV        g593(.A(new_new_n614_), .Y(new_new_n616_));
  NA3        g594(.A(new_new_n616_), .B(new_new_n605_), .C(new_new_n586_), .Y(new_new_n617_));
  NO3        g595(.A(new_new_n453_), .B(i_3_), .C(i_7_), .Y(new_new_n618_));
  OA210      g596(.A0(new_new_n618_), .A1(new_new_n232_), .B0(new_new_n79_), .Y(new_new_n619_));
  NA3        g597(.A(new_new_n150_), .B(new_new_n77_), .C(new_new_n79_), .Y(new_new_n620_));
  INV        g598(.A(new_new_n620_), .Y(new_new_n621_));
  OAI210     g599(.A0(new_new_n621_), .A1(new_new_n619_), .B0(i_1_), .Y(new_new_n622_));
  AOI210     g600(.A0(new_new_n249_), .A1(new_new_n90_), .B0(i_1_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n346_), .B(i_2_), .Y(new_new_n624_));
  NA2        g602(.A(new_new_n624_), .B(new_new_n623_), .Y(new_new_n625_));
  AOI210     g603(.A0(new_new_n625_), .A1(new_new_n622_), .B0(i_13_), .Y(new_new_n626_));
  OR2        g604(.A(i_11_), .B(i_7_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n99_), .B(new_new_n128_), .Y(new_new_n628_));
  AOI220     g606(.A0(new_new_n448_), .A1(new_new_n150_), .B0(i_2_), .B1(new_new_n128_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n629_), .B(new_new_n628_), .Y(new_new_n630_));
  NO2        g608(.A(new_new_n54_), .B(i_12_), .Y(new_new_n631_));
  INV        g609(.A(new_new_n631_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n454_), .B(new_new_n24_), .Y(new_new_n633_));
  NA2        g611(.A(new_new_n633_), .B(new_new_n606_), .Y(new_new_n634_));
  OAI220     g612(.A0(new_new_n634_), .A1(new_new_n41_), .B0(new_new_n632_), .B1(new_new_n87_), .Y(new_new_n635_));
  AOI210     g613(.A0(new_new_n630_), .A1(new_new_n312_), .B0(new_new_n635_), .Y(new_new_n636_));
  INV        g614(.A(new_new_n107_), .Y(new_new_n637_));
  AOI220     g615(.A0(new_new_n637_), .A1(new_new_n66_), .B0(new_new_n363_), .B1(new_new_n951_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n229_), .Y(new_new_n639_));
  AOI210     g617(.A0(new_new_n422_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n640_));
  NOi21      g618(.An(new_new_n640_), .B(new_new_n557_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n120_), .B(i_13_), .Y(new_new_n642_));
  NO2        g620(.A(new_new_n597_), .B(new_new_n107_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n642_), .B(new_new_n623_), .Y(new_new_n644_));
  AOI220     g622(.A0(new_new_n363_), .A1(new_new_n951_), .B0(new_new_n86_), .B1(new_new_n95_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n560_), .Y(new_new_n646_));
  NO4        g624(.A(new_new_n646_), .B(new_new_n644_), .C(new_new_n641_), .D(new_new_n639_), .Y(new_new_n647_));
  OR2        g625(.A(i_11_), .B(i_6_), .Y(new_new_n648_));
  NO2        g626(.A(new_new_n597_), .B(new_new_n648_), .Y(new_new_n649_));
  NA3        g627(.A(new_new_n386_), .B(new_new_n563_), .C(new_new_n90_), .Y(new_new_n650_));
  NA2        g628(.A(new_new_n589_), .B(i_13_), .Y(new_new_n651_));
  NAi21      g629(.An(i_11_), .B(i_12_), .Y(new_new_n652_));
  NA2        g630(.A(new_new_n651_), .B(new_new_n650_), .Y(new_new_n653_));
  OAI210     g631(.A0(new_new_n653_), .A1(new_new_n649_), .B0(new_new_n59_), .Y(new_new_n654_));
  NO2        g632(.A(i_2_), .B(i_12_), .Y(new_new_n655_));
  NA2        g633(.A(new_new_n345_), .B(new_new_n655_), .Y(new_new_n656_));
  NO3        g634(.A(i_9_), .B(new_new_n361_), .C(new_new_n559_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n657_), .B(new_new_n345_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n121_), .B(i_2_), .Y(new_new_n659_));
  NA2        g637(.A(new_new_n659_), .B(new_new_n584_), .Y(new_new_n660_));
  NA3        g638(.A(new_new_n660_), .B(new_new_n658_), .C(new_new_n656_), .Y(new_new_n661_));
  NA3        g639(.A(new_new_n661_), .B(new_new_n45_), .C(new_new_n212_), .Y(new_new_n662_));
  NA4        g640(.A(new_new_n662_), .B(new_new_n654_), .C(new_new_n647_), .D(new_new_n636_), .Y(new_new_n663_));
  OR4        g641(.A(new_new_n663_), .B(new_new_n626_), .C(new_new_n617_), .D(new_new_n574_), .Y(mai5));
  AN2        g642(.A(new_new_n24_), .B(i_10_), .Y(new_new_n665_));
  NA3        g643(.A(new_new_n665_), .B(new_new_n655_), .C(new_new_n101_), .Y(new_new_n666_));
  INV        g644(.A(new_new_n666_), .Y(new_new_n667_));
  NO3        g645(.A(i_11_), .B(new_new_n224_), .C(i_13_), .Y(new_new_n668_));
  NO2        g646(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n669_));
  NA2        g647(.A(i_12_), .B(i_8_), .Y(new_new_n670_));
  INV        g648(.A(new_new_n421_), .Y(new_new_n671_));
  NA2        g649(.A(i_2_), .B(new_new_n669_), .Y(new_new_n672_));
  INV        g650(.A(new_new_n672_), .Y(new_new_n673_));
  NO2        g651(.A(new_new_n673_), .B(new_new_n667_), .Y(new_new_n674_));
  INV        g652(.A(new_new_n160_), .Y(new_new_n675_));
  INV        g653(.A(new_new_n232_), .Y(new_new_n676_));
  OAI210     g654(.A0(new_new_n624_), .A1(new_new_n423_), .B0(new_new_n103_), .Y(new_new_n677_));
  AOI210     g655(.A0(new_new_n677_), .A1(new_new_n676_), .B0(new_new_n675_), .Y(new_new_n678_));
  NO2        g656(.A(new_new_n431_), .B(new_new_n26_), .Y(new_new_n679_));
  INV        g657(.A(new_new_n678_), .Y(new_new_n680_));
  INV        g658(.A(new_new_n161_), .Y(new_new_n681_));
  NO3        g659(.A(new_new_n576_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n682_));
  AOI210     g660(.A0(new_new_n681_), .A1(new_new_n82_), .B0(new_new_n682_), .Y(new_new_n683_));
  NO2        g661(.A(new_new_n683_), .B(new_new_n182_), .Y(new_new_n684_));
  OA210      g662(.A0(new_new_n577_), .A1(new_new_n119_), .B0(i_13_), .Y(new_new_n685_));
  INV        g663(.A(new_new_n141_), .Y(new_new_n686_));
  NO2        g664(.A(new_new_n686_), .B(new_new_n349_), .Y(new_new_n687_));
  NO2        g665(.A(new_new_n138_), .B(new_new_n490_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n688_), .B(new_new_n396_), .Y(new_new_n689_));
  NO2        g667(.A(new_new_n95_), .B(new_new_n44_), .Y(new_new_n690_));
  INV        g668(.A(new_new_n284_), .Y(new_new_n691_));
  NA4        g669(.A(new_new_n691_), .B(new_new_n288_), .C(new_new_n117_), .D(new_new_n42_), .Y(new_new_n692_));
  OAI210     g670(.A0(new_new_n692_), .A1(new_new_n690_), .B0(new_new_n689_), .Y(new_new_n693_));
  NO4        g671(.A(new_new_n693_), .B(new_new_n687_), .C(new_new_n685_), .D(new_new_n684_), .Y(new_new_n694_));
  INV        g672(.A(new_new_n542_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n668_), .B(new_new_n258_), .Y(new_new_n696_));
  NA2        g674(.A(new_new_n696_), .B(new_new_n695_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n58_), .B(i_12_), .Y(new_new_n698_));
  AOI220     g676(.A0(new_new_n698_), .A1(new_new_n36_), .B0(new_new_n697_), .B1(new_new_n46_), .Y(new_new_n699_));
  NA4        g677(.A(new_new_n699_), .B(new_new_n694_), .C(new_new_n680_), .D(new_new_n674_), .Y(mai6));
  NO3        g678(.A(i_9_), .B(new_new_n290_), .C(i_1_), .Y(new_new_n701_));
  NO2        g679(.A(new_new_n174_), .B(new_new_n129_), .Y(new_new_n702_));
  OAI210     g680(.A0(new_new_n702_), .A1(new_new_n701_), .B0(new_new_n659_), .Y(new_new_n703_));
  NA4        g681(.A(new_new_n367_), .B(new_new_n459_), .C(new_new_n65_), .D(new_new_n94_), .Y(new_new_n704_));
  INV        g682(.A(new_new_n704_), .Y(new_new_n705_));
  NO2        g683(.A(i_11_), .B(i_9_), .Y(new_new_n706_));
  NO2        g684(.A(new_new_n705_), .B(new_new_n308_), .Y(new_new_n707_));
  AO210      g685(.A0(new_new_n707_), .A1(new_new_n703_), .B0(i_12_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n350_), .B(new_new_n315_), .Y(new_new_n709_));
  NA2        g687(.A(new_new_n549_), .B(new_new_n59_), .Y(new_new_n710_));
  NA2        g688(.A(new_new_n618_), .B(new_new_n65_), .Y(new_new_n711_));
  BUFFER     g689(.A(new_new_n80_), .Y(new_new_n712_));
  NA4        g690(.A(new_new_n712_), .B(new_new_n711_), .C(new_new_n710_), .D(new_new_n709_), .Y(new_new_n713_));
  INV        g691(.A(new_new_n185_), .Y(new_new_n714_));
  AOI220     g692(.A0(new_new_n714_), .A1(new_new_n706_), .B0(new_new_n713_), .B1(new_new_n67_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n307_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n117_), .Y(new_new_n717_));
  NA2        g695(.A(new_new_n717_), .B(new_new_n46_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n718_), .B(new_new_n716_), .Y(new_new_n719_));
  NO2        g697(.A(new_new_n239_), .B(i_9_), .Y(new_new_n720_));
  NA2        g698(.A(new_new_n720_), .B(new_new_n698_), .Y(new_new_n721_));
  NO2        g699(.A(new_new_n721_), .B(new_new_n174_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n32_), .B(i_11_), .Y(new_new_n723_));
  NA3        g701(.A(new_new_n723_), .B(new_new_n452_), .C(new_new_n367_), .Y(new_new_n724_));
  OAI210     g702(.A0(new_new_n618_), .A1(new_new_n531_), .B0(new_new_n530_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(new_new_n724_), .Y(new_new_n726_));
  OR3        g704(.A(new_new_n726_), .B(new_new_n722_), .C(new_new_n719_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n627_), .B(i_2_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n729_));
  OAI210     g707(.A0(new_new_n729_), .A1(new_new_n385_), .B0(new_new_n339_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n730_), .B(new_new_n728_), .Y(new_new_n731_));
  AO220      g709(.A0(new_new_n338_), .A1(new_new_n329_), .B0(new_new_n375_), .B1(i_8_), .Y(new_new_n732_));
  NA3        g710(.A(new_new_n732_), .B(new_new_n242_), .C(i_7_), .Y(new_new_n733_));
  BUFFER     g711(.A(new_new_n423_), .Y(new_new_n734_));
  NA3        g712(.A(new_new_n734_), .B(new_new_n137_), .C(new_new_n63_), .Y(new_new_n735_));
  AO210      g713(.A0(new_new_n468_), .A1(new_new_n671_), .B0(new_new_n36_), .Y(new_new_n736_));
  NA4        g714(.A(new_new_n736_), .B(new_new_n735_), .C(new_new_n733_), .D(new_new_n731_), .Y(new_new_n737_));
  OAI210     g715(.A0(i_6_), .A1(i_11_), .B0(new_new_n80_), .Y(new_new_n738_));
  NA2        g716(.A(new_new_n738_), .B(new_new_n530_), .Y(new_new_n739_));
  OAI210     g717(.A0(new_new_n375_), .A1(new_new_n192_), .B0(new_new_n64_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n740_), .B(new_new_n739_), .Y(new_new_n741_));
  AO210      g719(.A0(new_new_n490_), .A1(new_new_n46_), .B0(new_new_n81_), .Y(new_new_n742_));
  NA3        g720(.A(new_new_n742_), .B(new_new_n460_), .C(new_new_n206_), .Y(new_new_n743_));
  AOI210     g721(.A0(new_new_n423_), .A1(new_new_n421_), .B0(new_new_n529_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n104_), .B(new_new_n383_), .Y(new_new_n745_));
  NA2        g723(.A(new_new_n231_), .B(new_new_n46_), .Y(new_new_n746_));
  NA3        g724(.A(new_new_n745_), .B(new_new_n744_), .C(new_new_n743_), .Y(new_new_n747_));
  NO4        g725(.A(new_new_n747_), .B(new_new_n741_), .C(new_new_n737_), .D(new_new_n727_), .Y(new_new_n748_));
  NA4        g726(.A(new_new_n748_), .B(new_new_n715_), .C(new_new_n708_), .D(new_new_n357_), .Y(mai3));
  NA2        g727(.A(i_6_), .B(i_7_), .Y(new_new_n750_));
  NO2        g728(.A(new_new_n750_), .B(i_0_), .Y(new_new_n751_));
  NO2        g729(.A(i_11_), .B(new_new_n224_), .Y(new_new_n752_));
  OAI210     g730(.A0(new_new_n751_), .A1(new_new_n272_), .B0(new_new_n752_), .Y(new_new_n753_));
  INV        g731(.A(new_new_n753_), .Y(new_new_n754_));
  NO3        g732(.A(new_new_n427_), .B(new_new_n84_), .C(new_new_n44_), .Y(new_new_n755_));
  OA210      g733(.A0(new_new_n755_), .A1(new_new_n754_), .B0(new_new_n163_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n386_), .B(new_new_n45_), .Y(new_new_n757_));
  NO4        g735(.A(new_new_n353_), .B(new_new_n360_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n758_));
  NA2        g736(.A(new_new_n174_), .B(new_new_n539_), .Y(new_new_n759_));
  NOi21      g737(.An(new_new_n759_), .B(new_new_n758_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n640_), .B(new_new_n611_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n313_), .B(i_5_), .Y(new_new_n762_));
  OAI220     g740(.A0(new_new_n762_), .A1(new_new_n761_), .B0(new_new_n760_), .B1(new_new_n59_), .Y(new_new_n763_));
  NOi21      g741(.An(i_5_), .B(i_9_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n764_), .B(new_new_n419_), .Y(new_new_n765_));
  NO2        g743(.A(new_new_n164_), .B(new_new_n138_), .Y(new_new_n766_));
  NA2        g744(.A(new_new_n766_), .B(new_new_n231_), .Y(new_new_n767_));
  NO2        g745(.A(new_new_n767_), .B(new_new_n170_), .Y(new_new_n768_));
  NO3        g746(.A(new_new_n768_), .B(new_new_n763_), .C(new_new_n756_), .Y(new_new_n769_));
  NA2        g747(.A(new_new_n174_), .B(new_new_n24_), .Y(new_new_n770_));
  NO2        g748(.A(new_new_n609_), .B(new_new_n556_), .Y(new_new_n771_));
  NO2        g749(.A(new_new_n771_), .B(new_new_n770_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n295_), .B(new_new_n122_), .Y(new_new_n773_));
  NAi21      g751(.An(new_new_n151_), .B(i_5_), .Y(new_new_n774_));
  OAI220     g752(.A0(new_new_n774_), .A1(new_new_n746_), .B0(new_new_n773_), .B1(new_new_n376_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n775_), .B(new_new_n772_), .Y(new_new_n776_));
  NO2        g754(.A(new_new_n367_), .B(new_new_n276_), .Y(new_new_n777_));
  NA2        g755(.A(new_new_n777_), .B(new_new_n643_), .Y(new_new_n778_));
  INV        g756(.A(new_new_n452_), .Y(new_new_n779_));
  AN2        g757(.A(new_new_n89_), .B(new_new_n230_), .Y(new_new_n780_));
  NA2        g758(.A(new_new_n668_), .B(new_new_n308_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n602_), .B(new_new_n508_), .Y(new_new_n782_));
  NO2        g760(.A(new_new_n241_), .B(new_new_n142_), .Y(new_new_n783_));
  NA2        g761(.A(i_0_), .B(i_10_), .Y(new_new_n784_));
  AN2        g762(.A(new_new_n783_), .B(i_6_), .Y(new_new_n785_));
  NA2        g763(.A(new_new_n174_), .B(new_new_n77_), .Y(new_new_n786_));
  NA2        g764(.A(new_new_n534_), .B(i_4_), .Y(new_new_n787_));
  NA2        g765(.A(new_new_n177_), .B(new_new_n191_), .Y(new_new_n788_));
  OAI220     g766(.A0(new_new_n788_), .A1(new_new_n781_), .B0(new_new_n787_), .B1(new_new_n786_), .Y(new_new_n789_));
  NO4        g767(.A(new_new_n789_), .B(new_new_n785_), .C(new_new_n782_), .D(new_new_n780_), .Y(new_new_n790_));
  NA3        g768(.A(new_new_n790_), .B(new_new_n778_), .C(new_new_n776_), .Y(new_new_n791_));
  NA2        g769(.A(i_11_), .B(i_9_), .Y(new_new_n792_));
  NO2        g770(.A(new_new_n48_), .B(i_7_), .Y(new_new_n793_));
  NA2        g771(.A(new_new_n372_), .B(new_new_n168_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n794_), .B(new_new_n149_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n792_), .B(new_new_n67_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n164_), .B(i_0_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n452_), .B(new_new_n218_), .Y(new_new_n798_));
  NA2        g776(.A(i_6_), .B(i_4_), .Y(new_new_n799_));
  OAI220     g777(.A0(new_new_n799_), .A1(new_new_n765_), .B0(new_new_n798_), .B1(new_new_n164_), .Y(new_new_n800_));
  NO2        g778(.A(new_new_n800_), .B(new_new_n795_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n601_), .B(new_new_n114_), .Y(new_new_n802_));
  NO2        g780(.A(i_6_), .B(new_new_n802_), .Y(new_new_n803_));
  AOI210     g781(.A0(new_new_n422_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n804_));
  NA2        g782(.A(new_new_n160_), .B(new_new_n96_), .Y(new_new_n805_));
  NOi32      g783(.An(new_new_n804_), .Bn(new_new_n177_), .C(new_new_n805_), .Y(new_new_n806_));
  NA2        g784(.A(new_new_n563_), .B(new_new_n308_), .Y(new_new_n807_));
  NO2        g785(.A(new_new_n807_), .B(new_new_n757_), .Y(new_new_n808_));
  NO3        g786(.A(new_new_n808_), .B(new_new_n806_), .C(new_new_n803_), .Y(new_new_n809_));
  NOi21      g787(.An(i_7_), .B(i_5_), .Y(new_new_n810_));
  NOi31      g788(.An(new_new_n810_), .B(i_0_), .C(new_new_n652_), .Y(new_new_n811_));
  NO3        g789(.A(new_new_n378_), .B(new_new_n341_), .C(new_new_n337_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n243_), .B(i_5_), .Y(new_new_n813_));
  INV        g791(.A(new_new_n652_), .Y(new_new_n814_));
  AOI210     g792(.A0(new_new_n814_), .A1(new_new_n813_), .B0(new_new_n812_), .Y(new_new_n815_));
  NA3        g793(.A(new_new_n815_), .B(new_new_n809_), .C(new_new_n801_), .Y(new_new_n816_));
  NO2        g794(.A(new_new_n770_), .B(new_new_n227_), .Y(new_new_n817_));
  AN2        g795(.A(new_new_n312_), .B(new_new_n308_), .Y(new_new_n818_));
  AN2        g796(.A(new_new_n818_), .B(new_new_n766_), .Y(new_new_n819_));
  OAI210     g797(.A0(new_new_n819_), .A1(new_new_n817_), .B0(i_10_), .Y(new_new_n820_));
  NA3        g798(.A(new_new_n451_), .B(new_new_n386_), .C(new_new_n45_), .Y(new_new_n821_));
  OAI210     g799(.A0(new_new_n774_), .A1(new_new_n779_), .B0(new_new_n821_), .Y(new_new_n822_));
  NO2        g800(.A(new_new_n242_), .B(new_new_n46_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n796_), .B(new_new_n288_), .Y(new_new_n824_));
  OAI210     g802(.A0(new_new_n823_), .A1(new_new_n176_), .B0(new_new_n824_), .Y(new_new_n825_));
  AOI220     g803(.A0(new_new_n825_), .A1(new_new_n452_), .B0(new_new_n822_), .B1(new_new_n67_), .Y(new_new_n826_));
  NA3        g804(.A(new_new_n729_), .B(new_new_n359_), .C(i_6_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n87_), .B(new_new_n44_), .Y(new_new_n828_));
  NO2        g806(.A(new_new_n69_), .B(new_new_n670_), .Y(new_new_n829_));
  AOI220     g807(.A0(new_new_n829_), .A1(new_new_n828_), .B0(new_new_n163_), .B1(new_new_n556_), .Y(new_new_n830_));
  AOI210     g808(.A0(new_new_n830_), .A1(new_new_n827_), .B0(new_new_n47_), .Y(new_new_n831_));
  NO3        g809(.A(new_new_n551_), .B(new_new_n336_), .C(new_new_n24_), .Y(new_new_n832_));
  AOI210     g810(.A0(new_new_n633_), .A1(new_new_n517_), .B0(new_new_n832_), .Y(new_new_n833_));
  NO2        g811(.A(new_new_n558_), .B(new_new_n98_), .Y(new_new_n834_));
  NA2        g812(.A(new_new_n834_), .B(i_0_), .Y(new_new_n835_));
  OAI220     g813(.A0(new_new_n835_), .A1(new_new_n79_), .B0(new_new_n833_), .B1(new_new_n161_), .Y(new_new_n836_));
  NO3        g814(.A(new_new_n836_), .B(new_new_n831_), .C(new_new_n492_), .Y(new_new_n837_));
  NA3        g815(.A(new_new_n837_), .B(new_new_n826_), .C(new_new_n820_), .Y(new_new_n838_));
  NO3        g816(.A(new_new_n838_), .B(new_new_n816_), .C(new_new_n791_), .Y(new_new_n839_));
  NO2        g817(.A(i_0_), .B(new_new_n652_), .Y(new_new_n840_));
  NO3        g818(.A(new_new_n98_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n841_));
  AO220      g819(.A0(new_new_n841_), .A1(new_new_n44_), .B0(new_new_n840_), .B1(new_new_n163_), .Y(new_new_n842_));
  NO2        g820(.A(new_new_n710_), .B(new_new_n805_), .Y(new_new_n843_));
  AOI210     g821(.A0(new_new_n842_), .A1(new_new_n327_), .B0(new_new_n843_), .Y(new_new_n844_));
  NA3        g822(.A(new_new_n136_), .B(new_new_n611_), .C(new_new_n67_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n725_), .B(new_new_n378_), .Y(new_new_n846_));
  NA3        g824(.A(new_new_n751_), .B(i_2_), .C(new_new_n48_), .Y(new_new_n847_));
  NA2        g825(.A(new_new_n752_), .B(i_9_), .Y(new_new_n848_));
  AOI210     g826(.A0(new_new_n847_), .A1(new_new_n471_), .B0(new_new_n848_), .Y(new_new_n849_));
  NO2        g827(.A(new_new_n849_), .B(new_new_n846_), .Y(new_new_n850_));
  NA3        g828(.A(new_new_n850_), .B(new_new_n845_), .C(new_new_n844_), .Y(new_new_n851_));
  NA2        g829(.A(new_new_n818_), .B(new_new_n349_), .Y(new_new_n852_));
  AOI210     g830(.A0(new_new_n283_), .A1(new_new_n151_), .B0(new_new_n852_), .Y(new_new_n853_));
  NA2        g831(.A(new_new_n40_), .B(new_new_n44_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n793_), .B(new_new_n462_), .Y(new_new_n855_));
  AOI210     g833(.A0(new_new_n854_), .A1(new_new_n151_), .B0(new_new_n855_), .Y(new_new_n856_));
  NO2        g834(.A(new_new_n856_), .B(new_new_n853_), .Y(new_new_n857_));
  NO3        g835(.A(new_new_n784_), .B(new_new_n764_), .C(new_new_n179_), .Y(new_new_n858_));
  AOI220     g836(.A0(new_new_n858_), .A1(i_11_), .B0(new_new_n535_), .B1(new_new_n69_), .Y(new_new_n859_));
  NO3        g837(.A(new_new_n198_), .B(new_new_n360_), .C(i_0_), .Y(new_new_n860_));
  OAI210     g838(.A0(new_new_n860_), .A1(new_new_n70_), .B0(i_13_), .Y(new_new_n861_));
  INV        g839(.A(new_new_n206_), .Y(new_new_n862_));
  OAI220     g840(.A0(new_new_n502_), .A1(new_new_n129_), .B0(new_new_n947_), .B1(new_new_n571_), .Y(new_new_n863_));
  NA2        g841(.A(new_new_n863_), .B(new_new_n862_), .Y(new_new_n864_));
  NA4        g842(.A(new_new_n864_), .B(new_new_n861_), .C(new_new_n859_), .D(new_new_n857_), .Y(new_new_n865_));
  NA2        g843(.A(new_new_n810_), .B(new_new_n462_), .Y(new_new_n866_));
  INV        g844(.A(new_new_n165_), .Y(new_new_n867_));
  OR2        g845(.A(new_new_n867_), .B(new_new_n866_), .Y(new_new_n868_));
  AOI210     g846(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n164_), .Y(new_new_n869_));
  NA3        g847(.A(new_new_n568_), .B(new_new_n174_), .C(new_new_n77_), .Y(new_new_n870_));
  NA2        g848(.A(new_new_n870_), .B(new_new_n515_), .Y(new_new_n871_));
  NO3        g849(.A(new_new_n757_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n872_));
  NA2        g850(.A(new_new_n467_), .B(new_new_n449_), .Y(new_new_n873_));
  NO3        g851(.A(new_new_n873_), .B(new_new_n872_), .C(new_new_n871_), .Y(new_new_n874_));
  NA3        g852(.A(new_new_n793_), .B(new_new_n272_), .C(new_new_n217_), .Y(new_new_n875_));
  INV        g853(.A(new_new_n875_), .Y(new_new_n876_));
  NA3        g854(.A(new_new_n367_), .B(new_new_n314_), .C(new_new_n209_), .Y(new_new_n877_));
  INV        g855(.A(new_new_n877_), .Y(new_new_n878_));
  NO3        g856(.A(new_new_n792_), .B(new_new_n206_), .C(new_new_n179_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n879_), .B(new_new_n878_), .C(new_new_n876_), .Y(new_new_n880_));
  NA3        g858(.A(new_new_n880_), .B(new_new_n874_), .C(new_new_n868_), .Y(new_new_n881_));
  INV        g859(.A(new_new_n570_), .Y(new_new_n882_));
  NO3        g860(.A(new_new_n882_), .B(new_new_n948_), .C(i_3_), .Y(new_new_n883_));
  INV        g861(.A(new_new_n883_), .Y(new_new_n884_));
  NA3        g862(.A(new_new_n288_), .B(i_5_), .C(new_new_n182_), .Y(new_new_n885_));
  NA2        g863(.A(new_new_n885_), .B(new_new_n229_), .Y(new_new_n886_));
  NO4        g864(.A(new_new_n227_), .B(new_new_n198_), .C(i_0_), .D(i_12_), .Y(new_new_n887_));
  AOI220     g865(.A0(new_new_n887_), .A1(new_new_n886_), .B0(new_new_n705_), .B1(new_new_n165_), .Y(new_new_n888_));
  AN2        g866(.A(new_new_n784_), .B(new_new_n142_), .Y(new_new_n889_));
  NO3        g867(.A(new_new_n889_), .B(i_12_), .C(new_new_n595_), .Y(new_new_n890_));
  NA2        g868(.A(new_new_n890_), .B(new_new_n206_), .Y(new_new_n891_));
  NA3        g869(.A(new_new_n91_), .B(new_new_n539_), .C(i_11_), .Y(new_new_n892_));
  NO2        g870(.A(new_new_n892_), .B(new_new_n144_), .Y(new_new_n893_));
  NA2        g871(.A(new_new_n810_), .B(new_new_n448_), .Y(new_new_n894_));
  NA2        g872(.A(new_new_n60_), .B(new_new_n94_), .Y(new_new_n895_));
  OAI220     g873(.A0(new_new_n895_), .A1(new_new_n885_), .B0(new_new_n894_), .B1(new_new_n612_), .Y(new_new_n896_));
  AOI210     g874(.A0(new_new_n896_), .A1(new_new_n797_), .B0(new_new_n893_), .Y(new_new_n897_));
  NA4        g875(.A(new_new_n897_), .B(new_new_n891_), .C(new_new_n888_), .D(new_new_n884_), .Y(new_new_n898_));
  NO4        g876(.A(new_new_n898_), .B(new_new_n881_), .C(new_new_n865_), .D(new_new_n851_), .Y(new_new_n899_));
  OAI210     g877(.A0(new_new_n728_), .A1(new_new_n723_), .B0(new_new_n37_), .Y(new_new_n900_));
  NA3        g878(.A(new_new_n804_), .B(new_new_n345_), .C(i_5_), .Y(new_new_n901_));
  NA3        g879(.A(new_new_n901_), .B(new_new_n900_), .C(new_new_n567_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n902_), .B(new_new_n195_), .Y(new_new_n903_));
  NA2        g881(.A(new_new_n175_), .B(new_new_n177_), .Y(new_new_n904_));
  AO210      g882(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n904_), .Y(new_new_n905_));
  NAi31      g883(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n906_));
  NO2        g884(.A(new_new_n64_), .B(new_new_n906_), .Y(new_new_n907_));
  NO2        g885(.A(new_new_n907_), .B(new_new_n593_), .Y(new_new_n908_));
  NA2        g886(.A(new_new_n908_), .B(new_new_n905_), .Y(new_new_n909_));
  NO2        g887(.A(new_new_n439_), .B(new_new_n249_), .Y(new_new_n910_));
  NO4        g888(.A(new_new_n220_), .B(new_new_n135_), .C(new_new_n615_), .D(new_new_n37_), .Y(new_new_n911_));
  NO2        g889(.A(new_new_n911_), .B(new_new_n910_), .Y(new_new_n912_));
  OAI210     g890(.A0(new_new_n892_), .A1(new_new_n138_), .B0(new_new_n912_), .Y(new_new_n913_));
  AOI210     g891(.A0(new_new_n909_), .A1(new_new_n48_), .B0(new_new_n913_), .Y(new_new_n914_));
  AOI210     g892(.A0(new_new_n914_), .A1(new_new_n903_), .B0(new_new_n67_), .Y(new_new_n915_));
  NO2        g893(.A(new_new_n532_), .B(new_new_n356_), .Y(new_new_n916_));
  NO2        g894(.A(new_new_n916_), .B(new_new_n675_), .Y(new_new_n917_));
  INV        g895(.A(new_new_n101_), .Y(new_new_n918_));
  NA2        g896(.A(new_new_n918_), .B(new_new_n70_), .Y(new_new_n919_));
  AOI210     g897(.A0(new_new_n869_), .A1(new_new_n793_), .B0(new_new_n811_), .Y(new_new_n920_));
  AOI210     g898(.A0(new_new_n920_), .A1(new_new_n919_), .B0(new_new_n615_), .Y(new_new_n921_));
  INV        g899(.A(new_new_n243_), .Y(new_new_n922_));
  NA2        g900(.A(new_new_n922_), .B(new_new_n70_), .Y(new_new_n923_));
  NO2        g901(.A(new_new_n923_), .B(new_new_n224_), .Y(new_new_n924_));
  NA3        g902(.A(new_new_n89_), .B(new_new_n290_), .C(new_new_n31_), .Y(new_new_n925_));
  INV        g903(.A(new_new_n925_), .Y(new_new_n926_));
  NO3        g904(.A(new_new_n926_), .B(new_new_n924_), .C(new_new_n921_), .Y(new_new_n927_));
  OAI210     g905(.A0(new_new_n251_), .A1(new_new_n147_), .B0(new_new_n82_), .Y(new_new_n928_));
  NA2        g906(.A(new_new_n679_), .B(new_new_n272_), .Y(new_new_n929_));
  AOI210     g907(.A0(new_new_n929_), .A1(new_new_n928_), .B0(i_11_), .Y(new_new_n930_));
  INV        g908(.A(new_new_n195_), .Y(new_new_n931_));
  NA2        g909(.A(new_new_n153_), .B(i_5_), .Y(new_new_n932_));
  NO2        g910(.A(new_new_n931_), .B(new_new_n932_), .Y(new_new_n933_));
  NO3        g911(.A(i_9_), .B(new_new_n453_), .C(new_new_n240_), .Y(new_new_n934_));
  NO2        g912(.A(new_new_n934_), .B(new_new_n529_), .Y(new_new_n935_));
  INV        g913(.A(new_new_n342_), .Y(new_new_n936_));
  AOI210     g914(.A0(new_new_n936_), .A1(new_new_n935_), .B0(new_new_n41_), .Y(new_new_n937_));
  NO3        g915(.A(new_new_n937_), .B(new_new_n933_), .C(new_new_n930_), .Y(new_new_n938_));
  OAI210     g916(.A0(new_new_n927_), .A1(i_4_), .B0(new_new_n938_), .Y(new_new_n939_));
  NO3        g917(.A(new_new_n939_), .B(new_new_n917_), .C(new_new_n915_), .Y(new_new_n940_));
  NA4        g918(.A(new_new_n940_), .B(new_new_n899_), .C(new_new_n839_), .D(new_new_n769_), .Y(mai4));
  INV        g919(.A(i_2_), .Y(new_new_n944_));
  INV        g920(.A(i_3_), .Y(new_new_n945_));
  INV        g921(.A(i_7_), .Y(new_new_n946_));
  INV        g922(.A(i_6_), .Y(new_new_n947_));
  INV        g923(.A(i_0_), .Y(new_new_n948_));
  INV        g924(.A(i_10_), .Y(new_new_n949_));
  INV        g925(.A(i_4_), .Y(new_new_n950_));
  INV        g926(.A(i_1_), .Y(new_new_n951_));
endmodule


