// Benchmark "top" written by ABC on Thu Jun 20 14:59:17 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n748_, new_new_n749_, new_new_n750_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1010_, new_new_n1011_,
    new_new_n1012_, new_new_n1013_, new_new_n1014_, new_new_n1015_,
    new_new_n1016_, new_new_n1017_, new_new_n1018_, new_new_n1019_,
    new_new_n1020_, new_new_n1021_, new_new_n1022_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(men1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  OAI210     g027(.A0(new_new_n49_), .A1(i_3_), .B0(new_new_n47_), .Y(new_new_n50_));
  AOI210     g028(.A0(new_new_n50_), .A1(new_new_n46_), .B0(new_new_n45_), .Y(new_new_n51_));
  NA2        g029(.A(i_0_), .B(i_2_), .Y(new_new_n52_));
  NA2        g030(.A(i_7_), .B(i_9_), .Y(new_new_n53_));
  NO2        g031(.A(new_new_n53_), .B(new_new_n52_), .Y(new_new_n54_));
  NA2        g032(.A(new_new_n51_), .B(new_new_n44_), .Y(new_new_n55_));
  NA3        g033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n56_));
  NO2        g034(.A(i_1_), .B(i_6_), .Y(new_new_n57_));
  NA2        g035(.A(i_8_), .B(i_7_), .Y(new_new_n58_));
  NA2        g036(.A(i_6_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NA3        g040(.A(new_new_n62_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(new_new_n59_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n49_), .B(i_2_), .Y(new_new_n65_));
  AOI210     g043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_6_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(new_new_n25_), .Y(new_new_n68_));
  INV        g046(.A(i_0_), .Y(new_new_n69_));
  NAi21      g047(.An(i_5_), .B(i_10_), .Y(new_new_n70_));
  NA2        g048(.A(i_5_), .B(i_9_), .Y(new_new_n71_));
  AOI210     g049(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n69_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n68_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n66_), .A1(new_new_n65_), .B0(new_new_n73_), .Y(new_new_n74_));
  OAI210     g052(.A0(new_new_n74_), .A1(new_new_n64_), .B0(i_0_), .Y(new_new_n75_));
  NA2        g053(.A(i_12_), .B(i_5_), .Y(new_new_n76_));
  NA2        g054(.A(i_2_), .B(i_8_), .Y(new_new_n77_));
  NO2        g055(.A(i_3_), .B(i_9_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n79_), .B(new_new_n61_), .Y(new_new_n80_));
  INV        g058(.A(i_6_), .Y(new_new_n81_));
  OR4        g059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n82_));
  INV        g060(.A(new_new_n82_), .Y(new_new_n83_));
  NO2        g061(.A(i_2_), .B(i_7_), .Y(new_new_n84_));
  NA2        g062(.A(new_new_n80_), .B(new_new_n82_), .Y(new_new_n85_));
  NAi21      g063(.An(i_6_), .B(i_10_), .Y(new_new_n86_));
  NA2        g064(.A(i_6_), .B(i_9_), .Y(new_new_n87_));
  NA2        g065(.A(i_2_), .B(i_6_), .Y(new_new_n88_));
  NO3        g066(.A(new_new_n88_), .B(new_new_n48_), .C(new_new_n25_), .Y(new_new_n89_));
  INV        g067(.A(new_new_n89_), .Y(new_new_n90_));
  AOI210     g068(.A0(new_new_n90_), .A1(new_new_n85_), .B0(new_new_n76_), .Y(new_new_n91_));
  AN3        g069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n92_));
  NAi21      g070(.An(i_6_), .B(i_11_), .Y(new_new_n93_));
  NO2        g071(.A(i_5_), .B(i_8_), .Y(new_new_n94_));
  NOi21      g072(.An(new_new_n94_), .B(new_new_n93_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n92_), .B(new_new_n32_), .Y(new_new_n96_));
  INV        g074(.A(i_7_), .Y(new_new_n97_));
  NO2        g075(.A(i_0_), .B(i_5_), .Y(new_new_n98_));
  NO2        g076(.A(new_new_n98_), .B(new_new_n81_), .Y(new_new_n99_));
  NA2        g077(.A(i_12_), .B(i_3_), .Y(new_new_n100_));
  NAi21      g078(.An(i_7_), .B(i_11_), .Y(new_new_n101_));
  NO3        g079(.A(new_new_n101_), .B(new_new_n86_), .C(new_new_n52_), .Y(new_new_n102_));
  AN2        g080(.A(i_2_), .B(i_10_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n103_), .B(i_7_), .Y(new_new_n104_));
  OR2        g082(.A(new_new_n76_), .B(new_new_n57_), .Y(new_new_n105_));
  NO2        g083(.A(i_8_), .B(new_new_n97_), .Y(new_new_n106_));
  NO3        g084(.A(new_new_n106_), .B(new_new_n105_), .C(new_new_n104_), .Y(new_new_n107_));
  NA2        g085(.A(i_12_), .B(i_7_), .Y(new_new_n108_));
  NA2        g086(.A(i_1_), .B(i_0_), .Y(new_new_n109_));
  NA2        g087(.A(i_11_), .B(i_12_), .Y(new_new_n110_));
  OAI210     g088(.A0(new_new_n109_), .A1(new_new_n108_), .B0(new_new_n110_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(new_new_n107_), .Y(new_new_n112_));
  NAi31      g090(.An(new_new_n102_), .B(new_new_n112_), .C(new_new_n96_), .Y(new_new_n113_));
  NOi21      g091(.An(i_1_), .B(i_5_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(i_11_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n116_));
  NA2        g094(.A(i_7_), .B(new_new_n25_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n117_), .B(new_new_n116_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n118_), .B(new_new_n45_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n87_), .B(new_new_n86_), .Y(new_new_n120_));
  NAi21      g098(.An(i_3_), .B(i_8_), .Y(new_new_n121_));
  NA2        g099(.A(new_new_n121_), .B(new_new_n60_), .Y(new_new_n122_));
  NOi31      g100(.An(new_new_n122_), .B(new_new_n120_), .C(new_new_n119_), .Y(new_new_n123_));
  NO2        g101(.A(i_1_), .B(new_new_n81_), .Y(new_new_n124_));
  NO2        g102(.A(i_6_), .B(i_5_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(i_3_), .Y(new_new_n126_));
  AO210      g104(.A0(new_new_n126_), .A1(new_new_n46_), .B0(new_new_n124_), .Y(new_new_n127_));
  OAI220     g105(.A0(new_new_n127_), .A1(new_new_n101_), .B0(new_new_n123_), .B1(new_new_n115_), .Y(new_new_n128_));
  NO3        g106(.A(new_new_n128_), .B(new_new_n113_), .C(new_new_n91_), .Y(new_new_n129_));
  NA3        g107(.A(new_new_n129_), .B(new_new_n75_), .C(new_new_n55_), .Y(men2));
  NA3        g108(.A(new_new_n73_), .B(new_new_n65_), .C(new_new_n30_), .Y(men0));
  AN2        g109(.A(i_8_), .B(i_7_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n132_), .B(i_6_), .Y(new_new_n133_));
  NO2        g111(.A(i_12_), .B(i_13_), .Y(new_new_n134_));
  NAi21      g112(.An(i_5_), .B(i_11_), .Y(new_new_n135_));
  NOi21      g113(.An(new_new_n134_), .B(new_new_n135_), .Y(new_new_n136_));
  NO2        g114(.A(i_0_), .B(i_1_), .Y(new_new_n137_));
  NA2        g115(.A(i_2_), .B(i_3_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n138_), .B(i_4_), .Y(new_new_n139_));
  NA3        g117(.A(new_new_n139_), .B(new_new_n137_), .C(new_new_n136_), .Y(new_new_n140_));
  OR2        g118(.A(new_new_n140_), .B(new_new_n25_), .Y(new_new_n141_));
  AN2        g119(.A(new_new_n134_), .B(new_new_n78_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n142_), .B(new_new_n27_), .Y(new_new_n143_));
  NA2        g121(.A(i_1_), .B(i_5_), .Y(new_new_n144_));
  NO2        g122(.A(new_new_n69_), .B(new_new_n45_), .Y(new_new_n145_));
  NA2        g123(.A(new_new_n145_), .B(new_new_n36_), .Y(new_new_n146_));
  NO3        g124(.A(new_new_n146_), .B(new_new_n144_), .C(new_new_n143_), .Y(new_new_n147_));
  OR2        g125(.A(i_0_), .B(i_1_), .Y(new_new_n148_));
  NO3        g126(.A(new_new_n148_), .B(new_new_n76_), .C(i_13_), .Y(new_new_n149_));
  NAi32      g127(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n150_));
  NAi21      g128(.An(new_new_n150_), .B(new_new_n149_), .Y(new_new_n151_));
  NOi21      g129(.An(i_4_), .B(i_10_), .Y(new_new_n152_));
  NA2        g130(.A(new_new_n152_), .B(new_new_n39_), .Y(new_new_n153_));
  NO2        g131(.A(i_3_), .B(i_5_), .Y(new_new_n154_));
  NO3        g132(.A(new_new_n69_), .B(i_2_), .C(i_1_), .Y(new_new_n155_));
  NA2        g133(.A(new_new_n155_), .B(new_new_n154_), .Y(new_new_n156_));
  OAI210     g134(.A0(new_new_n156_), .A1(new_new_n153_), .B0(new_new_n151_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(new_new_n147_), .Y(new_new_n158_));
  AOI210     g136(.A0(new_new_n158_), .A1(new_new_n141_), .B0(new_new_n133_), .Y(new_new_n159_));
  NA2        g137(.A(i_3_), .B(new_new_n47_), .Y(new_new_n160_));
  NOi21      g138(.An(i_4_), .B(i_9_), .Y(new_new_n161_));
  NOi21      g139(.An(i_11_), .B(i_13_), .Y(new_new_n162_));
  NA2        g140(.A(new_new_n162_), .B(new_new_n161_), .Y(new_new_n163_));
  OR2        g141(.A(new_new_n163_), .B(new_new_n160_), .Y(new_new_n164_));
  NO2        g142(.A(i_4_), .B(i_5_), .Y(new_new_n165_));
  NAi21      g143(.An(i_12_), .B(i_11_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n166_), .B(i_13_), .Y(new_new_n167_));
  NA3        g145(.A(new_new_n167_), .B(new_new_n165_), .C(new_new_n78_), .Y(new_new_n168_));
  AOI210     g146(.A0(new_new_n168_), .A1(new_new_n164_), .B0(new_new_n1011_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n69_), .B(new_new_n61_), .Y(new_new_n170_));
  NA2        g148(.A(new_new_n170_), .B(new_new_n45_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n36_), .B(i_5_), .Y(new_new_n172_));
  NAi31      g150(.An(new_new_n172_), .B(new_new_n142_), .C(i_11_), .Y(new_new_n173_));
  NA2        g151(.A(i_3_), .B(i_5_), .Y(new_new_n174_));
  OR2        g152(.A(new_new_n174_), .B(new_new_n163_), .Y(new_new_n175_));
  AOI210     g153(.A0(new_new_n175_), .A1(new_new_n173_), .B0(new_new_n171_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n69_), .B(i_5_), .Y(new_new_n177_));
  NO2        g155(.A(i_13_), .B(i_10_), .Y(new_new_n178_));
  NA3        g156(.A(new_new_n178_), .B(new_new_n177_), .C(new_new_n43_), .Y(new_new_n179_));
  NO2        g157(.A(i_2_), .B(i_1_), .Y(new_new_n180_));
  NA2        g158(.A(new_new_n180_), .B(i_3_), .Y(new_new_n181_));
  NAi21      g159(.An(i_4_), .B(i_12_), .Y(new_new_n182_));
  NO4        g160(.A(new_new_n182_), .B(new_new_n181_), .C(new_new_n179_), .D(new_new_n25_), .Y(new_new_n183_));
  NO3        g161(.A(new_new_n183_), .B(new_new_n176_), .C(new_new_n169_), .Y(new_new_n184_));
  INV        g162(.A(i_8_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(i_7_), .Y(new_new_n186_));
  NA2        g164(.A(new_new_n186_), .B(i_6_), .Y(new_new_n187_));
  NO3        g165(.A(i_3_), .B(new_new_n81_), .C(new_new_n47_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(new_new_n106_), .Y(new_new_n189_));
  NO3        g167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n190_));
  NA3        g168(.A(new_new_n190_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n191_));
  NO3        g169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n192_));
  NA2        g170(.A(i_12_), .B(new_new_n192_), .Y(new_new_n193_));
  AOI210     g171(.A0(new_new_n193_), .A1(new_new_n191_), .B0(new_new_n189_), .Y(new_new_n194_));
  NO2        g172(.A(i_3_), .B(i_8_), .Y(new_new_n195_));
  NO3        g173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n196_));
  NA3        g174(.A(new_new_n196_), .B(new_new_n195_), .C(new_new_n39_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n98_), .B(new_new_n57_), .Y(new_new_n198_));
  NO2        g176(.A(i_13_), .B(i_9_), .Y(new_new_n199_));
  NA3        g177(.A(new_new_n199_), .B(i_6_), .C(new_new_n185_), .Y(new_new_n200_));
  NAi21      g178(.An(i_12_), .B(i_3_), .Y(new_new_n201_));
  OR2        g179(.A(new_new_n201_), .B(new_new_n200_), .Y(new_new_n202_));
  NO2        g180(.A(new_new_n43_), .B(i_5_), .Y(new_new_n203_));
  NO3        g181(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n204_));
  OAI220     g182(.A0(i_2_), .A1(new_new_n202_), .B0(new_new_n98_), .B1(new_new_n197_), .Y(new_new_n205_));
  AOI210     g183(.A0(new_new_n205_), .A1(i_7_), .B0(new_new_n194_), .Y(new_new_n206_));
  OAI220     g184(.A0(new_new_n206_), .A1(i_4_), .B0(new_new_n187_), .B1(new_new_n184_), .Y(new_new_n207_));
  NAi21      g185(.An(i_12_), .B(i_7_), .Y(new_new_n208_));
  NA3        g186(.A(i_13_), .B(new_new_n185_), .C(i_10_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n210_));
  NA2        g188(.A(i_0_), .B(i_5_), .Y(new_new_n211_));
  NA2        g189(.A(new_new_n211_), .B(new_new_n99_), .Y(new_new_n212_));
  OAI220     g190(.A0(new_new_n212_), .A1(new_new_n181_), .B0(new_new_n171_), .B1(new_new_n126_), .Y(new_new_n213_));
  NAi31      g191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n36_), .B(i_13_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n69_), .B(new_new_n26_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n45_), .B(new_new_n61_), .Y(new_new_n217_));
  NA3        g195(.A(new_new_n217_), .B(new_new_n216_), .C(new_new_n215_), .Y(new_new_n218_));
  INV        g196(.A(i_13_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(new_new_n219_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n190_), .C(new_new_n188_), .Y(new_new_n221_));
  NA2        g199(.A(new_new_n218_), .B(new_new_n221_), .Y(new_new_n222_));
  AOI220     g200(.A0(new_new_n222_), .A1(new_new_n132_), .B0(new_new_n213_), .B1(new_new_n210_), .Y(new_new_n223_));
  NO2        g201(.A(i_12_), .B(new_new_n37_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n174_), .B(i_4_), .Y(new_new_n225_));
  INV        g203(.A(new_new_n225_), .Y(new_new_n226_));
  OR2        g204(.A(i_8_), .B(i_7_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n81_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n52_), .B(i_1_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n230_));
  INV        g208(.A(i_12_), .Y(new_new_n231_));
  NO3        g209(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n232_));
  NA2        g210(.A(i_2_), .B(i_1_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n230_), .B(new_new_n226_), .Y(new_new_n234_));
  NAi21      g212(.An(i_4_), .B(i_3_), .Y(new_new_n235_));
  NO2        g213(.A(new_new_n235_), .B(new_new_n71_), .Y(new_new_n236_));
  NO2        g214(.A(i_0_), .B(i_6_), .Y(new_new_n237_));
  NOi41      g215(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n238_), .B(new_new_n237_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n233_), .B(new_new_n174_), .Y(new_new_n240_));
  NAi21      g218(.An(new_new_n239_), .B(new_new_n240_), .Y(new_new_n241_));
  INV        g219(.A(new_new_n241_), .Y(new_new_n242_));
  AOI220     g220(.A0(new_new_n242_), .A1(new_new_n39_), .B0(new_new_n234_), .B1(new_new_n199_), .Y(new_new_n243_));
  NO2        g221(.A(i_11_), .B(new_new_n219_), .Y(new_new_n244_));
  NOi21      g222(.An(i_1_), .B(i_6_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n231_), .B(i_9_), .Y(new_new_n246_));
  OR4        g224(.A(new_new_n246_), .B(i_3_), .C(new_new_n245_), .D(new_new_n177_), .Y(new_new_n247_));
  NO2        g225(.A(new_new_n47_), .B(new_new_n25_), .Y(new_new_n248_));
  NO2        g226(.A(i_12_), .B(i_3_), .Y(new_new_n249_));
  NA2        g227(.A(new_new_n69_), .B(i_5_), .Y(new_new_n250_));
  NA2        g228(.A(i_3_), .B(i_9_), .Y(new_new_n251_));
  NAi21      g229(.An(i_7_), .B(i_10_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n252_), .B(new_new_n251_), .Y(new_new_n253_));
  NA3        g231(.A(new_new_n253_), .B(new_new_n250_), .C(new_new_n62_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n254_), .B(new_new_n247_), .Y(new_new_n255_));
  NA3        g233(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n255_), .B(new_new_n244_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n227_), .B(new_new_n37_), .Y(new_new_n258_));
  NA2        g236(.A(i_12_), .B(i_6_), .Y(new_new_n259_));
  OR2        g237(.A(i_13_), .B(i_9_), .Y(new_new_n260_));
  NO3        g238(.A(new_new_n260_), .B(new_new_n259_), .C(new_new_n47_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n235_), .B(i_2_), .Y(new_new_n262_));
  NA3        g240(.A(new_new_n262_), .B(new_new_n261_), .C(new_new_n43_), .Y(new_new_n263_));
  NA2        g241(.A(new_new_n244_), .B(i_9_), .Y(new_new_n264_));
  OAI210     g242(.A0(new_new_n69_), .A1(new_new_n264_), .B0(new_new_n263_), .Y(new_new_n265_));
  NA2        g243(.A(new_new_n145_), .B(new_new_n61_), .Y(new_new_n266_));
  NO3        g244(.A(i_11_), .B(new_new_n219_), .C(new_new_n25_), .Y(new_new_n267_));
  NO2        g245(.A(i_3_), .B(i_8_), .Y(new_new_n268_));
  NO2        g246(.A(i_6_), .B(new_new_n47_), .Y(new_new_n269_));
  NA3        g247(.A(new_new_n269_), .B(new_new_n268_), .C(new_new_n267_), .Y(new_new_n270_));
  NO3        g248(.A(new_new_n26_), .B(new_new_n81_), .C(i_5_), .Y(new_new_n271_));
  NA3        g249(.A(new_new_n271_), .B(new_new_n258_), .C(new_new_n220_), .Y(new_new_n272_));
  AOI210     g250(.A0(new_new_n272_), .A1(new_new_n270_), .B0(new_new_n266_), .Y(new_new_n273_));
  AOI210     g251(.A0(new_new_n265_), .A1(new_new_n258_), .B0(new_new_n273_), .Y(new_new_n274_));
  NA4        g252(.A(new_new_n274_), .B(new_new_n257_), .C(new_new_n243_), .D(new_new_n223_), .Y(new_new_n275_));
  NO3        g253(.A(i_12_), .B(new_new_n219_), .C(new_new_n37_), .Y(new_new_n276_));
  INV        g254(.A(new_new_n276_), .Y(new_new_n277_));
  NOi21      g255(.An(new_new_n154_), .B(new_new_n81_), .Y(new_new_n278_));
  NO3        g256(.A(i_0_), .B(new_new_n45_), .C(i_1_), .Y(new_new_n279_));
  AOI220     g257(.A0(new_new_n279_), .A1(new_new_n188_), .B0(new_new_n278_), .B1(new_new_n229_), .Y(new_new_n280_));
  NO2        g258(.A(new_new_n280_), .B(i_7_), .Y(new_new_n281_));
  NO3        g259(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n233_), .B(i_0_), .Y(new_new_n283_));
  AOI220     g261(.A0(new_new_n283_), .A1(new_new_n186_), .B0(new_new_n282_), .B1(new_new_n132_), .Y(new_new_n284_));
  NA2        g262(.A(new_new_n269_), .B(new_new_n26_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n285_), .B(new_new_n284_), .Y(new_new_n286_));
  NA2        g264(.A(i_0_), .B(i_1_), .Y(new_new_n287_));
  NO2        g265(.A(new_new_n287_), .B(i_2_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n58_), .B(i_6_), .Y(new_new_n289_));
  NA3        g267(.A(new_new_n289_), .B(new_new_n288_), .C(new_new_n154_), .Y(new_new_n290_));
  OAI210     g268(.A0(new_new_n156_), .A1(new_new_n133_), .B0(new_new_n290_), .Y(new_new_n291_));
  NO3        g269(.A(new_new_n291_), .B(new_new_n286_), .C(new_new_n281_), .Y(new_new_n292_));
  NO2        g270(.A(i_3_), .B(i_10_), .Y(new_new_n293_));
  NA3        g271(.A(new_new_n293_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n294_));
  NO2        g272(.A(i_2_), .B(new_new_n97_), .Y(new_new_n295_));
  NOi21      g273(.An(new_new_n211_), .B(new_new_n98_), .Y(new_new_n296_));
  NA3        g274(.A(new_new_n296_), .B(i_1_), .C(new_new_n295_), .Y(new_new_n297_));
  AN2        g275(.A(i_3_), .B(i_10_), .Y(new_new_n298_));
  NA3        g276(.A(new_new_n190_), .B(new_new_n167_), .C(new_new_n165_), .Y(new_new_n299_));
  NO2        g277(.A(i_5_), .B(new_new_n37_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n45_), .B(new_new_n26_), .Y(new_new_n301_));
  OR2        g279(.A(new_new_n297_), .B(new_new_n294_), .Y(new_new_n302_));
  OAI220     g280(.A0(new_new_n302_), .A1(i_6_), .B0(new_new_n292_), .B1(new_new_n277_), .Y(new_new_n303_));
  NO4        g281(.A(new_new_n303_), .B(new_new_n275_), .C(new_new_n207_), .D(new_new_n159_), .Y(new_new_n304_));
  NO3        g282(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n305_));
  NO3        g283(.A(i_6_), .B(new_new_n185_), .C(i_7_), .Y(new_new_n306_));
  NA2        g284(.A(new_new_n306_), .B(new_new_n190_), .Y(new_new_n307_));
  AOI210     g285(.A0(new_new_n307_), .A1(new_new_n233_), .B0(new_new_n160_), .Y(new_new_n308_));
  NO2        g286(.A(i_2_), .B(i_3_), .Y(new_new_n309_));
  OR2        g287(.A(i_0_), .B(i_5_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n211_), .B(new_new_n310_), .Y(new_new_n311_));
  NA4        g289(.A(new_new_n311_), .B(new_new_n228_), .C(new_new_n309_), .D(i_1_), .Y(new_new_n312_));
  NA3        g290(.A(new_new_n283_), .B(new_new_n278_), .C(new_new_n106_), .Y(new_new_n313_));
  NO2        g291(.A(i_8_), .B(i_6_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n148_), .B(new_new_n45_), .Y(new_new_n315_));
  NA3        g293(.A(new_new_n315_), .B(new_new_n314_), .C(new_new_n154_), .Y(new_new_n316_));
  NA3        g294(.A(new_new_n316_), .B(new_new_n313_), .C(new_new_n312_), .Y(new_new_n317_));
  OAI210     g295(.A0(new_new_n317_), .A1(new_new_n308_), .B0(i_4_), .Y(new_new_n318_));
  NO2        g296(.A(i_12_), .B(i_10_), .Y(new_new_n319_));
  NOi21      g297(.An(i_5_), .B(i_0_), .Y(new_new_n320_));
  AOI210     g298(.A0(i_2_), .A1(new_new_n47_), .B0(new_new_n97_), .Y(new_new_n321_));
  NO4        g299(.A(new_new_n321_), .B(i_4_), .C(new_new_n320_), .D(new_new_n121_), .Y(new_new_n322_));
  NA4        g300(.A(new_new_n79_), .B(new_new_n36_), .C(new_new_n81_), .D(i_8_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n322_), .B(new_new_n319_), .Y(new_new_n324_));
  NO2        g302(.A(i_6_), .B(i_8_), .Y(new_new_n325_));
  AN2        g303(.A(i_0_), .B(new_new_n325_), .Y(new_new_n326_));
  NO2        g304(.A(i_1_), .B(i_7_), .Y(new_new_n327_));
  NA3        g305(.A(new_new_n326_), .B(i_4_), .C(i_5_), .Y(new_new_n328_));
  NA3        g306(.A(new_new_n328_), .B(new_new_n324_), .C(new_new_n318_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n1016_), .B(i_6_), .Y(new_new_n330_));
  NA3        g308(.A(new_new_n245_), .B(new_new_n295_), .C(new_new_n185_), .Y(new_new_n331_));
  AOI210     g309(.A0(new_new_n331_), .A1(new_new_n330_), .B0(new_new_n311_), .Y(new_new_n332_));
  NOi21      g310(.An(new_new_n144_), .B(new_new_n99_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n333_), .B(new_new_n117_), .Y(new_new_n334_));
  OAI210     g312(.A0(new_new_n334_), .A1(new_new_n332_), .B0(i_3_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n287_), .B(new_new_n77_), .Y(new_new_n336_));
  NA2        g314(.A(new_new_n336_), .B(new_new_n125_), .Y(new_new_n337_));
  NO2        g315(.A(new_new_n88_), .B(new_new_n185_), .Y(new_new_n338_));
  NA3        g316(.A(new_new_n296_), .B(new_new_n338_), .C(new_new_n61_), .Y(new_new_n339_));
  AOI210     g317(.A0(new_new_n339_), .A1(new_new_n337_), .B0(i_3_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n185_), .B(i_9_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n198_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n340_), .B(new_new_n286_), .Y(new_new_n343_));
  AOI210     g321(.A0(new_new_n343_), .A1(new_new_n335_), .B0(new_new_n153_), .Y(new_new_n344_));
  AOI210     g322(.A0(new_new_n329_), .A1(new_new_n305_), .B0(new_new_n344_), .Y(new_new_n345_));
  NOi32      g323(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n346_));
  INV        g324(.A(new_new_n346_), .Y(new_new_n347_));
  NAi21      g325(.An(i_1_), .B(i_5_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n348_), .B(i_0_), .Y(new_new_n349_));
  NA2        g327(.A(new_new_n349_), .B(new_new_n25_), .Y(new_new_n350_));
  OAI210     g328(.A0(new_new_n350_), .A1(new_new_n150_), .B0(new_new_n239_), .Y(new_new_n351_));
  NAi41      g329(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n352_));
  OAI220     g330(.A0(new_new_n352_), .A1(new_new_n348_), .B0(new_new_n214_), .B1(new_new_n150_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n150_), .B(new_new_n148_), .Y(new_new_n354_));
  NOi32      g332(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n355_));
  NAi21      g333(.An(i_6_), .B(i_1_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n355_), .B(new_new_n45_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n357_), .B(i_0_), .Y(new_new_n358_));
  OR3        g336(.A(new_new_n358_), .B(new_new_n354_), .C(new_new_n353_), .Y(new_new_n359_));
  NO2        g337(.A(i_1_), .B(new_new_n97_), .Y(new_new_n360_));
  NAi21      g338(.An(i_3_), .B(i_4_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n361_), .B(i_9_), .Y(new_new_n362_));
  AN2        g340(.A(i_6_), .B(i_7_), .Y(new_new_n363_));
  OAI210     g341(.A0(new_new_n363_), .A1(new_new_n360_), .B0(new_new_n362_), .Y(new_new_n364_));
  NA2        g342(.A(i_2_), .B(i_7_), .Y(new_new_n365_));
  NO2        g343(.A(new_new_n361_), .B(i_10_), .Y(new_new_n366_));
  NA3        g344(.A(new_new_n366_), .B(new_new_n365_), .C(new_new_n237_), .Y(new_new_n367_));
  AOI210     g345(.A0(new_new_n367_), .A1(new_new_n364_), .B0(new_new_n177_), .Y(new_new_n368_));
  AOI210     g346(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n369_));
  OAI210     g347(.A0(new_new_n369_), .A1(new_new_n180_), .B0(new_new_n366_), .Y(new_new_n370_));
  AOI220     g348(.A0(new_new_n366_), .A1(new_new_n327_), .B0(new_new_n232_), .B1(new_new_n180_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n370_), .B(i_5_), .Y(new_new_n372_));
  NO4        g350(.A(new_new_n372_), .B(new_new_n368_), .C(new_new_n359_), .D(new_new_n351_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n373_), .B(new_new_n347_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n58_), .B(new_new_n25_), .Y(new_new_n375_));
  AN2        g353(.A(i_12_), .B(i_5_), .Y(new_new_n376_));
  NO2        g354(.A(i_4_), .B(new_new_n26_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n377_), .B(new_new_n376_), .Y(new_new_n378_));
  NO2        g356(.A(i_11_), .B(i_6_), .Y(new_new_n379_));
  NA3        g357(.A(new_new_n379_), .B(new_new_n315_), .C(new_new_n219_), .Y(new_new_n380_));
  NO2        g358(.A(new_new_n380_), .B(new_new_n378_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n235_), .B(i_5_), .Y(new_new_n382_));
  NO2        g360(.A(i_5_), .B(i_10_), .Y(new_new_n383_));
  AOI220     g361(.A0(new_new_n383_), .A1(new_new_n262_), .B0(new_new_n382_), .B1(new_new_n190_), .Y(new_new_n384_));
  INV        g362(.A(new_new_n44_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n385_), .B(new_new_n384_), .Y(new_new_n386_));
  OAI210     g364(.A0(new_new_n386_), .A1(new_new_n381_), .B0(new_new_n375_), .Y(new_new_n387_));
  NO2        g365(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n140_), .B(new_new_n81_), .Y(new_new_n389_));
  OAI210     g367(.A0(new_new_n389_), .A1(new_new_n381_), .B0(new_new_n388_), .Y(new_new_n390_));
  NO3        g368(.A(new_new_n81_), .B(new_new_n47_), .C(i_9_), .Y(new_new_n391_));
  NO2        g369(.A(i_11_), .B(i_12_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n392_), .B(new_new_n36_), .Y(new_new_n393_));
  NO2        g371(.A(i_3_), .B(new_new_n393_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n383_), .B(new_new_n231_), .Y(new_new_n395_));
  NA3        g373(.A(new_new_n106_), .B(i_4_), .C(i_11_), .Y(new_new_n396_));
  INV        g374(.A(new_new_n396_), .Y(new_new_n397_));
  NAi21      g375(.An(i_13_), .B(i_0_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n233_), .Y(new_new_n399_));
  OAI210     g377(.A0(new_new_n397_), .A1(new_new_n394_), .B0(new_new_n399_), .Y(new_new_n400_));
  NA3        g378(.A(new_new_n400_), .B(new_new_n390_), .C(new_new_n387_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n43_), .B(new_new_n219_), .Y(new_new_n402_));
  NO3        g380(.A(i_1_), .B(i_12_), .C(new_new_n81_), .Y(new_new_n403_));
  NO2        g381(.A(i_0_), .B(i_11_), .Y(new_new_n404_));
  AN2        g382(.A(i_1_), .B(i_6_), .Y(new_new_n405_));
  NOi21      g383(.An(i_2_), .B(i_12_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n406_), .B(new_new_n405_), .Y(new_new_n407_));
  NO2        g385(.A(new_new_n407_), .B(new_new_n1010_), .Y(new_new_n408_));
  NA2        g386(.A(new_new_n132_), .B(i_9_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n408_), .B(i_9_), .Y(new_new_n410_));
  NAi21      g388(.An(i_9_), .B(i_4_), .Y(new_new_n411_));
  OR2        g389(.A(i_13_), .B(i_10_), .Y(new_new_n412_));
  NO3        g390(.A(new_new_n412_), .B(new_new_n110_), .C(new_new_n411_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n163_), .B(new_new_n116_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n97_), .B(new_new_n25_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n276_), .B(new_new_n415_), .Y(new_new_n416_));
  NA2        g394(.A(new_new_n269_), .B(new_new_n204_), .Y(new_new_n417_));
  OAI220     g395(.A0(new_new_n417_), .A1(new_new_n209_), .B0(new_new_n416_), .B1(new_new_n333_), .Y(new_new_n418_));
  INV        g396(.A(new_new_n418_), .Y(new_new_n419_));
  AOI210     g397(.A0(new_new_n419_), .A1(new_new_n410_), .B0(new_new_n26_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n313_), .B(new_new_n312_), .Y(new_new_n421_));
  AOI220     g399(.A0(new_new_n289_), .A1(new_new_n279_), .B0(new_new_n283_), .B1(i_7_), .Y(new_new_n422_));
  NO2        g400(.A(new_new_n174_), .B(new_new_n81_), .Y(new_new_n423_));
  AOI220     g401(.A0(new_new_n423_), .A1(new_new_n288_), .B0(new_new_n271_), .B1(new_new_n204_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n424_), .B(i_7_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n425_), .B(new_new_n421_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n188_), .B(new_new_n92_), .Y(new_new_n427_));
  NA3        g405(.A(new_new_n315_), .B(new_new_n154_), .C(new_new_n81_), .Y(new_new_n428_));
  AOI210     g406(.A0(new_new_n428_), .A1(new_new_n427_), .B0(i_8_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n185_), .B(i_10_), .Y(new_new_n430_));
  NA3        g408(.A(new_new_n250_), .B(new_new_n62_), .C(i_2_), .Y(new_new_n431_));
  NA2        g409(.A(new_new_n289_), .B(new_new_n229_), .Y(new_new_n432_));
  OAI220     g410(.A0(new_new_n432_), .A1(new_new_n174_), .B0(new_new_n431_), .B1(new_new_n430_), .Y(new_new_n433_));
  NO2        g411(.A(i_3_), .B(new_new_n47_), .Y(new_new_n434_));
  NA3        g412(.A(new_new_n327_), .B(new_new_n326_), .C(new_new_n434_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n306_), .B(new_new_n311_), .Y(new_new_n436_));
  OAI210     g414(.A0(new_new_n436_), .A1(new_new_n181_), .B0(new_new_n435_), .Y(new_new_n437_));
  NO3        g415(.A(new_new_n437_), .B(new_new_n433_), .C(new_new_n429_), .Y(new_new_n438_));
  AOI210     g416(.A0(new_new_n438_), .A1(new_new_n426_), .B0(new_new_n264_), .Y(new_new_n439_));
  NO4        g417(.A(new_new_n439_), .B(new_new_n420_), .C(new_new_n401_), .D(new_new_n374_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n69_), .B(i_13_), .Y(new_new_n441_));
  NO2        g419(.A(i_10_), .B(i_9_), .Y(new_new_n442_));
  NAi21      g420(.An(i_12_), .B(i_8_), .Y(new_new_n443_));
  NO2        g421(.A(new_new_n443_), .B(i_3_), .Y(new_new_n444_));
  NA2        g422(.A(i_2_), .B(new_new_n99_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n445_), .B(new_new_n197_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n301_), .B(i_0_), .Y(new_new_n447_));
  NO3        g425(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n448_));
  NA2        g426(.A(new_new_n259_), .B(new_new_n93_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n449_), .B(new_new_n448_), .Y(new_new_n450_));
  NA2        g428(.A(i_8_), .B(i_9_), .Y(new_new_n451_));
  NA2        g429(.A(new_new_n276_), .B(new_new_n198_), .Y(new_new_n452_));
  OAI220     g430(.A0(new_new_n452_), .A1(new_new_n451_), .B0(new_new_n450_), .B1(new_new_n447_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n244_), .B(new_new_n300_), .Y(new_new_n454_));
  NO3        g432(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n455_));
  INV        g433(.A(new_new_n455_), .Y(new_new_n456_));
  NA3        g434(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n456_), .B(new_new_n454_), .Y(new_new_n458_));
  NO3        g436(.A(new_new_n458_), .B(new_new_n453_), .C(new_new_n446_), .Y(new_new_n459_));
  NA2        g437(.A(new_new_n288_), .B(new_new_n101_), .Y(new_new_n460_));
  OR2        g438(.A(new_new_n460_), .B(new_new_n200_), .Y(new_new_n461_));
  OA220      g439(.A0(new_new_n342_), .A1(new_new_n153_), .B0(new_new_n461_), .B1(new_new_n226_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n92_), .B(i_13_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n423_), .B(new_new_n375_), .Y(new_new_n464_));
  NO2        g442(.A(i_2_), .B(i_13_), .Y(new_new_n465_));
  NA3        g443(.A(new_new_n465_), .B(new_new_n152_), .C(new_new_n95_), .Y(new_new_n466_));
  OAI220     g444(.A0(new_new_n466_), .A1(new_new_n231_), .B0(new_new_n464_), .B1(new_new_n463_), .Y(new_new_n467_));
  NO3        g445(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n468_));
  NO2        g446(.A(i_6_), .B(i_7_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n69_), .B(i_3_), .Y(new_new_n470_));
  NOi21      g448(.An(i_2_), .B(i_7_), .Y(new_new_n471_));
  NAi31      g449(.An(i_11_), .B(new_new_n471_), .C(new_new_n470_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n412_), .B(i_6_), .Y(new_new_n473_));
  NA3        g451(.A(new_new_n473_), .B(i_1_), .C(new_new_n71_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n474_), .B(new_new_n472_), .Y(new_new_n475_));
  NO2        g453(.A(i_3_), .B(new_new_n185_), .Y(new_new_n476_));
  NO2        g454(.A(i_6_), .B(i_10_), .Y(new_new_n477_));
  NA4        g455(.A(new_new_n477_), .B(new_new_n305_), .C(new_new_n476_), .D(new_new_n231_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n478_), .B(new_new_n146_), .Y(new_new_n479_));
  NA3        g457(.A(new_new_n238_), .B(new_new_n162_), .C(new_new_n125_), .Y(new_new_n480_));
  NA2        g458(.A(new_new_n45_), .B(new_new_n43_), .Y(new_new_n481_));
  NO2        g459(.A(new_new_n148_), .B(i_3_), .Y(new_new_n482_));
  NAi31      g460(.An(new_new_n481_), .B(new_new_n482_), .C(new_new_n220_), .Y(new_new_n483_));
  NA3        g461(.A(new_new_n388_), .B(new_new_n170_), .C(new_new_n139_), .Y(new_new_n484_));
  NA3        g462(.A(new_new_n484_), .B(new_new_n483_), .C(new_new_n480_), .Y(new_new_n485_));
  NO4        g463(.A(new_new_n485_), .B(new_new_n479_), .C(new_new_n475_), .D(new_new_n467_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n448_), .B(new_new_n376_), .Y(new_new_n487_));
  NA2        g465(.A(new_new_n455_), .B(new_new_n383_), .Y(new_new_n488_));
  NO2        g466(.A(new_new_n488_), .B(new_new_n218_), .Y(new_new_n489_));
  NAi21      g467(.An(new_new_n209_), .B(new_new_n392_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n327_), .B(new_new_n211_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n26_), .B(i_5_), .Y(new_new_n492_));
  NA3        g470(.A(new_new_n1019_), .B(new_new_n492_), .C(new_new_n132_), .Y(new_new_n493_));
  OAI220     g471(.A0(new_new_n38_), .A1(new_new_n493_), .B0(new_new_n491_), .B1(new_new_n490_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n27_), .B(i_10_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n495_), .B(new_new_n463_), .Y(new_new_n496_));
  NO3        g474(.A(new_new_n496_), .B(new_new_n494_), .C(new_new_n489_), .Y(new_new_n497_));
  NA4        g475(.A(new_new_n497_), .B(new_new_n486_), .C(new_new_n462_), .D(new_new_n459_), .Y(new_new_n498_));
  NA2        g476(.A(new_new_n167_), .B(new_new_n165_), .Y(new_new_n499_));
  OAI210     g477(.A0(new_new_n294_), .A1(new_new_n172_), .B0(new_new_n499_), .Y(new_new_n500_));
  AN2        g478(.A(new_new_n279_), .B(new_new_n228_), .Y(new_new_n501_));
  NA2        g479(.A(new_new_n501_), .B(new_new_n500_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n115_), .B(new_new_n105_), .Y(new_new_n503_));
  AO220      g481(.A0(new_new_n503_), .A1(new_new_n448_), .B0(new_new_n413_), .B1(i_6_), .Y(new_new_n504_));
  NA2        g482(.A(new_new_n305_), .B(new_new_n155_), .Y(new_new_n505_));
  OAI210     g483(.A0(new_new_n505_), .A1(new_new_n226_), .B0(new_new_n299_), .Y(new_new_n506_));
  AOI220     g484(.A0(new_new_n506_), .A1(new_new_n314_), .B0(new_new_n504_), .B1(new_new_n301_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n376_), .B(new_new_n219_), .Y(new_new_n508_));
  NA2        g486(.A(new_new_n346_), .B(new_new_n69_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n363_), .B(new_new_n355_), .Y(new_new_n510_));
  AO210      g488(.A0(new_new_n509_), .A1(new_new_n508_), .B0(new_new_n510_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n36_), .B(i_8_), .Y(new_new_n512_));
  INV        g490(.A(new_new_n413_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n513_), .B(new_new_n511_), .Y(new_new_n514_));
  INV        g492(.A(new_new_n514_), .Y(new_new_n515_));
  OAI210     g493(.A0(i_8_), .A1(new_new_n61_), .B0(new_new_n127_), .Y(new_new_n516_));
  AOI210     g494(.A0(new_new_n186_), .A1(i_9_), .B0(new_new_n258_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n517_), .B(new_new_n191_), .Y(new_new_n518_));
  AOI220     g496(.A0(i_5_), .A1(new_new_n518_), .B0(new_new_n516_), .B1(new_new_n414_), .Y(new_new_n519_));
  NA4        g497(.A(new_new_n519_), .B(new_new_n515_), .C(new_new_n507_), .D(new_new_n502_), .Y(new_new_n520_));
  NO2        g498(.A(i_12_), .B(new_new_n185_), .Y(new_new_n521_));
  NA3        g499(.A(new_new_n477_), .B(new_new_n165_), .C(new_new_n27_), .Y(new_new_n522_));
  NO3        g500(.A(new_new_n522_), .B(i_13_), .C(new_new_n460_), .Y(new_new_n523_));
  NOi31      g501(.An(new_new_n306_), .B(new_new_n412_), .C(new_new_n38_), .Y(new_new_n524_));
  OAI210     g502(.A0(new_new_n524_), .A1(new_new_n523_), .B0(new_new_n377_), .Y(new_new_n525_));
  NO2        g503(.A(i_8_), .B(i_7_), .Y(new_new_n526_));
  AOI220     g504(.A0(new_new_n315_), .A1(new_new_n39_), .B0(new_new_n229_), .B1(new_new_n199_), .Y(new_new_n527_));
  OAI220     g505(.A0(new_new_n527_), .A1(new_new_n174_), .B0(i_5_), .B1(new_new_n235_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n43_), .B(i_10_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n529_), .B(i_6_), .Y(new_new_n530_));
  NA3        g508(.A(new_new_n530_), .B(new_new_n528_), .C(new_new_n526_), .Y(new_new_n531_));
  AOI220     g509(.A0(new_new_n423_), .A1(new_new_n315_), .B0(new_new_n240_), .B1(new_new_n237_), .Y(new_new_n532_));
  OAI220     g510(.A0(new_new_n532_), .A1(i_12_), .B0(new_new_n463_), .B1(new_new_n126_), .Y(new_new_n533_));
  NA2        g511(.A(new_new_n533_), .B(new_new_n258_), .Y(new_new_n534_));
  NOi31      g512(.An(new_new_n283_), .B(new_new_n294_), .C(new_new_n172_), .Y(new_new_n535_));
  NA3        g513(.A(new_new_n298_), .B(new_new_n165_), .C(new_new_n92_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n148_), .B(i_5_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n537_), .B(new_new_n402_), .C(new_new_n309_), .Y(new_new_n538_));
  NA2        g516(.A(new_new_n538_), .B(new_new_n536_), .Y(new_new_n539_));
  OAI210     g517(.A0(new_new_n539_), .A1(new_new_n535_), .B0(new_new_n455_), .Y(new_new_n540_));
  NA4        g518(.A(new_new_n540_), .B(new_new_n534_), .C(new_new_n531_), .D(new_new_n525_), .Y(new_new_n541_));
  NA3        g519(.A(new_new_n211_), .B(new_new_n67_), .C(new_new_n43_), .Y(new_new_n542_));
  NA2        g520(.A(new_new_n276_), .B(new_new_n79_), .Y(new_new_n543_));
  AOI210     g521(.A0(new_new_n542_), .A1(new_new_n337_), .B0(new_new_n543_), .Y(new_new_n544_));
  NA2        g522(.A(new_new_n289_), .B(new_new_n279_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n545_), .B(new_new_n164_), .Y(new_new_n546_));
  NA2        g524(.A(new_new_n217_), .B(new_new_n216_), .Y(new_new_n547_));
  NA2        g525(.A(new_new_n442_), .B(new_new_n215_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n547_), .B(new_new_n548_), .Y(new_new_n549_));
  NA2        g527(.A(i_0_), .B(new_new_n47_), .Y(new_new_n550_));
  NA3        g528(.A(new_new_n521_), .B(new_new_n267_), .C(new_new_n550_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n1017_), .B(new_new_n551_), .Y(new_new_n552_));
  NO4        g530(.A(new_new_n552_), .B(new_new_n549_), .C(new_new_n546_), .D(new_new_n544_), .Y(new_new_n553_));
  NO4        g531(.A(new_new_n245_), .B(new_new_n41_), .C(i_2_), .D(new_new_n47_), .Y(new_new_n554_));
  NO3        g532(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n227_), .B(new_new_n36_), .Y(new_new_n556_));
  AN2        g534(.A(new_new_n556_), .B(new_new_n555_), .Y(new_new_n557_));
  OA210      g535(.A0(new_new_n557_), .A1(new_new_n554_), .B0(new_new_n346_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n412_), .B(i_1_), .Y(new_new_n559_));
  NOi31      g537(.An(new_new_n559_), .B(new_new_n449_), .C(new_new_n69_), .Y(new_new_n560_));
  AN4        g538(.A(new_new_n560_), .B(i_9_), .C(new_new_n492_), .D(i_2_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n422_), .B(new_new_n168_), .Y(new_new_n562_));
  NO3        g540(.A(new_new_n562_), .B(new_new_n561_), .C(new_new_n558_), .Y(new_new_n563_));
  NOi21      g541(.An(i_10_), .B(i_6_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n81_), .B(new_new_n25_), .Y(new_new_n565_));
  AOI220     g543(.A0(new_new_n276_), .A1(new_new_n565_), .B0(new_new_n267_), .B1(new_new_n564_), .Y(new_new_n566_));
  NO2        g544(.A(new_new_n566_), .B(new_new_n447_), .Y(new_new_n567_));
  NO2        g545(.A(new_new_n108_), .B(new_new_n23_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n306_), .B(new_new_n155_), .Y(new_new_n569_));
  AOI220     g547(.A0(new_new_n569_), .A1(new_new_n432_), .B0(new_new_n175_), .B1(new_new_n173_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n190_), .B(new_new_n37_), .Y(new_new_n571_));
  NOi31      g549(.An(new_new_n136_), .B(new_new_n571_), .C(new_new_n323_), .Y(new_new_n572_));
  NO3        g550(.A(new_new_n572_), .B(new_new_n570_), .C(new_new_n567_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n509_), .B(new_new_n371_), .Y(new_new_n574_));
  INV        g552(.A(new_new_n309_), .Y(new_new_n575_));
  NO2        g553(.A(i_12_), .B(new_new_n81_), .Y(new_new_n576_));
  NA3        g554(.A(new_new_n379_), .B(new_new_n276_), .C(new_new_n211_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n577_), .B(new_new_n575_), .Y(new_new_n578_));
  NA2        g556(.A(new_new_n165_), .B(i_0_), .Y(new_new_n579_));
  NO3        g557(.A(new_new_n579_), .B(new_new_n330_), .C(new_new_n294_), .Y(new_new_n580_));
  OR2        g558(.A(i_2_), .B(i_5_), .Y(new_new_n581_));
  OR2        g559(.A(new_new_n581_), .B(new_new_n405_), .Y(new_new_n582_));
  INV        g560(.A(new_new_n190_), .Y(new_new_n583_));
  AOI210     g561(.A0(new_new_n583_), .A1(new_new_n582_), .B0(new_new_n490_), .Y(new_new_n584_));
  NO4        g562(.A(new_new_n584_), .B(new_new_n580_), .C(new_new_n578_), .D(new_new_n574_), .Y(new_new_n585_));
  NA4        g563(.A(new_new_n585_), .B(new_new_n573_), .C(new_new_n563_), .D(new_new_n553_), .Y(new_new_n586_));
  NO4        g564(.A(new_new_n586_), .B(new_new_n541_), .C(new_new_n520_), .D(new_new_n498_), .Y(new_new_n587_));
  NA4        g565(.A(new_new_n587_), .B(new_new_n440_), .C(new_new_n345_), .D(new_new_n304_), .Y(men7));
  NO2        g566(.A(new_new_n101_), .B(new_new_n86_), .Y(new_new_n589_));
  NA2        g567(.A(new_new_n477_), .B(new_new_n79_), .Y(new_new_n590_));
  NA2        g568(.A(i_11_), .B(new_new_n185_), .Y(new_new_n591_));
  NA3        g569(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n592_));
  NA2        g570(.A(i_12_), .B(i_8_), .Y(new_new_n593_));
  AOI210     g571(.A0(new_new_n593_), .A1(new_new_n100_), .B0(new_new_n592_), .Y(new_new_n594_));
  NA2        g572(.A(i_2_), .B(new_new_n81_), .Y(new_new_n595_));
  OAI210     g573(.A0(new_new_n84_), .A1(new_new_n195_), .B0(new_new_n196_), .Y(new_new_n596_));
  NO2        g574(.A(i_7_), .B(new_new_n37_), .Y(new_new_n597_));
  NA2        g575(.A(i_4_), .B(i_8_), .Y(new_new_n598_));
  NO2        g576(.A(new_new_n594_), .B(new_new_n589_), .Y(new_new_n599_));
  OR2        g577(.A(i_6_), .B(i_10_), .Y(new_new_n600_));
  NO2        g578(.A(new_new_n600_), .B(new_new_n23_), .Y(new_new_n601_));
  NO3        g579(.A(i_6_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n602_));
  INV        g580(.A(new_new_n192_), .Y(new_new_n603_));
  NO2        g581(.A(new_new_n599_), .B(new_new_n61_), .Y(new_new_n604_));
  NOi21      g582(.An(i_11_), .B(i_7_), .Y(new_new_n605_));
  AO210      g583(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n606_));
  NO2        g584(.A(new_new_n606_), .B(new_new_n605_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n607_), .B(new_new_n199_), .Y(new_new_n608_));
  NA3        g586(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n609_));
  NAi31      g587(.An(new_new_n609_), .B(new_new_n208_), .C(i_11_), .Y(new_new_n610_));
  AOI210     g588(.A0(new_new_n610_), .A1(new_new_n608_), .B0(new_new_n61_), .Y(new_new_n611_));
  NO3        g589(.A(new_new_n252_), .B(new_new_n201_), .C(new_new_n591_), .Y(new_new_n612_));
  OAI210     g590(.A0(new_new_n612_), .A1(new_new_n220_), .B0(new_new_n61_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n406_), .B(new_new_n31_), .Y(new_new_n614_));
  OR2        g592(.A(new_new_n201_), .B(new_new_n101_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n615_), .B(new_new_n614_), .Y(new_new_n616_));
  NO2        g594(.A(new_new_n61_), .B(i_9_), .Y(new_new_n617_));
  INV        g595(.A(i_4_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n618_), .B(new_new_n616_), .Y(new_new_n619_));
  NO2        g597(.A(i_1_), .B(i_12_), .Y(new_new_n620_));
  NA3        g598(.A(new_new_n620_), .B(new_new_n103_), .C(new_new_n24_), .Y(new_new_n621_));
  NA4        g599(.A(new_new_n621_), .B(new_new_n619_), .C(new_new_n613_), .D(new_new_n82_), .Y(new_new_n622_));
  OAI210     g600(.A0(new_new_n622_), .A1(new_new_n611_), .B0(i_6_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n609_), .B(new_new_n101_), .Y(new_new_n624_));
  NA2        g602(.A(new_new_n624_), .B(new_new_n576_), .Y(new_new_n625_));
  NO2        g603(.A(i_6_), .B(i_11_), .Y(new_new_n626_));
  NA2        g604(.A(new_new_n625_), .B(new_new_n450_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n1022_), .B(new_new_n617_), .Y(new_new_n628_));
  NO3        g606(.A(new_new_n600_), .B(new_new_n227_), .C(new_new_n23_), .Y(new_new_n629_));
  AOI210     g607(.A0(i_1_), .A1(new_new_n253_), .B0(new_new_n629_), .Y(new_new_n630_));
  OAI210     g608(.A0(new_new_n630_), .A1(new_new_n43_), .B0(new_new_n628_), .Y(new_new_n631_));
  NA3        g609(.A(new_new_n526_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n632_));
  NA3        g610(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n633_));
  NO2        g611(.A(new_new_n45_), .B(i_1_), .Y(new_new_n634_));
  NA3        g612(.A(new_new_n634_), .B(new_new_n259_), .C(new_new_n43_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n635_), .B(new_new_n633_), .Y(new_new_n636_));
  NO2        g614(.A(i_11_), .B(new_new_n37_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n637_), .B(new_new_n24_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(i_6_), .Y(new_new_n639_));
  OR2        g617(.A(new_new_n639_), .B(new_new_n636_), .Y(new_new_n640_));
  NO3        g618(.A(new_new_n640_), .B(new_new_n631_), .C(new_new_n627_), .Y(new_new_n641_));
  INV        g619(.A(new_new_n605_), .Y(new_new_n642_));
  NA2        g620(.A(new_new_n642_), .B(i_1_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n643_), .B(i_6_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n411_), .B(new_new_n81_), .Y(new_new_n645_));
  NA2        g623(.A(new_new_n644_), .B(new_new_n45_), .Y(new_new_n646_));
  NA2        g624(.A(i_3_), .B(new_new_n185_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n227_), .B(new_new_n43_), .Y(new_new_n648_));
  NO3        g626(.A(new_new_n648_), .B(new_new_n301_), .C(i_12_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n110_), .B(new_new_n37_), .Y(new_new_n650_));
  INV        g628(.A(i_6_), .Y(new_new_n651_));
  NO2        g629(.A(new_new_n81_), .B(i_9_), .Y(new_new_n652_));
  NO2        g630(.A(new_new_n652_), .B(new_new_n61_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n653_), .B(new_new_n620_), .Y(new_new_n654_));
  NO4        g632(.A(new_new_n654_), .B(new_new_n651_), .C(new_new_n649_), .D(i_4_), .Y(new_new_n655_));
  NA2        g633(.A(i_1_), .B(i_3_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n451_), .B(new_new_n88_), .Y(new_new_n657_));
  INV        g635(.A(new_new_n657_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n658_), .B(new_new_n656_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n659_), .B(new_new_n655_), .Y(new_new_n660_));
  NA4        g638(.A(new_new_n660_), .B(new_new_n646_), .C(new_new_n641_), .D(new_new_n623_), .Y(new_new_n661_));
  NO3        g639(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n662_));
  OA210      g640(.A0(new_new_n662_), .A1(new_new_n238_), .B0(new_new_n81_), .Y(new_new_n663_));
  NA2        g641(.A(new_new_n363_), .B(new_new_n362_), .Y(new_new_n664_));
  NO2        g642(.A(new_new_n598_), .B(new_new_n81_), .Y(new_new_n665_));
  NA2        g643(.A(new_new_n665_), .B(new_new_n25_), .Y(new_new_n666_));
  INV        g644(.A(new_new_n666_), .Y(new_new_n667_));
  OAI210     g645(.A0(new_new_n667_), .A1(new_new_n663_), .B0(i_1_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n259_), .B(new_new_n93_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n361_), .B(i_2_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n670_), .B(new_new_n669_), .Y(new_new_n671_));
  AOI210     g649(.A0(new_new_n671_), .A1(new_new_n668_), .B0(i_13_), .Y(new_new_n672_));
  OR2        g650(.A(i_11_), .B(i_7_), .Y(new_new_n673_));
  AOI220     g651(.A0(new_new_n465_), .A1(new_new_n152_), .B0(i_2_), .B1(i_1_), .Y(new_new_n674_));
  NO2        g652(.A(new_new_n674_), .B(new_new_n43_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n471_), .B(new_new_n24_), .Y(new_new_n676_));
  AOI210     g654(.A0(new_new_n676_), .A1(new_new_n645_), .B0(new_new_n238_), .Y(new_new_n677_));
  OAI220     g655(.A0(new_new_n677_), .A1(new_new_n40_), .B0(new_new_n53_), .B1(new_new_n88_), .Y(new_new_n678_));
  AOI210     g656(.A0(new_new_n675_), .A1(new_new_n325_), .B0(new_new_n678_), .Y(new_new_n679_));
  AOI220     g657(.A0(i_12_), .A1(new_new_n68_), .B0(new_new_n379_), .B1(new_new_n634_), .Y(new_new_n680_));
  NO2        g658(.A(new_new_n680_), .B(new_new_n235_), .Y(new_new_n681_));
  AOI210     g659(.A0(new_new_n443_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n682_));
  NO2        g660(.A(new_new_n590_), .B(new_new_n43_), .Y(new_new_n683_));
  NO2        g661(.A(new_new_n633_), .B(new_new_n108_), .Y(new_new_n684_));
  NO3        g662(.A(new_new_n67_), .B(new_new_n32_), .C(new_new_n97_), .Y(new_new_n685_));
  NA2        g663(.A(i_3_), .B(i_7_), .Y(new_new_n686_));
  NO3        g664(.A(new_new_n471_), .B(new_new_n231_), .C(new_new_n81_), .Y(new_new_n687_));
  AOI210     g665(.A0(new_new_n687_), .A1(new_new_n686_), .B0(new_new_n685_), .Y(new_new_n688_));
  NA2        g666(.A(new_new_n379_), .B(new_new_n634_), .Y(new_new_n689_));
  OAI220     g667(.A0(new_new_n689_), .A1(new_new_n593_), .B0(new_new_n688_), .B1(new_new_n603_), .Y(new_new_n690_));
  NO4        g668(.A(new_new_n690_), .B(new_new_n684_), .C(new_new_n683_), .D(new_new_n681_), .Y(new_new_n691_));
  NA3        g669(.A(new_new_n406_), .B(new_new_n597_), .C(new_new_n93_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n626_), .B(i_13_), .Y(new_new_n693_));
  NAi21      g671(.An(i_11_), .B(i_12_), .Y(new_new_n694_));
  NOi41      g672(.An(new_new_n104_), .B(new_new_n694_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n695_));
  NO3        g673(.A(new_new_n471_), .B(new_new_n576_), .C(new_new_n598_), .Y(new_new_n696_));
  AOI210     g674(.A0(new_new_n696_), .A1(new_new_n305_), .B0(new_new_n695_), .Y(new_new_n697_));
  NA3        g675(.A(new_new_n697_), .B(new_new_n693_), .C(new_new_n692_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n698_), .B(new_new_n61_), .Y(new_new_n699_));
  NA2        g677(.A(i_8_), .B(new_new_n25_), .Y(new_new_n700_));
  NO3        g678(.A(new_new_n700_), .B(new_new_n377_), .C(i_12_), .Y(new_new_n701_));
  OAI210     g679(.A0(new_new_n701_), .A1(new_new_n362_), .B0(new_new_n360_), .Y(new_new_n702_));
  NO2        g680(.A(new_new_n121_), .B(i_2_), .Y(new_new_n703_));
  INV        g681(.A(new_new_n703_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n704_), .B(new_new_n702_), .Y(new_new_n705_));
  NA3        g683(.A(new_new_n705_), .B(new_new_n44_), .C(new_new_n219_), .Y(new_new_n706_));
  NA4        g684(.A(new_new_n706_), .B(new_new_n699_), .C(new_new_n691_), .D(new_new_n679_), .Y(new_new_n707_));
  OR4        g685(.A(new_new_n707_), .B(new_new_n672_), .C(new_new_n661_), .D(new_new_n604_), .Y(men5));
  AOI210     g686(.A0(new_new_n642_), .A1(new_new_n262_), .B0(new_new_n414_), .Y(new_new_n709_));
  NO3        g687(.A(i_11_), .B(new_new_n231_), .C(i_13_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n117_), .B(new_new_n23_), .Y(new_new_n711_));
  NA2        g689(.A(i_12_), .B(i_8_), .Y(new_new_n712_));
  OAI210     g690(.A0(new_new_n45_), .A1(i_3_), .B0(new_new_n712_), .Y(new_new_n713_));
  INV        g691(.A(new_new_n442_), .Y(new_new_n714_));
  AOI220     g692(.A0(new_new_n309_), .A1(new_new_n568_), .B0(new_new_n713_), .B1(new_new_n711_), .Y(new_new_n715_));
  INV        g693(.A(new_new_n715_), .Y(new_new_n716_));
  NO2        g694(.A(new_new_n716_), .B(new_new_n1013_), .Y(new_new_n717_));
  INV        g695(.A(new_new_n162_), .Y(new_new_n718_));
  INV        g696(.A(new_new_n238_), .Y(new_new_n719_));
  OAI210     g697(.A0(new_new_n670_), .A1(new_new_n444_), .B0(new_new_n104_), .Y(new_new_n720_));
  AOI210     g698(.A0(new_new_n720_), .A1(new_new_n719_), .B0(new_new_n718_), .Y(new_new_n721_));
  NO2        g699(.A(new_new_n451_), .B(new_new_n26_), .Y(new_new_n722_));
  NO2        g700(.A(new_new_n722_), .B(new_new_n415_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n723_), .B(i_2_), .Y(new_new_n724_));
  INV        g702(.A(new_new_n724_), .Y(new_new_n725_));
  AOI210     g703(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n412_), .Y(new_new_n726_));
  AOI210     g704(.A0(new_new_n726_), .A1(new_new_n725_), .B0(new_new_n721_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n182_), .B(new_new_n118_), .Y(new_new_n728_));
  OAI210     g706(.A0(new_new_n728_), .A1(new_new_n711_), .B0(i_2_), .Y(new_new_n729_));
  INV        g707(.A(new_new_n163_), .Y(new_new_n730_));
  NO3        g708(.A(new_new_n606_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n731_));
  AOI210     g709(.A0(new_new_n730_), .A1(new_new_n84_), .B0(new_new_n731_), .Y(new_new_n732_));
  AOI210     g710(.A0(new_new_n732_), .A1(new_new_n729_), .B0(new_new_n185_), .Y(new_new_n733_));
  OA210      g711(.A0(new_new_n607_), .A1(new_new_n119_), .B0(i_13_), .Y(new_new_n734_));
  AOI210     g712(.A0(new_new_n201_), .A1(new_new_n138_), .B0(new_new_n512_), .Y(new_new_n735_));
  NA2        g713(.A(new_new_n735_), .B(new_new_n415_), .Y(new_new_n736_));
  NA3        g714(.A(new_new_n298_), .B(new_new_n117_), .C(new_new_n41_), .Y(new_new_n737_));
  OAI210     g715(.A0(new_new_n737_), .A1(i_11_), .B0(new_new_n736_), .Y(new_new_n738_));
  NO3        g716(.A(new_new_n738_), .B(new_new_n734_), .C(new_new_n733_), .Y(new_new_n739_));
  NA2        g717(.A(new_new_n568_), .B(new_new_n28_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n710_), .B(new_new_n268_), .Y(new_new_n741_));
  NA2        g719(.A(new_new_n741_), .B(new_new_n740_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n60_), .B(i_12_), .Y(new_new_n743_));
  NO2        g721(.A(new_new_n743_), .B(new_new_n119_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n744_), .B(new_new_n591_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n745_), .A1(new_new_n36_), .B0(new_new_n742_), .Y(new_new_n746_));
  NA4        g724(.A(new_new_n746_), .B(new_new_n739_), .C(new_new_n727_), .D(new_new_n717_), .Y(men6));
  NO2        g725(.A(new_new_n177_), .B(i_9_), .Y(new_new_n748_));
  OAI210     g726(.A0(new_new_n748_), .A1(i_5_), .B0(new_new_n703_), .Y(new_new_n749_));
  NA4        g727(.A(new_new_n383_), .B(new_new_n476_), .C(new_new_n67_), .D(new_new_n97_), .Y(new_new_n750_));
  INV        g728(.A(new_new_n750_), .Y(new_new_n751_));
  NO2        g729(.A(new_new_n214_), .B(new_new_n481_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n751_), .B(new_new_n320_), .Y(new_new_n753_));
  AO210      g731(.A0(new_new_n753_), .A1(new_new_n749_), .B0(i_12_), .Y(new_new_n754_));
  NA2        g732(.A(new_new_n366_), .B(new_new_n327_), .Y(new_new_n755_));
  NA2        g733(.A(new_new_n576_), .B(new_new_n61_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n756_), .B(new_new_n755_), .Y(new_new_n757_));
  INV        g735(.A(new_new_n189_), .Y(new_new_n758_));
  AOI210     g736(.A0(new_new_n757_), .A1(new_new_n69_), .B0(new_new_n758_), .Y(new_new_n759_));
  NA2        g737(.A(new_new_n1014_), .B(new_new_n743_), .Y(new_new_n760_));
  NO2        g738(.A(new_new_n760_), .B(new_new_n177_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n32_), .B(i_11_), .Y(new_new_n762_));
  OAI210     g740(.A0(new_new_n662_), .A1(new_new_n556_), .B0(new_new_n555_), .Y(new_new_n763_));
  INV        g741(.A(new_new_n763_), .Y(new_new_n764_));
  OR2        g742(.A(new_new_n764_), .B(new_new_n761_), .Y(new_new_n765_));
  NA2        g743(.A(new_new_n47_), .B(new_new_n37_), .Y(new_new_n766_));
  OAI210     g744(.A0(new_new_n766_), .A1(new_new_n405_), .B0(new_new_n350_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n767_), .B(new_new_n1021_), .Y(new_new_n768_));
  AO210      g746(.A0(new_new_n349_), .A1(new_new_n341_), .B0(new_new_n391_), .Y(new_new_n769_));
  NA2        g747(.A(new_new_n769_), .B(i_7_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n444_), .B(new_new_n137_), .C(new_new_n65_), .Y(new_new_n771_));
  AO210      g749(.A0(new_new_n488_), .A1(new_new_n714_), .B0(new_new_n36_), .Y(new_new_n772_));
  NA4        g750(.A(new_new_n772_), .B(new_new_n771_), .C(new_new_n770_), .D(new_new_n768_), .Y(new_new_n773_));
  INV        g751(.A(new_new_n752_), .Y(new_new_n774_));
  NA3        g752(.A(new_new_n365_), .B(new_new_n232_), .C(new_new_n137_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n391_), .B(new_new_n66_), .Y(new_new_n776_));
  NA4        g754(.A(new_new_n776_), .B(new_new_n775_), .C(new_new_n774_), .D(new_new_n596_), .Y(new_new_n777_));
  AO210      g755(.A0(new_new_n512_), .A1(new_new_n45_), .B0(new_new_n83_), .Y(new_new_n778_));
  NA3        g756(.A(new_new_n778_), .B(new_new_n477_), .C(new_new_n211_), .Y(new_new_n779_));
  AOI210     g757(.A0(new_new_n444_), .A1(new_new_n442_), .B0(new_new_n554_), .Y(new_new_n780_));
  NA2        g758(.A(new_new_n237_), .B(new_new_n45_), .Y(new_new_n781_));
  INV        g759(.A(new_new_n582_), .Y(new_new_n782_));
  NA3        g760(.A(new_new_n782_), .B(new_new_n319_), .C(i_7_), .Y(new_new_n783_));
  NA4        g761(.A(new_new_n783_), .B(new_new_n1020_), .C(new_new_n780_), .D(new_new_n779_), .Y(new_new_n784_));
  NO4        g762(.A(new_new_n784_), .B(new_new_n777_), .C(new_new_n773_), .D(new_new_n765_), .Y(new_new_n785_));
  NA4        g763(.A(new_new_n785_), .B(new_new_n759_), .C(new_new_n754_), .D(new_new_n373_), .Y(men3));
  NA2        g764(.A(i_12_), .B(i_10_), .Y(new_new_n787_));
  NA2        g765(.A(i_6_), .B(i_7_), .Y(new_new_n788_));
  NO2        g766(.A(new_new_n788_), .B(i_0_), .Y(new_new_n789_));
  NO2        g767(.A(i_11_), .B(new_new_n231_), .Y(new_new_n790_));
  OAI210     g768(.A0(new_new_n789_), .A1(new_new_n283_), .B0(new_new_n790_), .Y(new_new_n791_));
  NO2        g769(.A(new_new_n791_), .B(new_new_n185_), .Y(new_new_n792_));
  NO3        g770(.A(new_new_n447_), .B(new_new_n86_), .C(new_new_n43_), .Y(new_new_n793_));
  OA210      g771(.A0(new_new_n793_), .A1(new_new_n792_), .B0(new_new_n165_), .Y(new_new_n794_));
  NA3        g772(.A(new_new_n775_), .B(new_new_n596_), .C(new_new_n364_), .Y(new_new_n795_));
  NA2        g773(.A(new_new_n795_), .B(new_new_n39_), .Y(new_new_n796_));
  NOi21      g774(.An(new_new_n92_), .B(new_new_n723_), .Y(new_new_n797_));
  NO3        g775(.A(new_new_n615_), .B(new_new_n451_), .C(new_new_n124_), .Y(new_new_n798_));
  NA2        g776(.A(new_new_n406_), .B(new_new_n44_), .Y(new_new_n799_));
  AN2        g777(.A(new_new_n449_), .B(new_new_n54_), .Y(new_new_n800_));
  NO3        g778(.A(new_new_n800_), .B(new_new_n798_), .C(new_new_n797_), .Y(new_new_n801_));
  AOI210     g779(.A0(new_new_n801_), .A1(new_new_n796_), .B0(new_new_n47_), .Y(new_new_n802_));
  NO4        g780(.A(new_new_n369_), .B(new_new_n376_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n177_), .B(new_new_n564_), .Y(new_new_n804_));
  NOi21      g782(.An(new_new_n804_), .B(new_new_n803_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n682_), .B(new_new_n652_), .Y(new_new_n806_));
  NA2        g784(.A(i_0_), .B(new_new_n434_), .Y(new_new_n807_));
  OAI220     g785(.A0(new_new_n807_), .A1(new_new_n806_), .B0(new_new_n805_), .B1(new_new_n61_), .Y(new_new_n808_));
  NOi21      g786(.An(i_5_), .B(i_9_), .Y(new_new_n809_));
  NA2        g787(.A(new_new_n809_), .B(new_new_n441_), .Y(new_new_n810_));
  NO3        g788(.A(new_new_n409_), .B(new_new_n259_), .C(new_new_n69_), .Y(new_new_n811_));
  NO2        g789(.A(new_new_n166_), .B(new_new_n138_), .Y(new_new_n812_));
  AOI210     g790(.A0(new_new_n812_), .A1(new_new_n237_), .B0(new_new_n811_), .Y(new_new_n813_));
  OAI220     g791(.A0(new_new_n813_), .A1(new_new_n172_), .B0(new_new_n598_), .B1(new_new_n810_), .Y(new_new_n814_));
  NO4        g792(.A(new_new_n814_), .B(new_new_n808_), .C(new_new_n802_), .D(new_new_n794_), .Y(new_new_n815_));
  NA2        g793(.A(new_new_n177_), .B(new_new_n24_), .Y(new_new_n816_));
  NO2        g794(.A(new_new_n650_), .B(new_new_n589_), .Y(new_new_n817_));
  NO2        g795(.A(new_new_n817_), .B(new_new_n816_), .Y(new_new_n818_));
  NA2        g796(.A(new_new_n305_), .B(new_new_n122_), .Y(new_new_n819_));
  NAi21      g797(.An(new_new_n153_), .B(new_new_n434_), .Y(new_new_n820_));
  OAI220     g798(.A0(new_new_n820_), .A1(new_new_n781_), .B0(new_new_n819_), .B1(new_new_n395_), .Y(new_new_n821_));
  NO2        g799(.A(new_new_n821_), .B(new_new_n818_), .Y(new_new_n822_));
  INV        g800(.A(new_new_n287_), .Y(new_new_n823_));
  NA2        g801(.A(new_new_n823_), .B(new_new_n684_), .Y(new_new_n824_));
  NA2        g802(.A(new_new_n565_), .B(i_0_), .Y(new_new_n825_));
  NO3        g803(.A(new_new_n825_), .B(new_new_n378_), .C(new_new_n84_), .Y(new_new_n826_));
  NO4        g804(.A(new_new_n581_), .B(new_new_n208_), .C(new_new_n412_), .D(new_new_n405_), .Y(new_new_n827_));
  AOI210     g805(.A0(new_new_n827_), .A1(i_11_), .B0(new_new_n826_), .Y(new_new_n828_));
  AN2        g806(.A(new_new_n92_), .B(new_new_n236_), .Y(new_new_n829_));
  NA2        g807(.A(new_new_n710_), .B(new_new_n320_), .Y(new_new_n830_));
  AOI210     g808(.A0(new_new_n477_), .A1(new_new_n84_), .B0(new_new_n57_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n831_), .B(new_new_n830_), .Y(new_new_n832_));
  NO2        g810(.A(new_new_n246_), .B(new_new_n144_), .Y(new_new_n833_));
  NA2        g811(.A(i_0_), .B(i_10_), .Y(new_new_n834_));
  OAI210     g812(.A0(new_new_n834_), .A1(new_new_n81_), .B0(new_new_n529_), .Y(new_new_n835_));
  NO4        g813(.A(new_new_n108_), .B(new_new_n57_), .C(new_new_n647_), .D(i_5_), .Y(new_new_n836_));
  AO220      g814(.A0(new_new_n836_), .A1(new_new_n835_), .B0(new_new_n833_), .B1(i_6_), .Y(new_new_n837_));
  NA2        g815(.A(new_new_n559_), .B(i_4_), .Y(new_new_n838_));
  OAI220     g816(.A0(i_1_), .A1(new_new_n830_), .B0(new_new_n838_), .B1(new_new_n1018_), .Y(new_new_n839_));
  NO4        g817(.A(new_new_n839_), .B(new_new_n837_), .C(new_new_n832_), .D(new_new_n829_), .Y(new_new_n840_));
  NA4        g818(.A(new_new_n840_), .B(new_new_n828_), .C(new_new_n824_), .D(new_new_n822_), .Y(new_new_n841_));
  NO2        g819(.A(new_new_n98_), .B(new_new_n37_), .Y(new_new_n842_));
  NA2        g820(.A(i_11_), .B(i_9_), .Y(new_new_n843_));
  NO3        g821(.A(i_12_), .B(new_new_n843_), .C(new_new_n595_), .Y(new_new_n844_));
  AN2        g822(.A(new_new_n844_), .B(new_new_n842_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n47_), .B(i_7_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n454_), .B(new_new_n151_), .Y(new_new_n847_));
  NO2        g825(.A(new_new_n843_), .B(new_new_n69_), .Y(new_new_n848_));
  NO2        g826(.A(new_new_n166_), .B(i_0_), .Y(new_new_n849_));
  INV        g827(.A(new_new_n849_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n469_), .B(new_new_n225_), .Y(new_new_n851_));
  INV        g829(.A(new_new_n403_), .Y(new_new_n852_));
  OAI220     g830(.A0(new_new_n852_), .A1(new_new_n810_), .B0(new_new_n851_), .B1(new_new_n850_), .Y(new_new_n853_));
  NO3        g831(.A(new_new_n853_), .B(new_new_n847_), .C(new_new_n845_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n637_), .B(new_new_n114_), .Y(new_new_n855_));
  NO2        g833(.A(i_6_), .B(new_new_n855_), .Y(new_new_n856_));
  AOI210     g834(.A0(new_new_n443_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n857_));
  NA2        g835(.A(new_new_n162_), .B(new_new_n98_), .Y(new_new_n858_));
  NOi32      g836(.An(new_new_n857_), .Bn(new_new_n180_), .C(new_new_n858_), .Y(new_new_n859_));
  AOI210     g837(.A0(new_new_n597_), .A1(new_new_n320_), .B0(new_new_n236_), .Y(new_new_n860_));
  NO2        g838(.A(new_new_n860_), .B(new_new_n799_), .Y(new_new_n861_));
  NO3        g839(.A(new_new_n861_), .B(new_new_n859_), .C(new_new_n856_), .Y(new_new_n862_));
  NOi21      g840(.An(i_7_), .B(i_5_), .Y(new_new_n863_));
  NOi31      g841(.An(new_new_n863_), .B(i_0_), .C(new_new_n694_), .Y(new_new_n864_));
  NA3        g842(.A(new_new_n864_), .B(new_new_n377_), .C(i_6_), .Y(new_new_n865_));
  OA210      g843(.A0(new_new_n858_), .A1(new_new_n510_), .B0(new_new_n865_), .Y(new_new_n866_));
  INV        g844(.A(new_new_n310_), .Y(new_new_n867_));
  NA3        g845(.A(new_new_n866_), .B(new_new_n862_), .C(new_new_n854_), .Y(new_new_n868_));
  NO2        g846(.A(new_new_n816_), .B(new_new_n233_), .Y(new_new_n869_));
  AN2        g847(.A(new_new_n325_), .B(new_new_n320_), .Y(new_new_n870_));
  AN2        g848(.A(new_new_n870_), .B(new_new_n812_), .Y(new_new_n871_));
  OAI210     g849(.A0(new_new_n871_), .A1(new_new_n869_), .B0(i_10_), .Y(new_new_n872_));
  NO2        g850(.A(new_new_n787_), .B(new_new_n309_), .Y(new_new_n873_));
  OA210      g851(.A0(new_new_n469_), .A1(new_new_n217_), .B0(new_new_n468_), .Y(new_new_n874_));
  NA2        g852(.A(new_new_n873_), .B(new_new_n848_), .Y(new_new_n875_));
  NA3        g853(.A(new_new_n468_), .B(new_new_n406_), .C(new_new_n44_), .Y(new_new_n876_));
  OAI210     g854(.A0(new_new_n820_), .A1(i_7_), .B0(new_new_n876_), .Y(new_new_n877_));
  NO2        g855(.A(new_new_n249_), .B(new_new_n45_), .Y(new_new_n878_));
  NA2        g856(.A(new_new_n848_), .B(new_new_n298_), .Y(new_new_n879_));
  OAI210     g857(.A0(new_new_n878_), .A1(new_new_n179_), .B0(new_new_n879_), .Y(new_new_n880_));
  AOI220     g858(.A0(new_new_n880_), .A1(new_new_n469_), .B0(new_new_n877_), .B1(new_new_n69_), .Y(new_new_n881_));
  NA3        g859(.A(new_new_n766_), .B(new_new_n375_), .C(i_6_), .Y(new_new_n882_));
  NA2        g860(.A(new_new_n88_), .B(new_new_n43_), .Y(new_new_n883_));
  NO2        g861(.A(new_new_n71_), .B(new_new_n712_), .Y(new_new_n884_));
  AOI220     g862(.A0(new_new_n884_), .A1(new_new_n883_), .B0(new_new_n165_), .B1(new_new_n589_), .Y(new_new_n885_));
  AOI210     g863(.A0(new_new_n885_), .A1(new_new_n882_), .B0(new_new_n46_), .Y(new_new_n886_));
  NO3        g864(.A(new_new_n581_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n887_));
  AOI210     g865(.A0(new_new_n676_), .A1(new_new_n537_), .B0(new_new_n887_), .Y(new_new_n888_));
  NAi21      g866(.An(i_9_), .B(i_5_), .Y(new_new_n889_));
  NO2        g867(.A(new_new_n889_), .B(new_new_n398_), .Y(new_new_n890_));
  NO2        g868(.A(new_new_n592_), .B(new_new_n100_), .Y(new_new_n891_));
  AOI220     g869(.A0(new_new_n891_), .A1(i_0_), .B0(new_new_n890_), .B1(new_new_n607_), .Y(new_new_n892_));
  OAI220     g870(.A0(new_new_n892_), .A1(new_new_n81_), .B0(new_new_n888_), .B1(new_new_n163_), .Y(new_new_n893_));
  NO3        g871(.A(new_new_n893_), .B(new_new_n886_), .C(new_new_n514_), .Y(new_new_n894_));
  NA4        g872(.A(new_new_n894_), .B(new_new_n881_), .C(new_new_n875_), .D(new_new_n872_), .Y(new_new_n895_));
  NO3        g873(.A(new_new_n895_), .B(new_new_n868_), .C(new_new_n841_), .Y(new_new_n896_));
  NO2        g874(.A(i_0_), .B(new_new_n694_), .Y(new_new_n897_));
  NA2        g875(.A(new_new_n69_), .B(new_new_n43_), .Y(new_new_n898_));
  NO3        g876(.A(new_new_n100_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n899_));
  AO220      g877(.A0(new_new_n899_), .A1(new_new_n43_), .B0(new_new_n897_), .B1(new_new_n165_), .Y(new_new_n900_));
  AOI210     g878(.A0(new_new_n756_), .A1(new_new_n664_), .B0(new_new_n858_), .Y(new_new_n901_));
  AOI210     g879(.A0(new_new_n900_), .A1(new_new_n338_), .B0(new_new_n901_), .Y(new_new_n902_));
  NA2        g880(.A(new_new_n703_), .B(new_new_n136_), .Y(new_new_n903_));
  NO2        g881(.A(new_new_n763_), .B(new_new_n398_), .Y(new_new_n904_));
  NA3        g882(.A(new_new_n789_), .B(i_2_), .C(new_new_n47_), .Y(new_new_n905_));
  NA2        g883(.A(new_new_n790_), .B(i_9_), .Y(new_new_n906_));
  AOI210     g884(.A0(new_new_n905_), .A1(new_new_n493_), .B0(new_new_n906_), .Y(new_new_n907_));
  OAI210     g885(.A0(new_new_n237_), .A1(i_9_), .B0(new_new_n224_), .Y(new_new_n908_));
  AOI210     g886(.A0(new_new_n908_), .A1(new_new_n825_), .B0(new_new_n144_), .Y(new_new_n909_));
  NO3        g887(.A(new_new_n909_), .B(new_new_n907_), .C(new_new_n904_), .Y(new_new_n910_));
  NA3        g888(.A(new_new_n910_), .B(new_new_n903_), .C(new_new_n902_), .Y(new_new_n911_));
  NA2        g889(.A(new_new_n870_), .B(new_new_n365_), .Y(new_new_n912_));
  AOI210     g890(.A0(new_new_n294_), .A1(new_new_n153_), .B0(new_new_n912_), .Y(new_new_n913_));
  INV        g891(.A(new_new_n913_), .Y(new_new_n914_));
  NO2        g892(.A(new_new_n834_), .B(new_new_n182_), .Y(new_new_n915_));
  NA2        g893(.A(new_new_n915_), .B(i_11_), .Y(new_new_n916_));
  NA2        g894(.A(new_new_n72_), .B(i_13_), .Y(new_new_n917_));
  INV        g895(.A(new_new_n211_), .Y(new_new_n918_));
  NO2        g896(.A(i_12_), .B(new_new_n603_), .Y(new_new_n919_));
  NA3        g897(.A(new_new_n919_), .B(new_new_n1015_), .C(new_new_n918_), .Y(new_new_n920_));
  NA4        g898(.A(new_new_n920_), .B(new_new_n917_), .C(new_new_n916_), .D(new_new_n914_), .Y(new_new_n921_));
  NO2        g899(.A(new_new_n235_), .B(new_new_n88_), .Y(new_new_n922_));
  AOI210     g900(.A0(new_new_n922_), .A1(new_new_n897_), .B0(new_new_n102_), .Y(new_new_n923_));
  AOI220     g901(.A0(new_new_n863_), .A1(new_new_n482_), .B0(new_new_n789_), .B1(new_new_n154_), .Y(new_new_n924_));
  NA2        g902(.A(new_new_n341_), .B(new_new_n167_), .Y(new_new_n925_));
  OA220      g903(.A0(new_new_n925_), .A1(new_new_n924_), .B0(new_new_n923_), .B1(i_5_), .Y(new_new_n926_));
  AOI210     g904(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n166_), .Y(new_new_n927_));
  NA2        g905(.A(new_new_n927_), .B(new_new_n874_), .Y(new_new_n928_));
  NA3        g906(.A(new_new_n601_), .B(new_new_n177_), .C(new_new_n79_), .Y(new_new_n929_));
  NA2        g907(.A(new_new_n929_), .B(new_new_n536_), .Y(new_new_n930_));
  NO3        g908(.A(new_new_n799_), .B(new_new_n53_), .C(new_new_n47_), .Y(new_new_n931_));
  NA3        g909(.A(new_new_n487_), .B(new_new_n480_), .C(new_new_n466_), .Y(new_new_n932_));
  NO3        g910(.A(new_new_n932_), .B(new_new_n931_), .C(new_new_n930_), .Y(new_new_n933_));
  NA2        g911(.A(new_new_n383_), .B(new_new_n161_), .Y(new_new_n934_));
  NA3        g912(.A(new_new_n383_), .B(new_new_n326_), .C(new_new_n215_), .Y(new_new_n935_));
  INV        g913(.A(new_new_n935_), .Y(new_new_n936_));
  NOi31      g914(.An(new_new_n382_), .B(new_new_n898_), .C(new_new_n233_), .Y(new_new_n937_));
  NO3        g915(.A(new_new_n937_), .B(new_new_n936_), .C(new_new_n1012_), .Y(new_new_n938_));
  NA4        g916(.A(new_new_n938_), .B(new_new_n933_), .C(new_new_n928_), .D(new_new_n926_), .Y(new_new_n939_));
  INV        g917(.A(new_new_n602_), .Y(new_new_n940_));
  NO3        g918(.A(new_new_n940_), .B(new_new_n550_), .C(i_3_), .Y(new_new_n941_));
  NO2        g919(.A(new_new_n81_), .B(i_5_), .Y(new_new_n942_));
  NA3        g920(.A(new_new_n790_), .B(new_new_n103_), .C(new_new_n117_), .Y(new_new_n943_));
  INV        g921(.A(new_new_n943_), .Y(new_new_n944_));
  AOI210     g922(.A0(new_new_n944_), .A1(new_new_n942_), .B0(new_new_n941_), .Y(new_new_n945_));
  NA3        g923(.A(new_new_n298_), .B(i_5_), .C(new_new_n185_), .Y(new_new_n946_));
  NO4        g924(.A(new_new_n233_), .B(new_new_n203_), .C(i_0_), .D(i_12_), .Y(new_new_n947_));
  AOI220     g925(.A0(new_new_n947_), .A1(i_10_), .B0(new_new_n751_), .B1(new_new_n167_), .Y(new_new_n948_));
  AN2        g926(.A(new_new_n834_), .B(new_new_n144_), .Y(new_new_n949_));
  NO4        g927(.A(new_new_n949_), .B(i_12_), .C(new_new_n632_), .D(new_new_n124_), .Y(new_new_n950_));
  NA2        g928(.A(new_new_n950_), .B(new_new_n211_), .Y(new_new_n951_));
  NA3        g929(.A(new_new_n94_), .B(new_new_n564_), .C(i_11_), .Y(new_new_n952_));
  NO2        g930(.A(new_new_n952_), .B(new_new_n146_), .Y(new_new_n953_));
  NA2        g931(.A(new_new_n863_), .B(new_new_n465_), .Y(new_new_n954_));
  NA2        g932(.A(new_new_n62_), .B(new_new_n97_), .Y(new_new_n955_));
  OAI220     g933(.A0(new_new_n955_), .A1(new_new_n946_), .B0(new_new_n954_), .B1(new_new_n653_), .Y(new_new_n956_));
  AOI210     g934(.A0(new_new_n956_), .A1(new_new_n849_), .B0(new_new_n953_), .Y(new_new_n957_));
  NA4        g935(.A(new_new_n957_), .B(new_new_n951_), .C(new_new_n948_), .D(new_new_n945_), .Y(new_new_n958_));
  NO4        g936(.A(new_new_n958_), .B(new_new_n939_), .C(new_new_n921_), .D(new_new_n911_), .Y(new_new_n959_));
  NA2        g937(.A(new_new_n762_), .B(new_new_n37_), .Y(new_new_n960_));
  NA3        g938(.A(new_new_n857_), .B(new_new_n360_), .C(i_5_), .Y(new_new_n961_));
  NA2        g939(.A(new_new_n961_), .B(new_new_n960_), .Y(new_new_n962_));
  NA2        g940(.A(new_new_n962_), .B(new_new_n199_), .Y(new_new_n963_));
  AN2        g941(.A(new_new_n673_), .B(new_new_n361_), .Y(new_new_n964_));
  NA2        g942(.A(new_new_n178_), .B(new_new_n180_), .Y(new_new_n965_));
  AO210      g943(.A0(new_new_n964_), .A1(new_new_n33_), .B0(new_new_n965_), .Y(new_new_n966_));
  NA2        g944(.A(new_new_n601_), .B(new_new_n309_), .Y(new_new_n967_));
  NAi31      g945(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n968_));
  NO2        g946(.A(new_new_n66_), .B(new_new_n968_), .Y(new_new_n969_));
  NO2        g947(.A(new_new_n969_), .B(new_new_n629_), .Y(new_new_n970_));
  NA3        g948(.A(new_new_n970_), .B(new_new_n967_), .C(new_new_n966_), .Y(new_new_n971_));
  NO2        g949(.A(new_new_n457_), .B(new_new_n259_), .Y(new_new_n972_));
  NO4        g950(.A(new_new_n227_), .B(new_new_n135_), .C(new_new_n656_), .D(new_new_n37_), .Y(new_new_n973_));
  NO3        g951(.A(new_new_n973_), .B(new_new_n972_), .C(new_new_n827_), .Y(new_new_n974_));
  OAI210     g952(.A0(new_new_n952_), .A1(new_new_n138_), .B0(new_new_n974_), .Y(new_new_n975_));
  AOI210     g953(.A0(new_new_n971_), .A1(new_new_n47_), .B0(new_new_n975_), .Y(new_new_n976_));
  AOI210     g954(.A0(new_new_n976_), .A1(new_new_n963_), .B0(new_new_n69_), .Y(new_new_n977_));
  INV        g955(.A(new_new_n372_), .Y(new_new_n978_));
  NO2        g956(.A(new_new_n978_), .B(new_new_n718_), .Y(new_new_n979_));
  OAI210     g957(.A0(new_new_n76_), .A1(new_new_n53_), .B0(new_new_n101_), .Y(new_new_n980_));
  NA2        g958(.A(new_new_n980_), .B(new_new_n72_), .Y(new_new_n981_));
  AOI210     g959(.A0(new_new_n927_), .A1(new_new_n846_), .B0(new_new_n864_), .Y(new_new_n982_));
  AOI210     g960(.A0(new_new_n982_), .A1(new_new_n981_), .B0(new_new_n656_), .Y(new_new_n983_));
  NA2        g961(.A(new_new_n256_), .B(new_new_n56_), .Y(new_new_n984_));
  AOI220     g962(.A0(new_new_n984_), .A1(new_new_n72_), .B0(new_new_n336_), .B1(new_new_n248_), .Y(new_new_n985_));
  NO2        g963(.A(new_new_n985_), .B(new_new_n231_), .Y(new_new_n986_));
  NA3        g964(.A(new_new_n92_), .B(new_new_n300_), .C(new_new_n31_), .Y(new_new_n987_));
  INV        g965(.A(new_new_n987_), .Y(new_new_n988_));
  NO3        g966(.A(new_new_n988_), .B(new_new_n986_), .C(new_new_n983_), .Y(new_new_n989_));
  OAI210     g967(.A0(new_new_n261_), .A1(new_new_n149_), .B0(new_new_n84_), .Y(new_new_n990_));
  NA3        g968(.A(new_new_n722_), .B(new_new_n283_), .C(new_new_n76_), .Y(new_new_n991_));
  AOI210     g969(.A0(new_new_n991_), .A1(new_new_n990_), .B0(i_11_), .Y(new_new_n992_));
  NA2        g970(.A(new_new_n598_), .B(new_new_n208_), .Y(new_new_n993_));
  OAI210     g971(.A0(new_new_n993_), .A1(new_new_n857_), .B0(new_new_n199_), .Y(new_new_n994_));
  NA2        g972(.A(new_new_n155_), .B(i_5_), .Y(new_new_n995_));
  NO2        g973(.A(new_new_n994_), .B(new_new_n995_), .Y(new_new_n996_));
  NO3        g974(.A(new_new_n58_), .B(new_new_n57_), .C(i_4_), .Y(new_new_n997_));
  OAI210     g975(.A0(new_new_n867_), .A1(new_new_n300_), .B0(new_new_n997_), .Y(new_new_n998_));
  NO2        g976(.A(new_new_n998_), .B(new_new_n694_), .Y(new_new_n999_));
  NO4        g977(.A(new_new_n889_), .B(i_11_), .C(i_3_), .D(new_new_n245_), .Y(new_new_n1000_));
  NO2        g978(.A(new_new_n1000_), .B(new_new_n554_), .Y(new_new_n1001_));
  INV        g979(.A(new_new_n353_), .Y(new_new_n1002_));
  AOI210     g980(.A0(new_new_n1002_), .A1(new_new_n1001_), .B0(new_new_n40_), .Y(new_new_n1003_));
  NO4        g981(.A(new_new_n1003_), .B(new_new_n999_), .C(new_new_n996_), .D(new_new_n992_), .Y(new_new_n1004_));
  OAI210     g982(.A0(new_new_n989_), .A1(i_4_), .B0(new_new_n1004_), .Y(new_new_n1005_));
  NO3        g983(.A(new_new_n1005_), .B(new_new_n979_), .C(new_new_n977_), .Y(new_new_n1006_));
  NA4        g984(.A(new_new_n1006_), .B(new_new_n959_), .C(new_new_n896_), .D(new_new_n815_), .Y(men4));
  INV        g985(.A(i_5_), .Y(new_new_n1010_));
  INV        g986(.A(i_1_), .Y(new_new_n1011_));
  INV        g987(.A(new_new_n934_), .Y(new_new_n1012_));
  INV        g988(.A(new_new_n709_), .Y(new_new_n1013_));
  INV        g989(.A(i_9_), .Y(new_new_n1014_));
  INV        g990(.A(i_3_), .Y(new_new_n1015_));
  INV        g991(.A(i_1_), .Y(new_new_n1016_));
  INV        g992(.A(new_new_n356_), .Y(new_new_n1017_));
  INV        g993(.A(new_new_n94_), .Y(new_new_n1018_));
  INV        g994(.A(i_0_), .Y(new_new_n1019_));
  INV        g995(.A(new_new_n404_), .Y(new_new_n1020_));
  INV        g996(.A(i_11_), .Y(new_new_n1021_));
  INV        g997(.A(i_3_), .Y(new_new_n1022_));
endmodule


