// Benchmark "top" written by ABC on Fri Jun 21 17:49:22 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n123_,
    new_new_n124_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n259_, new_new_n260_, new_new_n261_,
    new_new_n262_, new_new_n263_, new_new_n264_, new_new_n265_,
    new_new_n266_, new_new_n267_, new_new_n268_, new_new_n269_,
    new_new_n270_, new_new_n271_, new_new_n272_, new_new_n273_,
    new_new_n274_, new_new_n275_, new_new_n276_, new_new_n277_,
    new_new_n278_, new_new_n279_, new_new_n280_, new_new_n281_,
    new_new_n282_, new_new_n283_, new_new_n284_, new_new_n285_,
    new_new_n286_, new_new_n287_, new_new_n288_, new_new_n289_,
    new_new_n290_, new_new_n291_, new_new_n292_, new_new_n293_,
    new_new_n294_, new_new_n295_, new_new_n296_, new_new_n297_,
    new_new_n298_, new_new_n299_, new_new_n300_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n314_, new_new_n315_, new_new_n316_, new_new_n317_,
    new_new_n318_, new_new_n319_, new_new_n320_, new_new_n321_,
    new_new_n322_, new_new_n323_, new_new_n324_, new_new_n325_,
    new_new_n326_, new_new_n327_, new_new_n328_, new_new_n329_,
    new_new_n330_, new_new_n331_, new_new_n332_, new_new_n333_,
    new_new_n334_, new_new_n335_, new_new_n336_, new_new_n337_,
    new_new_n338_, new_new_n339_, new_new_n340_, new_new_n341_,
    new_new_n342_, new_new_n343_, new_new_n344_, new_new_n345_,
    new_new_n346_, new_new_n347_, new_new_n348_, new_new_n349_,
    new_new_n351_, new_new_n352_, new_new_n353_, new_new_n354_,
    new_new_n355_, new_new_n356_, new_new_n357_, new_new_n358_,
    new_new_n359_, new_new_n360_, new_new_n361_, new_new_n362_,
    new_new_n363_, new_new_n364_, new_new_n365_, new_new_n366_,
    new_new_n367_, new_new_n368_, new_new_n369_, new_new_n370_,
    new_new_n371_, new_new_n372_, new_new_n373_, new_new_n374_,
    new_new_n375_, new_new_n376_, new_new_n377_, new_new_n378_,
    new_new_n379_, new_new_n380_, new_new_n381_, new_new_n382_,
    new_new_n383_, new_new_n384_, new_new_n385_, new_new_n386_,
    new_new_n387_, new_new_n388_, new_new_n389_, new_new_n390_,
    new_new_n391_, new_new_n392_, new_new_n393_, new_new_n394_,
    new_new_n395_, new_new_n397_, new_new_n398_, new_new_n399_,
    new_new_n400_, new_new_n401_, new_new_n402_, new_new_n403_,
    new_new_n404_, new_new_n405_, new_new_n406_, new_new_n407_,
    new_new_n408_, new_new_n409_, new_new_n410_, new_new_n411_,
    new_new_n412_, new_new_n413_, new_new_n414_, new_new_n415_,
    new_new_n416_, new_new_n417_, new_new_n418_, new_new_n419_,
    new_new_n420_, new_new_n421_, new_new_n422_, new_new_n423_,
    new_new_n424_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n504_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  OAI210     g027(.A0(new_new_n49_), .A1(i_3_), .B0(new_new_n47_), .Y(new_new_n50_));
  NO2        g028(.A(new_new_n50_), .B(new_new_n46_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NA2        g030(.A(new_new_n51_), .B(new_new_n45_), .Y(new_new_n53_));
  NO2        g031(.A(i_1_), .B(i_6_), .Y(new_new_n54_));
  NAi21      g032(.An(i_2_), .B(i_7_), .Y(new_new_n55_));
  INV        g033(.A(i_1_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n56_), .B(i_6_), .Y(new_new_n57_));
  NA3        g035(.A(new_new_n57_), .B(new_new_n55_), .C(new_new_n31_), .Y(new_new_n58_));
  NA2        g036(.A(i_1_), .B(i_10_), .Y(new_new_n59_));
  NO2        g037(.A(new_new_n59_), .B(i_6_), .Y(new_new_n60_));
  NAi21      g038(.An(new_new_n60_), .B(new_new_n58_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n49_), .B(i_2_), .Y(new_new_n62_));
  AOI210     g040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(i_1_), .B(i_6_), .Y(new_new_n64_));
  NO2        g042(.A(new_new_n64_), .B(new_new_n25_), .Y(new_new_n65_));
  INV        g043(.A(i_0_), .Y(new_new_n66_));
  NAi21      g044(.An(i_5_), .B(i_10_), .Y(new_new_n67_));
  NA2        g045(.A(i_5_), .B(i_9_), .Y(new_new_n68_));
  AOI210     g046(.A0(new_new_n68_), .A1(new_new_n67_), .B0(new_new_n66_), .Y(new_new_n69_));
  NO2        g047(.A(new_new_n69_), .B(new_new_n65_), .Y(new_new_n70_));
  OAI210     g048(.A0(new_new_n63_), .A1(new_new_n62_), .B0(new_new_n70_), .Y(new_new_n71_));
  OAI210     g049(.A0(new_new_n71_), .A1(new_new_n61_), .B0(i_0_), .Y(new_new_n72_));
  NA2        g050(.A(i_12_), .B(i_5_), .Y(new_new_n73_));
  INV        g051(.A(i_8_), .Y(new_new_n74_));
  NO2        g052(.A(new_new_n74_), .B(new_new_n54_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_9_), .Y(new_new_n76_));
  NO2        g054(.A(i_3_), .B(i_7_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n76_), .B(new_new_n56_), .Y(new_new_n78_));
  INV        g056(.A(i_6_), .Y(new_new_n79_));
  NO2        g057(.A(i_2_), .B(i_7_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n80_), .Y(new_new_n81_));
  OAI210     g059(.A0(new_new_n78_), .A1(new_new_n75_), .B0(new_new_n81_), .Y(new_new_n82_));
  NAi21      g060(.An(i_6_), .B(i_10_), .Y(new_new_n83_));
  NA2        g061(.A(i_6_), .B(i_9_), .Y(new_new_n84_));
  AOI210     g062(.A0(new_new_n84_), .A1(new_new_n83_), .B0(new_new_n56_), .Y(new_new_n85_));
  NA2        g063(.A(i_2_), .B(i_6_), .Y(new_new_n86_));
  NO2        g064(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n87_));
  NO2        g065(.A(new_new_n87_), .B(new_new_n85_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n88_), .A1(new_new_n82_), .B0(new_new_n73_), .Y(new_new_n89_));
  AN3        g067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n90_));
  NAi21      g068(.An(i_6_), .B(i_11_), .Y(new_new_n91_));
  NA2        g069(.A(new_new_n90_), .B(new_new_n32_), .Y(new_new_n92_));
  INV        g070(.A(i_7_), .Y(new_new_n93_));
  NA2        g071(.A(new_new_n46_), .B(new_new_n93_), .Y(new_new_n94_));
  NO2        g072(.A(i_0_), .B(i_5_), .Y(new_new_n95_));
  NO2        g073(.A(new_new_n95_), .B(new_new_n79_), .Y(new_new_n96_));
  NA2        g074(.A(i_12_), .B(i_3_), .Y(new_new_n97_));
  INV        g075(.A(new_new_n97_), .Y(new_new_n98_));
  NA3        g076(.A(new_new_n98_), .B(new_new_n96_), .C(new_new_n94_), .Y(new_new_n99_));
  NAi21      g077(.An(i_7_), .B(i_11_), .Y(new_new_n100_));
  AN2        g078(.A(i_2_), .B(i_10_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n101_), .B(i_7_), .Y(new_new_n102_));
  OR2        g080(.A(new_new_n73_), .B(new_new_n54_), .Y(new_new_n103_));
  NA2        g081(.A(i_12_), .B(i_7_), .Y(new_new_n104_));
  NA2        g082(.A(i_11_), .B(i_12_), .Y(new_new_n105_));
  NA3        g083(.A(new_new_n105_), .B(new_new_n99_), .C(new_new_n92_), .Y(new_new_n106_));
  NOi21      g084(.An(i_1_), .B(i_5_), .Y(new_new_n107_));
  NA2        g085(.A(new_new_n107_), .B(i_11_), .Y(new_new_n108_));
  NA2        g086(.A(new_new_n93_), .B(new_new_n37_), .Y(new_new_n109_));
  NA2        g087(.A(i_7_), .B(new_new_n25_), .Y(new_new_n110_));
  NA2        g088(.A(new_new_n110_), .B(new_new_n109_), .Y(new_new_n111_));
  NO2        g089(.A(new_new_n111_), .B(new_new_n46_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n84_), .B(new_new_n83_), .Y(new_new_n113_));
  NAi21      g091(.An(i_3_), .B(i_8_), .Y(new_new_n114_));
  NA2        g092(.A(new_new_n114_), .B(new_new_n55_), .Y(new_new_n115_));
  NOi31      g093(.An(new_new_n115_), .B(new_new_n113_), .C(new_new_n112_), .Y(new_new_n116_));
  NO2        g094(.A(i_1_), .B(new_new_n79_), .Y(new_new_n117_));
  NO2        g095(.A(i_6_), .B(i_5_), .Y(new_new_n118_));
  NA2        g096(.A(new_new_n118_), .B(i_3_), .Y(new_new_n119_));
  OAI220     g097(.A0(new_new_n119_), .A1(new_new_n100_), .B0(new_new_n116_), .B1(new_new_n108_), .Y(new_new_n120_));
  NO3        g098(.A(new_new_n120_), .B(new_new_n106_), .C(new_new_n89_), .Y(new_new_n121_));
  NA3        g099(.A(new_new_n121_), .B(new_new_n72_), .C(new_new_n53_), .Y(ori2));
  NO2        g100(.A(new_new_n56_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n504_), .B(new_new_n123_), .Y(new_new_n124_));
  NA4        g102(.A(new_new_n124_), .B(new_new_n70_), .C(new_new_n62_), .D(new_new_n30_), .Y(ori0));
  NO2        g103(.A(i_0_), .B(i_1_), .Y(new_new_n126_));
  NA2        g104(.A(i_2_), .B(i_3_), .Y(new_new_n127_));
  NO2        g105(.A(new_new_n127_), .B(i_4_), .Y(new_new_n128_));
  NA2        g106(.A(i_1_), .B(i_5_), .Y(new_new_n129_));
  OR2        g107(.A(i_0_), .B(i_1_), .Y(new_new_n130_));
  NO3        g108(.A(new_new_n130_), .B(new_new_n73_), .C(i_13_), .Y(new_new_n131_));
  NAi32      g109(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n132_));
  NAi21      g110(.An(new_new_n132_), .B(new_new_n131_), .Y(new_new_n133_));
  NOi21      g111(.An(i_4_), .B(i_10_), .Y(new_new_n134_));
  NOi21      g112(.An(i_4_), .B(i_9_), .Y(new_new_n135_));
  NOi21      g113(.An(i_11_), .B(i_13_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(new_new_n135_), .Y(new_new_n137_));
  NO2        g115(.A(new_new_n66_), .B(new_new_n56_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n66_), .B(i_5_), .Y(new_new_n139_));
  NO2        g117(.A(i_2_), .B(i_1_), .Y(new_new_n140_));
  NAi21      g118(.An(i_4_), .B(i_12_), .Y(new_new_n141_));
  INV        g119(.A(i_8_), .Y(new_new_n142_));
  NO2        g120(.A(i_3_), .B(i_8_), .Y(new_new_n143_));
  NO3        g121(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n144_));
  NO2        g122(.A(new_new_n95_), .B(new_new_n54_), .Y(new_new_n145_));
  NO2        g123(.A(i_13_), .B(i_9_), .Y(new_new_n146_));
  NAi21      g124(.An(i_12_), .B(i_3_), .Y(new_new_n147_));
  NO2        g125(.A(new_new_n44_), .B(i_5_), .Y(new_new_n148_));
  NA2        g126(.A(i_0_), .B(i_5_), .Y(new_new_n149_));
  INV        g127(.A(i_13_), .Y(new_new_n150_));
  NO2        g128(.A(i_12_), .B(new_new_n150_), .Y(new_new_n151_));
  NO2        g129(.A(i_12_), .B(new_new_n37_), .Y(new_new_n152_));
  OR2        g130(.A(i_8_), .B(i_7_), .Y(new_new_n153_));
  INV        g131(.A(i_12_), .Y(new_new_n154_));
  NO2        g132(.A(new_new_n44_), .B(new_new_n154_), .Y(new_new_n155_));
  NA2        g133(.A(i_2_), .B(i_1_), .Y(new_new_n156_));
  NO3        g134(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n157_));
  NAi21      g135(.An(i_4_), .B(i_3_), .Y(new_new_n158_));
  NO2        g136(.A(i_0_), .B(i_6_), .Y(new_new_n159_));
  NOi41      g137(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n160_));
  NO2        g138(.A(i_11_), .B(new_new_n150_), .Y(new_new_n161_));
  NOi21      g139(.An(i_1_), .B(i_6_), .Y(new_new_n162_));
  NAi21      g140(.An(i_3_), .B(i_7_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n154_), .B(i_9_), .Y(new_new_n164_));
  OR4        g142(.A(new_new_n164_), .B(new_new_n163_), .C(new_new_n162_), .D(new_new_n139_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n66_), .B(i_5_), .Y(new_new_n166_));
  NA2        g144(.A(i_3_), .B(i_9_), .Y(new_new_n167_));
  NAi21      g145(.An(i_7_), .B(i_10_), .Y(new_new_n168_));
  NO2        g146(.A(new_new_n168_), .B(new_new_n167_), .Y(new_new_n169_));
  NA3        g147(.A(new_new_n169_), .B(new_new_n166_), .C(new_new_n57_), .Y(new_new_n170_));
  NA2        g148(.A(new_new_n170_), .B(new_new_n165_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n171_), .B(new_new_n161_), .Y(new_new_n172_));
  NA2        g150(.A(i_12_), .B(i_6_), .Y(new_new_n173_));
  OR2        g151(.A(i_13_), .B(i_9_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n158_), .B(i_2_), .Y(new_new_n175_));
  NO2        g153(.A(new_new_n163_), .B(i_8_), .Y(new_new_n176_));
  NO3        g154(.A(i_12_), .B(new_new_n150_), .C(new_new_n37_), .Y(new_new_n177_));
  NO2        g155(.A(i_2_), .B(new_new_n93_), .Y(new_new_n178_));
  AN2        g156(.A(i_3_), .B(i_10_), .Y(new_new_n179_));
  NO2        g157(.A(i_5_), .B(new_new_n37_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n181_));
  NO2        g159(.A(i_2_), .B(i_3_), .Y(new_new_n182_));
  NO2        g160(.A(i_12_), .B(i_10_), .Y(new_new_n183_));
  NOi21      g161(.An(i_5_), .B(i_0_), .Y(new_new_n184_));
  NOi32      g162(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n185_));
  INV        g163(.A(new_new_n185_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n132_), .B(new_new_n130_), .Y(new_new_n187_));
  NOi32      g165(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n188_));
  NO2        g166(.A(i_1_), .B(new_new_n93_), .Y(new_new_n189_));
  NAi21      g167(.An(i_3_), .B(i_4_), .Y(new_new_n190_));
  NO2        g168(.A(new_new_n190_), .B(i_9_), .Y(new_new_n191_));
  AN2        g169(.A(i_6_), .B(i_7_), .Y(new_new_n192_));
  OAI210     g170(.A0(new_new_n192_), .A1(new_new_n189_), .B0(new_new_n191_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n190_), .B(i_10_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n193_), .B(new_new_n139_), .Y(new_new_n195_));
  AOI210     g173(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n196_));
  OAI210     g174(.A0(new_new_n196_), .A1(new_new_n140_), .B0(new_new_n194_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n197_), .B(i_5_), .Y(new_new_n198_));
  NO3        g176(.A(new_new_n198_), .B(new_new_n195_), .C(new_new_n187_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n199_), .B(new_new_n186_), .Y(new_new_n200_));
  AN2        g178(.A(i_12_), .B(i_5_), .Y(new_new_n201_));
  NO2        g179(.A(i_11_), .B(i_6_), .Y(new_new_n202_));
  NO2        g180(.A(i_5_), .B(i_10_), .Y(new_new_n203_));
  NO2        g181(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n204_));
  NO3        g182(.A(new_new_n79_), .B(new_new_n47_), .C(i_9_), .Y(new_new_n205_));
  NO2        g183(.A(i_0_), .B(i_11_), .Y(new_new_n206_));
  NOi21      g184(.An(i_2_), .B(i_12_), .Y(new_new_n207_));
  NAi21      g185(.An(i_9_), .B(i_4_), .Y(new_new_n208_));
  OR2        g186(.A(i_13_), .B(i_10_), .Y(new_new_n209_));
  NO3        g187(.A(new_new_n209_), .B(new_new_n105_), .C(new_new_n208_), .Y(new_new_n210_));
  NO2        g188(.A(new_new_n93_), .B(new_new_n25_), .Y(new_new_n211_));
  INV        g189(.A(new_new_n200_), .Y(new_new_n212_));
  NO2        g190(.A(new_new_n66_), .B(i_13_), .Y(new_new_n213_));
  NO2        g191(.A(i_10_), .B(i_9_), .Y(new_new_n214_));
  NAi21      g192(.An(i_12_), .B(i_8_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n215_), .B(i_3_), .Y(new_new_n216_));
  NO3        g194(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n217_));
  NA2        g195(.A(new_new_n173_), .B(new_new_n91_), .Y(new_new_n218_));
  NA2        g196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  NA2        g197(.A(i_8_), .B(i_9_), .Y(new_new_n220_));
  NO2        g198(.A(i_7_), .B(i_2_), .Y(new_new_n221_));
  OR2        g199(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n222_));
  NA2        g200(.A(new_new_n177_), .B(new_new_n145_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  NA2        g202(.A(new_new_n161_), .B(new_new_n180_), .Y(new_new_n225_));
  NO3        g203(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n226_));
  INV        g204(.A(new_new_n226_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n227_), .B(new_new_n225_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n228_), .B(new_new_n224_), .Y(new_new_n229_));
  NO2        g207(.A(i_11_), .B(i_1_), .Y(new_new_n230_));
  NOi21      g208(.An(i_2_), .B(i_7_), .Y(new_new_n231_));
  NA3        g209(.A(new_new_n160_), .B(new_new_n136_), .C(new_new_n118_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n130_), .B(i_3_), .Y(new_new_n234_));
  NAi31      g212(.An(new_new_n233_), .B(new_new_n234_), .C(new_new_n151_), .Y(new_new_n235_));
  NA3        g213(.A(new_new_n204_), .B(new_new_n138_), .C(new_new_n128_), .Y(new_new_n236_));
  NA3        g214(.A(new_new_n236_), .B(new_new_n235_), .C(new_new_n232_), .Y(new_new_n237_));
  INV        g215(.A(new_new_n237_), .Y(new_new_n238_));
  NA2        g216(.A(new_new_n217_), .B(new_new_n201_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n226_), .B(new_new_n203_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n238_), .B(new_new_n229_), .Y(new_new_n241_));
  NA2        g219(.A(new_new_n201_), .B(new_new_n150_), .Y(new_new_n242_));
  NA2        g220(.A(new_new_n192_), .B(new_new_n188_), .Y(new_new_n243_));
  OR2        g221(.A(new_new_n242_), .B(new_new_n243_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n36_), .B(i_8_), .Y(new_new_n245_));
  AOI210     g223(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n210_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n246_), .B(new_new_n244_), .Y(new_new_n247_));
  NA3        g225(.A(new_new_n149_), .B(new_new_n64_), .C(new_new_n44_), .Y(new_new_n248_));
  NA2        g226(.A(new_new_n177_), .B(new_new_n77_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n248_), .B(new_new_n249_), .Y(new_new_n250_));
  NO3        g228(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n251_));
  NO2        g229(.A(new_new_n209_), .B(i_1_), .Y(new_new_n252_));
  NOi31      g230(.An(new_new_n252_), .B(new_new_n218_), .C(new_new_n66_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n79_), .B(new_new_n25_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n104_), .B(new_new_n23_), .Y(new_new_n255_));
  NO2        g233(.A(i_12_), .B(new_new_n79_), .Y(new_new_n256_));
  NO3        g234(.A(new_new_n250_), .B(new_new_n247_), .C(new_new_n241_), .Y(new_new_n257_));
  NA3        g235(.A(new_new_n257_), .B(new_new_n212_), .C(new_new_n172_), .Y(ori7));
  NO2        g236(.A(new_new_n86_), .B(new_new_n52_), .Y(new_new_n259_));
  NA2        g237(.A(i_11_), .B(new_new_n142_), .Y(new_new_n260_));
  NA3        g238(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n154_), .B(i_4_), .Y(new_new_n262_));
  NA2        g240(.A(new_new_n262_), .B(i_8_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n97_), .B(new_new_n261_), .Y(new_new_n264_));
  NA2        g242(.A(i_2_), .B(new_new_n79_), .Y(new_new_n265_));
  OAI210     g243(.A0(new_new_n80_), .A1(new_new_n143_), .B0(new_new_n144_), .Y(new_new_n266_));
  NO2        g244(.A(i_7_), .B(new_new_n37_), .Y(new_new_n267_));
  NA2        g245(.A(i_4_), .B(i_8_), .Y(new_new_n268_));
  AOI210     g246(.A0(new_new_n268_), .A1(new_new_n179_), .B0(new_new_n267_), .Y(new_new_n269_));
  OAI220     g247(.A0(new_new_n269_), .A1(new_new_n265_), .B0(new_new_n266_), .B1(i_13_), .Y(new_new_n270_));
  NO3        g248(.A(new_new_n270_), .B(new_new_n264_), .C(new_new_n259_), .Y(new_new_n271_));
  AOI210     g249(.A0(new_new_n114_), .A1(new_new_n55_), .B0(i_10_), .Y(new_new_n272_));
  AOI210     g250(.A0(new_new_n272_), .A1(new_new_n154_), .B0(new_new_n134_), .Y(new_new_n273_));
  OR2        g251(.A(i_6_), .B(i_10_), .Y(new_new_n274_));
  OR3        g252(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n275_));
  OR2        g253(.A(new_new_n273_), .B(new_new_n174_), .Y(new_new_n276_));
  AOI210     g254(.A0(new_new_n276_), .A1(new_new_n271_), .B0(new_new_n56_), .Y(new_new_n277_));
  NOi21      g255(.An(i_11_), .B(i_7_), .Y(new_new_n278_));
  AO210      g256(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(new_new_n278_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n280_), .B(new_new_n146_), .Y(new_new_n281_));
  NO2        g259(.A(new_new_n281_), .B(new_new_n56_), .Y(new_new_n282_));
  NA2        g260(.A(new_new_n151_), .B(new_new_n56_), .Y(new_new_n283_));
  NO2        g261(.A(i_1_), .B(i_12_), .Y(new_new_n284_));
  INV        g262(.A(new_new_n283_), .Y(new_new_n285_));
  OAI210     g263(.A0(new_new_n285_), .A1(new_new_n282_), .B0(i_6_), .Y(new_new_n286_));
  NO2        g264(.A(i_6_), .B(i_11_), .Y(new_new_n287_));
  INV        g265(.A(new_new_n219_), .Y(new_new_n288_));
  NO3        g266(.A(new_new_n274_), .B(new_new_n153_), .C(new_new_n23_), .Y(new_new_n289_));
  AOI210     g267(.A0(i_1_), .A1(new_new_n169_), .B0(new_new_n289_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(new_new_n44_), .Y(new_new_n291_));
  INV        g269(.A(i_2_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n123_), .B(i_9_), .Y(new_new_n293_));
  NO2        g271(.A(new_new_n46_), .B(i_1_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n293_), .B(new_new_n292_), .Y(new_new_n295_));
  AOI210     g273(.A0(new_new_n230_), .A1(new_new_n211_), .B0(new_new_n157_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n296_), .B(new_new_n265_), .Y(new_new_n297_));
  NO2        g275(.A(i_11_), .B(new_new_n37_), .Y(new_new_n298_));
  OR2        g276(.A(new_new_n297_), .B(new_new_n295_), .Y(new_new_n299_));
  NO3        g277(.A(new_new_n299_), .B(new_new_n291_), .C(new_new_n288_), .Y(new_new_n300_));
  NO2        g278(.A(new_new_n154_), .B(new_new_n93_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(new_new_n278_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n302_), .B(i_1_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n303_), .B(new_new_n275_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n208_), .B(new_new_n79_), .Y(new_new_n305_));
  NA2        g283(.A(new_new_n304_), .B(new_new_n46_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n153_), .B(new_new_n44_), .Y(new_new_n307_));
  NO3        g285(.A(new_new_n307_), .B(new_new_n181_), .C(new_new_n155_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n309_), .B(i_6_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n79_), .B(i_9_), .Y(new_new_n311_));
  NO2        g289(.A(new_new_n311_), .B(new_new_n56_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n312_), .B(new_new_n284_), .Y(new_new_n313_));
  NO4        g291(.A(new_new_n313_), .B(new_new_n310_), .C(new_new_n308_), .D(i_4_), .Y(new_new_n314_));
  INV        g292(.A(new_new_n314_), .Y(new_new_n315_));
  NA4        g293(.A(new_new_n315_), .B(new_new_n306_), .C(new_new_n300_), .D(new_new_n286_), .Y(new_new_n316_));
  AOI210     g294(.A0(new_new_n173_), .A1(new_new_n91_), .B0(i_1_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n190_), .B(i_2_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n318_), .B(new_new_n317_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n319_), .B(i_13_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n52_), .B(i_12_), .Y(new_new_n321_));
  INV        g299(.A(new_new_n321_), .Y(new_new_n322_));
  NO2        g300(.A(new_new_n231_), .B(new_new_n24_), .Y(new_new_n323_));
  NA2        g301(.A(new_new_n323_), .B(new_new_n305_), .Y(new_new_n324_));
  OAI220     g302(.A0(new_new_n324_), .A1(new_new_n41_), .B0(new_new_n322_), .B1(new_new_n86_), .Y(new_new_n325_));
  INV        g303(.A(new_new_n325_), .Y(new_new_n326_));
  NA2        g304(.A(new_new_n202_), .B(new_new_n294_), .Y(new_new_n327_));
  NO2        g305(.A(new_new_n327_), .B(new_new_n158_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n113_), .B(i_13_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n329_), .B(new_new_n317_), .Y(new_new_n330_));
  NA2        g308(.A(new_new_n26_), .B(new_new_n142_), .Y(new_new_n331_));
  AOI220     g309(.A0(new_new_n202_), .A1(new_new_n294_), .B0(new_new_n85_), .B1(new_new_n94_), .Y(new_new_n332_));
  NO2        g310(.A(new_new_n332_), .B(new_new_n263_), .Y(new_new_n333_));
  NO3        g311(.A(new_new_n333_), .B(new_new_n330_), .C(new_new_n328_), .Y(new_new_n334_));
  OR2        g312(.A(i_11_), .B(i_6_), .Y(new_new_n335_));
  NA3        g313(.A(new_new_n262_), .B(new_new_n331_), .C(i_7_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n336_), .B(new_new_n335_), .Y(new_new_n337_));
  NA3        g315(.A(new_new_n207_), .B(new_new_n267_), .C(new_new_n91_), .Y(new_new_n338_));
  NA2        g316(.A(new_new_n287_), .B(i_13_), .Y(new_new_n339_));
  NAi21      g317(.An(i_11_), .B(i_12_), .Y(new_new_n340_));
  NOi41      g318(.An(new_new_n102_), .B(new_new_n340_), .C(i_13_), .D(new_new_n79_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n46_), .Y(new_new_n342_));
  NA3        g320(.A(new_new_n342_), .B(new_new_n339_), .C(new_new_n338_), .Y(new_new_n343_));
  OAI210     g321(.A0(new_new_n343_), .A1(new_new_n337_), .B0(new_new_n56_), .Y(new_new_n344_));
  NO2        g322(.A(i_2_), .B(i_12_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n189_), .B(new_new_n345_), .Y(new_new_n346_));
  INV        g324(.A(new_new_n346_), .Y(new_new_n347_));
  NA3        g325(.A(new_new_n347_), .B(new_new_n45_), .C(new_new_n150_), .Y(new_new_n348_));
  NA4        g326(.A(new_new_n348_), .B(new_new_n344_), .C(new_new_n334_), .D(new_new_n326_), .Y(new_new_n349_));
  OR4        g327(.A(new_new_n349_), .B(new_new_n320_), .C(new_new_n316_), .D(new_new_n277_), .Y(ori5));
  NA2        g328(.A(new_new_n302_), .B(new_new_n175_), .Y(new_new_n351_));
  AN2        g329(.A(new_new_n24_), .B(i_10_), .Y(new_new_n352_));
  NA3        g330(.A(new_new_n352_), .B(new_new_n345_), .C(new_new_n100_), .Y(new_new_n353_));
  NO2        g331(.A(new_new_n263_), .B(i_11_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n80_), .B(new_new_n354_), .Y(new_new_n355_));
  NA3        g333(.A(new_new_n355_), .B(new_new_n353_), .C(new_new_n351_), .Y(new_new_n356_));
  NO3        g334(.A(i_11_), .B(new_new_n154_), .C(i_13_), .Y(new_new_n357_));
  NO2        g335(.A(new_new_n110_), .B(new_new_n23_), .Y(new_new_n358_));
  NA2        g336(.A(i_12_), .B(i_8_), .Y(new_new_n359_));
  OAI210     g337(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n359_), .Y(new_new_n360_));
  INV        g338(.A(new_new_n214_), .Y(new_new_n361_));
  AOI220     g339(.A0(new_new_n182_), .A1(new_new_n255_), .B0(new_new_n360_), .B1(new_new_n358_), .Y(new_new_n362_));
  INV        g340(.A(new_new_n362_), .Y(new_new_n363_));
  NO2        g341(.A(new_new_n363_), .B(new_new_n356_), .Y(new_new_n364_));
  INV        g342(.A(new_new_n136_), .Y(new_new_n365_));
  INV        g343(.A(new_new_n160_), .Y(new_new_n366_));
  OAI210     g344(.A0(new_new_n318_), .A1(new_new_n216_), .B0(new_new_n102_), .Y(new_new_n367_));
  AOI210     g345(.A0(new_new_n367_), .A1(new_new_n366_), .B0(new_new_n365_), .Y(new_new_n368_));
  NO2        g346(.A(new_new_n220_), .B(new_new_n26_), .Y(new_new_n369_));
  NO2        g347(.A(new_new_n369_), .B(new_new_n211_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n370_), .B(i_2_), .Y(new_new_n371_));
  INV        g349(.A(new_new_n371_), .Y(new_new_n372_));
  AOI210     g350(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n209_), .Y(new_new_n373_));
  AOI210     g351(.A0(new_new_n373_), .A1(new_new_n372_), .B0(new_new_n368_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n141_), .B(new_new_n111_), .Y(new_new_n375_));
  OAI210     g353(.A0(new_new_n375_), .A1(new_new_n358_), .B0(i_2_), .Y(new_new_n376_));
  INV        g354(.A(new_new_n137_), .Y(new_new_n377_));
  NO3        g355(.A(new_new_n279_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n378_));
  AOI210     g356(.A0(new_new_n377_), .A1(new_new_n80_), .B0(new_new_n378_), .Y(new_new_n379_));
  AOI210     g357(.A0(new_new_n379_), .A1(new_new_n376_), .B0(new_new_n142_), .Y(new_new_n380_));
  OA210      g358(.A0(new_new_n280_), .A1(new_new_n112_), .B0(i_13_), .Y(new_new_n381_));
  AOI210     g359(.A0(new_new_n147_), .A1(new_new_n127_), .B0(new_new_n245_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n382_), .B(new_new_n211_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n94_), .B(new_new_n44_), .Y(new_new_n384_));
  INV        g362(.A(new_new_n178_), .Y(new_new_n385_));
  NA4        g363(.A(new_new_n385_), .B(new_new_n179_), .C(new_new_n110_), .D(new_new_n42_), .Y(new_new_n386_));
  OAI210     g364(.A0(new_new_n386_), .A1(new_new_n384_), .B0(new_new_n383_), .Y(new_new_n387_));
  NO3        g365(.A(new_new_n387_), .B(new_new_n381_), .C(new_new_n380_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n255_), .B(new_new_n28_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n357_), .B(new_new_n176_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n55_), .B(i_12_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n392_), .B(new_new_n112_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n393_), .B(new_new_n260_), .Y(new_new_n394_));
  AOI220     g372(.A0(new_new_n394_), .A1(new_new_n36_), .B0(new_new_n391_), .B1(new_new_n46_), .Y(new_new_n395_));
  NA4        g373(.A(new_new_n395_), .B(new_new_n388_), .C(new_new_n374_), .D(new_new_n364_), .Y(ori6));
  INV        g374(.A(new_new_n184_), .Y(new_new_n397_));
  OR2        g375(.A(new_new_n397_), .B(i_12_), .Y(new_new_n398_));
  NA2        g376(.A(new_new_n256_), .B(new_new_n56_), .Y(new_new_n399_));
  INV        g377(.A(new_new_n399_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n400_), .B(new_new_n66_), .Y(new_new_n401_));
  INV        g379(.A(new_new_n183_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n68_), .B(new_new_n117_), .Y(new_new_n403_));
  INV        g381(.A(new_new_n110_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n404_), .B(new_new_n46_), .Y(new_new_n405_));
  AOI210     g383(.A0(new_new_n405_), .A1(new_new_n403_), .B0(new_new_n402_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n162_), .B(i_9_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n407_), .B(new_new_n392_), .Y(new_new_n408_));
  AOI210     g386(.A0(new_new_n408_), .A1(new_new_n243_), .B0(new_new_n139_), .Y(new_new_n409_));
  NAi32      g387(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n335_), .B(new_new_n410_), .Y(new_new_n411_));
  OR3        g389(.A(new_new_n411_), .B(new_new_n409_), .C(new_new_n406_), .Y(new_new_n412_));
  BUFFER     g390(.A(new_new_n280_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n413_), .B(new_new_n126_), .Y(new_new_n414_));
  AO210      g392(.A0(new_new_n240_), .A1(new_new_n361_), .B0(new_new_n36_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(new_new_n414_), .Y(new_new_n416_));
  NO2        g394(.A(i_6_), .B(i_11_), .Y(new_new_n417_));
  NA2        g395(.A(new_new_n417_), .B(new_new_n251_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n205_), .B(new_new_n63_), .Y(new_new_n419_));
  NA3        g397(.A(new_new_n419_), .B(new_new_n418_), .C(new_new_n266_), .Y(new_new_n420_));
  NA2        g398(.A(new_new_n216_), .B(new_new_n214_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n103_), .B(new_new_n206_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n422_), .B(new_new_n421_), .Y(new_new_n423_));
  NO4        g401(.A(new_new_n423_), .B(new_new_n420_), .C(new_new_n416_), .D(new_new_n412_), .Y(new_new_n424_));
  NA4        g402(.A(new_new_n424_), .B(new_new_n401_), .C(new_new_n398_), .D(new_new_n199_), .Y(ori3));
  NA2        g403(.A(i_12_), .B(i_10_), .Y(new_new_n426_));
  NO2        g404(.A(i_11_), .B(new_new_n154_), .Y(new_new_n427_));
  NA2        g405(.A(new_new_n266_), .B(new_new_n193_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n428_), .B(new_new_n40_), .Y(new_new_n429_));
  NOi21      g407(.An(new_new_n90_), .B(new_new_n370_), .Y(new_new_n430_));
  INV        g408(.A(new_new_n430_), .Y(new_new_n431_));
  AOI210     g409(.A0(new_new_n431_), .A1(new_new_n429_), .B0(new_new_n47_), .Y(new_new_n432_));
  NO4        g410(.A(new_new_n196_), .B(new_new_n201_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n139_), .B(i_10_), .Y(new_new_n434_));
  NOi21      g412(.An(new_new_n434_), .B(new_new_n433_), .Y(new_new_n435_));
  NO2        g413(.A(new_new_n435_), .B(new_new_n56_), .Y(new_new_n436_));
  NOi21      g414(.An(i_5_), .B(i_9_), .Y(new_new_n437_));
  NA2        g415(.A(new_new_n437_), .B(new_new_n213_), .Y(new_new_n438_));
  BUFFER     g416(.A(new_new_n173_), .Y(new_new_n439_));
  NA2        g417(.A(new_new_n439_), .B(new_new_n230_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n440_), .B(new_new_n438_), .Y(new_new_n441_));
  NO3        g419(.A(new_new_n441_), .B(new_new_n436_), .C(new_new_n432_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n254_), .B(i_0_), .Y(new_new_n443_));
  NA2        g421(.A(new_new_n357_), .B(new_new_n184_), .Y(new_new_n444_));
  INV        g422(.A(new_new_n54_), .Y(new_new_n445_));
  NO2        g423(.A(new_new_n445_), .B(new_new_n444_), .Y(new_new_n446_));
  NO2        g424(.A(new_new_n164_), .B(new_new_n129_), .Y(new_new_n447_));
  NA2        g425(.A(i_0_), .B(i_10_), .Y(new_new_n448_));
  AN2        g426(.A(new_new_n447_), .B(i_6_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n449_), .B(new_new_n446_), .Y(new_new_n450_));
  INV        g428(.A(new_new_n450_), .Y(new_new_n451_));
  NA2        g429(.A(i_11_), .B(i_9_), .Y(new_new_n452_));
  NO3        g430(.A(i_12_), .B(new_new_n452_), .C(new_new_n265_), .Y(new_new_n453_));
  AN2        g431(.A(new_new_n453_), .B(i_5_), .Y(new_new_n454_));
  NA2        g432(.A(new_new_n204_), .B(new_new_n138_), .Y(new_new_n455_));
  NA2        g433(.A(new_new_n455_), .B(new_new_n133_), .Y(new_new_n456_));
  NO2        g434(.A(new_new_n452_), .B(new_new_n66_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n456_), .B(new_new_n454_), .Y(new_new_n458_));
  NA2        g436(.A(new_new_n298_), .B(new_new_n107_), .Y(new_new_n459_));
  NO2        g437(.A(i_6_), .B(new_new_n459_), .Y(new_new_n460_));
  NA2        g438(.A(new_new_n136_), .B(new_new_n95_), .Y(new_new_n461_));
  INV        g439(.A(new_new_n460_), .Y(new_new_n462_));
  NA2        g440(.A(new_new_n462_), .B(new_new_n458_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n426_), .B(new_new_n182_), .Y(new_new_n464_));
  NA2        g442(.A(new_new_n464_), .B(new_new_n457_), .Y(new_new_n465_));
  NA2        g443(.A(new_new_n244_), .B(new_new_n465_), .Y(new_new_n466_));
  NO3        g444(.A(new_new_n466_), .B(new_new_n463_), .C(new_new_n451_), .Y(new_new_n467_));
  NO2        g445(.A(new_new_n399_), .B(new_new_n461_), .Y(new_new_n468_));
  INV        g446(.A(new_new_n468_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n159_), .B(new_new_n152_), .Y(new_new_n470_));
  AOI210     g448(.A0(new_new_n470_), .A1(new_new_n443_), .B0(new_new_n129_), .Y(new_new_n471_));
  INV        g449(.A(new_new_n471_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n472_), .B(new_new_n469_), .Y(new_new_n473_));
  NO3        g451(.A(new_new_n448_), .B(new_new_n437_), .C(new_new_n141_), .Y(new_new_n474_));
  AOI220     g452(.A0(new_new_n474_), .A1(i_11_), .B0(new_new_n253_), .B1(new_new_n68_), .Y(new_new_n475_));
  NO3        g453(.A(new_new_n148_), .B(new_new_n201_), .C(i_0_), .Y(new_new_n476_));
  OAI210     g454(.A0(new_new_n476_), .A1(new_new_n69_), .B0(i_13_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n477_), .B(new_new_n475_), .Y(new_new_n478_));
  NA2        g456(.A(new_new_n239_), .B(new_new_n232_), .Y(new_new_n479_));
  INV        g457(.A(new_new_n479_), .Y(new_new_n480_));
  NA3        g458(.A(new_new_n203_), .B(new_new_n136_), .C(new_new_n135_), .Y(new_new_n481_));
  INV        g459(.A(new_new_n481_), .Y(new_new_n482_));
  NO3        g460(.A(new_new_n452_), .B(new_new_n149_), .C(new_new_n141_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n482_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n484_), .B(new_new_n480_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n79_), .B(i_5_), .Y(new_new_n486_));
  NA3        g464(.A(new_new_n427_), .B(new_new_n101_), .C(new_new_n110_), .Y(new_new_n487_));
  INV        g465(.A(new_new_n487_), .Y(new_new_n488_));
  NA2        g466(.A(new_new_n488_), .B(new_new_n486_), .Y(new_new_n489_));
  NAi21      g467(.An(new_new_n157_), .B(new_new_n158_), .Y(new_new_n490_));
  NO4        g468(.A(new_new_n156_), .B(new_new_n148_), .C(i_0_), .D(i_12_), .Y(new_new_n491_));
  NA2        g469(.A(new_new_n491_), .B(new_new_n490_), .Y(new_new_n492_));
  NA2        g470(.A(new_new_n492_), .B(new_new_n489_), .Y(new_new_n493_));
  NO4        g471(.A(new_new_n493_), .B(new_new_n485_), .C(new_new_n478_), .D(new_new_n473_), .Y(new_new_n494_));
  INV        g472(.A(new_new_n273_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n495_), .B(new_new_n146_), .Y(new_new_n496_));
  NO2        g474(.A(new_new_n496_), .B(new_new_n66_), .Y(new_new_n497_));
  INV        g475(.A(new_new_n198_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(new_new_n365_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n499_), .B(new_new_n497_), .Y(new_new_n500_));
  NA4        g478(.A(new_new_n500_), .B(new_new_n494_), .C(new_new_n467_), .D(new_new_n442_), .Y(ori4));
  INV        g479(.A(i_6_), .Y(new_new_n504_));
endmodule


