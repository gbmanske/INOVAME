library verilog;
use verilog.vl_types.all;
entity tb_average_comparator is
end tb_average_comparator;
