//Benchmark atmr_9sym_175_0.125

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n124_, mai_mai_n125_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, ori00, mai00, men00;
  INV        o00(.A(i_3_), .Y(ori_ori_n11_));
  INV        o01(.A(i_5_), .Y(ori_ori_n12_));
  NOi21      o02(.An(i_3_), .B(i_7_), .Y(ori_ori_n13_));
  INV        o03(.A(i_0_), .Y(ori_ori_n14_));
  NOi21      o04(.An(i_1_), .B(i_3_), .Y(ori_ori_n15_));
  INV        o05(.A(i_4_), .Y(ori_ori_n16_));
  INV        o06(.A(i_7_), .Y(ori_ori_n17_));
  NA3        o07(.A(i_6_), .B(i_5_), .C(ori_ori_n17_), .Y(ori_ori_n18_));
  INV        o08(.A(ori_ori_n18_), .Y(ori_ori_n19_));
  NA2        o09(.A(ori_ori_n19_), .B(ori_ori_n11_), .Y(ori_ori_n20_));
  NA2        o10(.A(ori_ori_n14_), .B(i_5_), .Y(ori_ori_n21_));
  INV        o11(.A(i_2_), .Y(ori_ori_n22_));
  NOi21      o12(.An(i_5_), .B(i_0_), .Y(ori_ori_n23_));
  NOi21      o13(.An(i_6_), .B(i_8_), .Y(ori_ori_n24_));
  NOi21      o14(.An(i_7_), .B(i_1_), .Y(ori_ori_n25_));
  NOi21      o15(.An(i_5_), .B(i_6_), .Y(ori_ori_n26_));
  AOI220     o16(.A0(ori_ori_n26_), .A1(ori_ori_n25_), .B0(ori_ori_n24_), .B1(ori_ori_n23_), .Y(ori_ori_n27_));
  NO3        o17(.A(ori_ori_n27_), .B(ori_ori_n22_), .C(i_4_), .Y(ori_ori_n28_));
  NOi21      o18(.An(i_0_), .B(i_4_), .Y(ori_ori_n29_));
  NOi21      o19(.An(i_7_), .B(i_5_), .Y(ori_ori_n30_));
  INV        o20(.A(i_1_), .Y(ori_ori_n31_));
  INV        o21(.A(ori_ori_n28_), .Y(ori_ori_n32_));
  NA2        o22(.A(i_1_), .B(ori_ori_n12_), .Y(ori_ori_n33_));
  NOi21      o23(.An(i_2_), .B(i_8_), .Y(ori_ori_n34_));
  NO2        o24(.A(ori_ori_n34_), .B(ori_ori_n29_), .Y(ori_ori_n35_));
  NO2        o25(.A(ori_ori_n35_), .B(ori_ori_n33_), .Y(ori_ori_n36_));
  INV        o26(.A(ori_ori_n36_), .Y(ori_ori_n37_));
  NOi21      o27(.An(i_4_), .B(i_3_), .Y(ori_ori_n38_));
  NOi21      o28(.An(i_1_), .B(i_4_), .Y(ori_ori_n39_));
  AN2        o29(.A(i_8_), .B(i_7_), .Y(ori_ori_n40_));
  NOi21      o30(.An(i_8_), .B(i_7_), .Y(ori_ori_n41_));
  NA2        o31(.A(ori_ori_n38_), .B(i_6_), .Y(ori_ori_n42_));
  INV        o32(.A(ori_ori_n42_), .Y(ori_ori_n43_));
  AOI220     o33(.A0(ori_ori_n43_), .A1(ori_ori_n22_), .B0(ori_ori_n38_), .B1(ori_ori_n26_), .Y(ori_ori_n44_));
  NA4        o34(.A(ori_ori_n44_), .B(ori_ori_n37_), .C(ori_ori_n32_), .D(ori_ori_n20_), .Y(ori_ori_n45_));
  NA2        o35(.A(i_8_), .B(ori_ori_n17_), .Y(ori_ori_n46_));
  AOI210     o36(.A0(i_3_), .A1(i_1_), .B0(i_2_), .Y(ori_ori_n47_));
  NOi21      o37(.An(i_1_), .B(i_2_), .Y(ori_ori_n48_));
  NO2        o38(.A(ori_ori_n47_), .B(ori_ori_n46_), .Y(ori_ori_n49_));
  NA2        o39(.A(ori_ori_n49_), .B(ori_ori_n12_), .Y(ori_ori_n50_));
  NA2        o40(.A(ori_ori_n41_), .B(i_2_), .Y(ori_ori_n51_));
  NOi32      o41(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n52_));
  INV        o42(.A(i_0_), .Y(ori_ori_n53_));
  NA2        o43(.A(ori_ori_n53_), .B(ori_ori_n52_), .Y(ori_ori_n54_));
  NA2        o44(.A(ori_ori_n54_), .B(ori_ori_n50_), .Y(ori_ori_n55_));
  NA2        o45(.A(ori_ori_n24_), .B(ori_ori_n23_), .Y(ori_ori_n56_));
  NOi21      o46(.An(i_7_), .B(i_8_), .Y(ori_ori_n57_));
  INV        o47(.A(ori_ori_n56_), .Y(ori_ori_n58_));
  NA2        o48(.A(ori_ori_n58_), .B(ori_ori_n48_), .Y(ori_ori_n59_));
  NA2        o49(.A(ori_ori_n15_), .B(ori_ori_n22_), .Y(ori_ori_n60_));
  NA3        o50(.A(ori_ori_n16_), .B(i_5_), .C(i_7_), .Y(ori_ori_n61_));
  NO2        o51(.A(ori_ori_n61_), .B(ori_ori_n60_), .Y(ori_ori_n62_));
  INV        o52(.A(ori_ori_n62_), .Y(ori_ori_n63_));
  NA3        o53(.A(ori_ori_n41_), .B(ori_ori_n22_), .C(i_3_), .Y(ori_ori_n64_));
  NA2        o54(.A(ori_ori_n31_), .B(i_6_), .Y(ori_ori_n65_));
  NO2        o55(.A(ori_ori_n65_), .B(ori_ori_n64_), .Y(ori_ori_n66_));
  NAi21      o56(.An(i_6_), .B(i_0_), .Y(ori_ori_n67_));
  NA2        o57(.A(ori_ori_n39_), .B(i_5_), .Y(ori_ori_n68_));
  NOi21      o58(.An(i_4_), .B(i_6_), .Y(ori_ori_n69_));
  NA2        o59(.A(ori_ori_n48_), .B(ori_ori_n69_), .Y(ori_ori_n70_));
  OAI210     o60(.A0(ori_ori_n68_), .A1(ori_ori_n67_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  NA2        o61(.A(ori_ori_n48_), .B(ori_ori_n24_), .Y(ori_ori_n72_));
  NOi21      o62(.An(ori_ori_n30_), .B(ori_ori_n72_), .Y(ori_ori_n73_));
  NO3        o63(.A(ori_ori_n73_), .B(ori_ori_n71_), .C(ori_ori_n66_), .Y(ori_ori_n74_));
  NOi21      o64(.An(i_3_), .B(i_1_), .Y(ori_ori_n75_));
  NA2        o65(.A(ori_ori_n75_), .B(i_4_), .Y(ori_ori_n76_));
  AOI210     o66(.A0(i_8_), .A1(i_6_), .B0(ori_ori_n76_), .Y(ori_ori_n77_));
  INV        o67(.A(ori_ori_n77_), .Y(ori_ori_n78_));
  NA4        o68(.A(ori_ori_n78_), .B(ori_ori_n74_), .C(ori_ori_n63_), .D(ori_ori_n59_), .Y(ori_ori_n79_));
  NA2        o69(.A(ori_ori_n34_), .B(ori_ori_n13_), .Y(ori_ori_n80_));
  NA2        o70(.A(ori_ori_n80_), .B(ori_ori_n72_), .Y(ori_ori_n81_));
  NA2        o71(.A(ori_ori_n81_), .B(ori_ori_n29_), .Y(ori_ori_n82_));
  INV        o72(.A(ori_ori_n38_), .Y(ori_ori_n83_));
  AOI210     o73(.A0(ori_ori_n83_), .A1(ori_ori_n51_), .B0(ori_ori_n21_), .Y(ori_ori_n84_));
  NOi21      o74(.An(i_0_), .B(i_2_), .Y(ori_ori_n85_));
  NA2        o75(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n86_));
  INV        o76(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  NA3        o77(.A(ori_ori_n39_), .B(ori_ori_n26_), .C(i_8_), .Y(ori_ori_n88_));
  INV        o78(.A(ori_ori_n88_), .Y(ori_ori_n89_));
  NO3        o79(.A(ori_ori_n89_), .B(ori_ori_n87_), .C(ori_ori_n84_), .Y(ori_ori_n90_));
  INV        o80(.A(ori_ori_n57_), .Y(ori_ori_n91_));
  AOI210     o81(.A0(ori_ori_n91_), .A1(ori_ori_n80_), .B0(ori_ori_n65_), .Y(ori_ori_n92_));
  NA2        o82(.A(ori_ori_n75_), .B(i_0_), .Y(ori_ori_n93_));
  NO2        o83(.A(ori_ori_n93_), .B(i_4_), .Y(ori_ori_n94_));
  NO2        o84(.A(ori_ori_n94_), .B(ori_ori_n92_), .Y(ori_ori_n95_));
  NO2        o85(.A(ori_ori_n64_), .B(ori_ori_n21_), .Y(ori_ori_n96_));
  NA3        o86(.A(ori_ori_n40_), .B(ori_ori_n31_), .C(ori_ori_n16_), .Y(ori_ori_n97_));
  NA3        o87(.A(ori_ori_n34_), .B(ori_ori_n23_), .C(ori_ori_n13_), .Y(ori_ori_n98_));
  NA2        o88(.A(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  NO2        o89(.A(ori_ori_n99_), .B(ori_ori_n96_), .Y(ori_ori_n100_));
  NA4        o90(.A(ori_ori_n100_), .B(ori_ori_n95_), .C(ori_ori_n90_), .D(ori_ori_n82_), .Y(ori_ori_n101_));
  OR4        o91(.A(ori_ori_n101_), .B(ori_ori_n79_), .C(ori_ori_n55_), .D(ori_ori_n45_), .Y(ori00));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NA3        m007(.A(i_1_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n18_));
  AOI210     m008(.A0(mai_mai_n18_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n19_));
  INV        m009(.A(i_4_), .Y(mai_mai_n20_));
  NA2        m010(.A(i_0_), .B(mai_mai_n20_), .Y(mai_mai_n21_));
  INV        m011(.A(i_7_), .Y(mai_mai_n22_));
  NOi21      m012(.An(i_8_), .B(i_6_), .Y(mai_mai_n23_));
  NO2        m013(.A(mai_mai_n124_), .B(mai_mai_n21_), .Y(mai_mai_n24_));
  AOI210     m014(.A0(mai_mai_n24_), .A1(mai_mai_n11_), .B0(mai_mai_n19_), .Y(mai_mai_n25_));
  NA2        m015(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n26_));
  INV        m016(.A(i_2_), .Y(mai_mai_n27_));
  NOi21      m017(.An(i_6_), .B(i_8_), .Y(mai_mai_n28_));
  NOi21      m018(.An(i_7_), .B(i_1_), .Y(mai_mai_n29_));
  NOi21      m019(.An(i_5_), .B(i_6_), .Y(mai_mai_n30_));
  AOI220     m020(.A0(mai_mai_n30_), .A1(mai_mai_n29_), .B0(mai_mai_n28_), .B1(i_5_), .Y(mai_mai_n31_));
  NO3        m021(.A(mai_mai_n31_), .B(mai_mai_n27_), .C(i_4_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_0_), .B(i_4_), .Y(mai_mai_n33_));
  XO2        m023(.A(i_1_), .B(i_3_), .Y(mai_mai_n34_));
  NOi21      m024(.An(i_3_), .B(i_0_), .Y(mai_mai_n35_));
  INV        m025(.A(mai_mai_n32_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_4_), .B(i_0_), .Y(mai_mai_n37_));
  INV        m027(.A(mai_mai_n15_), .Y(mai_mai_n38_));
  NA2        m028(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n39_));
  NOi21      m029(.An(i_2_), .B(i_8_), .Y(mai_mai_n40_));
  NO2        m030(.A(mai_mai_n40_), .B(mai_mai_n33_), .Y(mai_mai_n41_));
  NO3        m031(.A(mai_mai_n41_), .B(mai_mai_n39_), .C(mai_mai_n38_), .Y(mai_mai_n42_));
  INV        m032(.A(mai_mai_n42_), .Y(mai_mai_n43_));
  NOi31      m033(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n44_));
  NA2        m034(.A(mai_mai_n44_), .B(i_0_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_4_), .B(i_3_), .Y(mai_mai_n46_));
  NOi21      m036(.An(i_1_), .B(i_4_), .Y(mai_mai_n47_));
  OAI210     m037(.A0(mai_mai_n47_), .A1(mai_mai_n46_), .B0(mai_mai_n40_), .Y(mai_mai_n48_));
  NA2        m038(.A(mai_mai_n48_), .B(mai_mai_n45_), .Y(mai_mai_n49_));
  AN2        m039(.A(i_8_), .B(i_7_), .Y(mai_mai_n50_));
  INV        m040(.A(mai_mai_n50_), .Y(mai_mai_n51_));
  NOi21      m041(.An(i_8_), .B(i_7_), .Y(mai_mai_n52_));
  NA3        m042(.A(mai_mai_n52_), .B(mai_mai_n46_), .C(i_6_), .Y(mai_mai_n53_));
  OAI210     m043(.A0(mai_mai_n51_), .A1(mai_mai_n39_), .B0(mai_mai_n53_), .Y(mai_mai_n54_));
  AOI220     m044(.A0(mai_mai_n54_), .A1(mai_mai_n27_), .B0(mai_mai_n49_), .B1(mai_mai_n30_), .Y(mai_mai_n55_));
  NA4        m045(.A(mai_mai_n55_), .B(mai_mai_n43_), .C(mai_mai_n36_), .D(mai_mai_n25_), .Y(mai_mai_n56_));
  NA2        m046(.A(mai_mai_n34_), .B(i_2_), .Y(mai_mai_n57_));
  NOi21      m047(.An(i_1_), .B(i_2_), .Y(mai_mai_n58_));
  NO2        m048(.A(mai_mai_n57_), .B(mai_mai_n125_), .Y(mai_mai_n59_));
  NA2        m049(.A(mai_mai_n59_), .B(mai_mai_n14_), .Y(mai_mai_n60_));
  NA3        m050(.A(mai_mai_n52_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n61_));
  NA2        m051(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n62_));
  NA2        m052(.A(mai_mai_n62_), .B(mai_mai_n61_), .Y(mai_mai_n63_));
  NA2        m053(.A(i_8_), .B(i_3_), .Y(mai_mai_n64_));
  NA2        m054(.A(i_1_), .B(i_6_), .Y(mai_mai_n65_));
  NA2        m055(.A(mai_mai_n65_), .B(mai_mai_n64_), .Y(mai_mai_n66_));
  NO2        m056(.A(i_0_), .B(i_4_), .Y(mai_mai_n67_));
  AOI220     m057(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n63_), .B1(mai_mai_n46_), .Y(mai_mai_n68_));
  NA2        m058(.A(mai_mai_n68_), .B(mai_mai_n60_), .Y(mai_mai_n69_));
  NAi21      m059(.An(i_3_), .B(i_6_), .Y(mai_mai_n70_));
  NO2        m060(.A(mai_mai_n70_), .B(i_0_), .Y(mai_mai_n71_));
  NOi21      m061(.An(i_7_), .B(i_8_), .Y(mai_mai_n72_));
  NOi21      m062(.An(i_6_), .B(i_5_), .Y(mai_mai_n73_));
  AOI210     m063(.A0(mai_mai_n72_), .A1(mai_mai_n12_), .B0(mai_mai_n73_), .Y(mai_mai_n74_));
  NO2        m064(.A(mai_mai_n74_), .B(mai_mai_n11_), .Y(mai_mai_n75_));
  OAI210     m065(.A0(mai_mai_n75_), .A1(mai_mai_n71_), .B0(mai_mai_n58_), .Y(mai_mai_n76_));
  NA3        m066(.A(mai_mai_n20_), .B(i_5_), .C(i_7_), .Y(mai_mai_n77_));
  NO2        m067(.A(mai_mai_n77_), .B(i_2_), .Y(mai_mai_n78_));
  INV        m068(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  NA3        m069(.A(mai_mai_n52_), .B(mai_mai_n27_), .C(i_3_), .Y(mai_mai_n80_));
  INV        m070(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NOi21      m071(.An(i_2_), .B(i_1_), .Y(mai_mai_n82_));
  AN3        m072(.A(mai_mai_n72_), .B(mai_mai_n82_), .C(mai_mai_n37_), .Y(mai_mai_n83_));
  NAi21      m073(.An(i_6_), .B(i_0_), .Y(mai_mai_n84_));
  NOi21      m074(.An(i_4_), .B(i_6_), .Y(mai_mai_n85_));
  NOi21      m075(.An(i_5_), .B(i_3_), .Y(mai_mai_n86_));
  NA3        m076(.A(mai_mai_n86_), .B(mai_mai_n58_), .C(mai_mai_n85_), .Y(mai_mai_n87_));
  INV        m077(.A(mai_mai_n87_), .Y(mai_mai_n88_));
  NO3        m078(.A(mai_mai_n88_), .B(mai_mai_n83_), .C(mai_mai_n81_), .Y(mai_mai_n89_));
  NOi21      m079(.An(i_6_), .B(i_1_), .Y(mai_mai_n90_));
  AOI220     m080(.A0(mai_mai_n90_), .A1(i_7_), .B0(mai_mai_n23_), .B1(i_5_), .Y(mai_mai_n91_));
  NOi31      m081(.An(mai_mai_n37_), .B(mai_mai_n91_), .C(i_2_), .Y(mai_mai_n92_));
  NA2        m082(.A(mai_mai_n28_), .B(mai_mai_n14_), .Y(mai_mai_n93_));
  NOi21      m083(.An(i_3_), .B(i_1_), .Y(mai_mai_n94_));
  NA2        m084(.A(mai_mai_n94_), .B(i_4_), .Y(mai_mai_n95_));
  NO2        m085(.A(mai_mai_n93_), .B(mai_mai_n95_), .Y(mai_mai_n96_));
  NA2        m086(.A(mai_mai_n72_), .B(mai_mai_n14_), .Y(mai_mai_n97_));
  NOi31      m087(.An(mai_mai_n35_), .B(mai_mai_n97_), .C(mai_mai_n27_), .Y(mai_mai_n98_));
  NO3        m088(.A(mai_mai_n98_), .B(mai_mai_n96_), .C(mai_mai_n92_), .Y(mai_mai_n99_));
  NA4        m089(.A(mai_mai_n99_), .B(mai_mai_n89_), .C(mai_mai_n79_), .D(mai_mai_n76_), .Y(mai_mai_n100_));
  NA2        m090(.A(mai_mai_n28_), .B(mai_mai_n33_), .Y(mai_mai_n101_));
  NA2        m091(.A(mai_mai_n46_), .B(mai_mai_n29_), .Y(mai_mai_n102_));
  AOI210     m092(.A0(mai_mai_n102_), .A1(mai_mai_n61_), .B0(mai_mai_n26_), .Y(mai_mai_n103_));
  NAi31      m093(.An(mai_mai_n84_), .B(mai_mai_n72_), .C(mai_mai_n82_), .Y(mai_mai_n104_));
  NA3        m094(.A(mai_mai_n52_), .B(mai_mai_n44_), .C(i_6_), .Y(mai_mai_n105_));
  NA2        m095(.A(mai_mai_n105_), .B(mai_mai_n104_), .Y(mai_mai_n106_));
  NOi21      m096(.An(i_0_), .B(i_2_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n107_), .B(mai_mai_n29_), .C(mai_mai_n85_), .Y(mai_mai_n108_));
  NA3        m098(.A(mai_mai_n107_), .B(mai_mai_n46_), .C(mai_mai_n28_), .Y(mai_mai_n109_));
  NA2        m099(.A(mai_mai_n109_), .B(mai_mai_n108_), .Y(mai_mai_n110_));
  NO3        m100(.A(mai_mai_n110_), .B(mai_mai_n106_), .C(mai_mai_n103_), .Y(mai_mai_n111_));
  NO3        m101(.A(i_2_), .B(mai_mai_n11_), .C(mai_mai_n14_), .Y(mai_mai_n112_));
  NA2        m102(.A(i_2_), .B(i_4_), .Y(mai_mai_n113_));
  AOI210     m103(.A0(mai_mai_n84_), .A1(mai_mai_n70_), .B0(mai_mai_n113_), .Y(mai_mai_n114_));
  NO2        m104(.A(i_8_), .B(i_7_), .Y(mai_mai_n115_));
  OA210      m105(.A0(mai_mai_n114_), .A1(mai_mai_n112_), .B0(mai_mai_n115_), .Y(mai_mai_n116_));
  NA3        m106(.A(mai_mai_n94_), .B(i_5_), .C(mai_mai_n22_), .Y(mai_mai_n117_));
  INV        m107(.A(mai_mai_n117_), .Y(mai_mai_n118_));
  NO2        m108(.A(mai_mai_n118_), .B(mai_mai_n116_), .Y(mai_mai_n119_));
  NA3        m109(.A(mai_mai_n119_), .B(mai_mai_n111_), .C(mai_mai_n101_), .Y(mai_mai_n120_));
  OR4        m110(.A(mai_mai_n120_), .B(mai_mai_n100_), .C(mai_mai_n69_), .D(mai_mai_n56_), .Y(mai00));
  INV        m111(.A(i_8_), .Y(mai_mai_n124_));
  INV        m112(.A(i_8_), .Y(mai_mai_n125_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  INV        u005(.A(i_0_), .Y(men_men_n16_));
  NOi21      u006(.An(i_1_), .B(i_3_), .Y(men_men_n17_));
  INV        u007(.A(i_4_), .Y(men_men_n18_));
  INV        u008(.A(i_0_), .Y(men_men_n19_));
  INV        u009(.A(i_7_), .Y(men_men_n20_));
  NOi21      u010(.An(i_8_), .B(i_6_), .Y(men_men_n21_));
  NOi21      u011(.An(i_1_), .B(i_8_), .Y(men_men_n22_));
  NA2        u012(.A(men_men_n22_), .B(i_2_), .Y(men_men_n23_));
  NO2        u013(.A(men_men_n23_), .B(men_men_n19_), .Y(men_men_n24_));
  NA2        u014(.A(men_men_n24_), .B(men_men_n11_), .Y(men_men_n25_));
  NO2        u015(.A(i_2_), .B(i_4_), .Y(men_men_n26_));
  NA3        u016(.A(men_men_n26_), .B(i_6_), .C(i_8_), .Y(men_men_n27_));
  AOI210     u017(.A0(i_0_), .A1(i_5_), .B0(men_men_n27_), .Y(men_men_n28_));
  INV        u018(.A(i_2_), .Y(men_men_n29_));
  NOi21      u019(.An(i_6_), .B(i_8_), .Y(men_men_n30_));
  NOi21      u020(.An(i_5_), .B(i_6_), .Y(men_men_n31_));
  NOi21      u021(.An(i_0_), .B(i_4_), .Y(men_men_n32_));
  XO2        u022(.A(i_1_), .B(i_3_), .Y(men_men_n33_));
  NOi21      u023(.An(i_7_), .B(i_5_), .Y(men_men_n34_));
  AN3        u024(.A(men_men_n34_), .B(men_men_n33_), .C(men_men_n32_), .Y(men_men_n35_));
  INV        u025(.A(i_1_), .Y(men_men_n36_));
  NOi21      u026(.An(i_3_), .B(i_0_), .Y(men_men_n37_));
  NA2        u027(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  AOI210     u028(.A0(men_men_n123_), .A1(men_men_n125_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO3        u029(.A(men_men_n39_), .B(men_men_n35_), .C(men_men_n28_), .Y(men_men_n40_));
  NOi21      u030(.An(i_4_), .B(i_0_), .Y(men_men_n41_));
  INV        u031(.A(men_men_n15_), .Y(men_men_n42_));
  NA2        u032(.A(i_1_), .B(men_men_n14_), .Y(men_men_n43_));
  NO3        u033(.A(i_2_), .B(men_men_n43_), .C(men_men_n42_), .Y(men_men_n44_));
  INV        u034(.A(men_men_n44_), .Y(men_men_n45_));
  NOi31      u035(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n46_));
  NOi21      u036(.An(i_4_), .B(i_3_), .Y(men_men_n47_));
  NOi21      u037(.An(i_1_), .B(i_4_), .Y(men_men_n48_));
  NA2        u038(.A(i_8_), .B(men_men_n12_), .Y(men_men_n49_));
  NOi21      u039(.An(i_8_), .B(i_7_), .Y(men_men_n50_));
  NA3        u040(.A(men_men_n50_), .B(men_men_n47_), .C(i_6_), .Y(men_men_n51_));
  OAI210     u041(.A0(men_men_n49_), .A1(men_men_n43_), .B0(men_men_n51_), .Y(men_men_n52_));
  NA2        u042(.A(men_men_n52_), .B(men_men_n29_), .Y(men_men_n53_));
  NA4        u043(.A(men_men_n53_), .B(men_men_n45_), .C(men_men_n40_), .D(men_men_n25_), .Y(men_men_n54_));
  NA2        u044(.A(i_8_), .B(i_7_), .Y(men_men_n55_));
  NO3        u045(.A(men_men_n55_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n56_));
  NA2        u046(.A(i_8_), .B(men_men_n20_), .Y(men_men_n57_));
  AOI220     u047(.A0(men_men_n37_), .A1(i_1_), .B0(men_men_n33_), .B1(i_2_), .Y(men_men_n58_));
  NOi21      u048(.An(i_1_), .B(i_2_), .Y(men_men_n59_));
  NO2        u049(.A(men_men_n58_), .B(men_men_n57_), .Y(men_men_n60_));
  OAI210     u050(.A0(men_men_n60_), .A1(men_men_n56_), .B0(men_men_n14_), .Y(men_men_n61_));
  NOi32      u051(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n17_), .B(i_2_), .C(i_6_), .Y(men_men_n63_));
  INV        u053(.A(men_men_n63_), .Y(men_men_n64_));
  NO2        u054(.A(i_0_), .B(i_4_), .Y(men_men_n65_));
  NA2        u055(.A(men_men_n65_), .B(men_men_n64_), .Y(men_men_n66_));
  NA2        u056(.A(men_men_n66_), .B(men_men_n61_), .Y(men_men_n67_));
  NOi21      u057(.An(i_7_), .B(i_8_), .Y(men_men_n68_));
  NA2        u058(.A(men_men_n68_), .B(men_men_n59_), .Y(men_men_n69_));
  NA3        u059(.A(men_men_n21_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n70_));
  AOI210     u060(.A0(men_men_n19_), .A1(men_men_n124_), .B0(men_men_n70_), .Y(men_men_n71_));
  INV        u061(.A(i_5_), .Y(men_men_n72_));
  NA3        u062(.A(men_men_n55_), .B(men_men_n17_), .C(men_men_n16_), .Y(men_men_n73_));
  NO2        u063(.A(men_men_n73_), .B(men_men_n72_), .Y(men_men_n74_));
  NO2        u064(.A(men_men_n74_), .B(men_men_n71_), .Y(men_men_n75_));
  NA3        u065(.A(men_men_n48_), .B(i_5_), .C(men_men_n20_), .Y(men_men_n76_));
  NOi21      u066(.An(i_4_), .B(i_6_), .Y(men_men_n77_));
  NOi21      u067(.An(i_5_), .B(i_3_), .Y(men_men_n78_));
  NA3        u068(.A(men_men_n76_), .B(men_men_n75_), .C(men_men_n69_), .Y(men_men_n79_));
  NA2        u069(.A(i_2_), .B(men_men_n15_), .Y(men_men_n80_));
  NOi31      u070(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n81_));
  NOi31      u071(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n82_));
  OAI210     u072(.A0(men_men_n82_), .A1(men_men_n81_), .B0(i_7_), .Y(men_men_n83_));
  NA3        u073(.A(men_men_n30_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n84_));
  NA3        u074(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n80_), .Y(men_men_n85_));
  NA2        u075(.A(men_men_n85_), .B(men_men_n32_), .Y(men_men_n86_));
  NA3        u076(.A(men_men_n50_), .B(men_men_n46_), .C(i_6_), .Y(men_men_n87_));
  INV        u077(.A(men_men_n87_), .Y(men_men_n88_));
  NA3        u078(.A(men_men_n41_), .B(men_men_n34_), .C(men_men_n17_), .Y(men_men_n89_));
  NOi32      u079(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n90_));
  NA2        u080(.A(men_men_n90_), .B(men_men_n81_), .Y(men_men_n91_));
  NA3        u081(.A(i_0_), .B(men_men_n47_), .C(men_men_n30_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n92_), .B(men_men_n91_), .C(men_men_n89_), .Y(men_men_n93_));
  NA3        u083(.A(men_men_n46_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n94_));
  NA4        u084(.A(men_men_n48_), .B(men_men_n31_), .C(men_men_n16_), .D(i_8_), .Y(men_men_n95_));
  NA2        u085(.A(men_men_n95_), .B(men_men_n94_), .Y(men_men_n96_));
  NO3        u086(.A(men_men_n96_), .B(men_men_n93_), .C(men_men_n88_), .Y(men_men_n97_));
  NOi21      u087(.An(i_5_), .B(i_2_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n98_), .B(men_men_n68_), .Y(men_men_n99_));
  NO2        u089(.A(men_men_n99_), .B(men_men_n126_), .Y(men_men_n100_));
  NO4        u090(.A(i_2_), .B(men_men_n18_), .C(men_men_n11_), .D(men_men_n14_), .Y(men_men_n101_));
  NA2        u091(.A(i_2_), .B(i_4_), .Y(men_men_n102_));
  INV        u092(.A(men_men_n102_), .Y(men_men_n103_));
  NO2        u093(.A(i_8_), .B(i_7_), .Y(men_men_n104_));
  OA210      u094(.A0(men_men_n103_), .A1(men_men_n101_), .B0(men_men_n104_), .Y(men_men_n105_));
  NA3        u095(.A(i_0_), .B(i_5_), .C(men_men_n20_), .Y(men_men_n106_));
  NO2        u096(.A(men_men_n106_), .B(i_4_), .Y(men_men_n107_));
  NO3        u097(.A(men_men_n107_), .B(men_men_n105_), .C(men_men_n100_), .Y(men_men_n108_));
  NA2        u098(.A(men_men_n68_), .B(men_men_n12_), .Y(men_men_n109_));
  NO2        u099(.A(men_men_n122_), .B(men_men_n109_), .Y(men_men_n110_));
  NA2        u100(.A(men_men_n50_), .B(men_men_n77_), .Y(men_men_n111_));
  INV        u101(.A(men_men_n111_), .Y(men_men_n112_));
  NA3        u102(.A(men_men_n78_), .B(i_8_), .C(men_men_n36_), .Y(men_men_n113_));
  NOi31      u103(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n114_));
  OAI210     u104(.A0(men_men_n90_), .A1(men_men_n62_), .B0(men_men_n114_), .Y(men_men_n115_));
  NA2        u105(.A(men_men_n115_), .B(men_men_n113_), .Y(men_men_n116_));
  NO3        u106(.A(men_men_n116_), .B(men_men_n112_), .C(men_men_n110_), .Y(men_men_n117_));
  NA4        u107(.A(men_men_n117_), .B(men_men_n108_), .C(men_men_n97_), .D(men_men_n86_), .Y(men_men_n118_));
  OR4        u108(.A(men_men_n118_), .B(men_men_n79_), .C(men_men_n67_), .D(men_men_n54_), .Y(men00));
  INV        u109(.A(i_2_), .Y(men_men_n122_));
  INV        u110(.A(i_7_), .Y(men_men_n123_));
  INV        u111(.A(i_1_), .Y(men_men_n124_));
  INV        u112(.A(i_6_), .Y(men_men_n125_));
  INV        u113(.A(i_6_), .Y(men_men_n126_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule