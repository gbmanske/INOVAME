// Benchmark "top" written by ABC on Fri Jun 21 17:49:28 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n142_, new_new_n143_,
    new_new_n144_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n703_, new_new_n704_, new_new_n705_, new_new_n706_,
    new_new_n707_, new_new_n708_, new_new_n709_, new_new_n710_,
    new_new_n711_, new_new_n712_, new_new_n713_, new_new_n714_,
    new_new_n715_, new_new_n716_, new_new_n717_, new_new_n718_,
    new_new_n719_, new_new_n720_, new_new_n721_, new_new_n722_,
    new_new_n723_, new_new_n724_, new_new_n725_, new_new_n726_,
    new_new_n727_, new_new_n728_, new_new_n729_, new_new_n730_,
    new_new_n731_, new_new_n732_, new_new_n733_, new_new_n734_,
    new_new_n735_, new_new_n736_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n751_,
    new_new_n752_, new_new_n753_, new_new_n754_, new_new_n755_,
    new_new_n756_, new_new_n757_, new_new_n758_, new_new_n759_,
    new_new_n760_, new_new_n761_, new_new_n762_, new_new_n763_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_,
    new_new_n768_, new_new_n769_, new_new_n770_, new_new_n771_,
    new_new_n772_, new_new_n773_, new_new_n774_, new_new_n775_,
    new_new_n776_, new_new_n777_, new_new_n778_, new_new_n779_,
    new_new_n780_, new_new_n781_, new_new_n782_, new_new_n783_,
    new_new_n784_, new_new_n785_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g021(.A(new_new_n35_), .Y(mai1));
  INV        g022(.A(i_11_), .Y(new_new_n45_));
  NO2        g023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g024(.A(i_2_), .Y(new_new_n47_));
  NA2        g025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g026(.A(i_5_), .Y(new_new_n49_));
  NO2        g027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g041(.A(i_1_), .Y(new_new_n64_));
  NA2        g042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g064(.A(i_6_), .Y(new_new_n87_));
  OR4        g065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g082(.A(i_7_), .Y(new_new_n105_));
  NA2        g083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  AN2        g090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g092(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n115_));
  NO2        g093(.A(i_8_), .B(new_new_n105_), .Y(new_new_n116_));
  NO3        g094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_0_), .Y(new_new_n120_));
  NA2        g098(.A(i_11_), .B(i_12_), .Y(new_new_n121_));
  OAI210     g099(.A0(new_new_n120_), .A1(new_new_n118_), .B0(new_new_n121_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n122_), .B(new_new_n117_), .Y(new_new_n123_));
  NA3        g101(.A(new_new_n123_), .B(new_new_n111_), .C(new_new_n104_), .Y(new_new_n124_));
  NOi21      g102(.An(i_1_), .B(i_5_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(i_11_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g105(.A(i_7_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NO2        g107(.A(new_new_n129_), .B(new_new_n47_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n131_));
  NAi21      g109(.An(i_3_), .B(i_8_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n132_), .B(new_new_n63_), .Y(new_new_n133_));
  NOi31      g111(.An(new_new_n133_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n134_));
  NO2        g112(.A(i_1_), .B(new_new_n87_), .Y(new_new_n135_));
  NO2        g113(.A(i_6_), .B(i_5_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_3_), .Y(new_new_n137_));
  AO210      g115(.A0(new_new_n137_), .A1(new_new_n48_), .B0(new_new_n135_), .Y(new_new_n138_));
  OAI220     g116(.A0(new_new_n138_), .A1(new_new_n112_), .B0(new_new_n134_), .B1(new_new_n126_), .Y(new_new_n139_));
  NO3        g117(.A(new_new_n139_), .B(new_new_n124_), .C(new_new_n99_), .Y(new_new_n140_));
  NA3        g118(.A(new_new_n140_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g119(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n142_));
  INV        g120(.A(i_6_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NA4        g122(.A(new_new_n144_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g123(.A(i_8_), .B(i_7_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(i_6_), .Y(new_new_n147_));
  NO2        g125(.A(i_12_), .B(i_13_), .Y(new_new_n148_));
  NAi21      g126(.An(i_5_), .B(i_11_), .Y(new_new_n149_));
  NOi21      g127(.An(new_new_n148_), .B(new_new_n149_), .Y(new_new_n150_));
  NO2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NA2        g129(.A(i_2_), .B(i_3_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n152_), .B(i_4_), .Y(new_new_n153_));
  NA3        g131(.A(new_new_n153_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n154_));
  OR2        g132(.A(new_new_n154_), .B(new_new_n25_), .Y(new_new_n155_));
  AN2        g133(.A(new_new_n148_), .B(new_new_n84_), .Y(new_new_n156_));
  NA2        g134(.A(i_1_), .B(i_5_), .Y(new_new_n157_));
  OR2        g135(.A(i_0_), .B(i_1_), .Y(new_new_n158_));
  NAi32      g136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NOi21      g137(.An(i_4_), .B(i_10_), .Y(new_new_n160_));
  NA2        g138(.A(new_new_n160_), .B(new_new_n40_), .Y(new_new_n161_));
  NO2        g139(.A(i_3_), .B(i_5_), .Y(new_new_n162_));
  NO3        g140(.A(new_new_n74_), .B(i_2_), .C(i_1_), .Y(new_new_n163_));
  NA2        g141(.A(new_new_n163_), .B(new_new_n162_), .Y(new_new_n164_));
  NO2        g142(.A(new_new_n155_), .B(new_new_n147_), .Y(new_new_n165_));
  NA3        g143(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n166_));
  NA2        g144(.A(i_3_), .B(new_new_n49_), .Y(new_new_n167_));
  NOi21      g145(.An(i_4_), .B(i_9_), .Y(new_new_n168_));
  NOi21      g146(.An(i_11_), .B(i_13_), .Y(new_new_n169_));
  NA2        g147(.A(new_new_n169_), .B(new_new_n168_), .Y(new_new_n170_));
  OR2        g148(.A(new_new_n170_), .B(new_new_n167_), .Y(new_new_n171_));
  NO2        g149(.A(i_4_), .B(i_5_), .Y(new_new_n172_));
  NAi21      g150(.An(i_12_), .B(i_11_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n173_), .B(i_13_), .Y(new_new_n174_));
  NA3        g152(.A(new_new_n174_), .B(new_new_n172_), .C(new_new_n84_), .Y(new_new_n175_));
  AOI210     g153(.A0(new_new_n175_), .A1(new_new_n171_), .B0(new_new_n166_), .Y(new_new_n176_));
  NO2        g154(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n177_), .B(new_new_n47_), .Y(new_new_n178_));
  NA2        g156(.A(new_new_n36_), .B(i_5_), .Y(new_new_n179_));
  NA2        g157(.A(i_3_), .B(i_5_), .Y(new_new_n180_));
  NO2        g158(.A(new_new_n74_), .B(i_5_), .Y(new_new_n181_));
  NO2        g159(.A(i_2_), .B(i_1_), .Y(new_new_n182_));
  NA2        g160(.A(new_new_n182_), .B(i_3_), .Y(new_new_n183_));
  NAi21      g161(.An(i_4_), .B(i_12_), .Y(new_new_n184_));
  NO4        g162(.A(new_new_n184_), .B(new_new_n183_), .C(i_11_), .D(new_new_n25_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(new_new_n176_), .Y(new_new_n186_));
  INV        g164(.A(i_8_), .Y(new_new_n187_));
  NO2        g165(.A(new_new_n187_), .B(i_7_), .Y(new_new_n188_));
  NA2        g166(.A(new_new_n188_), .B(i_6_), .Y(new_new_n189_));
  NO3        g167(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n190_));
  NO3        g168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n191_));
  NO2        g169(.A(i_3_), .B(i_8_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n193_));
  NA3        g171(.A(new_new_n193_), .B(new_new_n192_), .C(new_new_n40_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n195_));
  INV        g173(.A(new_new_n195_), .Y(new_new_n196_));
  NO2        g174(.A(i_13_), .B(i_9_), .Y(new_new_n197_));
  NA3        g175(.A(new_new_n197_), .B(i_6_), .C(new_new_n187_), .Y(new_new_n198_));
  NAi21      g176(.An(i_12_), .B(i_3_), .Y(new_new_n199_));
  OR2        g177(.A(new_new_n199_), .B(new_new_n198_), .Y(new_new_n200_));
  NO2        g178(.A(new_new_n45_), .B(i_5_), .Y(new_new_n201_));
  NA3        g179(.A(i_1_), .B(new_new_n201_), .C(i_10_), .Y(new_new_n202_));
  OAI220     g180(.A0(new_new_n202_), .A1(new_new_n200_), .B0(new_new_n196_), .B1(new_new_n194_), .Y(new_new_n203_));
  NA2        g181(.A(new_new_n203_), .B(i_7_), .Y(new_new_n204_));
  OAI220     g182(.A0(new_new_n204_), .A1(i_4_), .B0(new_new_n189_), .B1(new_new_n186_), .Y(new_new_n205_));
  NAi21      g183(.An(i_12_), .B(i_7_), .Y(new_new_n206_));
  NA3        g184(.A(i_13_), .B(new_new_n187_), .C(i_10_), .Y(new_new_n207_));
  NO2        g185(.A(new_new_n207_), .B(new_new_n206_), .Y(new_new_n208_));
  NA2        g186(.A(i_0_), .B(i_5_), .Y(new_new_n209_));
  INV        g187(.A(new_new_n108_), .Y(new_new_n210_));
  OAI220     g188(.A0(new_new_n210_), .A1(new_new_n183_), .B0(new_new_n178_), .B1(new_new_n137_), .Y(new_new_n211_));
  NAi31      g189(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n212_));
  NO2        g190(.A(new_new_n36_), .B(i_13_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n214_));
  NO2        g192(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n215_));
  NA3        g193(.A(new_new_n215_), .B(new_new_n214_), .C(new_new_n213_), .Y(new_new_n216_));
  INV        g194(.A(i_13_), .Y(new_new_n217_));
  NO2        g195(.A(i_12_), .B(new_new_n217_), .Y(new_new_n218_));
  NA3        g196(.A(new_new_n218_), .B(new_new_n191_), .C(new_new_n190_), .Y(new_new_n219_));
  OAI210     g197(.A0(new_new_n216_), .A1(new_new_n212_), .B0(new_new_n219_), .Y(new_new_n220_));
  AOI220     g198(.A0(new_new_n220_), .A1(new_new_n146_), .B0(new_new_n211_), .B1(new_new_n208_), .Y(new_new_n221_));
  NO2        g199(.A(i_12_), .B(new_new_n37_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n180_), .B(i_4_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n223_), .B(new_new_n222_), .Y(new_new_n224_));
  OR2        g202(.A(i_8_), .B(i_7_), .Y(new_new_n225_));
  NO2        g203(.A(new_new_n225_), .B(new_new_n87_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n54_), .B(i_1_), .Y(new_new_n227_));
  INV        g205(.A(i_12_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n45_), .B(new_new_n228_), .Y(new_new_n229_));
  NO3        g207(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n230_));
  NA2        g208(.A(i_2_), .B(i_1_), .Y(new_new_n231_));
  NO3        g209(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n232_));
  NAi21      g210(.An(i_4_), .B(i_3_), .Y(new_new_n233_));
  NO2        g211(.A(i_0_), .B(i_6_), .Y(new_new_n234_));
  NOi41      g212(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n235_));
  NA2        g213(.A(new_new_n235_), .B(new_new_n234_), .Y(new_new_n236_));
  NO2        g214(.A(new_new_n231_), .B(new_new_n180_), .Y(new_new_n237_));
  NAi21      g215(.An(new_new_n236_), .B(new_new_n237_), .Y(new_new_n238_));
  INV        g216(.A(new_new_n238_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n239_), .B(new_new_n40_), .Y(new_new_n240_));
  NO2        g218(.A(i_11_), .B(new_new_n217_), .Y(new_new_n241_));
  NOi21      g219(.An(i_1_), .B(i_6_), .Y(new_new_n242_));
  NAi21      g220(.An(i_3_), .B(i_7_), .Y(new_new_n243_));
  NA2        g221(.A(new_new_n228_), .B(i_9_), .Y(new_new_n244_));
  OR4        g222(.A(new_new_n244_), .B(new_new_n243_), .C(new_new_n242_), .D(new_new_n181_), .Y(new_new_n245_));
  NO2        g223(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n74_), .B(i_5_), .Y(new_new_n247_));
  NA2        g225(.A(i_3_), .B(i_9_), .Y(new_new_n248_));
  NAi21      g226(.An(i_7_), .B(i_10_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n249_), .B(new_new_n248_), .Y(new_new_n250_));
  NA3        g228(.A(new_new_n250_), .B(new_new_n247_), .C(new_new_n65_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n251_), .B(new_new_n245_), .Y(new_new_n252_));
  NA3        g230(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n253_));
  INV        g231(.A(new_new_n147_), .Y(new_new_n254_));
  NA2        g232(.A(new_new_n228_), .B(i_13_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n255_), .B(new_new_n76_), .Y(new_new_n256_));
  AOI220     g234(.A0(new_new_n256_), .A1(new_new_n254_), .B0(new_new_n252_), .B1(new_new_n241_), .Y(new_new_n257_));
  NA2        g235(.A(i_12_), .B(i_6_), .Y(new_new_n258_));
  OR2        g236(.A(i_13_), .B(i_9_), .Y(new_new_n259_));
  NO2        g237(.A(new_new_n233_), .B(i_2_), .Y(new_new_n260_));
  NA2        g238(.A(new_new_n241_), .B(i_9_), .Y(new_new_n261_));
  NO3        g239(.A(i_11_), .B(new_new_n217_), .C(new_new_n25_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n243_), .B(i_8_), .Y(new_new_n263_));
  NO2        g241(.A(i_6_), .B(new_new_n49_), .Y(new_new_n264_));
  NA3        g242(.A(new_new_n257_), .B(new_new_n240_), .C(new_new_n221_), .Y(new_new_n265_));
  NO3        g243(.A(i_12_), .B(new_new_n217_), .C(new_new_n37_), .Y(new_new_n266_));
  INV        g244(.A(new_new_n266_), .Y(new_new_n267_));
  NA2        g245(.A(i_8_), .B(new_new_n105_), .Y(new_new_n268_));
  NOi21      g246(.An(new_new_n162_), .B(new_new_n87_), .Y(new_new_n269_));
  NO3        g247(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n270_));
  AOI220     g248(.A0(new_new_n270_), .A1(new_new_n190_), .B0(new_new_n269_), .B1(new_new_n227_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n271_), .B(new_new_n268_), .Y(new_new_n272_));
  NO3        g250(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n231_), .B(i_0_), .Y(new_new_n274_));
  AOI220     g252(.A0(new_new_n274_), .A1(new_new_n188_), .B0(new_new_n273_), .B1(new_new_n146_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n264_), .B(new_new_n26_), .Y(new_new_n276_));
  NO2        g254(.A(new_new_n276_), .B(new_new_n275_), .Y(new_new_n277_));
  NA2        g255(.A(i_0_), .B(i_1_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n278_), .B(i_2_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n60_), .B(i_6_), .Y(new_new_n280_));
  NA3        g258(.A(new_new_n280_), .B(new_new_n279_), .C(new_new_n162_), .Y(new_new_n281_));
  OAI210     g259(.A0(new_new_n164_), .A1(new_new_n147_), .B0(new_new_n281_), .Y(new_new_n282_));
  NO3        g260(.A(new_new_n282_), .B(new_new_n277_), .C(new_new_n272_), .Y(new_new_n283_));
  NO2        g261(.A(i_3_), .B(i_10_), .Y(new_new_n284_));
  NA3        g262(.A(new_new_n284_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n285_));
  NO2        g263(.A(i_2_), .B(new_new_n105_), .Y(new_new_n286_));
  NOi21      g264(.An(new_new_n209_), .B(new_new_n107_), .Y(new_new_n287_));
  NA3        g265(.A(new_new_n287_), .B(i_1_), .C(new_new_n286_), .Y(new_new_n288_));
  AN2        g266(.A(i_3_), .B(i_10_), .Y(new_new_n289_));
  NA4        g267(.A(new_new_n289_), .B(new_new_n191_), .C(new_new_n174_), .D(new_new_n172_), .Y(new_new_n290_));
  NO2        g268(.A(i_5_), .B(new_new_n37_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n292_));
  OR2        g270(.A(new_new_n288_), .B(new_new_n285_), .Y(new_new_n293_));
  OAI220     g271(.A0(new_new_n293_), .A1(i_6_), .B0(new_new_n283_), .B1(new_new_n267_), .Y(new_new_n294_));
  NO4        g272(.A(new_new_n294_), .B(new_new_n265_), .C(new_new_n205_), .D(new_new_n165_), .Y(new_new_n295_));
  NO3        g273(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n274_), .B(new_new_n297_), .Y(new_new_n298_));
  NO3        g276(.A(i_6_), .B(new_new_n187_), .C(i_7_), .Y(new_new_n299_));
  NO2        g277(.A(new_new_n298_), .B(new_new_n167_), .Y(new_new_n300_));
  NO2        g278(.A(i_2_), .B(i_3_), .Y(new_new_n301_));
  OR2        g279(.A(i_0_), .B(i_5_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n209_), .B(new_new_n302_), .Y(new_new_n303_));
  NA4        g281(.A(new_new_n303_), .B(new_new_n226_), .C(new_new_n301_), .D(i_1_), .Y(new_new_n304_));
  NA3        g282(.A(new_new_n274_), .B(new_new_n269_), .C(new_new_n116_), .Y(new_new_n305_));
  NAi21      g283(.An(i_8_), .B(i_7_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(i_6_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n158_), .B(new_new_n47_), .Y(new_new_n308_));
  NA3        g286(.A(new_new_n308_), .B(new_new_n307_), .C(new_new_n162_), .Y(new_new_n309_));
  NA3        g287(.A(new_new_n309_), .B(new_new_n305_), .C(new_new_n304_), .Y(new_new_n310_));
  OAI210     g288(.A0(new_new_n310_), .A1(new_new_n300_), .B0(i_4_), .Y(new_new_n311_));
  NO2        g289(.A(i_12_), .B(i_10_), .Y(new_new_n312_));
  NOi21      g290(.An(i_5_), .B(i_0_), .Y(new_new_n313_));
  NA4        g291(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n314_));
  NO2        g292(.A(i_6_), .B(i_8_), .Y(new_new_n315_));
  NOi21      g293(.An(i_0_), .B(i_2_), .Y(new_new_n316_));
  AN2        g294(.A(new_new_n316_), .B(new_new_n315_), .Y(new_new_n317_));
  NO2        g295(.A(i_1_), .B(i_7_), .Y(new_new_n318_));
  AO220      g296(.A0(new_new_n318_), .A1(new_new_n317_), .B0(new_new_n307_), .B1(new_new_n227_), .Y(new_new_n319_));
  NA2        g297(.A(new_new_n319_), .B(new_new_n42_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n320_), .B(new_new_n311_), .Y(new_new_n321_));
  NA3        g299(.A(new_new_n242_), .B(new_new_n286_), .C(new_new_n187_), .Y(new_new_n322_));
  INV        g300(.A(new_new_n85_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n278_), .B(new_new_n82_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n324_), .B(new_new_n136_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n96_), .B(new_new_n187_), .Y(new_new_n326_));
  NA3        g304(.A(new_new_n287_), .B(new_new_n326_), .C(new_new_n64_), .Y(new_new_n327_));
  AOI210     g305(.A0(new_new_n327_), .A1(new_new_n325_), .B0(new_new_n323_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n187_), .B(i_9_), .Y(new_new_n329_));
  NA2        g307(.A(new_new_n329_), .B(new_new_n195_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n328_), .B(new_new_n277_), .Y(new_new_n331_));
  AOI210     g309(.A0(new_new_n331_), .A1(new_new_n322_), .B0(new_new_n161_), .Y(new_new_n332_));
  AOI210     g310(.A0(new_new_n321_), .A1(new_new_n296_), .B0(new_new_n332_), .Y(new_new_n333_));
  NOi32      g311(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n334_));
  INV        g312(.A(new_new_n334_), .Y(new_new_n335_));
  NAi21      g313(.An(i_1_), .B(i_5_), .Y(new_new_n336_));
  INV        g314(.A(new_new_n236_), .Y(new_new_n337_));
  NAi41      g315(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n338_));
  OAI220     g316(.A0(new_new_n338_), .A1(new_new_n336_), .B0(new_new_n212_), .B1(new_new_n159_), .Y(new_new_n339_));
  AOI210     g317(.A0(new_new_n338_), .A1(new_new_n159_), .B0(new_new_n158_), .Y(new_new_n340_));
  NOi32      g318(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n341_));
  NAi21      g319(.An(i_6_), .B(i_1_), .Y(new_new_n342_));
  NA3        g320(.A(new_new_n342_), .B(new_new_n341_), .C(new_new_n47_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n343_), .B(i_0_), .Y(new_new_n344_));
  OR3        g322(.A(new_new_n344_), .B(new_new_n340_), .C(new_new_n339_), .Y(new_new_n345_));
  NO2        g323(.A(i_1_), .B(new_new_n105_), .Y(new_new_n346_));
  NAi21      g324(.An(i_3_), .B(i_4_), .Y(new_new_n347_));
  NO2        g325(.A(new_new_n347_), .B(i_9_), .Y(new_new_n348_));
  AN2        g326(.A(i_6_), .B(i_7_), .Y(new_new_n349_));
  OAI210     g327(.A0(new_new_n349_), .A1(new_new_n346_), .B0(new_new_n348_), .Y(new_new_n350_));
  NA2        g328(.A(i_2_), .B(i_7_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n347_), .B(i_10_), .Y(new_new_n352_));
  NA3        g330(.A(new_new_n352_), .B(new_new_n351_), .C(new_new_n234_), .Y(new_new_n353_));
  AOI210     g331(.A0(new_new_n353_), .A1(new_new_n350_), .B0(new_new_n181_), .Y(new_new_n354_));
  AOI210     g332(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n355_));
  OAI210     g333(.A0(new_new_n355_), .A1(new_new_n182_), .B0(new_new_n352_), .Y(new_new_n356_));
  AOI220     g334(.A0(new_new_n352_), .A1(new_new_n318_), .B0(new_new_n230_), .B1(new_new_n182_), .Y(new_new_n357_));
  AOI210     g335(.A0(new_new_n357_), .A1(new_new_n356_), .B0(i_5_), .Y(new_new_n358_));
  NO4        g336(.A(new_new_n358_), .B(new_new_n354_), .C(new_new_n345_), .D(new_new_n337_), .Y(new_new_n359_));
  NO2        g337(.A(new_new_n359_), .B(new_new_n335_), .Y(new_new_n360_));
  NO2        g338(.A(new_new_n60_), .B(new_new_n25_), .Y(new_new_n361_));
  AN2        g339(.A(i_12_), .B(i_5_), .Y(new_new_n362_));
  NO2        g340(.A(i_4_), .B(new_new_n26_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n363_), .B(new_new_n362_), .Y(new_new_n364_));
  NO2        g342(.A(i_11_), .B(i_6_), .Y(new_new_n365_));
  NA3        g343(.A(new_new_n365_), .B(new_new_n308_), .C(new_new_n217_), .Y(new_new_n366_));
  NO2        g344(.A(new_new_n366_), .B(new_new_n364_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n233_), .B(i_5_), .Y(new_new_n368_));
  NO2        g346(.A(i_5_), .B(i_10_), .Y(new_new_n369_));
  AOI220     g347(.A0(new_new_n369_), .A1(new_new_n260_), .B0(new_new_n368_), .B1(new_new_n191_), .Y(new_new_n370_));
  NA2        g348(.A(new_new_n148_), .B(new_new_n46_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n371_), .B(new_new_n370_), .Y(new_new_n372_));
  OAI210     g350(.A0(new_new_n372_), .A1(new_new_n367_), .B0(new_new_n361_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n374_));
  NO2        g352(.A(new_new_n154_), .B(new_new_n87_), .Y(new_new_n375_));
  OAI210     g353(.A0(new_new_n375_), .A1(new_new_n367_), .B0(new_new_n374_), .Y(new_new_n376_));
  NO3        g354(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n377_));
  NO2        g355(.A(i_11_), .B(i_12_), .Y(new_new_n378_));
  NA3        g356(.A(new_new_n116_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n212_), .Y(new_new_n380_));
  NAi21      g358(.An(i_13_), .B(i_0_), .Y(new_new_n381_));
  NO2        g359(.A(new_new_n381_), .B(new_new_n231_), .Y(new_new_n382_));
  NA2        g360(.A(new_new_n380_), .B(new_new_n382_), .Y(new_new_n383_));
  NA3        g361(.A(new_new_n383_), .B(new_new_n376_), .C(new_new_n373_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n45_), .B(new_new_n217_), .Y(new_new_n385_));
  NO3        g363(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n386_));
  NO2        g364(.A(i_0_), .B(i_11_), .Y(new_new_n387_));
  INV        g365(.A(i_5_), .Y(new_new_n388_));
  AN2        g366(.A(i_1_), .B(i_6_), .Y(new_new_n389_));
  NOi21      g367(.An(i_2_), .B(i_12_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n391_), .B(new_new_n388_), .Y(new_new_n392_));
  NA2        g370(.A(new_new_n146_), .B(i_9_), .Y(new_new_n393_));
  NO2        g371(.A(new_new_n393_), .B(i_4_), .Y(new_new_n394_));
  NA2        g372(.A(new_new_n392_), .B(new_new_n394_), .Y(new_new_n395_));
  NAi21      g373(.An(i_9_), .B(i_4_), .Y(new_new_n396_));
  OR2        g374(.A(i_13_), .B(i_10_), .Y(new_new_n397_));
  NO3        g375(.A(new_new_n397_), .B(new_new_n121_), .C(new_new_n396_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n170_), .B(new_new_n127_), .Y(new_new_n399_));
  NO2        g377(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n400_));
  NO2        g378(.A(new_new_n395_), .B(new_new_n26_), .Y(new_new_n401_));
  NA2        g379(.A(new_new_n305_), .B(new_new_n304_), .Y(new_new_n402_));
  AOI220     g380(.A0(new_new_n280_), .A1(new_new_n270_), .B0(new_new_n274_), .B1(new_new_n297_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n403_), .B(new_new_n167_), .Y(new_new_n404_));
  NO2        g382(.A(new_new_n180_), .B(new_new_n87_), .Y(new_new_n405_));
  NO2        g383(.A(new_new_n404_), .B(new_new_n402_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n190_), .B(new_new_n100_), .Y(new_new_n407_));
  NA3        g385(.A(new_new_n308_), .B(new_new_n162_), .C(new_new_n87_), .Y(new_new_n408_));
  AOI210     g386(.A0(new_new_n408_), .A1(new_new_n407_), .B0(new_new_n306_), .Y(new_new_n409_));
  NO2        g387(.A(i_3_), .B(new_new_n49_), .Y(new_new_n410_));
  NA3        g388(.A(new_new_n318_), .B(new_new_n317_), .C(new_new_n410_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n299_), .B(new_new_n303_), .Y(new_new_n412_));
  OAI210     g390(.A0(new_new_n412_), .A1(new_new_n183_), .B0(new_new_n411_), .Y(new_new_n413_));
  NO2        g391(.A(new_new_n413_), .B(new_new_n409_), .Y(new_new_n414_));
  AOI210     g392(.A0(new_new_n414_), .A1(new_new_n406_), .B0(new_new_n261_), .Y(new_new_n415_));
  NO4        g393(.A(new_new_n415_), .B(new_new_n401_), .C(new_new_n384_), .D(new_new_n360_), .Y(new_new_n416_));
  NO2        g394(.A(new_new_n64_), .B(i_4_), .Y(new_new_n417_));
  NO2        g395(.A(new_new_n74_), .B(i_13_), .Y(new_new_n418_));
  NA3        g396(.A(new_new_n418_), .B(new_new_n417_), .C(i_2_), .Y(new_new_n419_));
  NO2        g397(.A(i_10_), .B(i_9_), .Y(new_new_n420_));
  NAi21      g398(.An(i_12_), .B(i_8_), .Y(new_new_n421_));
  NO2        g399(.A(new_new_n421_), .B(i_3_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n422_), .B(new_new_n420_), .Y(new_new_n423_));
  NO2        g401(.A(new_new_n47_), .B(i_4_), .Y(new_new_n424_));
  NA2        g402(.A(new_new_n424_), .B(new_new_n108_), .Y(new_new_n425_));
  OAI220     g403(.A0(new_new_n425_), .A1(new_new_n194_), .B0(new_new_n423_), .B1(new_new_n419_), .Y(new_new_n426_));
  NA2        g404(.A(new_new_n292_), .B(i_0_), .Y(new_new_n427_));
  NO3        g405(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n428_));
  NA2        g406(.A(new_new_n258_), .B(new_new_n101_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NA2        g408(.A(i_8_), .B(i_9_), .Y(new_new_n431_));
  AOI210     g409(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n432_));
  OR2        g410(.A(new_new_n432_), .B(new_new_n431_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n266_), .B(new_new_n195_), .Y(new_new_n434_));
  OAI220     g412(.A0(new_new_n434_), .A1(new_new_n433_), .B0(new_new_n430_), .B1(new_new_n427_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n241_), .B(new_new_n291_), .Y(new_new_n436_));
  NO3        g414(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n437_));
  INV        g415(.A(new_new_n437_), .Y(new_new_n438_));
  NA3        g416(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n439_));
  NA4        g417(.A(new_new_n149_), .B(new_new_n119_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n440_));
  OAI220     g418(.A0(new_new_n440_), .A1(new_new_n439_), .B0(new_new_n438_), .B1(new_new_n436_), .Y(new_new_n441_));
  NO3        g419(.A(new_new_n441_), .B(new_new_n435_), .C(new_new_n426_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n279_), .B(new_new_n112_), .Y(new_new_n443_));
  OR2        g421(.A(new_new_n443_), .B(new_new_n198_), .Y(new_new_n444_));
  OR2        g422(.A(new_new_n330_), .B(new_new_n105_), .Y(new_new_n445_));
  OA220      g423(.A0(new_new_n445_), .A1(new_new_n161_), .B0(new_new_n444_), .B1(new_new_n224_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n100_), .B(i_13_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n405_), .B(new_new_n361_), .Y(new_new_n448_));
  NO2        g426(.A(i_2_), .B(i_13_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n448_), .B(new_new_n447_), .Y(new_new_n450_));
  NO3        g428(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n451_));
  NO2        g429(.A(i_6_), .B(i_7_), .Y(new_new_n452_));
  NA2        g430(.A(new_new_n452_), .B(new_new_n451_), .Y(new_new_n453_));
  NO2        g431(.A(i_11_), .B(i_1_), .Y(new_new_n454_));
  OR2        g432(.A(i_11_), .B(i_8_), .Y(new_new_n455_));
  NOi21      g433(.An(i_2_), .B(i_7_), .Y(new_new_n456_));
  NAi31      g434(.An(new_new_n455_), .B(new_new_n456_), .C(i_0_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n397_), .B(i_6_), .Y(new_new_n458_));
  NA3        g436(.A(new_new_n458_), .B(new_new_n417_), .C(new_new_n76_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n459_), .B(new_new_n457_), .Y(new_new_n460_));
  NO2        g438(.A(i_3_), .B(new_new_n187_), .Y(new_new_n461_));
  NO2        g439(.A(i_6_), .B(i_10_), .Y(new_new_n462_));
  NA3        g440(.A(new_new_n235_), .B(new_new_n169_), .C(new_new_n136_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n464_));
  NO2        g442(.A(new_new_n158_), .B(i_3_), .Y(new_new_n465_));
  NAi31      g443(.An(new_new_n464_), .B(new_new_n465_), .C(new_new_n218_), .Y(new_new_n466_));
  NA3        g444(.A(new_new_n374_), .B(new_new_n177_), .C(new_new_n153_), .Y(new_new_n467_));
  NA3        g445(.A(new_new_n467_), .B(new_new_n466_), .C(new_new_n463_), .Y(new_new_n468_));
  NO3        g446(.A(new_new_n468_), .B(new_new_n460_), .C(new_new_n450_), .Y(new_new_n469_));
  NA2        g447(.A(new_new_n437_), .B(new_new_n369_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n216_), .Y(new_new_n471_));
  NAi21      g449(.An(new_new_n207_), .B(new_new_n378_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n318_), .B(new_new_n209_), .Y(new_new_n473_));
  NO2        g451(.A(new_new_n473_), .B(new_new_n472_), .Y(new_new_n474_));
  NA2        g452(.A(new_new_n27_), .B(i_10_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n475_), .B(new_new_n447_), .Y(new_new_n476_));
  NA4        g454(.A(new_new_n289_), .B(new_new_n215_), .C(new_new_n74_), .D(new_new_n228_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n477_), .B(new_new_n453_), .Y(new_new_n478_));
  NO4        g456(.A(new_new_n478_), .B(new_new_n476_), .C(new_new_n474_), .D(new_new_n471_), .Y(new_new_n479_));
  NA4        g457(.A(new_new_n479_), .B(new_new_n469_), .C(new_new_n446_), .D(new_new_n442_), .Y(new_new_n480_));
  NA3        g458(.A(new_new_n289_), .B(new_new_n174_), .C(new_new_n172_), .Y(new_new_n481_));
  OAI210     g459(.A0(new_new_n285_), .A1(new_new_n179_), .B0(new_new_n481_), .Y(new_new_n482_));
  AN2        g460(.A(new_new_n270_), .B(new_new_n226_), .Y(new_new_n483_));
  NA2        g461(.A(new_new_n483_), .B(new_new_n482_), .Y(new_new_n484_));
  NA2        g462(.A(new_new_n126_), .B(new_new_n115_), .Y(new_new_n485_));
  AN2        g463(.A(new_new_n485_), .B(new_new_n428_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n296_), .B(new_new_n163_), .Y(new_new_n487_));
  OAI210     g465(.A0(new_new_n487_), .A1(new_new_n224_), .B0(new_new_n290_), .Y(new_new_n488_));
  AOI220     g466(.A0(new_new_n488_), .A1(new_new_n307_), .B0(new_new_n486_), .B1(new_new_n292_), .Y(new_new_n489_));
  NA2        g467(.A(new_new_n334_), .B(new_new_n74_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n349_), .B(new_new_n341_), .Y(new_new_n491_));
  NO2        g469(.A(new_new_n36_), .B(i_8_), .Y(new_new_n492_));
  NAi41      g470(.An(new_new_n490_), .B(new_new_n462_), .C(new_new_n492_), .D(new_new_n47_), .Y(new_new_n493_));
  AOI210     g471(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n398_), .Y(new_new_n494_));
  NA2        g472(.A(new_new_n494_), .B(new_new_n493_), .Y(new_new_n495_));
  NA2        g473(.A(new_new_n247_), .B(new_new_n65_), .Y(new_new_n496_));
  OAI210     g474(.A0(i_8_), .A1(new_new_n496_), .B0(new_new_n138_), .Y(new_new_n497_));
  NA2        g475(.A(new_new_n497_), .B(new_new_n399_), .Y(new_new_n498_));
  NA4        g476(.A(new_new_n498_), .B(new_new_n494_), .C(new_new_n489_), .D(new_new_n484_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n368_), .B(new_new_n279_), .Y(new_new_n500_));
  OAI210     g478(.A0(new_new_n364_), .A1(new_new_n166_), .B0(new_new_n500_), .Y(new_new_n501_));
  NO2        g479(.A(i_12_), .B(new_new_n187_), .Y(new_new_n502_));
  NA2        g480(.A(new_new_n462_), .B(new_new_n27_), .Y(new_new_n503_));
  NO3        g481(.A(new_new_n503_), .B(i_12_), .C(new_new_n443_), .Y(new_new_n504_));
  NOi31      g482(.An(new_new_n299_), .B(new_new_n397_), .C(new_new_n38_), .Y(new_new_n505_));
  OAI210     g483(.A0(new_new_n505_), .A1(new_new_n504_), .B0(new_new_n501_), .Y(new_new_n506_));
  NO2        g484(.A(i_8_), .B(i_7_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n45_), .B(i_10_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n508_), .B(i_6_), .Y(new_new_n509_));
  NOi31      g487(.An(new_new_n274_), .B(new_new_n285_), .C(new_new_n179_), .Y(new_new_n510_));
  NA3        g488(.A(new_new_n289_), .B(new_new_n172_), .C(new_new_n100_), .Y(new_new_n511_));
  NO2        g489(.A(new_new_n213_), .B(new_new_n45_), .Y(new_new_n512_));
  NO2        g490(.A(new_new_n158_), .B(i_5_), .Y(new_new_n513_));
  NA3        g491(.A(new_new_n513_), .B(new_new_n385_), .C(new_new_n301_), .Y(new_new_n514_));
  OAI210     g492(.A0(new_new_n514_), .A1(new_new_n512_), .B0(new_new_n511_), .Y(new_new_n515_));
  OAI210     g493(.A0(new_new_n515_), .A1(new_new_n510_), .B0(new_new_n437_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n516_), .B(new_new_n506_), .Y(new_new_n517_));
  NA3        g495(.A(new_new_n209_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n266_), .B(new_new_n85_), .Y(new_new_n519_));
  AOI210     g497(.A0(new_new_n518_), .A1(new_new_n325_), .B0(new_new_n519_), .Y(new_new_n520_));
  NA2        g498(.A(new_new_n280_), .B(new_new_n270_), .Y(new_new_n521_));
  NO2        g499(.A(new_new_n521_), .B(new_new_n171_), .Y(new_new_n522_));
  NA2        g500(.A(new_new_n215_), .B(new_new_n214_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n420_), .B(new_new_n213_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n523_), .B(new_new_n524_), .Y(new_new_n525_));
  AOI210     g503(.A0(new_new_n342_), .A1(new_new_n47_), .B0(new_new_n346_), .Y(new_new_n526_));
  NA2        g504(.A(i_0_), .B(new_new_n49_), .Y(new_new_n527_));
  NA3        g505(.A(new_new_n502_), .B(new_new_n262_), .C(new_new_n527_), .Y(new_new_n528_));
  NO2        g506(.A(new_new_n526_), .B(new_new_n528_), .Y(new_new_n529_));
  NO4        g507(.A(new_new_n529_), .B(new_new_n525_), .C(new_new_n522_), .D(new_new_n520_), .Y(new_new_n530_));
  NO4        g508(.A(new_new_n242_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n531_));
  NO3        g509(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n532_));
  NO2        g510(.A(new_new_n225_), .B(new_new_n36_), .Y(new_new_n533_));
  AN2        g511(.A(new_new_n533_), .B(new_new_n532_), .Y(new_new_n534_));
  OA210      g512(.A0(new_new_n534_), .A1(new_new_n531_), .B0(new_new_n334_), .Y(new_new_n535_));
  NO2        g513(.A(new_new_n397_), .B(i_1_), .Y(new_new_n536_));
  NOi31      g514(.An(new_new_n536_), .B(new_new_n429_), .C(new_new_n74_), .Y(new_new_n537_));
  AN4        g515(.A(new_new_n537_), .B(new_new_n394_), .C(i_3_), .D(i_2_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n403_), .B(new_new_n175_), .Y(new_new_n539_));
  NO3        g517(.A(new_new_n539_), .B(new_new_n538_), .C(new_new_n535_), .Y(new_new_n540_));
  NOi21      g518(.An(i_10_), .B(i_6_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n542_));
  AOI220     g520(.A0(new_new_n266_), .A1(new_new_n542_), .B0(new_new_n262_), .B1(new_new_n541_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n543_), .B(new_new_n427_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n191_), .B(new_new_n37_), .Y(new_new_n546_));
  NOi31      g524(.An(new_new_n150_), .B(new_new_n546_), .C(new_new_n314_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n547_), .B(new_new_n544_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n490_), .B(new_new_n357_), .Y(new_new_n549_));
  INV        g527(.A(new_new_n301_), .Y(new_new_n550_));
  NO2        g528(.A(i_12_), .B(new_new_n87_), .Y(new_new_n551_));
  OR2        g529(.A(i_2_), .B(i_5_), .Y(new_new_n552_));
  OR2        g530(.A(new_new_n552_), .B(new_new_n389_), .Y(new_new_n553_));
  NA2        g531(.A(new_new_n351_), .B(new_new_n234_), .Y(new_new_n554_));
  AOI210     g532(.A0(new_new_n554_), .A1(new_new_n553_), .B0(new_new_n472_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n555_), .B(new_new_n549_), .Y(new_new_n556_));
  NA4        g534(.A(new_new_n556_), .B(new_new_n548_), .C(new_new_n540_), .D(new_new_n530_), .Y(new_new_n557_));
  NO4        g535(.A(new_new_n557_), .B(new_new_n517_), .C(new_new_n499_), .D(new_new_n480_), .Y(new_new_n558_));
  NA4        g536(.A(new_new_n558_), .B(new_new_n416_), .C(new_new_n333_), .D(new_new_n295_), .Y(mai7));
  NO2        g537(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n560_));
  NA2        g538(.A(i_11_), .B(new_new_n187_), .Y(new_new_n561_));
  NA3        g539(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n562_));
  NO2        g540(.A(new_new_n228_), .B(i_4_), .Y(new_new_n563_));
  NA2        g541(.A(new_new_n563_), .B(i_8_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n109_), .B(new_new_n562_), .Y(new_new_n565_));
  NA2        g543(.A(i_2_), .B(new_new_n87_), .Y(new_new_n566_));
  OAI210     g544(.A0(new_new_n90_), .A1(new_new_n192_), .B0(new_new_n193_), .Y(new_new_n567_));
  NO2        g545(.A(i_7_), .B(new_new_n37_), .Y(new_new_n568_));
  NA2        g546(.A(i_4_), .B(i_8_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n569_), .A1(new_new_n289_), .B0(new_new_n568_), .Y(new_new_n570_));
  OAI220     g548(.A0(new_new_n570_), .A1(new_new_n566_), .B0(new_new_n567_), .B1(i_13_), .Y(new_new_n571_));
  NO3        g549(.A(new_new_n571_), .B(new_new_n565_), .C(new_new_n560_), .Y(new_new_n572_));
  AOI210     g550(.A0(new_new_n132_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n573_));
  AOI210     g551(.A0(new_new_n573_), .A1(new_new_n228_), .B0(new_new_n160_), .Y(new_new_n574_));
  OR2        g552(.A(i_6_), .B(i_10_), .Y(new_new_n575_));
  NO2        g553(.A(new_new_n575_), .B(new_new_n23_), .Y(new_new_n576_));
  OR3        g554(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n577_));
  NO3        g555(.A(new_new_n577_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n578_));
  NO2        g556(.A(new_new_n578_), .B(new_new_n576_), .Y(new_new_n579_));
  OA220      g557(.A0(new_new_n579_), .A1(new_new_n550_), .B0(new_new_n574_), .B1(new_new_n259_), .Y(new_new_n580_));
  AOI210     g558(.A0(new_new_n580_), .A1(new_new_n572_), .B0(new_new_n64_), .Y(new_new_n581_));
  NOi21      g559(.An(i_11_), .B(i_7_), .Y(new_new_n582_));
  AO210      g560(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n583_));
  NO2        g561(.A(new_new_n583_), .B(new_new_n582_), .Y(new_new_n584_));
  NA2        g562(.A(new_new_n584_), .B(new_new_n197_), .Y(new_new_n585_));
  NA3        g563(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n586_));
  NAi31      g564(.An(new_new_n586_), .B(new_new_n206_), .C(i_11_), .Y(new_new_n587_));
  AOI210     g565(.A0(new_new_n587_), .A1(new_new_n585_), .B0(new_new_n64_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n589_));
  AO210      g567(.A0(new_new_n589_), .A1(new_new_n357_), .B0(new_new_n41_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n218_), .B(new_new_n64_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n390_), .B(new_new_n31_), .Y(new_new_n592_));
  OR2        g570(.A(new_new_n199_), .B(new_new_n112_), .Y(new_new_n593_));
  NA2        g571(.A(new_new_n593_), .B(new_new_n592_), .Y(new_new_n594_));
  NO2        g572(.A(new_new_n64_), .B(i_9_), .Y(new_new_n595_));
  NO2        g573(.A(new_new_n595_), .B(i_4_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n596_), .B(new_new_n594_), .Y(new_new_n597_));
  NO2        g575(.A(i_1_), .B(i_12_), .Y(new_new_n598_));
  NA3        g576(.A(new_new_n598_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n599_));
  BUFFER     g577(.A(new_new_n599_), .Y(new_new_n600_));
  NA4        g578(.A(new_new_n600_), .B(new_new_n597_), .C(new_new_n591_), .D(new_new_n590_), .Y(new_new_n601_));
  OAI210     g579(.A0(new_new_n601_), .A1(new_new_n588_), .B0(i_6_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n586_), .B(new_new_n112_), .Y(new_new_n603_));
  NA2        g581(.A(new_new_n603_), .B(new_new_n551_), .Y(new_new_n604_));
  NO2        g582(.A(i_6_), .B(i_11_), .Y(new_new_n605_));
  NA2        g583(.A(new_new_n604_), .B(new_new_n430_), .Y(new_new_n606_));
  NO4        g584(.A(new_new_n206_), .B(new_new_n132_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n607_), .B(new_new_n595_), .Y(new_new_n608_));
  NO3        g586(.A(new_new_n575_), .B(new_new_n225_), .C(new_new_n23_), .Y(new_new_n609_));
  AOI210     g587(.A0(i_1_), .A1(new_new_n250_), .B0(new_new_n609_), .Y(new_new_n610_));
  OAI210     g588(.A0(new_new_n610_), .A1(new_new_n45_), .B0(new_new_n608_), .Y(new_new_n611_));
  NA3        g589(.A(new_new_n507_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n612_));
  INV        g590(.A(i_2_), .Y(new_new_n613_));
  NA2        g591(.A(new_new_n142_), .B(i_9_), .Y(new_new_n614_));
  NA3        g592(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n615_));
  NO2        g593(.A(new_new_n47_), .B(i_1_), .Y(new_new_n616_));
  NA3        g594(.A(new_new_n616_), .B(new_new_n258_), .C(new_new_n45_), .Y(new_new_n617_));
  OAI220     g595(.A0(new_new_n617_), .A1(new_new_n615_), .B0(new_new_n614_), .B1(new_new_n613_), .Y(new_new_n618_));
  AOI210     g596(.A0(new_new_n454_), .A1(new_new_n400_), .B0(new_new_n232_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n619_), .B(new_new_n566_), .Y(new_new_n620_));
  NAi21      g598(.An(new_new_n612_), .B(new_new_n95_), .Y(new_new_n621_));
  NO2        g599(.A(i_11_), .B(new_new_n37_), .Y(new_new_n622_));
  INV        g600(.A(new_new_n621_), .Y(new_new_n623_));
  OR3        g601(.A(new_new_n623_), .B(new_new_n620_), .C(new_new_n618_), .Y(new_new_n624_));
  NO3        g602(.A(new_new_n624_), .B(new_new_n611_), .C(new_new_n606_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n228_), .B(new_new_n105_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n626_), .B(new_new_n582_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n627_), .B(i_1_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n628_), .B(new_new_n577_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n396_), .B(new_new_n87_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n629_), .B(new_new_n47_), .Y(new_new_n631_));
  NA2        g609(.A(i_3_), .B(new_new_n187_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n118_), .Y(new_new_n633_));
  AN2        g611(.A(new_new_n633_), .B(new_new_n509_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n225_), .B(new_new_n45_), .Y(new_new_n635_));
  NO3        g613(.A(new_new_n635_), .B(new_new_n292_), .C(new_new_n229_), .Y(new_new_n636_));
  NO2        g614(.A(new_new_n121_), .B(new_new_n37_), .Y(new_new_n637_));
  NO2        g615(.A(new_new_n637_), .B(i_6_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n87_), .B(i_9_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n639_), .B(new_new_n64_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n640_), .B(new_new_n598_), .Y(new_new_n641_));
  NO4        g619(.A(new_new_n641_), .B(new_new_n638_), .C(new_new_n636_), .D(i_4_), .Y(new_new_n642_));
  NA2        g620(.A(i_1_), .B(i_3_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n642_), .B(new_new_n634_), .Y(new_new_n644_));
  NA4        g622(.A(new_new_n644_), .B(new_new_n631_), .C(new_new_n625_), .D(new_new_n602_), .Y(new_new_n645_));
  NO3        g623(.A(new_new_n455_), .B(i_3_), .C(i_7_), .Y(new_new_n646_));
  NOi21      g624(.An(new_new_n646_), .B(i_10_), .Y(new_new_n647_));
  OA210      g625(.A0(new_new_n647_), .A1(new_new_n235_), .B0(new_new_n87_), .Y(new_new_n648_));
  NA2        g626(.A(new_new_n349_), .B(new_new_n348_), .Y(new_new_n649_));
  NA3        g627(.A(new_new_n462_), .B(new_new_n492_), .C(new_new_n47_), .Y(new_new_n650_));
  NO3        g628(.A(new_new_n456_), .B(new_new_n569_), .C(new_new_n87_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n651_), .B(new_new_n25_), .Y(new_new_n652_));
  NA3        g630(.A(new_new_n160_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n653_));
  NA4        g631(.A(new_new_n653_), .B(new_new_n652_), .C(new_new_n650_), .D(new_new_n649_), .Y(new_new_n654_));
  OAI210     g632(.A0(new_new_n654_), .A1(new_new_n648_), .B0(i_1_), .Y(new_new_n655_));
  AOI210     g633(.A0(new_new_n258_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n347_), .B(i_2_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n657_), .B(new_new_n656_), .Y(new_new_n658_));
  AOI210     g636(.A0(new_new_n658_), .A1(new_new_n655_), .B0(i_13_), .Y(new_new_n659_));
  OR2        g637(.A(i_11_), .B(i_7_), .Y(new_new_n660_));
  NA3        g638(.A(new_new_n660_), .B(new_new_n110_), .C(new_new_n142_), .Y(new_new_n661_));
  AOI220     g639(.A0(new_new_n449_), .A1(new_new_n160_), .B0(new_new_n424_), .B1(new_new_n142_), .Y(new_new_n662_));
  OAI210     g640(.A0(new_new_n662_), .A1(new_new_n45_), .B0(new_new_n661_), .Y(new_new_n663_));
  NO2        g641(.A(new_new_n55_), .B(i_12_), .Y(new_new_n664_));
  INV        g642(.A(new_new_n664_), .Y(new_new_n665_));
  NO2        g643(.A(new_new_n456_), .B(new_new_n24_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n666_), .B(new_new_n630_), .Y(new_new_n667_));
  OAI220     g645(.A0(new_new_n667_), .A1(new_new_n41_), .B0(new_new_n665_), .B1(new_new_n96_), .Y(new_new_n668_));
  AOI210     g646(.A0(new_new_n663_), .A1(new_new_n315_), .B0(new_new_n668_), .Y(new_new_n669_));
  INV        g647(.A(new_new_n118_), .Y(new_new_n670_));
  AOI220     g648(.A0(new_new_n670_), .A1(new_new_n73_), .B0(new_new_n365_), .B1(new_new_n616_), .Y(new_new_n671_));
  NO2        g649(.A(new_new_n671_), .B(new_new_n233_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n131_), .B(i_13_), .Y(new_new_n673_));
  NO2        g651(.A(new_new_n615_), .B(new_new_n118_), .Y(new_new_n674_));
  INV        g652(.A(new_new_n674_), .Y(new_new_n675_));
  OAI220     g653(.A0(new_new_n675_), .A1(new_new_n72_), .B0(new_new_n673_), .B1(new_new_n656_), .Y(new_new_n676_));
  NA2        g654(.A(new_new_n26_), .B(new_new_n187_), .Y(new_new_n677_));
  NA2        g655(.A(new_new_n677_), .B(i_7_), .Y(new_new_n678_));
  AOI220     g656(.A0(new_new_n365_), .A1(new_new_n616_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n679_));
  NO2        g657(.A(new_new_n679_), .B(new_new_n564_), .Y(new_new_n680_));
  NO3        g658(.A(new_new_n680_), .B(new_new_n676_), .C(new_new_n672_), .Y(new_new_n681_));
  OR2        g659(.A(i_11_), .B(i_6_), .Y(new_new_n682_));
  NA3        g660(.A(new_new_n563_), .B(new_new_n677_), .C(i_7_), .Y(new_new_n683_));
  AOI210     g661(.A0(new_new_n683_), .A1(new_new_n675_), .B0(new_new_n682_), .Y(new_new_n684_));
  NA3        g662(.A(new_new_n390_), .B(new_new_n568_), .C(new_new_n101_), .Y(new_new_n685_));
  NA2        g663(.A(new_new_n605_), .B(i_13_), .Y(new_new_n686_));
  NA2        g664(.A(new_new_n106_), .B(new_new_n677_), .Y(new_new_n687_));
  NAi21      g665(.An(i_11_), .B(i_12_), .Y(new_new_n688_));
  NOi41      g666(.An(new_new_n114_), .B(new_new_n688_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n689_), .B(new_new_n687_), .Y(new_new_n690_));
  NA3        g668(.A(new_new_n690_), .B(new_new_n686_), .C(new_new_n685_), .Y(new_new_n691_));
  OAI210     g669(.A0(new_new_n691_), .A1(new_new_n684_), .B0(new_new_n64_), .Y(new_new_n692_));
  NO2        g670(.A(i_2_), .B(i_12_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n346_), .B(new_new_n693_), .Y(new_new_n694_));
  NA2        g672(.A(i_8_), .B(new_new_n25_), .Y(new_new_n695_));
  NO3        g673(.A(new_new_n695_), .B(new_new_n363_), .C(new_new_n563_), .Y(new_new_n696_));
  OAI210     g674(.A0(new_new_n696_), .A1(new_new_n348_), .B0(new_new_n346_), .Y(new_new_n697_));
  NO2        g675(.A(new_new_n132_), .B(i_2_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n697_), .B(new_new_n694_), .Y(new_new_n699_));
  NA3        g677(.A(new_new_n699_), .B(new_new_n46_), .C(new_new_n217_), .Y(new_new_n700_));
  NA4        g678(.A(new_new_n700_), .B(new_new_n692_), .C(new_new_n681_), .D(new_new_n669_), .Y(new_new_n701_));
  OR4        g679(.A(new_new_n701_), .B(new_new_n659_), .C(new_new_n645_), .D(new_new_n581_), .Y(mai5));
  NA2        g680(.A(new_new_n627_), .B(new_new_n260_), .Y(new_new_n703_));
  AN2        g681(.A(new_new_n24_), .B(i_10_), .Y(new_new_n704_));
  NA3        g682(.A(new_new_n704_), .B(new_new_n693_), .C(new_new_n112_), .Y(new_new_n705_));
  NO2        g683(.A(new_new_n564_), .B(i_11_), .Y(new_new_n706_));
  NA2        g684(.A(new_new_n90_), .B(new_new_n706_), .Y(new_new_n707_));
  NA3        g685(.A(new_new_n707_), .B(new_new_n705_), .C(new_new_n703_), .Y(new_new_n708_));
  NO3        g686(.A(i_11_), .B(new_new_n228_), .C(i_13_), .Y(new_new_n709_));
  NO2        g687(.A(new_new_n128_), .B(new_new_n23_), .Y(new_new_n710_));
  NA2        g688(.A(i_12_), .B(i_8_), .Y(new_new_n711_));
  OAI210     g689(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n711_), .Y(new_new_n712_));
  INV        g690(.A(new_new_n420_), .Y(new_new_n713_));
  AOI220     g691(.A0(new_new_n301_), .A1(new_new_n545_), .B0(new_new_n712_), .B1(new_new_n710_), .Y(new_new_n714_));
  INV        g692(.A(new_new_n714_), .Y(new_new_n715_));
  NO2        g693(.A(new_new_n715_), .B(new_new_n708_), .Y(new_new_n716_));
  INV        g694(.A(new_new_n169_), .Y(new_new_n717_));
  INV        g695(.A(new_new_n235_), .Y(new_new_n718_));
  OAI210     g696(.A0(new_new_n657_), .A1(new_new_n422_), .B0(new_new_n114_), .Y(new_new_n719_));
  AOI210     g697(.A0(new_new_n719_), .A1(new_new_n718_), .B0(new_new_n717_), .Y(new_new_n720_));
  NO2        g698(.A(new_new_n431_), .B(new_new_n26_), .Y(new_new_n721_));
  NO2        g699(.A(new_new_n721_), .B(new_new_n400_), .Y(new_new_n722_));
  NA2        g700(.A(new_new_n722_), .B(i_2_), .Y(new_new_n723_));
  INV        g701(.A(new_new_n723_), .Y(new_new_n724_));
  AOI210     g702(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n397_), .Y(new_new_n725_));
  AOI210     g703(.A0(new_new_n725_), .A1(new_new_n724_), .B0(new_new_n720_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n184_), .B(new_new_n129_), .Y(new_new_n727_));
  OAI210     g705(.A0(new_new_n727_), .A1(new_new_n710_), .B0(i_2_), .Y(new_new_n728_));
  INV        g706(.A(new_new_n170_), .Y(new_new_n729_));
  NO3        g707(.A(new_new_n583_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n730_));
  AOI210     g708(.A0(new_new_n729_), .A1(new_new_n90_), .B0(new_new_n730_), .Y(new_new_n731_));
  AOI210     g709(.A0(new_new_n731_), .A1(new_new_n728_), .B0(new_new_n187_), .Y(new_new_n732_));
  OA210      g710(.A0(new_new_n584_), .A1(new_new_n130_), .B0(i_13_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n156_), .B(new_new_n561_), .Y(new_new_n734_));
  NO2        g712(.A(new_new_n734_), .B(new_new_n351_), .Y(new_new_n735_));
  AOI210     g713(.A0(new_new_n199_), .A1(new_new_n152_), .B0(new_new_n492_), .Y(new_new_n736_));
  NA2        g714(.A(new_new_n736_), .B(new_new_n400_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n738_));
  INV        g716(.A(new_new_n286_), .Y(new_new_n739_));
  NA4        g717(.A(new_new_n739_), .B(new_new_n289_), .C(new_new_n128_), .D(new_new_n43_), .Y(new_new_n740_));
  OAI210     g718(.A0(new_new_n740_), .A1(new_new_n738_), .B0(new_new_n737_), .Y(new_new_n741_));
  NO4        g719(.A(new_new_n741_), .B(new_new_n735_), .C(new_new_n733_), .D(new_new_n732_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n545_), .B(new_new_n28_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n709_), .B(new_new_n263_), .Y(new_new_n744_));
  NA2        g722(.A(new_new_n744_), .B(new_new_n743_), .Y(new_new_n745_));
  NO2        g723(.A(new_new_n63_), .B(i_12_), .Y(new_new_n746_));
  NO2        g724(.A(new_new_n746_), .B(new_new_n130_), .Y(new_new_n747_));
  NO2        g725(.A(new_new_n747_), .B(new_new_n561_), .Y(new_new_n748_));
  AOI220     g726(.A0(new_new_n748_), .A1(new_new_n36_), .B0(new_new_n745_), .B1(new_new_n47_), .Y(new_new_n749_));
  NA4        g727(.A(new_new_n749_), .B(new_new_n742_), .C(new_new_n726_), .D(new_new_n716_), .Y(mai6));
  NA4        g728(.A(new_new_n369_), .B(new_new_n461_), .C(new_new_n72_), .D(new_new_n105_), .Y(new_new_n751_));
  INV        g729(.A(new_new_n751_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n212_), .B(new_new_n464_), .Y(new_new_n753_));
  NO2        g731(.A(new_new_n752_), .B(new_new_n313_), .Y(new_new_n754_));
  OR2        g732(.A(new_new_n754_), .B(i_12_), .Y(new_new_n755_));
  NA2        g733(.A(new_new_n352_), .B(new_new_n318_), .Y(new_new_n756_));
  NA2        g734(.A(new_new_n551_), .B(new_new_n64_), .Y(new_new_n757_));
  NA2        g735(.A(new_new_n647_), .B(new_new_n72_), .Y(new_new_n758_));
  BUFFER     g736(.A(new_new_n589_), .Y(new_new_n759_));
  NA4        g737(.A(new_new_n759_), .B(new_new_n758_), .C(new_new_n757_), .D(new_new_n756_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n760_), .B(new_new_n74_), .Y(new_new_n761_));
  INV        g739(.A(new_new_n312_), .Y(new_new_n762_));
  NA2        g740(.A(new_new_n76_), .B(new_new_n135_), .Y(new_new_n763_));
  INV        g741(.A(new_new_n128_), .Y(new_new_n764_));
  NA2        g742(.A(new_new_n764_), .B(new_new_n47_), .Y(new_new_n765_));
  AOI210     g743(.A0(new_new_n765_), .A1(new_new_n763_), .B0(new_new_n762_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n242_), .B(i_9_), .Y(new_new_n767_));
  NA2        g745(.A(new_new_n767_), .B(new_new_n746_), .Y(new_new_n768_));
  AOI210     g746(.A0(new_new_n768_), .A1(new_new_n491_), .B0(new_new_n181_), .Y(new_new_n769_));
  NO2        g747(.A(new_new_n32_), .B(i_11_), .Y(new_new_n770_));
  NA3        g748(.A(new_new_n770_), .B(new_new_n452_), .C(new_new_n369_), .Y(new_new_n771_));
  NAi32      g749(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n772_));
  NO2        g750(.A(new_new_n682_), .B(new_new_n772_), .Y(new_new_n773_));
  NAi21      g751(.An(new_new_n773_), .B(new_new_n771_), .Y(new_new_n774_));
  OR3        g752(.A(new_new_n774_), .B(new_new_n769_), .C(new_new_n766_), .Y(new_new_n775_));
  NO2        g753(.A(new_new_n660_), .B(i_2_), .Y(new_new_n776_));
  OR2        g754(.A(new_new_n584_), .B(new_new_n422_), .Y(new_new_n777_));
  NA3        g755(.A(new_new_n777_), .B(new_new_n151_), .C(new_new_n70_), .Y(new_new_n778_));
  AO210      g756(.A0(new_new_n470_), .A1(new_new_n713_), .B0(new_new_n36_), .Y(new_new_n779_));
  NA2        g757(.A(new_new_n779_), .B(new_new_n778_), .Y(new_new_n780_));
  OAI210     g758(.A0(i_6_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n781_));
  AOI220     g759(.A0(new_new_n781_), .A1(new_new_n532_), .B0(new_new_n753_), .B1(new_new_n678_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n377_), .B(new_new_n71_), .Y(new_new_n783_));
  NA3        g761(.A(new_new_n783_), .B(new_new_n782_), .C(new_new_n567_), .Y(new_new_n784_));
  AO210      g762(.A0(new_new_n492_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n785_));
  NA3        g763(.A(new_new_n785_), .B(new_new_n462_), .C(new_new_n209_), .Y(new_new_n786_));
  AOI210     g764(.A0(new_new_n422_), .A1(new_new_n420_), .B0(new_new_n531_), .Y(new_new_n787_));
  NA2        g765(.A(new_new_n115_), .B(new_new_n387_), .Y(new_new_n788_));
  NA2        g766(.A(new_new_n234_), .B(new_new_n47_), .Y(new_new_n789_));
  INV        g767(.A(new_new_n553_), .Y(new_new_n790_));
  NA3        g768(.A(new_new_n790_), .B(new_new_n312_), .C(i_7_), .Y(new_new_n791_));
  NA4        g769(.A(new_new_n791_), .B(new_new_n788_), .C(new_new_n787_), .D(new_new_n786_), .Y(new_new_n792_));
  NO4        g770(.A(new_new_n792_), .B(new_new_n784_), .C(new_new_n780_), .D(new_new_n775_), .Y(new_new_n793_));
  NA4        g771(.A(new_new_n793_), .B(new_new_n761_), .C(new_new_n755_), .D(new_new_n359_), .Y(mai3));
  NA2        g772(.A(i_12_), .B(i_10_), .Y(new_new_n795_));
  NA2        g773(.A(i_6_), .B(i_7_), .Y(new_new_n796_));
  NO2        g774(.A(new_new_n796_), .B(i_0_), .Y(new_new_n797_));
  NO2        g775(.A(i_11_), .B(new_new_n228_), .Y(new_new_n798_));
  OAI210     g776(.A0(new_new_n797_), .A1(new_new_n274_), .B0(new_new_n798_), .Y(new_new_n799_));
  NO2        g777(.A(new_new_n799_), .B(new_new_n187_), .Y(new_new_n800_));
  NO3        g778(.A(new_new_n427_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n801_));
  OA210      g779(.A0(new_new_n801_), .A1(new_new_n800_), .B0(new_new_n172_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n567_), .B(new_new_n350_), .Y(new_new_n803_));
  NA2        g781(.A(new_new_n803_), .B(new_new_n40_), .Y(new_new_n804_));
  NOi21      g782(.An(new_new_n100_), .B(new_new_n722_), .Y(new_new_n805_));
  NO3        g783(.A(new_new_n593_), .B(new_new_n431_), .C(new_new_n135_), .Y(new_new_n806_));
  AN2        g784(.A(new_new_n429_), .B(new_new_n56_), .Y(new_new_n807_));
  NO3        g785(.A(new_new_n807_), .B(new_new_n806_), .C(new_new_n805_), .Y(new_new_n808_));
  AOI210     g786(.A0(new_new_n808_), .A1(new_new_n804_), .B0(new_new_n49_), .Y(new_new_n809_));
  NO4        g787(.A(new_new_n355_), .B(new_new_n362_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n810_));
  NA2        g788(.A(new_new_n181_), .B(new_new_n541_), .Y(new_new_n811_));
  NOi21      g789(.An(new_new_n811_), .B(new_new_n810_), .Y(new_new_n812_));
  NO2        g790(.A(new_new_n812_), .B(new_new_n64_), .Y(new_new_n813_));
  NOi21      g791(.An(i_5_), .B(i_9_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n814_), .B(new_new_n418_), .Y(new_new_n815_));
  BUFFER     g793(.A(new_new_n258_), .Y(new_new_n816_));
  AOI210     g794(.A0(new_new_n816_), .A1(new_new_n454_), .B0(new_new_n651_), .Y(new_new_n817_));
  NO3        g795(.A(new_new_n393_), .B(new_new_n258_), .C(new_new_n74_), .Y(new_new_n818_));
  NO2        g796(.A(new_new_n173_), .B(new_new_n152_), .Y(new_new_n819_));
  AOI210     g797(.A0(new_new_n819_), .A1(new_new_n234_), .B0(new_new_n818_), .Y(new_new_n820_));
  OAI220     g798(.A0(new_new_n820_), .A1(new_new_n179_), .B0(new_new_n817_), .B1(new_new_n815_), .Y(new_new_n821_));
  NO4        g799(.A(new_new_n821_), .B(new_new_n813_), .C(new_new_n809_), .D(new_new_n802_), .Y(new_new_n822_));
  NA2        g800(.A(new_new_n181_), .B(new_new_n24_), .Y(new_new_n823_));
  NAi21      g801(.An(new_new_n161_), .B(new_new_n410_), .Y(new_new_n824_));
  NO2        g802(.A(new_new_n824_), .B(new_new_n789_), .Y(new_new_n825_));
  INV        g803(.A(new_new_n825_), .Y(new_new_n826_));
  NO2        g804(.A(new_new_n369_), .B(new_new_n278_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n827_), .B(new_new_n674_), .Y(new_new_n828_));
  NA2        g806(.A(new_new_n542_), .B(i_0_), .Y(new_new_n829_));
  NO4        g807(.A(new_new_n552_), .B(new_new_n206_), .C(new_new_n397_), .D(new_new_n389_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n830_), .B(i_11_), .Y(new_new_n831_));
  INV        g809(.A(new_new_n452_), .Y(new_new_n832_));
  NA2        g810(.A(new_new_n709_), .B(new_new_n313_), .Y(new_new_n833_));
  INV        g811(.A(new_new_n59_), .Y(new_new_n834_));
  NO2        g812(.A(new_new_n834_), .B(new_new_n833_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n244_), .B(new_new_n157_), .Y(new_new_n836_));
  NA2        g814(.A(i_0_), .B(i_10_), .Y(new_new_n837_));
  INV        g815(.A(new_new_n508_), .Y(new_new_n838_));
  NO4        g816(.A(new_new_n118_), .B(new_new_n59_), .C(new_new_n632_), .D(i_5_), .Y(new_new_n839_));
  AO220      g817(.A0(new_new_n839_), .A1(new_new_n838_), .B0(new_new_n836_), .B1(i_6_), .Y(new_new_n840_));
  AOI220     g818(.A0(new_new_n316_), .A1(new_new_n102_), .B0(new_new_n181_), .B1(new_new_n85_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n536_), .B(i_4_), .Y(new_new_n842_));
  NA2        g820(.A(new_new_n182_), .B(new_new_n192_), .Y(new_new_n843_));
  OAI220     g821(.A0(new_new_n843_), .A1(new_new_n833_), .B0(new_new_n842_), .B1(new_new_n841_), .Y(new_new_n844_));
  NO3        g822(.A(new_new_n844_), .B(new_new_n840_), .C(new_new_n835_), .Y(new_new_n845_));
  NA4        g823(.A(new_new_n845_), .B(new_new_n831_), .C(new_new_n828_), .D(new_new_n826_), .Y(new_new_n846_));
  NO2        g824(.A(new_new_n107_), .B(new_new_n37_), .Y(new_new_n847_));
  NA2        g825(.A(i_11_), .B(i_9_), .Y(new_new_n848_));
  NO3        g826(.A(i_12_), .B(new_new_n848_), .C(new_new_n566_), .Y(new_new_n849_));
  AN2        g827(.A(new_new_n849_), .B(new_new_n847_), .Y(new_new_n850_));
  NO2        g828(.A(new_new_n49_), .B(i_7_), .Y(new_new_n851_));
  NA2        g829(.A(new_new_n374_), .B(new_new_n177_), .Y(new_new_n852_));
  INV        g830(.A(new_new_n852_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n848_), .B(new_new_n74_), .Y(new_new_n854_));
  NO2        g832(.A(new_new_n173_), .B(i_0_), .Y(new_new_n855_));
  INV        g833(.A(new_new_n855_), .Y(new_new_n856_));
  NA2        g834(.A(new_new_n452_), .B(new_new_n223_), .Y(new_new_n857_));
  AOI210     g835(.A0(new_new_n349_), .A1(new_new_n42_), .B0(new_new_n386_), .Y(new_new_n858_));
  OAI220     g836(.A0(new_new_n858_), .A1(new_new_n815_), .B0(new_new_n857_), .B1(new_new_n856_), .Y(new_new_n859_));
  NO3        g837(.A(new_new_n859_), .B(new_new_n853_), .C(new_new_n850_), .Y(new_new_n860_));
  NA2        g838(.A(new_new_n622_), .B(new_new_n125_), .Y(new_new_n861_));
  NO2        g839(.A(i_6_), .B(new_new_n861_), .Y(new_new_n862_));
  NA2        g840(.A(new_new_n169_), .B(new_new_n107_), .Y(new_new_n863_));
  INV        g841(.A(new_new_n862_), .Y(new_new_n864_));
  NOi21      g842(.An(i_7_), .B(i_5_), .Y(new_new_n865_));
  NOi31      g843(.An(new_new_n865_), .B(i_0_), .C(new_new_n688_), .Y(new_new_n866_));
  NA3        g844(.A(new_new_n866_), .B(new_new_n363_), .C(i_6_), .Y(new_new_n867_));
  OA210      g845(.A0(new_new_n863_), .A1(new_new_n491_), .B0(new_new_n867_), .Y(new_new_n868_));
  NO3        g846(.A(new_new_n381_), .B(new_new_n338_), .C(new_new_n336_), .Y(new_new_n869_));
  NO2        g847(.A(new_new_n253_), .B(new_new_n302_), .Y(new_new_n870_));
  NO2        g848(.A(new_new_n688_), .B(new_new_n248_), .Y(new_new_n871_));
  AOI210     g849(.A0(new_new_n871_), .A1(new_new_n870_), .B0(new_new_n869_), .Y(new_new_n872_));
  NA4        g850(.A(new_new_n872_), .B(new_new_n868_), .C(new_new_n864_), .D(new_new_n860_), .Y(new_new_n873_));
  NO2        g851(.A(new_new_n823_), .B(new_new_n231_), .Y(new_new_n874_));
  AN2        g852(.A(new_new_n315_), .B(new_new_n313_), .Y(new_new_n875_));
  AN2        g853(.A(new_new_n875_), .B(new_new_n819_), .Y(new_new_n876_));
  OAI210     g854(.A0(new_new_n876_), .A1(new_new_n874_), .B0(i_10_), .Y(new_new_n877_));
  NO2        g855(.A(new_new_n795_), .B(new_new_n301_), .Y(new_new_n878_));
  OA210      g856(.A0(new_new_n452_), .A1(new_new_n215_), .B0(new_new_n451_), .Y(new_new_n879_));
  NA2        g857(.A(new_new_n878_), .B(new_new_n854_), .Y(new_new_n880_));
  NA3        g858(.A(new_new_n451_), .B(new_new_n390_), .C(new_new_n46_), .Y(new_new_n881_));
  OAI210     g859(.A0(new_new_n824_), .A1(new_new_n832_), .B0(new_new_n881_), .Y(new_new_n882_));
  NA2        g860(.A(new_new_n854_), .B(new_new_n289_), .Y(new_new_n883_));
  INV        g861(.A(new_new_n883_), .Y(new_new_n884_));
  AOI220     g862(.A0(new_new_n884_), .A1(new_new_n452_), .B0(new_new_n882_), .B1(new_new_n74_), .Y(new_new_n885_));
  NA2        g863(.A(new_new_n666_), .B(new_new_n513_), .Y(new_new_n886_));
  NAi21      g864(.An(i_9_), .B(i_5_), .Y(new_new_n887_));
  NO2        g865(.A(new_new_n887_), .B(new_new_n381_), .Y(new_new_n888_));
  NO2        g866(.A(new_new_n562_), .B(new_new_n109_), .Y(new_new_n889_));
  AOI220     g867(.A0(new_new_n889_), .A1(i_0_), .B0(new_new_n888_), .B1(new_new_n584_), .Y(new_new_n890_));
  OAI220     g868(.A0(new_new_n890_), .A1(new_new_n87_), .B0(new_new_n886_), .B1(new_new_n170_), .Y(new_new_n891_));
  NO2        g869(.A(new_new_n891_), .B(new_new_n495_), .Y(new_new_n892_));
  NA4        g870(.A(new_new_n892_), .B(new_new_n885_), .C(new_new_n880_), .D(new_new_n877_), .Y(new_new_n893_));
  NO3        g871(.A(new_new_n893_), .B(new_new_n873_), .C(new_new_n846_), .Y(new_new_n894_));
  NO2        g872(.A(i_0_), .B(new_new_n688_), .Y(new_new_n895_));
  NA2        g873(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n896_));
  INV        g874(.A(new_new_n896_), .Y(new_new_n897_));
  NO3        g875(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n898_));
  AO220      g876(.A0(new_new_n898_), .A1(new_new_n897_), .B0(new_new_n895_), .B1(new_new_n172_), .Y(new_new_n899_));
  AOI210     g877(.A0(new_new_n757_), .A1(new_new_n649_), .B0(new_new_n863_), .Y(new_new_n900_));
  AOI210     g878(.A0(new_new_n899_), .A1(new_new_n326_), .B0(new_new_n900_), .Y(new_new_n901_));
  NA2        g879(.A(new_new_n698_), .B(new_new_n150_), .Y(new_new_n902_));
  INV        g880(.A(new_new_n902_), .Y(new_new_n903_));
  NA3        g881(.A(new_new_n903_), .B(new_new_n639_), .C(new_new_n74_), .Y(new_new_n904_));
  NA3        g882(.A(new_new_n797_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n905_));
  NA2        g883(.A(new_new_n798_), .B(i_9_), .Y(new_new_n906_));
  NO2        g884(.A(new_new_n905_), .B(new_new_n906_), .Y(new_new_n907_));
  NA2        g885(.A(new_new_n234_), .B(new_new_n222_), .Y(new_new_n908_));
  AOI210     g886(.A0(new_new_n908_), .A1(new_new_n829_), .B0(new_new_n157_), .Y(new_new_n909_));
  NO2        g887(.A(new_new_n909_), .B(new_new_n907_), .Y(new_new_n910_));
  NA3        g888(.A(new_new_n910_), .B(new_new_n904_), .C(new_new_n901_), .Y(new_new_n911_));
  NA2        g889(.A(new_new_n875_), .B(new_new_n351_), .Y(new_new_n912_));
  AOI210     g890(.A0(new_new_n285_), .A1(new_new_n161_), .B0(new_new_n912_), .Y(new_new_n913_));
  NA3        g891(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n914_));
  NA2        g892(.A(new_new_n851_), .B(new_new_n465_), .Y(new_new_n915_));
  AOI210     g893(.A0(new_new_n914_), .A1(new_new_n161_), .B0(new_new_n915_), .Y(new_new_n916_));
  NO2        g894(.A(new_new_n916_), .B(new_new_n913_), .Y(new_new_n917_));
  NO3        g895(.A(new_new_n837_), .B(new_new_n814_), .C(new_new_n184_), .Y(new_new_n918_));
  AOI220     g896(.A0(new_new_n918_), .A1(i_11_), .B0(new_new_n537_), .B1(new_new_n76_), .Y(new_new_n919_));
  NO3        g897(.A(new_new_n201_), .B(new_new_n362_), .C(i_0_), .Y(new_new_n920_));
  OAI210     g898(.A0(new_new_n920_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n921_));
  NA3        g899(.A(new_new_n921_), .B(new_new_n919_), .C(new_new_n917_), .Y(new_new_n922_));
  AOI220     g900(.A0(new_new_n865_), .A1(new_new_n465_), .B0(new_new_n797_), .B1(new_new_n162_), .Y(new_new_n923_));
  NA2        g901(.A(new_new_n329_), .B(new_new_n174_), .Y(new_new_n924_));
  OR2        g902(.A(new_new_n924_), .B(new_new_n923_), .Y(new_new_n925_));
  AOI210     g903(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n173_), .Y(new_new_n926_));
  NA2        g904(.A(new_new_n926_), .B(new_new_n879_), .Y(new_new_n927_));
  NA3        g905(.A(new_new_n576_), .B(new_new_n181_), .C(new_new_n85_), .Y(new_new_n928_));
  NA2        g906(.A(new_new_n928_), .B(new_new_n511_), .Y(new_new_n929_));
  INV        g907(.A(new_new_n929_), .Y(new_new_n930_));
  NA3        g908(.A(new_new_n369_), .B(new_new_n169_), .C(new_new_n168_), .Y(new_new_n931_));
  NA3        g909(.A(new_new_n851_), .B(new_new_n274_), .C(new_new_n222_), .Y(new_new_n932_));
  NA2        g910(.A(new_new_n932_), .B(new_new_n931_), .Y(new_new_n933_));
  NA3        g911(.A(new_new_n369_), .B(new_new_n317_), .C(new_new_n213_), .Y(new_new_n934_));
  INV        g912(.A(new_new_n934_), .Y(new_new_n935_));
  NOi31      g913(.An(new_new_n368_), .B(new_new_n896_), .C(new_new_n231_), .Y(new_new_n936_));
  NO3        g914(.A(new_new_n848_), .B(new_new_n209_), .C(new_new_n184_), .Y(new_new_n937_));
  NO4        g915(.A(new_new_n937_), .B(new_new_n936_), .C(new_new_n935_), .D(new_new_n933_), .Y(new_new_n938_));
  NA4        g916(.A(new_new_n938_), .B(new_new_n930_), .C(new_new_n927_), .D(new_new_n925_), .Y(new_new_n939_));
  INV        g917(.A(new_new_n578_), .Y(new_new_n940_));
  NO3        g918(.A(new_new_n940_), .B(new_new_n527_), .C(new_new_n323_), .Y(new_new_n941_));
  NO2        g919(.A(new_new_n87_), .B(i_5_), .Y(new_new_n942_));
  NA3        g920(.A(new_new_n798_), .B(new_new_n113_), .C(new_new_n128_), .Y(new_new_n943_));
  INV        g921(.A(new_new_n943_), .Y(new_new_n944_));
  AOI210     g922(.A0(new_new_n944_), .A1(new_new_n942_), .B0(new_new_n941_), .Y(new_new_n945_));
  NA3        g923(.A(new_new_n289_), .B(i_5_), .C(new_new_n187_), .Y(new_new_n946_));
  NAi31      g924(.An(new_new_n232_), .B(new_new_n946_), .C(new_new_n233_), .Y(new_new_n947_));
  NO4        g925(.A(new_new_n231_), .B(new_new_n201_), .C(i_0_), .D(i_12_), .Y(new_new_n948_));
  AOI220     g926(.A0(new_new_n948_), .A1(new_new_n947_), .B0(new_new_n752_), .B1(new_new_n174_), .Y(new_new_n949_));
  AN2        g927(.A(new_new_n837_), .B(new_new_n157_), .Y(new_new_n950_));
  NO4        g928(.A(new_new_n950_), .B(i_12_), .C(new_new_n612_), .D(new_new_n135_), .Y(new_new_n951_));
  NA2        g929(.A(new_new_n951_), .B(new_new_n209_), .Y(new_new_n952_));
  NA2        g930(.A(new_new_n865_), .B(new_new_n449_), .Y(new_new_n953_));
  NA2        g931(.A(new_new_n65_), .B(new_new_n105_), .Y(new_new_n954_));
  OAI220     g932(.A0(new_new_n954_), .A1(new_new_n946_), .B0(new_new_n953_), .B1(new_new_n640_), .Y(new_new_n955_));
  NA2        g933(.A(new_new_n955_), .B(new_new_n855_), .Y(new_new_n956_));
  NA4        g934(.A(new_new_n956_), .B(new_new_n952_), .C(new_new_n949_), .D(new_new_n945_), .Y(new_new_n957_));
  NO4        g935(.A(new_new_n957_), .B(new_new_n939_), .C(new_new_n922_), .D(new_new_n911_), .Y(new_new_n958_));
  OAI210     g936(.A0(new_new_n776_), .A1(new_new_n770_), .B0(new_new_n37_), .Y(new_new_n959_));
  NA2        g937(.A(new_new_n959_), .B(new_new_n574_), .Y(new_new_n960_));
  NA2        g938(.A(new_new_n960_), .B(new_new_n197_), .Y(new_new_n961_));
  OAI210     g939(.A0(new_new_n578_), .A1(new_new_n576_), .B0(new_new_n301_), .Y(new_new_n962_));
  NAi31      g940(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n963_));
  AOI210     g941(.A0(new_new_n121_), .A1(new_new_n71_), .B0(new_new_n963_), .Y(new_new_n964_));
  NO2        g942(.A(new_new_n964_), .B(new_new_n609_), .Y(new_new_n965_));
  NA2        g943(.A(new_new_n965_), .B(new_new_n962_), .Y(new_new_n966_));
  NO2        g944(.A(new_new_n439_), .B(new_new_n258_), .Y(new_new_n967_));
  NO4        g945(.A(new_new_n225_), .B(new_new_n149_), .C(new_new_n643_), .D(new_new_n37_), .Y(new_new_n968_));
  NO3        g946(.A(new_new_n968_), .B(new_new_n967_), .C(new_new_n830_), .Y(new_new_n969_));
  INV        g947(.A(new_new_n969_), .Y(new_new_n970_));
  AOI210     g948(.A0(new_new_n966_), .A1(new_new_n49_), .B0(new_new_n970_), .Y(new_new_n971_));
  AOI210     g949(.A0(new_new_n971_), .A1(new_new_n961_), .B0(new_new_n74_), .Y(new_new_n972_));
  NO2        g950(.A(new_new_n534_), .B(new_new_n358_), .Y(new_new_n973_));
  NO2        g951(.A(new_new_n973_), .B(new_new_n717_), .Y(new_new_n974_));
  AOI210     g952(.A0(new_new_n926_), .A1(new_new_n851_), .B0(new_new_n866_), .Y(new_new_n975_));
  NO2        g953(.A(new_new_n975_), .B(new_new_n643_), .Y(new_new_n976_));
  NA2        g954(.A(new_new_n253_), .B(new_new_n58_), .Y(new_new_n977_));
  AOI220     g955(.A0(new_new_n977_), .A1(new_new_n77_), .B0(new_new_n324_), .B1(new_new_n246_), .Y(new_new_n978_));
  NO2        g956(.A(new_new_n978_), .B(new_new_n228_), .Y(new_new_n979_));
  NA3        g957(.A(new_new_n100_), .B(new_new_n291_), .C(new_new_n31_), .Y(new_new_n980_));
  INV        g958(.A(new_new_n980_), .Y(new_new_n981_));
  NO3        g959(.A(new_new_n981_), .B(new_new_n979_), .C(new_new_n976_), .Y(new_new_n982_));
  NA3        g960(.A(new_new_n721_), .B(new_new_n274_), .C(new_new_n81_), .Y(new_new_n983_));
  NO2        g961(.A(new_new_n983_), .B(i_11_), .Y(new_new_n984_));
  INV        g962(.A(new_new_n531_), .Y(new_new_n985_));
  INV        g963(.A(new_new_n339_), .Y(new_new_n986_));
  AOI210     g964(.A0(new_new_n986_), .A1(new_new_n985_), .B0(new_new_n41_), .Y(new_new_n987_));
  NO2        g965(.A(new_new_n987_), .B(new_new_n984_), .Y(new_new_n988_));
  OAI210     g966(.A0(new_new_n982_), .A1(i_4_), .B0(new_new_n988_), .Y(new_new_n989_));
  NO3        g967(.A(new_new_n989_), .B(new_new_n974_), .C(new_new_n972_), .Y(new_new_n990_));
  NA4        g968(.A(new_new_n990_), .B(new_new_n958_), .C(new_new_n894_), .D(new_new_n822_), .Y(mai4));
endmodule


