//Benchmark atmr_alu4_1266_0.25

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n120_, ori_ori_n121_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NOi21      o015(.An(i_12_), .B(i_13_), .Y(ori_ori_n38_));
  INV        o016(.A(ori_ori_n38_), .Y(ori_ori_n39_));
  NAi31      o017(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n35_), .Y(ori1));
  INV        o019(.A(i_11_), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n43_));
  INV        o021(.A(i_2_), .Y(ori_ori_n44_));
  NA2        o022(.A(i_0_), .B(i_3_), .Y(ori_ori_n45_));
  INV        o023(.A(i_5_), .Y(ori_ori_n46_));
  NO2        o024(.A(i_7_), .B(i_10_), .Y(ori_ori_n47_));
  AOI210     o025(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n47_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_5_), .B(ori_ori_n44_), .Y(ori_ori_n49_));
  NA2        o027(.A(i_0_), .B(i_2_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_7_), .B(i_9_), .Y(ori_ori_n51_));
  NO2        o029(.A(ori_ori_n51_), .B(ori_ori_n50_), .Y(ori_ori_n52_));
  NA2        o030(.A(ori_ori_n49_), .B(ori_ori_n43_), .Y(ori_ori_n53_));
  NA3        o031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n54_));
  NO2        o032(.A(i_1_), .B(i_6_), .Y(ori_ori_n55_));
  NA2        o033(.A(i_8_), .B(i_7_), .Y(ori_ori_n56_));
  OAI210     o034(.A0(ori_ori_n56_), .A1(ori_ori_n55_), .B0(ori_ori_n54_), .Y(ori_ori_n57_));
  NA2        o035(.A(ori_ori_n57_), .B(i_12_), .Y(ori_ori_n58_));
  NAi21      o036(.An(i_2_), .B(i_7_), .Y(ori_ori_n59_));
  INV        o037(.A(i_1_), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(i_6_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n59_), .B(ori_ori_n31_), .Y(ori_ori_n62_));
  NA2        o040(.A(i_1_), .B(i_10_), .Y(ori_ori_n63_));
  NO2        o041(.A(ori_ori_n63_), .B(i_6_), .Y(ori_ori_n64_));
  NAi31      o042(.An(ori_ori_n64_), .B(ori_ori_n62_), .C(ori_ori_n58_), .Y(ori_ori_n65_));
  NA2        o043(.A(ori_ori_n48_), .B(i_2_), .Y(ori_ori_n66_));
  AOI210     o044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n67_));
  NA2        o045(.A(i_1_), .B(i_6_), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n68_), .B(ori_ori_n25_), .Y(ori_ori_n69_));
  INV        o047(.A(i_0_), .Y(ori_ori_n70_));
  NAi21      o048(.An(i_5_), .B(i_10_), .Y(ori_ori_n71_));
  NA2        o049(.A(i_5_), .B(i_9_), .Y(ori_ori_n72_));
  AOI210     o050(.A0(ori_ori_n72_), .A1(ori_ori_n71_), .B0(ori_ori_n70_), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n73_), .B(ori_ori_n69_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n67_), .A1(ori_ori_n66_), .B0(ori_ori_n74_), .Y(ori_ori_n75_));
  OAI210     o053(.A0(ori_ori_n75_), .A1(ori_ori_n65_), .B0(i_0_), .Y(ori_ori_n76_));
  NA2        o054(.A(i_12_), .B(i_5_), .Y(ori_ori_n77_));
  INV        o055(.A(i_8_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n78_), .B(ori_ori_n55_), .Y(ori_ori_n79_));
  INV        o057(.A(i_3_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_3_), .B(i_7_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n80_), .B(ori_ori_n60_), .Y(ori_ori_n82_));
  INV        o060(.A(i_6_), .Y(ori_ori_n83_));
  NO2        o061(.A(i_2_), .B(i_7_), .Y(ori_ori_n84_));
  NO2        o062(.A(ori_ori_n82_), .B(ori_ori_n79_), .Y(ori_ori_n85_));
  NAi21      o063(.An(i_6_), .B(i_10_), .Y(ori_ori_n86_));
  NA2        o064(.A(i_6_), .B(i_9_), .Y(ori_ori_n87_));
  NA2        o065(.A(i_2_), .B(i_6_), .Y(ori_ori_n88_));
  AOI210     o066(.A0(ori_ori_n87_), .A1(ori_ori_n85_), .B0(ori_ori_n77_), .Y(ori_ori_n89_));
  AN3        o067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n90_));
  NAi21      o068(.An(i_6_), .B(i_11_), .Y(ori_ori_n91_));
  NA2        o069(.A(ori_ori_n90_), .B(ori_ori_n32_), .Y(ori_ori_n92_));
  INV        o070(.A(i_7_), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n44_), .B(ori_ori_n93_), .Y(ori_ori_n94_));
  NO2        o072(.A(i_0_), .B(i_5_), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n95_), .B(ori_ori_n83_), .Y(ori_ori_n96_));
  NAi21      o074(.An(i_7_), .B(i_11_), .Y(ori_ori_n97_));
  NO3        o075(.A(ori_ori_n97_), .B(ori_ori_n86_), .C(ori_ori_n50_), .Y(ori_ori_n98_));
  AN2        o076(.A(i_2_), .B(i_10_), .Y(ori_ori_n99_));
  NA2        o077(.A(i_12_), .B(i_7_), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n60_), .B(ori_ori_n26_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n101_), .B(i_0_), .Y(ori_ori_n102_));
  NA2        o080(.A(i_11_), .B(i_12_), .Y(ori_ori_n103_));
  OAI210     o081(.A0(ori_ori_n102_), .A1(ori_ori_n100_), .B0(ori_ori_n103_), .Y(ori_ori_n104_));
  INV        o082(.A(ori_ori_n104_), .Y(ori_ori_n105_));
  NAi31      o083(.An(ori_ori_n98_), .B(ori_ori_n105_), .C(ori_ori_n92_), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n93_), .B(ori_ori_n37_), .Y(ori_ori_n107_));
  NA2        o085(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n108_), .B(ori_ori_n107_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n109_), .B(ori_ori_n44_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n87_), .B(ori_ori_n86_), .Y(ori_ori_n111_));
  NAi21      o089(.An(i_3_), .B(i_8_), .Y(ori_ori_n112_));
  NO2        o090(.A(i_1_), .B(ori_ori_n83_), .Y(ori_ori_n113_));
  NO2        o091(.A(i_6_), .B(i_5_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(i_3_), .Y(ori_ori_n115_));
  AO210      o093(.A0(ori_ori_n115_), .A1(ori_ori_n45_), .B0(ori_ori_n113_), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n116_), .B(ori_ori_n97_), .Y(ori_ori_n117_));
  NO3        o095(.A(ori_ori_n117_), .B(ori_ori_n106_), .C(ori_ori_n89_), .Y(ori_ori_n118_));
  NA3        o096(.A(ori_ori_n118_), .B(ori_ori_n76_), .C(ori_ori_n53_), .Y(ori2));
  NO2        o097(.A(ori_ori_n60_), .B(ori_ori_n37_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n657_), .B(ori_ori_n120_), .Y(ori_ori_n121_));
  NA4        o099(.A(ori_ori_n121_), .B(ori_ori_n74_), .C(ori_ori_n66_), .D(ori_ori_n30_), .Y(ori0));
  NO2        o100(.A(i_12_), .B(i_13_), .Y(ori_ori_n123_));
  NAi21      o101(.An(i_5_), .B(i_11_), .Y(ori_ori_n124_));
  NOi21      o102(.An(ori_ori_n123_), .B(ori_ori_n124_), .Y(ori_ori_n125_));
  NO2        o103(.A(i_0_), .B(i_1_), .Y(ori_ori_n126_));
  NA2        o104(.A(i_1_), .B(i_5_), .Y(ori_ori_n127_));
  OR2        o105(.A(i_0_), .B(i_1_), .Y(ori_ori_n128_));
  NAi32      o106(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n129_));
  NOi21      o107(.An(i_4_), .B(i_10_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n130_), .B(ori_ori_n38_), .Y(ori_ori_n131_));
  NOi21      o109(.An(i_4_), .B(i_9_), .Y(ori_ori_n132_));
  NOi21      o110(.An(i_11_), .B(i_13_), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n133_), .B(ori_ori_n132_), .Y(ori_ori_n134_));
  NO2        o112(.A(i_4_), .B(i_5_), .Y(ori_ori_n135_));
  NAi21      o113(.An(i_12_), .B(i_11_), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n136_), .B(i_13_), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n70_), .B(i_5_), .Y(ori_ori_n138_));
  NO2        o116(.A(i_13_), .B(i_10_), .Y(ori_ori_n139_));
  NO2        o117(.A(i_2_), .B(i_1_), .Y(ori_ori_n140_));
  NAi21      o118(.An(i_4_), .B(i_12_), .Y(ori_ori_n141_));
  INV        o119(.A(i_8_), .Y(ori_ori_n142_));
  NO3        o120(.A(i_3_), .B(ori_ori_n83_), .C(ori_ori_n46_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(i_7_), .Y(ori_ori_n144_));
  NO3        o122(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_3_), .B(i_8_), .Y(ori_ori_n146_));
  NO3        o124(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n147_));
  NA3        o125(.A(ori_ori_n147_), .B(ori_ori_n146_), .C(ori_ori_n38_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n95_), .B(ori_ori_n55_), .Y(ori_ori_n149_));
  INV        o127(.A(ori_ori_n149_), .Y(ori_ori_n150_));
  NO2        o128(.A(i_13_), .B(i_9_), .Y(ori_ori_n151_));
  NAi21      o129(.An(i_12_), .B(i_3_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n42_), .B(i_5_), .Y(ori_ori_n153_));
  NO2        o131(.A(ori_ori_n150_), .B(ori_ori_n148_), .Y(ori_ori_n154_));
  INV        o132(.A(ori_ori_n154_), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n155_), .B(i_4_), .Y(ori_ori_n156_));
  NA3        o134(.A(i_13_), .B(ori_ori_n142_), .C(i_10_), .Y(ori_ori_n157_));
  NA2        o135(.A(i_0_), .B(i_5_), .Y(ori_ori_n158_));
  NAi31      o136(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n160_));
  NO2        o138(.A(ori_ori_n70_), .B(ori_ori_n26_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n44_), .B(ori_ori_n60_), .Y(ori_ori_n162_));
  INV        o140(.A(i_13_), .Y(ori_ori_n163_));
  NO2        o141(.A(i_12_), .B(ori_ori_n163_), .Y(ori_ori_n164_));
  NO2        o142(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n165_));
  OR2        o143(.A(i_8_), .B(i_7_), .Y(ori_ori_n166_));
  INV        o144(.A(i_12_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n42_), .B(ori_ori_n167_), .Y(ori_ori_n168_));
  NO3        o146(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n169_));
  NA2        o147(.A(i_2_), .B(i_1_), .Y(ori_ori_n170_));
  NO3        o148(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n171_));
  NAi21      o149(.An(i_4_), .B(i_3_), .Y(ori_ori_n172_));
  NO2        o150(.A(i_0_), .B(i_6_), .Y(ori_ori_n173_));
  NOi41      o151(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n174_), .B(ori_ori_n173_), .Y(ori_ori_n175_));
  NO2        o153(.A(i_11_), .B(ori_ori_n163_), .Y(ori_ori_n176_));
  NOi21      o154(.An(i_1_), .B(i_6_), .Y(ori_ori_n177_));
  NAi21      o155(.An(i_3_), .B(i_7_), .Y(ori_ori_n178_));
  NA2        o156(.A(ori_ori_n167_), .B(i_9_), .Y(ori_ori_n179_));
  OR4        o157(.A(ori_ori_n179_), .B(ori_ori_n178_), .C(ori_ori_n177_), .D(ori_ori_n138_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n70_), .B(i_5_), .Y(ori_ori_n181_));
  NA2        o159(.A(i_3_), .B(i_9_), .Y(ori_ori_n182_));
  NAi21      o160(.An(i_7_), .B(i_10_), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n183_), .B(ori_ori_n182_), .Y(ori_ori_n184_));
  NA3        o162(.A(ori_ori_n184_), .B(ori_ori_n181_), .C(ori_ori_n61_), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n185_), .B(ori_ori_n180_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n186_), .B(ori_ori_n176_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n166_), .B(ori_ori_n37_), .Y(ori_ori_n188_));
  NA2        o166(.A(i_12_), .B(i_6_), .Y(ori_ori_n189_));
  OR2        o167(.A(i_13_), .B(i_9_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n190_), .B(ori_ori_n46_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n172_), .B(i_2_), .Y(ori_ori_n192_));
  NA3        o170(.A(ori_ori_n192_), .B(ori_ori_n191_), .C(ori_ori_n42_), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n176_), .B(i_9_), .Y(ori_ori_n194_));
  OAI210     o172(.A0(ori_ori_n70_), .A1(ori_ori_n194_), .B0(ori_ori_n193_), .Y(ori_ori_n195_));
  NO3        o173(.A(i_11_), .B(ori_ori_n163_), .C(ori_ori_n25_), .Y(ori_ori_n196_));
  NA2        o174(.A(ori_ori_n195_), .B(ori_ori_n188_), .Y(ori_ori_n197_));
  NA2        o175(.A(ori_ori_n197_), .B(ori_ori_n187_), .Y(ori_ori_n198_));
  NO3        o176(.A(i_12_), .B(ori_ori_n163_), .C(ori_ori_n37_), .Y(ori_ori_n199_));
  AN2        o177(.A(i_3_), .B(i_10_), .Y(ori_ori_n200_));
  NO2        o178(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n44_), .B(ori_ori_n26_), .Y(ori_ori_n202_));
  NO2        o180(.A(ori_ori_n198_), .B(ori_ori_n156_), .Y(ori_ori_n203_));
  NO3        o181(.A(ori_ori_n42_), .B(i_13_), .C(i_9_), .Y(ori_ori_n204_));
  NO2        o182(.A(i_2_), .B(i_3_), .Y(ori_ori_n205_));
  NO2        o183(.A(i_12_), .B(i_10_), .Y(ori_ori_n206_));
  NOi21      o184(.An(i_5_), .B(i_0_), .Y(ori_ori_n207_));
  NA4        o185(.A(ori_ori_n81_), .B(ori_ori_n36_), .C(ori_ori_n83_), .D(i_8_), .Y(ori_ori_n208_));
  INV        o186(.A(i_6_), .Y(ori_ori_n209_));
  NO2        o187(.A(i_1_), .B(i_7_), .Y(ori_ori_n210_));
  NOi21      o188(.An(ori_ori_n127_), .B(ori_ori_n96_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(ori_ori_n108_), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n212_), .B(i_3_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n142_), .B(i_9_), .Y(ori_ori_n214_));
  NA2        o192(.A(ori_ori_n214_), .B(ori_ori_n149_), .Y(ori_ori_n215_));
  NO2        o193(.A(ori_ori_n215_), .B(ori_ori_n44_), .Y(ori_ori_n216_));
  INV        o194(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  AOI210     o195(.A0(ori_ori_n217_), .A1(ori_ori_n213_), .B0(ori_ori_n131_), .Y(ori_ori_n218_));
  INV        o196(.A(ori_ori_n218_), .Y(ori_ori_n219_));
  NOi32      o197(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n220_));
  INV        o198(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  NAi21      o199(.An(i_0_), .B(i_6_), .Y(ori_ori_n222_));
  NAi21      o200(.An(i_1_), .B(i_5_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n224_), .B(ori_ori_n25_), .Y(ori_ori_n225_));
  OAI210     o203(.A0(ori_ori_n225_), .A1(ori_ori_n129_), .B0(ori_ori_n175_), .Y(ori_ori_n226_));
  NAi41      o204(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n227_));
  OAI220     o205(.A0(ori_ori_n227_), .A1(ori_ori_n223_), .B0(ori_ori_n159_), .B1(ori_ori_n129_), .Y(ori_ori_n228_));
  NOi32      o206(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n229_));
  NAi21      o207(.An(i_6_), .B(i_1_), .Y(ori_ori_n230_));
  NA3        o208(.A(ori_ori_n230_), .B(ori_ori_n229_), .C(ori_ori_n44_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n231_), .B(i_0_), .Y(ori_ori_n232_));
  OR2        o210(.A(ori_ori_n232_), .B(ori_ori_n228_), .Y(ori_ori_n233_));
  NO2        o211(.A(i_1_), .B(ori_ori_n93_), .Y(ori_ori_n234_));
  NAi21      o212(.An(i_3_), .B(i_4_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n235_), .B(i_9_), .Y(ori_ori_n236_));
  AN2        o214(.A(i_6_), .B(i_7_), .Y(ori_ori_n237_));
  OAI210     o215(.A0(ori_ori_n237_), .A1(ori_ori_n234_), .B0(ori_ori_n236_), .Y(ori_ori_n238_));
  NA2        o216(.A(i_2_), .B(i_7_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n233_), .B(ori_ori_n226_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n240_), .B(ori_ori_n221_), .Y(ori_ori_n241_));
  AN2        o219(.A(i_12_), .B(i_5_), .Y(ori_ori_n242_));
  INV        o220(.A(ori_ori_n242_), .Y(ori_ori_n243_));
  NO2        o221(.A(i_11_), .B(i_6_), .Y(ori_ori_n244_));
  NO2        o222(.A(i_5_), .B(i_10_), .Y(ori_ori_n245_));
  NO2        o223(.A(i_11_), .B(i_12_), .Y(ori_ori_n246_));
  NA2        o224(.A(ori_ori_n246_), .B(ori_ori_n36_), .Y(ori_ori_n247_));
  NO2        o225(.A(i_3_), .B(ori_ori_n247_), .Y(ori_ori_n248_));
  NAi21      o226(.An(i_13_), .B(i_0_), .Y(ori_ori_n249_));
  NO2        o227(.A(ori_ori_n249_), .B(ori_ori_n170_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n248_), .B(ori_ori_n250_), .Y(ori_ori_n251_));
  INV        o229(.A(ori_ori_n251_), .Y(ori_ori_n252_));
  NO2        o230(.A(i_0_), .B(i_11_), .Y(ori_ori_n253_));
  AN2        o231(.A(i_1_), .B(i_6_), .Y(ori_ori_n254_));
  NOi21      o232(.An(i_2_), .B(i_12_), .Y(ori_ori_n255_));
  NAi21      o233(.An(i_9_), .B(i_4_), .Y(ori_ori_n256_));
  OR2        o234(.A(i_13_), .B(i_10_), .Y(ori_ori_n257_));
  NO3        o235(.A(ori_ori_n257_), .B(ori_ori_n103_), .C(ori_ori_n256_), .Y(ori_ori_n258_));
  NO2        o236(.A(ori_ori_n134_), .B(ori_ori_n107_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n93_), .B(ori_ori_n25_), .Y(ori_ori_n260_));
  NA2        o238(.A(ori_ori_n199_), .B(ori_ori_n260_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n261_), .B(ori_ori_n211_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n142_), .B(i_10_), .Y(ori_ori_n263_));
  NA3        o241(.A(ori_ori_n181_), .B(ori_ori_n61_), .C(i_2_), .Y(ori_ori_n264_));
  NO2        o242(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n265_));
  INV        o243(.A(ori_ori_n265_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n266_), .B(ori_ori_n194_), .Y(ori_ori_n267_));
  NO4        o245(.A(ori_ori_n267_), .B(ori_ori_n262_), .C(ori_ori_n252_), .D(ori_ori_n241_), .Y(ori_ori_n268_));
  NO2        o246(.A(ori_ori_n70_), .B(i_13_), .Y(ori_ori_n269_));
  NO2        o247(.A(i_10_), .B(i_9_), .Y(ori_ori_n270_));
  NAi21      o248(.An(i_12_), .B(i_8_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n271_), .B(i_3_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n202_), .B(i_0_), .Y(ori_ori_n273_));
  NO3        o251(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n274_));
  NA2        o252(.A(ori_ori_n189_), .B(ori_ori_n91_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n275_), .B(ori_ori_n274_), .Y(ori_ori_n276_));
  NA2        o254(.A(i_8_), .B(i_9_), .Y(ori_ori_n277_));
  NO2        o255(.A(i_7_), .B(i_2_), .Y(ori_ori_n278_));
  OR2        o256(.A(ori_ori_n278_), .B(ori_ori_n277_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n199_), .B(ori_ori_n149_), .Y(ori_ori_n280_));
  OAI220     o258(.A0(ori_ori_n280_), .A1(ori_ori_n279_), .B0(ori_ori_n276_), .B1(ori_ori_n273_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n176_), .B(ori_ori_n201_), .Y(ori_ori_n282_));
  NO3        o260(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n283_));
  INV        o261(.A(ori_ori_n283_), .Y(ori_ori_n284_));
  NA3        o262(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n285_));
  NA4        o263(.A(ori_ori_n124_), .B(ori_ori_n101_), .C(ori_ori_n77_), .D(ori_ori_n23_), .Y(ori_ori_n286_));
  OAI220     o264(.A0(ori_ori_n286_), .A1(ori_ori_n285_), .B0(ori_ori_n284_), .B1(ori_ori_n282_), .Y(ori_ori_n287_));
  NO2        o265(.A(ori_ori_n287_), .B(ori_ori_n281_), .Y(ori_ori_n288_));
  OR2        o266(.A(ori_ori_n215_), .B(ori_ori_n93_), .Y(ori_ori_n289_));
  OR2        o267(.A(ori_ori_n289_), .B(ori_ori_n131_), .Y(ori_ori_n290_));
  NO2        o268(.A(i_2_), .B(i_13_), .Y(ori_ori_n291_));
  NO3        o269(.A(i_4_), .B(ori_ori_n46_), .C(i_8_), .Y(ori_ori_n292_));
  NO2        o270(.A(i_6_), .B(i_7_), .Y(ori_ori_n293_));
  NO2        o271(.A(i_11_), .B(i_1_), .Y(ori_ori_n294_));
  NOi21      o272(.An(i_2_), .B(i_7_), .Y(ori_ori_n295_));
  NO2        o273(.A(i_3_), .B(ori_ori_n142_), .Y(ori_ori_n296_));
  NO2        o274(.A(i_6_), .B(i_10_), .Y(ori_ori_n297_));
  NA3        o275(.A(ori_ori_n174_), .B(ori_ori_n133_), .C(ori_ori_n114_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n44_), .B(ori_ori_n42_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n283_), .B(ori_ori_n245_), .Y(ori_ori_n300_));
  NAi21      o278(.An(ori_ori_n157_), .B(ori_ori_n246_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n210_), .B(ori_ori_n158_), .Y(ori_ori_n302_));
  NO2        o280(.A(ori_ori_n302_), .B(ori_ori_n301_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n204_), .B(ori_ori_n169_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n304_), .B(ori_ori_n264_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n305_), .B(ori_ori_n303_), .Y(ori_ori_n306_));
  NA4        o284(.A(ori_ori_n306_), .B(ori_ori_n298_), .C(ori_ori_n290_), .D(ori_ori_n288_), .Y(ori_ori_n307_));
  NA2        o285(.A(ori_ori_n242_), .B(ori_ori_n163_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n237_), .B(ori_ori_n229_), .Y(ori_ori_n309_));
  OR2        o287(.A(ori_ori_n308_), .B(ori_ori_n309_), .Y(ori_ori_n310_));
  INV        o288(.A(ori_ori_n258_), .Y(ori_ori_n311_));
  NA2        o289(.A(ori_ori_n311_), .B(ori_ori_n310_), .Y(ori_ori_n312_));
  INV        o290(.A(ori_ori_n312_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n181_), .B(ori_ori_n61_), .Y(ori_ori_n314_));
  OAI210     o292(.A0(i_8_), .A1(ori_ori_n314_), .B0(ori_ori_n116_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n315_), .B(ori_ori_n259_), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n316_), .B(ori_ori_n313_), .Y(ori_ori_n317_));
  NO2        o295(.A(i_12_), .B(ori_ori_n142_), .Y(ori_ori_n318_));
  NA3        o296(.A(ori_ori_n200_), .B(ori_ori_n135_), .C(ori_ori_n90_), .Y(ori_ori_n319_));
  NO2        o297(.A(ori_ori_n128_), .B(i_5_), .Y(ori_ori_n320_));
  NA2        o298(.A(ori_ori_n658_), .B(ori_ori_n283_), .Y(ori_ori_n321_));
  INV        o299(.A(ori_ori_n321_), .Y(ori_ori_n322_));
  NA3        o300(.A(ori_ori_n158_), .B(ori_ori_n68_), .C(ori_ori_n42_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n199_), .B(ori_ori_n81_), .Y(ori_ori_n324_));
  NO2        o302(.A(ori_ori_n323_), .B(ori_ori_n324_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n162_), .B(ori_ori_n161_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n270_), .B(ori_ori_n160_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n326_), .B(ori_ori_n327_), .Y(ori_ori_n328_));
  AOI210     o306(.A0(ori_ori_n230_), .A1(ori_ori_n44_), .B0(ori_ori_n234_), .Y(ori_ori_n329_));
  NA2        o307(.A(i_0_), .B(ori_ori_n46_), .Y(ori_ori_n330_));
  NA3        o308(.A(ori_ori_n318_), .B(ori_ori_n196_), .C(ori_ori_n330_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n329_), .B(ori_ori_n331_), .Y(ori_ori_n332_));
  NO3        o310(.A(ori_ori_n332_), .B(ori_ori_n328_), .C(ori_ori_n325_), .Y(ori_ori_n333_));
  NO4        o311(.A(ori_ori_n177_), .B(ori_ori_n40_), .C(i_2_), .D(ori_ori_n46_), .Y(ori_ori_n334_));
  NOi21      o312(.An(i_10_), .B(i_6_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n83_), .B(ori_ori_n25_), .Y(ori_ori_n336_));
  AOI220     o314(.A0(ori_ori_n199_), .A1(ori_ori_n336_), .B0(ori_ori_n196_), .B1(ori_ori_n335_), .Y(ori_ori_n337_));
  NO2        o315(.A(ori_ori_n337_), .B(ori_ori_n273_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n100_), .B(ori_ori_n23_), .Y(ori_ori_n339_));
  NOi31      o317(.An(ori_ori_n125_), .B(i_10_), .C(ori_ori_n208_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n340_), .B(ori_ori_n338_), .Y(ori_ori_n341_));
  INV        o319(.A(ori_ori_n205_), .Y(ori_ori_n342_));
  NO2        o320(.A(i_12_), .B(ori_ori_n83_), .Y(ori_ori_n343_));
  NA3        o321(.A(ori_ori_n343_), .B(ori_ori_n196_), .C(ori_ori_n330_), .Y(ori_ori_n344_));
  NA3        o322(.A(ori_ori_n244_), .B(ori_ori_n199_), .C(ori_ori_n158_), .Y(ori_ori_n345_));
  AOI210     o323(.A0(ori_ori_n345_), .A1(ori_ori_n344_), .B0(ori_ori_n342_), .Y(ori_ori_n346_));
  OR2        o324(.A(i_2_), .B(i_5_), .Y(ori_ori_n347_));
  OR2        o325(.A(ori_ori_n347_), .B(ori_ori_n254_), .Y(ori_ori_n348_));
  NA2        o326(.A(ori_ori_n239_), .B(ori_ori_n173_), .Y(ori_ori_n349_));
  AOI210     o327(.A0(ori_ori_n349_), .A1(ori_ori_n348_), .B0(ori_ori_n301_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n350_), .B(ori_ori_n346_), .Y(ori_ori_n351_));
  NA3        o329(.A(ori_ori_n351_), .B(ori_ori_n341_), .C(ori_ori_n333_), .Y(ori_ori_n352_));
  NO4        o330(.A(ori_ori_n352_), .B(ori_ori_n322_), .C(ori_ori_n317_), .D(ori_ori_n307_), .Y(ori_ori_n353_));
  NA4        o331(.A(ori_ori_n353_), .B(ori_ori_n268_), .C(ori_ori_n219_), .D(ori_ori_n203_), .Y(ori7));
  NO2        o332(.A(ori_ori_n88_), .B(ori_ori_n51_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n97_), .B(ori_ori_n86_), .Y(ori_ori_n356_));
  INV        o334(.A(ori_ori_n356_), .Y(ori_ori_n357_));
  NA2        o335(.A(ori_ori_n297_), .B(ori_ori_n81_), .Y(ori_ori_n358_));
  NA2        o336(.A(i_11_), .B(ori_ori_n142_), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n123_), .B(ori_ori_n359_), .Y(ori_ori_n360_));
  OAI210     o338(.A0(ori_ori_n360_), .A1(ori_ori_n358_), .B0(ori_ori_n357_), .Y(ori_ori_n361_));
  NA2        o339(.A(i_2_), .B(ori_ori_n83_), .Y(ori_ori_n362_));
  OAI210     o340(.A0(ori_ori_n84_), .A1(ori_ori_n146_), .B0(ori_ori_n147_), .Y(ori_ori_n363_));
  NO2        o341(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n364_));
  NA2        o342(.A(i_4_), .B(i_8_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n361_), .B(ori_ori_n355_), .Y(ori_ori_n366_));
  AOI210     o344(.A0(ori_ori_n112_), .A1(ori_ori_n59_), .B0(i_10_), .Y(ori_ori_n367_));
  AOI210     o345(.A0(ori_ori_n367_), .A1(ori_ori_n167_), .B0(ori_ori_n130_), .Y(ori_ori_n368_));
  OR2        o346(.A(i_6_), .B(i_10_), .Y(ori_ori_n369_));
  OR3        o347(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n370_));
  INV        o348(.A(ori_ori_n145_), .Y(ori_ori_n371_));
  OR2        o349(.A(ori_ori_n368_), .B(ori_ori_n190_), .Y(ori_ori_n372_));
  AOI210     o350(.A0(ori_ori_n372_), .A1(ori_ori_n366_), .B0(ori_ori_n60_), .Y(ori_ori_n373_));
  NOi21      o351(.An(i_11_), .B(i_7_), .Y(ori_ori_n374_));
  AO210      o352(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n375_));
  NO2        o353(.A(ori_ori_n375_), .B(ori_ori_n374_), .Y(ori_ori_n376_));
  NA2        o354(.A(ori_ori_n376_), .B(ori_ori_n151_), .Y(ori_ori_n377_));
  NA3        o355(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n378_));
  NAi31      o356(.An(ori_ori_n378_), .B(i_12_), .C(i_11_), .Y(ori_ori_n379_));
  AOI210     o357(.A0(ori_ori_n379_), .A1(ori_ori_n377_), .B0(ori_ori_n60_), .Y(ori_ori_n380_));
  NO3        o358(.A(ori_ori_n183_), .B(ori_ori_n152_), .C(ori_ori_n359_), .Y(ori_ori_n381_));
  OAI210     o359(.A0(ori_ori_n381_), .A1(ori_ori_n164_), .B0(ori_ori_n60_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n255_), .B(ori_ori_n31_), .Y(ori_ori_n383_));
  OR2        o361(.A(ori_ori_n152_), .B(ori_ori_n97_), .Y(ori_ori_n384_));
  NA2        o362(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n385_));
  NO2        o363(.A(i_1_), .B(i_4_), .Y(ori_ori_n386_));
  NA2        o364(.A(ori_ori_n386_), .B(ori_ori_n385_), .Y(ori_ori_n387_));
  NO2        o365(.A(i_1_), .B(i_12_), .Y(ori_ori_n388_));
  NA3        o366(.A(ori_ori_n388_), .B(ori_ori_n99_), .C(ori_ori_n24_), .Y(ori_ori_n389_));
  BUFFER     o367(.A(ori_ori_n389_), .Y(ori_ori_n390_));
  NA3        o368(.A(ori_ori_n390_), .B(ori_ori_n387_), .C(ori_ori_n382_), .Y(ori_ori_n391_));
  OAI210     o369(.A0(ori_ori_n391_), .A1(ori_ori_n380_), .B0(i_6_), .Y(ori_ori_n392_));
  NO2        o370(.A(ori_ori_n378_), .B(ori_ori_n97_), .Y(ori_ori_n393_));
  NA2        o371(.A(ori_ori_n393_), .B(ori_ori_n343_), .Y(ori_ori_n394_));
  NO2        o372(.A(i_6_), .B(i_11_), .Y(ori_ori_n395_));
  NA2        o373(.A(ori_ori_n394_), .B(ori_ori_n276_), .Y(ori_ori_n396_));
  NO3        o374(.A(ori_ori_n369_), .B(ori_ori_n166_), .C(ori_ori_n23_), .Y(ori_ori_n397_));
  AOI210     o375(.A0(i_1_), .A1(ori_ori_n184_), .B0(ori_ori_n397_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n398_), .B(ori_ori_n42_), .Y(ori_ori_n399_));
  NA3        o377(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n400_));
  NO2        o378(.A(ori_ori_n44_), .B(i_1_), .Y(ori_ori_n401_));
  NA3        o379(.A(ori_ori_n401_), .B(ori_ori_n189_), .C(ori_ori_n42_), .Y(ori_ori_n402_));
  NO2        o380(.A(ori_ori_n402_), .B(ori_ori_n400_), .Y(ori_ori_n403_));
  AOI210     o381(.A0(ori_ori_n294_), .A1(ori_ori_n260_), .B0(ori_ori_n171_), .Y(ori_ori_n404_));
  NO2        o382(.A(ori_ori_n404_), .B(ori_ori_n362_), .Y(ori_ori_n405_));
  OR2        o383(.A(ori_ori_n405_), .B(ori_ori_n403_), .Y(ori_ori_n406_));
  NO3        o384(.A(ori_ori_n406_), .B(ori_ori_n399_), .C(ori_ori_n396_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n167_), .B(ori_ori_n93_), .Y(ori_ori_n408_));
  NO2        o386(.A(ori_ori_n408_), .B(ori_ori_n374_), .Y(ori_ori_n409_));
  NA2        o387(.A(ori_ori_n409_), .B(i_1_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n410_), .B(ori_ori_n370_), .Y(ori_ori_n411_));
  NO2        o389(.A(ori_ori_n256_), .B(ori_ori_n83_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n411_), .B(ori_ori_n44_), .Y(ori_ori_n413_));
  NA2        o391(.A(i_3_), .B(ori_ori_n142_), .Y(ori_ori_n414_));
  NO2        o392(.A(ori_ori_n166_), .B(ori_ori_n42_), .Y(ori_ori_n415_));
  NO3        o393(.A(ori_ori_n415_), .B(ori_ori_n202_), .C(ori_ori_n168_), .Y(ori_ori_n416_));
  NO2        o394(.A(ori_ori_n103_), .B(ori_ori_n37_), .Y(ori_ori_n417_));
  INV        o395(.A(i_6_), .Y(ori_ori_n418_));
  NO2        o396(.A(ori_ori_n83_), .B(i_9_), .Y(ori_ori_n419_));
  NO2        o397(.A(ori_ori_n419_), .B(ori_ori_n60_), .Y(ori_ori_n420_));
  NO2        o398(.A(ori_ori_n420_), .B(ori_ori_n388_), .Y(ori_ori_n421_));
  NO4        o399(.A(ori_ori_n421_), .B(ori_ori_n418_), .C(ori_ori_n416_), .D(i_4_), .Y(ori_ori_n422_));
  NA2        o400(.A(i_1_), .B(i_3_), .Y(ori_ori_n423_));
  NO2        o401(.A(ori_ori_n277_), .B(ori_ori_n88_), .Y(ori_ori_n424_));
  INV        o402(.A(ori_ori_n424_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n425_), .B(ori_ori_n423_), .Y(ori_ori_n426_));
  NO2        o404(.A(ori_ori_n426_), .B(ori_ori_n422_), .Y(ori_ori_n427_));
  NA4        o405(.A(ori_ori_n427_), .B(ori_ori_n413_), .C(ori_ori_n407_), .D(ori_ori_n392_), .Y(ori_ori_n428_));
  NA2        o406(.A(ori_ori_n237_), .B(ori_ori_n236_), .Y(ori_ori_n429_));
  NO3        o407(.A(ori_ori_n295_), .B(ori_ori_n365_), .C(ori_ori_n83_), .Y(ori_ori_n430_));
  NA2        o408(.A(ori_ori_n430_), .B(ori_ori_n25_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n431_), .B(ori_ori_n429_), .Y(ori_ori_n432_));
  NA2        o410(.A(ori_ori_n432_), .B(i_1_), .Y(ori_ori_n433_));
  INV        o411(.A(i_1_), .Y(ori_ori_n434_));
  NO2        o412(.A(ori_ori_n433_), .B(i_13_), .Y(ori_ori_n435_));
  NA3        o413(.A(i_7_), .B(i_12_), .C(ori_ori_n120_), .Y(ori_ori_n436_));
  AOI220     o414(.A0(ori_ori_n291_), .A1(ori_ori_n130_), .B0(i_2_), .B1(ori_ori_n120_), .Y(ori_ori_n437_));
  NA2        o415(.A(ori_ori_n437_), .B(ori_ori_n436_), .Y(ori_ori_n438_));
  NO2        o416(.A(ori_ori_n295_), .B(ori_ori_n24_), .Y(ori_ori_n439_));
  AOI220     o417(.A0(ori_ori_n439_), .A1(ori_ori_n412_), .B0(ori_ori_n174_), .B1(ori_ori_n113_), .Y(ori_ori_n440_));
  NO2        o418(.A(ori_ori_n440_), .B(ori_ori_n39_), .Y(ori_ori_n441_));
  AOI210     o419(.A0(ori_ori_n438_), .A1(ori_ori_n209_), .B0(ori_ori_n441_), .Y(ori_ori_n442_));
  INV        o420(.A(ori_ori_n100_), .Y(ori_ori_n443_));
  AOI220     o421(.A0(ori_ori_n443_), .A1(ori_ori_n69_), .B0(ori_ori_n244_), .B1(ori_ori_n401_), .Y(ori_ori_n444_));
  NO2        o422(.A(ori_ori_n444_), .B(ori_ori_n172_), .Y(ori_ori_n445_));
  NA2        o423(.A(ori_ori_n111_), .B(i_13_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n400_), .B(ori_ori_n100_), .Y(ori_ori_n447_));
  INV        o425(.A(ori_ori_n447_), .Y(ori_ori_n448_));
  OAI220     o426(.A0(ori_ori_n448_), .A1(ori_ori_n68_), .B0(ori_ori_n446_), .B1(ori_ori_n434_), .Y(ori_ori_n449_));
  NO3        o427(.A(ori_ori_n68_), .B(ori_ori_n32_), .C(ori_ori_n93_), .Y(ori_ori_n450_));
  NA2        o428(.A(ori_ori_n26_), .B(ori_ori_n142_), .Y(ori_ori_n451_));
  NO2        o429(.A(ori_ori_n660_), .B(ori_ori_n371_), .Y(ori_ori_n452_));
  NO3        o430(.A(ori_ori_n452_), .B(ori_ori_n449_), .C(ori_ori_n445_), .Y(ori_ori_n453_));
  OR2        o431(.A(i_11_), .B(i_6_), .Y(ori_ori_n454_));
  NA3        o432(.A(i_12_), .B(ori_ori_n451_), .C(i_7_), .Y(ori_ori_n455_));
  NO2        o433(.A(ori_ori_n455_), .B(ori_ori_n454_), .Y(ori_ori_n456_));
  NA2        o434(.A(ori_ori_n395_), .B(i_13_), .Y(ori_ori_n457_));
  NA2        o435(.A(ori_ori_n94_), .B(ori_ori_n451_), .Y(ori_ori_n458_));
  NAi21      o436(.An(i_11_), .B(i_12_), .Y(ori_ori_n459_));
  NO3        o437(.A(ori_ori_n459_), .B(i_13_), .C(ori_ori_n83_), .Y(ori_ori_n460_));
  NO3        o438(.A(ori_ori_n295_), .B(ori_ori_n343_), .C(ori_ori_n365_), .Y(ori_ori_n461_));
  AOI220     o439(.A0(ori_ori_n461_), .A1(ori_ori_n204_), .B0(ori_ori_n460_), .B1(ori_ori_n458_), .Y(ori_ori_n462_));
  NA2        o440(.A(ori_ori_n462_), .B(ori_ori_n457_), .Y(ori_ori_n463_));
  OAI210     o441(.A0(ori_ori_n463_), .A1(ori_ori_n456_), .B0(ori_ori_n60_), .Y(ori_ori_n464_));
  NO2        o442(.A(i_2_), .B(i_12_), .Y(ori_ori_n465_));
  INV        o443(.A(i_2_), .Y(ori_ori_n466_));
  NA2        o444(.A(ori_ori_n466_), .B(ori_ori_n388_), .Y(ori_ori_n467_));
  INV        o445(.A(ori_ori_n467_), .Y(ori_ori_n468_));
  NA3        o446(.A(ori_ori_n468_), .B(ori_ori_n43_), .C(ori_ori_n163_), .Y(ori_ori_n469_));
  NA4        o447(.A(ori_ori_n469_), .B(ori_ori_n464_), .C(ori_ori_n453_), .D(ori_ori_n442_), .Y(ori_ori_n470_));
  OR4        o448(.A(ori_ori_n470_), .B(ori_ori_n435_), .C(ori_ori_n428_), .D(ori_ori_n373_), .Y(ori5));
  NA2        o449(.A(ori_ori_n409_), .B(ori_ori_n192_), .Y(ori_ori_n472_));
  AN2        o450(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n473_), .B(ori_ori_n465_), .Y(ori_ori_n474_));
  NA2        o452(.A(ori_ori_n474_), .B(ori_ori_n472_), .Y(ori_ori_n475_));
  NO3        o453(.A(i_11_), .B(ori_ori_n167_), .C(i_13_), .Y(ori_ori_n476_));
  NO2        o454(.A(ori_ori_n108_), .B(ori_ori_n23_), .Y(ori_ori_n477_));
  INV        o455(.A(ori_ori_n270_), .Y(ori_ori_n478_));
  INV        o456(.A(ori_ori_n475_), .Y(ori_ori_n479_));
  INV        o457(.A(ori_ori_n133_), .Y(ori_ori_n480_));
  INV        o458(.A(ori_ori_n174_), .Y(ori_ori_n481_));
  NO2        o459(.A(ori_ori_n481_), .B(ori_ori_n480_), .Y(ori_ori_n482_));
  NO2        o460(.A(ori_ori_n277_), .B(ori_ori_n26_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n483_), .B(ori_ori_n260_), .Y(ori_ori_n484_));
  NA2        o462(.A(ori_ori_n484_), .B(i_2_), .Y(ori_ori_n485_));
  INV        o463(.A(ori_ori_n485_), .Y(ori_ori_n486_));
  AOI210     o464(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n257_), .Y(ori_ori_n487_));
  AOI210     o465(.A0(ori_ori_n487_), .A1(ori_ori_n486_), .B0(ori_ori_n482_), .Y(ori_ori_n488_));
  NO2        o466(.A(ori_ori_n141_), .B(ori_ori_n109_), .Y(ori_ori_n489_));
  OAI210     o467(.A0(ori_ori_n489_), .A1(ori_ori_n477_), .B0(i_2_), .Y(ori_ori_n490_));
  AOI210     o468(.A0(ori_ori_n134_), .A1(ori_ori_n490_), .B0(ori_ori_n142_), .Y(ori_ori_n491_));
  OA210      o469(.A0(ori_ori_n376_), .A1(ori_ori_n110_), .B0(i_13_), .Y(ori_ori_n492_));
  NA2        o470(.A(ori_ori_n145_), .B(ori_ori_n146_), .Y(ori_ori_n493_));
  NO2        o471(.A(ori_ori_n493_), .B(ori_ori_n239_), .Y(ori_ori_n494_));
  NO2        o472(.A(ori_ori_n152_), .B(ori_ori_n661_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n495_), .B(ori_ori_n260_), .Y(ori_ori_n496_));
  NA2        o474(.A(ori_ori_n93_), .B(ori_ori_n200_), .Y(ori_ori_n497_));
  OAI210     o475(.A0(ori_ori_n497_), .A1(i_11_), .B0(ori_ori_n496_), .Y(ori_ori_n498_));
  NO4        o476(.A(ori_ori_n498_), .B(ori_ori_n494_), .C(ori_ori_n492_), .D(ori_ori_n491_), .Y(ori_ori_n499_));
  NA2        o477(.A(ori_ori_n339_), .B(ori_ori_n28_), .Y(ori_ori_n500_));
  INV        o478(.A(ori_ori_n500_), .Y(ori_ori_n501_));
  NO2        o479(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n502_));
  NO2        o480(.A(ori_ori_n502_), .B(ori_ori_n110_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n503_), .B(ori_ori_n359_), .Y(ori_ori_n504_));
  AOI220     o482(.A0(ori_ori_n504_), .A1(ori_ori_n36_), .B0(ori_ori_n501_), .B1(ori_ori_n44_), .Y(ori_ori_n505_));
  NA4        o483(.A(ori_ori_n505_), .B(ori_ori_n499_), .C(ori_ori_n488_), .D(ori_ori_n479_), .Y(ori6));
  NA4        o484(.A(ori_ori_n245_), .B(ori_ori_n296_), .C(ori_ori_n68_), .D(ori_ori_n93_), .Y(ori_ori_n507_));
  INV        o485(.A(ori_ori_n507_), .Y(ori_ori_n508_));
  NO2        o486(.A(ori_ori_n159_), .B(ori_ori_n299_), .Y(ori_ori_n509_));
  NO2        o487(.A(i_11_), .B(i_9_), .Y(ori_ori_n510_));
  NO2        o488(.A(ori_ori_n508_), .B(ori_ori_n207_), .Y(ori_ori_n511_));
  OR2        o489(.A(ori_ori_n511_), .B(i_12_), .Y(ori_ori_n512_));
  NA2        o490(.A(ori_ori_n343_), .B(ori_ori_n60_), .Y(ori_ori_n513_));
  INV        o491(.A(ori_ori_n513_), .Y(ori_ori_n514_));
  INV        o492(.A(ori_ori_n144_), .Y(ori_ori_n515_));
  AOI220     o493(.A0(ori_ori_n515_), .A1(ori_ori_n510_), .B0(ori_ori_n514_), .B1(ori_ori_n70_), .Y(ori_ori_n516_));
  NO2        o494(.A(ori_ori_n177_), .B(i_9_), .Y(ori_ori_n517_));
  NA2        o495(.A(ori_ori_n517_), .B(ori_ori_n502_), .Y(ori_ori_n518_));
  AOI210     o496(.A0(ori_ori_n518_), .A1(ori_ori_n309_), .B0(ori_ori_n138_), .Y(ori_ori_n519_));
  NAi32      o497(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n520_));
  NO2        o498(.A(ori_ori_n454_), .B(ori_ori_n520_), .Y(ori_ori_n521_));
  OR2        o499(.A(ori_ori_n521_), .B(ori_ori_n519_), .Y(ori_ori_n522_));
  BUFFER     o500(.A(ori_ori_n272_), .Y(ori_ori_n523_));
  NA3        o501(.A(ori_ori_n523_), .B(ori_ori_n126_), .C(ori_ori_n66_), .Y(ori_ori_n524_));
  AO210      o502(.A0(ori_ori_n300_), .A1(ori_ori_n478_), .B0(ori_ori_n36_), .Y(ori_ori_n525_));
  NA2        o503(.A(ori_ori_n525_), .B(ori_ori_n524_), .Y(ori_ori_n526_));
  INV        o504(.A(ori_ori_n509_), .Y(ori_ori_n527_));
  NA3        o505(.A(ori_ori_n239_), .B(ori_ori_n169_), .C(ori_ori_n126_), .Y(ori_ori_n528_));
  NA3        o506(.A(ori_ori_n528_), .B(ori_ori_n527_), .C(ori_ori_n363_), .Y(ori_ori_n529_));
  NA2        o507(.A(ori_ori_n272_), .B(ori_ori_n270_), .Y(ori_ori_n530_));
  NO2        o508(.A(ori_ori_n369_), .B(ori_ori_n94_), .Y(ori_ori_n531_));
  OAI210     o509(.A0(ori_ori_n531_), .A1(ori_ori_n77_), .B0(ori_ori_n253_), .Y(ori_ori_n532_));
  INV        o510(.A(ori_ori_n348_), .Y(ori_ori_n533_));
  NA3        o511(.A(ori_ori_n533_), .B(ori_ori_n206_), .C(i_7_), .Y(ori_ori_n534_));
  NA3        o512(.A(ori_ori_n534_), .B(ori_ori_n532_), .C(ori_ori_n530_), .Y(ori_ori_n535_));
  NO4        o513(.A(ori_ori_n535_), .B(ori_ori_n529_), .C(ori_ori_n526_), .D(ori_ori_n522_), .Y(ori_ori_n536_));
  NA4        o514(.A(ori_ori_n536_), .B(ori_ori_n516_), .C(ori_ori_n512_), .D(ori_ori_n240_), .Y(ori3));
  NA2        o515(.A(i_12_), .B(i_10_), .Y(ori_ori_n538_));
  NO2        o516(.A(i_11_), .B(ori_ori_n167_), .Y(ori_ori_n539_));
  NA3        o517(.A(ori_ori_n528_), .B(ori_ori_n363_), .C(ori_ori_n238_), .Y(ori_ori_n540_));
  NA2        o518(.A(ori_ori_n540_), .B(ori_ori_n38_), .Y(ori_ori_n541_));
  NOi21      o519(.An(ori_ori_n90_), .B(ori_ori_n484_), .Y(ori_ori_n542_));
  NO3        o520(.A(ori_ori_n384_), .B(ori_ori_n277_), .C(ori_ori_n113_), .Y(ori_ori_n543_));
  NA2        o521(.A(ori_ori_n255_), .B(ori_ori_n43_), .Y(ori_ori_n544_));
  AN2        o522(.A(ori_ori_n275_), .B(ori_ori_n52_), .Y(ori_ori_n545_));
  NO3        o523(.A(ori_ori_n545_), .B(ori_ori_n543_), .C(ori_ori_n542_), .Y(ori_ori_n546_));
  AOI210     o524(.A0(ori_ori_n546_), .A1(ori_ori_n541_), .B0(ori_ori_n46_), .Y(ori_ori_n547_));
  NA2        o525(.A(ori_ori_n138_), .B(ori_ori_n335_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n548_), .B(ori_ori_n60_), .Y(ori_ori_n549_));
  NOi21      o527(.An(i_5_), .B(i_9_), .Y(ori_ori_n550_));
  NA2        o528(.A(ori_ori_n550_), .B(ori_ori_n269_), .Y(ori_ori_n551_));
  BUFFER     o529(.A(ori_ori_n189_), .Y(ori_ori_n552_));
  AOI210     o530(.A0(ori_ori_n552_), .A1(ori_ori_n294_), .B0(ori_ori_n430_), .Y(ori_ori_n553_));
  NO2        o531(.A(ori_ori_n553_), .B(ori_ori_n551_), .Y(ori_ori_n554_));
  NO3        o532(.A(ori_ori_n554_), .B(ori_ori_n549_), .C(ori_ori_n547_), .Y(ori_ori_n555_));
  BUFFER     o533(.A(i_0_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n138_), .B(ori_ori_n24_), .Y(ori_ori_n557_));
  NO2        o535(.A(ori_ori_n417_), .B(ori_ori_n356_), .Y(ori_ori_n558_));
  NO2        o536(.A(ori_ori_n558_), .B(ori_ori_n557_), .Y(ori_ori_n559_));
  INV        o537(.A(ori_ori_n559_), .Y(ori_ori_n560_));
  NA2        o538(.A(ori_ori_n336_), .B(i_0_), .Y(ori_ori_n561_));
  NO3        o539(.A(ori_ori_n561_), .B(ori_ori_n243_), .C(ori_ori_n84_), .Y(ori_ori_n562_));
  NO4        o540(.A(ori_ori_n347_), .B(i_12_), .C(ori_ori_n257_), .D(ori_ori_n254_), .Y(ori_ori_n563_));
  AOI210     o541(.A0(ori_ori_n563_), .A1(i_11_), .B0(ori_ori_n562_), .Y(ori_ori_n564_));
  NA2        o542(.A(ori_ori_n476_), .B(ori_ori_n207_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n297_), .A1(ori_ori_n84_), .B0(ori_ori_n55_), .Y(ori_ori_n566_));
  NO2        o544(.A(ori_ori_n566_), .B(ori_ori_n565_), .Y(ori_ori_n567_));
  NO2        o545(.A(ori_ori_n179_), .B(ori_ori_n127_), .Y(ori_ori_n568_));
  NO4        o546(.A(ori_ori_n100_), .B(ori_ori_n55_), .C(ori_ori_n414_), .D(i_5_), .Y(ori_ori_n569_));
  AO220      o547(.A0(ori_ori_n569_), .A1(i_10_), .B0(ori_ori_n568_), .B1(i_6_), .Y(ori_ori_n570_));
  NO2        o548(.A(ori_ori_n570_), .B(ori_ori_n567_), .Y(ori_ori_n571_));
  NA3        o549(.A(ori_ori_n571_), .B(ori_ori_n564_), .C(ori_ori_n560_), .Y(ori_ori_n572_));
  NA2        o550(.A(i_11_), .B(i_9_), .Y(ori_ori_n573_));
  NO3        o551(.A(i_12_), .B(ori_ori_n573_), .C(ori_ori_n362_), .Y(ori_ori_n574_));
  AN2        o552(.A(ori_ori_n574_), .B(i_10_), .Y(ori_ori_n575_));
  NO2        o553(.A(ori_ori_n573_), .B(ori_ori_n70_), .Y(ori_ori_n576_));
  NO2        o554(.A(ori_ori_n136_), .B(i_0_), .Y(ori_ori_n577_));
  INV        o555(.A(ori_ori_n575_), .Y(ori_ori_n578_));
  NA2        o556(.A(ori_ori_n133_), .B(ori_ori_n95_), .Y(ori_ori_n579_));
  NA2        o557(.A(ori_ori_n364_), .B(ori_ori_n207_), .Y(ori_ori_n580_));
  NO2        o558(.A(ori_ori_n580_), .B(ori_ori_n544_), .Y(ori_ori_n581_));
  INV        o559(.A(ori_ori_n581_), .Y(ori_ori_n582_));
  NOi21      o560(.An(i_7_), .B(i_5_), .Y(ori_ori_n583_));
  NA2        o561(.A(ori_ori_n582_), .B(ori_ori_n578_), .Y(ori_ori_n584_));
  INV        o562(.A(ori_ori_n538_), .Y(ori_ori_n585_));
  OA210      o563(.A0(ori_ori_n293_), .A1(ori_ori_n162_), .B0(ori_ori_n292_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n585_), .B(ori_ori_n576_), .Y(ori_ori_n587_));
  NA2        o565(.A(ori_ori_n576_), .B(ori_ori_n200_), .Y(ori_ori_n588_));
  INV        o566(.A(ori_ori_n588_), .Y(ori_ori_n589_));
  NA2        o567(.A(ori_ori_n589_), .B(ori_ori_n293_), .Y(ori_ori_n590_));
  NO3        o568(.A(ori_ori_n347_), .B(ori_ori_n222_), .C(ori_ori_n24_), .Y(ori_ori_n591_));
  AOI210     o569(.A0(ori_ori_n439_), .A1(ori_ori_n320_), .B0(ori_ori_n591_), .Y(ori_ori_n592_));
  NAi21      o570(.An(i_9_), .B(i_5_), .Y(ori_ori_n593_));
  NO2        o571(.A(ori_ori_n593_), .B(ori_ori_n249_), .Y(ori_ori_n594_));
  NA2        o572(.A(ori_ori_n594_), .B(ori_ori_n376_), .Y(ori_ori_n595_));
  OAI220     o573(.A0(ori_ori_n595_), .A1(ori_ori_n83_), .B0(ori_ori_n592_), .B1(ori_ori_n134_), .Y(ori_ori_n596_));
  NO2        o574(.A(ori_ori_n596_), .B(ori_ori_n312_), .Y(ori_ori_n597_));
  NA3        o575(.A(ori_ori_n597_), .B(ori_ori_n590_), .C(ori_ori_n587_), .Y(ori_ori_n598_));
  NO3        o576(.A(ori_ori_n598_), .B(ori_ori_n584_), .C(ori_ori_n572_), .Y(ori_ori_n599_));
  NO2        o577(.A(ori_ori_n556_), .B(ori_ori_n459_), .Y(ori_ori_n600_));
  AOI210     o578(.A0(ori_ori_n513_), .A1(ori_ori_n429_), .B0(ori_ori_n579_), .Y(ori_ori_n601_));
  INV        o579(.A(ori_ori_n601_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n173_), .B(ori_ori_n165_), .Y(ori_ori_n603_));
  AOI210     o581(.A0(ori_ori_n603_), .A1(ori_ori_n561_), .B0(ori_ori_n127_), .Y(ori_ori_n604_));
  INV        o582(.A(ori_ori_n604_), .Y(ori_ori_n605_));
  NA2        o583(.A(ori_ori_n605_), .B(ori_ori_n602_), .Y(ori_ori_n606_));
  NO3        o584(.A(ori_ori_n153_), .B(ori_ori_n242_), .C(i_0_), .Y(ori_ori_n607_));
  OAI210     o585(.A0(ori_ori_n607_), .A1(ori_ori_n73_), .B0(i_13_), .Y(ori_ori_n608_));
  INV        o586(.A(ori_ori_n608_), .Y(ori_ori_n609_));
  NO2        o587(.A(ori_ori_n172_), .B(ori_ori_n88_), .Y(ori_ori_n610_));
  AOI210     o588(.A0(ori_ori_n610_), .A1(ori_ori_n600_), .B0(ori_ori_n98_), .Y(ori_ori_n611_));
  OR2        o589(.A(ori_ori_n611_), .B(i_5_), .Y(ori_ori_n612_));
  AOI210     o590(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n136_), .Y(ori_ori_n613_));
  NA2        o591(.A(ori_ori_n613_), .B(ori_ori_n586_), .Y(ori_ori_n614_));
  NO3        o592(.A(ori_ori_n544_), .B(ori_ori_n51_), .C(ori_ori_n46_), .Y(ori_ori_n615_));
  NO3        o593(.A(ori_ori_n659_), .B(ori_ori_n615_), .C(ori_ori_n656_), .Y(ori_ori_n616_));
  NO3        o594(.A(ori_ori_n573_), .B(ori_ori_n158_), .C(ori_ori_n141_), .Y(ori_ori_n617_));
  INV        o595(.A(ori_ori_n617_), .Y(ori_ori_n618_));
  NA4        o596(.A(ori_ori_n618_), .B(ori_ori_n616_), .C(ori_ori_n614_), .D(ori_ori_n612_), .Y(ori_ori_n619_));
  NO2        o597(.A(ori_ori_n83_), .B(i_5_), .Y(ori_ori_n620_));
  NA3        o598(.A(ori_ori_n539_), .B(ori_ori_n99_), .C(ori_ori_n108_), .Y(ori_ori_n621_));
  INV        o599(.A(ori_ori_n621_), .Y(ori_ori_n622_));
  NA2        o600(.A(ori_ori_n622_), .B(ori_ori_n620_), .Y(ori_ori_n623_));
  NAi21      o601(.An(ori_ori_n171_), .B(ori_ori_n172_), .Y(ori_ori_n624_));
  NO4        o602(.A(ori_ori_n170_), .B(ori_ori_n153_), .C(i_0_), .D(i_12_), .Y(ori_ori_n625_));
  AOI220     o603(.A0(ori_ori_n625_), .A1(ori_ori_n624_), .B0(ori_ori_n508_), .B1(ori_ori_n137_), .Y(ori_ori_n626_));
  NA2        o604(.A(ori_ori_n583_), .B(ori_ori_n291_), .Y(ori_ori_n627_));
  NO2        o605(.A(ori_ori_n627_), .B(ori_ori_n420_), .Y(ori_ori_n628_));
  NA2        o606(.A(ori_ori_n628_), .B(ori_ori_n577_), .Y(ori_ori_n629_));
  NA3        o607(.A(ori_ori_n629_), .B(ori_ori_n626_), .C(ori_ori_n623_), .Y(ori_ori_n630_));
  NO4        o608(.A(ori_ori_n630_), .B(ori_ori_n619_), .C(ori_ori_n609_), .D(ori_ori_n606_), .Y(ori_ori_n631_));
  INV        o609(.A(ori_ori_n368_), .Y(ori_ori_n632_));
  NA2        o610(.A(ori_ori_n632_), .B(ori_ori_n151_), .Y(ori_ori_n633_));
  BUFFER     o611(.A(i_7_), .Y(ori_ori_n634_));
  NA2        o612(.A(ori_ori_n139_), .B(ori_ori_n140_), .Y(ori_ori_n635_));
  AO210      o613(.A0(ori_ori_n634_), .A1(ori_ori_n33_), .B0(ori_ori_n635_), .Y(ori_ori_n636_));
  NAi31      o614(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n637_));
  NO2        o615(.A(ori_ori_n67_), .B(ori_ori_n637_), .Y(ori_ori_n638_));
  NO2        o616(.A(ori_ori_n638_), .B(ori_ori_n397_), .Y(ori_ori_n639_));
  NA2        o617(.A(ori_ori_n639_), .B(ori_ori_n636_), .Y(ori_ori_n640_));
  AOI210     o618(.A0(ori_ori_n640_), .A1(ori_ori_n46_), .B0(ori_ori_n563_), .Y(ori_ori_n641_));
  AOI210     o619(.A0(ori_ori_n641_), .A1(ori_ori_n633_), .B0(ori_ori_n70_), .Y(ori_ori_n642_));
  NO3        o620(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(i_4_), .Y(ori_ori_n643_));
  OAI210     o621(.A0(ori_ori_n662_), .A1(ori_ori_n201_), .B0(ori_ori_n643_), .Y(ori_ori_n644_));
  NO2        o622(.A(ori_ori_n644_), .B(ori_ori_n459_), .Y(ori_ori_n645_));
  NO4        o623(.A(ori_ori_n593_), .B(i_11_), .C(ori_ori_n178_), .D(ori_ori_n177_), .Y(ori_ori_n646_));
  NO2        o624(.A(ori_ori_n646_), .B(ori_ori_n334_), .Y(ori_ori_n647_));
  INV        o625(.A(ori_ori_n228_), .Y(ori_ori_n648_));
  AOI210     o626(.A0(ori_ori_n648_), .A1(ori_ori_n647_), .B0(ori_ori_n39_), .Y(ori_ori_n649_));
  NO2        o627(.A(ori_ori_n649_), .B(ori_ori_n645_), .Y(ori_ori_n650_));
  INV        o628(.A(ori_ori_n650_), .Y(ori_ori_n651_));
  NO2        o629(.A(ori_ori_n651_), .B(ori_ori_n642_), .Y(ori_ori_n652_));
  NA4        o630(.A(ori_ori_n652_), .B(ori_ori_n631_), .C(ori_ori_n599_), .D(ori_ori_n555_), .Y(ori4));
  INV        o631(.A(ori_ori_n319_), .Y(ori_ori_n656_));
  INV        o632(.A(i_6_), .Y(ori_ori_n657_));
  INV        o633(.A(ori_ori_n319_), .Y(ori_ori_n658_));
  INV        o634(.A(ori_ori_n298_), .Y(ori_ori_n659_));
  INV        o635(.A(ori_ori_n450_), .Y(ori_ori_n660_));
  INV        o636(.A(i_8_), .Y(ori_ori_n661_));
  INV        o637(.A(i_0_), .Y(ori_ori_n662_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NO2        m028(.A(mai_mai_n47_), .B(mai_mai_n46_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_0_), .B(i_2_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_7_), .B(i_9_), .Y(mai_mai_n53_));
  NA2        m031(.A(mai_mai_n51_), .B(mai_mai_n45_), .Y(mai_mai_n54_));
  NA3        m032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n55_));
  NO2        m033(.A(i_1_), .B(i_6_), .Y(mai_mai_n56_));
  NA2        m034(.A(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  OAI210     m035(.A0(mai_mai_n57_), .A1(mai_mai_n56_), .B0(mai_mai_n55_), .Y(mai_mai_n58_));
  NA2        m036(.A(mai_mai_n58_), .B(i_12_), .Y(mai_mai_n59_));
  NAi21      m037(.An(i_2_), .B(i_7_), .Y(mai_mai_n60_));
  INV        m038(.A(i_1_), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n61_), .B(i_6_), .Y(mai_mai_n62_));
  NA3        m040(.A(mai_mai_n62_), .B(mai_mai_n60_), .C(mai_mai_n31_), .Y(mai_mai_n63_));
  NA2        m041(.A(i_1_), .B(i_10_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NAi31      m043(.An(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n59_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n67_));
  AOI210     m045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n68_));
  NA2        m046(.A(i_1_), .B(i_6_), .Y(mai_mai_n69_));
  NO2        m047(.A(mai_mai_n69_), .B(mai_mai_n25_), .Y(mai_mai_n70_));
  INV        m048(.A(i_0_), .Y(mai_mai_n71_));
  NAi21      m049(.An(i_5_), .B(i_10_), .Y(mai_mai_n72_));
  NA2        m050(.A(i_5_), .B(i_9_), .Y(mai_mai_n73_));
  AOI210     m051(.A0(mai_mai_n73_), .A1(mai_mai_n72_), .B0(mai_mai_n71_), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n74_), .B(mai_mai_n70_), .Y(mai_mai_n75_));
  INV        m053(.A(mai_mai_n75_), .Y(mai_mai_n76_));
  OAI210     m054(.A0(mai_mai_n76_), .A1(mai_mai_n66_), .B0(i_0_), .Y(mai_mai_n77_));
  NA2        m055(.A(i_12_), .B(i_5_), .Y(mai_mai_n78_));
  NA2        m056(.A(i_2_), .B(i_8_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_3_), .B(i_9_), .Y(mai_mai_n80_));
  NO2        m058(.A(i_3_), .B(i_7_), .Y(mai_mai_n81_));
  INV        m059(.A(i_6_), .Y(mai_mai_n82_));
  OR4        m060(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n83_));
  INV        m061(.A(mai_mai_n83_), .Y(mai_mai_n84_));
  NO2        m062(.A(i_2_), .B(i_7_), .Y(mai_mai_n85_));
  NO2        m063(.A(mai_mai_n84_), .B(mai_mai_n85_), .Y(mai_mai_n86_));
  NA2        m064(.A(i_1_), .B(mai_mai_n86_), .Y(mai_mai_n87_));
  NAi21      m065(.An(i_6_), .B(i_10_), .Y(mai_mai_n88_));
  NA2        m066(.A(i_6_), .B(i_9_), .Y(mai_mai_n89_));
  AOI210     m067(.A0(mai_mai_n89_), .A1(mai_mai_n88_), .B0(mai_mai_n61_), .Y(mai_mai_n90_));
  NA2        m068(.A(i_2_), .B(i_6_), .Y(mai_mai_n91_));
  INV        m069(.A(mai_mai_n90_), .Y(mai_mai_n92_));
  AOI210     m070(.A0(mai_mai_n92_), .A1(mai_mai_n87_), .B0(mai_mai_n78_), .Y(mai_mai_n93_));
  AN3        m071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n94_));
  NAi21      m072(.An(i_6_), .B(i_11_), .Y(mai_mai_n95_));
  NO2        m073(.A(i_5_), .B(i_8_), .Y(mai_mai_n96_));
  NOi21      m074(.An(mai_mai_n96_), .B(mai_mai_n95_), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n97_), .B(mai_mai_n60_), .Y(mai_mai_n98_));
  INV        m076(.A(i_7_), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n46_), .B(mai_mai_n99_), .Y(mai_mai_n100_));
  NO2        m078(.A(i_0_), .B(i_5_), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n101_), .B(mai_mai_n82_), .Y(mai_mai_n102_));
  NA2        m080(.A(i_12_), .B(i_3_), .Y(mai_mai_n103_));
  INV        m081(.A(mai_mai_n103_), .Y(mai_mai_n104_));
  NA3        m082(.A(mai_mai_n104_), .B(mai_mai_n102_), .C(mai_mai_n100_), .Y(mai_mai_n105_));
  NAi21      m083(.An(i_7_), .B(i_11_), .Y(mai_mai_n106_));
  AN2        m084(.A(i_2_), .B(i_10_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(i_7_), .Y(mai_mai_n108_));
  OR2        m086(.A(mai_mai_n78_), .B(mai_mai_n56_), .Y(mai_mai_n109_));
  NO2        m087(.A(i_8_), .B(mai_mai_n99_), .Y(mai_mai_n110_));
  NO3        m088(.A(mai_mai_n110_), .B(mai_mai_n109_), .C(mai_mai_n108_), .Y(mai_mai_n111_));
  NA2        m089(.A(i_12_), .B(i_7_), .Y(mai_mai_n112_));
  NA2        m090(.A(i_11_), .B(i_12_), .Y(mai_mai_n113_));
  INV        m091(.A(mai_mai_n113_), .Y(mai_mai_n114_));
  NO2        m092(.A(mai_mai_n114_), .B(mai_mai_n111_), .Y(mai_mai_n115_));
  NA3        m093(.A(mai_mai_n115_), .B(mai_mai_n105_), .C(mai_mai_n98_), .Y(mai_mai_n116_));
  NOi21      m094(.An(i_1_), .B(i_5_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(i_11_), .Y(mai_mai_n118_));
  NA2        m096(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(i_10_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(mai_mai_n46_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n122_));
  NAi21      m100(.An(i_3_), .B(i_8_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(mai_mai_n60_), .Y(mai_mai_n124_));
  NOi31      m102(.An(mai_mai_n124_), .B(mai_mai_n122_), .C(mai_mai_n121_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_1_), .B(mai_mai_n82_), .Y(mai_mai_n126_));
  NO2        m104(.A(i_6_), .B(i_5_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(i_3_), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n125_), .B(mai_mai_n118_), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n116_), .C(mai_mai_n93_), .Y(mai_mai_n130_));
  NA3        m108(.A(mai_mai_n130_), .B(mai_mai_n77_), .C(mai_mai_n54_), .Y(mai2));
  NO2        m109(.A(mai_mai_n61_), .B(mai_mai_n37_), .Y(mai_mai_n132_));
  NA2        m110(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NA4        m112(.A(mai_mai_n134_), .B(mai_mai_n75_), .C(mai_mai_n67_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m113(.A(i_8_), .B(i_7_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n136_), .B(i_6_), .Y(mai_mai_n137_));
  NO2        m115(.A(i_12_), .B(i_13_), .Y(mai_mai_n138_));
  NAi21      m116(.An(i_5_), .B(i_11_), .Y(mai_mai_n139_));
  NOi21      m117(.An(mai_mai_n138_), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m118(.A(i_0_), .B(i_1_), .Y(mai_mai_n141_));
  NA2        m119(.A(i_2_), .B(i_3_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n142_), .B(i_4_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(mai_mai_n140_), .Y(mai_mai_n144_));
  AN2        m122(.A(mai_mai_n138_), .B(mai_mai_n80_), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n145_), .B(mai_mai_n27_), .Y(mai_mai_n146_));
  NA2        m124(.A(i_1_), .B(i_5_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n71_), .B(mai_mai_n46_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n150_));
  OR2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n78_), .C(i_13_), .Y(mai_mai_n152_));
  NAi32      m130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n153_));
  NAi21      m131(.An(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m132(.An(i_4_), .B(i_10_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NO2        m134(.A(i_3_), .B(i_5_), .Y(mai_mai_n157_));
  NO3        m135(.A(mai_mai_n71_), .B(i_2_), .C(i_1_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n154_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(mai_mai_n150_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(mai_mai_n161_), .A1(mai_mai_n144_), .B0(mai_mai_n137_), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n163_));
  NOi21      m141(.An(i_4_), .B(i_9_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_11_), .B(i_13_), .Y(mai_mai_n165_));
  NA2        m143(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  BUFFER     m144(.A(mai_mai_n166_), .Y(mai_mai_n167_));
  NO2        m145(.A(i_4_), .B(i_5_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_12_), .B(i_11_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(i_13_), .Y(mai_mai_n170_));
  NA3        m148(.A(mai_mai_n170_), .B(mai_mai_n168_), .C(mai_mai_n80_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n167_), .B0(mai_mai_n163_), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n71_), .B(mai_mai_n61_), .Y(mai_mai_n173_));
  INV        m151(.A(mai_mai_n173_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n175_));
  NAi31      m153(.An(mai_mai_n175_), .B(mai_mai_n145_), .C(i_11_), .Y(mai_mai_n176_));
  NA2        m154(.A(i_3_), .B(i_5_), .Y(mai_mai_n177_));
  NO2        m155(.A(mai_mai_n176_), .B(mai_mai_n174_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n71_), .B(i_5_), .Y(mai_mai_n179_));
  NO2        m157(.A(i_13_), .B(i_10_), .Y(mai_mai_n180_));
  NA3        m158(.A(mai_mai_n180_), .B(mai_mai_n179_), .C(mai_mai_n44_), .Y(mai_mai_n181_));
  NO2        m159(.A(i_2_), .B(i_1_), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n182_), .B(i_3_), .Y(mai_mai_n183_));
  NAi21      m161(.An(i_4_), .B(i_12_), .Y(mai_mai_n184_));
  NO3        m162(.A(mai_mai_n184_), .B(mai_mai_n183_), .C(mai_mai_n181_), .Y(mai_mai_n185_));
  NO3        m163(.A(mai_mai_n185_), .B(mai_mai_n178_), .C(mai_mai_n172_), .Y(mai_mai_n186_));
  INV        m164(.A(i_8_), .Y(mai_mai_n187_));
  NA2        m165(.A(i_8_), .B(i_6_), .Y(mai_mai_n188_));
  NO3        m166(.A(i_3_), .B(mai_mai_n82_), .C(mai_mai_n48_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n110_), .Y(mai_mai_n190_));
  NO3        m168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n191_));
  NA3        m169(.A(mai_mai_n191_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n192_));
  NO3        m170(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n193_));
  INV        m171(.A(mai_mai_n193_), .Y(mai_mai_n194_));
  AOI210     m172(.A0(mai_mai_n194_), .A1(mai_mai_n192_), .B0(mai_mai_n190_), .Y(mai_mai_n195_));
  NO2        m173(.A(i_3_), .B(i_8_), .Y(mai_mai_n196_));
  NO3        m174(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n197_));
  NO2        m175(.A(i_13_), .B(i_9_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n198_), .B(i_6_), .Y(mai_mai_n199_));
  NAi21      m177(.An(i_12_), .B(i_3_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n201_));
  NO3        m179(.A(i_0_), .B(i_2_), .C(mai_mai_n61_), .Y(mai_mai_n202_));
  INV        m180(.A(mai_mai_n195_), .Y(mai_mai_n203_));
  OAI220     m181(.A0(mai_mai_n203_), .A1(i_4_), .B0(mai_mai_n188_), .B1(mai_mai_n186_), .Y(mai_mai_n204_));
  NA3        m182(.A(i_13_), .B(mai_mai_n187_), .C(i_10_), .Y(mai_mai_n205_));
  NO2        m183(.A(mai_mai_n205_), .B(i_12_), .Y(mai_mai_n206_));
  NA2        m184(.A(i_0_), .B(i_5_), .Y(mai_mai_n207_));
  NA2        m185(.A(mai_mai_n207_), .B(mai_mai_n102_), .Y(mai_mai_n208_));
  OAI220     m186(.A0(mai_mai_n208_), .A1(mai_mai_n183_), .B0(mai_mai_n174_), .B1(mai_mai_n128_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n71_), .B(mai_mai_n26_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n46_), .B(mai_mai_n61_), .Y(mai_mai_n212_));
  NA3        m190(.A(mai_mai_n212_), .B(mai_mai_n211_), .C(mai_mai_n210_), .Y(mai_mai_n213_));
  INV        m191(.A(i_13_), .Y(mai_mai_n214_));
  NO2        m192(.A(i_12_), .B(mai_mai_n214_), .Y(mai_mai_n215_));
  NA3        m193(.A(mai_mai_n215_), .B(mai_mai_n191_), .C(mai_mai_n189_), .Y(mai_mai_n216_));
  OAI210     m194(.A0(mai_mai_n213_), .A1(i_9_), .B0(mai_mai_n216_), .Y(mai_mai_n217_));
  AOI220     m195(.A0(mai_mai_n217_), .A1(mai_mai_n136_), .B0(mai_mai_n209_), .B1(mai_mai_n206_), .Y(mai_mai_n218_));
  NO2        m196(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n219_));
  NA2        m197(.A(mai_mai_n219_), .B(mai_mai_n934_), .Y(mai_mai_n220_));
  OR2        m198(.A(i_8_), .B(i_7_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n52_), .B(i_1_), .Y(mai_mai_n222_));
  NA2        m200(.A(mai_mai_n222_), .B(i_6_), .Y(mai_mai_n223_));
  INV        m201(.A(i_12_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n44_), .B(mai_mai_n224_), .Y(mai_mai_n225_));
  NO3        m203(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n226_));
  NA2        m204(.A(i_2_), .B(i_1_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n223_), .B(mai_mai_n220_), .Y(mai_mai_n228_));
  NAi21      m206(.An(i_4_), .B(i_3_), .Y(mai_mai_n229_));
  NO2        m207(.A(mai_mai_n229_), .B(mai_mai_n73_), .Y(mai_mai_n230_));
  NO2        m208(.A(i_0_), .B(i_6_), .Y(mai_mai_n231_));
  NOi41      m209(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n232_));
  NA2        m210(.A(mai_mai_n232_), .B(mai_mai_n231_), .Y(mai_mai_n233_));
  AOI210     m211(.A0(mai_mai_n932_), .A1(mai_mai_n40_), .B0(mai_mai_n228_), .Y(mai_mai_n234_));
  NO2        m212(.A(i_11_), .B(mai_mai_n214_), .Y(mai_mai_n235_));
  NOi21      m213(.An(i_1_), .B(i_6_), .Y(mai_mai_n236_));
  NAi21      m214(.An(i_3_), .B(i_7_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n224_), .B(i_9_), .Y(mai_mai_n238_));
  OR4        m216(.A(mai_mai_n238_), .B(mai_mai_n237_), .C(mai_mai_n236_), .D(mai_mai_n179_), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n48_), .B(mai_mai_n25_), .Y(mai_mai_n240_));
  NO2        m218(.A(i_12_), .B(i_3_), .Y(mai_mai_n241_));
  NA2        m219(.A(mai_mai_n71_), .B(i_5_), .Y(mai_mai_n242_));
  NA2        m220(.A(i_3_), .B(i_9_), .Y(mai_mai_n243_));
  NAi21      m221(.An(i_7_), .B(i_10_), .Y(mai_mai_n244_));
  NO2        m222(.A(mai_mai_n244_), .B(mai_mai_n243_), .Y(mai_mai_n245_));
  NA3        m223(.A(mai_mai_n245_), .B(mai_mai_n242_), .C(mai_mai_n62_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n246_), .B(mai_mai_n239_), .Y(mai_mai_n247_));
  NA3        m225(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n248_));
  INV        m226(.A(mai_mai_n137_), .Y(mai_mai_n249_));
  NA2        m227(.A(mai_mai_n224_), .B(i_13_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n250_), .B(mai_mai_n73_), .Y(mai_mai_n251_));
  AOI220     m229(.A0(mai_mai_n251_), .A1(mai_mai_n249_), .B0(mai_mai_n247_), .B1(mai_mai_n235_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n221_), .B(mai_mai_n37_), .Y(mai_mai_n253_));
  NA2        m231(.A(i_12_), .B(i_6_), .Y(mai_mai_n254_));
  NO3        m232(.A(i_9_), .B(mai_mai_n254_), .C(mai_mai_n48_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n229_), .B(i_2_), .Y(mai_mai_n256_));
  NA2        m234(.A(mai_mai_n235_), .B(i_9_), .Y(mai_mai_n257_));
  NA2        m235(.A(mai_mai_n148_), .B(mai_mai_n61_), .Y(mai_mai_n258_));
  NO2        m236(.A(mai_mai_n237_), .B(i_8_), .Y(mai_mai_n259_));
  NO2        m237(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n260_));
  NA3        m238(.A(mai_mai_n260_), .B(mai_mai_n259_), .C(i_9_), .Y(mai_mai_n261_));
  NA3        m239(.A(i_6_), .B(mai_mai_n253_), .C(mai_mai_n215_), .Y(mai_mai_n262_));
  AOI210     m240(.A0(mai_mai_n262_), .A1(mai_mai_n261_), .B0(mai_mai_n258_), .Y(mai_mai_n263_));
  INV        m241(.A(mai_mai_n263_), .Y(mai_mai_n264_));
  NA4        m242(.A(mai_mai_n264_), .B(mai_mai_n252_), .C(mai_mai_n234_), .D(mai_mai_n218_), .Y(mai_mai_n265_));
  NO3        m243(.A(i_12_), .B(mai_mai_n214_), .C(mai_mai_n37_), .Y(mai_mai_n266_));
  INV        m244(.A(mai_mai_n266_), .Y(mai_mai_n267_));
  NA2        m245(.A(i_8_), .B(mai_mai_n99_), .Y(mai_mai_n268_));
  NO3        m246(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n269_));
  AOI220     m247(.A0(mai_mai_n269_), .A1(mai_mai_n189_), .B0(i_6_), .B1(mai_mai_n222_), .Y(mai_mai_n270_));
  NO2        m248(.A(mai_mai_n270_), .B(mai_mai_n268_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n227_), .B(i_0_), .Y(mai_mai_n272_));
  AOI220     m250(.A0(mai_mai_n272_), .A1(i_8_), .B0(i_1_), .B1(mai_mai_n136_), .Y(mai_mai_n273_));
  NA2        m251(.A(mai_mai_n260_), .B(mai_mai_n26_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n274_), .B(mai_mai_n273_), .Y(mai_mai_n275_));
  NA2        m253(.A(i_0_), .B(i_1_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(i_2_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n57_), .B(i_6_), .Y(mai_mai_n278_));
  NA3        m256(.A(mai_mai_n278_), .B(mai_mai_n277_), .C(mai_mai_n157_), .Y(mai_mai_n279_));
  OAI210     m257(.A0(mai_mai_n159_), .A1(mai_mai_n137_), .B0(mai_mai_n279_), .Y(mai_mai_n280_));
  NO3        m258(.A(mai_mai_n280_), .B(mai_mai_n275_), .C(mai_mai_n271_), .Y(mai_mai_n281_));
  NO2        m259(.A(i_3_), .B(i_10_), .Y(mai_mai_n282_));
  NA3        m260(.A(mai_mai_n282_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n283_));
  NA2        m261(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n284_));
  NO2        m262(.A(mai_mai_n284_), .B(i_8_), .Y(mai_mai_n285_));
  NA2        m263(.A(mai_mai_n285_), .B(i_7_), .Y(mai_mai_n286_));
  AN2        m264(.A(i_3_), .B(i_10_), .Y(mai_mai_n287_));
  NA3        m265(.A(mai_mai_n287_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n288_));
  NO2        m266(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n289_));
  NO2        m267(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n290_));
  OR2        m268(.A(mai_mai_n286_), .B(mai_mai_n283_), .Y(mai_mai_n291_));
  OAI220     m269(.A0(mai_mai_n291_), .A1(i_6_), .B0(mai_mai_n281_), .B1(mai_mai_n267_), .Y(mai_mai_n292_));
  NO4        m270(.A(mai_mai_n292_), .B(mai_mai_n265_), .C(mai_mai_n204_), .D(mai_mai_n162_), .Y(mai_mai_n293_));
  NO3        m271(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n57_), .B(mai_mai_n82_), .Y(mai_mai_n295_));
  NA2        m273(.A(mai_mai_n272_), .B(mai_mai_n295_), .Y(mai_mai_n296_));
  NO3        m274(.A(i_6_), .B(mai_mai_n187_), .C(i_7_), .Y(mai_mai_n297_));
  NA2        m275(.A(mai_mai_n297_), .B(mai_mai_n191_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n298_), .B(mai_mai_n296_), .Y(mai_mai_n299_));
  NO2        m277(.A(i_2_), .B(i_3_), .Y(mai_mai_n300_));
  OR2        m278(.A(i_0_), .B(i_5_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n207_), .B(mai_mai_n301_), .Y(mai_mai_n302_));
  NA4        m280(.A(mai_mai_n302_), .B(i_6_), .C(mai_mai_n300_), .D(i_1_), .Y(mai_mai_n303_));
  NA3        m281(.A(mai_mai_n272_), .B(i_6_), .C(mai_mai_n110_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n151_), .B(mai_mai_n46_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n305_), .B(i_7_), .C(mai_mai_n157_), .Y(mai_mai_n306_));
  NA3        m284(.A(mai_mai_n306_), .B(mai_mai_n304_), .C(mai_mai_n303_), .Y(mai_mai_n307_));
  OAI210     m285(.A0(mai_mai_n307_), .A1(mai_mai_n299_), .B0(i_4_), .Y(mai_mai_n308_));
  NO2        m286(.A(i_12_), .B(i_10_), .Y(mai_mai_n309_));
  NOi21      m287(.An(i_5_), .B(i_0_), .Y(mai_mai_n310_));
  NO3        m288(.A(mai_mai_n284_), .B(mai_mai_n310_), .C(mai_mai_n123_), .Y(mai_mai_n311_));
  NA4        m289(.A(mai_mai_n81_), .B(mai_mai_n36_), .C(mai_mai_n82_), .D(i_8_), .Y(mai_mai_n312_));
  NA2        m290(.A(mai_mai_n311_), .B(mai_mai_n309_), .Y(mai_mai_n313_));
  NO2        m291(.A(i_6_), .B(i_8_), .Y(mai_mai_n314_));
  NOi21      m292(.An(i_0_), .B(i_2_), .Y(mai_mai_n315_));
  AN2        m293(.A(mai_mai_n315_), .B(mai_mai_n314_), .Y(mai_mai_n316_));
  NO2        m294(.A(i_1_), .B(i_7_), .Y(mai_mai_n317_));
  AO220      m295(.A0(mai_mai_n317_), .A1(mai_mai_n316_), .B0(i_7_), .B1(mai_mai_n222_), .Y(mai_mai_n318_));
  NA3        m296(.A(mai_mai_n318_), .B(i_4_), .C(i_5_), .Y(mai_mai_n319_));
  NA3        m297(.A(mai_mai_n319_), .B(mai_mai_n313_), .C(mai_mai_n308_), .Y(mai_mai_n320_));
  NO3        m298(.A(mai_mai_n221_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n321_));
  OAI210     m299(.A0(i_7_), .A1(mai_mai_n321_), .B0(i_6_), .Y(mai_mai_n322_));
  AOI210     m300(.A0(mai_mai_n99_), .A1(mai_mai_n322_), .B0(mai_mai_n302_), .Y(mai_mai_n323_));
  NOi21      m301(.An(mai_mai_n147_), .B(mai_mai_n102_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n324_), .B(mai_mai_n119_), .Y(mai_mai_n325_));
  OAI210     m303(.A0(mai_mai_n325_), .A1(mai_mai_n323_), .B0(i_3_), .Y(mai_mai_n326_));
  INV        m304(.A(mai_mai_n81_), .Y(mai_mai_n327_));
  NO2        m305(.A(mai_mai_n276_), .B(mai_mai_n79_), .Y(mai_mai_n328_));
  INV        m306(.A(mai_mai_n328_), .Y(mai_mai_n329_));
  NO2        m307(.A(mai_mai_n91_), .B(mai_mai_n187_), .Y(mai_mai_n330_));
  NA2        m308(.A(mai_mai_n330_), .B(mai_mai_n61_), .Y(mai_mai_n331_));
  AOI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n329_), .B0(mai_mai_n327_), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n187_), .B(i_9_), .Y(mai_mai_n333_));
  NO2        m311(.A(mai_mai_n332_), .B(mai_mai_n275_), .Y(mai_mai_n334_));
  AOI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n326_), .B0(mai_mai_n156_), .Y(mai_mai_n335_));
  AOI210     m313(.A0(mai_mai_n320_), .A1(mai_mai_n294_), .B0(mai_mai_n335_), .Y(mai_mai_n336_));
  NOi32      m314(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n337_));
  INV        m315(.A(mai_mai_n337_), .Y(mai_mai_n338_));
  NAi21      m316(.An(i_0_), .B(i_6_), .Y(mai_mai_n339_));
  NAi21      m317(.An(i_1_), .B(i_5_), .Y(mai_mai_n340_));
  NA2        m318(.A(mai_mai_n340_), .B(mai_mai_n339_), .Y(mai_mai_n341_));
  NA2        m319(.A(mai_mai_n341_), .B(mai_mai_n25_), .Y(mai_mai_n342_));
  NO2        m320(.A(mai_mai_n342_), .B(mai_mai_n153_), .Y(mai_mai_n343_));
  NAi41      m321(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n344_));
  AOI210     m322(.A0(mai_mai_n344_), .A1(mai_mai_n153_), .B0(mai_mai_n151_), .Y(mai_mai_n345_));
  NOi32      m323(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n346_));
  NO2        m324(.A(i_1_), .B(mai_mai_n99_), .Y(mai_mai_n347_));
  NAi21      m325(.An(i_3_), .B(i_4_), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(i_9_), .Y(mai_mai_n349_));
  AN2        m327(.A(i_6_), .B(i_7_), .Y(mai_mai_n350_));
  OAI210     m328(.A0(mai_mai_n350_), .A1(mai_mai_n347_), .B0(mai_mai_n349_), .Y(mai_mai_n351_));
  NA2        m329(.A(i_2_), .B(i_7_), .Y(mai_mai_n352_));
  NO2        m330(.A(mai_mai_n348_), .B(i_10_), .Y(mai_mai_n353_));
  NA3        m331(.A(mai_mai_n353_), .B(mai_mai_n352_), .C(mai_mai_n231_), .Y(mai_mai_n354_));
  AOI210     m332(.A0(mai_mai_n354_), .A1(mai_mai_n351_), .B0(mai_mai_n179_), .Y(mai_mai_n355_));
  AOI210     m333(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n356_), .A1(mai_mai_n182_), .B0(mai_mai_n353_), .Y(mai_mai_n357_));
  AOI220     m335(.A0(mai_mai_n353_), .A1(mai_mai_n317_), .B0(mai_mai_n226_), .B1(mai_mai_n182_), .Y(mai_mai_n358_));
  AOI210     m336(.A0(mai_mai_n358_), .A1(mai_mai_n357_), .B0(i_5_), .Y(mai_mai_n359_));
  NO4        m337(.A(mai_mai_n359_), .B(mai_mai_n355_), .C(mai_mai_n345_), .D(mai_mai_n343_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n360_), .B(mai_mai_n338_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n57_), .B(mai_mai_n25_), .Y(mai_mai_n362_));
  AN2        m340(.A(i_12_), .B(i_5_), .Y(mai_mai_n363_));
  NA2        m341(.A(mai_mai_n937_), .B(mai_mai_n363_), .Y(mai_mai_n364_));
  NO2        m342(.A(i_11_), .B(i_6_), .Y(mai_mai_n365_));
  NA3        m343(.A(mai_mai_n365_), .B(mai_mai_n305_), .C(mai_mai_n214_), .Y(mai_mai_n366_));
  NO2        m344(.A(mai_mai_n366_), .B(mai_mai_n364_), .Y(mai_mai_n367_));
  NO2        m345(.A(i_5_), .B(i_10_), .Y(mai_mai_n368_));
  NA2        m346(.A(mai_mai_n138_), .B(mai_mai_n45_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n369_), .B(mai_mai_n229_), .Y(mai_mai_n370_));
  OAI210     m348(.A0(mai_mai_n370_), .A1(mai_mai_n367_), .B0(mai_mai_n362_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n372_));
  NA2        m350(.A(mai_mai_n367_), .B(mai_mai_n372_), .Y(mai_mai_n373_));
  NO3        m351(.A(mai_mai_n82_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n374_));
  NO2        m352(.A(i_11_), .B(i_12_), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n368_), .B(mai_mai_n224_), .Y(mai_mai_n376_));
  NA3        m354(.A(mai_mai_n110_), .B(i_4_), .C(i_11_), .Y(mai_mai_n377_));
  INV        m355(.A(mai_mai_n377_), .Y(mai_mai_n378_));
  NAi21      m356(.An(i_13_), .B(i_0_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(mai_mai_n227_), .Y(mai_mai_n380_));
  NA2        m358(.A(mai_mai_n378_), .B(mai_mai_n380_), .Y(mai_mai_n381_));
  NA3        m359(.A(mai_mai_n381_), .B(mai_mai_n373_), .C(mai_mai_n371_), .Y(mai_mai_n382_));
  NO3        m360(.A(i_1_), .B(i_12_), .C(mai_mai_n82_), .Y(mai_mai_n383_));
  NO2        m361(.A(i_0_), .B(i_11_), .Y(mai_mai_n384_));
  AN2        m362(.A(i_1_), .B(i_6_), .Y(mai_mai_n385_));
  NOi21      m363(.An(i_2_), .B(i_12_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n386_), .B(mai_mai_n385_), .Y(mai_mai_n387_));
  INV        m365(.A(mai_mai_n387_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n389_), .B(i_4_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n388_), .B(mai_mai_n390_), .Y(mai_mai_n391_));
  NAi21      m369(.An(i_9_), .B(i_4_), .Y(mai_mai_n392_));
  OR2        m370(.A(i_13_), .B(i_10_), .Y(mai_mai_n393_));
  NO3        m371(.A(mai_mai_n393_), .B(mai_mai_n113_), .C(mai_mai_n392_), .Y(mai_mai_n394_));
  BUFFER     m372(.A(mai_mai_n205_), .Y(mai_mai_n395_));
  NO2        m373(.A(mai_mai_n99_), .B(mai_mai_n25_), .Y(mai_mai_n396_));
  NA2        m374(.A(mai_mai_n266_), .B(mai_mai_n396_), .Y(mai_mai_n397_));
  NA2        m375(.A(mai_mai_n260_), .B(mai_mai_n202_), .Y(mai_mai_n398_));
  OAI220     m376(.A0(mai_mai_n398_), .A1(mai_mai_n395_), .B0(mai_mai_n397_), .B1(mai_mai_n324_), .Y(mai_mai_n399_));
  INV        m377(.A(mai_mai_n399_), .Y(mai_mai_n400_));
  AOI210     m378(.A0(mai_mai_n400_), .A1(mai_mai_n391_), .B0(mai_mai_n26_), .Y(mai_mai_n401_));
  NA2        m379(.A(mai_mai_n304_), .B(mai_mai_n303_), .Y(mai_mai_n402_));
  AOI220     m380(.A0(mai_mai_n278_), .A1(mai_mai_n269_), .B0(mai_mai_n272_), .B1(mai_mai_n295_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n403_), .B(i_5_), .Y(mai_mai_n404_));
  NO2        m382(.A(mai_mai_n177_), .B(mai_mai_n82_), .Y(mai_mai_n405_));
  AOI220     m383(.A0(mai_mai_n405_), .A1(mai_mai_n277_), .B0(i_6_), .B1(mai_mai_n202_), .Y(mai_mai_n406_));
  NO2        m384(.A(mai_mai_n406_), .B(mai_mai_n268_), .Y(mai_mai_n407_));
  NO3        m385(.A(mai_mai_n407_), .B(mai_mai_n404_), .C(mai_mai_n402_), .Y(mai_mai_n408_));
  NA2        m386(.A(mai_mai_n189_), .B(mai_mai_n94_), .Y(mai_mai_n409_));
  NA3        m387(.A(mai_mai_n305_), .B(mai_mai_n157_), .C(mai_mai_n82_), .Y(mai_mai_n410_));
  AOI210     m388(.A0(mai_mai_n410_), .A1(mai_mai_n409_), .B0(i_8_), .Y(mai_mai_n411_));
  INV        m389(.A(i_10_), .Y(mai_mai_n412_));
  NA3        m390(.A(mai_mai_n242_), .B(mai_mai_n62_), .C(i_2_), .Y(mai_mai_n413_));
  NA2        m391(.A(mai_mai_n278_), .B(mai_mai_n222_), .Y(mai_mai_n414_));
  OAI220     m392(.A0(mai_mai_n414_), .A1(mai_mai_n177_), .B0(mai_mai_n413_), .B1(mai_mai_n412_), .Y(mai_mai_n415_));
  NA3        m393(.A(mai_mai_n317_), .B(mai_mai_n316_), .C(i_5_), .Y(mai_mai_n416_));
  NA2        m394(.A(mai_mai_n297_), .B(mai_mai_n302_), .Y(mai_mai_n417_));
  OAI210     m395(.A0(mai_mai_n417_), .A1(mai_mai_n183_), .B0(mai_mai_n416_), .Y(mai_mai_n418_));
  NO3        m396(.A(mai_mai_n418_), .B(mai_mai_n415_), .C(mai_mai_n411_), .Y(mai_mai_n419_));
  AOI210     m397(.A0(mai_mai_n419_), .A1(mai_mai_n408_), .B0(mai_mai_n257_), .Y(mai_mai_n420_));
  NO4        m398(.A(mai_mai_n420_), .B(mai_mai_n401_), .C(mai_mai_n382_), .D(mai_mai_n361_), .Y(mai_mai_n421_));
  NO2        m399(.A(mai_mai_n71_), .B(i_13_), .Y(mai_mai_n422_));
  NO2        m400(.A(i_10_), .B(i_9_), .Y(mai_mai_n423_));
  NAi21      m401(.An(i_12_), .B(i_8_), .Y(mai_mai_n424_));
  NO2        m402(.A(mai_mai_n424_), .B(i_3_), .Y(mai_mai_n425_));
  NO3        m403(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n254_), .B(mai_mai_n95_), .Y(mai_mai_n427_));
  NA2        m405(.A(i_8_), .B(i_9_), .Y(mai_mai_n428_));
  NO3        m406(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n429_));
  NA3        m407(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n430_));
  OR2        m408(.A(mai_mai_n276_), .B(mai_mai_n199_), .Y(mai_mai_n431_));
  BUFFER     m409(.A(mai_mai_n279_), .Y(mai_mai_n432_));
  OA220      m410(.A0(mai_mai_n432_), .A1(mai_mai_n156_), .B0(mai_mai_n431_), .B1(mai_mai_n220_), .Y(mai_mai_n433_));
  NA2        m411(.A(mai_mai_n94_), .B(i_13_), .Y(mai_mai_n434_));
  INV        m412(.A(mai_mai_n362_), .Y(mai_mai_n435_));
  NO2        m413(.A(i_2_), .B(i_13_), .Y(mai_mai_n436_));
  NO2        m414(.A(mai_mai_n435_), .B(mai_mai_n434_), .Y(mai_mai_n437_));
  NO3        m415(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n438_));
  NO2        m416(.A(i_6_), .B(i_7_), .Y(mai_mai_n439_));
  NA2        m417(.A(mai_mai_n439_), .B(mai_mai_n438_), .Y(mai_mai_n440_));
  NO2        m418(.A(i_11_), .B(i_1_), .Y(mai_mai_n441_));
  NOi21      m419(.An(i_2_), .B(i_7_), .Y(mai_mai_n442_));
  NAi31      m420(.An(i_11_), .B(mai_mai_n442_), .C(mai_mai_n930_), .Y(mai_mai_n443_));
  NO2        m421(.A(mai_mai_n393_), .B(i_6_), .Y(mai_mai_n444_));
  NA3        m422(.A(mai_mai_n444_), .B(mai_mai_n935_), .C(mai_mai_n73_), .Y(mai_mai_n445_));
  NO2        m423(.A(mai_mai_n445_), .B(mai_mai_n443_), .Y(mai_mai_n446_));
  NO2        m424(.A(i_6_), .B(i_10_), .Y(mai_mai_n447_));
  NA3        m425(.A(mai_mai_n447_), .B(mai_mai_n294_), .C(i_8_), .Y(mai_mai_n448_));
  NO2        m426(.A(mai_mai_n448_), .B(mai_mai_n149_), .Y(mai_mai_n449_));
  NA3        m427(.A(mai_mai_n232_), .B(mai_mai_n165_), .C(mai_mai_n127_), .Y(mai_mai_n450_));
  NA2        m428(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n451_));
  NO2        m429(.A(mai_mai_n151_), .B(i_3_), .Y(mai_mai_n452_));
  NAi31      m430(.An(mai_mai_n451_), .B(mai_mai_n452_), .C(mai_mai_n215_), .Y(mai_mai_n453_));
  NA3        m431(.A(mai_mai_n372_), .B(mai_mai_n173_), .C(mai_mai_n143_), .Y(mai_mai_n454_));
  NA3        m432(.A(mai_mai_n454_), .B(mai_mai_n453_), .C(mai_mai_n450_), .Y(mai_mai_n455_));
  NO4        m433(.A(mai_mai_n455_), .B(mai_mai_n449_), .C(mai_mai_n446_), .D(mai_mai_n437_), .Y(mai_mai_n456_));
  NA2        m434(.A(mai_mai_n426_), .B(mai_mai_n363_), .Y(mai_mai_n457_));
  NO2        m435(.A(i_8_), .B(mai_mai_n213_), .Y(mai_mai_n458_));
  NAi21      m436(.An(mai_mai_n205_), .B(mai_mai_n375_), .Y(mai_mai_n459_));
  NO2        m437(.A(i_0_), .B(mai_mai_n82_), .Y(mai_mai_n460_));
  NA3        m438(.A(mai_mai_n460_), .B(mai_mai_n931_), .C(mai_mai_n136_), .Y(mai_mai_n461_));
  OR3        m439(.A(mai_mai_n284_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n462_));
  NO2        m440(.A(mai_mai_n462_), .B(mai_mai_n461_), .Y(mai_mai_n463_));
  NA2        m441(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n464_));
  NA2        m442(.A(mai_mai_n294_), .B(mai_mai_n226_), .Y(mai_mai_n465_));
  OAI220     m443(.A0(mai_mai_n465_), .A1(mai_mai_n413_), .B0(mai_mai_n464_), .B1(mai_mai_n434_), .Y(mai_mai_n466_));
  NA2        m444(.A(mai_mai_n287_), .B(mai_mai_n212_), .Y(mai_mai_n467_));
  NO2        m445(.A(mai_mai_n467_), .B(mai_mai_n440_), .Y(mai_mai_n468_));
  NO4        m446(.A(mai_mai_n468_), .B(mai_mai_n466_), .C(mai_mai_n463_), .D(mai_mai_n458_), .Y(mai_mai_n469_));
  NA3        m447(.A(mai_mai_n469_), .B(mai_mai_n456_), .C(mai_mai_n433_), .Y(mai_mai_n470_));
  NA3        m448(.A(mai_mai_n287_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n471_));
  OAI210     m449(.A0(mai_mai_n283_), .A1(mai_mai_n175_), .B0(mai_mai_n471_), .Y(mai_mai_n472_));
  BUFFER     m450(.A(mai_mai_n269_), .Y(mai_mai_n473_));
  NA2        m451(.A(mai_mai_n473_), .B(mai_mai_n472_), .Y(mai_mai_n474_));
  NA2        m452(.A(mai_mai_n118_), .B(mai_mai_n109_), .Y(mai_mai_n475_));
  AN2        m453(.A(mai_mai_n475_), .B(mai_mai_n426_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n294_), .B(mai_mai_n158_), .Y(mai_mai_n477_));
  OAI210     m455(.A0(mai_mai_n477_), .A1(mai_mai_n220_), .B0(mai_mai_n288_), .Y(mai_mai_n478_));
  AOI220     m456(.A0(mai_mai_n478_), .A1(i_7_), .B0(mai_mai_n476_), .B1(mai_mai_n290_), .Y(mai_mai_n479_));
  NA2        m457(.A(mai_mai_n363_), .B(mai_mai_n214_), .Y(mai_mai_n480_));
  NA2        m458(.A(mai_mai_n337_), .B(mai_mai_n71_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n350_), .B(mai_mai_n346_), .Y(mai_mai_n482_));
  OR2        m460(.A(mai_mai_n480_), .B(mai_mai_n482_), .Y(mai_mai_n483_));
  NO2        m461(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n484_));
  NAi41      m462(.An(mai_mai_n481_), .B(mai_mai_n447_), .C(mai_mai_n484_), .D(mai_mai_n46_), .Y(mai_mai_n485_));
  AOI210     m463(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n394_), .Y(mai_mai_n486_));
  NA3        m464(.A(mai_mai_n486_), .B(mai_mai_n485_), .C(mai_mai_n483_), .Y(mai_mai_n487_));
  INV        m465(.A(mai_mai_n487_), .Y(mai_mai_n488_));
  INV        m466(.A(mai_mai_n192_), .Y(mai_mai_n489_));
  OR2        m467(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n490_));
  NO2        m468(.A(mai_mai_n490_), .B(mai_mai_n82_), .Y(mai_mai_n491_));
  NA2        m469(.A(mai_mai_n491_), .B(mai_mai_n489_), .Y(mai_mai_n492_));
  NA4        m470(.A(mai_mai_n492_), .B(mai_mai_n488_), .C(mai_mai_n479_), .D(mai_mai_n474_), .Y(mai_mai_n493_));
  INV        m471(.A(mai_mai_n277_), .Y(mai_mai_n494_));
  OAI210     m472(.A0(mai_mai_n364_), .A1(mai_mai_n163_), .B0(mai_mai_n494_), .Y(mai_mai_n495_));
  NA2        m473(.A(mai_mai_n926_), .B(mai_mai_n214_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n447_), .B(mai_mai_n27_), .Y(mai_mai_n497_));
  NO2        m475(.A(mai_mai_n497_), .B(mai_mai_n496_), .Y(mai_mai_n498_));
  NOi31      m476(.An(mai_mai_n297_), .B(mai_mai_n393_), .C(mai_mai_n38_), .Y(mai_mai_n499_));
  OAI210     m477(.A0(mai_mai_n499_), .A1(mai_mai_n498_), .B0(mai_mai_n495_), .Y(mai_mai_n500_));
  NO2        m478(.A(i_8_), .B(i_7_), .Y(mai_mai_n501_));
  NO2        m479(.A(mai_mai_n46_), .B(mai_mai_n229_), .Y(mai_mai_n502_));
  NA2        m480(.A(mai_mai_n44_), .B(i_10_), .Y(mai_mai_n503_));
  NO2        m481(.A(mai_mai_n503_), .B(i_6_), .Y(mai_mai_n504_));
  NA3        m482(.A(mai_mai_n504_), .B(mai_mai_n502_), .C(mai_mai_n501_), .Y(mai_mai_n505_));
  OAI210     m483(.A0(mai_mai_n177_), .A1(mai_mai_n250_), .B0(mai_mai_n434_), .Y(mai_mai_n506_));
  NA2        m484(.A(mai_mai_n506_), .B(mai_mai_n253_), .Y(mai_mai_n507_));
  NOi31      m485(.An(mai_mai_n272_), .B(mai_mai_n283_), .C(mai_mai_n175_), .Y(mai_mai_n508_));
  NO2        m486(.A(mai_mai_n210_), .B(mai_mai_n44_), .Y(mai_mai_n509_));
  NO2        m487(.A(mai_mai_n151_), .B(i_5_), .Y(mai_mai_n510_));
  NA2        m488(.A(mai_mai_n510_), .B(mai_mai_n300_), .Y(mai_mai_n511_));
  NO2        m489(.A(mai_mai_n511_), .B(mai_mai_n509_), .Y(mai_mai_n512_));
  OAI210     m490(.A0(mai_mai_n512_), .A1(mai_mai_n508_), .B0(mai_mai_n429_), .Y(mai_mai_n513_));
  NA4        m491(.A(mai_mai_n513_), .B(mai_mai_n507_), .C(mai_mai_n505_), .D(mai_mai_n500_), .Y(mai_mai_n514_));
  NA2        m492(.A(mai_mai_n69_), .B(mai_mai_n44_), .Y(mai_mai_n515_));
  NA2        m493(.A(mai_mai_n266_), .B(mai_mai_n81_), .Y(mai_mai_n516_));
  AOI210     m494(.A0(mai_mai_n515_), .A1(mai_mai_n329_), .B0(mai_mai_n516_), .Y(mai_mai_n517_));
  NA2        m495(.A(mai_mai_n278_), .B(mai_mai_n269_), .Y(mai_mai_n518_));
  NO2        m496(.A(mai_mai_n518_), .B(mai_mai_n167_), .Y(mai_mai_n519_));
  NA2        m497(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n520_));
  NA2        m498(.A(mai_mai_n423_), .B(mai_mai_n210_), .Y(mai_mai_n521_));
  NO2        m499(.A(mai_mai_n520_), .B(mai_mai_n521_), .Y(mai_mai_n522_));
  NO3        m500(.A(mai_mai_n522_), .B(mai_mai_n519_), .C(mai_mai_n517_), .Y(mai_mai_n523_));
  NO4        m501(.A(mai_mai_n236_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n524_));
  NO3        m502(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n221_), .B(mai_mai_n36_), .Y(mai_mai_n526_));
  AN2        m504(.A(mai_mai_n526_), .B(mai_mai_n525_), .Y(mai_mai_n527_));
  OA210      m505(.A0(mai_mai_n527_), .A1(mai_mai_n524_), .B0(mai_mai_n337_), .Y(mai_mai_n528_));
  NO2        m506(.A(mai_mai_n393_), .B(i_1_), .Y(mai_mai_n529_));
  NOi31      m507(.An(mai_mai_n529_), .B(mai_mai_n427_), .C(mai_mai_n71_), .Y(mai_mai_n530_));
  AN3        m508(.A(mai_mai_n530_), .B(mai_mai_n390_), .C(i_2_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n403_), .B(mai_mai_n171_), .Y(mai_mai_n532_));
  NO3        m510(.A(mai_mai_n532_), .B(mai_mai_n531_), .C(mai_mai_n528_), .Y(mai_mai_n533_));
  NOi21      m511(.An(i_10_), .B(i_6_), .Y(mai_mai_n534_));
  NO2        m512(.A(mai_mai_n112_), .B(mai_mai_n23_), .Y(mai_mai_n535_));
  NA2        m513(.A(mai_mai_n297_), .B(mai_mai_n158_), .Y(mai_mai_n536_));
  AOI220     m514(.A0(mai_mai_n536_), .A1(mai_mai_n414_), .B0(mai_mai_n166_), .B1(mai_mai_n176_), .Y(mai_mai_n537_));
  NOi31      m515(.An(mai_mai_n140_), .B(i_1_), .C(mai_mai_n312_), .Y(mai_mai_n538_));
  NO2        m516(.A(mai_mai_n538_), .B(mai_mai_n537_), .Y(mai_mai_n539_));
  NO2        m517(.A(mai_mai_n481_), .B(mai_mai_n358_), .Y(mai_mai_n540_));
  NO2        m518(.A(i_12_), .B(mai_mai_n82_), .Y(mai_mai_n541_));
  NA2        m519(.A(mai_mai_n168_), .B(i_0_), .Y(mai_mai_n542_));
  NO3        m520(.A(mai_mai_n542_), .B(mai_mai_n322_), .C(mai_mai_n283_), .Y(mai_mai_n543_));
  NA2        m521(.A(mai_mai_n352_), .B(mai_mai_n231_), .Y(mai_mai_n544_));
  AOI210     m522(.A0(mai_mai_n544_), .A1(i_5_), .B0(mai_mai_n459_), .Y(mai_mai_n545_));
  NO3        m523(.A(mai_mai_n545_), .B(mai_mai_n543_), .C(mai_mai_n540_), .Y(mai_mai_n546_));
  NA4        m524(.A(mai_mai_n546_), .B(mai_mai_n539_), .C(mai_mai_n533_), .D(mai_mai_n523_), .Y(mai_mai_n547_));
  NO4        m525(.A(mai_mai_n547_), .B(mai_mai_n514_), .C(mai_mai_n493_), .D(mai_mai_n470_), .Y(mai_mai_n548_));
  NA4        m526(.A(mai_mai_n548_), .B(mai_mai_n421_), .C(mai_mai_n336_), .D(mai_mai_n293_), .Y(mai7));
  NO2        m527(.A(mai_mai_n91_), .B(mai_mai_n53_), .Y(mai_mai_n550_));
  NA2        m528(.A(mai_mai_n447_), .B(mai_mai_n81_), .Y(mai_mai_n551_));
  NA3        m529(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n552_));
  NO2        m530(.A(mai_mai_n224_), .B(i_4_), .Y(mai_mai_n553_));
  NA2        m531(.A(mai_mai_n553_), .B(i_8_), .Y(mai_mai_n554_));
  NO2        m532(.A(mai_mai_n103_), .B(mai_mai_n552_), .Y(mai_mai_n555_));
  NA2        m533(.A(i_2_), .B(mai_mai_n82_), .Y(mai_mai_n556_));
  OAI210     m534(.A0(mai_mai_n85_), .A1(mai_mai_n196_), .B0(mai_mai_n197_), .Y(mai_mai_n557_));
  NO2        m535(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n558_));
  NA2        m536(.A(i_4_), .B(i_8_), .Y(mai_mai_n559_));
  AOI210     m537(.A0(mai_mai_n559_), .A1(mai_mai_n287_), .B0(mai_mai_n558_), .Y(mai_mai_n560_));
  OAI220     m538(.A0(mai_mai_n560_), .A1(mai_mai_n556_), .B0(mai_mai_n557_), .B1(i_13_), .Y(mai_mai_n561_));
  NO3        m539(.A(mai_mai_n561_), .B(mai_mai_n555_), .C(mai_mai_n550_), .Y(mai_mai_n562_));
  OR2        m540(.A(i_6_), .B(i_10_), .Y(mai_mai_n563_));
  NO2        m541(.A(mai_mai_n563_), .B(mai_mai_n23_), .Y(mai_mai_n564_));
  OR3        m542(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n565_));
  NO3        m543(.A(mai_mai_n565_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n566_));
  INV        m544(.A(mai_mai_n193_), .Y(mai_mai_n567_));
  NO2        m545(.A(mai_mai_n566_), .B(mai_mai_n564_), .Y(mai_mai_n568_));
  OR2        m546(.A(mai_mai_n568_), .B(i_3_), .Y(mai_mai_n569_));
  AOI210     m547(.A0(mai_mai_n569_), .A1(mai_mai_n562_), .B0(mai_mai_n61_), .Y(mai_mai_n570_));
  NOi21      m548(.An(i_11_), .B(i_7_), .Y(mai_mai_n571_));
  AO210      m549(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n572_));
  NO2        m550(.A(mai_mai_n572_), .B(mai_mai_n571_), .Y(mai_mai_n573_));
  NA2        m551(.A(mai_mai_n573_), .B(mai_mai_n198_), .Y(mai_mai_n574_));
  NA3        m552(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n575_));
  NO2        m553(.A(mai_mai_n574_), .B(mai_mai_n61_), .Y(mai_mai_n576_));
  NA2        m554(.A(mai_mai_n84_), .B(mai_mai_n61_), .Y(mai_mai_n577_));
  AO210      m555(.A0(mai_mai_n577_), .A1(mai_mai_n358_), .B0(mai_mai_n41_), .Y(mai_mai_n578_));
  NA2        m556(.A(mai_mai_n215_), .B(mai_mai_n61_), .Y(mai_mai_n579_));
  OR2        m557(.A(mai_mai_n200_), .B(mai_mai_n106_), .Y(mai_mai_n580_));
  NO2        m558(.A(mai_mai_n61_), .B(i_9_), .Y(mai_mai_n581_));
  NO2        m559(.A(i_1_), .B(i_12_), .Y(mai_mai_n582_));
  NA2        m560(.A(mai_mai_n579_), .B(mai_mai_n578_), .Y(mai_mai_n583_));
  OAI210     m561(.A0(mai_mai_n583_), .A1(mai_mai_n576_), .B0(i_6_), .Y(mai_mai_n584_));
  NO2        m562(.A(mai_mai_n575_), .B(mai_mai_n106_), .Y(mai_mai_n585_));
  NA2        m563(.A(mai_mai_n585_), .B(mai_mai_n541_), .Y(mai_mai_n586_));
  NO2        m564(.A(i_6_), .B(i_11_), .Y(mai_mai_n587_));
  INV        m565(.A(mai_mai_n586_), .Y(mai_mai_n588_));
  NO4        m566(.A(i_12_), .B(mai_mai_n123_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n589_));
  NA2        m567(.A(mai_mai_n589_), .B(mai_mai_n581_), .Y(mai_mai_n590_));
  NA2        m568(.A(mai_mai_n224_), .B(i_6_), .Y(mai_mai_n591_));
  NO3        m569(.A(mai_mai_n563_), .B(mai_mai_n221_), .C(mai_mai_n23_), .Y(mai_mai_n592_));
  AOI210     m570(.A0(i_1_), .A1(mai_mai_n245_), .B0(mai_mai_n592_), .Y(mai_mai_n593_));
  OAI210     m571(.A0(mai_mai_n593_), .A1(mai_mai_n44_), .B0(mai_mai_n590_), .Y(mai_mai_n594_));
  NA3        m572(.A(mai_mai_n501_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n132_), .B(i_9_), .Y(mai_mai_n596_));
  NA3        m574(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n597_));
  NA3        m575(.A(i_2_), .B(mai_mai_n254_), .C(mai_mai_n44_), .Y(mai_mai_n598_));
  OAI220     m576(.A0(mai_mai_n598_), .A1(mai_mai_n597_), .B0(mai_mai_n596_), .B1(mai_mai_n925_), .Y(mai_mai_n599_));
  NA3        m577(.A(mai_mai_n581_), .B(mai_mai_n300_), .C(i_6_), .Y(mai_mai_n600_));
  NO2        m578(.A(mai_mai_n600_), .B(mai_mai_n23_), .Y(mai_mai_n601_));
  NA2        m579(.A(i_2_), .B(mai_mai_n254_), .Y(mai_mai_n602_));
  NO2        m580(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n603_));
  NA2        m581(.A(mai_mai_n603_), .B(mai_mai_n24_), .Y(mai_mai_n604_));
  NO2        m582(.A(mai_mai_n604_), .B(mai_mai_n602_), .Y(mai_mai_n605_));
  OR3        m583(.A(mai_mai_n605_), .B(mai_mai_n601_), .C(mai_mai_n599_), .Y(mai_mai_n606_));
  NO3        m584(.A(mai_mai_n606_), .B(mai_mai_n594_), .C(mai_mai_n588_), .Y(mai_mai_n607_));
  NO2        m585(.A(mai_mai_n224_), .B(mai_mai_n99_), .Y(mai_mai_n608_));
  NO2        m586(.A(mai_mai_n608_), .B(mai_mai_n571_), .Y(mai_mai_n609_));
  NA2        m587(.A(mai_mai_n609_), .B(i_1_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n610_), .B(mai_mai_n565_), .Y(mai_mai_n611_));
  NO2        m589(.A(mai_mai_n392_), .B(mai_mai_n82_), .Y(mai_mai_n612_));
  INV        m590(.A(mai_mai_n611_), .Y(mai_mai_n613_));
  NO2        m591(.A(mai_mai_n221_), .B(mai_mai_n44_), .Y(mai_mai_n614_));
  NO3        m592(.A(mai_mai_n614_), .B(mai_mai_n290_), .C(mai_mai_n225_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n113_), .B(mai_mai_n37_), .Y(mai_mai_n616_));
  NO2        m594(.A(mai_mai_n616_), .B(i_6_), .Y(mai_mai_n617_));
  NO2        m595(.A(mai_mai_n82_), .B(i_9_), .Y(mai_mai_n618_));
  NO2        m596(.A(mai_mai_n618_), .B(mai_mai_n61_), .Y(mai_mai_n619_));
  NO2        m597(.A(mai_mai_n619_), .B(mai_mai_n582_), .Y(mai_mai_n620_));
  NO4        m598(.A(mai_mai_n620_), .B(mai_mai_n617_), .C(mai_mai_n615_), .D(i_4_), .Y(mai_mai_n621_));
  NA2        m599(.A(i_1_), .B(i_3_), .Y(mai_mai_n622_));
  NO2        m600(.A(mai_mai_n428_), .B(mai_mai_n91_), .Y(mai_mai_n623_));
  AOI210     m601(.A0(mai_mai_n614_), .A1(mai_mai_n534_), .B0(mai_mai_n623_), .Y(mai_mai_n624_));
  NO2        m602(.A(mai_mai_n624_), .B(mai_mai_n622_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n625_), .B(mai_mai_n621_), .Y(mai_mai_n626_));
  NA4        m604(.A(mai_mai_n626_), .B(mai_mai_n613_), .C(mai_mai_n607_), .D(mai_mai_n584_), .Y(mai_mai_n627_));
  NO3        m605(.A(i_11_), .B(i_3_), .C(i_7_), .Y(mai_mai_n628_));
  NOi21      m606(.An(mai_mai_n628_), .B(i_10_), .Y(mai_mai_n629_));
  NA2        m607(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n630_));
  NA2        m608(.A(mai_mai_n447_), .B(mai_mai_n484_), .Y(mai_mai_n631_));
  NA2        m609(.A(mai_mai_n631_), .B(mai_mai_n630_), .Y(mai_mai_n632_));
  NA2        m610(.A(mai_mai_n632_), .B(i_1_), .Y(mai_mai_n633_));
  AOI210     m611(.A0(mai_mai_n254_), .A1(mai_mai_n95_), .B0(i_1_), .Y(mai_mai_n634_));
  NO2        m612(.A(mai_mai_n348_), .B(i_2_), .Y(mai_mai_n635_));
  NA2        m613(.A(mai_mai_n635_), .B(mai_mai_n634_), .Y(mai_mai_n636_));
  AOI210     m614(.A0(mai_mai_n636_), .A1(mai_mai_n633_), .B0(i_13_), .Y(mai_mai_n637_));
  OR2        m615(.A(i_11_), .B(i_7_), .Y(mai_mai_n638_));
  NO2        m616(.A(mai_mai_n53_), .B(i_12_), .Y(mai_mai_n639_));
  INV        m617(.A(mai_mai_n639_), .Y(mai_mai_n640_));
  AOI220     m618(.A0(i_7_), .A1(mai_mai_n612_), .B0(mai_mai_n232_), .B1(mai_mai_n126_), .Y(mai_mai_n641_));
  OAI220     m619(.A0(mai_mai_n641_), .A1(mai_mai_n41_), .B0(mai_mai_n640_), .B1(mai_mai_n91_), .Y(mai_mai_n642_));
  INV        m620(.A(mai_mai_n642_), .Y(mai_mai_n643_));
  AOI210     m621(.A0(mai_mai_n424_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n644_));
  NOi31      m622(.An(mai_mai_n644_), .B(mai_mai_n551_), .C(mai_mai_n44_), .Y(mai_mai_n645_));
  NA2        m623(.A(mai_mai_n122_), .B(i_13_), .Y(mai_mai_n646_));
  NO2        m624(.A(mai_mai_n597_), .B(mai_mai_n112_), .Y(mai_mai_n647_));
  INV        m625(.A(mai_mai_n647_), .Y(mai_mai_n648_));
  OAI220     m626(.A0(mai_mai_n648_), .A1(mai_mai_n69_), .B0(mai_mai_n646_), .B1(mai_mai_n634_), .Y(mai_mai_n649_));
  AOI220     m627(.A0(mai_mai_n365_), .A1(i_2_), .B0(mai_mai_n90_), .B1(mai_mai_n100_), .Y(mai_mai_n650_));
  NO2        m628(.A(mai_mai_n650_), .B(mai_mai_n554_), .Y(mai_mai_n651_));
  NO3        m629(.A(mai_mai_n651_), .B(mai_mai_n649_), .C(mai_mai_n645_), .Y(mai_mai_n652_));
  OR2        m630(.A(i_11_), .B(i_6_), .Y(mai_mai_n653_));
  NA2        m631(.A(mai_mai_n553_), .B(i_7_), .Y(mai_mai_n654_));
  AOI210     m632(.A0(mai_mai_n654_), .A1(mai_mai_n648_), .B0(mai_mai_n653_), .Y(mai_mai_n655_));
  NA3        m633(.A(mai_mai_n386_), .B(mai_mai_n558_), .C(mai_mai_n95_), .Y(mai_mai_n656_));
  NA2        m634(.A(mai_mai_n587_), .B(i_13_), .Y(mai_mai_n657_));
  NAi21      m635(.An(i_11_), .B(i_12_), .Y(mai_mai_n658_));
  NOi41      m636(.An(mai_mai_n108_), .B(mai_mai_n658_), .C(i_13_), .D(mai_mai_n82_), .Y(mai_mai_n659_));
  INV        m637(.A(mai_mai_n659_), .Y(mai_mai_n660_));
  NA3        m638(.A(mai_mai_n660_), .B(mai_mai_n657_), .C(mai_mai_n656_), .Y(mai_mai_n661_));
  OAI210     m639(.A0(mai_mai_n661_), .A1(mai_mai_n655_), .B0(mai_mai_n61_), .Y(mai_mai_n662_));
  NA2        m640(.A(mai_mai_n936_), .B(mai_mai_n347_), .Y(mai_mai_n663_));
  NO2        m641(.A(mai_mai_n123_), .B(i_2_), .Y(mai_mai_n664_));
  NA2        m642(.A(mai_mai_n664_), .B(mai_mai_n582_), .Y(mai_mai_n665_));
  NA2        m643(.A(mai_mai_n665_), .B(mai_mai_n663_), .Y(mai_mai_n666_));
  NA3        m644(.A(mai_mai_n666_), .B(mai_mai_n45_), .C(mai_mai_n214_), .Y(mai_mai_n667_));
  NA4        m645(.A(mai_mai_n667_), .B(mai_mai_n662_), .C(mai_mai_n652_), .D(mai_mai_n643_), .Y(mai_mai_n668_));
  OR4        m646(.A(mai_mai_n668_), .B(mai_mai_n637_), .C(mai_mai_n627_), .D(mai_mai_n570_), .Y(mai5));
  NA2        m647(.A(mai_mai_n609_), .B(mai_mai_n256_), .Y(mai_mai_n670_));
  NO2        m648(.A(mai_mai_n554_), .B(i_11_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n85_), .B(mai_mai_n671_), .Y(mai_mai_n672_));
  NA2        m650(.A(mai_mai_n672_), .B(mai_mai_n670_), .Y(mai_mai_n673_));
  NO3        m651(.A(i_11_), .B(mai_mai_n224_), .C(i_13_), .Y(mai_mai_n674_));
  NA2        m652(.A(i_12_), .B(i_8_), .Y(mai_mai_n675_));
  INV        m653(.A(mai_mai_n423_), .Y(mai_mai_n676_));
  NO2        m654(.A(mai_mai_n535_), .B(mai_mai_n673_), .Y(mai_mai_n677_));
  INV        m655(.A(mai_mai_n165_), .Y(mai_mai_n678_));
  INV        m656(.A(mai_mai_n232_), .Y(mai_mai_n679_));
  OAI210     m657(.A0(mai_mai_n635_), .A1(mai_mai_n425_), .B0(mai_mai_n108_), .Y(mai_mai_n680_));
  AOI210     m658(.A0(mai_mai_n680_), .A1(mai_mai_n679_), .B0(mai_mai_n678_), .Y(mai_mai_n681_));
  NO2        m659(.A(mai_mai_n428_), .B(mai_mai_n26_), .Y(mai_mai_n682_));
  NO2        m660(.A(mai_mai_n682_), .B(mai_mai_n396_), .Y(mai_mai_n683_));
  AOI210     m661(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n393_), .Y(mai_mai_n684_));
  AOI210     m662(.A0(mai_mai_n684_), .A1(i_2_), .B0(mai_mai_n681_), .Y(mai_mai_n685_));
  NO3        m663(.A(mai_mai_n572_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n686_));
  OA210      m664(.A0(mai_mai_n573_), .A1(mai_mai_n121_), .B0(i_13_), .Y(mai_mai_n687_));
  INV        m665(.A(mai_mai_n145_), .Y(mai_mai_n688_));
  NO2        m666(.A(mai_mai_n688_), .B(mai_mai_n352_), .Y(mai_mai_n689_));
  NA2        m667(.A(i_2_), .B(mai_mai_n396_), .Y(mai_mai_n690_));
  NA3        m668(.A(mai_mai_n287_), .B(mai_mai_n119_), .C(mai_mai_n42_), .Y(mai_mai_n691_));
  OAI210     m669(.A0(mai_mai_n691_), .A1(mai_mai_n46_), .B0(mai_mai_n690_), .Y(mai_mai_n692_));
  NO4        m670(.A(mai_mai_n692_), .B(mai_mai_n689_), .C(mai_mai_n687_), .D(mai_mai_n686_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n674_), .B(mai_mai_n259_), .Y(mai_mai_n694_));
  NO2        m672(.A(mai_mai_n60_), .B(i_12_), .Y(mai_mai_n695_));
  NA4        m673(.A(mai_mai_n694_), .B(mai_mai_n693_), .C(mai_mai_n685_), .D(mai_mai_n677_), .Y(mai6));
  NO3        m674(.A(mai_mai_n240_), .B(mai_mai_n289_), .C(i_1_), .Y(mai_mai_n697_));
  NO2        m675(.A(mai_mai_n179_), .B(mai_mai_n133_), .Y(mai_mai_n698_));
  OAI210     m676(.A0(mai_mai_n698_), .A1(mai_mai_n697_), .B0(mai_mai_n664_), .Y(mai_mai_n699_));
  INV        m677(.A(mai_mai_n310_), .Y(mai_mai_n700_));
  AO210      m678(.A0(mai_mai_n700_), .A1(mai_mai_n699_), .B0(i_12_), .Y(mai_mai_n701_));
  NA2        m679(.A(mai_mai_n353_), .B(mai_mai_n317_), .Y(mai_mai_n702_));
  NA2        m680(.A(mai_mai_n541_), .B(mai_mai_n61_), .Y(mai_mai_n703_));
  NA2        m681(.A(mai_mai_n629_), .B(mai_mai_n69_), .Y(mai_mai_n704_));
  BUFFER     m682(.A(mai_mai_n577_), .Y(mai_mai_n705_));
  NA4        m683(.A(mai_mai_n705_), .B(mai_mai_n704_), .C(mai_mai_n703_), .D(mai_mai_n702_), .Y(mai_mai_n706_));
  NA2        m684(.A(mai_mai_n706_), .B(mai_mai_n71_), .Y(mai_mai_n707_));
  INV        m685(.A(mai_mai_n309_), .Y(mai_mai_n708_));
  NA2        m686(.A(mai_mai_n73_), .B(mai_mai_n126_), .Y(mai_mai_n709_));
  AOI210     m687(.A0(mai_mai_n119_), .A1(mai_mai_n709_), .B0(mai_mai_n708_), .Y(mai_mai_n710_));
  NO2        m688(.A(mai_mai_n236_), .B(i_9_), .Y(mai_mai_n711_));
  NA2        m689(.A(mai_mai_n711_), .B(mai_mai_n695_), .Y(mai_mai_n712_));
  AOI210     m690(.A0(mai_mai_n712_), .A1(mai_mai_n482_), .B0(mai_mai_n179_), .Y(mai_mai_n713_));
  NO2        m691(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n714_));
  NA3        m692(.A(mai_mai_n714_), .B(mai_mai_n439_), .C(mai_mai_n368_), .Y(mai_mai_n715_));
  NAi32      m693(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n716_));
  NO2        m694(.A(mai_mai_n653_), .B(mai_mai_n716_), .Y(mai_mai_n717_));
  OAI210     m695(.A0(mai_mai_n628_), .A1(mai_mai_n526_), .B0(mai_mai_n525_), .Y(mai_mai_n718_));
  NAi31      m696(.An(mai_mai_n717_), .B(mai_mai_n718_), .C(mai_mai_n715_), .Y(mai_mai_n719_));
  OR3        m697(.A(mai_mai_n719_), .B(mai_mai_n713_), .C(mai_mai_n710_), .Y(mai_mai_n720_));
  NO2        m698(.A(mai_mai_n638_), .B(i_2_), .Y(mai_mai_n721_));
  NA2        m699(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n722_));
  NO2        m700(.A(mai_mai_n722_), .B(mai_mai_n385_), .Y(mai_mai_n723_));
  NA2        m701(.A(mai_mai_n723_), .B(mai_mai_n721_), .Y(mai_mai_n724_));
  AO210      m702(.A0(mai_mai_n341_), .A1(mai_mai_n333_), .B0(mai_mai_n374_), .Y(mai_mai_n725_));
  NA3        m703(.A(mai_mai_n725_), .B(mai_mai_n241_), .C(i_7_), .Y(mai_mai_n726_));
  OR2        m704(.A(mai_mai_n573_), .B(mai_mai_n425_), .Y(mai_mai_n727_));
  NA2        m705(.A(mai_mai_n727_), .B(mai_mai_n141_), .Y(mai_mai_n728_));
  OR2        m706(.A(mai_mai_n676_), .B(mai_mai_n36_), .Y(mai_mai_n729_));
  NA4        m707(.A(mai_mai_n729_), .B(mai_mai_n728_), .C(mai_mai_n726_), .D(mai_mai_n724_), .Y(mai_mai_n730_));
  NA2        m708(.A(mai_mai_n933_), .B(mai_mai_n525_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n374_), .B(mai_mai_n68_), .Y(mai_mai_n732_));
  NA3        m710(.A(mai_mai_n732_), .B(mai_mai_n731_), .C(mai_mai_n557_), .Y(mai_mai_n733_));
  OR2        m711(.A(mai_mai_n484_), .B(mai_mai_n84_), .Y(mai_mai_n734_));
  NA3        m712(.A(mai_mai_n734_), .B(mai_mai_n447_), .C(mai_mai_n207_), .Y(mai_mai_n735_));
  AOI210     m713(.A0(mai_mai_n425_), .A1(mai_mai_n423_), .B0(mai_mai_n524_), .Y(mai_mai_n736_));
  OAI210     m714(.A0(mai_mai_n939_), .A1(mai_mai_n109_), .B0(mai_mai_n384_), .Y(mai_mai_n737_));
  NA3        m715(.A(mai_mai_n737_), .B(mai_mai_n736_), .C(mai_mai_n735_), .Y(mai_mai_n738_));
  NO4        m716(.A(mai_mai_n738_), .B(mai_mai_n733_), .C(mai_mai_n730_), .D(mai_mai_n720_), .Y(mai_mai_n739_));
  NA4        m717(.A(mai_mai_n739_), .B(mai_mai_n707_), .C(mai_mai_n701_), .D(mai_mai_n360_), .Y(mai3));
  NA2        m718(.A(i_12_), .B(i_10_), .Y(mai_mai_n741_));
  INV        m719(.A(i_0_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n272_), .B(mai_mai_n940_), .Y(mai_mai_n743_));
  INV        m721(.A(mai_mai_n743_), .Y(mai_mai_n744_));
  NO3        m722(.A(mai_mai_n928_), .B(mai_mai_n88_), .C(mai_mai_n44_), .Y(mai_mai_n745_));
  OA210      m723(.A0(mai_mai_n745_), .A1(mai_mai_n744_), .B0(mai_mai_n168_), .Y(mai_mai_n746_));
  NOi21      m724(.An(mai_mai_n94_), .B(mai_mai_n683_), .Y(mai_mai_n747_));
  NO3        m725(.A(mai_mai_n580_), .B(mai_mai_n428_), .C(mai_mai_n126_), .Y(mai_mai_n748_));
  NO2        m726(.A(mai_mai_n748_), .B(mai_mai_n747_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n749_), .B(mai_mai_n48_), .Y(mai_mai_n750_));
  NO4        m728(.A(mai_mai_n356_), .B(mai_mai_n363_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n751_));
  INV        m729(.A(mai_mai_n751_), .Y(mai_mai_n752_));
  NA2        m730(.A(mai_mai_n644_), .B(mai_mai_n618_), .Y(mai_mai_n753_));
  NA2        m731(.A(mai_mai_n315_), .B(i_5_), .Y(mai_mai_n754_));
  OAI220     m732(.A0(mai_mai_n754_), .A1(mai_mai_n753_), .B0(mai_mai_n752_), .B1(mai_mai_n61_), .Y(mai_mai_n755_));
  NOi21      m733(.An(i_5_), .B(i_9_), .Y(mai_mai_n756_));
  NA2        m734(.A(mai_mai_n756_), .B(mai_mai_n422_), .Y(mai_mai_n757_));
  BUFFER     m735(.A(mai_mai_n254_), .Y(mai_mai_n758_));
  NA2        m736(.A(mai_mai_n758_), .B(mai_mai_n441_), .Y(mai_mai_n759_));
  NO2        m737(.A(mai_mai_n169_), .B(mai_mai_n142_), .Y(mai_mai_n760_));
  INV        m738(.A(mai_mai_n760_), .Y(mai_mai_n761_));
  OAI220     m739(.A0(mai_mai_n761_), .A1(mai_mai_n175_), .B0(mai_mai_n759_), .B1(mai_mai_n757_), .Y(mai_mai_n762_));
  NO4        m740(.A(mai_mai_n762_), .B(mai_mai_n755_), .C(mai_mai_n750_), .D(mai_mai_n746_), .Y(mai_mai_n763_));
  NA2        m741(.A(mai_mai_n179_), .B(mai_mai_n24_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n294_), .B(mai_mai_n124_), .Y(mai_mai_n765_));
  NAi21      m743(.An(mai_mai_n156_), .B(i_5_), .Y(mai_mai_n766_));
  NO2        m744(.A(mai_mai_n765_), .B(mai_mai_n376_), .Y(mai_mai_n767_));
  INV        m745(.A(mai_mai_n767_), .Y(mai_mai_n768_));
  NO2        m746(.A(mai_mai_n368_), .B(mai_mai_n276_), .Y(mai_mai_n769_));
  NA2        m747(.A(mai_mai_n769_), .B(mai_mai_n647_), .Y(mai_mai_n770_));
  AN2        m748(.A(mai_mai_n94_), .B(mai_mai_n230_), .Y(mai_mai_n771_));
  NA2        m749(.A(mai_mai_n674_), .B(mai_mai_n310_), .Y(mai_mai_n772_));
  AOI210     m750(.A0(mai_mai_n447_), .A1(mai_mai_n85_), .B0(mai_mai_n56_), .Y(mai_mai_n773_));
  NO2        m751(.A(mai_mai_n773_), .B(mai_mai_n772_), .Y(mai_mai_n774_));
  NO2        m752(.A(mai_mai_n238_), .B(mai_mai_n147_), .Y(mai_mai_n775_));
  NA2        m753(.A(i_0_), .B(i_10_), .Y(mai_mai_n776_));
  AN2        m754(.A(mai_mai_n775_), .B(i_6_), .Y(mai_mai_n777_));
  NA2        m755(.A(mai_mai_n315_), .B(mai_mai_n96_), .Y(mai_mai_n778_));
  NA2        m756(.A(mai_mai_n529_), .B(i_4_), .Y(mai_mai_n779_));
  NA2        m757(.A(mai_mai_n182_), .B(mai_mai_n196_), .Y(mai_mai_n780_));
  OAI220     m758(.A0(mai_mai_n780_), .A1(mai_mai_n772_), .B0(mai_mai_n779_), .B1(mai_mai_n778_), .Y(mai_mai_n781_));
  NO4        m759(.A(mai_mai_n781_), .B(mai_mai_n777_), .C(mai_mai_n774_), .D(mai_mai_n771_), .Y(mai_mai_n782_));
  NA3        m760(.A(mai_mai_n782_), .B(mai_mai_n770_), .C(mai_mai_n768_), .Y(mai_mai_n783_));
  NA2        m761(.A(i_11_), .B(i_9_), .Y(mai_mai_n784_));
  NO2        m762(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n785_));
  NA2        m763(.A(mai_mai_n372_), .B(mai_mai_n173_), .Y(mai_mai_n786_));
  NA2        m764(.A(mai_mai_n786_), .B(mai_mai_n154_), .Y(mai_mai_n787_));
  NO2        m765(.A(mai_mai_n784_), .B(mai_mai_n71_), .Y(mai_mai_n788_));
  NO2        m766(.A(mai_mai_n169_), .B(i_0_), .Y(mai_mai_n789_));
  NA2        m767(.A(mai_mai_n439_), .B(mai_mai_n219_), .Y(mai_mai_n790_));
  INV        m768(.A(mai_mai_n383_), .Y(mai_mai_n791_));
  OAI220     m769(.A0(mai_mai_n791_), .A1(mai_mai_n757_), .B0(mai_mai_n790_), .B1(mai_mai_n169_), .Y(mai_mai_n792_));
  NO2        m770(.A(mai_mai_n792_), .B(mai_mai_n787_), .Y(mai_mai_n793_));
  NA2        m771(.A(mai_mai_n603_), .B(mai_mai_n117_), .Y(mai_mai_n794_));
  NO2        m772(.A(i_6_), .B(mai_mai_n794_), .Y(mai_mai_n795_));
  AOI210     m773(.A0(mai_mai_n424_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n796_));
  NA2        m774(.A(mai_mai_n165_), .B(mai_mai_n101_), .Y(mai_mai_n797_));
  NOi32      m775(.An(mai_mai_n796_), .Bn(mai_mai_n182_), .C(mai_mai_n797_), .Y(mai_mai_n798_));
  NO2        m776(.A(mai_mai_n798_), .B(mai_mai_n795_), .Y(mai_mai_n799_));
  NOi21      m777(.An(i_7_), .B(i_5_), .Y(mai_mai_n800_));
  NOi31      m778(.An(mai_mai_n800_), .B(i_0_), .C(mai_mai_n658_), .Y(mai_mai_n801_));
  NA3        m779(.A(mai_mai_n801_), .B(mai_mai_n937_), .C(i_6_), .Y(mai_mai_n802_));
  OA210      m780(.A0(mai_mai_n797_), .A1(mai_mai_n482_), .B0(mai_mai_n802_), .Y(mai_mai_n803_));
  NO3        m781(.A(mai_mai_n379_), .B(mai_mai_n344_), .C(mai_mai_n340_), .Y(mai_mai_n804_));
  NO2        m782(.A(mai_mai_n248_), .B(mai_mai_n301_), .Y(mai_mai_n805_));
  NO2        m783(.A(mai_mai_n658_), .B(mai_mai_n243_), .Y(mai_mai_n806_));
  AOI210     m784(.A0(mai_mai_n806_), .A1(mai_mai_n805_), .B0(mai_mai_n804_), .Y(mai_mai_n807_));
  NA4        m785(.A(mai_mai_n807_), .B(mai_mai_n803_), .C(mai_mai_n799_), .D(mai_mai_n793_), .Y(mai_mai_n808_));
  NO2        m786(.A(mai_mai_n764_), .B(mai_mai_n227_), .Y(mai_mai_n809_));
  AN2        m787(.A(mai_mai_n314_), .B(mai_mai_n310_), .Y(mai_mai_n810_));
  AN2        m788(.A(mai_mai_n810_), .B(mai_mai_n760_), .Y(mai_mai_n811_));
  OAI210     m789(.A0(mai_mai_n811_), .A1(mai_mai_n809_), .B0(i_10_), .Y(mai_mai_n812_));
  NO2        m790(.A(mai_mai_n741_), .B(mai_mai_n300_), .Y(mai_mai_n813_));
  OA210      m791(.A0(mai_mai_n439_), .A1(mai_mai_n212_), .B0(mai_mai_n438_), .Y(mai_mai_n814_));
  NA2        m792(.A(mai_mai_n813_), .B(mai_mai_n788_), .Y(mai_mai_n815_));
  NA3        m793(.A(mai_mai_n438_), .B(mai_mai_n386_), .C(mai_mai_n45_), .Y(mai_mai_n816_));
  OAI210     m794(.A0(mai_mai_n766_), .A1(i_6_), .B0(mai_mai_n816_), .Y(mai_mai_n817_));
  NO2        m795(.A(mai_mai_n241_), .B(mai_mai_n46_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n818_), .B(mai_mai_n181_), .Y(mai_mai_n819_));
  AOI220     m797(.A0(mai_mai_n819_), .A1(mai_mai_n439_), .B0(mai_mai_n817_), .B1(mai_mai_n71_), .Y(mai_mai_n820_));
  NA3        m798(.A(mai_mai_n722_), .B(mai_mai_n362_), .C(i_6_), .Y(mai_mai_n821_));
  NA2        m799(.A(mai_mai_n91_), .B(mai_mai_n44_), .Y(mai_mai_n822_));
  NO2        m800(.A(mai_mai_n73_), .B(mai_mai_n675_), .Y(mai_mai_n823_));
  NA2        m801(.A(mai_mai_n823_), .B(mai_mai_n822_), .Y(mai_mai_n824_));
  AOI210     m802(.A0(mai_mai_n824_), .A1(mai_mai_n821_), .B0(mai_mai_n47_), .Y(mai_mai_n825_));
  NO2        m803(.A(mai_mai_n552_), .B(mai_mai_n103_), .Y(mai_mai_n826_));
  NA2        m804(.A(mai_mai_n826_), .B(i_0_), .Y(mai_mai_n827_));
  NO2        m805(.A(mai_mai_n827_), .B(mai_mai_n82_), .Y(mai_mai_n828_));
  NO3        m806(.A(mai_mai_n828_), .B(mai_mai_n825_), .C(mai_mai_n487_), .Y(mai_mai_n829_));
  NA4        m807(.A(mai_mai_n829_), .B(mai_mai_n820_), .C(mai_mai_n815_), .D(mai_mai_n812_), .Y(mai_mai_n830_));
  NO3        m808(.A(mai_mai_n830_), .B(mai_mai_n808_), .C(mai_mai_n783_), .Y(mai_mai_n831_));
  AOI210     m809(.A0(mai_mai_n703_), .A1(mai_mai_n630_), .B0(mai_mai_n797_), .Y(mai_mai_n832_));
  AOI210     m810(.A0(mai_mai_n168_), .A1(mai_mai_n330_), .B0(mai_mai_n832_), .Y(mai_mai_n833_));
  NO2        m811(.A(mai_mai_n718_), .B(mai_mai_n379_), .Y(mai_mai_n834_));
  NA3        m812(.A(mai_mai_n742_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n835_));
  NA2        m813(.A(mai_mai_n940_), .B(i_9_), .Y(mai_mai_n836_));
  AOI210     m814(.A0(mai_mai_n835_), .A1(mai_mai_n461_), .B0(mai_mai_n836_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n837_), .B(mai_mai_n834_), .Y(mai_mai_n838_));
  NA2        m816(.A(mai_mai_n838_), .B(mai_mai_n833_), .Y(mai_mai_n839_));
  NA2        m817(.A(mai_mai_n810_), .B(mai_mai_n352_), .Y(mai_mai_n840_));
  AOI210     m818(.A0(mai_mai_n283_), .A1(mai_mai_n156_), .B0(mai_mai_n840_), .Y(mai_mai_n841_));
  NA2        m819(.A(mai_mai_n785_), .B(mai_mai_n452_), .Y(mai_mai_n842_));
  AOI210     m820(.A0(i_11_), .A1(mai_mai_n156_), .B0(mai_mai_n842_), .Y(mai_mai_n843_));
  NO2        m821(.A(mai_mai_n843_), .B(mai_mai_n841_), .Y(mai_mai_n844_));
  NO3        m822(.A(mai_mai_n776_), .B(mai_mai_n756_), .C(mai_mai_n184_), .Y(mai_mai_n845_));
  AOI220     m823(.A0(mai_mai_n845_), .A1(i_11_), .B0(mai_mai_n530_), .B1(mai_mai_n73_), .Y(mai_mai_n846_));
  NO3        m824(.A(mai_mai_n201_), .B(mai_mai_n363_), .C(i_0_), .Y(mai_mai_n847_));
  OAI210     m825(.A0(mai_mai_n847_), .A1(mai_mai_n74_), .B0(i_13_), .Y(mai_mai_n848_));
  OAI220     m826(.A0(mai_mai_n496_), .A1(mai_mai_n133_), .B0(mai_mai_n591_), .B1(mai_mai_n567_), .Y(mai_mai_n849_));
  NA3        m827(.A(mai_mai_n849_), .B(i_7_), .C(i_0_), .Y(mai_mai_n850_));
  NA4        m828(.A(mai_mai_n850_), .B(mai_mai_n848_), .C(mai_mai_n846_), .D(mai_mai_n844_), .Y(mai_mai_n851_));
  NA2        m829(.A(mai_mai_n333_), .B(mai_mai_n170_), .Y(mai_mai_n852_));
  OR2        m830(.A(mai_mai_n852_), .B(mai_mai_n929_), .Y(mai_mai_n853_));
  AOI210     m831(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n169_), .Y(mai_mai_n854_));
  NA2        m832(.A(mai_mai_n854_), .B(mai_mai_n814_), .Y(mai_mai_n855_));
  NA3        m833(.A(mai_mai_n564_), .B(mai_mai_n179_), .C(mai_mai_n81_), .Y(mai_mai_n856_));
  INV        m834(.A(mai_mai_n856_), .Y(mai_mai_n857_));
  NO3        m835(.A(mai_mai_n938_), .B(mai_mai_n53_), .C(mai_mai_n48_), .Y(mai_mai_n858_));
  NA2        m836(.A(mai_mai_n457_), .B(mai_mai_n450_), .Y(mai_mai_n859_));
  NO3        m837(.A(mai_mai_n859_), .B(mai_mai_n858_), .C(mai_mai_n857_), .Y(mai_mai_n860_));
  NA3        m838(.A(mai_mai_n368_), .B(mai_mai_n165_), .C(mai_mai_n164_), .Y(mai_mai_n861_));
  INV        m839(.A(mai_mai_n861_), .Y(mai_mai_n862_));
  NA3        m840(.A(mai_mai_n368_), .B(mai_mai_n316_), .C(mai_mai_n210_), .Y(mai_mai_n863_));
  INV        m841(.A(mai_mai_n863_), .Y(mai_mai_n864_));
  NO3        m842(.A(mai_mai_n784_), .B(mai_mai_n207_), .C(mai_mai_n184_), .Y(mai_mai_n865_));
  NO3        m843(.A(mai_mai_n865_), .B(mai_mai_n864_), .C(mai_mai_n862_), .Y(mai_mai_n866_));
  NA4        m844(.A(mai_mai_n866_), .B(mai_mai_n860_), .C(mai_mai_n855_), .D(mai_mai_n853_), .Y(mai_mai_n867_));
  INV        m845(.A(mai_mai_n566_), .Y(mai_mai_n868_));
  NO3        m846(.A(mai_mai_n868_), .B(i_5_), .C(mai_mai_n327_), .Y(mai_mai_n869_));
  INV        m847(.A(mai_mai_n869_), .Y(mai_mai_n870_));
  NA2        m848(.A(mai_mai_n287_), .B(i_5_), .Y(mai_mai_n871_));
  NO4        m849(.A(mai_mai_n227_), .B(mai_mai_n201_), .C(i_0_), .D(i_12_), .Y(mai_mai_n872_));
  NA2        m850(.A(mai_mai_n872_), .B(i_10_), .Y(mai_mai_n873_));
  AN2        m851(.A(mai_mai_n776_), .B(mai_mai_n147_), .Y(mai_mai_n874_));
  NO4        m852(.A(mai_mai_n874_), .B(i_12_), .C(mai_mai_n595_), .D(mai_mai_n126_), .Y(mai_mai_n875_));
  INV        m853(.A(mai_mai_n875_), .Y(mai_mai_n876_));
  NA3        m854(.A(mai_mai_n96_), .B(mai_mai_n534_), .C(i_11_), .Y(mai_mai_n877_));
  NA2        m855(.A(mai_mai_n800_), .B(mai_mai_n436_), .Y(mai_mai_n878_));
  OAI220     m856(.A0(i_7_), .A1(mai_mai_n871_), .B0(mai_mai_n878_), .B1(mai_mai_n619_), .Y(mai_mai_n879_));
  NA2        m857(.A(mai_mai_n879_), .B(mai_mai_n789_), .Y(mai_mai_n880_));
  NA4        m858(.A(mai_mai_n880_), .B(mai_mai_n876_), .C(mai_mai_n873_), .D(mai_mai_n870_), .Y(mai_mai_n881_));
  NO4        m859(.A(mai_mai_n881_), .B(mai_mai_n867_), .C(mai_mai_n851_), .D(mai_mai_n839_), .Y(mai_mai_n882_));
  OAI210     m860(.A0(mai_mai_n721_), .A1(mai_mai_n714_), .B0(mai_mai_n37_), .Y(mai_mai_n883_));
  NA3        m861(.A(mai_mai_n796_), .B(mai_mai_n347_), .C(i_5_), .Y(mai_mai_n884_));
  NA2        m862(.A(mai_mai_n884_), .B(mai_mai_n883_), .Y(mai_mai_n885_));
  NA2        m863(.A(mai_mai_n885_), .B(mai_mai_n198_), .Y(mai_mai_n886_));
  BUFFER     m864(.A(mai_mai_n348_), .Y(mai_mai_n887_));
  NA2        m865(.A(mai_mai_n180_), .B(mai_mai_n182_), .Y(mai_mai_n888_));
  AO210      m866(.A0(mai_mai_n887_), .A1(mai_mai_n33_), .B0(mai_mai_n888_), .Y(mai_mai_n889_));
  OAI210     m867(.A0(mai_mai_n566_), .A1(mai_mai_n564_), .B0(mai_mai_n300_), .Y(mai_mai_n890_));
  NAi31      m868(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n891_));
  NO2        m869(.A(mai_mai_n68_), .B(mai_mai_n891_), .Y(mai_mai_n892_));
  NO2        m870(.A(mai_mai_n892_), .B(mai_mai_n592_), .Y(mai_mai_n893_));
  NA3        m871(.A(mai_mai_n893_), .B(mai_mai_n890_), .C(mai_mai_n889_), .Y(mai_mai_n894_));
  NO2        m872(.A(mai_mai_n430_), .B(mai_mai_n254_), .Y(mai_mai_n895_));
  NO4        m873(.A(mai_mai_n221_), .B(mai_mai_n139_), .C(mai_mai_n622_), .D(mai_mai_n37_), .Y(mai_mai_n896_));
  NO2        m874(.A(mai_mai_n896_), .B(mai_mai_n895_), .Y(mai_mai_n897_));
  OAI210     m875(.A0(mai_mai_n877_), .A1(mai_mai_n142_), .B0(mai_mai_n897_), .Y(mai_mai_n898_));
  AOI210     m876(.A0(mai_mai_n894_), .A1(mai_mai_n48_), .B0(mai_mai_n898_), .Y(mai_mai_n899_));
  AOI210     m877(.A0(mai_mai_n899_), .A1(mai_mai_n886_), .B0(mai_mai_n71_), .Y(mai_mai_n900_));
  NO2        m878(.A(mai_mai_n527_), .B(mai_mai_n359_), .Y(mai_mai_n901_));
  NO2        m879(.A(mai_mai_n901_), .B(mai_mai_n678_), .Y(mai_mai_n902_));
  NA2        m880(.A(mai_mai_n53_), .B(mai_mai_n106_), .Y(mai_mai_n903_));
  NA2        m881(.A(mai_mai_n903_), .B(mai_mai_n74_), .Y(mai_mai_n904_));
  AOI210     m882(.A0(mai_mai_n854_), .A1(mai_mai_n785_), .B0(mai_mai_n801_), .Y(mai_mai_n905_));
  AOI210     m883(.A0(mai_mai_n905_), .A1(mai_mai_n904_), .B0(mai_mai_n622_), .Y(mai_mai_n906_));
  NA2        m884(.A(mai_mai_n248_), .B(mai_mai_n55_), .Y(mai_mai_n907_));
  AOI220     m885(.A0(mai_mai_n907_), .A1(mai_mai_n74_), .B0(mai_mai_n328_), .B1(mai_mai_n240_), .Y(mai_mai_n908_));
  NO2        m886(.A(mai_mai_n908_), .B(mai_mai_n224_), .Y(mai_mai_n909_));
  NA3        m887(.A(mai_mai_n94_), .B(mai_mai_n289_), .C(mai_mai_n31_), .Y(mai_mai_n910_));
  INV        m888(.A(mai_mai_n910_), .Y(mai_mai_n911_));
  NO3        m889(.A(mai_mai_n911_), .B(mai_mai_n909_), .C(mai_mai_n906_), .Y(mai_mai_n912_));
  OAI210     m890(.A0(mai_mai_n255_), .A1(mai_mai_n152_), .B0(mai_mai_n85_), .Y(mai_mai_n913_));
  NA3        m891(.A(mai_mai_n682_), .B(mai_mai_n272_), .C(mai_mai_n78_), .Y(mai_mai_n914_));
  AOI210     m892(.A0(mai_mai_n914_), .A1(mai_mai_n913_), .B0(i_11_), .Y(mai_mai_n915_));
  OAI210     m893(.A0(mai_mai_n927_), .A1(mai_mai_n796_), .B0(mai_mai_n198_), .Y(mai_mai_n916_));
  NA2        m894(.A(mai_mai_n158_), .B(i_5_), .Y(mai_mai_n917_));
  NO2        m895(.A(mai_mai_n916_), .B(mai_mai_n917_), .Y(mai_mai_n918_));
  NO2        m896(.A(mai_mai_n918_), .B(mai_mai_n915_), .Y(mai_mai_n919_));
  OAI210     m897(.A0(mai_mai_n912_), .A1(i_4_), .B0(mai_mai_n919_), .Y(mai_mai_n920_));
  NO3        m898(.A(mai_mai_n920_), .B(mai_mai_n902_), .C(mai_mai_n900_), .Y(mai_mai_n921_));
  NA4        m899(.A(mai_mai_n921_), .B(mai_mai_n882_), .C(mai_mai_n831_), .D(mai_mai_n763_), .Y(mai4));
  INV        m900(.A(i_2_), .Y(mai_mai_n925_));
  INV        m901(.A(i_12_), .Y(mai_mai_n926_));
  INV        m902(.A(i_12_), .Y(mai_mai_n927_));
  INV        m903(.A(i_0_), .Y(mai_mai_n928_));
  INV        m904(.A(mai_mai_n157_), .Y(mai_mai_n929_));
  INV        m905(.A(i_3_), .Y(mai_mai_n930_));
  INV        m906(.A(i_5_), .Y(mai_mai_n931_));
  INV        m907(.A(mai_mai_n233_), .Y(mai_mai_n932_));
  INV        m908(.A(i_11_), .Y(mai_mai_n933_));
  INV        m909(.A(i_12_), .Y(mai_mai_n934_));
  INV        m910(.A(i_4_), .Y(mai_mai_n935_));
  INV        m911(.A(i_9_), .Y(mai_mai_n936_));
  INV        m912(.A(i_4_), .Y(mai_mai_n937_));
  INV        m913(.A(mai_mai_n386_), .Y(mai_mai_n938_));
  INV        m914(.A(mai_mai_n563_), .Y(mai_mai_n939_));
  INV        m915(.A(i_11_), .Y(mai_mai_n940_));
  NAi21      u000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u002(.A(i_9_), .Y(men_men_n25_));
  INV        u003(.A(i_3_), .Y(men_men_n26_));
  NO2        u004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u013(.A(i_4_), .Y(men_men_n36_));
  INV        u014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u021(.A(men_men_n35_), .Y(men1));
  INV        u022(.A(i_11_), .Y(men_men_n45_));
  NO2        u023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u024(.A(i_2_), .Y(men_men_n47_));
  NA2        u025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u026(.A(i_5_), .Y(men_men_n49_));
  NO2        u027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NO2        u033(.A(men_men_n55_), .B(men_men_n54_), .Y(men_men_n56_));
  NA2        u034(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n57_));
  NO2        u035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  NAi21      u037(.An(i_2_), .B(i_7_), .Y(men_men_n60_));
  INV        u038(.A(i_1_), .Y(men_men_n61_));
  NA2        u039(.A(men_men_n61_), .B(i_6_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n51_), .B(i_2_), .Y(men_men_n63_));
  AOI210     u041(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n64_));
  NA2        u042(.A(i_1_), .B(i_6_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n65_), .B(men_men_n25_), .Y(men_men_n66_));
  INV        u044(.A(i_0_), .Y(men_men_n67_));
  NAi21      u045(.An(i_5_), .B(i_10_), .Y(men_men_n68_));
  NA2        u046(.A(i_5_), .B(i_9_), .Y(men_men_n69_));
  AOI210     u047(.A0(men_men_n69_), .A1(men_men_n68_), .B0(men_men_n67_), .Y(men_men_n70_));
  NO2        u048(.A(men_men_n70_), .B(men_men_n66_), .Y(men_men_n71_));
  OAI210     u049(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n71_), .Y(men_men_n72_));
  NA2        u050(.A(men_men_n72_), .B(i_0_), .Y(men_men_n73_));
  NA2        u051(.A(i_12_), .B(i_5_), .Y(men_men_n74_));
  NA2        u052(.A(i_2_), .B(i_8_), .Y(men_men_n75_));
  NO2        u053(.A(i_3_), .B(i_9_), .Y(men_men_n76_));
  NO2        u054(.A(i_3_), .B(i_7_), .Y(men_men_n77_));
  NO3        u055(.A(men_men_n77_), .B(men_men_n76_), .C(men_men_n61_), .Y(men_men_n78_));
  INV        u056(.A(i_6_), .Y(men_men_n79_));
  OR4        u057(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n80_));
  INV        u058(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u059(.A(i_2_), .B(i_7_), .Y(men_men_n82_));
  OAI210     u060(.A0(men_men_n78_), .A1(i_8_), .B0(i_2_), .Y(men_men_n83_));
  NAi21      u061(.An(i_6_), .B(i_10_), .Y(men_men_n84_));
  NA2        u062(.A(i_6_), .B(i_9_), .Y(men_men_n85_));
  AOI210     u063(.A0(men_men_n85_), .A1(men_men_n84_), .B0(men_men_n61_), .Y(men_men_n86_));
  NA2        u064(.A(i_2_), .B(i_6_), .Y(men_men_n87_));
  NO3        u065(.A(men_men_n87_), .B(men_men_n50_), .C(men_men_n25_), .Y(men_men_n88_));
  NO2        u066(.A(men_men_n88_), .B(men_men_n86_), .Y(men_men_n89_));
  AOI210     u067(.A0(men_men_n89_), .A1(men_men_n83_), .B0(men_men_n74_), .Y(men_men_n90_));
  AN3        u068(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n91_));
  NAi21      u069(.An(i_6_), .B(i_11_), .Y(men_men_n92_));
  NO2        u070(.A(i_5_), .B(i_8_), .Y(men_men_n93_));
  NOi21      u071(.An(men_men_n93_), .B(men_men_n92_), .Y(men_men_n94_));
  AOI220     u072(.A0(men_men_n94_), .A1(men_men_n60_), .B0(men_men_n91_), .B1(men_men_n32_), .Y(men_men_n95_));
  INV        u073(.A(i_7_), .Y(men_men_n96_));
  NA2        u074(.A(men_men_n47_), .B(men_men_n96_), .Y(men_men_n97_));
  NO2        u075(.A(i_0_), .B(i_5_), .Y(men_men_n98_));
  NO2        u076(.A(men_men_n98_), .B(men_men_n79_), .Y(men_men_n99_));
  NA2        u077(.A(i_12_), .B(i_3_), .Y(men_men_n100_));
  INV        u078(.A(men_men_n100_), .Y(men_men_n101_));
  NA3        u079(.A(men_men_n101_), .B(men_men_n99_), .C(men_men_n97_), .Y(men_men_n102_));
  NAi21      u080(.An(i_7_), .B(i_11_), .Y(men_men_n103_));
  NO3        u081(.A(men_men_n103_), .B(men_men_n84_), .C(men_men_n54_), .Y(men_men_n104_));
  AN2        u082(.A(i_2_), .B(i_10_), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n105_), .B(i_7_), .Y(men_men_n106_));
  OR2        u084(.A(men_men_n74_), .B(men_men_n58_), .Y(men_men_n107_));
  NO2        u085(.A(i_8_), .B(men_men_n96_), .Y(men_men_n108_));
  NO3        u086(.A(men_men_n108_), .B(men_men_n107_), .C(men_men_n106_), .Y(men_men_n109_));
  NA2        u087(.A(i_12_), .B(i_7_), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n61_), .B(men_men_n26_), .Y(men_men_n111_));
  NA2        u089(.A(men_men_n111_), .B(i_0_), .Y(men_men_n112_));
  NA2        u090(.A(i_11_), .B(i_12_), .Y(men_men_n113_));
  OAI210     u091(.A0(men_men_n112_), .A1(men_men_n110_), .B0(men_men_n113_), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n114_), .B(men_men_n109_), .Y(men_men_n115_));
  NAi41      u093(.An(men_men_n104_), .B(men_men_n115_), .C(men_men_n102_), .D(men_men_n95_), .Y(men_men_n116_));
  NOi21      u094(.An(i_1_), .B(i_5_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n117_), .B(i_11_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n96_), .B(men_men_n37_), .Y(men_men_n119_));
  NA2        u097(.A(i_7_), .B(men_men_n25_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n120_), .B(men_men_n119_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(men_men_n47_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n85_), .B(men_men_n84_), .Y(men_men_n123_));
  NAi21      u101(.An(i_3_), .B(i_8_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n124_), .B(men_men_n60_), .Y(men_men_n125_));
  NOi31      u103(.An(men_men_n125_), .B(men_men_n123_), .C(men_men_n122_), .Y(men_men_n126_));
  NO2        u104(.A(i_1_), .B(men_men_n79_), .Y(men_men_n127_));
  NO2        u105(.A(i_6_), .B(i_5_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n128_), .B(i_3_), .Y(men_men_n129_));
  AO210      u107(.A0(men_men_n129_), .A1(men_men_n48_), .B0(men_men_n127_), .Y(men_men_n130_));
  OAI220     u108(.A0(men_men_n130_), .A1(men_men_n103_), .B0(men_men_n126_), .B1(men_men_n118_), .Y(men_men_n131_));
  NO3        u109(.A(men_men_n131_), .B(men_men_n116_), .C(men_men_n90_), .Y(men_men_n132_));
  NA3        u110(.A(men_men_n132_), .B(men_men_n73_), .C(men_men_n57_), .Y(men2));
  NO2        u111(.A(men_men_n61_), .B(men_men_n37_), .Y(men_men_n134_));
  NA2        u112(.A(i_6_), .B(men_men_n25_), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(men_men_n134_), .Y(men_men_n136_));
  NA4        u114(.A(men_men_n136_), .B(men_men_n71_), .C(men_men_n63_), .D(men_men_n30_), .Y(men0));
  AN2        u115(.A(i_8_), .B(i_7_), .Y(men_men_n138_));
  NA2        u116(.A(men_men_n138_), .B(i_6_), .Y(men_men_n139_));
  NO2        u117(.A(i_12_), .B(i_13_), .Y(men_men_n140_));
  NAi21      u118(.An(i_5_), .B(i_11_), .Y(men_men_n141_));
  NOi21      u119(.An(men_men_n140_), .B(men_men_n141_), .Y(men_men_n142_));
  NO2        u120(.A(i_0_), .B(i_1_), .Y(men_men_n143_));
  NA2        u121(.A(i_2_), .B(i_3_), .Y(men_men_n144_));
  NO2        u122(.A(men_men_n144_), .B(i_4_), .Y(men_men_n145_));
  NA3        u123(.A(men_men_n145_), .B(men_men_n143_), .C(men_men_n142_), .Y(men_men_n146_));
  OR2        u124(.A(men_men_n146_), .B(men_men_n25_), .Y(men_men_n147_));
  AN2        u125(.A(men_men_n140_), .B(men_men_n76_), .Y(men_men_n148_));
  NO2        u126(.A(men_men_n148_), .B(men_men_n27_), .Y(men_men_n149_));
  NA2        u127(.A(i_1_), .B(i_5_), .Y(men_men_n150_));
  NO2        u128(.A(men_men_n67_), .B(men_men_n47_), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n151_), .B(men_men_n36_), .Y(men_men_n152_));
  NO3        u130(.A(men_men_n152_), .B(men_men_n150_), .C(men_men_n149_), .Y(men_men_n153_));
  OR2        u131(.A(i_0_), .B(i_1_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n154_), .B(men_men_n74_), .C(i_13_), .Y(men_men_n155_));
  NAi32      u133(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n156_));
  NAi21      u134(.An(men_men_n156_), .B(men_men_n155_), .Y(men_men_n157_));
  NOi21      u135(.An(i_4_), .B(i_10_), .Y(men_men_n158_));
  NA2        u136(.A(men_men_n158_), .B(men_men_n40_), .Y(men_men_n159_));
  NO2        u137(.A(i_3_), .B(i_5_), .Y(men_men_n160_));
  NO3        u138(.A(men_men_n67_), .B(i_2_), .C(i_1_), .Y(men_men_n161_));
  OAI210     u139(.A0(i_3_), .A1(men_men_n159_), .B0(men_men_n157_), .Y(men_men_n162_));
  NO2        u140(.A(men_men_n162_), .B(men_men_n153_), .Y(men_men_n163_));
  AOI210     u141(.A0(men_men_n163_), .A1(men_men_n147_), .B0(men_men_n139_), .Y(men_men_n164_));
  NA2        u142(.A(i_3_), .B(men_men_n49_), .Y(men_men_n165_));
  NOi21      u143(.An(i_4_), .B(i_9_), .Y(men_men_n166_));
  NOi21      u144(.An(i_11_), .B(i_13_), .Y(men_men_n167_));
  NA2        u145(.A(men_men_n167_), .B(men_men_n166_), .Y(men_men_n168_));
  OR2        u146(.A(men_men_n168_), .B(men_men_n165_), .Y(men_men_n169_));
  NO2        u147(.A(i_4_), .B(i_5_), .Y(men_men_n170_));
  NAi21      u148(.An(i_12_), .B(i_11_), .Y(men_men_n171_));
  NO2        u149(.A(men_men_n171_), .B(i_13_), .Y(men_men_n172_));
  NA3        u150(.A(men_men_n172_), .B(men_men_n170_), .C(men_men_n76_), .Y(men_men_n173_));
  AOI210     u151(.A0(men_men_n173_), .A1(men_men_n169_), .B0(i_0_), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n67_), .B(men_men_n61_), .Y(men_men_n175_));
  NA2        u153(.A(men_men_n175_), .B(men_men_n47_), .Y(men_men_n176_));
  NA2        u154(.A(men_men_n36_), .B(i_5_), .Y(men_men_n177_));
  NAi31      u155(.An(men_men_n177_), .B(men_men_n148_), .C(i_11_), .Y(men_men_n178_));
  NA2        u156(.A(i_3_), .B(i_5_), .Y(men_men_n179_));
  OR2        u157(.A(men_men_n179_), .B(men_men_n168_), .Y(men_men_n180_));
  AOI210     u158(.A0(men_men_n180_), .A1(men_men_n178_), .B0(men_men_n176_), .Y(men_men_n181_));
  NO2        u159(.A(men_men_n67_), .B(i_5_), .Y(men_men_n182_));
  NO2        u160(.A(i_13_), .B(i_10_), .Y(men_men_n183_));
  NA3        u161(.A(men_men_n183_), .B(men_men_n182_), .C(men_men_n45_), .Y(men_men_n184_));
  NO2        u162(.A(i_2_), .B(i_1_), .Y(men_men_n185_));
  NA2        u163(.A(men_men_n185_), .B(i_3_), .Y(men_men_n186_));
  NAi21      u164(.An(i_4_), .B(i_12_), .Y(men_men_n187_));
  NO3        u165(.A(men_men_n187_), .B(men_men_n186_), .C(men_men_n25_), .Y(men_men_n188_));
  NO3        u166(.A(men_men_n188_), .B(men_men_n181_), .C(men_men_n174_), .Y(men_men_n189_));
  INV        u167(.A(i_8_), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n190_), .B(i_7_), .Y(men_men_n191_));
  NA2        u169(.A(men_men_n191_), .B(i_6_), .Y(men_men_n192_));
  NO3        u170(.A(i_3_), .B(men_men_n79_), .C(men_men_n49_), .Y(men_men_n193_));
  NA2        u171(.A(men_men_n193_), .B(men_men_n108_), .Y(men_men_n194_));
  NO3        u172(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n195_));
  NA3        u173(.A(men_men_n195_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n196_));
  NO3        u174(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n197_));
  OAI210     u175(.A0(men_men_n91_), .A1(i_12_), .B0(men_men_n197_), .Y(men_men_n198_));
  AOI210     u176(.A0(men_men_n198_), .A1(men_men_n196_), .B0(men_men_n194_), .Y(men_men_n199_));
  NO2        u177(.A(i_3_), .B(i_8_), .Y(men_men_n200_));
  NO3        u178(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n201_));
  NA3        u179(.A(men_men_n201_), .B(men_men_n200_), .C(men_men_n40_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n98_), .B(men_men_n58_), .Y(men_men_n203_));
  INV        u181(.A(men_men_n203_), .Y(men_men_n204_));
  NO2        u182(.A(i_13_), .B(i_9_), .Y(men_men_n205_));
  NA3        u183(.A(men_men_n205_), .B(i_6_), .C(men_men_n190_), .Y(men_men_n206_));
  NAi21      u184(.An(i_12_), .B(i_3_), .Y(men_men_n207_));
  OR2        u185(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n45_), .B(i_5_), .Y(men_men_n209_));
  NO3        u187(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n210_));
  NA2        u188(.A(men_men_n210_), .B(i_10_), .Y(men_men_n211_));
  OAI220     u189(.A0(men_men_n211_), .A1(men_men_n208_), .B0(men_men_n204_), .B1(men_men_n202_), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n212_), .A1(i_7_), .B0(men_men_n199_), .Y(men_men_n213_));
  OAI220     u191(.A0(men_men_n213_), .A1(i_4_), .B0(men_men_n192_), .B1(men_men_n189_), .Y(men_men_n214_));
  NAi21      u192(.An(i_12_), .B(i_7_), .Y(men_men_n215_));
  NA3        u193(.A(i_13_), .B(men_men_n190_), .C(i_10_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n217_));
  NA2        u195(.A(i_0_), .B(i_5_), .Y(men_men_n218_));
  OAI220     u196(.A0(men_men_n79_), .A1(men_men_n186_), .B0(men_men_n176_), .B1(men_men_n129_), .Y(men_men_n219_));
  NAi31      u197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n220_));
  NO2        u198(.A(men_men_n47_), .B(men_men_n61_), .Y(men_men_n221_));
  NA3        u199(.A(men_men_n221_), .B(i_0_), .C(i_4_), .Y(men_men_n222_));
  INV        u200(.A(i_13_), .Y(men_men_n223_));
  NO2        u201(.A(i_12_), .B(men_men_n223_), .Y(men_men_n224_));
  NA3        u202(.A(men_men_n224_), .B(men_men_n195_), .C(men_men_n193_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n222_), .A1(men_men_n220_), .B0(men_men_n225_), .Y(men_men_n226_));
  AOI220     u204(.A0(men_men_n226_), .A1(men_men_n138_), .B0(men_men_n219_), .B1(men_men_n217_), .Y(men_men_n227_));
  NO2        u205(.A(i_12_), .B(men_men_n37_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n179_), .B(i_4_), .Y(men_men_n229_));
  NA2        u207(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  OR2        u208(.A(i_8_), .B(i_7_), .Y(men_men_n231_));
  NO2        u209(.A(men_men_n231_), .B(men_men_n79_), .Y(men_men_n232_));
  NO2        u210(.A(men_men_n54_), .B(i_1_), .Y(men_men_n233_));
  NA2        u211(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  INV        u212(.A(i_12_), .Y(men_men_n235_));
  NO3        u213(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n236_));
  NA2        u214(.A(i_2_), .B(i_1_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n234_), .B(men_men_n230_), .Y(men_men_n238_));
  NO3        u216(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n239_));
  NAi21      u217(.An(i_4_), .B(i_3_), .Y(men_men_n240_));
  NO2        u218(.A(i_0_), .B(i_6_), .Y(men_men_n241_));
  NOi41      u219(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n242_));
  NA2        u220(.A(men_men_n242_), .B(men_men_n241_), .Y(men_men_n243_));
  NO2        u221(.A(men_men_n237_), .B(men_men_n179_), .Y(men_men_n244_));
  NAi21      u222(.An(men_men_n243_), .B(men_men_n244_), .Y(men_men_n245_));
  INV        u223(.A(men_men_n245_), .Y(men_men_n246_));
  AOI220     u224(.A0(men_men_n246_), .A1(men_men_n40_), .B0(men_men_n238_), .B1(men_men_n205_), .Y(men_men_n247_));
  NO2        u225(.A(i_11_), .B(men_men_n223_), .Y(men_men_n248_));
  NOi21      u226(.An(i_1_), .B(i_6_), .Y(men_men_n249_));
  NAi21      u227(.An(i_3_), .B(i_7_), .Y(men_men_n250_));
  NO2        u228(.A(i_12_), .B(i_3_), .Y(men_men_n251_));
  NA3        u229(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n252_));
  INV        u230(.A(men_men_n139_), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n235_), .B(i_13_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n254_), .B(men_men_n69_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n255_), .B(men_men_n253_), .Y(men_men_n256_));
  NO2        u234(.A(men_men_n231_), .B(men_men_n37_), .Y(men_men_n257_));
  NA2        u235(.A(i_12_), .B(i_6_), .Y(men_men_n258_));
  OR2        u236(.A(i_13_), .B(i_9_), .Y(men_men_n259_));
  NO3        u237(.A(men_men_n259_), .B(men_men_n258_), .C(men_men_n49_), .Y(men_men_n260_));
  NO2        u238(.A(men_men_n240_), .B(i_2_), .Y(men_men_n261_));
  NA3        u239(.A(men_men_n261_), .B(men_men_n260_), .C(men_men_n45_), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n248_), .B(i_9_), .Y(men_men_n263_));
  NA2        u241(.A(i_0_), .B(men_men_n62_), .Y(men_men_n264_));
  OAI210     u242(.A0(men_men_n264_), .A1(men_men_n263_), .B0(men_men_n262_), .Y(men_men_n265_));
  NA2        u243(.A(men_men_n151_), .B(men_men_n61_), .Y(men_men_n266_));
  NO3        u244(.A(i_11_), .B(men_men_n223_), .C(men_men_n25_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n250_), .B(i_8_), .Y(men_men_n268_));
  NA3        u246(.A(i_5_), .B(men_men_n268_), .C(men_men_n267_), .Y(men_men_n269_));
  NO3        u247(.A(men_men_n26_), .B(men_men_n79_), .C(i_5_), .Y(men_men_n270_));
  NA3        u248(.A(men_men_n270_), .B(men_men_n257_), .C(men_men_n224_), .Y(men_men_n271_));
  AOI210     u249(.A0(men_men_n271_), .A1(men_men_n269_), .B0(men_men_n266_), .Y(men_men_n272_));
  AOI210     u250(.A0(men_men_n265_), .A1(men_men_n257_), .B0(men_men_n272_), .Y(men_men_n273_));
  NA4        u251(.A(men_men_n273_), .B(men_men_n256_), .C(men_men_n247_), .D(men_men_n227_), .Y(men_men_n274_));
  NO3        u252(.A(i_12_), .B(men_men_n223_), .C(men_men_n37_), .Y(men_men_n275_));
  INV        u253(.A(men_men_n275_), .Y(men_men_n276_));
  NO3        u254(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n277_));
  AOI220     u255(.A0(men_men_n277_), .A1(men_men_n193_), .B0(men_men_n160_), .B1(men_men_n233_), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n278_), .B(men_men_n969_), .Y(men_men_n279_));
  NO3        u257(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n280_));
  NO2        u258(.A(men_men_n237_), .B(i_0_), .Y(men_men_n281_));
  AOI220     u259(.A0(men_men_n281_), .A1(men_men_n191_), .B0(men_men_n280_), .B1(men_men_n138_), .Y(men_men_n282_));
  NO2        u260(.A(i_3_), .B(men_men_n282_), .Y(men_men_n283_));
  NA2        u261(.A(i_0_), .B(i_1_), .Y(men_men_n284_));
  NO2        u262(.A(men_men_n284_), .B(i_2_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n59_), .B(i_6_), .Y(men_men_n286_));
  NA3        u264(.A(men_men_n286_), .B(men_men_n285_), .C(men_men_n160_), .Y(men_men_n287_));
  OAI210     u265(.A0(i_3_), .A1(men_men_n139_), .B0(men_men_n287_), .Y(men_men_n288_));
  NO3        u266(.A(men_men_n288_), .B(men_men_n283_), .C(men_men_n279_), .Y(men_men_n289_));
  NO2        u267(.A(i_3_), .B(i_10_), .Y(men_men_n290_));
  NA3        u268(.A(men_men_n290_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n291_));
  NO2        u269(.A(i_2_), .B(men_men_n96_), .Y(men_men_n292_));
  NOi21      u270(.An(men_men_n218_), .B(men_men_n98_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n294_));
  AN2        u272(.A(i_3_), .B(i_10_), .Y(men_men_n295_));
  NA4        u273(.A(men_men_n295_), .B(men_men_n195_), .C(men_men_n172_), .D(men_men_n170_), .Y(men_men_n296_));
  NO2        u274(.A(i_5_), .B(men_men_n37_), .Y(men_men_n297_));
  NO2        u275(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n298_));
  OR2        u276(.A(men_men_n294_), .B(men_men_n291_), .Y(men_men_n299_));
  OAI220     u277(.A0(men_men_n299_), .A1(i_6_), .B0(men_men_n289_), .B1(men_men_n276_), .Y(men_men_n300_));
  NO4        u278(.A(men_men_n300_), .B(men_men_n274_), .C(men_men_n214_), .D(men_men_n164_), .Y(men_men_n301_));
  NO3        u279(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n302_));
  NA2        u280(.A(men_men_n281_), .B(i_8_), .Y(men_men_n303_));
  NO3        u281(.A(i_6_), .B(men_men_n190_), .C(i_7_), .Y(men_men_n304_));
  AOI210     u282(.A0(men_men_n971_), .A1(men_men_n303_), .B0(men_men_n165_), .Y(men_men_n305_));
  NO2        u283(.A(i_2_), .B(i_3_), .Y(men_men_n306_));
  OR2        u284(.A(i_0_), .B(i_5_), .Y(men_men_n307_));
  NA3        u285(.A(men_men_n232_), .B(men_men_n306_), .C(i_1_), .Y(men_men_n308_));
  NA3        u286(.A(men_men_n281_), .B(men_men_n160_), .C(men_men_n108_), .Y(men_men_n309_));
  NAi21      u287(.An(i_8_), .B(i_7_), .Y(men_men_n310_));
  NO2        u288(.A(men_men_n310_), .B(i_6_), .Y(men_men_n311_));
  NO2        u289(.A(men_men_n154_), .B(men_men_n47_), .Y(men_men_n312_));
  NA3        u290(.A(men_men_n312_), .B(men_men_n311_), .C(men_men_n160_), .Y(men_men_n313_));
  NA3        u291(.A(men_men_n313_), .B(men_men_n309_), .C(men_men_n308_), .Y(men_men_n314_));
  OAI210     u292(.A0(men_men_n314_), .A1(men_men_n305_), .B0(i_4_), .Y(men_men_n315_));
  NO2        u293(.A(i_12_), .B(i_10_), .Y(men_men_n316_));
  NOi21      u294(.An(i_5_), .B(i_0_), .Y(men_men_n317_));
  AOI210     u295(.A0(i_2_), .A1(men_men_n49_), .B0(men_men_n96_), .Y(men_men_n318_));
  NO3        u296(.A(men_men_n318_), .B(i_4_), .C(men_men_n124_), .Y(men_men_n319_));
  NA4        u297(.A(men_men_n77_), .B(men_men_n36_), .C(men_men_n79_), .D(i_8_), .Y(men_men_n320_));
  NA2        u298(.A(men_men_n319_), .B(men_men_n316_), .Y(men_men_n321_));
  NO2        u299(.A(i_6_), .B(i_8_), .Y(men_men_n322_));
  NO2        u300(.A(i_1_), .B(i_7_), .Y(men_men_n323_));
  AO220      u301(.A0(men_men_n323_), .A1(men_men_n322_), .B0(men_men_n311_), .B1(men_men_n233_), .Y(men_men_n324_));
  NA2        u302(.A(men_men_n324_), .B(men_men_n42_), .Y(men_men_n325_));
  NA3        u303(.A(men_men_n325_), .B(men_men_n321_), .C(men_men_n315_), .Y(men_men_n326_));
  NO3        u304(.A(men_men_n231_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n327_));
  NO3        u305(.A(men_men_n310_), .B(i_2_), .C(i_1_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n328_), .A1(men_men_n327_), .B0(i_6_), .Y(men_men_n329_));
  NA3        u307(.A(men_men_n249_), .B(men_men_n292_), .C(men_men_n190_), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(men_men_n329_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n331_), .B(i_3_), .Y(men_men_n332_));
  NO2        u310(.A(men_men_n284_), .B(men_men_n75_), .Y(men_men_n333_));
  NA2        u311(.A(men_men_n333_), .B(men_men_n128_), .Y(men_men_n334_));
  NO2        u312(.A(men_men_n87_), .B(men_men_n190_), .Y(men_men_n335_));
  NA3        u313(.A(men_men_n293_), .B(men_men_n335_), .C(men_men_n61_), .Y(men_men_n336_));
  AOI210     u314(.A0(men_men_n336_), .A1(men_men_n334_), .B0(i_7_), .Y(men_men_n337_));
  NO2        u315(.A(men_men_n190_), .B(i_9_), .Y(men_men_n338_));
  NA2        u316(.A(men_men_n338_), .B(men_men_n203_), .Y(men_men_n339_));
  NO2        u317(.A(men_men_n337_), .B(men_men_n283_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n340_), .A1(men_men_n332_), .B0(men_men_n159_), .Y(men_men_n341_));
  AOI210     u319(.A0(men_men_n326_), .A1(men_men_n302_), .B0(men_men_n341_), .Y(men_men_n342_));
  NOi32      u320(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n343_));
  INV        u321(.A(men_men_n343_), .Y(men_men_n344_));
  NAi21      u322(.An(i_0_), .B(i_6_), .Y(men_men_n345_));
  NAi21      u323(.An(i_1_), .B(i_5_), .Y(men_men_n346_));
  NAi41      u324(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n347_));
  OAI220     u325(.A0(men_men_n347_), .A1(men_men_n346_), .B0(men_men_n220_), .B1(men_men_n156_), .Y(men_men_n348_));
  AOI210     u326(.A0(men_men_n347_), .A1(men_men_n156_), .B0(men_men_n154_), .Y(men_men_n349_));
  NOi32      u327(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n350_));
  NA2        u328(.A(men_men_n350_), .B(men_men_n47_), .Y(men_men_n351_));
  NO2        u329(.A(men_men_n351_), .B(i_0_), .Y(men_men_n352_));
  OR3        u330(.A(men_men_n352_), .B(men_men_n349_), .C(men_men_n348_), .Y(men_men_n353_));
  NO2        u331(.A(i_1_), .B(men_men_n96_), .Y(men_men_n354_));
  NAi21      u332(.An(i_3_), .B(i_4_), .Y(men_men_n355_));
  NO2        u333(.A(men_men_n355_), .B(i_9_), .Y(men_men_n356_));
  AN2        u334(.A(i_6_), .B(i_7_), .Y(men_men_n357_));
  OAI210     u335(.A0(men_men_n357_), .A1(men_men_n354_), .B0(men_men_n356_), .Y(men_men_n358_));
  NA2        u336(.A(i_2_), .B(i_7_), .Y(men_men_n359_));
  NO2        u337(.A(men_men_n355_), .B(i_10_), .Y(men_men_n360_));
  NA3        u338(.A(men_men_n360_), .B(men_men_n359_), .C(men_men_n241_), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n361_), .A1(men_men_n358_), .B0(men_men_n182_), .Y(men_men_n362_));
  AOI210     u340(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n363_));
  OAI210     u341(.A0(men_men_n363_), .A1(men_men_n185_), .B0(men_men_n360_), .Y(men_men_n364_));
  AOI220     u342(.A0(men_men_n360_), .A1(men_men_n323_), .B0(men_men_n236_), .B1(men_men_n185_), .Y(men_men_n365_));
  AOI210     u343(.A0(men_men_n365_), .A1(men_men_n364_), .B0(i_5_), .Y(men_men_n366_));
  NO3        u344(.A(men_men_n366_), .B(men_men_n362_), .C(men_men_n353_), .Y(men_men_n367_));
  NO2        u345(.A(men_men_n367_), .B(men_men_n344_), .Y(men_men_n368_));
  NO2        u346(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n369_));
  AN2        u347(.A(i_12_), .B(i_5_), .Y(men_men_n370_));
  NO2        u348(.A(i_4_), .B(men_men_n26_), .Y(men_men_n371_));
  NA2        u349(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  NO2        u350(.A(i_11_), .B(i_6_), .Y(men_men_n373_));
  NA3        u351(.A(men_men_n373_), .B(men_men_n312_), .C(men_men_n223_), .Y(men_men_n374_));
  NO2        u352(.A(men_men_n374_), .B(men_men_n372_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n240_), .B(i_5_), .Y(men_men_n376_));
  NO2        u354(.A(i_5_), .B(i_10_), .Y(men_men_n377_));
  AOI220     u355(.A0(men_men_n377_), .A1(men_men_n261_), .B0(men_men_n376_), .B1(men_men_n195_), .Y(men_men_n378_));
  NA2        u356(.A(men_men_n140_), .B(men_men_n46_), .Y(men_men_n379_));
  NO2        u357(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n380_));
  OAI210     u358(.A0(men_men_n380_), .A1(men_men_n375_), .B0(men_men_n369_), .Y(men_men_n381_));
  NO2        u359(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n382_));
  NO2        u360(.A(men_men_n146_), .B(men_men_n79_), .Y(men_men_n383_));
  OAI210     u361(.A0(men_men_n383_), .A1(men_men_n375_), .B0(men_men_n382_), .Y(men_men_n384_));
  NO3        u362(.A(men_men_n79_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n385_));
  NO2        u363(.A(i_11_), .B(i_12_), .Y(men_men_n386_));
  NA2        u364(.A(men_men_n377_), .B(men_men_n235_), .Y(men_men_n387_));
  NA2        u365(.A(men_men_n42_), .B(i_11_), .Y(men_men_n388_));
  OAI220     u366(.A0(men_men_n388_), .A1(men_men_n220_), .B0(men_men_n387_), .B1(men_men_n320_), .Y(men_men_n389_));
  NAi21      u367(.An(i_13_), .B(i_0_), .Y(men_men_n390_));
  NO2        u368(.A(men_men_n390_), .B(men_men_n237_), .Y(men_men_n391_));
  NA2        u369(.A(men_men_n389_), .B(men_men_n391_), .Y(men_men_n392_));
  NA3        u370(.A(men_men_n392_), .B(men_men_n384_), .C(men_men_n381_), .Y(men_men_n393_));
  NA2        u371(.A(men_men_n45_), .B(men_men_n223_), .Y(men_men_n394_));
  NO3        u372(.A(i_1_), .B(i_12_), .C(men_men_n79_), .Y(men_men_n395_));
  NO2        u373(.A(i_0_), .B(i_11_), .Y(men_men_n396_));
  INV        u374(.A(i_5_), .Y(men_men_n397_));
  AN2        u375(.A(i_1_), .B(i_6_), .Y(men_men_n398_));
  NOi21      u376(.An(i_2_), .B(i_12_), .Y(men_men_n399_));
  NA2        u377(.A(men_men_n399_), .B(men_men_n398_), .Y(men_men_n400_));
  NO2        u378(.A(men_men_n400_), .B(men_men_n397_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n138_), .B(i_9_), .Y(men_men_n402_));
  NO2        u380(.A(men_men_n402_), .B(i_4_), .Y(men_men_n403_));
  NA2        u381(.A(men_men_n401_), .B(men_men_n403_), .Y(men_men_n404_));
  OR2        u382(.A(i_13_), .B(i_10_), .Y(men_men_n405_));
  NO2        u383(.A(men_men_n168_), .B(men_men_n119_), .Y(men_men_n406_));
  OR2        u384(.A(men_men_n216_), .B(men_men_n215_), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n96_), .B(men_men_n25_), .Y(men_men_n408_));
  NA2        u386(.A(i_5_), .B(men_men_n210_), .Y(men_men_n409_));
  NO2        u387(.A(men_men_n409_), .B(men_men_n407_), .Y(men_men_n410_));
  INV        u388(.A(men_men_n410_), .Y(men_men_n411_));
  AOI210     u389(.A0(men_men_n411_), .A1(men_men_n404_), .B0(men_men_n26_), .Y(men_men_n412_));
  NA2        u390(.A(men_men_n309_), .B(men_men_n308_), .Y(men_men_n413_));
  AOI220     u391(.A0(men_men_n286_), .A1(men_men_n277_), .B0(men_men_n281_), .B1(i_8_), .Y(men_men_n414_));
  NO2        u392(.A(men_men_n414_), .B(men_men_n165_), .Y(men_men_n415_));
  NO2        u393(.A(men_men_n179_), .B(men_men_n79_), .Y(men_men_n416_));
  AOI220     u394(.A0(men_men_n416_), .A1(men_men_n285_), .B0(men_men_n270_), .B1(men_men_n210_), .Y(men_men_n417_));
  INV        u395(.A(men_men_n417_), .Y(men_men_n418_));
  NO3        u396(.A(men_men_n418_), .B(men_men_n415_), .C(men_men_n413_), .Y(men_men_n419_));
  INV        u397(.A(men_men_n91_), .Y(men_men_n420_));
  AOI210     u398(.A0(men_men_n154_), .A1(men_men_n420_), .B0(men_men_n310_), .Y(men_men_n421_));
  NA2        u399(.A(men_men_n286_), .B(men_men_n233_), .Y(men_men_n422_));
  NO2        u400(.A(men_men_n422_), .B(men_men_n179_), .Y(men_men_n423_));
  NO2        u401(.A(i_3_), .B(men_men_n49_), .Y(men_men_n424_));
  NA3        u402(.A(men_men_n323_), .B(men_men_n322_), .C(men_men_n424_), .Y(men_men_n425_));
  OAI210     u403(.A0(men_men_n190_), .A1(men_men_n186_), .B0(men_men_n425_), .Y(men_men_n426_));
  NO3        u404(.A(men_men_n426_), .B(men_men_n423_), .C(men_men_n421_), .Y(men_men_n427_));
  AOI210     u405(.A0(men_men_n427_), .A1(men_men_n419_), .B0(men_men_n263_), .Y(men_men_n428_));
  NO4        u406(.A(men_men_n428_), .B(men_men_n412_), .C(men_men_n393_), .D(men_men_n368_), .Y(men_men_n429_));
  NO2        u407(.A(men_men_n67_), .B(i_13_), .Y(men_men_n430_));
  NA3        u408(.A(men_men_n430_), .B(i_1_), .C(i_2_), .Y(men_men_n431_));
  NO2        u409(.A(i_10_), .B(i_9_), .Y(men_men_n432_));
  NAi21      u410(.An(i_12_), .B(i_8_), .Y(men_men_n433_));
  NO2        u411(.A(men_men_n433_), .B(i_3_), .Y(men_men_n434_));
  NA2        u412(.A(men_men_n434_), .B(men_men_n432_), .Y(men_men_n435_));
  NO2        u413(.A(men_men_n47_), .B(i_4_), .Y(men_men_n436_));
  NA2        u414(.A(men_men_n436_), .B(men_men_n99_), .Y(men_men_n437_));
  OAI220     u415(.A0(men_men_n437_), .A1(men_men_n202_), .B0(men_men_n435_), .B1(men_men_n431_), .Y(men_men_n438_));
  NA2        u416(.A(men_men_n298_), .B(i_0_), .Y(men_men_n439_));
  NO3        u417(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n440_));
  NA2        u418(.A(men_men_n258_), .B(men_men_n92_), .Y(men_men_n441_));
  NA2        u419(.A(men_men_n441_), .B(men_men_n440_), .Y(men_men_n442_));
  NA2        u420(.A(i_8_), .B(i_9_), .Y(men_men_n443_));
  NA2        u421(.A(men_men_n275_), .B(men_men_n203_), .Y(men_men_n444_));
  OAI220     u422(.A0(men_men_n444_), .A1(men_men_n443_), .B0(men_men_n442_), .B1(men_men_n439_), .Y(men_men_n445_));
  NA2        u423(.A(men_men_n248_), .B(men_men_n297_), .Y(men_men_n446_));
  NO3        u424(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n447_));
  INV        u425(.A(men_men_n447_), .Y(men_men_n448_));
  NA3        u426(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n449_));
  NA4        u427(.A(men_men_n141_), .B(men_men_n111_), .C(men_men_n74_), .D(men_men_n23_), .Y(men_men_n450_));
  OAI220     u428(.A0(men_men_n450_), .A1(men_men_n449_), .B0(men_men_n448_), .B1(men_men_n446_), .Y(men_men_n451_));
  NO3        u429(.A(men_men_n451_), .B(men_men_n445_), .C(men_men_n438_), .Y(men_men_n452_));
  NA2        u430(.A(men_men_n285_), .B(men_men_n103_), .Y(men_men_n453_));
  OR2        u431(.A(men_men_n453_), .B(men_men_n206_), .Y(men_men_n454_));
  OA220      u432(.A0(men_men_n339_), .A1(men_men_n159_), .B0(men_men_n454_), .B1(men_men_n230_), .Y(men_men_n455_));
  NA2        u433(.A(men_men_n91_), .B(i_13_), .Y(men_men_n456_));
  NA2        u434(.A(men_men_n416_), .B(men_men_n369_), .Y(men_men_n457_));
  NO2        u435(.A(i_2_), .B(i_13_), .Y(men_men_n458_));
  NA3        u436(.A(men_men_n458_), .B(men_men_n158_), .C(men_men_n94_), .Y(men_men_n459_));
  NO2        u437(.A(men_men_n457_), .B(men_men_n456_), .Y(men_men_n460_));
  NO2        u438(.A(i_6_), .B(i_7_), .Y(men_men_n461_));
  NA2        u439(.A(men_men_n461_), .B(i_5_), .Y(men_men_n462_));
  NO2        u440(.A(i_11_), .B(i_1_), .Y(men_men_n463_));
  OR2        u441(.A(i_11_), .B(i_8_), .Y(men_men_n464_));
  NOi21      u442(.An(i_2_), .B(i_7_), .Y(men_men_n465_));
  NAi31      u443(.An(men_men_n464_), .B(men_men_n465_), .C(i_0_), .Y(men_men_n466_));
  NO2        u444(.A(men_men_n405_), .B(i_6_), .Y(men_men_n467_));
  NA3        u445(.A(men_men_n467_), .B(i_1_), .C(men_men_n69_), .Y(men_men_n468_));
  NO2        u446(.A(men_men_n468_), .B(men_men_n466_), .Y(men_men_n469_));
  NO2        u447(.A(i_3_), .B(men_men_n190_), .Y(men_men_n470_));
  NO2        u448(.A(i_6_), .B(i_10_), .Y(men_men_n471_));
  NA2        u449(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n472_));
  NO2        u450(.A(men_men_n154_), .B(i_3_), .Y(men_men_n473_));
  NAi31      u451(.An(men_men_n472_), .B(men_men_n473_), .C(men_men_n224_), .Y(men_men_n474_));
  NA3        u452(.A(men_men_n382_), .B(men_men_n175_), .C(men_men_n145_), .Y(men_men_n475_));
  NA2        u453(.A(men_men_n475_), .B(men_men_n474_), .Y(men_men_n476_));
  NO3        u454(.A(men_men_n476_), .B(men_men_n469_), .C(men_men_n460_), .Y(men_men_n477_));
  NA2        u455(.A(men_men_n440_), .B(men_men_n370_), .Y(men_men_n478_));
  NA2        u456(.A(men_men_n447_), .B(men_men_n377_), .Y(men_men_n479_));
  NO2        u457(.A(men_men_n479_), .B(men_men_n222_), .Y(men_men_n480_));
  NAi21      u458(.An(men_men_n216_), .B(men_men_n386_), .Y(men_men_n481_));
  NA2        u459(.A(men_men_n323_), .B(men_men_n218_), .Y(men_men_n482_));
  NO2        u460(.A(men_men_n26_), .B(i_5_), .Y(men_men_n483_));
  NO2        u461(.A(i_0_), .B(men_men_n79_), .Y(men_men_n484_));
  NA3        u462(.A(men_men_n484_), .B(men_men_n483_), .C(men_men_n138_), .Y(men_men_n485_));
  OAI220     u463(.A0(men_men_n38_), .A1(men_men_n485_), .B0(men_men_n482_), .B1(men_men_n481_), .Y(men_men_n486_));
  NA2        u464(.A(men_men_n27_), .B(i_10_), .Y(men_men_n487_));
  NO2        u465(.A(men_men_n487_), .B(men_men_n456_), .Y(men_men_n488_));
  NA4        u466(.A(men_men_n295_), .B(men_men_n221_), .C(men_men_n67_), .D(men_men_n235_), .Y(men_men_n489_));
  NO2        u467(.A(men_men_n489_), .B(men_men_n462_), .Y(men_men_n490_));
  NO4        u468(.A(men_men_n490_), .B(men_men_n488_), .C(men_men_n486_), .D(men_men_n480_), .Y(men_men_n491_));
  NA4        u469(.A(men_men_n491_), .B(men_men_n477_), .C(men_men_n455_), .D(men_men_n452_), .Y(men_men_n492_));
  AN2        u470(.A(men_men_n277_), .B(men_men_n232_), .Y(men_men_n493_));
  NA2        u471(.A(men_men_n493_), .B(men_men_n172_), .Y(men_men_n494_));
  NA2        u472(.A(men_men_n118_), .B(men_men_n107_), .Y(men_men_n495_));
  AN2        u473(.A(men_men_n495_), .B(men_men_n440_), .Y(men_men_n496_));
  OAI210     u474(.A0(i_2_), .A1(men_men_n230_), .B0(men_men_n296_), .Y(men_men_n497_));
  AOI220     u475(.A0(men_men_n497_), .A1(men_men_n311_), .B0(men_men_n496_), .B1(men_men_n298_), .Y(men_men_n498_));
  NA4        u476(.A(men_men_n430_), .B(i_1_), .C(men_men_n200_), .D(i_2_), .Y(men_men_n499_));
  INV        u477(.A(men_men_n499_), .Y(men_men_n500_));
  NA2        u478(.A(men_men_n343_), .B(men_men_n67_), .Y(men_men_n501_));
  NA2        u479(.A(men_men_n357_), .B(men_men_n350_), .Y(men_men_n502_));
  NO2        u480(.A(men_men_n36_), .B(i_8_), .Y(men_men_n503_));
  NA2        u481(.A(men_men_n39_), .B(i_13_), .Y(men_men_n504_));
  INV        u482(.A(men_men_n504_), .Y(men_men_n505_));
  AOI210     u483(.A0(men_men_n500_), .A1(men_men_n201_), .B0(men_men_n505_), .Y(men_men_n506_));
  OAI210     u484(.A0(i_8_), .A1(men_men_n61_), .B0(men_men_n130_), .Y(men_men_n507_));
  AOI210     u485(.A0(men_men_n191_), .A1(i_9_), .B0(men_men_n257_), .Y(men_men_n508_));
  NO2        u486(.A(men_men_n508_), .B(men_men_n196_), .Y(men_men_n509_));
  AOI220     u487(.A0(i_6_), .A1(men_men_n509_), .B0(men_men_n507_), .B1(men_men_n406_), .Y(men_men_n510_));
  NA4        u488(.A(men_men_n510_), .B(men_men_n506_), .C(men_men_n498_), .D(men_men_n494_), .Y(men_men_n511_));
  INV        u489(.A(men_men_n376_), .Y(men_men_n512_));
  OAI210     u490(.A0(men_men_n372_), .A1(i_0_), .B0(men_men_n512_), .Y(men_men_n513_));
  NO2        u491(.A(i_12_), .B(men_men_n190_), .Y(men_men_n514_));
  NA2        u492(.A(men_men_n514_), .B(men_men_n223_), .Y(men_men_n515_));
  NO3        u493(.A(i_10_), .B(men_men_n515_), .C(men_men_n453_), .Y(men_men_n516_));
  NOi21      u494(.An(men_men_n304_), .B(men_men_n38_), .Y(men_men_n517_));
  OAI210     u495(.A0(men_men_n517_), .A1(men_men_n516_), .B0(men_men_n513_), .Y(men_men_n518_));
  NO2        u496(.A(i_8_), .B(i_7_), .Y(men_men_n519_));
  OAI210     u497(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n520_));
  NA2        u498(.A(men_men_n520_), .B(men_men_n221_), .Y(men_men_n521_));
  AOI220     u499(.A0(men_men_n312_), .A1(men_men_n40_), .B0(men_men_n233_), .B1(men_men_n205_), .Y(men_men_n522_));
  OAI220     u500(.A0(men_men_n522_), .A1(men_men_n179_), .B0(men_men_n521_), .B1(men_men_n240_), .Y(men_men_n523_));
  NO2        u501(.A(men_men_n974_), .B(i_6_), .Y(men_men_n524_));
  NA3        u502(.A(men_men_n524_), .B(men_men_n523_), .C(men_men_n519_), .Y(men_men_n525_));
  NA2        u503(.A(men_men_n416_), .B(men_men_n312_), .Y(men_men_n526_));
  OAI220     u504(.A0(men_men_n526_), .A1(men_men_n254_), .B0(men_men_n456_), .B1(men_men_n129_), .Y(men_men_n527_));
  NA2        u505(.A(men_men_n527_), .B(men_men_n257_), .Y(men_men_n528_));
  NOi31      u506(.An(men_men_n281_), .B(men_men_n291_), .C(men_men_n177_), .Y(men_men_n529_));
  NA3        u507(.A(men_men_n295_), .B(men_men_n170_), .C(men_men_n91_), .Y(men_men_n530_));
  NO2        u508(.A(men_men_n154_), .B(i_5_), .Y(men_men_n531_));
  NA3        u509(.A(men_men_n531_), .B(men_men_n394_), .C(men_men_n306_), .Y(men_men_n532_));
  INV        u510(.A(men_men_n532_), .Y(men_men_n533_));
  OAI210     u511(.A0(men_men_n533_), .A1(men_men_n529_), .B0(men_men_n447_), .Y(men_men_n534_));
  NA4        u512(.A(men_men_n534_), .B(men_men_n528_), .C(men_men_n525_), .D(men_men_n518_), .Y(men_men_n535_));
  NA2        u513(.A(men_men_n275_), .B(men_men_n77_), .Y(men_men_n536_));
  NO2        u514(.A(men_men_n334_), .B(men_men_n536_), .Y(men_men_n537_));
  INV        u515(.A(men_men_n277_), .Y(men_men_n538_));
  NO2        u516(.A(men_men_n538_), .B(men_men_n169_), .Y(men_men_n539_));
  NO2        u517(.A(men_men_n47_), .B(men_men_n354_), .Y(men_men_n540_));
  NA2        u518(.A(men_men_n514_), .B(men_men_n267_), .Y(men_men_n541_));
  NO2        u519(.A(men_men_n540_), .B(men_men_n541_), .Y(men_men_n542_));
  NO3        u520(.A(men_men_n542_), .B(men_men_n539_), .C(men_men_n537_), .Y(men_men_n543_));
  NO3        u521(.A(men_men_n43_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n544_));
  NO3        u522(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n545_));
  NO2        u523(.A(men_men_n231_), .B(men_men_n36_), .Y(men_men_n546_));
  AN2        u524(.A(men_men_n546_), .B(men_men_n545_), .Y(men_men_n547_));
  OA210      u525(.A0(men_men_n547_), .A1(men_men_n544_), .B0(men_men_n343_), .Y(men_men_n548_));
  NO2        u526(.A(men_men_n405_), .B(i_1_), .Y(men_men_n549_));
  NOi31      u527(.An(men_men_n549_), .B(men_men_n441_), .C(men_men_n67_), .Y(men_men_n550_));
  AN4        u528(.A(men_men_n550_), .B(men_men_n403_), .C(men_men_n483_), .D(i_2_), .Y(men_men_n551_));
  NO2        u529(.A(men_men_n414_), .B(men_men_n173_), .Y(men_men_n552_));
  NO3        u530(.A(men_men_n552_), .B(men_men_n551_), .C(men_men_n548_), .Y(men_men_n553_));
  NOi21      u531(.An(i_10_), .B(i_6_), .Y(men_men_n554_));
  NO2        u532(.A(men_men_n79_), .B(men_men_n25_), .Y(men_men_n555_));
  AOI220     u533(.A0(men_men_n275_), .A1(men_men_n555_), .B0(men_men_n267_), .B1(men_men_n554_), .Y(men_men_n556_));
  NO2        u534(.A(men_men_n556_), .B(men_men_n439_), .Y(men_men_n557_));
  NO2        u535(.A(men_men_n110_), .B(men_men_n23_), .Y(men_men_n558_));
  NA2        u536(.A(men_men_n304_), .B(men_men_n161_), .Y(men_men_n559_));
  AOI220     u537(.A0(men_men_n559_), .A1(men_men_n422_), .B0(men_men_n180_), .B1(men_men_n178_), .Y(men_men_n560_));
  NO2        u538(.A(men_men_n195_), .B(men_men_n37_), .Y(men_men_n561_));
  NOi31      u539(.An(men_men_n142_), .B(men_men_n561_), .C(men_men_n320_), .Y(men_men_n562_));
  NO3        u540(.A(men_men_n562_), .B(men_men_n560_), .C(men_men_n557_), .Y(men_men_n563_));
  NO2        u541(.A(men_men_n501_), .B(men_men_n365_), .Y(men_men_n564_));
  INV        u542(.A(men_men_n306_), .Y(men_men_n565_));
  NA2        u543(.A(men_men_n973_), .B(men_men_n267_), .Y(men_men_n566_));
  NA3        u544(.A(men_men_n373_), .B(men_men_n275_), .C(men_men_n218_), .Y(men_men_n567_));
  AOI210     u545(.A0(men_men_n567_), .A1(men_men_n566_), .B0(men_men_n565_), .Y(men_men_n568_));
  NO3        u546(.A(i_4_), .B(men_men_n329_), .C(men_men_n291_), .Y(men_men_n569_));
  OR2        u547(.A(i_2_), .B(i_5_), .Y(men_men_n570_));
  BUFFER     u548(.A(men_men_n570_), .Y(men_men_n571_));
  NO3        u549(.A(men_men_n569_), .B(men_men_n568_), .C(men_men_n564_), .Y(men_men_n572_));
  NA4        u550(.A(men_men_n572_), .B(men_men_n563_), .C(men_men_n553_), .D(men_men_n543_), .Y(men_men_n573_));
  NO4        u551(.A(men_men_n573_), .B(men_men_n535_), .C(men_men_n511_), .D(men_men_n492_), .Y(men_men_n574_));
  NA4        u552(.A(men_men_n574_), .B(men_men_n429_), .C(men_men_n342_), .D(men_men_n301_), .Y(men7));
  NO2        u553(.A(men_men_n103_), .B(men_men_n84_), .Y(men_men_n576_));
  NA2        u554(.A(men_men_n371_), .B(men_men_n576_), .Y(men_men_n577_));
  NA2        u555(.A(men_men_n471_), .B(men_men_n77_), .Y(men_men_n578_));
  NA2        u556(.A(i_11_), .B(men_men_n190_), .Y(men_men_n579_));
  OAI210     u557(.A0(men_men_n970_), .A1(men_men_n578_), .B0(men_men_n577_), .Y(men_men_n580_));
  NA3        u558(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n581_));
  NO2        u559(.A(men_men_n235_), .B(i_4_), .Y(men_men_n582_));
  NA2        u560(.A(men_men_n582_), .B(i_8_), .Y(men_men_n583_));
  NO2        u561(.A(men_men_n100_), .B(men_men_n581_), .Y(men_men_n584_));
  NA2        u562(.A(i_2_), .B(men_men_n79_), .Y(men_men_n585_));
  OAI210     u563(.A0(men_men_n82_), .A1(men_men_n200_), .B0(men_men_n201_), .Y(men_men_n586_));
  NO2        u564(.A(i_7_), .B(men_men_n37_), .Y(men_men_n587_));
  NA2        u565(.A(i_4_), .B(i_8_), .Y(men_men_n588_));
  AOI210     u566(.A0(men_men_n588_), .A1(men_men_n295_), .B0(men_men_n587_), .Y(men_men_n589_));
  OAI220     u567(.A0(men_men_n589_), .A1(men_men_n585_), .B0(men_men_n586_), .B1(i_13_), .Y(men_men_n590_));
  NO3        u568(.A(men_men_n590_), .B(men_men_n584_), .C(men_men_n580_), .Y(men_men_n591_));
  AOI210     u569(.A0(men_men_n124_), .A1(men_men_n60_), .B0(i_10_), .Y(men_men_n592_));
  AOI210     u570(.A0(men_men_n592_), .A1(men_men_n235_), .B0(men_men_n158_), .Y(men_men_n593_));
  NO2        u571(.A(i_10_), .B(men_men_n23_), .Y(men_men_n594_));
  OR3        u572(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n595_));
  NO3        u573(.A(men_men_n595_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n596_));
  INV        u574(.A(men_men_n197_), .Y(men_men_n597_));
  OA220      u575(.A0(men_men_n595_), .A1(men_men_n565_), .B0(men_men_n593_), .B1(men_men_n259_), .Y(men_men_n598_));
  AOI210     u576(.A0(men_men_n598_), .A1(men_men_n591_), .B0(men_men_n61_), .Y(men_men_n599_));
  NOi21      u577(.An(i_11_), .B(i_7_), .Y(men_men_n600_));
  AO210      u578(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n601_));
  NO2        u579(.A(men_men_n601_), .B(men_men_n600_), .Y(men_men_n602_));
  NA3        u580(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n603_));
  NO2        u581(.A(men_men_n603_), .B(men_men_n61_), .Y(men_men_n604_));
  AO210      u582(.A0(men_men_n80_), .A1(men_men_n365_), .B0(men_men_n41_), .Y(men_men_n605_));
  NA2        u583(.A(men_men_n61_), .B(men_men_n977_), .Y(men_men_n606_));
  NA2        u584(.A(men_men_n606_), .B(men_men_n605_), .Y(men_men_n607_));
  OAI210     u585(.A0(men_men_n607_), .A1(men_men_n604_), .B0(i_6_), .Y(men_men_n608_));
  NO2        u586(.A(i_6_), .B(i_11_), .Y(men_men_n609_));
  NO4        u587(.A(men_men_n215_), .B(men_men_n124_), .C(i_13_), .D(men_men_n79_), .Y(men_men_n610_));
  NA3        u588(.A(men_men_n519_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n611_));
  NA2        u589(.A(men_men_n134_), .B(i_9_), .Y(men_men_n612_));
  NO2        u590(.A(men_men_n612_), .B(men_men_n964_), .Y(men_men_n613_));
  NA3        u591(.A(i_1_), .B(men_men_n306_), .C(i_6_), .Y(men_men_n614_));
  AOI210     u592(.A0(men_men_n463_), .A1(men_men_n408_), .B0(men_men_n239_), .Y(men_men_n615_));
  NO2        u593(.A(men_men_n615_), .B(men_men_n585_), .Y(men_men_n616_));
  NAi21      u594(.An(men_men_n611_), .B(men_men_n86_), .Y(men_men_n617_));
  NO2        u595(.A(i_11_), .B(men_men_n37_), .Y(men_men_n618_));
  NA2        u596(.A(men_men_n618_), .B(men_men_n24_), .Y(men_men_n619_));
  OAI210     u597(.A0(men_men_n619_), .A1(i_6_), .B0(men_men_n617_), .Y(men_men_n620_));
  OR3        u598(.A(men_men_n620_), .B(men_men_n616_), .C(men_men_n613_), .Y(men_men_n621_));
  NO2        u599(.A(men_men_n621_), .B(men_men_n610_), .Y(men_men_n622_));
  NA2        u600(.A(i_3_), .B(men_men_n190_), .Y(men_men_n623_));
  NO2        u601(.A(men_men_n113_), .B(men_men_n37_), .Y(men_men_n624_));
  NO2        u602(.A(men_men_n79_), .B(i_9_), .Y(men_men_n625_));
  NA2        u603(.A(i_1_), .B(i_3_), .Y(men_men_n626_));
  NA2        u604(.A(men_men_n622_), .B(men_men_n608_), .Y(men_men_n627_));
  NO3        u605(.A(men_men_n464_), .B(i_3_), .C(i_7_), .Y(men_men_n628_));
  OA210      u606(.A0(men_men_n628_), .A1(men_men_n242_), .B0(men_men_n79_), .Y(men_men_n629_));
  NA3        u607(.A(men_men_n471_), .B(men_men_n503_), .C(men_men_n47_), .Y(men_men_n630_));
  NO3        u608(.A(men_men_n465_), .B(men_men_n588_), .C(men_men_n79_), .Y(men_men_n631_));
  NA2        u609(.A(men_men_n631_), .B(men_men_n25_), .Y(men_men_n632_));
  NA3        u610(.A(men_men_n158_), .B(men_men_n77_), .C(men_men_n79_), .Y(men_men_n633_));
  NA3        u611(.A(men_men_n633_), .B(men_men_n632_), .C(men_men_n630_), .Y(men_men_n634_));
  OAI210     u612(.A0(men_men_n634_), .A1(men_men_n629_), .B0(i_1_), .Y(men_men_n635_));
  AOI210     u613(.A0(men_men_n258_), .A1(men_men_n92_), .B0(i_1_), .Y(men_men_n636_));
  NO2        u614(.A(men_men_n355_), .B(i_2_), .Y(men_men_n637_));
  NA2        u615(.A(men_men_n637_), .B(men_men_n636_), .Y(men_men_n638_));
  NA2        u616(.A(men_men_n614_), .B(men_men_n638_), .Y(men_men_n639_));
  INV        u617(.A(men_men_n639_), .Y(men_men_n640_));
  AOI210     u618(.A0(men_men_n640_), .A1(men_men_n635_), .B0(i_13_), .Y(men_men_n641_));
  OR2        u619(.A(i_11_), .B(i_7_), .Y(men_men_n642_));
  NA2        u620(.A(men_men_n101_), .B(men_men_n134_), .Y(men_men_n643_));
  AOI220     u621(.A0(men_men_n458_), .A1(men_men_n158_), .B0(men_men_n436_), .B1(men_men_n134_), .Y(men_men_n644_));
  OAI210     u622(.A0(men_men_n644_), .A1(men_men_n45_), .B0(men_men_n643_), .Y(men_men_n645_));
  NO2        u623(.A(men_men_n55_), .B(i_12_), .Y(men_men_n646_));
  NO2        u624(.A(men_men_n465_), .B(men_men_n24_), .Y(men_men_n647_));
  NO2        u625(.A(men_men_n963_), .B(men_men_n87_), .Y(men_men_n648_));
  AOI210     u626(.A0(men_men_n645_), .A1(men_men_n322_), .B0(men_men_n648_), .Y(men_men_n649_));
  AOI220     u627(.A0(i_12_), .A1(men_men_n66_), .B0(men_men_n373_), .B1(men_men_n975_), .Y(men_men_n650_));
  NO2        u628(.A(men_men_n650_), .B(men_men_n240_), .Y(men_men_n651_));
  AOI210     u629(.A0(men_men_n433_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n652_));
  NOi31      u630(.An(men_men_n652_), .B(men_men_n578_), .C(men_men_n45_), .Y(men_men_n653_));
  NA2        u631(.A(men_men_n123_), .B(i_13_), .Y(men_men_n654_));
  NO2        u632(.A(men_men_n654_), .B(men_men_n636_), .Y(men_men_n655_));
  NO3        u633(.A(men_men_n65_), .B(men_men_n32_), .C(men_men_n96_), .Y(men_men_n656_));
  NA2        u634(.A(men_men_n26_), .B(men_men_n190_), .Y(men_men_n657_));
  NA2        u635(.A(men_men_n657_), .B(i_7_), .Y(men_men_n658_));
  NO3        u636(.A(men_men_n465_), .B(men_men_n235_), .C(men_men_n79_), .Y(men_men_n659_));
  AOI210     u637(.A0(men_men_n659_), .A1(men_men_n658_), .B0(men_men_n656_), .Y(men_men_n660_));
  AOI220     u638(.A0(men_men_n373_), .A1(men_men_n975_), .B0(men_men_n86_), .B1(men_men_n97_), .Y(men_men_n661_));
  OAI220     u639(.A0(men_men_n661_), .A1(men_men_n583_), .B0(men_men_n660_), .B1(men_men_n597_), .Y(men_men_n662_));
  NO4        u640(.A(men_men_n662_), .B(men_men_n655_), .C(men_men_n653_), .D(men_men_n651_), .Y(men_men_n663_));
  NA2        u641(.A(men_men_n609_), .B(i_13_), .Y(men_men_n664_));
  NAi21      u642(.An(i_11_), .B(i_12_), .Y(men_men_n665_));
  NA2        u643(.A(men_men_n972_), .B(men_men_n302_), .Y(men_men_n666_));
  NA2        u644(.A(men_men_n666_), .B(men_men_n664_), .Y(men_men_n667_));
  NA2        u645(.A(men_men_n667_), .B(men_men_n61_), .Y(men_men_n668_));
  NO2        u646(.A(i_2_), .B(i_12_), .Y(men_men_n669_));
  NA2        u647(.A(men_men_n354_), .B(men_men_n669_), .Y(men_men_n670_));
  NA2        u648(.A(i_8_), .B(men_men_n25_), .Y(men_men_n671_));
  NO3        u649(.A(men_men_n671_), .B(men_men_n371_), .C(men_men_n582_), .Y(men_men_n672_));
  OAI210     u650(.A0(men_men_n672_), .A1(men_men_n356_), .B0(men_men_n354_), .Y(men_men_n673_));
  NA2        u651(.A(men_men_n673_), .B(men_men_n670_), .Y(men_men_n674_));
  NA3        u652(.A(men_men_n674_), .B(men_men_n46_), .C(men_men_n223_), .Y(men_men_n675_));
  NA4        u653(.A(men_men_n675_), .B(men_men_n668_), .C(men_men_n663_), .D(men_men_n649_), .Y(men_men_n676_));
  OR4        u654(.A(men_men_n676_), .B(men_men_n641_), .C(men_men_n627_), .D(men_men_n599_), .Y(men5));
  AN2        u655(.A(men_men_n24_), .B(i_10_), .Y(men_men_n678_));
  NA3        u656(.A(men_men_n678_), .B(men_men_n669_), .C(men_men_n103_), .Y(men_men_n679_));
  NO2        u657(.A(men_men_n583_), .B(i_11_), .Y(men_men_n680_));
  NA2        u658(.A(men_men_n82_), .B(men_men_n680_), .Y(men_men_n681_));
  NA2        u659(.A(men_men_n681_), .B(men_men_n679_), .Y(men_men_n682_));
  NO3        u660(.A(i_11_), .B(men_men_n235_), .C(i_13_), .Y(men_men_n683_));
  NO2        u661(.A(men_men_n120_), .B(men_men_n23_), .Y(men_men_n684_));
  NA2        u662(.A(i_12_), .B(i_8_), .Y(men_men_n685_));
  OAI210     u663(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n685_), .Y(men_men_n686_));
  INV        u664(.A(men_men_n432_), .Y(men_men_n687_));
  AOI220     u665(.A0(men_men_n306_), .A1(men_men_n558_), .B0(men_men_n686_), .B1(men_men_n684_), .Y(men_men_n688_));
  INV        u666(.A(men_men_n688_), .Y(men_men_n689_));
  NO2        u667(.A(men_men_n689_), .B(men_men_n682_), .Y(men_men_n690_));
  INV        u668(.A(men_men_n167_), .Y(men_men_n691_));
  OAI210     u669(.A0(men_men_n637_), .A1(men_men_n434_), .B0(men_men_n106_), .Y(men_men_n692_));
  NO2        u670(.A(men_men_n692_), .B(men_men_n691_), .Y(men_men_n693_));
  NO2        u671(.A(men_men_n443_), .B(men_men_n26_), .Y(men_men_n694_));
  NO2        u672(.A(men_men_n187_), .B(men_men_n121_), .Y(men_men_n695_));
  OAI210     u673(.A0(men_men_n695_), .A1(men_men_n684_), .B0(i_2_), .Y(men_men_n696_));
  INV        u674(.A(men_men_n168_), .Y(men_men_n697_));
  NO3        u675(.A(men_men_n601_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n698_));
  AOI210     u676(.A0(men_men_n697_), .A1(men_men_n82_), .B0(men_men_n698_), .Y(men_men_n699_));
  AOI210     u677(.A0(men_men_n699_), .A1(men_men_n696_), .B0(men_men_n190_), .Y(men_men_n700_));
  OA210      u678(.A0(men_men_n602_), .A1(men_men_n122_), .B0(i_13_), .Y(men_men_n701_));
  NA2        u679(.A(men_men_n197_), .B(men_men_n200_), .Y(men_men_n702_));
  NA2        u680(.A(men_men_n148_), .B(men_men_n579_), .Y(men_men_n703_));
  AOI210     u681(.A0(men_men_n703_), .A1(men_men_n702_), .B0(men_men_n359_), .Y(men_men_n704_));
  AOI210     u682(.A0(men_men_n207_), .A1(men_men_n144_), .B0(men_men_n503_), .Y(men_men_n705_));
  NA2        u683(.A(men_men_n705_), .B(men_men_n408_), .Y(men_men_n706_));
  NO2        u684(.A(men_men_n97_), .B(men_men_n45_), .Y(men_men_n707_));
  INV        u685(.A(men_men_n292_), .Y(men_men_n708_));
  NA4        u686(.A(men_men_n708_), .B(men_men_n295_), .C(men_men_n120_), .D(men_men_n43_), .Y(men_men_n709_));
  OAI210     u687(.A0(men_men_n709_), .A1(men_men_n707_), .B0(men_men_n706_), .Y(men_men_n710_));
  NO4        u688(.A(men_men_n710_), .B(men_men_n704_), .C(men_men_n701_), .D(men_men_n700_), .Y(men_men_n711_));
  NA2        u689(.A(men_men_n558_), .B(men_men_n28_), .Y(men_men_n712_));
  NA2        u690(.A(men_men_n683_), .B(men_men_n268_), .Y(men_men_n713_));
  NA2        u691(.A(men_men_n713_), .B(men_men_n712_), .Y(men_men_n714_));
  NO2        u692(.A(men_men_n60_), .B(i_12_), .Y(men_men_n715_));
  NO2        u693(.A(men_men_n715_), .B(men_men_n122_), .Y(men_men_n716_));
  NO2        u694(.A(men_men_n716_), .B(men_men_n579_), .Y(men_men_n717_));
  AOI220     u695(.A0(men_men_n717_), .A1(men_men_n36_), .B0(men_men_n714_), .B1(men_men_n47_), .Y(men_men_n718_));
  NA4        u696(.A(men_men_n718_), .B(men_men_n711_), .C(men_men_n976_), .D(men_men_n690_), .Y(men6));
  NO3        u697(.A(i_9_), .B(men_men_n297_), .C(i_1_), .Y(men_men_n720_));
  NO2        u698(.A(men_men_n182_), .B(men_men_n135_), .Y(men_men_n721_));
  OAI210     u699(.A0(men_men_n721_), .A1(men_men_n720_), .B0(men_men_n967_), .Y(men_men_n722_));
  NA4        u700(.A(men_men_n377_), .B(men_men_n470_), .C(men_men_n65_), .D(men_men_n96_), .Y(men_men_n723_));
  INV        u701(.A(men_men_n723_), .Y(men_men_n724_));
  NO2        u702(.A(men_men_n220_), .B(men_men_n472_), .Y(men_men_n725_));
  NO2        u703(.A(i_11_), .B(i_9_), .Y(men_men_n726_));
  NO2        u704(.A(men_men_n724_), .B(men_men_n317_), .Y(men_men_n727_));
  AO210      u705(.A0(men_men_n727_), .A1(men_men_n722_), .B0(i_12_), .Y(men_men_n728_));
  NA2        u706(.A(men_men_n360_), .B(men_men_n323_), .Y(men_men_n729_));
  NA2        u707(.A(men_men_n628_), .B(men_men_n65_), .Y(men_men_n730_));
  NA3        u708(.A(men_men_n80_), .B(men_men_n730_), .C(men_men_n729_), .Y(men_men_n731_));
  INV        u709(.A(men_men_n194_), .Y(men_men_n732_));
  AOI220     u710(.A0(men_men_n732_), .A1(men_men_n726_), .B0(men_men_n731_), .B1(men_men_n67_), .Y(men_men_n733_));
  INV        u711(.A(men_men_n316_), .Y(men_men_n734_));
  NA2        u712(.A(men_men_n69_), .B(men_men_n127_), .Y(men_men_n735_));
  NA2        u713(.A(men_men_n25_), .B(men_men_n47_), .Y(men_men_n736_));
  AOI210     u714(.A0(men_men_n736_), .A1(men_men_n735_), .B0(men_men_n734_), .Y(men_men_n737_));
  NO2        u715(.A(men_men_n32_), .B(i_11_), .Y(men_men_n738_));
  NA3        u716(.A(men_men_n738_), .B(men_men_n461_), .C(men_men_n377_), .Y(men_men_n739_));
  OAI210     u717(.A0(men_men_n628_), .A1(men_men_n546_), .B0(men_men_n545_), .Y(men_men_n740_));
  NA2        u718(.A(men_men_n740_), .B(men_men_n739_), .Y(men_men_n741_));
  OR2        u719(.A(men_men_n741_), .B(men_men_n737_), .Y(men_men_n742_));
  NO2        u720(.A(men_men_n642_), .B(i_2_), .Y(men_men_n743_));
  NA2        u721(.A(men_men_n37_), .B(men_men_n743_), .Y(men_men_n744_));
  NA3        u722(.A(men_men_n338_), .B(men_men_n251_), .C(i_7_), .Y(men_men_n745_));
  BUFFER     u723(.A(men_men_n602_), .Y(men_men_n746_));
  NA2        u724(.A(men_men_n746_), .B(men_men_n143_), .Y(men_men_n747_));
  AO210      u725(.A0(men_men_n479_), .A1(men_men_n687_), .B0(men_men_n36_), .Y(men_men_n748_));
  NA4        u726(.A(men_men_n748_), .B(men_men_n747_), .C(men_men_n745_), .D(men_men_n744_), .Y(men_men_n749_));
  OAI210     u727(.A0(i_6_), .A1(i_11_), .B0(men_men_n80_), .Y(men_men_n750_));
  AOI220     u728(.A0(men_men_n750_), .A1(men_men_n545_), .B0(men_men_n725_), .B1(men_men_n658_), .Y(men_men_n751_));
  NA3        u729(.A(men_men_n359_), .B(men_men_n236_), .C(men_men_n143_), .Y(men_men_n752_));
  NA2        u730(.A(men_men_n385_), .B(men_men_n64_), .Y(men_men_n753_));
  NA3        u731(.A(men_men_n753_), .B(men_men_n752_), .C(men_men_n751_), .Y(men_men_n754_));
  AO210      u732(.A0(men_men_n503_), .A1(men_men_n47_), .B0(men_men_n81_), .Y(men_men_n755_));
  NA3        u733(.A(men_men_n755_), .B(men_men_n471_), .C(men_men_n218_), .Y(men_men_n756_));
  INV        u734(.A(men_men_n544_), .Y(men_men_n757_));
  NA2        u735(.A(men_men_n107_), .B(men_men_n396_), .Y(men_men_n758_));
  NA2        u736(.A(men_men_n241_), .B(men_men_n47_), .Y(men_men_n759_));
  INV        u737(.A(men_men_n571_), .Y(men_men_n760_));
  NA3        u738(.A(men_men_n760_), .B(men_men_n316_), .C(i_7_), .Y(men_men_n761_));
  NA4        u739(.A(men_men_n761_), .B(men_men_n758_), .C(men_men_n757_), .D(men_men_n756_), .Y(men_men_n762_));
  NO4        u740(.A(men_men_n762_), .B(men_men_n754_), .C(men_men_n749_), .D(men_men_n742_), .Y(men_men_n763_));
  NA4        u741(.A(men_men_n763_), .B(men_men_n733_), .C(men_men_n728_), .D(men_men_n367_), .Y(men3));
  NA2        u742(.A(i_6_), .B(i_7_), .Y(men_men_n765_));
  NO2        u743(.A(men_men_n765_), .B(i_0_), .Y(men_men_n766_));
  NO2        u744(.A(i_11_), .B(men_men_n235_), .Y(men_men_n767_));
  OAI210     u745(.A0(men_men_n766_), .A1(men_men_n281_), .B0(men_men_n767_), .Y(men_men_n768_));
  NO2        u746(.A(men_men_n768_), .B(men_men_n190_), .Y(men_men_n769_));
  NO3        u747(.A(men_men_n439_), .B(men_men_n84_), .C(men_men_n45_), .Y(men_men_n770_));
  OA210      u748(.A0(men_men_n770_), .A1(men_men_n769_), .B0(men_men_n170_), .Y(men_men_n771_));
  NA3        u749(.A(men_men_n752_), .B(men_men_n586_), .C(men_men_n358_), .Y(men_men_n772_));
  NA2        u750(.A(men_men_n772_), .B(men_men_n40_), .Y(men_men_n773_));
  AN2        u751(.A(men_men_n441_), .B(men_men_n56_), .Y(men_men_n774_));
  AOI210     u752(.A0(men_men_n965_), .A1(men_men_n773_), .B0(men_men_n49_), .Y(men_men_n775_));
  NO4        u753(.A(men_men_n363_), .B(men_men_n370_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n776_));
  NA2        u754(.A(men_men_n182_), .B(men_men_n554_), .Y(men_men_n777_));
  NOi21      u755(.An(men_men_n777_), .B(men_men_n776_), .Y(men_men_n778_));
  NA2        u756(.A(men_men_n652_), .B(men_men_n625_), .Y(men_men_n779_));
  NA2        u757(.A(i_0_), .B(men_men_n424_), .Y(men_men_n780_));
  OAI220     u758(.A0(men_men_n780_), .A1(men_men_n779_), .B0(men_men_n778_), .B1(men_men_n61_), .Y(men_men_n781_));
  NOi21      u759(.An(i_5_), .B(i_9_), .Y(men_men_n782_));
  NA2        u760(.A(men_men_n782_), .B(men_men_n430_), .Y(men_men_n783_));
  NO3        u761(.A(men_men_n402_), .B(men_men_n258_), .C(men_men_n67_), .Y(men_men_n784_));
  INV        u762(.A(men_men_n784_), .Y(men_men_n785_));
  OAI220     u763(.A0(men_men_n785_), .A1(men_men_n177_), .B0(men_men_n588_), .B1(men_men_n783_), .Y(men_men_n786_));
  NO4        u764(.A(men_men_n786_), .B(men_men_n781_), .C(men_men_n775_), .D(men_men_n771_), .Y(men_men_n787_));
  NA2        u765(.A(men_men_n182_), .B(men_men_n24_), .Y(men_men_n788_));
  NO2        u766(.A(men_men_n624_), .B(men_men_n576_), .Y(men_men_n789_));
  NO2        u767(.A(men_men_n789_), .B(men_men_n788_), .Y(men_men_n790_));
  NA2        u768(.A(men_men_n302_), .B(men_men_n125_), .Y(men_men_n791_));
  NAi21      u769(.An(men_men_n159_), .B(men_men_n424_), .Y(men_men_n792_));
  OAI220     u770(.A0(men_men_n792_), .A1(men_men_n759_), .B0(men_men_n791_), .B1(men_men_n387_), .Y(men_men_n793_));
  NO2        u771(.A(men_men_n793_), .B(men_men_n790_), .Y(men_men_n794_));
  NA2        u772(.A(men_men_n555_), .B(i_0_), .Y(men_men_n795_));
  NO3        u773(.A(men_men_n795_), .B(men_men_n372_), .C(men_men_n82_), .Y(men_men_n796_));
  NO3        u774(.A(men_men_n570_), .B(men_men_n215_), .C(men_men_n405_), .Y(men_men_n797_));
  AOI210     u775(.A0(men_men_n797_), .A1(i_11_), .B0(men_men_n796_), .Y(men_men_n798_));
  NA2        u776(.A(men_men_n683_), .B(men_men_n317_), .Y(men_men_n799_));
  NO2        u777(.A(men_men_n619_), .B(men_men_n521_), .Y(men_men_n800_));
  NA2        u778(.A(i_0_), .B(i_10_), .Y(men_men_n801_));
  NO4        u779(.A(men_men_n110_), .B(men_men_n58_), .C(men_men_n623_), .D(i_5_), .Y(men_men_n802_));
  AN2        u780(.A(men_men_n802_), .B(men_men_n45_), .Y(men_men_n803_));
  NA2        u781(.A(men_men_n182_), .B(men_men_n77_), .Y(men_men_n804_));
  NA2        u782(.A(men_men_n549_), .B(i_4_), .Y(men_men_n805_));
  NA2        u783(.A(men_men_n185_), .B(men_men_n200_), .Y(men_men_n806_));
  OAI220     u784(.A0(men_men_n806_), .A1(men_men_n799_), .B0(men_men_n805_), .B1(men_men_n804_), .Y(men_men_n807_));
  NO3        u785(.A(men_men_n807_), .B(men_men_n803_), .C(men_men_n800_), .Y(men_men_n808_));
  NA3        u786(.A(men_men_n808_), .B(men_men_n798_), .C(men_men_n794_), .Y(men_men_n809_));
  NA2        u787(.A(i_11_), .B(i_9_), .Y(men_men_n810_));
  NO3        u788(.A(i_12_), .B(men_men_n810_), .C(men_men_n585_), .Y(men_men_n811_));
  AN2        u789(.A(men_men_n811_), .B(i_0_), .Y(men_men_n812_));
  NO2        u790(.A(men_men_n49_), .B(i_7_), .Y(men_men_n813_));
  NA2        u791(.A(men_men_n382_), .B(men_men_n175_), .Y(men_men_n814_));
  NA2        u792(.A(men_men_n814_), .B(men_men_n157_), .Y(men_men_n815_));
  NO2        u793(.A(men_men_n810_), .B(men_men_n67_), .Y(men_men_n816_));
  NO2        u794(.A(men_men_n171_), .B(i_0_), .Y(men_men_n817_));
  INV        u795(.A(men_men_n817_), .Y(men_men_n818_));
  NA2        u796(.A(men_men_n461_), .B(men_men_n229_), .Y(men_men_n819_));
  AOI210     u797(.A0(men_men_n357_), .A1(men_men_n42_), .B0(men_men_n395_), .Y(men_men_n820_));
  OAI220     u798(.A0(men_men_n820_), .A1(men_men_n783_), .B0(men_men_n819_), .B1(men_men_n818_), .Y(men_men_n821_));
  NO3        u799(.A(men_men_n821_), .B(men_men_n815_), .C(men_men_n812_), .Y(men_men_n822_));
  NA2        u800(.A(men_men_n618_), .B(men_men_n117_), .Y(men_men_n823_));
  NO2        u801(.A(i_6_), .B(men_men_n823_), .Y(men_men_n824_));
  AOI210     u802(.A0(men_men_n433_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n825_));
  NA2        u803(.A(men_men_n167_), .B(men_men_n98_), .Y(men_men_n826_));
  NOi32      u804(.An(men_men_n825_), .Bn(men_men_n185_), .C(men_men_n826_), .Y(men_men_n827_));
  NO2        u805(.A(men_men_n827_), .B(men_men_n824_), .Y(men_men_n828_));
  OR2        u806(.A(men_men_n826_), .B(men_men_n502_), .Y(men_men_n829_));
  NO2        u807(.A(men_men_n252_), .B(men_men_n307_), .Y(men_men_n830_));
  INV        u808(.A(men_men_n665_), .Y(men_men_n831_));
  NA2        u809(.A(men_men_n831_), .B(men_men_n830_), .Y(men_men_n832_));
  NA4        u810(.A(men_men_n832_), .B(men_men_n829_), .C(men_men_n828_), .D(men_men_n822_), .Y(men_men_n833_));
  NO2        u811(.A(men_men_n788_), .B(men_men_n237_), .Y(men_men_n834_));
  AN2        u812(.A(men_men_n322_), .B(men_men_n317_), .Y(men_men_n835_));
  NA2        u813(.A(men_men_n834_), .B(i_10_), .Y(men_men_n836_));
  NA3        u814(.A(i_5_), .B(men_men_n399_), .C(men_men_n46_), .Y(men_men_n837_));
  OAI210     u815(.A0(men_men_n792_), .A1(i_7_), .B0(men_men_n837_), .Y(men_men_n838_));
  NA2        u816(.A(men_men_n816_), .B(men_men_n295_), .Y(men_men_n839_));
  NA2        u817(.A(men_men_n184_), .B(men_men_n839_), .Y(men_men_n840_));
  AOI220     u818(.A0(men_men_n840_), .A1(men_men_n461_), .B0(men_men_n838_), .B1(men_men_n67_), .Y(men_men_n841_));
  NO2        u819(.A(men_men_n69_), .B(men_men_n685_), .Y(men_men_n842_));
  AOI210     u820(.A0(men_men_n170_), .A1(men_men_n576_), .B0(men_men_n842_), .Y(men_men_n843_));
  NO2        u821(.A(men_men_n843_), .B(men_men_n48_), .Y(men_men_n844_));
  NO3        u822(.A(men_men_n570_), .B(men_men_n345_), .C(men_men_n24_), .Y(men_men_n845_));
  AOI210     u823(.A0(men_men_n647_), .A1(men_men_n531_), .B0(men_men_n845_), .Y(men_men_n846_));
  NAi21      u824(.An(i_9_), .B(i_5_), .Y(men_men_n847_));
  NO2        u825(.A(men_men_n847_), .B(men_men_n390_), .Y(men_men_n848_));
  NO2        u826(.A(men_men_n581_), .B(men_men_n100_), .Y(men_men_n849_));
  AOI220     u827(.A0(men_men_n849_), .A1(i_0_), .B0(men_men_n848_), .B1(men_men_n602_), .Y(men_men_n850_));
  OAI220     u828(.A0(men_men_n850_), .A1(men_men_n79_), .B0(men_men_n846_), .B1(men_men_n168_), .Y(men_men_n851_));
  NO2        u829(.A(men_men_n851_), .B(men_men_n844_), .Y(men_men_n852_));
  NA3        u830(.A(men_men_n852_), .B(men_men_n841_), .C(men_men_n836_), .Y(men_men_n853_));
  NO3        u831(.A(men_men_n853_), .B(men_men_n833_), .C(men_men_n809_), .Y(men_men_n854_));
  NO2        u832(.A(i_0_), .B(men_men_n665_), .Y(men_men_n855_));
  NA2        u833(.A(men_men_n67_), .B(men_men_n45_), .Y(men_men_n856_));
  NA2        u834(.A(men_men_n801_), .B(men_men_n856_), .Y(men_men_n857_));
  NO3        u835(.A(men_men_n100_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n858_));
  AO220      u836(.A0(men_men_n858_), .A1(men_men_n857_), .B0(men_men_n855_), .B1(men_men_n170_), .Y(men_men_n859_));
  NA2        u837(.A(men_men_n859_), .B(men_men_n335_), .Y(men_men_n860_));
  NA2        u838(.A(men_men_n967_), .B(men_men_n142_), .Y(men_men_n861_));
  INV        u839(.A(men_men_n861_), .Y(men_men_n862_));
  NA3        u840(.A(men_men_n862_), .B(men_men_n625_), .C(men_men_n67_), .Y(men_men_n863_));
  NO2        u841(.A(men_men_n740_), .B(men_men_n390_), .Y(men_men_n864_));
  NA3        u842(.A(men_men_n766_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n865_));
  NA2        u843(.A(men_men_n767_), .B(i_9_), .Y(men_men_n866_));
  AOI210     u844(.A0(men_men_n865_), .A1(men_men_n485_), .B0(men_men_n866_), .Y(men_men_n867_));
  OAI210     u845(.A0(men_men_n241_), .A1(i_9_), .B0(men_men_n228_), .Y(men_men_n868_));
  AOI210     u846(.A0(men_men_n868_), .A1(men_men_n795_), .B0(men_men_n150_), .Y(men_men_n869_));
  NO3        u847(.A(men_men_n869_), .B(men_men_n867_), .C(men_men_n864_), .Y(men_men_n870_));
  NA3        u848(.A(men_men_n870_), .B(men_men_n863_), .C(men_men_n860_), .Y(men_men_n871_));
  NA2        u849(.A(men_men_n835_), .B(men_men_n359_), .Y(men_men_n872_));
  AOI210     u850(.A0(men_men_n291_), .A1(men_men_n159_), .B0(men_men_n872_), .Y(men_men_n873_));
  NA3        u851(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n874_));
  NA2        u852(.A(men_men_n813_), .B(men_men_n473_), .Y(men_men_n875_));
  AOI210     u853(.A0(men_men_n874_), .A1(men_men_n159_), .B0(men_men_n875_), .Y(men_men_n876_));
  NO2        u854(.A(men_men_n876_), .B(men_men_n873_), .Y(men_men_n877_));
  NO3        u855(.A(men_men_n801_), .B(men_men_n782_), .C(men_men_n187_), .Y(men_men_n878_));
  AOI220     u856(.A0(men_men_n878_), .A1(i_11_), .B0(men_men_n550_), .B1(men_men_n69_), .Y(men_men_n879_));
  NO3        u857(.A(men_men_n209_), .B(men_men_n370_), .C(i_0_), .Y(men_men_n880_));
  OAI210     u858(.A0(men_men_n880_), .A1(men_men_n70_), .B0(i_13_), .Y(men_men_n881_));
  INV        u859(.A(men_men_n218_), .Y(men_men_n882_));
  NO2        u860(.A(i_12_), .B(men_men_n597_), .Y(men_men_n883_));
  NA3        u861(.A(men_men_n883_), .B(men_men_n968_), .C(men_men_n882_), .Y(men_men_n884_));
  NA4        u862(.A(men_men_n884_), .B(men_men_n881_), .C(men_men_n879_), .D(men_men_n877_), .Y(men_men_n885_));
  NO2        u863(.A(men_men_n240_), .B(men_men_n87_), .Y(men_men_n886_));
  AOI210     u864(.A0(men_men_n886_), .A1(men_men_n855_), .B0(men_men_n104_), .Y(men_men_n887_));
  AOI220     u865(.A0(i_7_), .A1(men_men_n473_), .B0(men_men_n766_), .B1(men_men_n160_), .Y(men_men_n888_));
  NA2        u866(.A(men_men_n338_), .B(men_men_n172_), .Y(men_men_n889_));
  OA220      u867(.A0(men_men_n889_), .A1(men_men_n888_), .B0(men_men_n887_), .B1(i_5_), .Y(men_men_n890_));
  AOI210     u868(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n171_), .Y(men_men_n891_));
  INV        u869(.A(men_men_n530_), .Y(men_men_n892_));
  NA2        u870(.A(men_men_n478_), .B(men_men_n459_), .Y(men_men_n893_));
  NO2        u871(.A(men_men_n893_), .B(men_men_n892_), .Y(men_men_n894_));
  NA3        u872(.A(men_men_n377_), .B(men_men_n167_), .C(men_men_n166_), .Y(men_men_n895_));
  NA3        u873(.A(men_men_n813_), .B(men_men_n281_), .C(men_men_n228_), .Y(men_men_n896_));
  NA2        u874(.A(men_men_n896_), .B(men_men_n895_), .Y(men_men_n897_));
  NOi31      u875(.An(men_men_n376_), .B(men_men_n856_), .C(men_men_n237_), .Y(men_men_n898_));
  NO2        u876(.A(men_men_n898_), .B(men_men_n897_), .Y(men_men_n899_));
  NA3        u877(.A(men_men_n899_), .B(men_men_n894_), .C(men_men_n890_), .Y(men_men_n900_));
  NO2        u878(.A(men_men_n79_), .B(i_5_), .Y(men_men_n901_));
  NA3        u879(.A(men_men_n767_), .B(men_men_n105_), .C(men_men_n120_), .Y(men_men_n902_));
  INV        u880(.A(men_men_n902_), .Y(men_men_n903_));
  NA2        u881(.A(men_men_n903_), .B(men_men_n901_), .Y(men_men_n904_));
  NA3        u882(.A(men_men_n295_), .B(i_5_), .C(men_men_n190_), .Y(men_men_n905_));
  INV        u883(.A(men_men_n240_), .Y(men_men_n906_));
  NO4        u884(.A(men_men_n237_), .B(men_men_n209_), .C(i_0_), .D(i_12_), .Y(men_men_n907_));
  AOI220     u885(.A0(men_men_n907_), .A1(men_men_n906_), .B0(men_men_n724_), .B1(men_men_n172_), .Y(men_men_n908_));
  AN2        u886(.A(men_men_n801_), .B(men_men_n150_), .Y(men_men_n909_));
  NO3        u887(.A(men_men_n909_), .B(i_12_), .C(men_men_n611_), .Y(men_men_n910_));
  NA2        u888(.A(men_men_n910_), .B(men_men_n218_), .Y(men_men_n911_));
  NA3        u889(.A(men_men_n93_), .B(men_men_n554_), .C(i_11_), .Y(men_men_n912_));
  NO2        u890(.A(men_men_n912_), .B(men_men_n152_), .Y(men_men_n913_));
  INV        u891(.A(men_men_n62_), .Y(men_men_n914_));
  NO2        u892(.A(men_men_n914_), .B(men_men_n905_), .Y(men_men_n915_));
  AOI210     u893(.A0(men_men_n915_), .A1(men_men_n817_), .B0(men_men_n913_), .Y(men_men_n916_));
  NA4        u894(.A(men_men_n916_), .B(men_men_n911_), .C(men_men_n908_), .D(men_men_n904_), .Y(men_men_n917_));
  NO4        u895(.A(men_men_n917_), .B(men_men_n900_), .C(men_men_n885_), .D(men_men_n871_), .Y(men_men_n918_));
  OAI210     u896(.A0(men_men_n743_), .A1(men_men_n738_), .B0(men_men_n37_), .Y(men_men_n919_));
  NA3        u897(.A(men_men_n825_), .B(men_men_n354_), .C(i_5_), .Y(men_men_n920_));
  NA3        u898(.A(men_men_n920_), .B(men_men_n919_), .C(men_men_n593_), .Y(men_men_n921_));
  NA2        u899(.A(men_men_n921_), .B(men_men_n205_), .Y(men_men_n922_));
  NA2        u900(.A(men_men_n183_), .B(men_men_n185_), .Y(men_men_n923_));
  AO210      u901(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n923_), .Y(men_men_n924_));
  OAI210     u902(.A0(men_men_n596_), .A1(men_men_n594_), .B0(men_men_n306_), .Y(men_men_n925_));
  NA2        u903(.A(men_men_n925_), .B(men_men_n924_), .Y(men_men_n926_));
  NO2        u904(.A(men_men_n449_), .B(men_men_n258_), .Y(men_men_n927_));
  NO4        u905(.A(men_men_n231_), .B(men_men_n141_), .C(men_men_n626_), .D(men_men_n37_), .Y(men_men_n928_));
  NO3        u906(.A(men_men_n928_), .B(men_men_n927_), .C(men_men_n797_), .Y(men_men_n929_));
  OAI210     u907(.A0(men_men_n912_), .A1(men_men_n144_), .B0(men_men_n929_), .Y(men_men_n930_));
  AOI210     u908(.A0(men_men_n926_), .A1(men_men_n49_), .B0(men_men_n930_), .Y(men_men_n931_));
  AOI210     u909(.A0(men_men_n931_), .A1(men_men_n922_), .B0(men_men_n67_), .Y(men_men_n932_));
  NO2        u910(.A(men_men_n547_), .B(men_men_n366_), .Y(men_men_n933_));
  NO2        u911(.A(men_men_n933_), .B(men_men_n691_), .Y(men_men_n934_));
  NA2        u912(.A(men_men_n966_), .B(men_men_n70_), .Y(men_men_n935_));
  NA2        u913(.A(men_men_n891_), .B(men_men_n813_), .Y(men_men_n936_));
  AOI210     u914(.A0(men_men_n936_), .A1(men_men_n935_), .B0(men_men_n626_), .Y(men_men_n937_));
  NA2        u915(.A(i_1_), .B(men_men_n70_), .Y(men_men_n938_));
  NO2        u916(.A(men_men_n938_), .B(men_men_n235_), .Y(men_men_n939_));
  NA3        u917(.A(men_men_n91_), .B(men_men_n297_), .C(men_men_n31_), .Y(men_men_n940_));
  INV        u918(.A(men_men_n940_), .Y(men_men_n941_));
  NO3        u919(.A(men_men_n941_), .B(men_men_n939_), .C(men_men_n937_), .Y(men_men_n942_));
  OAI210     u920(.A0(men_men_n260_), .A1(men_men_n155_), .B0(men_men_n82_), .Y(men_men_n943_));
  NA3        u921(.A(men_men_n694_), .B(men_men_n281_), .C(men_men_n74_), .Y(men_men_n944_));
  AOI210     u922(.A0(men_men_n944_), .A1(men_men_n943_), .B0(i_11_), .Y(men_men_n945_));
  NA2        u923(.A(men_men_n588_), .B(men_men_n215_), .Y(men_men_n946_));
  OAI210     u924(.A0(men_men_n946_), .A1(men_men_n825_), .B0(men_men_n205_), .Y(men_men_n947_));
  NA2        u925(.A(men_men_n161_), .B(i_5_), .Y(men_men_n948_));
  NO2        u926(.A(men_men_n947_), .B(men_men_n948_), .Y(men_men_n949_));
  NO3        u927(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n950_));
  NA2        u928(.A(men_men_n297_), .B(men_men_n950_), .Y(men_men_n951_));
  NO2        u929(.A(men_men_n951_), .B(men_men_n665_), .Y(men_men_n952_));
  NO3        u930(.A(men_men_n847_), .B(men_men_n464_), .C(men_men_n250_), .Y(men_men_n953_));
  NO2        u931(.A(men_men_n953_), .B(men_men_n544_), .Y(men_men_n954_));
  INV        u932(.A(men_men_n348_), .Y(men_men_n955_));
  AOI210     u933(.A0(men_men_n955_), .A1(men_men_n954_), .B0(men_men_n41_), .Y(men_men_n956_));
  NO4        u934(.A(men_men_n956_), .B(men_men_n952_), .C(men_men_n949_), .D(men_men_n945_), .Y(men_men_n957_));
  OAI210     u935(.A0(men_men_n942_), .A1(i_4_), .B0(men_men_n957_), .Y(men_men_n958_));
  NO3        u936(.A(men_men_n958_), .B(men_men_n934_), .C(men_men_n932_), .Y(men_men_n959_));
  NA4        u937(.A(men_men_n959_), .B(men_men_n918_), .C(men_men_n854_), .D(men_men_n787_), .Y(men4));
  INV        u938(.A(men_men_n646_), .Y(men_men_n963_));
  INV        u939(.A(i_2_), .Y(men_men_n964_));
  INV        u940(.A(men_men_n774_), .Y(men_men_n965_));
  INV        u941(.A(i_7_), .Y(men_men_n966_));
  INV        u942(.A(i_2_), .Y(men_men_n967_));
  INV        u943(.A(i_3_), .Y(men_men_n968_));
  INV        u944(.A(i_8_), .Y(men_men_n969_));
  INV        u945(.A(men_men_n140_), .Y(men_men_n970_));
  INV        u946(.A(men_men_n195_), .Y(men_men_n971_));
  INV        u947(.A(men_men_n588_), .Y(men_men_n972_));
  INV        u948(.A(i_12_), .Y(men_men_n973_));
  INV        u949(.A(i_10_), .Y(men_men_n974_));
  INV        u950(.A(i_1_), .Y(men_men_n975_));
  INV        u951(.A(men_men_n693_), .Y(men_men_n976_));
  INV        u952(.A(i_12_), .Y(men_men_n977_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule