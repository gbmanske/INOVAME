// Benchmark "top" written by ABC on Thu Jun 20 14:59:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n128_, new_new_n129_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n617_, new_new_n618_,
    new_new_n619_, new_new_n620_, new_new_n621_, new_new_n622_,
    new_new_n623_, new_new_n624_, new_new_n625_, new_new_n626_,
    new_new_n627_, new_new_n628_, new_new_n629_, new_new_n630_,
    new_new_n631_, new_new_n632_, new_new_n633_, new_new_n634_,
    new_new_n635_, new_new_n636_, new_new_n637_, new_new_n638_,
    new_new_n639_, new_new_n640_, new_new_n641_, new_new_n642_,
    new_new_n643_, new_new_n644_, new_new_n645_, new_new_n646_,
    new_new_n647_, new_new_n648_, new_new_n649_, new_new_n650_,
    new_new_n651_, new_new_n652_, new_new_n653_, new_new_n654_,
    new_new_n655_, new_new_n656_, new_new_n657_, new_new_n658_,
    new_new_n659_, new_new_n660_, new_new_n662_, new_new_n663_,
    new_new_n664_, new_new_n665_, new_new_n666_, new_new_n667_,
    new_new_n668_, new_new_n669_, new_new_n670_, new_new_n671_,
    new_new_n672_, new_new_n673_, new_new_n674_, new_new_n675_,
    new_new_n676_, new_new_n677_, new_new_n678_, new_new_n679_,
    new_new_n680_, new_new_n681_, new_new_n682_, new_new_n683_,
    new_new_n684_, new_new_n685_, new_new_n686_, new_new_n687_,
    new_new_n688_, new_new_n689_, new_new_n690_, new_new_n691_,
    new_new_n692_, new_new_n693_, new_new_n694_, new_new_n695_,
    new_new_n696_, new_new_n697_, new_new_n698_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n863_,
    new_new_n864_, new_new_n865_, new_new_n866_, new_new_n867_,
    new_new_n868_, new_new_n869_, new_new_n870_, new_new_n871_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(mai1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  NO2        g027(.A(new_new_n46_), .B(new_new_n45_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n50_), .B(new_new_n44_), .Y(new_new_n54_));
  NA3        g032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n55_));
  NO2        g033(.A(i_1_), .B(i_6_), .Y(new_new_n56_));
  NA2        g034(.A(i_8_), .B(i_7_), .Y(new_new_n57_));
  NO2        g035(.A(new_new_n57_), .B(new_new_n56_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_12_), .Y(new_new_n59_));
  NAi21      g037(.An(i_2_), .B(i_7_), .Y(new_new_n60_));
  INV        g038(.A(i_1_), .Y(new_new_n61_));
  NA3        g039(.A(i_1_), .B(new_new_n60_), .C(new_new_n31_), .Y(new_new_n62_));
  NA2        g040(.A(new_new_n62_), .B(new_new_n59_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n49_), .B(i_2_), .Y(new_new_n64_));
  NA2        g042(.A(i_1_), .B(i_6_), .Y(new_new_n65_));
  NO2        g043(.A(new_new_n65_), .B(new_new_n25_), .Y(new_new_n66_));
  INV        g044(.A(i_0_), .Y(new_new_n67_));
  NAi21      g045(.An(i_5_), .B(i_10_), .Y(new_new_n68_));
  NA2        g046(.A(i_5_), .B(i_9_), .Y(new_new_n69_));
  AOI210     g047(.A0(new_new_n69_), .A1(new_new_n68_), .B0(new_new_n67_), .Y(new_new_n70_));
  NO2        g048(.A(new_new_n70_), .B(new_new_n66_), .Y(new_new_n71_));
  NA2        g049(.A(new_new_n64_), .B(new_new_n71_), .Y(new_new_n72_));
  OAI210     g050(.A0(new_new_n72_), .A1(new_new_n63_), .B0(i_0_), .Y(new_new_n73_));
  NA2        g051(.A(i_12_), .B(i_5_), .Y(new_new_n74_));
  NO2        g052(.A(i_3_), .B(i_9_), .Y(new_new_n75_));
  NO2        g053(.A(i_3_), .B(i_7_), .Y(new_new_n76_));
  INV        g054(.A(i_6_), .Y(new_new_n77_));
  OR4        g055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n78_));
  INV        g056(.A(new_new_n78_), .Y(new_new_n79_));
  NO2        g057(.A(i_2_), .B(i_7_), .Y(new_new_n80_));
  NAi21      g058(.An(i_6_), .B(i_10_), .Y(new_new_n81_));
  NA2        g059(.A(i_6_), .B(i_9_), .Y(new_new_n82_));
  AOI210     g060(.A0(new_new_n82_), .A1(new_new_n81_), .B0(new_new_n61_), .Y(new_new_n83_));
  NA2        g061(.A(i_2_), .B(i_6_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n83_), .Y(new_new_n85_));
  NO2        g063(.A(new_new_n85_), .B(new_new_n74_), .Y(new_new_n86_));
  AN3        g064(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n87_));
  NAi21      g065(.An(i_6_), .B(i_11_), .Y(new_new_n88_));
  NO2        g066(.A(i_5_), .B(i_8_), .Y(new_new_n89_));
  NOi21      g067(.An(new_new_n89_), .B(new_new_n88_), .Y(new_new_n90_));
  AOI220     g068(.A0(new_new_n90_), .A1(new_new_n60_), .B0(new_new_n87_), .B1(new_new_n32_), .Y(new_new_n91_));
  INV        g069(.A(i_7_), .Y(new_new_n92_));
  NA2        g070(.A(new_new_n45_), .B(new_new_n92_), .Y(new_new_n93_));
  NO2        g071(.A(i_0_), .B(i_5_), .Y(new_new_n94_));
  NO2        g072(.A(new_new_n94_), .B(new_new_n77_), .Y(new_new_n95_));
  NA2        g073(.A(i_12_), .B(i_3_), .Y(new_new_n96_));
  INV        g074(.A(new_new_n96_), .Y(new_new_n97_));
  NA3        g075(.A(new_new_n97_), .B(new_new_n95_), .C(new_new_n93_), .Y(new_new_n98_));
  NAi21      g076(.An(i_7_), .B(i_11_), .Y(new_new_n99_));
  AN2        g077(.A(i_2_), .B(i_10_), .Y(new_new_n100_));
  NO2        g078(.A(new_new_n100_), .B(i_7_), .Y(new_new_n101_));
  OR2        g079(.A(new_new_n74_), .B(new_new_n56_), .Y(new_new_n102_));
  NO2        g080(.A(i_8_), .B(new_new_n92_), .Y(new_new_n103_));
  NO3        g081(.A(new_new_n103_), .B(new_new_n102_), .C(new_new_n101_), .Y(new_new_n104_));
  NA2        g082(.A(i_12_), .B(i_7_), .Y(new_new_n105_));
  NO2        g083(.A(new_new_n61_), .B(new_new_n26_), .Y(new_new_n106_));
  NA2        g084(.A(new_new_n106_), .B(i_0_), .Y(new_new_n107_));
  NA2        g085(.A(i_11_), .B(i_12_), .Y(new_new_n108_));
  OAI210     g086(.A0(new_new_n107_), .A1(new_new_n105_), .B0(new_new_n108_), .Y(new_new_n109_));
  NO2        g087(.A(new_new_n109_), .B(new_new_n104_), .Y(new_new_n110_));
  NA3        g088(.A(new_new_n110_), .B(new_new_n98_), .C(new_new_n91_), .Y(new_new_n111_));
  NOi21      g089(.An(i_1_), .B(i_5_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(i_11_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n92_), .B(new_new_n37_), .Y(new_new_n114_));
  NA2        g092(.A(i_7_), .B(new_new_n25_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n115_), .B(new_new_n114_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n116_), .B(new_new_n45_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n82_), .B(new_new_n81_), .Y(new_new_n118_));
  NAi21      g096(.An(i_3_), .B(i_8_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n60_), .Y(new_new_n120_));
  NO2        g098(.A(i_1_), .B(new_new_n77_), .Y(new_new_n121_));
  NO2        g099(.A(i_6_), .B(i_5_), .Y(new_new_n122_));
  NA2        g100(.A(new_new_n122_), .B(i_3_), .Y(new_new_n123_));
  AO210      g101(.A0(new_new_n123_), .A1(new_new_n46_), .B0(new_new_n121_), .Y(new_new_n124_));
  OAI220     g102(.A0(new_new_n124_), .A1(new_new_n99_), .B0(new_new_n120_), .B1(new_new_n113_), .Y(new_new_n125_));
  NO3        g103(.A(new_new_n125_), .B(new_new_n111_), .C(new_new_n86_), .Y(new_new_n126_));
  NA3        g104(.A(new_new_n126_), .B(new_new_n73_), .C(new_new_n54_), .Y(mai2));
  NO2        g105(.A(new_new_n61_), .B(new_new_n37_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n868_), .B(new_new_n128_), .Y(new_new_n129_));
  NA4        g107(.A(new_new_n129_), .B(new_new_n71_), .C(new_new_n64_), .D(new_new_n30_), .Y(mai0));
  AN2        g108(.A(i_8_), .B(i_7_), .Y(new_new_n131_));
  NA2        g109(.A(new_new_n131_), .B(i_6_), .Y(new_new_n132_));
  NO2        g110(.A(i_12_), .B(i_13_), .Y(new_new_n133_));
  NAi21      g111(.An(i_5_), .B(i_11_), .Y(new_new_n134_));
  NOi21      g112(.An(new_new_n133_), .B(new_new_n134_), .Y(new_new_n135_));
  NO2        g113(.A(i_0_), .B(i_1_), .Y(new_new_n136_));
  AN2        g114(.A(new_new_n133_), .B(new_new_n75_), .Y(new_new_n137_));
  NA2        g115(.A(i_1_), .B(i_5_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n67_), .B(new_new_n45_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(new_new_n36_), .Y(new_new_n140_));
  NO3        g118(.A(new_new_n140_), .B(new_new_n138_), .C(i_13_), .Y(new_new_n141_));
  OR2        g119(.A(i_0_), .B(i_1_), .Y(new_new_n142_));
  NO3        g120(.A(new_new_n142_), .B(new_new_n74_), .C(i_13_), .Y(new_new_n143_));
  NAi32      g121(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n144_));
  NAi21      g122(.An(new_new_n144_), .B(new_new_n143_), .Y(new_new_n145_));
  NOi21      g123(.An(i_4_), .B(i_10_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(new_new_n39_), .Y(new_new_n147_));
  NO2        g125(.A(i_3_), .B(i_5_), .Y(new_new_n148_));
  NA2        g126(.A(i_0_), .B(new_new_n148_), .Y(new_new_n149_));
  OAI210     g127(.A0(new_new_n149_), .A1(new_new_n147_), .B0(new_new_n145_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n150_), .B(new_new_n141_), .Y(new_new_n151_));
  NO2        g129(.A(new_new_n151_), .B(new_new_n132_), .Y(new_new_n152_));
  NOi21      g130(.An(i_4_), .B(i_9_), .Y(new_new_n153_));
  NOi21      g131(.An(i_11_), .B(i_13_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n154_), .B(new_new_n153_), .Y(new_new_n155_));
  NO2        g133(.A(i_4_), .B(i_5_), .Y(new_new_n156_));
  NAi21      g134(.An(i_12_), .B(i_11_), .Y(new_new_n157_));
  NO2        g135(.A(new_new_n157_), .B(i_13_), .Y(new_new_n158_));
  NO2        g136(.A(new_new_n67_), .B(new_new_n61_), .Y(new_new_n159_));
  NAi31      g137(.An(i_4_), .B(new_new_n137_), .C(i_11_), .Y(new_new_n160_));
  NA2        g138(.A(i_3_), .B(i_5_), .Y(new_new_n161_));
  BUFFER     g139(.A(new_new_n155_), .Y(new_new_n162_));
  AOI210     g140(.A0(new_new_n162_), .A1(new_new_n160_), .B0(new_new_n61_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n67_), .B(i_5_), .Y(new_new_n164_));
  NO2        g142(.A(i_13_), .B(i_10_), .Y(new_new_n165_));
  NA3        g143(.A(new_new_n165_), .B(new_new_n164_), .C(new_new_n43_), .Y(new_new_n166_));
  NO2        g144(.A(i_2_), .B(i_1_), .Y(new_new_n167_));
  NA2        g145(.A(new_new_n167_), .B(i_3_), .Y(new_new_n168_));
  NAi21      g146(.An(i_4_), .B(i_12_), .Y(new_new_n169_));
  NO4        g147(.A(new_new_n169_), .B(new_new_n168_), .C(new_new_n166_), .D(new_new_n25_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n170_), .B(new_new_n163_), .Y(new_new_n171_));
  INV        g149(.A(i_8_), .Y(new_new_n172_));
  NA2        g150(.A(i_8_), .B(i_6_), .Y(new_new_n173_));
  NO3        g151(.A(i_3_), .B(new_new_n77_), .C(new_new_n47_), .Y(new_new_n174_));
  NA2        g152(.A(new_new_n174_), .B(new_new_n103_), .Y(new_new_n175_));
  NO3        g153(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n176_));
  NA3        g154(.A(new_new_n176_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n177_));
  NO3        g155(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n178_));
  NA2        g156(.A(i_12_), .B(new_new_n178_), .Y(new_new_n179_));
  AOI210     g157(.A0(new_new_n179_), .A1(new_new_n177_), .B0(new_new_n175_), .Y(new_new_n180_));
  NO2        g158(.A(i_3_), .B(i_8_), .Y(new_new_n181_));
  NO3        g159(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n94_), .B(new_new_n56_), .Y(new_new_n183_));
  NO2        g161(.A(i_13_), .B(i_9_), .Y(new_new_n184_));
  NA2        g162(.A(new_new_n184_), .B(new_new_n172_), .Y(new_new_n185_));
  NAi21      g163(.An(i_12_), .B(i_3_), .Y(new_new_n186_));
  NO2        g164(.A(new_new_n43_), .B(i_5_), .Y(new_new_n187_));
  NO3        g165(.A(i_0_), .B(i_2_), .C(new_new_n61_), .Y(new_new_n188_));
  INV        g166(.A(new_new_n180_), .Y(new_new_n189_));
  OAI220     g167(.A0(new_new_n189_), .A1(i_4_), .B0(new_new_n173_), .B1(new_new_n171_), .Y(new_new_n190_));
  NAi21      g168(.An(i_12_), .B(i_7_), .Y(new_new_n191_));
  NA3        g169(.A(i_13_), .B(new_new_n172_), .C(i_10_), .Y(new_new_n192_));
  NO2        g170(.A(new_new_n192_), .B(new_new_n191_), .Y(new_new_n193_));
  NA2        g171(.A(i_0_), .B(i_5_), .Y(new_new_n194_));
  OAI220     g172(.A0(new_new_n77_), .A1(new_new_n168_), .B0(new_new_n61_), .B1(new_new_n123_), .Y(new_new_n195_));
  NAi31      g173(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n36_), .B(i_13_), .Y(new_new_n197_));
  NO2        g175(.A(new_new_n45_), .B(new_new_n61_), .Y(new_new_n198_));
  NA2        g176(.A(new_new_n198_), .B(new_new_n197_), .Y(new_new_n199_));
  INV        g177(.A(i_13_), .Y(new_new_n200_));
  NO2        g178(.A(i_12_), .B(new_new_n200_), .Y(new_new_n201_));
  NA3        g179(.A(new_new_n201_), .B(new_new_n176_), .C(new_new_n174_), .Y(new_new_n202_));
  INV        g180(.A(new_new_n202_), .Y(new_new_n203_));
  AOI220     g181(.A0(new_new_n203_), .A1(new_new_n131_), .B0(new_new_n195_), .B1(new_new_n193_), .Y(new_new_n204_));
  NO2        g182(.A(i_12_), .B(new_new_n37_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n161_), .B(i_4_), .Y(new_new_n206_));
  NA2        g184(.A(new_new_n206_), .B(new_new_n205_), .Y(new_new_n207_));
  OR2        g185(.A(i_8_), .B(i_7_), .Y(new_new_n208_));
  NO2        g186(.A(new_new_n208_), .B(new_new_n77_), .Y(new_new_n209_));
  INV        g187(.A(i_12_), .Y(new_new_n210_));
  NO3        g188(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n211_));
  NA2        g189(.A(i_2_), .B(i_1_), .Y(new_new_n212_));
  NAi21      g190(.An(i_4_), .B(i_3_), .Y(new_new_n213_));
  NO2        g191(.A(i_0_), .B(i_6_), .Y(new_new_n214_));
  NOi41      g192(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n215_));
  NO2        g193(.A(i_11_), .B(new_new_n200_), .Y(new_new_n216_));
  NAi21      g194(.An(i_3_), .B(i_7_), .Y(new_new_n217_));
  NA2        g195(.A(new_new_n210_), .B(i_9_), .Y(new_new_n218_));
  OR2        g196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  NO2        g197(.A(i_12_), .B(i_3_), .Y(new_new_n220_));
  NA2        g198(.A(i_3_), .B(i_9_), .Y(new_new_n221_));
  NAi21      g199(.An(i_7_), .B(i_10_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n223_));
  INV        g201(.A(new_new_n219_), .Y(new_new_n224_));
  INV        g202(.A(new_new_n132_), .Y(new_new_n225_));
  NA2        g203(.A(new_new_n210_), .B(i_13_), .Y(new_new_n226_));
  NO2        g204(.A(new_new_n226_), .B(new_new_n69_), .Y(new_new_n227_));
  AOI220     g205(.A0(new_new_n227_), .A1(new_new_n225_), .B0(new_new_n224_), .B1(new_new_n216_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n208_), .B(new_new_n37_), .Y(new_new_n229_));
  NA2        g207(.A(i_12_), .B(i_6_), .Y(new_new_n230_));
  OR2        g208(.A(i_13_), .B(i_9_), .Y(new_new_n231_));
  NO3        g209(.A(new_new_n231_), .B(new_new_n230_), .C(new_new_n47_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n213_), .B(i_2_), .Y(new_new_n233_));
  NA3        g211(.A(new_new_n233_), .B(new_new_n232_), .C(new_new_n43_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n216_), .B(i_9_), .Y(new_new_n235_));
  OAI210     g213(.A0(new_new_n61_), .A1(new_new_n235_), .B0(new_new_n234_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n139_), .B(new_new_n61_), .Y(new_new_n237_));
  NO3        g215(.A(i_11_), .B(new_new_n200_), .C(new_new_n25_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n217_), .B(i_8_), .Y(new_new_n239_));
  NO2        g217(.A(i_6_), .B(new_new_n47_), .Y(new_new_n240_));
  NA2        g218(.A(new_new_n239_), .B(new_new_n238_), .Y(new_new_n241_));
  NA3        g219(.A(i_3_), .B(new_new_n229_), .C(new_new_n201_), .Y(new_new_n242_));
  AOI210     g220(.A0(new_new_n242_), .A1(new_new_n241_), .B0(new_new_n237_), .Y(new_new_n243_));
  AOI210     g221(.A0(new_new_n236_), .A1(new_new_n229_), .B0(new_new_n243_), .Y(new_new_n244_));
  NA3        g222(.A(new_new_n244_), .B(new_new_n228_), .C(new_new_n204_), .Y(new_new_n245_));
  NO3        g223(.A(i_12_), .B(new_new_n200_), .C(new_new_n37_), .Y(new_new_n246_));
  INV        g224(.A(new_new_n246_), .Y(new_new_n247_));
  NA2        g225(.A(i_8_), .B(new_new_n92_), .Y(new_new_n248_));
  NO2        g226(.A(i_3_), .B(new_new_n248_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n212_), .B(i_0_), .Y(new_new_n250_));
  AOI220     g228(.A0(new_new_n250_), .A1(i_8_), .B0(i_1_), .B1(new_new_n131_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n240_), .B(new_new_n26_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n252_), .B(new_new_n251_), .Y(new_new_n253_));
  NA2        g231(.A(i_0_), .B(i_1_), .Y(new_new_n254_));
  NO2        g232(.A(new_new_n254_), .B(i_2_), .Y(new_new_n255_));
  NO2        g233(.A(new_new_n57_), .B(i_6_), .Y(new_new_n256_));
  NA2        g234(.A(new_new_n256_), .B(new_new_n255_), .Y(new_new_n257_));
  OAI210     g235(.A0(new_new_n149_), .A1(new_new_n132_), .B0(new_new_n257_), .Y(new_new_n258_));
  NO3        g236(.A(new_new_n258_), .B(new_new_n253_), .C(new_new_n249_), .Y(new_new_n259_));
  NO2        g237(.A(i_3_), .B(i_10_), .Y(new_new_n260_));
  NA3        g238(.A(new_new_n260_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n261_));
  AN2        g239(.A(i_3_), .B(i_10_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n45_), .B(new_new_n26_), .Y(new_new_n263_));
  NO2        g241(.A(new_new_n259_), .B(new_new_n247_), .Y(new_new_n264_));
  NO4        g242(.A(new_new_n264_), .B(new_new_n245_), .C(new_new_n190_), .D(new_new_n152_), .Y(new_new_n265_));
  NO3        g243(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n266_));
  NO3        g244(.A(i_6_), .B(new_new_n172_), .C(i_7_), .Y(new_new_n267_));
  NO2        g245(.A(i_2_), .B(i_3_), .Y(new_new_n268_));
  INV        g246(.A(new_new_n194_), .Y(new_new_n269_));
  NA3        g247(.A(new_new_n209_), .B(new_new_n268_), .C(i_1_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n45_), .B(new_new_n270_), .Y(new_new_n271_));
  NA2        g249(.A(new_new_n271_), .B(i_4_), .Y(new_new_n272_));
  NO2        g250(.A(i_12_), .B(i_10_), .Y(new_new_n273_));
  NOi21      g251(.An(i_5_), .B(i_0_), .Y(new_new_n274_));
  NA4        g252(.A(new_new_n76_), .B(new_new_n36_), .C(new_new_n77_), .D(i_8_), .Y(new_new_n275_));
  NO2        g253(.A(i_6_), .B(i_8_), .Y(new_new_n276_));
  AN2        g254(.A(i_0_), .B(new_new_n276_), .Y(new_new_n277_));
  NO2        g255(.A(i_1_), .B(i_7_), .Y(new_new_n278_));
  NA2        g256(.A(new_new_n277_), .B(i_4_), .Y(new_new_n279_));
  NA2        g257(.A(new_new_n279_), .B(new_new_n272_), .Y(new_new_n280_));
  NO2        g258(.A(i_8_), .B(new_new_n269_), .Y(new_new_n281_));
  OAI210     g259(.A0(new_new_n25_), .A1(new_new_n281_), .B0(i_3_), .Y(new_new_n282_));
  NO2        g260(.A(new_new_n84_), .B(new_new_n172_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n172_), .B(i_9_), .Y(new_new_n284_));
  NO3        g262(.A(new_new_n284_), .B(new_new_n283_), .C(new_new_n253_), .Y(new_new_n285_));
  AOI210     g263(.A0(new_new_n285_), .A1(new_new_n282_), .B0(new_new_n147_), .Y(new_new_n286_));
  AOI210     g264(.A0(new_new_n280_), .A1(new_new_n266_), .B0(new_new_n286_), .Y(new_new_n287_));
  NOi32      g265(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n288_));
  INV        g266(.A(new_new_n288_), .Y(new_new_n289_));
  NAi21      g267(.An(i_1_), .B(i_5_), .Y(new_new_n290_));
  NA2        g268(.A(new_new_n290_), .B(i_0_), .Y(new_new_n291_));
  NA2        g269(.A(new_new_n291_), .B(new_new_n25_), .Y(new_new_n292_));
  NO2        g270(.A(new_new_n292_), .B(new_new_n144_), .Y(new_new_n293_));
  NO2        g271(.A(new_new_n196_), .B(new_new_n144_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n144_), .B(new_new_n142_), .Y(new_new_n295_));
  NOi32      g273(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n296_));
  NA2        g274(.A(new_new_n296_), .B(new_new_n45_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n297_), .B(i_0_), .Y(new_new_n298_));
  OR3        g276(.A(new_new_n298_), .B(new_new_n295_), .C(new_new_n294_), .Y(new_new_n299_));
  NO2        g277(.A(i_1_), .B(new_new_n92_), .Y(new_new_n300_));
  NAi21      g278(.An(i_3_), .B(i_4_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(i_9_), .Y(new_new_n302_));
  NA2        g280(.A(i_7_), .B(new_new_n302_), .Y(new_new_n303_));
  NA2        g281(.A(i_2_), .B(i_7_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n301_), .B(i_10_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n305_), .B(new_new_n304_), .C(new_new_n214_), .Y(new_new_n306_));
  AOI210     g284(.A0(new_new_n306_), .A1(new_new_n303_), .B0(new_new_n164_), .Y(new_new_n307_));
  AOI210     g285(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n308_));
  OAI210     g286(.A0(new_new_n308_), .A1(new_new_n167_), .B0(new_new_n305_), .Y(new_new_n309_));
  AOI220     g287(.A0(new_new_n305_), .A1(new_new_n278_), .B0(new_new_n211_), .B1(new_new_n167_), .Y(new_new_n310_));
  AOI210     g288(.A0(new_new_n310_), .A1(new_new_n309_), .B0(i_5_), .Y(new_new_n311_));
  NO4        g289(.A(new_new_n311_), .B(new_new_n307_), .C(new_new_n299_), .D(new_new_n293_), .Y(new_new_n312_));
  NO2        g290(.A(new_new_n312_), .B(new_new_n289_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n57_), .B(new_new_n25_), .Y(new_new_n314_));
  AN2        g292(.A(i_12_), .B(i_5_), .Y(new_new_n315_));
  NO2        g293(.A(i_4_), .B(new_new_n26_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n315_), .Y(new_new_n317_));
  NO2        g295(.A(i_11_), .B(i_6_), .Y(new_new_n318_));
  NA3        g296(.A(new_new_n318_), .B(i_2_), .C(new_new_n200_), .Y(new_new_n319_));
  NO2        g297(.A(new_new_n319_), .B(new_new_n317_), .Y(new_new_n320_));
  NO2        g298(.A(new_new_n213_), .B(i_5_), .Y(new_new_n321_));
  NO2        g299(.A(i_5_), .B(i_10_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n133_), .B(new_new_n44_), .Y(new_new_n323_));
  NO2        g301(.A(new_new_n323_), .B(new_new_n213_), .Y(new_new_n324_));
  NA2        g302(.A(new_new_n324_), .B(new_new_n314_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n326_));
  INV        g304(.A(new_new_n320_), .Y(new_new_n327_));
  NO2        g305(.A(i_11_), .B(i_12_), .Y(new_new_n328_));
  NA2        g306(.A(new_new_n322_), .B(new_new_n210_), .Y(new_new_n329_));
  NO2        g307(.A(new_new_n92_), .B(new_new_n196_), .Y(new_new_n330_));
  NO2        g308(.A(i_13_), .B(new_new_n212_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n330_), .B(new_new_n331_), .Y(new_new_n332_));
  NA3        g310(.A(new_new_n332_), .B(new_new_n327_), .C(new_new_n325_), .Y(new_new_n333_));
  NO2        g311(.A(i_0_), .B(i_11_), .Y(new_new_n334_));
  NOi21      g312(.An(i_2_), .B(i_12_), .Y(new_new_n335_));
  NA2        g313(.A(new_new_n131_), .B(i_9_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n336_), .B(i_4_), .Y(new_new_n337_));
  NA2        g315(.A(new_new_n335_), .B(new_new_n337_), .Y(new_new_n338_));
  NAi21      g316(.An(i_9_), .B(i_4_), .Y(new_new_n339_));
  OR2        g317(.A(i_13_), .B(i_10_), .Y(new_new_n340_));
  NO2        g318(.A(new_new_n155_), .B(new_new_n114_), .Y(new_new_n341_));
  BUFFER     g319(.A(new_new_n192_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n92_), .B(new_new_n25_), .Y(new_new_n343_));
  NA2        g321(.A(new_new_n246_), .B(new_new_n343_), .Y(new_new_n344_));
  NA2        g322(.A(new_new_n240_), .B(new_new_n188_), .Y(new_new_n345_));
  OAI220     g323(.A0(new_new_n345_), .A1(new_new_n342_), .B0(new_new_n344_), .B1(new_new_n94_), .Y(new_new_n346_));
  INV        g324(.A(new_new_n346_), .Y(new_new_n347_));
  AOI210     g325(.A0(new_new_n347_), .A1(new_new_n338_), .B0(new_new_n26_), .Y(new_new_n348_));
  INV        g326(.A(new_new_n270_), .Y(new_new_n349_));
  AOI220     g327(.A0(new_new_n256_), .A1(i_2_), .B0(new_new_n250_), .B1(i_7_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n350_), .B(i_5_), .Y(new_new_n351_));
  AOI220     g329(.A0(i_3_), .A1(new_new_n255_), .B0(i_3_), .B1(new_new_n188_), .Y(new_new_n352_));
  NO2        g330(.A(new_new_n352_), .B(new_new_n248_), .Y(new_new_n353_));
  NO3        g331(.A(new_new_n353_), .B(new_new_n351_), .C(new_new_n349_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n174_), .B(new_new_n87_), .Y(new_new_n355_));
  NA3        g333(.A(i_2_), .B(new_new_n148_), .C(new_new_n77_), .Y(new_new_n356_));
  AOI210     g334(.A0(new_new_n356_), .A1(new_new_n355_), .B0(i_8_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n172_), .B(i_10_), .Y(new_new_n358_));
  NA2        g336(.A(i_1_), .B(i_2_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n256_), .B(i_2_), .Y(new_new_n360_));
  OAI220     g338(.A0(new_new_n360_), .A1(new_new_n161_), .B0(new_new_n359_), .B1(new_new_n358_), .Y(new_new_n361_));
  NA3        g339(.A(new_new_n278_), .B(new_new_n277_), .C(i_5_), .Y(new_new_n362_));
  INV        g340(.A(new_new_n267_), .Y(new_new_n363_));
  OAI210     g341(.A0(new_new_n363_), .A1(new_new_n168_), .B0(new_new_n362_), .Y(new_new_n364_));
  NO3        g342(.A(new_new_n364_), .B(new_new_n361_), .C(new_new_n357_), .Y(new_new_n365_));
  AOI210     g343(.A0(new_new_n365_), .A1(new_new_n354_), .B0(new_new_n235_), .Y(new_new_n366_));
  NO4        g344(.A(new_new_n366_), .B(new_new_n348_), .C(new_new_n333_), .D(new_new_n313_), .Y(new_new_n367_));
  NO2        g345(.A(new_new_n67_), .B(i_13_), .Y(new_new_n368_));
  NA3        g346(.A(new_new_n368_), .B(i_1_), .C(i_2_), .Y(new_new_n369_));
  NO2        g347(.A(i_10_), .B(i_9_), .Y(new_new_n370_));
  NAi21      g348(.An(i_12_), .B(i_8_), .Y(new_new_n371_));
  NO2        g349(.A(new_new_n371_), .B(i_3_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n372_), .B(new_new_n370_), .Y(new_new_n373_));
  NO2        g351(.A(new_new_n373_), .B(new_new_n369_), .Y(new_new_n374_));
  INV        g352(.A(new_new_n263_), .Y(new_new_n375_));
  NO3        g353(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n376_));
  NA2        g354(.A(new_new_n230_), .B(new_new_n88_), .Y(new_new_n377_));
  NA2        g355(.A(i_8_), .B(i_9_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n246_), .B(new_new_n183_), .Y(new_new_n379_));
  NO2        g357(.A(new_new_n379_), .B(new_new_n378_), .Y(new_new_n380_));
  NO3        g358(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n381_));
  NA3        g359(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n382_));
  NA4        g360(.A(new_new_n134_), .B(new_new_n106_), .C(new_new_n74_), .D(new_new_n23_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n382_), .Y(new_new_n384_));
  NO3        g362(.A(new_new_n384_), .B(new_new_n380_), .C(new_new_n374_), .Y(new_new_n385_));
  BUFFER     g363(.A(new_new_n257_), .Y(new_new_n386_));
  OA220      g364(.A0(new_new_n386_), .A1(new_new_n147_), .B0(new_new_n185_), .B1(new_new_n207_), .Y(new_new_n387_));
  NA2        g365(.A(new_new_n87_), .B(i_13_), .Y(new_new_n388_));
  NA2        g366(.A(i_3_), .B(new_new_n314_), .Y(new_new_n389_));
  NO2        g367(.A(i_2_), .B(i_13_), .Y(new_new_n390_));
  NA3        g368(.A(new_new_n390_), .B(new_new_n146_), .C(new_new_n90_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n389_), .B(new_new_n388_), .Y(new_new_n392_));
  NO3        g370(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n393_));
  NO2        g371(.A(i_6_), .B(i_7_), .Y(new_new_n394_));
  NOi21      g372(.An(i_2_), .B(i_7_), .Y(new_new_n395_));
  NAi31      g373(.An(i_11_), .B(new_new_n395_), .C(i_0_), .Y(new_new_n396_));
  NO2        g374(.A(new_new_n340_), .B(i_6_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n397_), .B(i_1_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n396_), .Y(new_new_n399_));
  NO2        g377(.A(i_3_), .B(new_new_n172_), .Y(new_new_n400_));
  NO2        g378(.A(i_6_), .B(i_10_), .Y(new_new_n401_));
  NA3        g379(.A(new_new_n215_), .B(new_new_n154_), .C(new_new_n122_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n45_), .B(new_new_n43_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n142_), .B(i_3_), .Y(new_new_n404_));
  NAi31      g382(.An(new_new_n403_), .B(new_new_n404_), .C(new_new_n201_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n405_), .B(new_new_n402_), .Y(new_new_n406_));
  NO3        g384(.A(new_new_n406_), .B(new_new_n399_), .C(new_new_n392_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n381_), .B(new_new_n322_), .Y(new_new_n408_));
  NO2        g386(.A(new_new_n408_), .B(new_new_n199_), .Y(new_new_n409_));
  NAi21      g387(.An(new_new_n192_), .B(new_new_n328_), .Y(new_new_n410_));
  NO2        g388(.A(new_new_n26_), .B(i_5_), .Y(new_new_n411_));
  NA3        g389(.A(i_6_), .B(new_new_n411_), .C(new_new_n131_), .Y(new_new_n412_));
  OAI220     g390(.A0(new_new_n38_), .A1(new_new_n412_), .B0(i_7_), .B1(new_new_n410_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n27_), .B(i_10_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n414_), .B(new_new_n388_), .Y(new_new_n415_));
  NO3        g393(.A(new_new_n415_), .B(new_new_n413_), .C(new_new_n409_), .Y(new_new_n416_));
  NA4        g394(.A(new_new_n416_), .B(new_new_n407_), .C(new_new_n387_), .D(new_new_n385_), .Y(new_new_n417_));
  NA3        g395(.A(new_new_n262_), .B(new_new_n158_), .C(new_new_n156_), .Y(new_new_n418_));
  NA2        g396(.A(new_new_n376_), .B(new_new_n263_), .Y(new_new_n419_));
  NA4        g397(.A(new_new_n368_), .B(i_1_), .C(new_new_n181_), .D(i_2_), .Y(new_new_n420_));
  INV        g398(.A(new_new_n420_), .Y(new_new_n421_));
  NA2        g399(.A(new_new_n315_), .B(new_new_n200_), .Y(new_new_n422_));
  NA2        g400(.A(new_new_n288_), .B(new_new_n67_), .Y(new_new_n423_));
  NA2        g401(.A(i_7_), .B(new_new_n296_), .Y(new_new_n424_));
  AO210      g402(.A0(new_new_n423_), .A1(new_new_n422_), .B0(new_new_n424_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n36_), .B(i_8_), .Y(new_new_n426_));
  INV        g404(.A(new_new_n425_), .Y(new_new_n427_));
  AOI210     g405(.A0(new_new_n421_), .A1(new_new_n182_), .B0(new_new_n427_), .Y(new_new_n428_));
  NO2        g406(.A(i_7_), .B(new_new_n177_), .Y(new_new_n429_));
  INV        g407(.A(new_new_n161_), .Y(new_new_n430_));
  AOI210     g408(.A0(new_new_n430_), .A1(new_new_n429_), .B0(new_new_n341_), .Y(new_new_n431_));
  NA4        g409(.A(new_new_n431_), .B(new_new_n428_), .C(new_new_n419_), .D(new_new_n418_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n321_), .B(new_new_n255_), .Y(new_new_n433_));
  NA2        g411(.A(new_new_n317_), .B(new_new_n433_), .Y(new_new_n434_));
  NO2        g412(.A(i_12_), .B(new_new_n172_), .Y(new_new_n435_));
  NOi31      g413(.An(new_new_n267_), .B(new_new_n340_), .C(new_new_n38_), .Y(new_new_n436_));
  OAI210     g414(.A0(new_new_n436_), .A1(new_new_n435_), .B0(new_new_n434_), .Y(new_new_n437_));
  NO2        g415(.A(i_8_), .B(i_7_), .Y(new_new_n438_));
  NA2        g416(.A(new_new_n43_), .B(i_10_), .Y(new_new_n439_));
  NO2        g417(.A(new_new_n439_), .B(i_6_), .Y(new_new_n440_));
  NA3        g418(.A(new_new_n440_), .B(new_new_n865_), .C(new_new_n438_), .Y(new_new_n441_));
  OAI220     g419(.A0(new_new_n161_), .A1(new_new_n226_), .B0(new_new_n388_), .B1(new_new_n123_), .Y(new_new_n442_));
  NA2        g420(.A(new_new_n442_), .B(new_new_n229_), .Y(new_new_n443_));
  NA3        g421(.A(new_new_n262_), .B(new_new_n156_), .C(new_new_n87_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n142_), .B(i_5_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n445_), .B(new_new_n268_), .Y(new_new_n446_));
  NA2        g424(.A(new_new_n446_), .B(new_new_n444_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n447_), .B(new_new_n381_), .Y(new_new_n448_));
  NA4        g426(.A(new_new_n448_), .B(new_new_n443_), .C(new_new_n441_), .D(new_new_n437_), .Y(new_new_n449_));
  NA2        g427(.A(new_new_n435_), .B(new_new_n238_), .Y(new_new_n450_));
  NO2        g428(.A(i_2_), .B(new_new_n450_), .Y(new_new_n451_));
  INV        g429(.A(new_new_n451_), .Y(new_new_n452_));
  NO3        g430(.A(new_new_n41_), .B(i_2_), .C(new_new_n47_), .Y(new_new_n453_));
  NO3        g431(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n208_), .B(new_new_n36_), .Y(new_new_n455_));
  AN2        g433(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n456_));
  OA210      g434(.A0(new_new_n456_), .A1(new_new_n453_), .B0(new_new_n288_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n340_), .B(i_1_), .Y(new_new_n458_));
  AN3        g436(.A(new_new_n458_), .B(new_new_n337_), .C(i_2_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n459_), .B(new_new_n457_), .Y(new_new_n460_));
  NO2        g438(.A(new_new_n77_), .B(new_new_n25_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n238_), .B(i_10_), .Y(new_new_n462_));
  NO2        g440(.A(new_new_n462_), .B(new_new_n375_), .Y(new_new_n463_));
  NO2        g441(.A(new_new_n105_), .B(new_new_n23_), .Y(new_new_n464_));
  INV        g442(.A(new_new_n267_), .Y(new_new_n465_));
  AOI220     g443(.A0(new_new_n465_), .A1(new_new_n360_), .B0(new_new_n162_), .B1(new_new_n160_), .Y(new_new_n466_));
  NOi21      g444(.An(new_new_n135_), .B(new_new_n275_), .Y(new_new_n467_));
  NO3        g445(.A(new_new_n467_), .B(new_new_n466_), .C(new_new_n463_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n423_), .B(new_new_n310_), .Y(new_new_n469_));
  INV        g447(.A(new_new_n268_), .Y(new_new_n470_));
  NO2        g448(.A(i_12_), .B(new_new_n77_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n471_), .B(new_new_n238_), .Y(new_new_n472_));
  NA2        g450(.A(new_new_n318_), .B(new_new_n246_), .Y(new_new_n473_));
  AOI210     g451(.A0(new_new_n473_), .A1(new_new_n472_), .B0(new_new_n470_), .Y(new_new_n474_));
  NO3        g452(.A(i_4_), .B(i_8_), .C(new_new_n261_), .Y(new_new_n475_));
  OR2        g453(.A(i_2_), .B(i_5_), .Y(new_new_n476_));
  NO2        g454(.A(i_2_), .B(new_new_n410_), .Y(new_new_n477_));
  NO4        g455(.A(new_new_n477_), .B(new_new_n475_), .C(new_new_n474_), .D(new_new_n469_), .Y(new_new_n478_));
  NA4        g456(.A(new_new_n478_), .B(new_new_n468_), .C(new_new_n460_), .D(new_new_n452_), .Y(new_new_n479_));
  NO4        g457(.A(new_new_n479_), .B(new_new_n449_), .C(new_new_n432_), .D(new_new_n417_), .Y(new_new_n480_));
  NA4        g458(.A(new_new_n480_), .B(new_new_n367_), .C(new_new_n287_), .D(new_new_n265_), .Y(mai7));
  NO2        g459(.A(new_new_n99_), .B(new_new_n81_), .Y(new_new_n482_));
  NA2        g460(.A(new_new_n401_), .B(new_new_n76_), .Y(new_new_n483_));
  NA2        g461(.A(i_11_), .B(new_new_n172_), .Y(new_new_n484_));
  NA3        g462(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n485_));
  NO2        g463(.A(new_new_n210_), .B(i_4_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n486_), .B(i_8_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n487_), .A1(new_new_n96_), .B0(new_new_n485_), .Y(new_new_n488_));
  OAI210     g466(.A0(new_new_n80_), .A1(new_new_n181_), .B0(new_new_n182_), .Y(new_new_n489_));
  NA2        g467(.A(i_4_), .B(i_8_), .Y(new_new_n490_));
  NO2        g468(.A(new_new_n489_), .B(i_13_), .Y(new_new_n491_));
  NO3        g469(.A(new_new_n491_), .B(new_new_n488_), .C(new_new_n482_), .Y(new_new_n492_));
  AOI210     g470(.A0(new_new_n119_), .A1(new_new_n60_), .B0(i_10_), .Y(new_new_n493_));
  AOI210     g471(.A0(new_new_n493_), .A1(new_new_n210_), .B0(new_new_n146_), .Y(new_new_n494_));
  OR2        g472(.A(i_6_), .B(i_10_), .Y(new_new_n495_));
  NO2        g473(.A(new_new_n495_), .B(new_new_n23_), .Y(new_new_n496_));
  OR3        g474(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n497_));
  NO3        g475(.A(new_new_n497_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n498_));
  INV        g476(.A(new_new_n178_), .Y(new_new_n499_));
  NO2        g477(.A(new_new_n498_), .B(new_new_n496_), .Y(new_new_n500_));
  OA220      g478(.A0(new_new_n500_), .A1(new_new_n470_), .B0(new_new_n494_), .B1(new_new_n231_), .Y(new_new_n501_));
  AOI210     g479(.A0(new_new_n501_), .A1(new_new_n492_), .B0(new_new_n61_), .Y(new_new_n502_));
  NOi21      g480(.An(i_11_), .B(i_7_), .Y(new_new_n503_));
  AO210      g481(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n504_));
  NO2        g482(.A(new_new_n504_), .B(new_new_n503_), .Y(new_new_n505_));
  NA2        g483(.A(new_new_n505_), .B(new_new_n184_), .Y(new_new_n506_));
  NA3        g484(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n507_));
  NAi21      g485(.An(new_new_n507_), .B(i_11_), .Y(new_new_n508_));
  AOI210     g486(.A0(new_new_n508_), .A1(new_new_n506_), .B0(new_new_n61_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n79_), .B(new_new_n61_), .Y(new_new_n510_));
  AO210      g488(.A0(new_new_n510_), .A1(new_new_n310_), .B0(new_new_n40_), .Y(new_new_n511_));
  NO3        g489(.A(new_new_n222_), .B(new_new_n186_), .C(new_new_n484_), .Y(new_new_n512_));
  OAI210     g490(.A0(new_new_n512_), .A1(new_new_n201_), .B0(new_new_n61_), .Y(new_new_n513_));
  NA2        g491(.A(new_new_n335_), .B(new_new_n31_), .Y(new_new_n514_));
  OR2        g492(.A(new_new_n186_), .B(new_new_n99_), .Y(new_new_n515_));
  NA2        g493(.A(new_new_n515_), .B(new_new_n514_), .Y(new_new_n516_));
  NO2        g494(.A(new_new_n61_), .B(i_9_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n517_), .B(i_4_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n518_), .B(new_new_n516_), .Y(new_new_n519_));
  NO2        g497(.A(i_1_), .B(i_12_), .Y(new_new_n520_));
  NA3        g498(.A(new_new_n519_), .B(new_new_n513_), .C(new_new_n511_), .Y(new_new_n521_));
  OAI210     g499(.A0(new_new_n521_), .A1(new_new_n509_), .B0(i_6_), .Y(new_new_n522_));
  NO2        g500(.A(new_new_n507_), .B(new_new_n99_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n523_), .B(new_new_n471_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n210_), .B(new_new_n77_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n525_), .B(i_11_), .Y(new_new_n526_));
  INV        g504(.A(new_new_n524_), .Y(new_new_n527_));
  NO3        g505(.A(new_new_n191_), .B(i_13_), .C(new_new_n77_), .Y(new_new_n528_));
  NA2        g506(.A(new_new_n528_), .B(new_new_n517_), .Y(new_new_n529_));
  NO3        g507(.A(new_new_n495_), .B(new_new_n208_), .C(new_new_n23_), .Y(new_new_n530_));
  AOI210     g508(.A0(i_1_), .A1(new_new_n223_), .B0(new_new_n530_), .Y(new_new_n531_));
  OAI210     g509(.A0(new_new_n531_), .A1(new_new_n43_), .B0(new_new_n529_), .Y(new_new_n532_));
  NA3        g510(.A(new_new_n438_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n533_));
  INV        g511(.A(i_2_), .Y(new_new_n534_));
  NA2        g512(.A(new_new_n128_), .B(i_9_), .Y(new_new_n535_));
  NA3        g513(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n536_));
  NO2        g514(.A(new_new_n45_), .B(i_1_), .Y(new_new_n537_));
  NA3        g515(.A(new_new_n537_), .B(new_new_n230_), .C(new_new_n43_), .Y(new_new_n538_));
  OAI220     g516(.A0(new_new_n538_), .A1(new_new_n536_), .B0(new_new_n535_), .B1(new_new_n534_), .Y(new_new_n539_));
  NA3        g517(.A(new_new_n517_), .B(new_new_n268_), .C(i_6_), .Y(new_new_n540_));
  NO2        g518(.A(new_new_n540_), .B(new_new_n23_), .Y(new_new_n541_));
  NO2        g519(.A(i_11_), .B(new_new_n37_), .Y(new_new_n542_));
  OR2        g520(.A(new_new_n541_), .B(new_new_n539_), .Y(new_new_n543_));
  NO3        g521(.A(new_new_n543_), .B(new_new_n532_), .C(new_new_n527_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n210_), .B(new_new_n92_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n545_), .B(new_new_n503_), .Y(new_new_n546_));
  NA2        g524(.A(new_new_n546_), .B(i_1_), .Y(new_new_n547_));
  NO2        g525(.A(new_new_n547_), .B(new_new_n497_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n339_), .B(new_new_n77_), .Y(new_new_n549_));
  NA2        g527(.A(new_new_n548_), .B(new_new_n45_), .Y(new_new_n550_));
  NA2        g528(.A(i_3_), .B(new_new_n172_), .Y(new_new_n551_));
  NO2        g529(.A(new_new_n551_), .B(new_new_n105_), .Y(new_new_n552_));
  AN2        g530(.A(new_new_n552_), .B(new_new_n440_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n77_), .B(i_9_), .Y(new_new_n554_));
  NA2        g532(.A(i_1_), .B(i_3_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n378_), .B(new_new_n84_), .Y(new_new_n556_));
  INV        g534(.A(new_new_n556_), .Y(new_new_n557_));
  NO2        g535(.A(new_new_n557_), .B(new_new_n555_), .Y(new_new_n558_));
  NO2        g536(.A(new_new_n558_), .B(new_new_n553_), .Y(new_new_n559_));
  NA4        g537(.A(new_new_n559_), .B(new_new_n550_), .C(new_new_n544_), .D(new_new_n522_), .Y(new_new_n560_));
  NO3        g538(.A(i_11_), .B(i_3_), .C(i_7_), .Y(new_new_n561_));
  NOi21      g539(.An(new_new_n561_), .B(i_10_), .Y(new_new_n562_));
  OA210      g540(.A0(new_new_n562_), .A1(new_new_n215_), .B0(new_new_n77_), .Y(new_new_n563_));
  NA2        g541(.A(i_7_), .B(new_new_n302_), .Y(new_new_n564_));
  NA3        g542(.A(new_new_n401_), .B(new_new_n426_), .C(new_new_n45_), .Y(new_new_n565_));
  NO2        g543(.A(new_new_n490_), .B(new_new_n77_), .Y(new_new_n566_));
  NA2        g544(.A(new_new_n566_), .B(new_new_n25_), .Y(new_new_n567_));
  NA2        g545(.A(new_new_n567_), .B(new_new_n565_), .Y(new_new_n568_));
  OAI210     g546(.A0(new_new_n568_), .A1(new_new_n563_), .B0(i_1_), .Y(new_new_n569_));
  AOI210     g547(.A0(new_new_n230_), .A1(new_new_n88_), .B0(i_1_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n301_), .B(i_2_), .Y(new_new_n571_));
  NA2        g549(.A(new_new_n571_), .B(new_new_n570_), .Y(new_new_n572_));
  OAI210     g550(.A0(new_new_n540_), .A1(new_new_n371_), .B0(new_new_n572_), .Y(new_new_n573_));
  INV        g551(.A(new_new_n573_), .Y(new_new_n574_));
  AOI210     g552(.A0(new_new_n574_), .A1(new_new_n569_), .B0(i_13_), .Y(new_new_n575_));
  NA2        g553(.A(new_new_n97_), .B(new_new_n128_), .Y(new_new_n576_));
  AOI220     g554(.A0(new_new_n390_), .A1(new_new_n146_), .B0(i_2_), .B1(new_new_n128_), .Y(new_new_n577_));
  OAI210     g555(.A0(new_new_n577_), .A1(new_new_n43_), .B0(new_new_n576_), .Y(new_new_n578_));
  AOI220     g556(.A0(i_7_), .A1(new_new_n549_), .B0(new_new_n215_), .B1(new_new_n121_), .Y(new_new_n579_));
  NO2        g557(.A(new_new_n579_), .B(new_new_n40_), .Y(new_new_n580_));
  AOI210     g558(.A0(new_new_n578_), .A1(new_new_n276_), .B0(new_new_n580_), .Y(new_new_n581_));
  NA2        g559(.A(new_new_n318_), .B(new_new_n537_), .Y(new_new_n582_));
  NO2        g560(.A(new_new_n582_), .B(new_new_n213_), .Y(new_new_n583_));
  AOI210     g561(.A0(new_new_n371_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n584_));
  NOi31      g562(.An(new_new_n584_), .B(new_new_n483_), .C(new_new_n43_), .Y(new_new_n585_));
  NA2        g563(.A(new_new_n118_), .B(i_13_), .Y(new_new_n586_));
  NO2        g564(.A(new_new_n536_), .B(new_new_n105_), .Y(new_new_n587_));
  INV        g565(.A(new_new_n587_), .Y(new_new_n588_));
  OAI220     g566(.A0(new_new_n588_), .A1(new_new_n65_), .B0(new_new_n586_), .B1(new_new_n570_), .Y(new_new_n589_));
  NA2        g567(.A(i_3_), .B(i_7_), .Y(new_new_n590_));
  NO3        g568(.A(new_new_n395_), .B(new_new_n210_), .C(new_new_n77_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n590_), .Y(new_new_n592_));
  AOI220     g570(.A0(new_new_n318_), .A1(new_new_n537_), .B0(new_new_n83_), .B1(new_new_n93_), .Y(new_new_n593_));
  OAI220     g571(.A0(new_new_n593_), .A1(new_new_n487_), .B0(new_new_n592_), .B1(new_new_n499_), .Y(new_new_n594_));
  NO4        g572(.A(new_new_n594_), .B(new_new_n589_), .C(new_new_n585_), .D(new_new_n583_), .Y(new_new_n595_));
  OR2        g573(.A(i_11_), .B(i_6_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n486_), .B(i_7_), .Y(new_new_n597_));
  AOI210     g575(.A0(new_new_n597_), .A1(new_new_n588_), .B0(new_new_n596_), .Y(new_new_n598_));
  NA3        g576(.A(new_new_n335_), .B(i_10_), .C(new_new_n88_), .Y(new_new_n599_));
  NA2        g577(.A(new_new_n526_), .B(i_13_), .Y(new_new_n600_));
  NAi21      g578(.An(i_11_), .B(i_12_), .Y(new_new_n601_));
  NOi41      g579(.An(new_new_n101_), .B(new_new_n601_), .C(i_13_), .D(new_new_n77_), .Y(new_new_n602_));
  NO2        g580(.A(new_new_n471_), .B(new_new_n490_), .Y(new_new_n603_));
  AOI210     g581(.A0(new_new_n603_), .A1(new_new_n266_), .B0(new_new_n602_), .Y(new_new_n604_));
  NA3        g582(.A(new_new_n604_), .B(new_new_n600_), .C(new_new_n599_), .Y(new_new_n605_));
  OAI210     g583(.A0(new_new_n605_), .A1(new_new_n598_), .B0(new_new_n61_), .Y(new_new_n606_));
  NO2        g584(.A(i_2_), .B(i_12_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n300_), .B(new_new_n607_), .Y(new_new_n608_));
  NO3        g586(.A(i_9_), .B(new_new_n316_), .C(new_new_n486_), .Y(new_new_n609_));
  NA2        g587(.A(new_new_n609_), .B(new_new_n300_), .Y(new_new_n610_));
  NO2        g588(.A(new_new_n119_), .B(i_2_), .Y(new_new_n611_));
  NA2        g589(.A(new_new_n611_), .B(new_new_n520_), .Y(new_new_n612_));
  NA3        g590(.A(new_new_n612_), .B(new_new_n610_), .C(new_new_n608_), .Y(new_new_n613_));
  NA3        g591(.A(new_new_n613_), .B(new_new_n44_), .C(new_new_n200_), .Y(new_new_n614_));
  NA4        g592(.A(new_new_n614_), .B(new_new_n606_), .C(new_new_n595_), .D(new_new_n581_), .Y(new_new_n615_));
  OR4        g593(.A(new_new_n615_), .B(new_new_n575_), .C(new_new_n560_), .D(new_new_n502_), .Y(mai5));
  AOI210     g594(.A0(new_new_n546_), .A1(new_new_n233_), .B0(new_new_n341_), .Y(new_new_n617_));
  AO210      g595(.A0(new_new_n24_), .A1(i_10_), .B0(new_new_n216_), .Y(new_new_n618_));
  NA3        g596(.A(new_new_n618_), .B(new_new_n607_), .C(new_new_n99_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n487_), .B(i_11_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n80_), .B(new_new_n620_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n621_), .B(new_new_n619_), .C(new_new_n617_), .Y(new_new_n622_));
  NO3        g600(.A(i_11_), .B(new_new_n210_), .C(i_13_), .Y(new_new_n623_));
  NO2        g601(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n624_));
  NA2        g602(.A(i_12_), .B(i_8_), .Y(new_new_n625_));
  OAI210     g603(.A0(new_new_n45_), .A1(i_3_), .B0(new_new_n625_), .Y(new_new_n626_));
  INV        g604(.A(new_new_n370_), .Y(new_new_n627_));
  AOI220     g605(.A0(new_new_n268_), .A1(new_new_n464_), .B0(new_new_n626_), .B1(new_new_n624_), .Y(new_new_n628_));
  INV        g606(.A(new_new_n628_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n622_), .Y(new_new_n630_));
  INV        g608(.A(new_new_n154_), .Y(new_new_n631_));
  INV        g609(.A(new_new_n215_), .Y(new_new_n632_));
  OAI210     g610(.A0(new_new_n571_), .A1(new_new_n372_), .B0(new_new_n101_), .Y(new_new_n633_));
  AOI210     g611(.A0(new_new_n633_), .A1(new_new_n632_), .B0(new_new_n631_), .Y(new_new_n634_));
  NO2        g612(.A(new_new_n378_), .B(new_new_n26_), .Y(new_new_n635_));
  NO2        g613(.A(new_new_n635_), .B(new_new_n343_), .Y(new_new_n636_));
  NA2        g614(.A(new_new_n636_), .B(i_2_), .Y(new_new_n637_));
  INV        g615(.A(new_new_n637_), .Y(new_new_n638_));
  AOI210     g616(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n340_), .Y(new_new_n639_));
  AOI210     g617(.A0(new_new_n639_), .A1(new_new_n638_), .B0(new_new_n634_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n169_), .B(new_new_n116_), .Y(new_new_n641_));
  NA2        g619(.A(new_new_n641_), .B(i_2_), .Y(new_new_n642_));
  INV        g620(.A(new_new_n155_), .Y(new_new_n643_));
  NO3        g621(.A(new_new_n504_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n644_));
  AOI210     g622(.A0(new_new_n643_), .A1(new_new_n80_), .B0(new_new_n644_), .Y(new_new_n645_));
  AOI210     g623(.A0(new_new_n645_), .A1(new_new_n642_), .B0(new_new_n172_), .Y(new_new_n646_));
  OA210      g624(.A0(new_new_n505_), .A1(new_new_n117_), .B0(i_13_), .Y(new_new_n647_));
  NA2        g625(.A(new_new_n178_), .B(new_new_n181_), .Y(new_new_n648_));
  INV        g626(.A(new_new_n137_), .Y(new_new_n649_));
  AOI210     g627(.A0(new_new_n649_), .A1(new_new_n648_), .B0(new_new_n304_), .Y(new_new_n650_));
  NA3        g628(.A(i_2_), .B(new_new_n262_), .C(new_new_n115_), .Y(new_new_n651_));
  INV        g629(.A(new_new_n651_), .Y(new_new_n652_));
  NO4        g630(.A(new_new_n652_), .B(new_new_n650_), .C(new_new_n647_), .D(new_new_n646_), .Y(new_new_n653_));
  NA2        g631(.A(new_new_n464_), .B(new_new_n28_), .Y(new_new_n654_));
  NA2        g632(.A(new_new_n623_), .B(new_new_n239_), .Y(new_new_n655_));
  NA2        g633(.A(new_new_n655_), .B(new_new_n654_), .Y(new_new_n656_));
  NO2        g634(.A(new_new_n60_), .B(i_12_), .Y(new_new_n657_));
  NO2        g635(.A(new_new_n657_), .B(new_new_n117_), .Y(new_new_n658_));
  NO2        g636(.A(new_new_n658_), .B(new_new_n484_), .Y(new_new_n659_));
  AOI220     g637(.A0(new_new_n659_), .A1(new_new_n36_), .B0(new_new_n656_), .B1(new_new_n45_), .Y(new_new_n660_));
  NA4        g638(.A(new_new_n660_), .B(new_new_n653_), .C(new_new_n640_), .D(new_new_n630_), .Y(mai6));
  NO2        g639(.A(i_9_), .B(new_new_n871_), .Y(new_new_n662_));
  OAI210     g640(.A0(new_new_n67_), .A1(new_new_n662_), .B0(new_new_n611_), .Y(new_new_n663_));
  NA4        g641(.A(new_new_n322_), .B(new_new_n400_), .C(new_new_n65_), .D(new_new_n92_), .Y(new_new_n664_));
  INV        g642(.A(new_new_n664_), .Y(new_new_n665_));
  NO2        g643(.A(new_new_n196_), .B(new_new_n403_), .Y(new_new_n666_));
  NO2        g644(.A(i_11_), .B(i_9_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n665_), .B(new_new_n274_), .Y(new_new_n668_));
  AO210      g646(.A0(new_new_n668_), .A1(new_new_n663_), .B0(i_12_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n305_), .B(new_new_n278_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n471_), .B(new_new_n61_), .Y(new_new_n671_));
  NA2        g649(.A(new_new_n562_), .B(new_new_n65_), .Y(new_new_n672_));
  NA4        g650(.A(new_new_n510_), .B(new_new_n672_), .C(new_new_n671_), .D(new_new_n670_), .Y(new_new_n673_));
  INV        g651(.A(new_new_n175_), .Y(new_new_n674_));
  AOI220     g652(.A0(new_new_n674_), .A1(new_new_n667_), .B0(new_new_n673_), .B1(new_new_n67_), .Y(new_new_n675_));
  NA2        g653(.A(new_new_n864_), .B(new_new_n657_), .Y(new_new_n676_));
  AOI210     g654(.A0(new_new_n676_), .A1(new_new_n424_), .B0(new_new_n164_), .Y(new_new_n677_));
  NO2        g655(.A(new_new_n32_), .B(i_11_), .Y(new_new_n678_));
  NA3        g656(.A(new_new_n678_), .B(new_new_n394_), .C(new_new_n322_), .Y(new_new_n679_));
  NA2        g657(.A(new_new_n455_), .B(new_new_n454_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n680_), .B(new_new_n679_), .Y(new_new_n681_));
  OR2        g659(.A(new_new_n681_), .B(new_new_n677_), .Y(new_new_n682_));
  NO2        g660(.A(i_11_), .B(i_2_), .Y(new_new_n683_));
  NA2        g661(.A(new_new_n47_), .B(new_new_n37_), .Y(new_new_n684_));
  NA2        g662(.A(new_new_n867_), .B(new_new_n683_), .Y(new_new_n685_));
  NA3        g663(.A(new_new_n284_), .B(new_new_n220_), .C(i_7_), .Y(new_new_n686_));
  OR2        g664(.A(new_new_n627_), .B(new_new_n36_), .Y(new_new_n687_));
  NA3        g665(.A(new_new_n687_), .B(new_new_n686_), .C(new_new_n685_), .Y(new_new_n688_));
  AOI220     g666(.A0(new_new_n866_), .A1(new_new_n454_), .B0(new_new_n666_), .B1(new_new_n590_), .Y(new_new_n689_));
  NA3        g667(.A(new_new_n304_), .B(new_new_n211_), .C(new_new_n136_), .Y(new_new_n690_));
  NA3        g668(.A(new_new_n690_), .B(new_new_n689_), .C(new_new_n489_), .Y(new_new_n691_));
  NA3        g669(.A(new_new_n426_), .B(new_new_n401_), .C(new_new_n194_), .Y(new_new_n692_));
  AOI210     g670(.A0(new_new_n372_), .A1(new_new_n370_), .B0(new_new_n453_), .Y(new_new_n693_));
  OAI210     g671(.A0(new_new_n870_), .A1(new_new_n102_), .B0(new_new_n334_), .Y(new_new_n694_));
  INV        g672(.A(new_new_n476_), .Y(new_new_n695_));
  NA3        g673(.A(new_new_n695_), .B(new_new_n273_), .C(i_7_), .Y(new_new_n696_));
  NA4        g674(.A(new_new_n696_), .B(new_new_n694_), .C(new_new_n693_), .D(new_new_n692_), .Y(new_new_n697_));
  NO4        g675(.A(new_new_n697_), .B(new_new_n691_), .C(new_new_n688_), .D(new_new_n682_), .Y(new_new_n698_));
  NA4        g676(.A(new_new_n698_), .B(new_new_n675_), .C(new_new_n669_), .D(new_new_n312_), .Y(mai3));
  NO2        g677(.A(i_11_), .B(new_new_n210_), .Y(new_new_n700_));
  NA2        g678(.A(new_new_n250_), .B(new_new_n700_), .Y(new_new_n701_));
  NO2        g679(.A(new_new_n701_), .B(new_new_n172_), .Y(new_new_n702_));
  AN2        g680(.A(new_new_n702_), .B(new_new_n156_), .Y(new_new_n703_));
  NA3        g681(.A(new_new_n690_), .B(new_new_n489_), .C(new_new_n303_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n704_), .B(new_new_n39_), .Y(new_new_n705_));
  NO3        g683(.A(new_new_n515_), .B(new_new_n378_), .C(new_new_n121_), .Y(new_new_n706_));
  NA2        g684(.A(new_new_n335_), .B(new_new_n44_), .Y(new_new_n707_));
  AN2        g685(.A(new_new_n377_), .B(new_new_n53_), .Y(new_new_n708_));
  NO2        g686(.A(new_new_n708_), .B(new_new_n706_), .Y(new_new_n709_));
  AOI210     g687(.A0(new_new_n709_), .A1(new_new_n705_), .B0(new_new_n47_), .Y(new_new_n710_));
  NOi21      g688(.An(i_5_), .B(i_9_), .Y(new_new_n711_));
  NA2        g689(.A(new_new_n711_), .B(new_new_n368_), .Y(new_new_n712_));
  NO3        g690(.A(new_new_n336_), .B(new_new_n230_), .C(new_new_n67_), .Y(new_new_n713_));
  INV        g691(.A(new_new_n713_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n714_), .B(i_4_), .Y(new_new_n715_));
  NO3        g693(.A(new_new_n715_), .B(new_new_n710_), .C(new_new_n703_), .Y(new_new_n716_));
  NA2        g694(.A(new_new_n266_), .B(new_new_n120_), .Y(new_new_n717_));
  NAi21      g695(.An(new_new_n147_), .B(i_5_), .Y(new_new_n718_));
  NO2        g696(.A(new_new_n717_), .B(new_new_n329_), .Y(new_new_n719_));
  INV        g697(.A(new_new_n719_), .Y(new_new_n720_));
  NA2        g698(.A(new_new_n461_), .B(i_0_), .Y(new_new_n721_));
  NO3        g699(.A(new_new_n721_), .B(new_new_n317_), .C(new_new_n80_), .Y(new_new_n722_));
  NO3        g700(.A(new_new_n476_), .B(new_new_n191_), .C(new_new_n340_), .Y(new_new_n723_));
  AOI210     g701(.A0(new_new_n723_), .A1(i_11_), .B0(new_new_n722_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n623_), .B(new_new_n274_), .Y(new_new_n725_));
  NO2        g703(.A(new_new_n401_), .B(new_new_n56_), .Y(new_new_n726_));
  NO2        g704(.A(new_new_n726_), .B(new_new_n725_), .Y(new_new_n727_));
  NO2        g705(.A(new_new_n218_), .B(new_new_n138_), .Y(new_new_n728_));
  INV        g706(.A(new_new_n439_), .Y(new_new_n729_));
  NO4        g707(.A(new_new_n105_), .B(new_new_n56_), .C(new_new_n551_), .D(i_5_), .Y(new_new_n730_));
  AO220      g708(.A0(new_new_n730_), .A1(new_new_n729_), .B0(new_new_n728_), .B1(i_6_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n167_), .B(new_new_n181_), .Y(new_new_n732_));
  NO2        g710(.A(new_new_n732_), .B(new_new_n725_), .Y(new_new_n733_));
  NO3        g711(.A(new_new_n733_), .B(new_new_n731_), .C(new_new_n727_), .Y(new_new_n734_));
  NA3        g712(.A(new_new_n734_), .B(new_new_n724_), .C(new_new_n720_), .Y(new_new_n735_));
  NA2        g713(.A(i_11_), .B(i_9_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n47_), .B(i_7_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n326_), .B(new_new_n159_), .Y(new_new_n738_));
  NAi31      g716(.An(new_new_n227_), .B(new_new_n738_), .C(new_new_n145_), .Y(new_new_n739_));
  NO2        g717(.A(new_new_n157_), .B(i_0_), .Y(new_new_n740_));
  NA2        g718(.A(new_new_n394_), .B(new_new_n206_), .Y(new_new_n741_));
  OAI220     g719(.A0(i_12_), .A1(new_new_n712_), .B0(new_new_n741_), .B1(new_new_n157_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n742_), .B(new_new_n739_), .Y(new_new_n743_));
  NA2        g721(.A(new_new_n542_), .B(new_new_n112_), .Y(new_new_n744_));
  NO2        g722(.A(i_6_), .B(new_new_n744_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n371_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n746_));
  NA2        g724(.A(new_new_n154_), .B(new_new_n94_), .Y(new_new_n747_));
  NOi32      g725(.An(new_new_n746_), .Bn(new_new_n167_), .C(new_new_n747_), .Y(new_new_n748_));
  NO2        g726(.A(new_new_n869_), .B(new_new_n707_), .Y(new_new_n749_));
  NO3        g727(.A(new_new_n749_), .B(new_new_n748_), .C(new_new_n745_), .Y(new_new_n750_));
  NOi21      g728(.An(i_7_), .B(i_5_), .Y(new_new_n751_));
  NOi31      g729(.An(new_new_n751_), .B(i_0_), .C(new_new_n601_), .Y(new_new_n752_));
  NA3        g730(.A(new_new_n752_), .B(new_new_n316_), .C(i_6_), .Y(new_new_n753_));
  BUFFER     g731(.A(new_new_n753_), .Y(new_new_n754_));
  NA3        g732(.A(new_new_n754_), .B(new_new_n750_), .C(new_new_n743_), .Y(new_new_n755_));
  OA210      g733(.A0(new_new_n394_), .A1(new_new_n198_), .B0(new_new_n393_), .Y(new_new_n756_));
  NA3        g734(.A(new_new_n393_), .B(new_new_n335_), .C(new_new_n44_), .Y(new_new_n757_));
  OAI210     g735(.A0(new_new_n718_), .A1(i_6_), .B0(new_new_n757_), .Y(new_new_n758_));
  INV        g736(.A(new_new_n166_), .Y(new_new_n759_));
  AOI220     g737(.A0(new_new_n759_), .A1(new_new_n394_), .B0(new_new_n758_), .B1(new_new_n67_), .Y(new_new_n760_));
  NA2        g738(.A(new_new_n314_), .B(new_new_n525_), .Y(new_new_n761_));
  NA2        g739(.A(new_new_n84_), .B(new_new_n43_), .Y(new_new_n762_));
  NO2        g740(.A(new_new_n69_), .B(new_new_n625_), .Y(new_new_n763_));
  NA2        g741(.A(new_new_n763_), .B(new_new_n762_), .Y(new_new_n764_));
  AOI210     g742(.A0(new_new_n764_), .A1(new_new_n761_), .B0(new_new_n46_), .Y(new_new_n765_));
  NO3        g743(.A(new_new_n476_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n766_));
  NO2        g744(.A(new_new_n445_), .B(new_new_n766_), .Y(new_new_n767_));
  NAi21      g745(.An(i_9_), .B(i_5_), .Y(new_new_n768_));
  NO2        g746(.A(new_new_n485_), .B(new_new_n96_), .Y(new_new_n769_));
  NA2        g747(.A(new_new_n769_), .B(i_0_), .Y(new_new_n770_));
  OAI220     g748(.A0(new_new_n770_), .A1(new_new_n77_), .B0(new_new_n767_), .B1(new_new_n155_), .Y(new_new_n771_));
  NO3        g749(.A(new_new_n771_), .B(new_new_n765_), .C(new_new_n427_), .Y(new_new_n772_));
  NA2        g750(.A(new_new_n772_), .B(new_new_n760_), .Y(new_new_n773_));
  NO3        g751(.A(new_new_n773_), .B(new_new_n755_), .C(new_new_n735_), .Y(new_new_n774_));
  NO2        g752(.A(i_0_), .B(new_new_n601_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n67_), .B(new_new_n43_), .Y(new_new_n776_));
  NO3        g754(.A(new_new_n96_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n777_));
  AO220      g755(.A0(new_new_n777_), .A1(new_new_n43_), .B0(new_new_n775_), .B1(new_new_n156_), .Y(new_new_n778_));
  AOI210     g756(.A0(new_new_n671_), .A1(new_new_n564_), .B0(new_new_n747_), .Y(new_new_n779_));
  AOI210     g757(.A0(new_new_n778_), .A1(new_new_n283_), .B0(new_new_n779_), .Y(new_new_n780_));
  NA3        g758(.A(new_new_n135_), .B(new_new_n554_), .C(new_new_n67_), .Y(new_new_n781_));
  NA3        g759(.A(i_6_), .B(i_2_), .C(new_new_n47_), .Y(new_new_n782_));
  NA2        g760(.A(new_new_n700_), .B(i_9_), .Y(new_new_n783_));
  AOI210     g761(.A0(new_new_n782_), .A1(new_new_n412_), .B0(new_new_n783_), .Y(new_new_n784_));
  NA2        g762(.A(new_new_n214_), .B(new_new_n205_), .Y(new_new_n785_));
  AOI210     g763(.A0(new_new_n785_), .A1(new_new_n721_), .B0(new_new_n138_), .Y(new_new_n786_));
  NO2        g764(.A(new_new_n786_), .B(new_new_n784_), .Y(new_new_n787_));
  NA3        g765(.A(new_new_n787_), .B(new_new_n781_), .C(new_new_n780_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n39_), .B(new_new_n28_), .C(new_new_n43_), .Y(new_new_n789_));
  NA2        g767(.A(new_new_n737_), .B(new_new_n404_), .Y(new_new_n790_));
  AOI210     g768(.A0(new_new_n789_), .A1(new_new_n147_), .B0(new_new_n790_), .Y(new_new_n791_));
  INV        g769(.A(new_new_n791_), .Y(new_new_n792_));
  NO3        g770(.A(new_new_n187_), .B(new_new_n315_), .C(i_0_), .Y(new_new_n793_));
  OAI210     g771(.A0(new_new_n793_), .A1(new_new_n70_), .B0(i_13_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n794_), .B(new_new_n792_), .Y(new_new_n795_));
  NO2        g773(.A(new_new_n213_), .B(new_new_n84_), .Y(new_new_n796_));
  NA2        g774(.A(new_new_n796_), .B(new_new_n775_), .Y(new_new_n797_));
  NA2        g775(.A(new_new_n751_), .B(new_new_n404_), .Y(new_new_n798_));
  INV        g776(.A(new_new_n158_), .Y(new_new_n799_));
  OA220      g777(.A0(new_new_n799_), .A1(new_new_n798_), .B0(new_new_n797_), .B1(i_5_), .Y(new_new_n800_));
  AOI210     g778(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n157_), .Y(new_new_n801_));
  NA2        g779(.A(new_new_n801_), .B(new_new_n756_), .Y(new_new_n802_));
  NA2        g780(.A(new_new_n402_), .B(new_new_n391_), .Y(new_new_n803_));
  INV        g781(.A(new_new_n803_), .Y(new_new_n804_));
  NA3        g782(.A(new_new_n322_), .B(new_new_n277_), .C(new_new_n197_), .Y(new_new_n805_));
  INV        g783(.A(new_new_n805_), .Y(new_new_n806_));
  NOi31      g784(.An(new_new_n321_), .B(new_new_n776_), .C(new_new_n212_), .Y(new_new_n807_));
  NO3        g785(.A(new_new_n736_), .B(new_new_n194_), .C(new_new_n169_), .Y(new_new_n808_));
  NO3        g786(.A(new_new_n808_), .B(new_new_n807_), .C(new_new_n806_), .Y(new_new_n809_));
  NA4        g787(.A(new_new_n809_), .B(new_new_n804_), .C(new_new_n802_), .D(new_new_n800_), .Y(new_new_n810_));
  NO2        g788(.A(new_new_n77_), .B(i_5_), .Y(new_new_n811_));
  NA3        g789(.A(new_new_n700_), .B(new_new_n100_), .C(new_new_n115_), .Y(new_new_n812_));
  INV        g790(.A(new_new_n812_), .Y(new_new_n813_));
  NA2        g791(.A(new_new_n813_), .B(new_new_n811_), .Y(new_new_n814_));
  NA2        g792(.A(new_new_n262_), .B(i_5_), .Y(new_new_n815_));
  NO4        g793(.A(new_new_n212_), .B(new_new_n187_), .C(i_0_), .D(i_12_), .Y(new_new_n816_));
  AOI220     g794(.A0(new_new_n816_), .A1(new_new_n863_), .B0(new_new_n665_), .B1(new_new_n158_), .Y(new_new_n817_));
  BUFFER     g795(.A(new_new_n138_), .Y(new_new_n818_));
  NO4        g796(.A(new_new_n818_), .B(i_12_), .C(new_new_n533_), .D(new_new_n121_), .Y(new_new_n819_));
  NA2        g797(.A(new_new_n819_), .B(new_new_n194_), .Y(new_new_n820_));
  NA2        g798(.A(new_new_n751_), .B(new_new_n390_), .Y(new_new_n821_));
  OAI220     g799(.A0(i_6_), .A1(new_new_n815_), .B0(new_new_n821_), .B1(i_1_), .Y(new_new_n822_));
  NA2        g800(.A(new_new_n822_), .B(new_new_n740_), .Y(new_new_n823_));
  NA4        g801(.A(new_new_n823_), .B(new_new_n820_), .C(new_new_n817_), .D(new_new_n814_), .Y(new_new_n824_));
  NO4        g802(.A(new_new_n824_), .B(new_new_n810_), .C(new_new_n795_), .D(new_new_n788_), .Y(new_new_n825_));
  OAI210     g803(.A0(new_new_n683_), .A1(new_new_n678_), .B0(new_new_n37_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n826_), .B(new_new_n494_), .Y(new_new_n827_));
  NA2        g805(.A(new_new_n827_), .B(new_new_n184_), .Y(new_new_n828_));
  NA2        g806(.A(new_new_n165_), .B(new_new_n167_), .Y(new_new_n829_));
  OAI210     g807(.A0(new_new_n498_), .A1(new_new_n496_), .B0(new_new_n268_), .Y(new_new_n830_));
  NA2        g808(.A(new_new_n830_), .B(new_new_n829_), .Y(new_new_n831_));
  NO2        g809(.A(new_new_n382_), .B(new_new_n230_), .Y(new_new_n832_));
  NO2        g810(.A(new_new_n832_), .B(new_new_n723_), .Y(new_new_n833_));
  INV        g811(.A(new_new_n833_), .Y(new_new_n834_));
  AOI210     g812(.A0(new_new_n831_), .A1(new_new_n47_), .B0(new_new_n834_), .Y(new_new_n835_));
  AOI210     g813(.A0(new_new_n835_), .A1(new_new_n828_), .B0(new_new_n67_), .Y(new_new_n836_));
  NO2        g814(.A(new_new_n456_), .B(new_new_n311_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n837_), .B(new_new_n631_), .Y(new_new_n838_));
  AOI210     g816(.A0(new_new_n801_), .A1(new_new_n737_), .B0(new_new_n752_), .Y(new_new_n839_));
  NO2        g817(.A(new_new_n839_), .B(new_new_n555_), .Y(new_new_n840_));
  INV        g818(.A(new_new_n55_), .Y(new_new_n841_));
  NA2        g819(.A(new_new_n841_), .B(new_new_n70_), .Y(new_new_n842_));
  NO2        g820(.A(new_new_n842_), .B(new_new_n210_), .Y(new_new_n843_));
  NO2        g821(.A(new_new_n843_), .B(new_new_n840_), .Y(new_new_n844_));
  OAI210     g822(.A0(new_new_n232_), .A1(new_new_n143_), .B0(new_new_n80_), .Y(new_new_n845_));
  NO2        g823(.A(new_new_n845_), .B(i_11_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n746_), .B(new_new_n184_), .Y(new_new_n847_));
  NA2        g825(.A(i_0_), .B(i_5_), .Y(new_new_n848_));
  AOI210     g826(.A0(new_new_n847_), .A1(new_new_n648_), .B0(new_new_n848_), .Y(new_new_n849_));
  NO3        g827(.A(new_new_n57_), .B(new_new_n56_), .C(i_4_), .Y(new_new_n850_));
  NA2        g828(.A(new_new_n871_), .B(new_new_n850_), .Y(new_new_n851_));
  NO2        g829(.A(new_new_n851_), .B(new_new_n601_), .Y(new_new_n852_));
  NO3        g830(.A(new_new_n768_), .B(i_11_), .C(new_new_n217_), .Y(new_new_n853_));
  NO2        g831(.A(new_new_n853_), .B(new_new_n453_), .Y(new_new_n854_));
  INV        g832(.A(new_new_n294_), .Y(new_new_n855_));
  AOI210     g833(.A0(new_new_n855_), .A1(new_new_n854_), .B0(new_new_n40_), .Y(new_new_n856_));
  NO4        g834(.A(new_new_n856_), .B(new_new_n852_), .C(new_new_n849_), .D(new_new_n846_), .Y(new_new_n857_));
  OAI210     g835(.A0(new_new_n844_), .A1(i_4_), .B0(new_new_n857_), .Y(new_new_n858_));
  NO3        g836(.A(new_new_n858_), .B(new_new_n838_), .C(new_new_n836_), .Y(new_new_n859_));
  NA4        g837(.A(new_new_n859_), .B(new_new_n825_), .C(new_new_n774_), .D(new_new_n716_), .Y(mai4));
  INV        g838(.A(new_new_n213_), .Y(new_new_n863_));
  INV        g839(.A(i_9_), .Y(new_new_n864_));
  INV        g840(.A(new_new_n213_), .Y(new_new_n865_));
  INV        g841(.A(i_11_), .Y(new_new_n866_));
  INV        g842(.A(new_new_n684_), .Y(new_new_n867_));
  INV        g843(.A(i_6_), .Y(new_new_n868_));
  INV        g844(.A(new_new_n274_), .Y(new_new_n869_));
  INV        g845(.A(new_new_n495_), .Y(new_new_n870_));
  INV        g846(.A(i_5_), .Y(new_new_n871_));
endmodule


