//Benchmark atmr_max1024_476_0.0156

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n62_), .B(ori_ori_n36_), .Y(ori_ori_n63_));
  NO2        o047(.A(x7), .B(x6), .Y(ori_ori_n64_));
  NO2        o048(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n65_));
  NO2        o049(.A(x8), .B(x2), .Y(ori_ori_n66_));
  INV        o050(.A(ori_ori_n66_), .Y(ori_ori_n67_));
  NO2        o051(.A(ori_ori_n67_), .B(x1), .Y(ori_ori_n68_));
  OA210      o052(.A0(ori_ori_n68_), .A1(ori_ori_n65_), .B0(ori_ori_n64_), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n70_));
  OAI210     o054(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  NO2        o055(.A(ori_ori_n71_), .B(ori_ori_n69_), .Y(ori_ori_n72_));
  NA2        o056(.A(ori_ori_n72_), .B(x4), .Y(ori_ori_n73_));
  NA2        o057(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n74_));
  OAI210     o058(.A0(ori_ori_n74_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n75_));
  NA2        o059(.A(x5), .B(x3), .Y(ori_ori_n76_));
  NO2        o060(.A(x8), .B(x6), .Y(ori_ori_n77_));
  NO4        o061(.A(ori_ori_n77_), .B(ori_ori_n76_), .C(ori_ori_n64_), .D(ori_ori_n54_), .Y(ori_ori_n78_));
  NAi21      o062(.An(x4), .B(x3), .Y(ori_ori_n79_));
  INV        o063(.A(ori_ori_n79_), .Y(ori_ori_n80_));
  NO2        o064(.A(ori_ori_n80_), .B(ori_ori_n22_), .Y(ori_ori_n81_));
  NO2        o065(.A(x4), .B(x2), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n82_), .B(x3), .Y(ori_ori_n83_));
  NO3        o067(.A(ori_ori_n83_), .B(ori_ori_n81_), .C(ori_ori_n18_), .Y(ori_ori_n84_));
  NO3        o068(.A(ori_ori_n84_), .B(ori_ori_n78_), .C(ori_ori_n75_), .Y(ori_ori_n85_));
  NA2        o069(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n86_));
  NO2        o070(.A(ori_ori_n86_), .B(ori_ori_n25_), .Y(ori_ori_n87_));
  INV        o071(.A(x8), .Y(ori_ori_n88_));
  NA2        o072(.A(x2), .B(x1), .Y(ori_ori_n89_));
  INV        o073(.A(ori_ori_n87_), .Y(ori_ori_n90_));
  NO2        o074(.A(ori_ori_n90_), .B(ori_ori_n26_), .Y(ori_ori_n91_));
  AOI210     o075(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n92_));
  OAI210     o076(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n93_));
  NO3        o077(.A(ori_ori_n93_), .B(ori_ori_n92_), .C(ori_ori_n91_), .Y(ori_ori_n94_));
  NA2        o078(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n95_));
  NO2        o079(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n96_));
  OAI210     o080(.A0(ori_ori_n96_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n97_));
  AOI210     o081(.A0(ori_ori_n95_), .A1(ori_ori_n52_), .B0(ori_ori_n97_), .Y(ori_ori_n98_));
  NO2        o082(.A(x3), .B(x2), .Y(ori_ori_n99_));
  NA3        o083(.A(ori_ori_n99_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n100_));
  AOI210     o084(.A0(x8), .A1(x6), .B0(ori_ori_n100_), .Y(ori_ori_n101_));
  NA2        o085(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n102_));
  OAI210     o086(.A0(ori_ori_n102_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n103_));
  NO4        o087(.A(ori_ori_n103_), .B(ori_ori_n101_), .C(ori_ori_n98_), .D(ori_ori_n94_), .Y(ori_ori_n104_));
  AO210      o088(.A0(ori_ori_n85_), .A1(ori_ori_n73_), .B0(ori_ori_n104_), .Y(ori02));
  NO2        o089(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n106_));
  NO2        o090(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n107_));
  NA2        o091(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n108_));
  NA2        o092(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n109_));
  INV        o093(.A(ori_ori_n109_), .Y(ori_ori_n110_));
  AOI220     o094(.A0(ori_ori_n110_), .A1(ori_ori_n107_), .B0(ori_ori_n106_), .B1(x4), .Y(ori_ori_n111_));
  NO3        o095(.A(ori_ori_n111_), .B(x7), .C(x5), .Y(ori_ori_n112_));
  NA2        o096(.A(x9), .B(x2), .Y(ori_ori_n113_));
  OR2        o097(.A(x8), .B(x0), .Y(ori_ori_n114_));
  INV        o098(.A(ori_ori_n114_), .Y(ori_ori_n115_));
  NAi21      o099(.An(x2), .B(x8), .Y(ori_ori_n116_));
  INV        o100(.A(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o101(.A(x4), .B(x1), .Y(ori_ori_n118_));
  NA3        o102(.A(ori_ori_n118_), .B(x2), .C(ori_ori_n60_), .Y(ori_ori_n119_));
  NOi21      o103(.An(x0), .B(x1), .Y(ori_ori_n120_));
  NO3        o104(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n121_));
  NOi21      o105(.An(x0), .B(x4), .Y(ori_ori_n122_));
  NAi21      o106(.An(x8), .B(x7), .Y(ori_ori_n123_));
  NO2        o107(.A(ori_ori_n123_), .B(ori_ori_n62_), .Y(ori_ori_n124_));
  AOI220     o108(.A0(ori_ori_n124_), .A1(ori_ori_n122_), .B0(ori_ori_n121_), .B1(ori_ori_n120_), .Y(ori_ori_n125_));
  AOI210     o109(.A0(ori_ori_n125_), .A1(ori_ori_n119_), .B0(ori_ori_n76_), .Y(ori_ori_n126_));
  NO2        o110(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n127_));
  NA2        o111(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n128_));
  AOI210     o112(.A0(ori_ori_n128_), .A1(ori_ori_n102_), .B0(ori_ori_n109_), .Y(ori_ori_n129_));
  OAI210     o113(.A0(ori_ori_n129_), .A1(ori_ori_n35_), .B0(ori_ori_n127_), .Y(ori_ori_n130_));
  NAi21      o114(.An(x0), .B(x4), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n131_), .B(x1), .Y(ori_ori_n132_));
  NO2        o116(.A(x7), .B(x0), .Y(ori_ori_n133_));
  NO2        o117(.A(ori_ori_n82_), .B(ori_ori_n96_), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n134_), .B(x3), .Y(ori_ori_n135_));
  OAI210     o119(.A0(ori_ori_n133_), .A1(ori_ori_n132_), .B0(ori_ori_n135_), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n137_));
  NA2        o121(.A(x5), .B(x0), .Y(ori_ori_n138_));
  NO2        o122(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n139_));
  NA3        o123(.A(ori_ori_n139_), .B(ori_ori_n138_), .C(ori_ori_n137_), .Y(ori_ori_n140_));
  NA4        o124(.A(ori_ori_n140_), .B(ori_ori_n136_), .C(ori_ori_n130_), .D(ori_ori_n36_), .Y(ori_ori_n141_));
  NO3        o125(.A(ori_ori_n141_), .B(ori_ori_n126_), .C(ori_ori_n112_), .Y(ori_ori_n142_));
  NO3        o126(.A(ori_ori_n76_), .B(ori_ori_n74_), .C(ori_ori_n24_), .Y(ori_ori_n143_));
  NO2        o127(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n144_));
  NA2        o128(.A(x7), .B(x3), .Y(ori_ori_n145_));
  NO2        o129(.A(ori_ori_n95_), .B(x5), .Y(ori_ori_n146_));
  NO2        o130(.A(x9), .B(x7), .Y(ori_ori_n147_));
  NOi21      o131(.An(x8), .B(x0), .Y(ori_ori_n148_));
  OA210      o132(.A0(ori_ori_n147_), .A1(x1), .B0(ori_ori_n148_), .Y(ori_ori_n149_));
  NO2        o133(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n150_));
  INV        o134(.A(x7), .Y(ori_ori_n151_));
  NA2        o135(.A(ori_ori_n151_), .B(ori_ori_n18_), .Y(ori_ori_n152_));
  AOI220     o136(.A0(ori_ori_n152_), .A1(ori_ori_n150_), .B0(ori_ori_n106_), .B1(ori_ori_n38_), .Y(ori_ori_n153_));
  NO2        o137(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n154_));
  NO2        o138(.A(ori_ori_n154_), .B(ori_ori_n122_), .Y(ori_ori_n155_));
  NO2        o139(.A(ori_ori_n155_), .B(ori_ori_n153_), .Y(ori_ori_n156_));
  AOI210     o140(.A0(ori_ori_n149_), .A1(ori_ori_n146_), .B0(ori_ori_n156_), .Y(ori_ori_n157_));
  OAI210     o141(.A0(ori_ori_n145_), .A1(ori_ori_n50_), .B0(ori_ori_n157_), .Y(ori_ori_n158_));
  NA2        o142(.A(x5), .B(x1), .Y(ori_ori_n159_));
  INV        o143(.A(ori_ori_n159_), .Y(ori_ori_n160_));
  AOI210     o144(.A0(ori_ori_n160_), .A1(ori_ori_n122_), .B0(ori_ori_n36_), .Y(ori_ori_n161_));
  NO2        o145(.A(ori_ori_n62_), .B(ori_ori_n88_), .Y(ori_ori_n162_));
  NAi21      o146(.An(x2), .B(x7), .Y(ori_ori_n163_));
  NO2        o147(.A(ori_ori_n163_), .B(ori_ori_n48_), .Y(ori_ori_n164_));
  NA2        o148(.A(ori_ori_n164_), .B(ori_ori_n65_), .Y(ori_ori_n165_));
  NAi31      o149(.An(ori_ori_n76_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n166_));
  NA3        o150(.A(ori_ori_n166_), .B(ori_ori_n165_), .C(ori_ori_n161_), .Y(ori_ori_n167_));
  NO3        o151(.A(ori_ori_n167_), .B(ori_ori_n158_), .C(ori_ori_n143_), .Y(ori_ori_n168_));
  NO2        o152(.A(ori_ori_n168_), .B(ori_ori_n142_), .Y(ori_ori_n169_));
  NO2        o153(.A(ori_ori_n138_), .B(ori_ori_n134_), .Y(ori_ori_n170_));
  NA2        o154(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n171_));
  NA2        o155(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n172_));
  NA3        o156(.A(ori_ori_n172_), .B(ori_ori_n171_), .C(ori_ori_n24_), .Y(ori_ori_n173_));
  AN2        o157(.A(ori_ori_n173_), .B(ori_ori_n139_), .Y(ori_ori_n174_));
  NA2        o158(.A(x8), .B(x0), .Y(ori_ori_n175_));
  NO2        o159(.A(ori_ori_n151_), .B(ori_ori_n25_), .Y(ori_ori_n176_));
  NO2        o160(.A(ori_ori_n120_), .B(x4), .Y(ori_ori_n177_));
  NA2        o161(.A(ori_ori_n177_), .B(ori_ori_n176_), .Y(ori_ori_n178_));
  AOI210     o162(.A0(ori_ori_n175_), .A1(ori_ori_n128_), .B0(ori_ori_n178_), .Y(ori_ori_n179_));
  NA2        o163(.A(x2), .B(x0), .Y(ori_ori_n180_));
  NA2        o164(.A(x4), .B(x1), .Y(ori_ori_n181_));
  NAi21      o165(.An(ori_ori_n118_), .B(ori_ori_n181_), .Y(ori_ori_n182_));
  NOi31      o166(.An(ori_ori_n182_), .B(ori_ori_n154_), .C(ori_ori_n180_), .Y(ori_ori_n183_));
  NO4        o167(.A(ori_ori_n183_), .B(ori_ori_n179_), .C(ori_ori_n174_), .D(ori_ori_n170_), .Y(ori_ori_n184_));
  NO2        o168(.A(ori_ori_n184_), .B(ori_ori_n43_), .Y(ori_ori_n185_));
  NO2        o169(.A(ori_ori_n173_), .B(ori_ori_n74_), .Y(ori_ori_n186_));
  INV        o170(.A(ori_ori_n127_), .Y(ori_ori_n187_));
  NO2        o171(.A(ori_ori_n102_), .B(ori_ori_n17_), .Y(ori_ori_n188_));
  AOI210     o172(.A0(ori_ori_n35_), .A1(ori_ori_n88_), .B0(ori_ori_n188_), .Y(ori_ori_n189_));
  NO3        o173(.A(ori_ori_n189_), .B(ori_ori_n187_), .C(x7), .Y(ori_ori_n190_));
  NA3        o174(.A(ori_ori_n182_), .B(ori_ori_n187_), .C(ori_ori_n42_), .Y(ori_ori_n191_));
  OAI210     o175(.A0(ori_ori_n172_), .A1(ori_ori_n134_), .B0(ori_ori_n191_), .Y(ori_ori_n192_));
  NO3        o176(.A(ori_ori_n192_), .B(ori_ori_n190_), .C(ori_ori_n186_), .Y(ori_ori_n193_));
  NO2        o177(.A(ori_ori_n193_), .B(x3), .Y(ori_ori_n194_));
  NO3        o178(.A(ori_ori_n194_), .B(ori_ori_n185_), .C(ori_ori_n169_), .Y(ori03));
  NO2        o179(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n196_));
  NO2        o180(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n197_));
  NO2        o181(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n198_));
  NO2        o182(.A(ori_ori_n76_), .B(x6), .Y(ori_ori_n199_));
  NA2        o183(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n200_));
  NO2        o184(.A(ori_ori_n200_), .B(x4), .Y(ori_ori_n201_));
  NO2        o185(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n202_));
  AO220      o186(.A0(ori_ori_n202_), .A1(ori_ori_n201_), .B0(ori_ori_n199_), .B1(ori_ori_n55_), .Y(ori_ori_n203_));
  NA2        o187(.A(ori_ori_n203_), .B(ori_ori_n62_), .Y(ori_ori_n204_));
  NA2        o188(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n205_));
  NO2        o189(.A(ori_ori_n205_), .B(ori_ori_n200_), .Y(ori_ori_n206_));
  NA2        o190(.A(x9), .B(ori_ori_n54_), .Y(ori_ori_n207_));
  NA2        o191(.A(ori_ori_n207_), .B(x4), .Y(ori_ori_n208_));
  NA2        o192(.A(ori_ori_n200_), .B(ori_ori_n79_), .Y(ori_ori_n209_));
  AOI210     o193(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n180_), .Y(ori_ori_n210_));
  AOI220     o194(.A0(ori_ori_n210_), .A1(ori_ori_n209_), .B0(ori_ori_n208_), .B1(ori_ori_n206_), .Y(ori_ori_n211_));
  NO3        o195(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n212_));
  NO2        o196(.A(x5), .B(x1), .Y(ori_ori_n213_));
  NO2        o197(.A(ori_ori_n205_), .B(ori_ori_n171_), .Y(ori_ori_n214_));
  NO3        o198(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n215_));
  NO2        o199(.A(ori_ori_n215_), .B(ori_ori_n214_), .Y(ori_ori_n216_));
  INV        o200(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  AOI220     o201(.A0(ori_ori_n217_), .A1(ori_ori_n48_), .B0(ori_ori_n212_), .B1(ori_ori_n127_), .Y(ori_ori_n218_));
  NA3        o202(.A(ori_ori_n218_), .B(ori_ori_n211_), .C(ori_ori_n204_), .Y(ori_ori_n219_));
  NO2        o203(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n220_));
  NA2        o204(.A(ori_ori_n220_), .B(ori_ori_n19_), .Y(ori_ori_n221_));
  NO2        o205(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n222_));
  NO2        o206(.A(ori_ori_n222_), .B(x6), .Y(ori_ori_n223_));
  NOi21      o207(.An(ori_ori_n82_), .B(ori_ori_n223_), .Y(ori_ori_n224_));
  NA2        o208(.A(ori_ori_n62_), .B(ori_ori_n88_), .Y(ori_ori_n225_));
  NA3        o209(.A(ori_ori_n225_), .B(ori_ori_n222_), .C(x6), .Y(ori_ori_n226_));
  AOI210     o210(.A0(ori_ori_n226_), .A1(ori_ori_n224_), .B0(ori_ori_n151_), .Y(ori_ori_n227_));
  AO210      o211(.A0(ori_ori_n227_), .A1(ori_ori_n221_), .B0(ori_ori_n176_), .Y(ori_ori_n228_));
  NA2        o212(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n229_));
  OAI210     o213(.A0(ori_ori_n229_), .A1(ori_ori_n25_), .B0(ori_ori_n172_), .Y(ori_ori_n230_));
  NO3        o214(.A(ori_ori_n181_), .B(ori_ori_n62_), .C(x6), .Y(ori_ori_n231_));
  AOI220     o215(.A0(ori_ori_n231_), .A1(ori_ori_n230_), .B0(ori_ori_n139_), .B1(ori_ori_n87_), .Y(ori_ori_n232_));
  NA2        o216(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n233_));
  OAI210     o217(.A0(ori_ori_n115_), .A1(ori_ori_n77_), .B0(x4), .Y(ori_ori_n234_));
  AOI210     o218(.A0(ori_ori_n234_), .A1(ori_ori_n233_), .B0(ori_ori_n76_), .Y(ori_ori_n235_));
  NO2        o219(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n236_));
  NO2        o220(.A(ori_ori_n159_), .B(ori_ori_n43_), .Y(ori_ori_n237_));
  OAI210     o221(.A0(ori_ori_n237_), .A1(ori_ori_n214_), .B0(ori_ori_n236_), .Y(ori_ori_n238_));
  NA2        o222(.A(ori_ori_n197_), .B(ori_ori_n132_), .Y(ori_ori_n239_));
  NA3        o223(.A(ori_ori_n205_), .B(ori_ori_n127_), .C(x6), .Y(ori_ori_n240_));
  OAI210     o224(.A0(ori_ori_n88_), .A1(ori_ori_n36_), .B0(ori_ori_n65_), .Y(ori_ori_n241_));
  NA4        o225(.A(ori_ori_n241_), .B(ori_ori_n240_), .C(ori_ori_n239_), .D(ori_ori_n238_), .Y(ori_ori_n242_));
  OAI210     o226(.A0(ori_ori_n242_), .A1(ori_ori_n235_), .B0(x2), .Y(ori_ori_n243_));
  NA3        o227(.A(ori_ori_n243_), .B(ori_ori_n232_), .C(ori_ori_n228_), .Y(ori_ori_n244_));
  AOI210     o228(.A0(ori_ori_n219_), .A1(x8), .B0(ori_ori_n244_), .Y(ori_ori_n245_));
  NO2        o229(.A(ori_ori_n88_), .B(x3), .Y(ori_ori_n246_));
  NA2        o230(.A(ori_ori_n246_), .B(ori_ori_n201_), .Y(ori_ori_n247_));
  NO3        o231(.A(ori_ori_n86_), .B(ori_ori_n77_), .C(ori_ori_n25_), .Y(ori_ori_n248_));
  AOI210     o232(.A0(ori_ori_n223_), .A1(ori_ori_n154_), .B0(ori_ori_n248_), .Y(ori_ori_n249_));
  AOI210     o233(.A0(ori_ori_n249_), .A1(ori_ori_n247_), .B0(x2), .Y(ori_ori_n250_));
  NO2        o234(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n251_));
  AOI220     o235(.A0(ori_ori_n201_), .A1(ori_ori_n188_), .B0(ori_ori_n251_), .B1(ori_ori_n65_), .Y(ori_ori_n252_));
  NA2        o236(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n253_));
  NA3        o237(.A(ori_ori_n25_), .B(x3), .C(x2), .Y(ori_ori_n254_));
  AOI210     o238(.A0(ori_ori_n254_), .A1(ori_ori_n138_), .B0(ori_ori_n253_), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n256_));
  NO2        o240(.A(ori_ori_n256_), .B(ori_ori_n25_), .Y(ori_ori_n257_));
  OAI210     o241(.A0(ori_ori_n257_), .A1(ori_ori_n255_), .B0(ori_ori_n118_), .Y(ori_ori_n258_));
  NA2        o242(.A(ori_ori_n205_), .B(x6), .Y(ori_ori_n259_));
  NO2        o243(.A(ori_ori_n205_), .B(x6), .Y(ori_ori_n260_));
  NAi21      o244(.An(ori_ori_n162_), .B(ori_ori_n260_), .Y(ori_ori_n261_));
  NA3        o245(.A(ori_ori_n261_), .B(ori_ori_n259_), .C(ori_ori_n144_), .Y(ori_ori_n262_));
  NA4        o246(.A(ori_ori_n262_), .B(ori_ori_n258_), .C(ori_ori_n252_), .D(ori_ori_n151_), .Y(ori_ori_n263_));
  NA2        o247(.A(ori_ori_n197_), .B(ori_ori_n222_), .Y(ori_ori_n264_));
  NO2        o248(.A(x9), .B(x6), .Y(ori_ori_n265_));
  NO2        o249(.A(ori_ori_n138_), .B(ori_ori_n18_), .Y(ori_ori_n266_));
  NAi21      o250(.An(ori_ori_n266_), .B(ori_ori_n254_), .Y(ori_ori_n267_));
  NAi21      o251(.An(x1), .B(x4), .Y(ori_ori_n268_));
  AOI210     o252(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n269_));
  OAI210     o253(.A0(ori_ori_n138_), .A1(x3), .B0(ori_ori_n269_), .Y(ori_ori_n270_));
  AOI220     o254(.A0(ori_ori_n270_), .A1(ori_ori_n268_), .B0(ori_ori_n267_), .B1(ori_ori_n265_), .Y(ori_ori_n271_));
  NA2        o255(.A(ori_ori_n271_), .B(ori_ori_n264_), .Y(ori_ori_n272_));
  NA2        o256(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n273_));
  NO3        o257(.A(x9), .B(x6), .C(x0), .Y(ori_ori_n274_));
  NA2        o258(.A(x6), .B(x2), .Y(ori_ori_n275_));
  NO2        o259(.A(ori_ori_n177_), .B(ori_ori_n46_), .Y(ori_ori_n276_));
  NA2        o260(.A(ori_ori_n276_), .B(ori_ori_n272_), .Y(ori_ori_n277_));
  NA2        o261(.A(x9), .B(ori_ori_n43_), .Y(ori_ori_n278_));
  NO2        o262(.A(ori_ori_n278_), .B(ori_ori_n200_), .Y(ori_ori_n279_));
  OR3        o263(.A(ori_ori_n279_), .B(ori_ori_n199_), .C(ori_ori_n146_), .Y(ori_ori_n280_));
  NA2        o264(.A(x4), .B(x0), .Y(ori_ori_n281_));
  NA2        o265(.A(ori_ori_n280_), .B(ori_ori_n42_), .Y(ori_ori_n282_));
  AOI210     o266(.A0(ori_ori_n282_), .A1(ori_ori_n277_), .B0(x8), .Y(ori_ori_n283_));
  INV        o267(.A(ori_ori_n253_), .Y(ori_ori_n284_));
  OAI210     o268(.A0(ori_ori_n266_), .A1(ori_ori_n213_), .B0(ori_ori_n284_), .Y(ori_ori_n285_));
  INV        o269(.A(ori_ori_n175_), .Y(ori_ori_n286_));
  OAI210     o270(.A0(ori_ori_n286_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n287_));
  AOI210     o271(.A0(ori_ori_n287_), .A1(ori_ori_n285_), .B0(ori_ori_n229_), .Y(ori_ori_n288_));
  NO4        o272(.A(ori_ori_n288_), .B(ori_ori_n283_), .C(ori_ori_n263_), .D(ori_ori_n250_), .Y(ori_ori_n289_));
  NO2        o273(.A(ori_ori_n162_), .B(x1), .Y(ori_ori_n290_));
  NO3        o274(.A(ori_ori_n290_), .B(x3), .C(ori_ori_n36_), .Y(ori_ori_n291_));
  OAI210     o275(.A0(ori_ori_n291_), .A1(ori_ori_n260_), .B0(x2), .Y(ori_ori_n292_));
  OAI210     o276(.A0(ori_ori_n286_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n293_));
  AOI210     o277(.A0(ori_ori_n293_), .A1(ori_ori_n292_), .B0(ori_ori_n187_), .Y(ori_ori_n294_));
  NOi21      o278(.An(ori_ori_n275_), .B(ori_ori_n17_), .Y(ori_ori_n295_));
  NA3        o279(.A(ori_ori_n295_), .B(ori_ori_n213_), .C(ori_ori_n40_), .Y(ori_ori_n296_));
  AOI210     o280(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n297_));
  NA3        o281(.A(ori_ori_n297_), .B(ori_ori_n160_), .C(ori_ori_n32_), .Y(ori_ori_n298_));
  NA2        o282(.A(x3), .B(x2), .Y(ori_ori_n299_));
  AOI220     o283(.A0(ori_ori_n299_), .A1(ori_ori_n229_), .B0(ori_ori_n298_), .B1(ori_ori_n296_), .Y(ori_ori_n300_));
  NAi21      o284(.An(x4), .B(x0), .Y(ori_ori_n301_));
  NO3        o285(.A(ori_ori_n301_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n302_));
  OAI210     o286(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n302_), .Y(ori_ori_n303_));
  OAI220     o287(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n304_));
  NO2        o288(.A(x9), .B(x8), .Y(ori_ori_n305_));
  NO2        o289(.A(ori_ori_n297_), .B(ori_ori_n295_), .Y(ori_ori_n306_));
  AOI220     o290(.A0(ori_ori_n306_), .A1(ori_ori_n80_), .B0(ori_ori_n304_), .B1(ori_ori_n31_), .Y(ori_ori_n307_));
  AOI210     o291(.A0(ori_ori_n307_), .A1(ori_ori_n303_), .B0(ori_ori_n25_), .Y(ori_ori_n308_));
  NA3        o292(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n309_));
  OAI210     o293(.A0(ori_ori_n297_), .A1(ori_ori_n295_), .B0(ori_ori_n309_), .Y(ori_ori_n310_));
  INV        o294(.A(ori_ori_n214_), .Y(ori_ori_n311_));
  NA2        o295(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n312_));
  OR2        o296(.A(ori_ori_n312_), .B(ori_ori_n281_), .Y(ori_ori_n313_));
  OAI220     o297(.A0(ori_ori_n313_), .A1(ori_ori_n159_), .B0(ori_ori_n233_), .B1(ori_ori_n311_), .Y(ori_ori_n314_));
  AO210      o298(.A0(ori_ori_n310_), .A1(ori_ori_n146_), .B0(ori_ori_n314_), .Y(ori_ori_n315_));
  NO4        o299(.A(ori_ori_n315_), .B(ori_ori_n308_), .C(ori_ori_n300_), .D(ori_ori_n294_), .Y(ori_ori_n316_));
  OAI210     o300(.A0(ori_ori_n289_), .A1(ori_ori_n245_), .B0(ori_ori_n316_), .Y(ori04));
  OAI210     o301(.A0(x8), .A1(ori_ori_n18_), .B0(x4), .Y(ori_ori_n318_));
  NA3        o302(.A(ori_ori_n318_), .B(ori_ori_n274_), .C(ori_ori_n83_), .Y(ori_ori_n319_));
  NO2        o303(.A(x2), .B(x1), .Y(ori_ori_n320_));
  OAI210     o304(.A0(ori_ori_n256_), .A1(ori_ori_n320_), .B0(ori_ori_n36_), .Y(ori_ori_n321_));
  NO2        o305(.A(ori_ori_n320_), .B(ori_ori_n301_), .Y(ori_ori_n322_));
  AOI210     o306(.A0(ori_ori_n62_), .A1(x4), .B0(ori_ori_n108_), .Y(ori_ori_n323_));
  OAI210     o307(.A0(ori_ori_n323_), .A1(ori_ori_n322_), .B0(ori_ori_n246_), .Y(ori_ori_n324_));
  NO2        o308(.A(ori_ori_n273_), .B(ori_ori_n86_), .Y(ori_ori_n325_));
  NO2        o309(.A(ori_ori_n325_), .B(ori_ori_n36_), .Y(ori_ori_n326_));
  NO2        o310(.A(ori_ori_n299_), .B(ori_ori_n202_), .Y(ori_ori_n327_));
  NA2        o311(.A(x9), .B(x0), .Y(ori_ori_n328_));
  AOI210     o312(.A0(ori_ori_n86_), .A1(ori_ori_n74_), .B0(ori_ori_n328_), .Y(ori_ori_n329_));
  OAI210     o313(.A0(ori_ori_n329_), .A1(ori_ori_n327_), .B0(ori_ori_n88_), .Y(ori_ori_n330_));
  NA3        o314(.A(ori_ori_n330_), .B(ori_ori_n326_), .C(ori_ori_n324_), .Y(ori_ori_n331_));
  NA2        o315(.A(ori_ori_n331_), .B(ori_ori_n321_), .Y(ori_ori_n332_));
  NO2        o316(.A(ori_ori_n207_), .B(ori_ori_n109_), .Y(ori_ori_n333_));
  NO3        o317(.A(ori_ori_n253_), .B(ori_ori_n116_), .C(ori_ori_n18_), .Y(ori_ori_n334_));
  NO2        o318(.A(ori_ori_n334_), .B(ori_ori_n333_), .Y(ori_ori_n335_));
  OAI210     o319(.A0(ori_ori_n114_), .A1(ori_ori_n102_), .B0(ori_ori_n175_), .Y(ori_ori_n336_));
  NA3        o320(.A(ori_ori_n336_), .B(x6), .C(x3), .Y(ori_ori_n337_));
  NOi21      o321(.An(ori_ori_n148_), .B(ori_ori_n128_), .Y(ori_ori_n338_));
  AOI210     o322(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n339_));
  OAI220     o323(.A0(ori_ori_n339_), .A1(ori_ori_n312_), .B0(ori_ori_n273_), .B1(ori_ori_n309_), .Y(ori_ori_n340_));
  AOI210     o324(.A0(ori_ori_n338_), .A1(ori_ori_n63_), .B0(ori_ori_n340_), .Y(ori_ori_n341_));
  NA2        o325(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n342_));
  OAI210     o326(.A0(ori_ori_n102_), .A1(ori_ori_n17_), .B0(ori_ori_n342_), .Y(ori_ori_n343_));
  AOI220     o327(.A0(ori_ori_n343_), .A1(ori_ori_n77_), .B0(ori_ori_n325_), .B1(ori_ori_n88_), .Y(ori_ori_n344_));
  NA4        o328(.A(ori_ori_n344_), .B(ori_ori_n341_), .C(ori_ori_n337_), .D(ori_ori_n335_), .Y(ori_ori_n345_));
  OAI210     o329(.A0(ori_ori_n107_), .A1(x3), .B0(ori_ori_n302_), .Y(ori_ori_n346_));
  NA2        o330(.A(ori_ori_n212_), .B(ori_ori_n82_), .Y(ori_ori_n347_));
  NA3        o331(.A(ori_ori_n347_), .B(ori_ori_n346_), .C(ori_ori_n151_), .Y(ori_ori_n348_));
  AOI210     o332(.A0(ori_ori_n345_), .A1(x4), .B0(ori_ori_n348_), .Y(ori_ori_n349_));
  NA3        o333(.A(ori_ori_n322_), .B(ori_ori_n207_), .C(ori_ori_n88_), .Y(ori_ori_n350_));
  NOi21      o334(.An(x4), .B(x0), .Y(ori_ori_n351_));
  XO2        o335(.A(x4), .B(x0), .Y(ori_ori_n352_));
  OAI210     o336(.A0(ori_ori_n352_), .A1(ori_ori_n113_), .B0(ori_ori_n268_), .Y(ori_ori_n353_));
  AOI220     o337(.A0(ori_ori_n353_), .A1(x8), .B0(ori_ori_n351_), .B1(ori_ori_n89_), .Y(ori_ori_n354_));
  AOI210     o338(.A0(ori_ori_n354_), .A1(ori_ori_n350_), .B0(x3), .Y(ori_ori_n355_));
  INV        o339(.A(ori_ori_n89_), .Y(ori_ori_n356_));
  NO2        o340(.A(ori_ori_n88_), .B(x4), .Y(ori_ori_n357_));
  AOI220     o341(.A0(ori_ori_n357_), .A1(ori_ori_n44_), .B0(ori_ori_n122_), .B1(ori_ori_n356_), .Y(ori_ori_n358_));
  NO3        o342(.A(ori_ori_n352_), .B(ori_ori_n162_), .C(x2), .Y(ori_ori_n359_));
  NO3        o343(.A(ori_ori_n225_), .B(ori_ori_n28_), .C(ori_ori_n24_), .Y(ori_ori_n360_));
  NO2        o344(.A(ori_ori_n360_), .B(ori_ori_n359_), .Y(ori_ori_n361_));
  NA4        o345(.A(ori_ori_n361_), .B(ori_ori_n358_), .C(ori_ori_n221_), .D(x6), .Y(ori_ori_n362_));
  OAI220     o346(.A0(ori_ori_n301_), .A1(ori_ori_n86_), .B0(ori_ori_n180_), .B1(ori_ori_n88_), .Y(ori_ori_n363_));
  NO2        o347(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n364_));
  OR2        o348(.A(ori_ori_n357_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  NO2        o349(.A(ori_ori_n148_), .B(ori_ori_n102_), .Y(ori_ori_n366_));
  AOI220     o350(.A0(ori_ori_n366_), .A1(ori_ori_n365_), .B0(ori_ori_n363_), .B1(ori_ori_n61_), .Y(ori_ori_n367_));
  NO2        o351(.A(ori_ori_n148_), .B(ori_ori_n79_), .Y(ori_ori_n368_));
  NO2        o352(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n369_));
  NOi21      o353(.An(ori_ori_n118_), .B(ori_ori_n27_), .Y(ori_ori_n370_));
  AOI210     o354(.A0(ori_ori_n369_), .A1(ori_ori_n368_), .B0(ori_ori_n370_), .Y(ori_ori_n371_));
  OAI210     o355(.A0(ori_ori_n367_), .A1(ori_ori_n62_), .B0(ori_ori_n371_), .Y(ori_ori_n372_));
  OAI220     o356(.A0(ori_ori_n372_), .A1(x6), .B0(ori_ori_n362_), .B1(ori_ori_n355_), .Y(ori_ori_n373_));
  OAI210     o357(.A0(ori_ori_n63_), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n374_));
  OAI210     o358(.A0(ori_ori_n374_), .A1(ori_ori_n88_), .B0(ori_ori_n313_), .Y(ori_ori_n375_));
  AOI210     o359(.A0(ori_ori_n375_), .A1(ori_ori_n18_), .B0(ori_ori_n151_), .Y(ori_ori_n376_));
  AO220      o360(.A0(ori_ori_n376_), .A1(ori_ori_n373_), .B0(ori_ori_n349_), .B1(ori_ori_n332_), .Y(ori_ori_n377_));
  NA2        o361(.A(ori_ori_n369_), .B(x6), .Y(ori_ori_n378_));
  AOI210     o362(.A0(x6), .A1(x1), .B0(ori_ori_n150_), .Y(ori_ori_n379_));
  NA2        o363(.A(ori_ori_n357_), .B(x0), .Y(ori_ori_n380_));
  NA2        o364(.A(ori_ori_n82_), .B(x6), .Y(ori_ori_n381_));
  OAI210     o365(.A0(ori_ori_n380_), .A1(ori_ori_n379_), .B0(ori_ori_n381_), .Y(ori_ori_n382_));
  AOI220     o366(.A0(ori_ori_n382_), .A1(ori_ori_n378_), .B0(ori_ori_n215_), .B1(ori_ori_n49_), .Y(ori_ori_n383_));
  NA3        o367(.A(ori_ori_n383_), .B(ori_ori_n377_), .C(ori_ori_n319_), .Y(ori_ori_n384_));
  AOI210     o368(.A0(ori_ori_n198_), .A1(x8), .B0(ori_ori_n107_), .Y(ori_ori_n385_));
  NA2        o369(.A(ori_ori_n385_), .B(ori_ori_n342_), .Y(ori_ori_n386_));
  NA3        o370(.A(ori_ori_n386_), .B(ori_ori_n196_), .C(ori_ori_n151_), .Y(ori_ori_n387_));
  OAI210     o371(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n229_), .Y(ori_ori_n388_));
  AO220      o372(.A0(ori_ori_n388_), .A1(ori_ori_n147_), .B0(ori_ori_n106_), .B1(x4), .Y(ori_ori_n389_));
  NA3        o373(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n390_));
  NA2        o374(.A(ori_ori_n220_), .B(x0), .Y(ori_ori_n391_));
  OAI220     o375(.A0(ori_ori_n391_), .A1(ori_ori_n207_), .B0(ori_ori_n390_), .B1(ori_ori_n356_), .Y(ori_ori_n392_));
  AOI210     o376(.A0(ori_ori_n389_), .A1(ori_ori_n115_), .B0(ori_ori_n392_), .Y(ori_ori_n393_));
  AOI210     o377(.A0(ori_ori_n393_), .A1(ori_ori_n387_), .B0(ori_ori_n25_), .Y(ori_ori_n394_));
  NA3        o378(.A(ori_ori_n117_), .B(ori_ori_n220_), .C(x0), .Y(ori_ori_n395_));
  OAI210     o379(.A0(ori_ori_n196_), .A1(ori_ori_n66_), .B0(ori_ori_n202_), .Y(ori_ori_n396_));
  NA3        o380(.A(ori_ori_n198_), .B(ori_ori_n222_), .C(x8), .Y(ori_ori_n397_));
  AOI210     o381(.A0(ori_ori_n397_), .A1(ori_ori_n396_), .B0(ori_ori_n25_), .Y(ori_ori_n398_));
  AOI210     o382(.A0(ori_ori_n116_), .A1(ori_ori_n114_), .B0(ori_ori_n42_), .Y(ori_ori_n399_));
  NOi31      o383(.An(ori_ori_n399_), .B(ori_ori_n364_), .C(ori_ori_n181_), .Y(ori_ori_n400_));
  OAI210     o384(.A0(ori_ori_n400_), .A1(ori_ori_n398_), .B0(ori_ori_n147_), .Y(ori_ori_n401_));
  NAi31      o385(.An(ori_ori_n50_), .B(ori_ori_n290_), .C(ori_ori_n176_), .Y(ori_ori_n402_));
  NA3        o386(.A(ori_ori_n402_), .B(ori_ori_n401_), .C(ori_ori_n395_), .Y(ori_ori_n403_));
  OAI210     o387(.A0(ori_ori_n403_), .A1(ori_ori_n394_), .B0(x6), .Y(ori_ori_n404_));
  OAI210     o388(.A0(ori_ori_n162_), .A1(ori_ori_n48_), .B0(ori_ori_n133_), .Y(ori_ori_n405_));
  NA3        o389(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n406_));
  AOI220     o390(.A0(ori_ori_n406_), .A1(ori_ori_n405_), .B0(ori_ori_n40_), .B1(ori_ori_n32_), .Y(ori_ori_n407_));
  NO2        o391(.A(ori_ori_n151_), .B(x0), .Y(ori_ori_n408_));
  AOI220     o392(.A0(ori_ori_n408_), .A1(ori_ori_n220_), .B0(ori_ori_n196_), .B1(ori_ori_n151_), .Y(ori_ori_n409_));
  AOI210     o393(.A0(ori_ori_n124_), .A1(ori_ori_n251_), .B0(x1), .Y(ori_ori_n410_));
  OAI210     o394(.A0(ori_ori_n409_), .A1(x8), .B0(ori_ori_n410_), .Y(ori_ori_n411_));
  NAi31      o395(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n412_));
  OAI210     o396(.A0(ori_ori_n412_), .A1(x4), .B0(ori_ori_n163_), .Y(ori_ori_n413_));
  NA3        o397(.A(ori_ori_n413_), .B(ori_ori_n145_), .C(x9), .Y(ori_ori_n414_));
  NO3        o398(.A(x9), .B(ori_ori_n151_), .C(x0), .Y(ori_ori_n415_));
  AOI220     o399(.A0(ori_ori_n415_), .A1(ori_ori_n246_), .B0(ori_ori_n368_), .B1(ori_ori_n151_), .Y(ori_ori_n416_));
  NA4        o400(.A(ori_ori_n416_), .B(x1), .C(ori_ori_n414_), .D(ori_ori_n50_), .Y(ori_ori_n417_));
  OAI210     o401(.A0(ori_ori_n411_), .A1(ori_ori_n407_), .B0(ori_ori_n417_), .Y(ori_ori_n418_));
  NOi31      o402(.An(ori_ori_n408_), .B(ori_ori_n32_), .C(x8), .Y(ori_ori_n419_));
  AOI210     o403(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n131_), .Y(ori_ori_n420_));
  NO3        o404(.A(ori_ori_n420_), .B(ori_ori_n121_), .C(ori_ori_n43_), .Y(ori_ori_n421_));
  NOi31      o405(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n422_));
  AOI220     o406(.A0(ori_ori_n422_), .A1(ori_ori_n351_), .B0(ori_ori_n122_), .B1(x3), .Y(ori_ori_n423_));
  AOI210     o407(.A0(ori_ori_n268_), .A1(ori_ori_n60_), .B0(ori_ori_n120_), .Y(ori_ori_n424_));
  OAI210     o408(.A0(ori_ori_n424_), .A1(x3), .B0(ori_ori_n423_), .Y(ori_ori_n425_));
  NO3        o409(.A(ori_ori_n425_), .B(ori_ori_n421_), .C(x2), .Y(ori_ori_n426_));
  OAI220     o410(.A0(ori_ori_n352_), .A1(ori_ori_n305_), .B0(ori_ori_n301_), .B1(ori_ori_n43_), .Y(ori_ori_n427_));
  AOI210     o411(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n390_), .Y(ori_ori_n428_));
  AOI220     o412(.A0(ori_ori_n428_), .A1(ori_ori_n88_), .B0(ori_ori_n427_), .B1(ori_ori_n151_), .Y(ori_ori_n429_));
  NO2        o413(.A(ori_ori_n429_), .B(ori_ori_n54_), .Y(ori_ori_n430_));
  NO3        o414(.A(ori_ori_n430_), .B(ori_ori_n426_), .C(ori_ori_n419_), .Y(ori_ori_n431_));
  AOI210     o415(.A0(ori_ori_n431_), .A1(ori_ori_n418_), .B0(ori_ori_n25_), .Y(ori_ori_n432_));
  NA4        o416(.A(ori_ori_n31_), .B(ori_ori_n88_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n433_));
  NO3        o417(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n434_));
  NO3        o418(.A(ori_ori_n66_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n435_));
  AOI220     o419(.A0(ori_ori_n435_), .A1(ori_ori_n269_), .B0(ori_ori_n434_), .B1(ori_ori_n399_), .Y(ori_ori_n436_));
  NO2        o420(.A(ori_ori_n436_), .B(ori_ori_n99_), .Y(ori_ori_n437_));
  NO3        o421(.A(ori_ori_n273_), .B(ori_ori_n175_), .C(ori_ori_n40_), .Y(ori_ori_n438_));
  OAI210     o422(.A0(ori_ori_n438_), .A1(ori_ori_n437_), .B0(x7), .Y(ori_ori_n439_));
  NA2        o423(.A(ori_ori_n225_), .B(x7), .Y(ori_ori_n440_));
  NA3        o424(.A(ori_ori_n440_), .B(ori_ori_n150_), .C(ori_ori_n132_), .Y(ori_ori_n441_));
  NA3        o425(.A(ori_ori_n441_), .B(ori_ori_n439_), .C(ori_ori_n433_), .Y(ori_ori_n442_));
  OAI210     o426(.A0(ori_ori_n442_), .A1(ori_ori_n432_), .B0(ori_ori_n36_), .Y(ori_ori_n443_));
  NO2        o427(.A(ori_ori_n415_), .B(ori_ori_n202_), .Y(ori_ori_n444_));
  NO4        o428(.A(ori_ori_n444_), .B(ori_ori_n76_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n445_));
  NA2        o429(.A(ori_ori_n256_), .B(ori_ori_n21_), .Y(ori_ori_n446_));
  NO2        o430(.A(ori_ori_n159_), .B(ori_ori_n133_), .Y(ori_ori_n447_));
  NA2        o431(.A(ori_ori_n447_), .B(ori_ori_n446_), .Y(ori_ori_n448_));
  AOI210     o432(.A0(ori_ori_n448_), .A1(ori_ori_n166_), .B0(ori_ori_n28_), .Y(ori_ori_n449_));
  AOI220     o433(.A0(ori_ori_n364_), .A1(ori_ori_n88_), .B0(ori_ori_n148_), .B1(ori_ori_n198_), .Y(ori_ori_n450_));
  NA3        o434(.A(ori_ori_n450_), .B(ori_ori_n412_), .C(ori_ori_n86_), .Y(ori_ori_n451_));
  NA2        o435(.A(ori_ori_n451_), .B(ori_ori_n176_), .Y(ori_ori_n452_));
  OAI220     o436(.A0(ori_ori_n278_), .A1(ori_ori_n67_), .B0(ori_ori_n159_), .B1(ori_ori_n43_), .Y(ori_ori_n453_));
  NA2        o437(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n454_));
  OAI210     o438(.A0(ori_ori_n147_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n455_));
  NO3        o439(.A(ori_ori_n422_), .B(x3), .C(ori_ori_n54_), .Y(ori_ori_n456_));
  NA2        o440(.A(ori_ori_n456_), .B(ori_ori_n455_), .Y(ori_ori_n457_));
  OAI210     o441(.A0(ori_ori_n152_), .A1(ori_ori_n454_), .B0(ori_ori_n457_), .Y(ori_ori_n458_));
  AOI220     o442(.A0(ori_ori_n458_), .A1(x0), .B0(ori_ori_n453_), .B1(ori_ori_n133_), .Y(ori_ori_n459_));
  AOI210     o443(.A0(ori_ori_n459_), .A1(ori_ori_n452_), .B0(ori_ori_n233_), .Y(ori_ori_n460_));
  NO3        o444(.A(ori_ori_n460_), .B(ori_ori_n449_), .C(ori_ori_n445_), .Y(ori_ori_n461_));
  NA3        o445(.A(ori_ori_n461_), .B(ori_ori_n443_), .C(ori_ori_n404_), .Y(ori_ori_n462_));
  AOI210     o446(.A0(ori_ori_n384_), .A1(ori_ori_n25_), .B0(ori_ori_n462_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  NO4        m012(.A(mai_mai_n28_), .B(mai_mai_n27_), .C(mai_mai_n26_), .D(mai_mai_n25_), .Y(mai_mai_n29_));
  NO2        m013(.A(mai_mai_n29_), .B(mai_mai_n24_), .Y(mai_mai_n30_));
  NO2        m014(.A(x4), .B(x3), .Y(mai_mai_n31_));
  INV        m015(.A(mai_mai_n31_), .Y(mai_mai_n32_));
  OA210      m016(.A0(mai_mai_n32_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n33_));
  NOi31      m017(.An(mai_mai_n23_), .B(mai_mai_n33_), .C(mai_mai_n30_), .Y(mai00));
  NO2        m018(.A(x1), .B(x0), .Y(mai_mai_n35_));
  INV        m019(.A(x6), .Y(mai_mai_n36_));
  NO2        m020(.A(mai_mai_n36_), .B(mai_mai_n25_), .Y(mai_mai_n37_));
  AN2        m021(.A(x8), .B(x7), .Y(mai_mai_n38_));
  NA3        m022(.A(mai_mai_n38_), .B(mai_mai_n37_), .C(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m023(.A(x4), .B(x3), .Y(mai_mai_n40_));
  AOI210     m024(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m025(.A(x2), .B(x0), .Y(mai_mai_n42_));
  INV        m026(.A(x3), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n44_));
  INV        m028(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO2        m029(.A(mai_mai_n37_), .B(x4), .Y(mai_mai_n46_));
  OAI210     m030(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n42_), .Y(mai_mai_n47_));
  INV        m031(.A(x4), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n49_), .B(x2), .Y(mai_mai_n50_));
  OAI210     m034(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n47_), .Y(mai_mai_n51_));
  NA2        m035(.A(mai_mai_n38_), .B(mai_mai_n37_), .Y(mai_mai_n52_));
  AOI220     m036(.A0(mai_mai_n52_), .A1(mai_mai_n35_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n53_));
  INV        m037(.A(x2), .Y(mai_mai_n54_));
  NO2        m038(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n55_));
  NA2        m039(.A(mai_mai_n43_), .B(mai_mai_n18_), .Y(mai_mai_n56_));
  NA2        m040(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  OAI210     m041(.A0(mai_mai_n53_), .A1(mai_mai_n32_), .B0(mai_mai_n57_), .Y(mai_mai_n58_));
  NO3        m042(.A(mai_mai_n58_), .B(mai_mai_n51_), .C(mai_mai_n41_), .Y(mai01));
  NA2        m043(.A(x8), .B(x7), .Y(mai_mai_n60_));
  NA2        m044(.A(mai_mai_n43_), .B(x1), .Y(mai_mai_n61_));
  INV        m045(.A(x9), .Y(mai_mai_n62_));
  NO2        m046(.A(mai_mai_n62_), .B(mai_mai_n36_), .Y(mai_mai_n63_));
  INV        m047(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  NO3        m048(.A(mai_mai_n64_), .B(mai_mai_n61_), .C(mai_mai_n60_), .Y(mai_mai_n65_));
  NO2        m049(.A(x7), .B(x6), .Y(mai_mai_n66_));
  NO2        m050(.A(mai_mai_n61_), .B(x5), .Y(mai_mai_n67_));
  NO2        m051(.A(x8), .B(x2), .Y(mai_mai_n68_));
  INV        m052(.A(mai_mai_n68_), .Y(mai_mai_n69_));
  AN2        m053(.A(mai_mai_n67_), .B(mai_mai_n66_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n44_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n71_));
  OAI210     m055(.A0(mai_mai_n56_), .A1(mai_mai_n20_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  NAi31      m056(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n73_));
  NO2        m057(.A(mai_mai_n72_), .B(mai_mai_n70_), .Y(mai_mai_n74_));
  OAI210     m058(.A0(mai_mai_n74_), .A1(mai_mai_n65_), .B0(x4), .Y(mai_mai_n75_));
  NA2        m059(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n76_));
  OAI210     m060(.A0(mai_mai_n76_), .A1(mai_mai_n56_), .B0(x0), .Y(mai_mai_n77_));
  NA2        m061(.A(x5), .B(x3), .Y(mai_mai_n78_));
  NO2        m062(.A(x8), .B(x6), .Y(mai_mai_n79_));
  NO4        m063(.A(mai_mai_n79_), .B(mai_mai_n78_), .C(mai_mai_n66_), .D(mai_mai_n54_), .Y(mai_mai_n80_));
  NAi21      m064(.An(x4), .B(x3), .Y(mai_mai_n81_));
  INV        m065(.A(mai_mai_n81_), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(mai_mai_n22_), .Y(mai_mai_n83_));
  NO2        m067(.A(x4), .B(x2), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(x3), .Y(mai_mai_n85_));
  NO3        m069(.A(mai_mai_n85_), .B(mai_mai_n83_), .C(mai_mai_n18_), .Y(mai_mai_n86_));
  NO3        m070(.A(mai_mai_n86_), .B(mai_mai_n80_), .C(mai_mai_n77_), .Y(mai_mai_n87_));
  NO4        m071(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n43_), .D(x1), .Y(mai_mai_n88_));
  NA2        m072(.A(mai_mai_n62_), .B(mai_mai_n48_), .Y(mai_mai_n89_));
  INV        m073(.A(mai_mai_n89_), .Y(mai_mai_n90_));
  OAI210     m074(.A0(mai_mai_n88_), .A1(mai_mai_n67_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  NA2        m075(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n92_));
  NO2        m076(.A(mai_mai_n92_), .B(mai_mai_n25_), .Y(mai_mai_n93_));
  INV        m077(.A(x8), .Y(mai_mai_n94_));
  NA2        m078(.A(x2), .B(x1), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n94_), .Y(mai_mai_n96_));
  NO2        m080(.A(mai_mai_n96_), .B(mai_mai_n93_), .Y(mai_mai_n97_));
  NO2        m081(.A(mai_mai_n97_), .B(mai_mai_n26_), .Y(mai_mai_n98_));
  AOI210     m082(.A0(mai_mai_n56_), .A1(mai_mai_n25_), .B0(mai_mai_n54_), .Y(mai_mai_n99_));
  OAI210     m083(.A0(mai_mai_n45_), .A1(mai_mai_n37_), .B0(mai_mai_n48_), .Y(mai_mai_n100_));
  NO3        m084(.A(mai_mai_n100_), .B(mai_mai_n99_), .C(mai_mai_n98_), .Y(mai_mai_n101_));
  NA2        m085(.A(x4), .B(mai_mai_n43_), .Y(mai_mai_n102_));
  NO2        m086(.A(mai_mai_n48_), .B(mai_mai_n54_), .Y(mai_mai_n103_));
  OAI210     m087(.A0(mai_mai_n103_), .A1(mai_mai_n43_), .B0(mai_mai_n18_), .Y(mai_mai_n104_));
  AOI210     m088(.A0(mai_mai_n102_), .A1(mai_mai_n52_), .B0(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m089(.A(x3), .B(x2), .Y(mai_mai_n106_));
  NA3        m090(.A(mai_mai_n106_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n107_));
  AOI210     m091(.A0(x8), .A1(x6), .B0(mai_mai_n107_), .Y(mai_mai_n108_));
  NA2        m092(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n109_));
  OAI210     m093(.A0(mai_mai_n109_), .A1(mai_mai_n40_), .B0(mai_mai_n17_), .Y(mai_mai_n110_));
  NO4        m094(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n105_), .D(mai_mai_n101_), .Y(mai_mai_n111_));
  AO220      m095(.A0(mai_mai_n111_), .A1(mai_mai_n91_), .B0(mai_mai_n87_), .B1(mai_mai_n75_), .Y(mai02));
  NO2        m096(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n113_));
  NO2        m097(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n114_));
  NA2        m098(.A(mai_mai_n54_), .B(mai_mai_n17_), .Y(mai_mai_n115_));
  NA2        m099(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n116_));
  OAI210     m100(.A0(mai_mai_n89_), .A1(mai_mai_n115_), .B0(mai_mai_n116_), .Y(mai_mai_n117_));
  AOI220     m101(.A0(mai_mai_n117_), .A1(mai_mai_n114_), .B0(mai_mai_n113_), .B1(x4), .Y(mai_mai_n118_));
  NO3        m102(.A(mai_mai_n118_), .B(x7), .C(x5), .Y(mai_mai_n119_));
  NA2        m103(.A(x9), .B(x2), .Y(mai_mai_n120_));
  OR2        m104(.A(x8), .B(x0), .Y(mai_mai_n121_));
  INV        m105(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  NAi21      m106(.An(x2), .B(x8), .Y(mai_mai_n123_));
  INV        m107(.A(mai_mai_n123_), .Y(mai_mai_n124_));
  OAI220     m108(.A0(mai_mai_n124_), .A1(mai_mai_n122_), .B0(mai_mai_n120_), .B1(x7), .Y(mai_mai_n125_));
  NO2        m109(.A(x4), .B(x1), .Y(mai_mai_n126_));
  NA3        m110(.A(mai_mai_n126_), .B(mai_mai_n125_), .C(mai_mai_n60_), .Y(mai_mai_n127_));
  NOi21      m111(.An(x0), .B(x1), .Y(mai_mai_n128_));
  NO3        m112(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n129_));
  NOi21      m113(.An(x0), .B(x4), .Y(mai_mai_n130_));
  NAi21      m114(.An(x8), .B(x7), .Y(mai_mai_n131_));
  NO2        m115(.A(mai_mai_n131_), .B(mai_mai_n62_), .Y(mai_mai_n132_));
  AOI220     m116(.A0(mai_mai_n132_), .A1(mai_mai_n130_), .B0(mai_mai_n129_), .B1(mai_mai_n128_), .Y(mai_mai_n133_));
  AOI210     m117(.A0(mai_mai_n133_), .A1(mai_mai_n127_), .B0(mai_mai_n78_), .Y(mai_mai_n134_));
  NO2        m118(.A(x5), .B(mai_mai_n48_), .Y(mai_mai_n135_));
  NA2        m119(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n136_));
  AOI210     m120(.A0(mai_mai_n136_), .A1(mai_mai_n109_), .B0(mai_mai_n116_), .Y(mai_mai_n137_));
  OAI210     m121(.A0(mai_mai_n137_), .A1(mai_mai_n35_), .B0(mai_mai_n135_), .Y(mai_mai_n138_));
  NAi21      m122(.An(x0), .B(x4), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n139_), .B(x1), .Y(mai_mai_n140_));
  NO2        m124(.A(x7), .B(x0), .Y(mai_mai_n141_));
  NO2        m125(.A(mai_mai_n84_), .B(mai_mai_n103_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n142_), .B(x3), .Y(mai_mai_n143_));
  OAI210     m127(.A0(mai_mai_n141_), .A1(mai_mai_n140_), .B0(mai_mai_n143_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n21_), .B(mai_mai_n43_), .Y(mai_mai_n145_));
  NA2        m129(.A(x5), .B(x0), .Y(mai_mai_n146_));
  NO2        m130(.A(mai_mai_n48_), .B(x2), .Y(mai_mai_n147_));
  NA3        m131(.A(mai_mai_n147_), .B(mai_mai_n146_), .C(mai_mai_n145_), .Y(mai_mai_n148_));
  NA4        m132(.A(mai_mai_n148_), .B(mai_mai_n144_), .C(mai_mai_n138_), .D(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m133(.A(mai_mai_n149_), .B(mai_mai_n134_), .C(mai_mai_n119_), .Y(mai_mai_n150_));
  NO3        m134(.A(mai_mai_n78_), .B(mai_mai_n76_), .C(mai_mai_n24_), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n152_));
  AOI220     m136(.A0(mai_mai_n128_), .A1(mai_mai_n152_), .B0(mai_mai_n67_), .B1(mai_mai_n17_), .Y(mai_mai_n153_));
  NO3        m137(.A(mai_mai_n153_), .B(mai_mai_n60_), .C(mai_mai_n62_), .Y(mai_mai_n154_));
  NA2        m138(.A(x7), .B(x3), .Y(mai_mai_n155_));
  NO2        m139(.A(mai_mai_n102_), .B(x5), .Y(mai_mai_n156_));
  NO2        m140(.A(x9), .B(x7), .Y(mai_mai_n157_));
  NOi21      m141(.An(x8), .B(x0), .Y(mai_mai_n158_));
  OA210      m142(.A0(mai_mai_n157_), .A1(x1), .B0(mai_mai_n158_), .Y(mai_mai_n159_));
  NO2        m143(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n160_));
  INV        m144(.A(x7), .Y(mai_mai_n161_));
  NA2        m145(.A(mai_mai_n161_), .B(mai_mai_n18_), .Y(mai_mai_n162_));
  AOI220     m146(.A0(mai_mai_n162_), .A1(mai_mai_n160_), .B0(mai_mai_n113_), .B1(mai_mai_n38_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n164_));
  NO2        m148(.A(mai_mai_n164_), .B(mai_mai_n130_), .Y(mai_mai_n165_));
  NO2        m149(.A(mai_mai_n165_), .B(mai_mai_n163_), .Y(mai_mai_n166_));
  AOI210     m150(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n166_), .Y(mai_mai_n167_));
  OAI210     m151(.A0(mai_mai_n155_), .A1(mai_mai_n50_), .B0(mai_mai_n167_), .Y(mai_mai_n168_));
  NA2        m152(.A(x5), .B(x1), .Y(mai_mai_n169_));
  INV        m153(.A(mai_mai_n169_), .Y(mai_mai_n170_));
  AOI210     m154(.A0(mai_mai_n170_), .A1(mai_mai_n130_), .B0(mai_mai_n36_), .Y(mai_mai_n171_));
  NO2        m155(.A(mai_mai_n62_), .B(mai_mai_n94_), .Y(mai_mai_n172_));
  NAi21      m156(.An(x2), .B(x7), .Y(mai_mai_n173_));
  NO3        m157(.A(mai_mai_n173_), .B(mai_mai_n172_), .C(mai_mai_n48_), .Y(mai_mai_n174_));
  NA2        m158(.A(mai_mai_n174_), .B(mai_mai_n67_), .Y(mai_mai_n175_));
  NAi31      m159(.An(mai_mai_n78_), .B(mai_mai_n38_), .C(mai_mai_n35_), .Y(mai_mai_n176_));
  NA3        m160(.A(mai_mai_n176_), .B(mai_mai_n175_), .C(mai_mai_n171_), .Y(mai_mai_n177_));
  NO4        m161(.A(mai_mai_n177_), .B(mai_mai_n168_), .C(mai_mai_n154_), .D(mai_mai_n151_), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n178_), .B(mai_mai_n150_), .Y(mai_mai_n179_));
  NO2        m163(.A(mai_mai_n146_), .B(mai_mai_n142_), .Y(mai_mai_n180_));
  NA2        m164(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n181_));
  NA2        m165(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n182_));
  NA3        m166(.A(mai_mai_n182_), .B(mai_mai_n181_), .C(mai_mai_n24_), .Y(mai_mai_n183_));
  AN2        m167(.A(mai_mai_n183_), .B(mai_mai_n147_), .Y(mai_mai_n184_));
  NA2        m168(.A(x8), .B(x0), .Y(mai_mai_n185_));
  NO2        m169(.A(mai_mai_n161_), .B(mai_mai_n25_), .Y(mai_mai_n186_));
  NO2        m170(.A(mai_mai_n128_), .B(x4), .Y(mai_mai_n187_));
  NA2        m171(.A(mai_mai_n187_), .B(mai_mai_n186_), .Y(mai_mai_n188_));
  AOI210     m172(.A0(mai_mai_n185_), .A1(mai_mai_n136_), .B0(mai_mai_n188_), .Y(mai_mai_n189_));
  NA2        m173(.A(x2), .B(x0), .Y(mai_mai_n190_));
  NA2        m174(.A(x4), .B(x1), .Y(mai_mai_n191_));
  NAi21      m175(.An(mai_mai_n126_), .B(mai_mai_n191_), .Y(mai_mai_n192_));
  NOi31      m176(.An(mai_mai_n192_), .B(mai_mai_n164_), .C(mai_mai_n190_), .Y(mai_mai_n193_));
  NO4        m177(.A(mai_mai_n193_), .B(mai_mai_n189_), .C(mai_mai_n184_), .D(mai_mai_n180_), .Y(mai_mai_n194_));
  NO2        m178(.A(mai_mai_n194_), .B(mai_mai_n43_), .Y(mai_mai_n195_));
  NO2        m179(.A(mai_mai_n183_), .B(mai_mai_n76_), .Y(mai_mai_n196_));
  INV        m180(.A(mai_mai_n135_), .Y(mai_mai_n197_));
  NO2        m181(.A(mai_mai_n109_), .B(mai_mai_n17_), .Y(mai_mai_n198_));
  AOI210     m182(.A0(mai_mai_n35_), .A1(mai_mai_n94_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  NO3        m183(.A(mai_mai_n199_), .B(mai_mai_n197_), .C(x7), .Y(mai_mai_n200_));
  NA3        m184(.A(mai_mai_n192_), .B(mai_mai_n197_), .C(mai_mai_n42_), .Y(mai_mai_n201_));
  OAI210     m185(.A0(mai_mai_n182_), .A1(mai_mai_n142_), .B0(mai_mai_n201_), .Y(mai_mai_n202_));
  NO3        m186(.A(mai_mai_n202_), .B(mai_mai_n200_), .C(mai_mai_n196_), .Y(mai_mai_n203_));
  NO2        m187(.A(mai_mai_n203_), .B(x3), .Y(mai_mai_n204_));
  NO3        m188(.A(mai_mai_n204_), .B(mai_mai_n195_), .C(mai_mai_n179_), .Y(mai03));
  NO2        m189(.A(mai_mai_n48_), .B(x3), .Y(mai_mai_n206_));
  NO2        m190(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n207_));
  INV        m191(.A(mai_mai_n207_), .Y(mai_mai_n208_));
  NO2        m192(.A(mai_mai_n54_), .B(x1), .Y(mai_mai_n209_));
  OAI210     m193(.A0(mai_mai_n209_), .A1(mai_mai_n25_), .B0(mai_mai_n63_), .Y(mai_mai_n210_));
  OAI220     m194(.A0(mai_mai_n210_), .A1(mai_mai_n17_), .B0(mai_mai_n208_), .B1(mai_mai_n109_), .Y(mai_mai_n211_));
  NA2        m195(.A(mai_mai_n211_), .B(mai_mai_n206_), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n78_), .B(x6), .Y(mai_mai_n213_));
  NA2        m197(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n214_));
  NO2        m198(.A(mai_mai_n214_), .B(x4), .Y(mai_mai_n215_));
  NO2        m199(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n216_));
  AO220      m200(.A0(mai_mai_n216_), .A1(mai_mai_n215_), .B0(mai_mai_n213_), .B1(mai_mai_n55_), .Y(mai_mai_n217_));
  NA2        m201(.A(mai_mai_n217_), .B(mai_mai_n62_), .Y(mai_mai_n218_));
  NA2        m202(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n219_));
  NO2        m203(.A(mai_mai_n219_), .B(mai_mai_n214_), .Y(mai_mai_n220_));
  NA2        m204(.A(x9), .B(mai_mai_n54_), .Y(mai_mai_n221_));
  NA2        m205(.A(mai_mai_n221_), .B(x4), .Y(mai_mai_n222_));
  NA2        m206(.A(mai_mai_n214_), .B(mai_mai_n81_), .Y(mai_mai_n223_));
  AOI210     m207(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n190_), .Y(mai_mai_n224_));
  AOI220     m208(.A0(mai_mai_n224_), .A1(mai_mai_n223_), .B0(mai_mai_n222_), .B1(mai_mai_n220_), .Y(mai_mai_n225_));
  NO3        m209(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n226_));
  NO2        m210(.A(x5), .B(x1), .Y(mai_mai_n227_));
  AOI220     m211(.A0(mai_mai_n227_), .A1(mai_mai_n17_), .B0(mai_mai_n106_), .B1(x5), .Y(mai_mai_n228_));
  NO2        m212(.A(mai_mai_n219_), .B(mai_mai_n181_), .Y(mai_mai_n229_));
  NO3        m213(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n230_));
  NO2        m214(.A(mai_mai_n230_), .B(mai_mai_n229_), .Y(mai_mai_n231_));
  OAI210     m215(.A0(mai_mai_n228_), .A1(mai_mai_n64_), .B0(mai_mai_n231_), .Y(mai_mai_n232_));
  AOI220     m216(.A0(mai_mai_n232_), .A1(mai_mai_n48_), .B0(mai_mai_n226_), .B1(mai_mai_n135_), .Y(mai_mai_n233_));
  NA4        m217(.A(mai_mai_n233_), .B(mai_mai_n225_), .C(mai_mai_n218_), .D(mai_mai_n212_), .Y(mai_mai_n234_));
  NO2        m218(.A(mai_mai_n48_), .B(mai_mai_n43_), .Y(mai_mai_n235_));
  NA2        m219(.A(mai_mai_n235_), .B(mai_mai_n19_), .Y(mai_mai_n236_));
  NO2        m220(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n237_));
  NO2        m221(.A(mai_mai_n237_), .B(x6), .Y(mai_mai_n238_));
  NOi21      m222(.An(mai_mai_n84_), .B(mai_mai_n238_), .Y(mai_mai_n239_));
  NA2        m223(.A(mai_mai_n62_), .B(mai_mai_n94_), .Y(mai_mai_n240_));
  NA3        m224(.A(mai_mai_n240_), .B(mai_mai_n237_), .C(x6), .Y(mai_mai_n241_));
  AOI210     m225(.A0(mai_mai_n241_), .A1(mai_mai_n239_), .B0(mai_mai_n161_), .Y(mai_mai_n242_));
  AO210      m226(.A0(mai_mai_n242_), .A1(mai_mai_n236_), .B0(mai_mai_n186_), .Y(mai_mai_n243_));
  NA2        m227(.A(mai_mai_n43_), .B(mai_mai_n54_), .Y(mai_mai_n244_));
  NA2        m228(.A(mai_mai_n147_), .B(mai_mai_n93_), .Y(mai_mai_n245_));
  NA2        m229(.A(x6), .B(mai_mai_n48_), .Y(mai_mai_n246_));
  OAI210     m230(.A0(mai_mai_n122_), .A1(mai_mai_n79_), .B0(x4), .Y(mai_mai_n247_));
  AOI210     m231(.A0(mai_mai_n247_), .A1(mai_mai_n246_), .B0(mai_mai_n78_), .Y(mai_mai_n248_));
  NO2        m232(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n249_));
  NO2        m233(.A(mai_mai_n169_), .B(mai_mai_n43_), .Y(mai_mai_n250_));
  NA2        m234(.A(mai_mai_n250_), .B(mai_mai_n249_), .Y(mai_mai_n251_));
  NA2        m235(.A(mai_mai_n207_), .B(mai_mai_n140_), .Y(mai_mai_n252_));
  NA3        m236(.A(mai_mai_n219_), .B(mai_mai_n135_), .C(x6), .Y(mai_mai_n253_));
  OAI210     m237(.A0(mai_mai_n94_), .A1(mai_mai_n36_), .B0(mai_mai_n67_), .Y(mai_mai_n254_));
  NA4        m238(.A(mai_mai_n254_), .B(mai_mai_n253_), .C(mai_mai_n252_), .D(mai_mai_n251_), .Y(mai_mai_n255_));
  OAI210     m239(.A0(mai_mai_n255_), .A1(mai_mai_n248_), .B0(x2), .Y(mai_mai_n256_));
  NA3        m240(.A(mai_mai_n256_), .B(mai_mai_n245_), .C(mai_mai_n243_), .Y(mai_mai_n257_));
  AOI210     m241(.A0(mai_mai_n234_), .A1(x8), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  NO2        m242(.A(mai_mai_n94_), .B(x3), .Y(mai_mai_n259_));
  NA2        m243(.A(mai_mai_n259_), .B(mai_mai_n215_), .Y(mai_mai_n260_));
  NO3        m244(.A(mai_mai_n92_), .B(mai_mai_n79_), .C(mai_mai_n25_), .Y(mai_mai_n261_));
  AOI210     m245(.A0(mai_mai_n238_), .A1(mai_mai_n164_), .B0(mai_mai_n261_), .Y(mai_mai_n262_));
  AOI210     m246(.A0(mai_mai_n262_), .A1(mai_mai_n260_), .B0(x2), .Y(mai_mai_n263_));
  NO2        m247(.A(x4), .B(mai_mai_n54_), .Y(mai_mai_n264_));
  AOI220     m248(.A0(mai_mai_n215_), .A1(mai_mai_n198_), .B0(mai_mai_n264_), .B1(mai_mai_n67_), .Y(mai_mai_n265_));
  NA2        m249(.A(mai_mai_n62_), .B(x6), .Y(mai_mai_n266_));
  NA2        m250(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n267_));
  NO2        m251(.A(mai_mai_n267_), .B(mai_mai_n25_), .Y(mai_mai_n268_));
  NA2        m252(.A(mai_mai_n268_), .B(mai_mai_n126_), .Y(mai_mai_n269_));
  NA2        m253(.A(mai_mai_n219_), .B(x6), .Y(mai_mai_n270_));
  NO2        m254(.A(mai_mai_n219_), .B(x6), .Y(mai_mai_n271_));
  NAi21      m255(.An(mai_mai_n172_), .B(mai_mai_n271_), .Y(mai_mai_n272_));
  NA3        m256(.A(mai_mai_n272_), .B(mai_mai_n270_), .C(mai_mai_n152_), .Y(mai_mai_n273_));
  NA4        m257(.A(mai_mai_n273_), .B(mai_mai_n269_), .C(mai_mai_n265_), .D(mai_mai_n161_), .Y(mai_mai_n274_));
  NA2        m258(.A(mai_mai_n207_), .B(mai_mai_n237_), .Y(mai_mai_n275_));
  NAi21      m259(.An(x1), .B(x4), .Y(mai_mai_n276_));
  AOI210     m260(.A0(x3), .A1(x2), .B0(mai_mai_n48_), .Y(mai_mai_n277_));
  OAI210     m261(.A0(mai_mai_n146_), .A1(x3), .B0(mai_mai_n277_), .Y(mai_mai_n278_));
  NA2        m262(.A(mai_mai_n278_), .B(mai_mai_n276_), .Y(mai_mai_n279_));
  NA2        m263(.A(mai_mai_n279_), .B(mai_mai_n275_), .Y(mai_mai_n280_));
  NA2        m264(.A(mai_mai_n62_), .B(x2), .Y(mai_mai_n281_));
  NO2        m265(.A(mai_mai_n281_), .B(mai_mai_n275_), .Y(mai_mai_n282_));
  NO3        m266(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n283_));
  NA2        m267(.A(mai_mai_n109_), .B(mai_mai_n25_), .Y(mai_mai_n284_));
  NA2        m268(.A(x6), .B(x2), .Y(mai_mai_n285_));
  NO2        m269(.A(mai_mai_n285_), .B(mai_mai_n181_), .Y(mai_mai_n286_));
  AOI210     m270(.A0(mai_mai_n284_), .A1(mai_mai_n283_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  OAI220     m271(.A0(mai_mai_n287_), .A1(mai_mai_n43_), .B0(mai_mai_n187_), .B1(mai_mai_n46_), .Y(mai_mai_n288_));
  OAI210     m272(.A0(mai_mai_n288_), .A1(mai_mai_n282_), .B0(mai_mai_n280_), .Y(mai_mai_n289_));
  NA2        m273(.A(x9), .B(mai_mai_n43_), .Y(mai_mai_n290_));
  NO2        m274(.A(mai_mai_n290_), .B(mai_mai_n214_), .Y(mai_mai_n291_));
  OR3        m275(.A(mai_mai_n291_), .B(mai_mai_n213_), .C(mai_mai_n156_), .Y(mai_mai_n292_));
  NA2        m276(.A(x4), .B(x0), .Y(mai_mai_n293_));
  NO3        m277(.A(mai_mai_n73_), .B(mai_mai_n293_), .C(x6), .Y(mai_mai_n294_));
  AOI210     m278(.A0(mai_mai_n292_), .A1(mai_mai_n42_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  AOI210     m279(.A0(mai_mai_n295_), .A1(mai_mai_n289_), .B0(x8), .Y(mai_mai_n296_));
  INV        m280(.A(mai_mai_n266_), .Y(mai_mai_n297_));
  NA2        m281(.A(mai_mai_n227_), .B(mai_mai_n297_), .Y(mai_mai_n298_));
  INV        m282(.A(mai_mai_n185_), .Y(mai_mai_n299_));
  OAI210     m283(.A0(mai_mai_n299_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n300_));
  AOI210     m284(.A0(mai_mai_n300_), .A1(mai_mai_n298_), .B0(mai_mai_n244_), .Y(mai_mai_n301_));
  NO4        m285(.A(mai_mai_n301_), .B(mai_mai_n296_), .C(mai_mai_n274_), .D(mai_mai_n263_), .Y(mai_mai_n302_));
  NO2        m286(.A(mai_mai_n172_), .B(x1), .Y(mai_mai_n303_));
  NO3        m287(.A(mai_mai_n303_), .B(x3), .C(mai_mai_n36_), .Y(mai_mai_n304_));
  OAI210     m288(.A0(mai_mai_n304_), .A1(mai_mai_n271_), .B0(x2), .Y(mai_mai_n305_));
  OAI210     m289(.A0(mai_mai_n299_), .A1(x6), .B0(mai_mai_n44_), .Y(mai_mai_n306_));
  AOI210     m290(.A0(mai_mai_n306_), .A1(mai_mai_n305_), .B0(mai_mai_n197_), .Y(mai_mai_n307_));
  NOi21      m291(.An(mai_mai_n285_), .B(mai_mai_n17_), .Y(mai_mai_n308_));
  NA3        m292(.A(mai_mai_n308_), .B(mai_mai_n227_), .C(mai_mai_n40_), .Y(mai_mai_n309_));
  AOI210     m293(.A0(mai_mai_n36_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n170_), .C(mai_mai_n32_), .Y(mai_mai_n311_));
  NA2        m295(.A(x3), .B(x2), .Y(mai_mai_n312_));
  AOI220     m296(.A0(mai_mai_n312_), .A1(mai_mai_n244_), .B0(mai_mai_n311_), .B1(mai_mai_n309_), .Y(mai_mai_n313_));
  NAi21      m297(.An(x4), .B(x0), .Y(mai_mai_n314_));
  NO3        m298(.A(mai_mai_n314_), .B(mai_mai_n44_), .C(x2), .Y(mai_mai_n315_));
  OAI210     m299(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n315_), .Y(mai_mai_n316_));
  OAI220     m300(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n317_));
  NO2        m301(.A(x9), .B(x8), .Y(mai_mai_n318_));
  NA3        m302(.A(mai_mai_n318_), .B(mai_mai_n36_), .C(mai_mai_n54_), .Y(mai_mai_n319_));
  OAI210     m303(.A0(mai_mai_n310_), .A1(mai_mai_n308_), .B0(mai_mai_n319_), .Y(mai_mai_n320_));
  AOI220     m304(.A0(mai_mai_n320_), .A1(mai_mai_n82_), .B0(mai_mai_n317_), .B1(mai_mai_n31_), .Y(mai_mai_n321_));
  AOI210     m305(.A0(mai_mai_n321_), .A1(mai_mai_n316_), .B0(mai_mai_n25_), .Y(mai_mai_n322_));
  NA3        m306(.A(mai_mai_n36_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n323_));
  OAI210     m307(.A0(mai_mai_n310_), .A1(mai_mai_n308_), .B0(mai_mai_n323_), .Y(mai_mai_n324_));
  INV        m308(.A(mai_mai_n229_), .Y(mai_mai_n325_));
  NA2        m309(.A(mai_mai_n36_), .B(mai_mai_n43_), .Y(mai_mai_n326_));
  OR2        m310(.A(mai_mai_n326_), .B(mai_mai_n293_), .Y(mai_mai_n327_));
  OAI220     m311(.A0(mai_mai_n327_), .A1(mai_mai_n169_), .B0(mai_mai_n246_), .B1(mai_mai_n325_), .Y(mai_mai_n328_));
  AO210      m312(.A0(mai_mai_n324_), .A1(mai_mai_n156_), .B0(mai_mai_n328_), .Y(mai_mai_n329_));
  NO4        m313(.A(mai_mai_n329_), .B(mai_mai_n322_), .C(mai_mai_n313_), .D(mai_mai_n307_), .Y(mai_mai_n330_));
  OAI210     m314(.A0(mai_mai_n302_), .A1(mai_mai_n258_), .B0(mai_mai_n330_), .Y(mai04));
  OAI210     m315(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n332_));
  NA3        m316(.A(mai_mai_n332_), .B(mai_mai_n283_), .C(mai_mai_n85_), .Y(mai_mai_n333_));
  NO2        m317(.A(x2), .B(x1), .Y(mai_mai_n334_));
  OAI210     m318(.A0(mai_mai_n267_), .A1(mai_mai_n334_), .B0(mai_mai_n36_), .Y(mai_mai_n335_));
  NO2        m319(.A(mai_mai_n334_), .B(mai_mai_n314_), .Y(mai_mai_n336_));
  AOI210     m320(.A0(mai_mai_n62_), .A1(x4), .B0(mai_mai_n115_), .Y(mai_mai_n337_));
  OAI210     m321(.A0(mai_mai_n337_), .A1(mai_mai_n336_), .B0(mai_mai_n259_), .Y(mai_mai_n338_));
  NO2        m322(.A(mai_mai_n281_), .B(mai_mai_n92_), .Y(mai_mai_n339_));
  NO2        m323(.A(mai_mai_n339_), .B(mai_mai_n36_), .Y(mai_mai_n340_));
  NO2        m324(.A(mai_mai_n312_), .B(mai_mai_n216_), .Y(mai_mai_n341_));
  NA2        m325(.A(x9), .B(x0), .Y(mai_mai_n342_));
  AOI210     m326(.A0(mai_mai_n92_), .A1(mai_mai_n76_), .B0(mai_mai_n342_), .Y(mai_mai_n343_));
  OAI210     m327(.A0(mai_mai_n343_), .A1(mai_mai_n341_), .B0(mai_mai_n94_), .Y(mai_mai_n344_));
  NA3        m328(.A(mai_mai_n344_), .B(mai_mai_n340_), .C(mai_mai_n338_), .Y(mai_mai_n345_));
  NA2        m329(.A(mai_mai_n345_), .B(mai_mai_n335_), .Y(mai_mai_n346_));
  NO2        m330(.A(mai_mai_n221_), .B(mai_mai_n116_), .Y(mai_mai_n347_));
  NO3        m331(.A(mai_mai_n266_), .B(mai_mai_n123_), .C(mai_mai_n18_), .Y(mai_mai_n348_));
  NO2        m332(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  OAI210     m333(.A0(mai_mai_n121_), .A1(mai_mai_n109_), .B0(mai_mai_n185_), .Y(mai_mai_n350_));
  NA3        m334(.A(mai_mai_n350_), .B(x6), .C(x3), .Y(mai_mai_n351_));
  NOi21      m335(.An(mai_mai_n158_), .B(mai_mai_n136_), .Y(mai_mai_n352_));
  AOI210     m336(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n353_));
  OAI220     m337(.A0(mai_mai_n353_), .A1(mai_mai_n326_), .B0(mai_mai_n281_), .B1(mai_mai_n323_), .Y(mai_mai_n354_));
  AOI210     m338(.A0(mai_mai_n352_), .A1(mai_mai_n63_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NA2        m339(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n109_), .A1(mai_mai_n17_), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  NA2        m341(.A(mai_mai_n357_), .B(mai_mai_n79_), .Y(mai_mai_n358_));
  NA4        m342(.A(mai_mai_n358_), .B(mai_mai_n355_), .C(mai_mai_n351_), .D(mai_mai_n349_), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n114_), .A1(x3), .B0(mai_mai_n315_), .Y(mai_mai_n360_));
  NA3        m344(.A(mai_mai_n240_), .B(mai_mai_n226_), .C(mai_mai_n84_), .Y(mai_mai_n361_));
  NA3        m345(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n161_), .Y(mai_mai_n362_));
  AOI210     m346(.A0(mai_mai_n359_), .A1(x4), .B0(mai_mai_n362_), .Y(mai_mai_n363_));
  NA3        m347(.A(mai_mai_n336_), .B(mai_mai_n221_), .C(mai_mai_n94_), .Y(mai_mai_n364_));
  NOi21      m348(.An(x4), .B(x0), .Y(mai_mai_n365_));
  XO2        m349(.A(x4), .B(x0), .Y(mai_mai_n366_));
  OAI210     m350(.A0(mai_mai_n366_), .A1(mai_mai_n120_), .B0(mai_mai_n276_), .Y(mai_mai_n367_));
  AOI220     m351(.A0(mai_mai_n367_), .A1(x8), .B0(mai_mai_n365_), .B1(mai_mai_n95_), .Y(mai_mai_n368_));
  AOI210     m352(.A0(mai_mai_n368_), .A1(mai_mai_n364_), .B0(x3), .Y(mai_mai_n369_));
  INV        m353(.A(mai_mai_n95_), .Y(mai_mai_n370_));
  NO2        m354(.A(mai_mai_n94_), .B(x4), .Y(mai_mai_n371_));
  AOI220     m355(.A0(mai_mai_n371_), .A1(mai_mai_n44_), .B0(mai_mai_n130_), .B1(mai_mai_n370_), .Y(mai_mai_n372_));
  NO3        m356(.A(mai_mai_n366_), .B(mai_mai_n172_), .C(x2), .Y(mai_mai_n373_));
  INV        m357(.A(mai_mai_n373_), .Y(mai_mai_n374_));
  NA4        m358(.A(mai_mai_n374_), .B(mai_mai_n372_), .C(mai_mai_n236_), .D(x6), .Y(mai_mai_n375_));
  OAI220     m359(.A0(mai_mai_n314_), .A1(mai_mai_n92_), .B0(mai_mai_n190_), .B1(mai_mai_n94_), .Y(mai_mai_n376_));
  NO2        m360(.A(mai_mai_n43_), .B(x0), .Y(mai_mai_n377_));
  NA2        m361(.A(mai_mai_n376_), .B(mai_mai_n61_), .Y(mai_mai_n378_));
  NO2        m362(.A(mai_mai_n158_), .B(mai_mai_n81_), .Y(mai_mai_n379_));
  NO2        m363(.A(mai_mai_n35_), .B(x2), .Y(mai_mai_n380_));
  NOi21      m364(.An(mai_mai_n126_), .B(mai_mai_n27_), .Y(mai_mai_n381_));
  AOI210     m365(.A0(mai_mai_n380_), .A1(mai_mai_n379_), .B0(mai_mai_n381_), .Y(mai_mai_n382_));
  OAI210     m366(.A0(mai_mai_n378_), .A1(mai_mai_n62_), .B0(mai_mai_n382_), .Y(mai_mai_n383_));
  OAI220     m367(.A0(mai_mai_n383_), .A1(x6), .B0(mai_mai_n375_), .B1(mai_mai_n369_), .Y(mai_mai_n384_));
  OAI210     m368(.A0(mai_mai_n63_), .A1(mai_mai_n48_), .B0(mai_mai_n42_), .Y(mai_mai_n385_));
  OAI210     m369(.A0(mai_mai_n385_), .A1(mai_mai_n94_), .B0(mai_mai_n327_), .Y(mai_mai_n386_));
  AOI210     m370(.A0(mai_mai_n386_), .A1(mai_mai_n18_), .B0(mai_mai_n161_), .Y(mai_mai_n387_));
  AO220      m371(.A0(mai_mai_n387_), .A1(mai_mai_n384_), .B0(mai_mai_n363_), .B1(mai_mai_n346_), .Y(mai_mai_n388_));
  NA2        m372(.A(mai_mai_n380_), .B(x6), .Y(mai_mai_n389_));
  AOI210     m373(.A0(x6), .A1(x1), .B0(mai_mai_n160_), .Y(mai_mai_n390_));
  NA2        m374(.A(mai_mai_n371_), .B(x0), .Y(mai_mai_n391_));
  NA2        m375(.A(mai_mai_n84_), .B(x6), .Y(mai_mai_n392_));
  OAI210     m376(.A0(mai_mai_n391_), .A1(mai_mai_n390_), .B0(mai_mai_n392_), .Y(mai_mai_n393_));
  AOI220     m377(.A0(mai_mai_n393_), .A1(mai_mai_n389_), .B0(mai_mai_n230_), .B1(mai_mai_n49_), .Y(mai_mai_n394_));
  NA3        m378(.A(mai_mai_n394_), .B(mai_mai_n388_), .C(mai_mai_n333_), .Y(mai_mai_n395_));
  AOI210     m379(.A0(mai_mai_n209_), .A1(x8), .B0(mai_mai_n114_), .Y(mai_mai_n396_));
  NA2        m380(.A(mai_mai_n396_), .B(mai_mai_n356_), .Y(mai_mai_n397_));
  NA3        m381(.A(mai_mai_n397_), .B(mai_mai_n206_), .C(mai_mai_n161_), .Y(mai_mai_n398_));
  OAI210     m382(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n244_), .Y(mai_mai_n399_));
  AO220      m383(.A0(mai_mai_n399_), .A1(mai_mai_n157_), .B0(mai_mai_n113_), .B1(x4), .Y(mai_mai_n400_));
  NA3        m384(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n401_));
  NA2        m385(.A(mai_mai_n235_), .B(x0), .Y(mai_mai_n402_));
  OAI220     m386(.A0(mai_mai_n402_), .A1(mai_mai_n221_), .B0(mai_mai_n401_), .B1(mai_mai_n370_), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n400_), .A1(mai_mai_n122_), .B0(mai_mai_n403_), .Y(mai_mai_n404_));
  AOI210     m388(.A0(mai_mai_n404_), .A1(mai_mai_n398_), .B0(mai_mai_n25_), .Y(mai_mai_n405_));
  NA3        m389(.A(mai_mai_n124_), .B(mai_mai_n235_), .C(x0), .Y(mai_mai_n406_));
  NAi31      m390(.An(mai_mai_n50_), .B(mai_mai_n303_), .C(mai_mai_n186_), .Y(mai_mai_n407_));
  NA2        m391(.A(mai_mai_n407_), .B(mai_mai_n406_), .Y(mai_mai_n408_));
  OAI210     m392(.A0(mai_mai_n408_), .A1(mai_mai_n405_), .B0(x6), .Y(mai_mai_n409_));
  OAI210     m393(.A0(mai_mai_n172_), .A1(mai_mai_n48_), .B0(mai_mai_n141_), .Y(mai_mai_n410_));
  NA3        m394(.A(mai_mai_n55_), .B(mai_mai_n38_), .C(mai_mai_n31_), .Y(mai_mai_n411_));
  AOI220     m395(.A0(mai_mai_n411_), .A1(mai_mai_n410_), .B0(mai_mai_n40_), .B1(mai_mai_n32_), .Y(mai_mai_n412_));
  NO2        m396(.A(mai_mai_n161_), .B(x0), .Y(mai_mai_n413_));
  AOI220     m397(.A0(mai_mai_n413_), .A1(mai_mai_n235_), .B0(mai_mai_n206_), .B1(mai_mai_n161_), .Y(mai_mai_n414_));
  AOI210     m398(.A0(mai_mai_n132_), .A1(mai_mai_n264_), .B0(x1), .Y(mai_mai_n415_));
  OAI210     m399(.A0(mai_mai_n414_), .A1(x8), .B0(mai_mai_n415_), .Y(mai_mai_n416_));
  NAi31      m400(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n417_));
  OAI210     m401(.A0(mai_mai_n417_), .A1(x4), .B0(mai_mai_n173_), .Y(mai_mai_n418_));
  NA3        m402(.A(mai_mai_n418_), .B(mai_mai_n155_), .C(x9), .Y(mai_mai_n419_));
  NO4        m403(.A(mai_mai_n131_), .B(mai_mai_n314_), .C(x9), .D(x2), .Y(mai_mai_n420_));
  NOi21      m404(.An(mai_mai_n129_), .B(mai_mai_n190_), .Y(mai_mai_n421_));
  NO3        m405(.A(mai_mai_n421_), .B(mai_mai_n420_), .C(mai_mai_n18_), .Y(mai_mai_n422_));
  NO3        m406(.A(x9), .B(mai_mai_n161_), .C(x0), .Y(mai_mai_n423_));
  AOI220     m407(.A0(mai_mai_n423_), .A1(mai_mai_n259_), .B0(mai_mai_n379_), .B1(mai_mai_n161_), .Y(mai_mai_n424_));
  NA4        m408(.A(mai_mai_n424_), .B(mai_mai_n422_), .C(mai_mai_n419_), .D(mai_mai_n50_), .Y(mai_mai_n425_));
  OAI210     m409(.A0(mai_mai_n416_), .A1(mai_mai_n412_), .B0(mai_mai_n425_), .Y(mai_mai_n426_));
  NOi31      m410(.An(mai_mai_n413_), .B(mai_mai_n32_), .C(x8), .Y(mai_mai_n427_));
  AOI210     m411(.A0(mai_mai_n38_), .A1(x9), .B0(mai_mai_n139_), .Y(mai_mai_n428_));
  NO3        m412(.A(mai_mai_n428_), .B(mai_mai_n129_), .C(mai_mai_n43_), .Y(mai_mai_n429_));
  NOi31      m413(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n430_));
  AOI220     m414(.A0(mai_mai_n430_), .A1(mai_mai_n365_), .B0(mai_mai_n130_), .B1(x3), .Y(mai_mai_n431_));
  AOI210     m415(.A0(mai_mai_n276_), .A1(mai_mai_n60_), .B0(mai_mai_n128_), .Y(mai_mai_n432_));
  OAI210     m416(.A0(mai_mai_n432_), .A1(x3), .B0(mai_mai_n431_), .Y(mai_mai_n433_));
  NO3        m417(.A(mai_mai_n433_), .B(mai_mai_n429_), .C(x2), .Y(mai_mai_n434_));
  OAI220     m418(.A0(mai_mai_n366_), .A1(mai_mai_n318_), .B0(mai_mai_n314_), .B1(mai_mai_n43_), .Y(mai_mai_n435_));
  AOI210     m419(.A0(x9), .A1(mai_mai_n48_), .B0(mai_mai_n401_), .Y(mai_mai_n436_));
  AOI220     m420(.A0(mai_mai_n436_), .A1(mai_mai_n94_), .B0(mai_mai_n435_), .B1(mai_mai_n161_), .Y(mai_mai_n437_));
  NO2        m421(.A(mai_mai_n437_), .B(mai_mai_n54_), .Y(mai_mai_n438_));
  NO3        m422(.A(mai_mai_n438_), .B(mai_mai_n434_), .C(mai_mai_n427_), .Y(mai_mai_n439_));
  AOI210     m423(.A0(mai_mai_n439_), .A1(mai_mai_n426_), .B0(mai_mai_n25_), .Y(mai_mai_n440_));
  NA4        m424(.A(mai_mai_n31_), .B(mai_mai_n94_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n441_));
  NO3        m425(.A(mai_mai_n68_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n442_));
  NA2        m426(.A(mai_mai_n442_), .B(mai_mai_n277_), .Y(mai_mai_n443_));
  NO2        m427(.A(mai_mai_n443_), .B(mai_mai_n106_), .Y(mai_mai_n444_));
  NO3        m428(.A(mai_mai_n281_), .B(mai_mai_n185_), .C(mai_mai_n40_), .Y(mai_mai_n445_));
  OAI210     m429(.A0(mai_mai_n445_), .A1(mai_mai_n444_), .B0(x7), .Y(mai_mai_n446_));
  NA2        m430(.A(mai_mai_n240_), .B(x7), .Y(mai_mai_n447_));
  NA3        m431(.A(mai_mai_n447_), .B(mai_mai_n160_), .C(mai_mai_n140_), .Y(mai_mai_n448_));
  NA3        m432(.A(mai_mai_n448_), .B(mai_mai_n446_), .C(mai_mai_n441_), .Y(mai_mai_n449_));
  OAI210     m433(.A0(mai_mai_n449_), .A1(mai_mai_n440_), .B0(mai_mai_n36_), .Y(mai_mai_n450_));
  NO2        m434(.A(mai_mai_n423_), .B(mai_mai_n216_), .Y(mai_mai_n451_));
  NO4        m435(.A(mai_mai_n451_), .B(mai_mai_n78_), .C(x4), .D(mai_mai_n54_), .Y(mai_mai_n452_));
  NA2        m436(.A(mai_mai_n267_), .B(mai_mai_n21_), .Y(mai_mai_n453_));
  NO2        m437(.A(mai_mai_n169_), .B(mai_mai_n141_), .Y(mai_mai_n454_));
  NA2        m438(.A(mai_mai_n454_), .B(mai_mai_n453_), .Y(mai_mai_n455_));
  AOI210     m439(.A0(mai_mai_n455_), .A1(mai_mai_n176_), .B0(mai_mai_n28_), .Y(mai_mai_n456_));
  AOI220     m440(.A0(mai_mai_n377_), .A1(mai_mai_n94_), .B0(mai_mai_n158_), .B1(mai_mai_n209_), .Y(mai_mai_n457_));
  NA3        m441(.A(mai_mai_n457_), .B(mai_mai_n417_), .C(mai_mai_n92_), .Y(mai_mai_n458_));
  NA2        m442(.A(mai_mai_n458_), .B(mai_mai_n186_), .Y(mai_mai_n459_));
  OAI220     m443(.A0(mai_mai_n290_), .A1(mai_mai_n69_), .B0(mai_mai_n169_), .B1(mai_mai_n43_), .Y(mai_mai_n460_));
  NA2        m444(.A(x3), .B(mai_mai_n54_), .Y(mai_mai_n461_));
  AOI210     m445(.A0(mai_mai_n173_), .A1(mai_mai_n27_), .B0(mai_mai_n73_), .Y(mai_mai_n462_));
  OAI210     m446(.A0(mai_mai_n157_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n463_));
  NO3        m447(.A(mai_mai_n430_), .B(x3), .C(mai_mai_n54_), .Y(mai_mai_n464_));
  AOI210     m448(.A0(mai_mai_n464_), .A1(mai_mai_n463_), .B0(mai_mai_n462_), .Y(mai_mai_n465_));
  OAI210     m449(.A0(mai_mai_n162_), .A1(mai_mai_n461_), .B0(mai_mai_n465_), .Y(mai_mai_n466_));
  AOI220     m450(.A0(mai_mai_n466_), .A1(x0), .B0(mai_mai_n460_), .B1(mai_mai_n141_), .Y(mai_mai_n467_));
  AOI210     m451(.A0(mai_mai_n467_), .A1(mai_mai_n459_), .B0(mai_mai_n246_), .Y(mai_mai_n468_));
  NA2        m452(.A(x9), .B(x5), .Y(mai_mai_n469_));
  NO4        m453(.A(mai_mai_n109_), .B(mai_mai_n469_), .C(mai_mai_n60_), .D(mai_mai_n32_), .Y(mai_mai_n470_));
  NO4        m454(.A(mai_mai_n470_), .B(mai_mai_n468_), .C(mai_mai_n456_), .D(mai_mai_n452_), .Y(mai_mai_n471_));
  NA3        m455(.A(mai_mai_n471_), .B(mai_mai_n450_), .C(mai_mai_n409_), .Y(mai_mai_n472_));
  AOI210     m456(.A0(mai_mai_n395_), .A1(mai_mai_n25_), .B0(mai_mai_n472_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  INV        u012(.A(men_men_n24_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  OA210      u015(.A0(men_men_n31_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n32_));
  NOi31      u016(.An(men_men_n23_), .B(men_men_n32_), .C(men_men_n29_), .Y(men00));
  NO2        u017(.A(x1), .B(x0), .Y(men_men_n34_));
  INV        u018(.A(x6), .Y(men_men_n35_));
  NO2        u019(.A(men_men_n35_), .B(men_men_n25_), .Y(men_men_n36_));
  AN2        u020(.A(x8), .B(x7), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  NO2        u022(.A(men_men_n23_), .B(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n36_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n50_));
  AOI220     u034(.A0(men_men_n50_), .A1(men_men_n34_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n35_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO3        u046(.A(men_men_n62_), .B(men_men_n59_), .C(men_men_n58_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  NO2        u051(.A(men_men_n67_), .B(x1), .Y(men_men_n68_));
  OA210      u052(.A0(men_men_n68_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n42_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n70_), .Y(men_men_n71_));
  NAi31      u055(.An(x1), .B(x9), .C(x5), .Y(men_men_n72_));
  OAI220     u056(.A0(men_men_n72_), .A1(men_men_n41_), .B0(men_men_n71_), .B1(men_men_n69_), .Y(men_men_n73_));
  OAI210     u057(.A0(men_men_n73_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n46_), .B(x2), .Y(men_men_n75_));
  OAI210     u059(.A0(men_men_n75_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n76_));
  NA2        u060(.A(x5), .B(x3), .Y(men_men_n77_));
  NO2        u061(.A(x8), .B(x6), .Y(men_men_n78_));
  NO4        u062(.A(men_men_n78_), .B(men_men_n77_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n79_));
  NAi21      u063(.An(x4), .B(x3), .Y(men_men_n80_));
  INV        u064(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(men_men_n22_), .Y(men_men_n82_));
  NO2        u066(.A(x4), .B(x2), .Y(men_men_n83_));
  NO2        u067(.A(men_men_n83_), .B(x3), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n84_), .B(men_men_n82_), .C(men_men_n18_), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n79_), .C(men_men_n76_), .Y(men_men_n86_));
  NO4        u070(.A(men_men_n21_), .B(x6), .C(men_men_n41_), .D(x1), .Y(men_men_n87_));
  NA2        u071(.A(men_men_n60_), .B(men_men_n46_), .Y(men_men_n88_));
  INV        u072(.A(men_men_n88_), .Y(men_men_n89_));
  OAI210     u073(.A0(men_men_n87_), .A1(men_men_n65_), .B0(men_men_n89_), .Y(men_men_n90_));
  NA2        u074(.A(x3), .B(men_men_n18_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n25_), .Y(men_men_n92_));
  INV        u076(.A(x8), .Y(men_men_n93_));
  NA2        u077(.A(x2), .B(x1), .Y(men_men_n94_));
  NO2        u078(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n92_), .Y(men_men_n96_));
  NO2        u080(.A(men_men_n96_), .B(men_men_n26_), .Y(men_men_n97_));
  AOI210     u081(.A0(men_men_n54_), .A1(men_men_n25_), .B0(men_men_n52_), .Y(men_men_n98_));
  OAI210     u082(.A0(men_men_n43_), .A1(men_men_n36_), .B0(men_men_n46_), .Y(men_men_n99_));
  NO3        u083(.A(men_men_n99_), .B(men_men_n98_), .C(men_men_n97_), .Y(men_men_n100_));
  NA2        u084(.A(x4), .B(men_men_n41_), .Y(men_men_n101_));
  NO2        u085(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n102_));
  NA2        u086(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n103_));
  AOI210     u087(.A0(men_men_n101_), .A1(men_men_n50_), .B0(men_men_n103_), .Y(men_men_n104_));
  NO2        u088(.A(x3), .B(x2), .Y(men_men_n105_));
  NA3        u089(.A(men_men_n105_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n106_));
  AOI210     u090(.A0(x8), .A1(x6), .B0(men_men_n106_), .Y(men_men_n107_));
  NA2        u091(.A(men_men_n52_), .B(x1), .Y(men_men_n108_));
  OAI210     u092(.A0(men_men_n108_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n109_));
  NO4        u093(.A(men_men_n109_), .B(men_men_n107_), .C(men_men_n104_), .D(men_men_n100_), .Y(men_men_n110_));
  AO220      u094(.A0(men_men_n110_), .A1(men_men_n90_), .B0(men_men_n86_), .B1(men_men_n74_), .Y(men02));
  NO2        u095(.A(x3), .B(men_men_n52_), .Y(men_men_n112_));
  NO2        u096(.A(x8), .B(men_men_n18_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n114_));
  NA2        u098(.A(men_men_n41_), .B(x0), .Y(men_men_n115_));
  OAI210     u099(.A0(men_men_n88_), .A1(men_men_n114_), .B0(men_men_n115_), .Y(men_men_n116_));
  AOI220     u100(.A0(men_men_n116_), .A1(men_men_n113_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n117_));
  NO3        u101(.A(men_men_n117_), .B(x7), .C(x5), .Y(men_men_n118_));
  NA2        u102(.A(x9), .B(x2), .Y(men_men_n119_));
  OR2        u103(.A(x8), .B(x0), .Y(men_men_n120_));
  INV        u104(.A(men_men_n120_), .Y(men_men_n121_));
  NAi21      u105(.An(x2), .B(x8), .Y(men_men_n122_));
  INV        u106(.A(men_men_n122_), .Y(men_men_n123_));
  OAI220     u107(.A0(men_men_n123_), .A1(men_men_n121_), .B0(men_men_n119_), .B1(x7), .Y(men_men_n124_));
  NO2        u108(.A(x4), .B(x1), .Y(men_men_n125_));
  NA3        u109(.A(men_men_n125_), .B(men_men_n124_), .C(men_men_n58_), .Y(men_men_n126_));
  NOi21      u110(.An(x0), .B(x1), .Y(men_men_n127_));
  NO3        u111(.A(x9), .B(x8), .C(x7), .Y(men_men_n128_));
  NOi21      u112(.An(x0), .B(x4), .Y(men_men_n129_));
  NAi21      u113(.An(x8), .B(x7), .Y(men_men_n130_));
  NO2        u114(.A(men_men_n130_), .B(men_men_n60_), .Y(men_men_n131_));
  NO2        u115(.A(men_men_n126_), .B(men_men_n77_), .Y(men_men_n132_));
  NO2        u116(.A(x5), .B(men_men_n46_), .Y(men_men_n133_));
  NA2        u117(.A(x2), .B(men_men_n18_), .Y(men_men_n134_));
  AOI210     u118(.A0(men_men_n134_), .A1(men_men_n108_), .B0(men_men_n115_), .Y(men_men_n135_));
  OAI210     u119(.A0(men_men_n135_), .A1(men_men_n34_), .B0(men_men_n133_), .Y(men_men_n136_));
  NAi21      u120(.An(x0), .B(x4), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x1), .Y(men_men_n138_));
  NO2        u122(.A(x7), .B(x0), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n83_), .B(men_men_n102_), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n140_), .B(x3), .Y(men_men_n141_));
  OAI210     u125(.A0(men_men_n139_), .A1(men_men_n138_), .B0(men_men_n141_), .Y(men_men_n142_));
  NO2        u126(.A(men_men_n21_), .B(men_men_n41_), .Y(men_men_n143_));
  NA2        u127(.A(x5), .B(x0), .Y(men_men_n144_));
  NO2        u128(.A(men_men_n46_), .B(x2), .Y(men_men_n145_));
  NA3        u129(.A(men_men_n145_), .B(men_men_n144_), .C(men_men_n143_), .Y(men_men_n146_));
  NA4        u130(.A(men_men_n146_), .B(men_men_n142_), .C(men_men_n136_), .D(men_men_n35_), .Y(men_men_n147_));
  NO3        u131(.A(men_men_n147_), .B(men_men_n132_), .C(men_men_n118_), .Y(men_men_n148_));
  NO3        u132(.A(men_men_n77_), .B(men_men_n75_), .C(men_men_n24_), .Y(men_men_n149_));
  NO2        u133(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n150_));
  AOI220     u134(.A0(men_men_n127_), .A1(men_men_n150_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n151_));
  NO3        u135(.A(men_men_n151_), .B(men_men_n58_), .C(men_men_n60_), .Y(men_men_n152_));
  NA2        u136(.A(x7), .B(x3), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n101_), .B(x5), .Y(men_men_n154_));
  NO2        u138(.A(x9), .B(x7), .Y(men_men_n155_));
  NOi21      u139(.An(x8), .B(x0), .Y(men_men_n156_));
  OA210      u140(.A0(men_men_n155_), .A1(x1), .B0(men_men_n156_), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n41_), .B(x2), .Y(men_men_n158_));
  INV        u142(.A(x7), .Y(men_men_n159_));
  NA2        u143(.A(men_men_n159_), .B(men_men_n18_), .Y(men_men_n160_));
  AOI220     u144(.A0(men_men_n160_), .A1(men_men_n158_), .B0(men_men_n112_), .B1(men_men_n37_), .Y(men_men_n161_));
  NO2        u145(.A(men_men_n25_), .B(x4), .Y(men_men_n162_));
  NO2        u146(.A(men_men_n162_), .B(men_men_n129_), .Y(men_men_n163_));
  NO2        u147(.A(men_men_n163_), .B(men_men_n161_), .Y(men_men_n164_));
  AOI210     u148(.A0(men_men_n157_), .A1(men_men_n154_), .B0(men_men_n164_), .Y(men_men_n165_));
  OAI210     u149(.A0(men_men_n153_), .A1(men_men_n48_), .B0(men_men_n165_), .Y(men_men_n166_));
  NA2        u150(.A(x5), .B(x1), .Y(men_men_n167_));
  INV        u151(.A(men_men_n167_), .Y(men_men_n168_));
  AOI210     u152(.A0(men_men_n168_), .A1(men_men_n129_), .B0(men_men_n35_), .Y(men_men_n169_));
  NO2        u153(.A(men_men_n60_), .B(men_men_n93_), .Y(men_men_n170_));
  NAi21      u154(.An(x2), .B(x7), .Y(men_men_n171_));
  NO3        u155(.A(men_men_n171_), .B(men_men_n170_), .C(men_men_n46_), .Y(men_men_n172_));
  NA2        u156(.A(men_men_n172_), .B(men_men_n65_), .Y(men_men_n173_));
  NA2        u157(.A(men_men_n173_), .B(men_men_n169_), .Y(men_men_n174_));
  NO4        u158(.A(men_men_n174_), .B(men_men_n166_), .C(men_men_n152_), .D(men_men_n149_), .Y(men_men_n175_));
  NO2        u159(.A(men_men_n175_), .B(men_men_n148_), .Y(men_men_n176_));
  NO2        u160(.A(men_men_n144_), .B(men_men_n140_), .Y(men_men_n177_));
  NA2        u161(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n178_));
  NA2        u162(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n179_));
  NA3        u163(.A(men_men_n179_), .B(men_men_n178_), .C(men_men_n24_), .Y(men_men_n180_));
  AN2        u164(.A(men_men_n180_), .B(men_men_n145_), .Y(men_men_n181_));
  NA2        u165(.A(x8), .B(x0), .Y(men_men_n182_));
  NO2        u166(.A(men_men_n159_), .B(men_men_n25_), .Y(men_men_n183_));
  NO2        u167(.A(men_men_n127_), .B(x4), .Y(men_men_n184_));
  NA2        u168(.A(men_men_n184_), .B(men_men_n183_), .Y(men_men_n185_));
  AOI210     u169(.A0(men_men_n182_), .A1(men_men_n134_), .B0(men_men_n185_), .Y(men_men_n186_));
  NA2        u170(.A(x2), .B(x0), .Y(men_men_n187_));
  NA2        u171(.A(x4), .B(x1), .Y(men_men_n188_));
  NAi21      u172(.An(men_men_n125_), .B(men_men_n188_), .Y(men_men_n189_));
  NOi31      u173(.An(men_men_n189_), .B(men_men_n162_), .C(men_men_n187_), .Y(men_men_n190_));
  NO4        u174(.A(men_men_n190_), .B(men_men_n186_), .C(men_men_n181_), .D(men_men_n177_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n191_), .B(men_men_n41_), .Y(men_men_n192_));
  NO2        u176(.A(men_men_n180_), .B(men_men_n75_), .Y(men_men_n193_));
  INV        u177(.A(men_men_n133_), .Y(men_men_n194_));
  NO2        u178(.A(men_men_n108_), .B(men_men_n17_), .Y(men_men_n195_));
  AOI210     u179(.A0(men_men_n34_), .A1(men_men_n93_), .B0(men_men_n195_), .Y(men_men_n196_));
  NO3        u180(.A(men_men_n196_), .B(men_men_n194_), .C(x7), .Y(men_men_n197_));
  NA3        u181(.A(men_men_n189_), .B(men_men_n194_), .C(men_men_n40_), .Y(men_men_n198_));
  OAI210     u182(.A0(men_men_n179_), .A1(men_men_n140_), .B0(men_men_n198_), .Y(men_men_n199_));
  NO3        u183(.A(men_men_n199_), .B(men_men_n197_), .C(men_men_n193_), .Y(men_men_n200_));
  NO2        u184(.A(men_men_n200_), .B(x3), .Y(men_men_n201_));
  NO3        u185(.A(men_men_n201_), .B(men_men_n192_), .C(men_men_n176_), .Y(men03));
  NO2        u186(.A(men_men_n46_), .B(x3), .Y(men_men_n203_));
  NO2        u187(.A(x6), .B(men_men_n25_), .Y(men_men_n204_));
  INV        u188(.A(men_men_n204_), .Y(men_men_n205_));
  NO2        u189(.A(men_men_n52_), .B(x1), .Y(men_men_n206_));
  OAI210     u190(.A0(men_men_n206_), .A1(men_men_n25_), .B0(men_men_n61_), .Y(men_men_n207_));
  OAI220     u191(.A0(men_men_n207_), .A1(men_men_n17_), .B0(men_men_n205_), .B1(men_men_n108_), .Y(men_men_n208_));
  NA2        u192(.A(men_men_n208_), .B(men_men_n203_), .Y(men_men_n209_));
  NO2        u193(.A(men_men_n77_), .B(x6), .Y(men_men_n210_));
  NA2        u194(.A(x6), .B(men_men_n25_), .Y(men_men_n211_));
  NO2        u195(.A(men_men_n211_), .B(x4), .Y(men_men_n212_));
  NO2        u196(.A(men_men_n18_), .B(x0), .Y(men_men_n213_));
  AO220      u197(.A0(men_men_n213_), .A1(men_men_n212_), .B0(men_men_n210_), .B1(men_men_n53_), .Y(men_men_n214_));
  INV        u198(.A(men_men_n214_), .Y(men_men_n215_));
  NA2        u199(.A(x3), .B(men_men_n17_), .Y(men_men_n216_));
  NA2        u200(.A(x9), .B(men_men_n52_), .Y(men_men_n217_));
  NA2        u201(.A(men_men_n211_), .B(men_men_n80_), .Y(men_men_n218_));
  AOI210     u202(.A0(men_men_n25_), .A1(x3), .B0(men_men_n187_), .Y(men_men_n219_));
  NA2        u203(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n220_));
  NO3        u204(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n221_));
  NO2        u205(.A(x5), .B(x1), .Y(men_men_n222_));
  AOI220     u206(.A0(men_men_n222_), .A1(men_men_n17_), .B0(men_men_n105_), .B1(x5), .Y(men_men_n223_));
  NO2        u207(.A(men_men_n216_), .B(men_men_n178_), .Y(men_men_n224_));
  NO3        u208(.A(x3), .B(x2), .C(x1), .Y(men_men_n225_));
  NO2        u209(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  OAI210     u210(.A0(men_men_n223_), .A1(men_men_n62_), .B0(men_men_n226_), .Y(men_men_n227_));
  AOI220     u211(.A0(men_men_n227_), .A1(men_men_n46_), .B0(men_men_n221_), .B1(men_men_n133_), .Y(men_men_n228_));
  NA4        u212(.A(men_men_n228_), .B(men_men_n220_), .C(men_men_n215_), .D(men_men_n209_), .Y(men_men_n229_));
  NO2        u213(.A(men_men_n46_), .B(men_men_n41_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n230_), .B(men_men_n19_), .Y(men_men_n231_));
  NO2        u215(.A(x3), .B(men_men_n17_), .Y(men_men_n232_));
  NO2        u216(.A(men_men_n232_), .B(x6), .Y(men_men_n233_));
  NOi21      u217(.An(men_men_n83_), .B(men_men_n233_), .Y(men_men_n234_));
  NA2        u218(.A(men_men_n60_), .B(men_men_n93_), .Y(men_men_n235_));
  NA3        u219(.A(men_men_n235_), .B(men_men_n232_), .C(x6), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n236_), .A1(men_men_n234_), .B0(men_men_n159_), .Y(men_men_n237_));
  AO210      u221(.A0(men_men_n237_), .A1(men_men_n231_), .B0(men_men_n183_), .Y(men_men_n238_));
  NA2        u222(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n239_), .A1(men_men_n25_), .B0(men_men_n179_), .Y(men_men_n240_));
  NO3        u224(.A(men_men_n188_), .B(men_men_n60_), .C(x6), .Y(men_men_n241_));
  AOI220     u225(.A0(men_men_n241_), .A1(men_men_n240_), .B0(men_men_n145_), .B1(men_men_n92_), .Y(men_men_n242_));
  NA2        u226(.A(x6), .B(men_men_n46_), .Y(men_men_n243_));
  OAI210     u227(.A0(men_men_n121_), .A1(men_men_n78_), .B0(x4), .Y(men_men_n244_));
  AOI210     u228(.A0(men_men_n244_), .A1(men_men_n243_), .B0(men_men_n77_), .Y(men_men_n245_));
  NO2        u229(.A(men_men_n60_), .B(x6), .Y(men_men_n246_));
  NA2        u230(.A(men_men_n224_), .B(men_men_n246_), .Y(men_men_n247_));
  NA2        u231(.A(men_men_n204_), .B(men_men_n138_), .Y(men_men_n248_));
  NA3        u232(.A(men_men_n216_), .B(men_men_n133_), .C(x6), .Y(men_men_n249_));
  OAI210     u233(.A0(men_men_n93_), .A1(men_men_n35_), .B0(men_men_n65_), .Y(men_men_n250_));
  NA4        u234(.A(men_men_n250_), .B(men_men_n249_), .C(men_men_n248_), .D(men_men_n247_), .Y(men_men_n251_));
  OAI210     u235(.A0(men_men_n251_), .A1(men_men_n245_), .B0(x2), .Y(men_men_n252_));
  NA3        u236(.A(men_men_n252_), .B(men_men_n242_), .C(men_men_n238_), .Y(men_men_n253_));
  AOI210     u237(.A0(men_men_n229_), .A1(x8), .B0(men_men_n253_), .Y(men_men_n254_));
  NO2        u238(.A(men_men_n93_), .B(x3), .Y(men_men_n255_));
  NA2        u239(.A(men_men_n255_), .B(men_men_n212_), .Y(men_men_n256_));
  NO2        u240(.A(men_men_n91_), .B(men_men_n25_), .Y(men_men_n257_));
  AOI210     u241(.A0(men_men_n233_), .A1(men_men_n162_), .B0(men_men_n257_), .Y(men_men_n258_));
  AOI210     u242(.A0(men_men_n258_), .A1(men_men_n256_), .B0(x2), .Y(men_men_n259_));
  NO2        u243(.A(x4), .B(men_men_n52_), .Y(men_men_n260_));
  AOI220     u244(.A0(men_men_n212_), .A1(men_men_n195_), .B0(men_men_n260_), .B1(men_men_n65_), .Y(men_men_n261_));
  NA2        u245(.A(men_men_n60_), .B(x6), .Y(men_men_n262_));
  NA3        u246(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n263_));
  AOI210     u247(.A0(men_men_n263_), .A1(men_men_n144_), .B0(men_men_n262_), .Y(men_men_n264_));
  NA2        u248(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n265_));
  NO2        u249(.A(men_men_n265_), .B(men_men_n25_), .Y(men_men_n266_));
  OAI210     u250(.A0(men_men_n266_), .A1(men_men_n264_), .B0(men_men_n125_), .Y(men_men_n267_));
  NA2        u251(.A(men_men_n216_), .B(x6), .Y(men_men_n268_));
  NO2        u252(.A(men_men_n216_), .B(x6), .Y(men_men_n269_));
  NAi21      u253(.An(men_men_n170_), .B(men_men_n269_), .Y(men_men_n270_));
  NA3        u254(.A(men_men_n270_), .B(men_men_n268_), .C(men_men_n150_), .Y(men_men_n271_));
  NA4        u255(.A(men_men_n271_), .B(men_men_n267_), .C(men_men_n261_), .D(men_men_n159_), .Y(men_men_n272_));
  NA2        u256(.A(men_men_n204_), .B(men_men_n232_), .Y(men_men_n273_));
  NO2        u257(.A(x9), .B(x6), .Y(men_men_n274_));
  NO2        u258(.A(men_men_n144_), .B(men_men_n18_), .Y(men_men_n275_));
  NAi21      u259(.An(men_men_n275_), .B(men_men_n263_), .Y(men_men_n276_));
  NAi21      u260(.An(x1), .B(x4), .Y(men_men_n277_));
  AOI210     u261(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n278_));
  OAI210     u262(.A0(men_men_n144_), .A1(x3), .B0(men_men_n278_), .Y(men_men_n279_));
  AOI220     u263(.A0(men_men_n279_), .A1(men_men_n277_), .B0(men_men_n276_), .B1(men_men_n274_), .Y(men_men_n280_));
  NA2        u264(.A(men_men_n280_), .B(men_men_n273_), .Y(men_men_n281_));
  NA2        u265(.A(men_men_n60_), .B(x2), .Y(men_men_n282_));
  NO2        u266(.A(men_men_n282_), .B(men_men_n273_), .Y(men_men_n283_));
  NO3        u267(.A(x9), .B(x6), .C(x0), .Y(men_men_n284_));
  NA2        u268(.A(men_men_n108_), .B(men_men_n25_), .Y(men_men_n285_));
  NA2        u269(.A(x6), .B(x2), .Y(men_men_n286_));
  NO2        u270(.A(men_men_n286_), .B(men_men_n178_), .Y(men_men_n287_));
  AOI210     u271(.A0(men_men_n285_), .A1(men_men_n284_), .B0(men_men_n287_), .Y(men_men_n288_));
  OAI220     u272(.A0(men_men_n288_), .A1(men_men_n41_), .B0(men_men_n184_), .B1(men_men_n44_), .Y(men_men_n289_));
  OAI210     u273(.A0(men_men_n289_), .A1(men_men_n283_), .B0(men_men_n281_), .Y(men_men_n290_));
  NA2        u274(.A(x9), .B(men_men_n41_), .Y(men_men_n291_));
  NO2        u275(.A(men_men_n291_), .B(men_men_n211_), .Y(men_men_n292_));
  OR3        u276(.A(men_men_n292_), .B(men_men_n210_), .C(men_men_n154_), .Y(men_men_n293_));
  NA2        u277(.A(x4), .B(x0), .Y(men_men_n294_));
  NA2        u278(.A(men_men_n293_), .B(men_men_n40_), .Y(men_men_n295_));
  AOI210     u279(.A0(men_men_n295_), .A1(men_men_n290_), .B0(x8), .Y(men_men_n296_));
  INV        u280(.A(men_men_n262_), .Y(men_men_n297_));
  OAI210     u281(.A0(men_men_n275_), .A1(men_men_n222_), .B0(men_men_n297_), .Y(men_men_n298_));
  INV        u282(.A(men_men_n182_), .Y(men_men_n299_));
  OAI210     u283(.A0(men_men_n299_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n300_));
  AOI210     u284(.A0(men_men_n300_), .A1(men_men_n298_), .B0(men_men_n239_), .Y(men_men_n301_));
  NO4        u285(.A(men_men_n301_), .B(men_men_n296_), .C(men_men_n272_), .D(men_men_n259_), .Y(men_men_n302_));
  NO2        u286(.A(men_men_n170_), .B(x1), .Y(men_men_n303_));
  NO3        u287(.A(men_men_n303_), .B(x3), .C(men_men_n35_), .Y(men_men_n304_));
  OAI210     u288(.A0(men_men_n304_), .A1(men_men_n269_), .B0(x2), .Y(men_men_n305_));
  OAI210     u289(.A0(men_men_n299_), .A1(x6), .B0(men_men_n42_), .Y(men_men_n306_));
  AOI210     u290(.A0(men_men_n306_), .A1(men_men_n305_), .B0(men_men_n194_), .Y(men_men_n307_));
  NOi21      u291(.An(men_men_n286_), .B(men_men_n17_), .Y(men_men_n308_));
  NA3        u292(.A(men_men_n308_), .B(men_men_n222_), .C(men_men_n38_), .Y(men_men_n309_));
  AOI210     u293(.A0(men_men_n35_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n310_));
  NA3        u294(.A(men_men_n310_), .B(men_men_n168_), .C(men_men_n31_), .Y(men_men_n311_));
  NA2        u295(.A(x3), .B(x2), .Y(men_men_n312_));
  AOI220     u296(.A0(men_men_n312_), .A1(men_men_n239_), .B0(men_men_n311_), .B1(men_men_n309_), .Y(men_men_n313_));
  NAi21      u297(.An(x4), .B(x0), .Y(men_men_n314_));
  NO3        u298(.A(men_men_n314_), .B(men_men_n42_), .C(x2), .Y(men_men_n315_));
  OAI210     u299(.A0(x6), .A1(men_men_n18_), .B0(men_men_n315_), .Y(men_men_n316_));
  OAI220     u300(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n317_));
  NO2        u301(.A(x9), .B(x8), .Y(men_men_n318_));
  NA3        u302(.A(men_men_n318_), .B(men_men_n35_), .C(men_men_n52_), .Y(men_men_n319_));
  OAI210     u303(.A0(men_men_n310_), .A1(men_men_n308_), .B0(men_men_n319_), .Y(men_men_n320_));
  AOI220     u304(.A0(men_men_n320_), .A1(men_men_n81_), .B0(men_men_n317_), .B1(men_men_n30_), .Y(men_men_n321_));
  AOI210     u305(.A0(men_men_n321_), .A1(men_men_n316_), .B0(men_men_n25_), .Y(men_men_n322_));
  NA3        u306(.A(men_men_n35_), .B(x1), .C(men_men_n17_), .Y(men_men_n323_));
  OAI210     u307(.A0(men_men_n310_), .A1(men_men_n308_), .B0(men_men_n323_), .Y(men_men_n324_));
  INV        u308(.A(men_men_n224_), .Y(men_men_n325_));
  NA2        u309(.A(men_men_n35_), .B(men_men_n41_), .Y(men_men_n326_));
  OR2        u310(.A(men_men_n326_), .B(men_men_n294_), .Y(men_men_n327_));
  OAI220     u311(.A0(men_men_n327_), .A1(men_men_n167_), .B0(men_men_n243_), .B1(men_men_n325_), .Y(men_men_n328_));
  AO210      u312(.A0(men_men_n324_), .A1(men_men_n154_), .B0(men_men_n328_), .Y(men_men_n329_));
  NO4        u313(.A(men_men_n329_), .B(men_men_n322_), .C(men_men_n313_), .D(men_men_n307_), .Y(men_men_n330_));
  OAI210     u314(.A0(men_men_n302_), .A1(men_men_n254_), .B0(men_men_n330_), .Y(men04));
  OAI210     u315(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n332_));
  NA3        u316(.A(men_men_n332_), .B(men_men_n284_), .C(men_men_n84_), .Y(men_men_n333_));
  NO2        u317(.A(x2), .B(x1), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n265_), .A1(men_men_n334_), .B0(men_men_n35_), .Y(men_men_n335_));
  NO2        u319(.A(men_men_n334_), .B(men_men_n314_), .Y(men_men_n336_));
  AOI210     u320(.A0(men_men_n60_), .A1(x4), .B0(men_men_n114_), .Y(men_men_n337_));
  OAI210     u321(.A0(men_men_n337_), .A1(men_men_n336_), .B0(men_men_n255_), .Y(men_men_n338_));
  NO2        u322(.A(men_men_n282_), .B(men_men_n91_), .Y(men_men_n339_));
  NO2        u323(.A(men_men_n339_), .B(men_men_n35_), .Y(men_men_n340_));
  NO2        u324(.A(men_men_n312_), .B(men_men_n213_), .Y(men_men_n341_));
  NA2        u325(.A(men_men_n341_), .B(men_men_n93_), .Y(men_men_n342_));
  NA3        u326(.A(men_men_n342_), .B(men_men_n340_), .C(men_men_n338_), .Y(men_men_n343_));
  NA2        u327(.A(men_men_n343_), .B(men_men_n335_), .Y(men_men_n344_));
  NO2        u328(.A(men_men_n217_), .B(men_men_n115_), .Y(men_men_n345_));
  NO3        u329(.A(men_men_n262_), .B(men_men_n122_), .C(men_men_n18_), .Y(men_men_n346_));
  NO2        u330(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  OAI210     u331(.A0(men_men_n120_), .A1(men_men_n108_), .B0(men_men_n182_), .Y(men_men_n348_));
  NA3        u332(.A(men_men_n348_), .B(x6), .C(x3), .Y(men_men_n349_));
  AOI210     u333(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n350_));
  OAI220     u334(.A0(men_men_n350_), .A1(men_men_n326_), .B0(men_men_n282_), .B1(men_men_n323_), .Y(men_men_n351_));
  INV        u335(.A(men_men_n351_), .Y(men_men_n352_));
  NA2        u336(.A(x2), .B(men_men_n17_), .Y(men_men_n353_));
  OAI210     u337(.A0(men_men_n108_), .A1(men_men_n17_), .B0(men_men_n353_), .Y(men_men_n354_));
  AOI220     u338(.A0(men_men_n354_), .A1(men_men_n78_), .B0(men_men_n339_), .B1(men_men_n93_), .Y(men_men_n355_));
  NA4        u339(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n349_), .D(men_men_n347_), .Y(men_men_n356_));
  OAI210     u340(.A0(men_men_n113_), .A1(x3), .B0(men_men_n315_), .Y(men_men_n357_));
  NA3        u341(.A(men_men_n235_), .B(men_men_n221_), .C(men_men_n83_), .Y(men_men_n358_));
  NA3        u342(.A(men_men_n358_), .B(men_men_n357_), .C(men_men_n159_), .Y(men_men_n359_));
  AOI210     u343(.A0(men_men_n356_), .A1(x4), .B0(men_men_n359_), .Y(men_men_n360_));
  NA3        u344(.A(men_men_n336_), .B(men_men_n217_), .C(men_men_n93_), .Y(men_men_n361_));
  NOi21      u345(.An(x4), .B(x0), .Y(men_men_n362_));
  XO2        u346(.A(x4), .B(x0), .Y(men_men_n363_));
  OAI210     u347(.A0(men_men_n363_), .A1(men_men_n119_), .B0(men_men_n277_), .Y(men_men_n364_));
  AOI220     u348(.A0(men_men_n364_), .A1(x8), .B0(men_men_n362_), .B1(men_men_n94_), .Y(men_men_n365_));
  AOI210     u349(.A0(men_men_n365_), .A1(men_men_n361_), .B0(x3), .Y(men_men_n366_));
  INV        u350(.A(men_men_n94_), .Y(men_men_n367_));
  NO2        u351(.A(men_men_n93_), .B(x4), .Y(men_men_n368_));
  AOI220     u352(.A0(men_men_n368_), .A1(men_men_n42_), .B0(men_men_n129_), .B1(men_men_n367_), .Y(men_men_n369_));
  NO3        u353(.A(men_men_n363_), .B(men_men_n170_), .C(x2), .Y(men_men_n370_));
  NO3        u354(.A(men_men_n235_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n371_));
  NO2        u355(.A(men_men_n371_), .B(men_men_n370_), .Y(men_men_n372_));
  NA4        u356(.A(men_men_n372_), .B(men_men_n369_), .C(men_men_n231_), .D(x6), .Y(men_men_n373_));
  OAI220     u357(.A0(men_men_n314_), .A1(men_men_n91_), .B0(men_men_n187_), .B1(men_men_n93_), .Y(men_men_n374_));
  NO2        u358(.A(men_men_n41_), .B(x0), .Y(men_men_n375_));
  OR2        u359(.A(men_men_n368_), .B(men_men_n375_), .Y(men_men_n376_));
  NO2        u360(.A(men_men_n156_), .B(men_men_n108_), .Y(men_men_n377_));
  AOI220     u361(.A0(men_men_n377_), .A1(men_men_n376_), .B0(men_men_n374_), .B1(men_men_n59_), .Y(men_men_n378_));
  NO2        u362(.A(men_men_n156_), .B(men_men_n80_), .Y(men_men_n379_));
  NO2        u363(.A(men_men_n34_), .B(x2), .Y(men_men_n380_));
  NOi21      u364(.An(men_men_n125_), .B(men_men_n27_), .Y(men_men_n381_));
  AOI210     u365(.A0(men_men_n380_), .A1(men_men_n379_), .B0(men_men_n381_), .Y(men_men_n382_));
  OAI210     u366(.A0(men_men_n378_), .A1(men_men_n60_), .B0(men_men_n382_), .Y(men_men_n383_));
  OAI220     u367(.A0(men_men_n383_), .A1(x6), .B0(men_men_n373_), .B1(men_men_n366_), .Y(men_men_n384_));
  NA2        u368(.A(men_men_n46_), .B(men_men_n40_), .Y(men_men_n385_));
  OAI210     u369(.A0(men_men_n385_), .A1(men_men_n93_), .B0(men_men_n327_), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n386_), .A1(men_men_n18_), .B0(men_men_n159_), .Y(men_men_n387_));
  AO220      u371(.A0(men_men_n387_), .A1(men_men_n384_), .B0(men_men_n360_), .B1(men_men_n344_), .Y(men_men_n388_));
  NA2        u372(.A(men_men_n380_), .B(x6), .Y(men_men_n389_));
  AOI210     u373(.A0(x6), .A1(x1), .B0(men_men_n158_), .Y(men_men_n390_));
  NA2        u374(.A(men_men_n368_), .B(x0), .Y(men_men_n391_));
  NA2        u375(.A(men_men_n83_), .B(x6), .Y(men_men_n392_));
  OAI210     u376(.A0(men_men_n391_), .A1(men_men_n390_), .B0(men_men_n392_), .Y(men_men_n393_));
  AOI220     u377(.A0(men_men_n393_), .A1(men_men_n389_), .B0(men_men_n225_), .B1(men_men_n47_), .Y(men_men_n394_));
  NA3        u378(.A(men_men_n394_), .B(men_men_n388_), .C(men_men_n333_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n206_), .A1(x8), .B0(men_men_n113_), .Y(men_men_n396_));
  NA2        u380(.A(men_men_n396_), .B(men_men_n353_), .Y(men_men_n397_));
  NA3        u381(.A(men_men_n397_), .B(men_men_n203_), .C(men_men_n159_), .Y(men_men_n398_));
  OAI210     u382(.A0(men_men_n28_), .A1(x1), .B0(men_men_n239_), .Y(men_men_n399_));
  AO220      u383(.A0(men_men_n399_), .A1(men_men_n155_), .B0(men_men_n112_), .B1(x4), .Y(men_men_n400_));
  NA3        u384(.A(x7), .B(x3), .C(x0), .Y(men_men_n401_));
  NA2        u385(.A(men_men_n230_), .B(x0), .Y(men_men_n402_));
  OAI220     u386(.A0(men_men_n402_), .A1(men_men_n217_), .B0(men_men_n401_), .B1(men_men_n367_), .Y(men_men_n403_));
  AOI210     u387(.A0(men_men_n400_), .A1(men_men_n121_), .B0(men_men_n403_), .Y(men_men_n404_));
  AOI210     u388(.A0(men_men_n404_), .A1(men_men_n398_), .B0(men_men_n25_), .Y(men_men_n405_));
  NA3        u389(.A(men_men_n123_), .B(men_men_n230_), .C(x0), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n203_), .A1(men_men_n66_), .B0(men_men_n213_), .Y(men_men_n407_));
  NA3        u391(.A(men_men_n206_), .B(men_men_n232_), .C(x8), .Y(men_men_n408_));
  AOI210     u392(.A0(men_men_n408_), .A1(men_men_n407_), .B0(men_men_n25_), .Y(men_men_n409_));
  AOI210     u393(.A0(men_men_n122_), .A1(men_men_n120_), .B0(men_men_n40_), .Y(men_men_n410_));
  NOi31      u394(.An(men_men_n410_), .B(men_men_n375_), .C(men_men_n188_), .Y(men_men_n411_));
  OAI210     u395(.A0(men_men_n411_), .A1(men_men_n409_), .B0(men_men_n155_), .Y(men_men_n412_));
  NAi31      u396(.An(men_men_n48_), .B(men_men_n303_), .C(men_men_n183_), .Y(men_men_n413_));
  NA3        u397(.A(men_men_n413_), .B(men_men_n412_), .C(men_men_n406_), .Y(men_men_n414_));
  OAI210     u398(.A0(men_men_n414_), .A1(men_men_n405_), .B0(x6), .Y(men_men_n415_));
  OAI210     u399(.A0(men_men_n170_), .A1(men_men_n46_), .B0(men_men_n139_), .Y(men_men_n416_));
  NA3        u400(.A(men_men_n53_), .B(men_men_n37_), .C(men_men_n30_), .Y(men_men_n417_));
  AOI220     u401(.A0(men_men_n417_), .A1(men_men_n416_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n418_));
  NO2        u402(.A(men_men_n159_), .B(x0), .Y(men_men_n419_));
  AOI220     u403(.A0(men_men_n419_), .A1(men_men_n230_), .B0(men_men_n203_), .B1(men_men_n159_), .Y(men_men_n420_));
  AOI210     u404(.A0(men_men_n131_), .A1(men_men_n260_), .B0(x1), .Y(men_men_n421_));
  OAI210     u405(.A0(men_men_n420_), .A1(x8), .B0(men_men_n421_), .Y(men_men_n422_));
  NAi31      u406(.An(x2), .B(x8), .C(x0), .Y(men_men_n423_));
  OAI210     u407(.A0(men_men_n423_), .A1(x4), .B0(men_men_n171_), .Y(men_men_n424_));
  NA3        u408(.A(men_men_n424_), .B(men_men_n153_), .C(x9), .Y(men_men_n425_));
  NO4        u409(.A(men_men_n130_), .B(men_men_n314_), .C(x9), .D(x2), .Y(men_men_n426_));
  NOi21      u410(.An(men_men_n128_), .B(men_men_n187_), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n427_), .B(men_men_n426_), .C(men_men_n18_), .Y(men_men_n428_));
  NO3        u412(.A(x9), .B(men_men_n159_), .C(x0), .Y(men_men_n429_));
  AOI220     u413(.A0(men_men_n429_), .A1(men_men_n255_), .B0(men_men_n379_), .B1(men_men_n159_), .Y(men_men_n430_));
  NA4        u414(.A(men_men_n430_), .B(men_men_n428_), .C(men_men_n425_), .D(men_men_n48_), .Y(men_men_n431_));
  OAI210     u415(.A0(men_men_n422_), .A1(men_men_n418_), .B0(men_men_n431_), .Y(men_men_n432_));
  NOi31      u416(.An(men_men_n419_), .B(men_men_n31_), .C(x8), .Y(men_men_n433_));
  AOI210     u417(.A0(men_men_n37_), .A1(x9), .B0(men_men_n137_), .Y(men_men_n434_));
  NO3        u418(.A(men_men_n434_), .B(men_men_n128_), .C(men_men_n41_), .Y(men_men_n435_));
  NOi31      u419(.An(x1), .B(x8), .C(x7), .Y(men_men_n436_));
  AOI220     u420(.A0(men_men_n436_), .A1(men_men_n362_), .B0(men_men_n129_), .B1(x3), .Y(men_men_n437_));
  AOI210     u421(.A0(men_men_n277_), .A1(men_men_n58_), .B0(men_men_n127_), .Y(men_men_n438_));
  OAI210     u422(.A0(men_men_n438_), .A1(x3), .B0(men_men_n437_), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n439_), .B(men_men_n435_), .C(x2), .Y(men_men_n440_));
  OAI220     u424(.A0(men_men_n363_), .A1(men_men_n318_), .B0(men_men_n314_), .B1(men_men_n41_), .Y(men_men_n441_));
  AOI210     u425(.A0(x9), .A1(men_men_n46_), .B0(men_men_n401_), .Y(men_men_n442_));
  AOI220     u426(.A0(men_men_n442_), .A1(men_men_n93_), .B0(men_men_n441_), .B1(men_men_n159_), .Y(men_men_n443_));
  NO2        u427(.A(men_men_n443_), .B(men_men_n52_), .Y(men_men_n444_));
  NO3        u428(.A(men_men_n444_), .B(men_men_n440_), .C(men_men_n433_), .Y(men_men_n445_));
  AOI210     u429(.A0(men_men_n445_), .A1(men_men_n432_), .B0(men_men_n25_), .Y(men_men_n446_));
  NO3        u430(.A(men_men_n60_), .B(x4), .C(x1), .Y(men_men_n447_));
  NO3        u431(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n448_));
  AOI220     u432(.A0(men_men_n448_), .A1(men_men_n278_), .B0(men_men_n447_), .B1(men_men_n410_), .Y(men_men_n449_));
  NO2        u433(.A(men_men_n449_), .B(men_men_n105_), .Y(men_men_n450_));
  NO3        u434(.A(men_men_n282_), .B(men_men_n182_), .C(men_men_n38_), .Y(men_men_n451_));
  OAI210     u435(.A0(men_men_n451_), .A1(men_men_n450_), .B0(x7), .Y(men_men_n452_));
  NA2        u436(.A(men_men_n235_), .B(x7), .Y(men_men_n453_));
  NA3        u437(.A(men_men_n453_), .B(men_men_n158_), .C(men_men_n138_), .Y(men_men_n454_));
  NA2        u438(.A(men_men_n454_), .B(men_men_n452_), .Y(men_men_n455_));
  OAI210     u439(.A0(men_men_n455_), .A1(men_men_n446_), .B0(men_men_n35_), .Y(men_men_n456_));
  NO2        u440(.A(men_men_n429_), .B(men_men_n213_), .Y(men_men_n457_));
  NO4        u441(.A(men_men_n457_), .B(men_men_n77_), .C(x4), .D(men_men_n52_), .Y(men_men_n458_));
  NA2        u442(.A(men_men_n265_), .B(men_men_n21_), .Y(men_men_n459_));
  NO2        u443(.A(men_men_n167_), .B(men_men_n139_), .Y(men_men_n460_));
  NA2        u444(.A(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  NO2        u445(.A(men_men_n461_), .B(men_men_n28_), .Y(men_men_n462_));
  AOI220     u446(.A0(men_men_n375_), .A1(men_men_n93_), .B0(men_men_n156_), .B1(men_men_n206_), .Y(men_men_n463_));
  NA3        u447(.A(men_men_n463_), .B(men_men_n423_), .C(men_men_n91_), .Y(men_men_n464_));
  NA2        u448(.A(men_men_n464_), .B(men_men_n183_), .Y(men_men_n465_));
  OAI220     u449(.A0(men_men_n291_), .A1(men_men_n67_), .B0(men_men_n167_), .B1(men_men_n41_), .Y(men_men_n466_));
  NA2        u450(.A(x3), .B(men_men_n52_), .Y(men_men_n467_));
  AOI210     u451(.A0(men_men_n171_), .A1(men_men_n27_), .B0(men_men_n72_), .Y(men_men_n468_));
  OAI210     u452(.A0(men_men_n155_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n469_));
  NO3        u453(.A(men_men_n436_), .B(x3), .C(men_men_n52_), .Y(men_men_n470_));
  AOI210     u454(.A0(men_men_n470_), .A1(men_men_n469_), .B0(men_men_n468_), .Y(men_men_n471_));
  OAI210     u455(.A0(men_men_n160_), .A1(men_men_n467_), .B0(men_men_n471_), .Y(men_men_n472_));
  AOI220     u456(.A0(men_men_n472_), .A1(x0), .B0(men_men_n466_), .B1(men_men_n139_), .Y(men_men_n473_));
  AOI210     u457(.A0(men_men_n473_), .A1(men_men_n465_), .B0(men_men_n243_), .Y(men_men_n474_));
  NA2        u458(.A(x9), .B(x5), .Y(men_men_n475_));
  NO4        u459(.A(men_men_n108_), .B(men_men_n475_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n476_));
  NO4        u460(.A(men_men_n476_), .B(men_men_n474_), .C(men_men_n462_), .D(men_men_n458_), .Y(men_men_n477_));
  NA3        u461(.A(men_men_n477_), .B(men_men_n456_), .C(men_men_n415_), .Y(men_men_n478_));
  AOI210     u462(.A0(men_men_n395_), .A1(men_men_n25_), .B0(men_men_n478_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule