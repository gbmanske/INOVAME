library verilog;
use verilog.vl_types.all;
entity freqdiv4_vlg_vec_tst is
end freqdiv4_vlg_vec_tst;
