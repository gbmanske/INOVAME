//Benchmark atmr_intb_466_0.0625

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n316_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n361_, ori_ori_n362_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n352_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n368_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n442_, men_men_n443_, men_men_n444_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  AOI220     o035(.A0(x11), .A1(ori_ori_n48_), .B0(x10), .B1(ori_ori_n57_), .Y(ori_ori_n58_));
  INV        o036(.A(ori_ori_n55_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n60_));
  NA2        o038(.A(ori_ori_n60_), .B(ori_ori_n24_), .Y(ori_ori_n61_));
  OAI220     o039(.A0(ori_ori_n61_), .A1(ori_ori_n59_), .B0(ori_ori_n58_), .B1(ori_ori_n56_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n63_));
  OAI210     o041(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n63_), .Y(ori_ori_n64_));
  AOI220     o042(.A0(ori_ori_n64_), .A1(ori_ori_n55_), .B0(ori_ori_n62_), .B1(ori_ori_n31_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(x05), .Y(ori_ori_n66_));
  NO2        o044(.A(ori_ori_n57_), .B(ori_ori_n23_), .Y(ori_ori_n67_));
  NA2        o045(.A(x09), .B(x05), .Y(ori_ori_n68_));
  NA2        o046(.A(x10), .B(x06), .Y(ori_ori_n69_));
  NA3        o047(.A(ori_ori_n69_), .B(ori_ori_n68_), .C(ori_ori_n28_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n57_), .B(ori_ori_n41_), .Y(ori_ori_n71_));
  OAI210     o049(.A0(ori_ori_n70_), .A1(ori_ori_n67_), .B0(x03), .Y(ori_ori_n72_));
  NOi31      o050(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n73_));
  NO2        o051(.A(x05), .B(ori_ori_n36_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n75_));
  NO2        o053(.A(x08), .B(x01), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n76_), .A1(ori_ori_n75_), .B0(ori_ori_n35_), .Y(ori_ori_n77_));
  NA2        o055(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n77_), .B(x02), .Y(ori_ori_n79_));
  AN2        o057(.A(ori_ori_n79_), .B(ori_ori_n72_), .Y(ori_ori_n80_));
  INV        o058(.A(ori_ori_n77_), .Y(ori_ori_n81_));
  NA2        o059(.A(x11), .B(x00), .Y(ori_ori_n82_));
  NO2        o060(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n83_));
  NOi21      o061(.An(ori_ori_n82_), .B(ori_ori_n83_), .Y(ori_ori_n84_));
  NOi21      o062(.An(x01), .B(x10), .Y(ori_ori_n85_));
  NO2        o063(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n86_));
  NO3        o064(.A(ori_ori_n86_), .B(ori_ori_n85_), .C(x06), .Y(ori_ori_n87_));
  NA2        o065(.A(ori_ori_n87_), .B(ori_ori_n27_), .Y(ori_ori_n88_));
  OAI210     o066(.A0(ori_ori_n361_), .A1(x07), .B0(ori_ori_n88_), .Y(ori_ori_n89_));
  NO3        o067(.A(ori_ori_n89_), .B(ori_ori_n80_), .C(ori_ori_n66_), .Y(ori01));
  INV        o068(.A(x12), .Y(ori_ori_n91_));
  INV        o069(.A(x13), .Y(ori_ori_n92_));
  NA2        o070(.A(ori_ori_n85_), .B(ori_ori_n28_), .Y(ori_ori_n93_));
  NO2        o071(.A(x10), .B(x01), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n95_));
  NO2        o073(.A(ori_ori_n95_), .B(ori_ori_n94_), .Y(ori_ori_n96_));
  NA2        o074(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n97_));
  NO2        o075(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n99_));
  NA2        o077(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n100_), .B(x05), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n102_));
  NA2        o080(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n103_));
  NA2        o081(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n104_), .B(ori_ori_n103_), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n107_));
  NA3        o085(.A(ori_ori_n107_), .B(ori_ori_n106_), .C(x13), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n109_));
  NOi31      o087(.An(ori_ori_n108_), .B(ori_ori_n109_), .C(ori_ori_n105_), .Y(ori_ori_n110_));
  NO3        o088(.A(ori_ori_n110_), .B(x06), .C(x03), .Y(ori_ori_n111_));
  INV        o089(.A(ori_ori_n111_), .Y(ori_ori_n112_));
  NA2        o090(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n113_));
  OAI210     o091(.A0(ori_ori_n76_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(ori_ori_n113_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n117_));
  AOI210     o095(.A0(ori_ori_n117_), .A1(ori_ori_n49_), .B0(ori_ori_n116_), .Y(ori_ori_n118_));
  AN2        o096(.A(ori_ori_n118_), .B(ori_ori_n115_), .Y(ori_ori_n119_));
  NO2        o097(.A(x09), .B(x05), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n47_), .Y(ori_ori_n121_));
  NO2        o099(.A(ori_ori_n96_), .B(ori_ori_n49_), .Y(ori_ori_n122_));
  NA2        o100(.A(x09), .B(x00), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n98_), .B(ori_ori_n123_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n122_), .B(ori_ori_n119_), .Y(ori_ori_n125_));
  NO2        o103(.A(x03), .B(x02), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n77_), .B(ori_ori_n92_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(ori_ori_n126_), .Y(ori_ori_n128_));
  OA210      o106(.A0(ori_ori_n125_), .A1(x11), .B0(ori_ori_n128_), .Y(ori_ori_n129_));
  OAI210     o107(.A0(ori_ori_n112_), .A1(ori_ori_n23_), .B0(ori_ori_n129_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n96_), .B(ori_ori_n40_), .Y(ori_ori_n131_));
  NOi21      o109(.An(x01), .B(x13), .Y(ori_ori_n132_));
  INV        o110(.A(ori_ori_n132_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n131_), .B(ori_ori_n41_), .Y(ori_ori_n134_));
  NO2        o112(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n92_), .B(x01), .Y(ori_ori_n136_));
  NO2        o114(.A(ori_ori_n136_), .B(x08), .Y(ori_ori_n137_));
  NO2        o115(.A(ori_ori_n135_), .B(ori_ori_n48_), .Y(ori_ori_n138_));
  AOI210     o116(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n139_));
  OAI210     o117(.A0(ori_ori_n138_), .A1(ori_ori_n134_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NA2        o118(.A(x10), .B(x05), .Y(ori_ori_n141_));
  NO2        o119(.A(x09), .B(x01), .Y(ori_ori_n142_));
  INV        o120(.A(ori_ori_n25_), .Y(ori_ori_n143_));
  NAi21      o121(.An(x13), .B(x00), .Y(ori_ori_n144_));
  AN2        o122(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n86_), .B(x06), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n144_), .B(ori_ori_n36_), .Y(ori_ori_n147_));
  INV        o125(.A(ori_ori_n147_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n146_), .B(ori_ori_n145_), .Y(ori_ori_n149_));
  NA2        o127(.A(ori_ori_n149_), .B(ori_ori_n143_), .Y(ori_ori_n150_));
  NOi21      o128(.An(x09), .B(x00), .Y(ori_ori_n151_));
  NO3        o129(.A(ori_ori_n75_), .B(ori_ori_n151_), .C(ori_ori_n47_), .Y(ori_ori_n152_));
  NA2        o130(.A(ori_ori_n152_), .B(ori_ori_n104_), .Y(ori_ori_n153_));
  NA2        o131(.A(x06), .B(x05), .Y(ori_ori_n154_));
  OAI210     o132(.A0(ori_ori_n154_), .A1(ori_ori_n35_), .B0(ori_ori_n91_), .Y(ori_ori_n155_));
  AOI210     o133(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n155_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n156_), .B(ori_ori_n153_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n92_), .B(x12), .Y(ori_ori_n158_));
  AOI210     o136(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n158_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n160_), .B(x02), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n159_), .B(ori_ori_n157_), .Y(ori_ori_n162_));
  NA3        o140(.A(ori_ori_n162_), .B(ori_ori_n150_), .C(ori_ori_n140_), .Y(ori_ori_n163_));
  AOI210     o141(.A0(ori_ori_n130_), .A1(ori_ori_n91_), .B0(ori_ori_n163_), .Y(ori_ori_n164_));
  INV        o142(.A(ori_ori_n70_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n165_), .B(ori_ori_n115_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n103_), .B(x06), .Y(ori_ori_n168_));
  INV        o146(.A(ori_ori_n168_), .Y(ori_ori_n169_));
  AOI210     o147(.A0(ori_ori_n169_), .A1(ori_ori_n166_), .B0(x12), .Y(ori_ori_n170_));
  INV        o148(.A(ori_ori_n73_), .Y(ori_ori_n171_));
  NO2        o149(.A(x05), .B(ori_ori_n50_), .Y(ori_ori_n172_));
  OAI210     o150(.A0(ori_ori_n172_), .A1(ori_ori_n133_), .B0(ori_ori_n53_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n173_), .B(ori_ori_n171_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n85_), .B(x06), .Y(ori_ori_n175_));
  AOI210     o153(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n176_));
  NO3        o154(.A(ori_ori_n176_), .B(ori_ori_n175_), .C(ori_ori_n41_), .Y(ori_ori_n177_));
  INV        o155(.A(ori_ori_n117_), .Y(ori_ori_n178_));
  OAI210     o156(.A0(ori_ori_n178_), .A1(ori_ori_n177_), .B0(x02), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n179_), .A1(ori_ori_n174_), .B0(ori_ori_n23_), .Y(ori_ori_n180_));
  OAI210     o158(.A0(ori_ori_n170_), .A1(ori_ori_n53_), .B0(ori_ori_n180_), .Y(ori_ori_n181_));
  INV        o159(.A(ori_ori_n117_), .Y(ori_ori_n182_));
  NO2        o160(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n92_), .B(x03), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n73_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NA2        o163(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n186_));
  NOi21      o164(.An(x13), .B(x04), .Y(ori_ori_n187_));
  NO3        o165(.A(ori_ori_n187_), .B(ori_ori_n73_), .C(ori_ori_n151_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n188_), .B(x05), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n189_), .B(ori_ori_n186_), .Y(ori_ori_n190_));
  NA2        o168(.A(ori_ori_n185_), .B(ori_ori_n190_), .Y(ori_ori_n191_));
  INV        o169(.A(ori_ori_n83_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n192_), .B(x12), .Y(ori_ori_n193_));
  NA2        o171(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n195_));
  AOI210     o173(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n196_));
  NO2        o174(.A(ori_ori_n196_), .B(ori_ori_n41_), .Y(ori_ori_n197_));
  INV        o175(.A(ori_ori_n69_), .Y(ori_ori_n198_));
  NO2        o176(.A(ori_ori_n198_), .B(ori_ori_n197_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n200_));
  NA2        o178(.A(ori_ori_n200_), .B(x03), .Y(ori_ori_n201_));
  OR2        o179(.A(ori_ori_n201_), .B(ori_ori_n199_), .Y(ori_ori_n202_));
  NA2        o180(.A(x13), .B(ori_ori_n91_), .Y(ori_ori_n203_));
  NA3        o181(.A(ori_ori_n203_), .B(ori_ori_n155_), .C(ori_ori_n84_), .Y(ori_ori_n204_));
  OAI210     o182(.A0(ori_ori_n202_), .A1(ori_ori_n194_), .B0(ori_ori_n204_), .Y(ori_ori_n205_));
  AOI210     o183(.A0(ori_ori_n193_), .A1(ori_ori_n191_), .B0(ori_ori_n205_), .Y(ori_ori_n206_));
  AOI210     o184(.A0(ori_ori_n206_), .A1(ori_ori_n181_), .B0(x07), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n68_), .B(ori_ori_n29_), .Y(ori_ori_n208_));
  NOi31      o186(.An(ori_ori_n113_), .B(ori_ori_n187_), .C(ori_ori_n151_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n209_), .B(ori_ori_n208_), .Y(ori_ori_n210_));
  NO2        o188(.A(x08), .B(x05), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(ori_ori_n196_), .Y(ori_ori_n212_));
  OAI210     o190(.A0(ori_ori_n73_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n213_));
  INV        o191(.A(ori_ori_n213_), .Y(ori_ori_n214_));
  NO2        o192(.A(x12), .B(x02), .Y(ori_ori_n215_));
  INV        o193(.A(ori_ori_n215_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n216_), .B(ori_ori_n192_), .Y(ori_ori_n217_));
  OA210      o195(.A0(ori_ori_n214_), .A1(ori_ori_n210_), .B0(ori_ori_n217_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n219_));
  NO2        o197(.A(ori_ori_n219_), .B(x01), .Y(ori_ori_n220_));
  INV        o198(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  AOI210     o199(.A0(ori_ori_n221_), .A1(ori_ori_n108_), .B0(ori_ori_n29_), .Y(ori_ori_n222_));
  NA2        o200(.A(ori_ori_n92_), .B(x04), .Y(ori_ori_n223_));
  NO3        o201(.A(ori_ori_n82_), .B(x12), .C(x03), .Y(ori_ori_n224_));
  NA2        o202(.A(ori_ori_n222_), .B(ori_ori_n224_), .Y(ori_ori_n225_));
  NOi21      o203(.An(ori_ori_n208_), .B(ori_ori_n175_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n226_), .B(ori_ori_n227_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n229_));
  NO3        o207(.A(ori_ori_n229_), .B(ori_ori_n176_), .C(ori_ori_n146_), .Y(ori_ori_n230_));
  NO2        o208(.A(ori_ori_n194_), .B(ori_ori_n28_), .Y(ori_ori_n231_));
  OAI210     o209(.A0(ori_ori_n230_), .A1(ori_ori_n182_), .B0(ori_ori_n231_), .Y(ori_ori_n232_));
  NA3        o210(.A(ori_ori_n232_), .B(ori_ori_n228_), .C(ori_ori_n225_), .Y(ori_ori_n233_));
  NO3        o211(.A(ori_ori_n233_), .B(ori_ori_n218_), .C(ori_ori_n207_), .Y(ori_ori_n234_));
  OAI210     o212(.A0(ori_ori_n164_), .A1(ori_ori_n57_), .B0(ori_ori_n234_), .Y(ori02));
  AOI210     o213(.A0(ori_ori_n113_), .A1(ori_ori_n77_), .B0(ori_ori_n106_), .Y(ori_ori_n236_));
  NOi21      o214(.An(ori_ori_n188_), .B(ori_ori_n142_), .Y(ori_ori_n237_));
  NO2        o215(.A(ori_ori_n237_), .B(ori_ori_n32_), .Y(ori_ori_n238_));
  OAI210     o216(.A0(ori_ori_n238_), .A1(ori_ori_n236_), .B0(ori_ori_n141_), .Y(ori_ori_n239_));
  INV        o217(.A(ori_ori_n141_), .Y(ori_ori_n240_));
  AOI210     o218(.A0(ori_ori_n99_), .A1(ori_ori_n78_), .B0(ori_ori_n176_), .Y(ori_ori_n241_));
  OAI220     o219(.A0(ori_ori_n241_), .A1(ori_ori_n92_), .B0(ori_ori_n77_), .B1(ori_ori_n50_), .Y(ori_ori_n242_));
  AOI220     o220(.A0(ori_ori_n242_), .A1(ori_ori_n240_), .B0(ori_ori_n127_), .B1(ori_ori_n126_), .Y(ori_ori_n243_));
  AOI210     o221(.A0(ori_ori_n243_), .A1(ori_ori_n239_), .B0(ori_ori_n48_), .Y(ori_ori_n244_));
  NO2        o222(.A(x05), .B(x02), .Y(ori_ori_n245_));
  OAI210     o223(.A0(ori_ori_n47_), .A1(ori_ori_n151_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  AOI220     o224(.A0(ori_ori_n211_), .A1(ori_ori_n54_), .B0(ori_ori_n52_), .B1(ori_ori_n36_), .Y(ori_ori_n247_));
  NO2        o225(.A(ori_ori_n246_), .B(ori_ori_n117_), .Y(ori_ori_n248_));
  NAi21      o226(.An(ori_ori_n189_), .B(ori_ori_n185_), .Y(ori_ori_n249_));
  NO2        o227(.A(ori_ori_n200_), .B(ori_ori_n47_), .Y(ori_ori_n250_));
  NA2        o228(.A(ori_ori_n250_), .B(ori_ori_n249_), .Y(ori_ori_n251_));
  OAI210     o229(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n252_));
  NA2        o230(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n253_));
  OA210      o231(.A0(ori_ori_n253_), .A1(x08), .B0(ori_ori_n121_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n254_), .A1(ori_ori_n114_), .B0(ori_ori_n252_), .Y(ori_ori_n255_));
  NA2        o233(.A(ori_ori_n255_), .B(ori_ori_n86_), .Y(ori_ori_n256_));
  INV        o234(.A(ori_ori_n126_), .Y(ori_ori_n257_));
  OAI220     o235(.A0(ori_ori_n212_), .A1(ori_ori_n93_), .B0(ori_ori_n257_), .B1(ori_ori_n105_), .Y(ori_ori_n258_));
  NA2        o236(.A(ori_ori_n258_), .B(x13), .Y(ori_ori_n259_));
  NA3        o237(.A(ori_ori_n259_), .B(ori_ori_n256_), .C(ori_ori_n251_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n260_), .B(ori_ori_n248_), .C(ori_ori_n244_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n116_), .B(x03), .Y(ori_ori_n262_));
  INV        o240(.A(ori_ori_n144_), .Y(ori_ori_n263_));
  NA2        o241(.A(ori_ori_n35_), .B(ori_ori_n36_), .Y(ori_ori_n264_));
  AOI220     o242(.A0(ori_ori_n264_), .A1(ori_ori_n263_), .B0(ori_ori_n160_), .B1(x08), .Y(ori_ori_n265_));
  OAI210     o243(.A0(ori_ori_n265_), .A1(ori_ori_n229_), .B0(ori_ori_n262_), .Y(ori_ori_n266_));
  NA2        o244(.A(ori_ori_n266_), .B(ori_ori_n94_), .Y(ori_ori_n267_));
  INV        o245(.A(ori_ori_n52_), .Y(ori_ori_n268_));
  OAI220     o246(.A0(ori_ori_n223_), .A1(ori_ori_n268_), .B0(ori_ori_n106_), .B1(ori_ori_n28_), .Y(ori_ori_n269_));
  NA2        o247(.A(ori_ori_n269_), .B(ori_ori_n95_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n223_), .B(ori_ori_n91_), .Y(ori_ori_n271_));
  NA2        o249(.A(ori_ori_n91_), .B(ori_ori_n41_), .Y(ori_ori_n272_));
  NA3        o250(.A(ori_ori_n272_), .B(ori_ori_n271_), .C(ori_ori_n105_), .Y(ori_ori_n273_));
  NA4        o251(.A(ori_ori_n273_), .B(ori_ori_n270_), .C(ori_ori_n267_), .D(ori_ori_n48_), .Y(ori_ori_n274_));
  INV        o252(.A(ori_ori_n160_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n276_));
  OAI210     o254(.A0(ori_ori_n275_), .A1(ori_ori_n55_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n277_), .B(x02), .Y(ori_ori_n278_));
  INV        o256(.A(ori_ori_n195_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n158_), .B(x04), .Y(ori_ori_n280_));
  NO3        o258(.A(ori_ori_n158_), .B(ori_ori_n135_), .C(ori_ori_n51_), .Y(ori_ori_n281_));
  OAI210     o259(.A0(ori_ori_n123_), .A1(ori_ori_n36_), .B0(ori_ori_n91_), .Y(ori_ori_n282_));
  OAI210     o260(.A0(ori_ori_n282_), .A1(ori_ori_n152_), .B0(ori_ori_n281_), .Y(ori_ori_n283_));
  NA3        o261(.A(ori_ori_n283_), .B(ori_ori_n278_), .C(x06), .Y(ori_ori_n284_));
  NA2        o262(.A(x09), .B(x03), .Y(ori_ori_n285_));
  OAI220     o263(.A0(ori_ori_n285_), .A1(ori_ori_n104_), .B0(ori_ori_n167_), .B1(ori_ori_n60_), .Y(ori_ori_n286_));
  NO3        o264(.A(ori_ori_n229_), .B(ori_ori_n103_), .C(x08), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n287_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n289_));
  NO3        o267(.A(ori_ori_n98_), .B(ori_ori_n104_), .C(ori_ori_n38_), .Y(ori_ori_n290_));
  AOI210     o268(.A0(ori_ori_n281_), .A1(ori_ori_n289_), .B0(ori_ori_n290_), .Y(ori_ori_n291_));
  OAI210     o269(.A0(ori_ori_n288_), .A1(ori_ori_n28_), .B0(ori_ori_n291_), .Y(ori_ori_n292_));
  AO220      o270(.A0(ori_ori_n292_), .A1(x04), .B0(ori_ori_n286_), .B1(x05), .Y(ori_ori_n293_));
  AOI210     o271(.A0(ori_ori_n284_), .A1(ori_ori_n274_), .B0(ori_ori_n293_), .Y(ori_ori_n294_));
  OAI210     o272(.A0(ori_ori_n261_), .A1(x12), .B0(ori_ori_n294_), .Y(ori03));
  OR2        o273(.A(ori_ori_n42_), .B(ori_ori_n183_), .Y(ori_ori_n296_));
  AOI210     o274(.A0(ori_ori_n127_), .A1(ori_ori_n91_), .B0(ori_ori_n296_), .Y(ori_ori_n297_));
  AO210      o275(.A0(ori_ori_n279_), .A1(ori_ori_n78_), .B0(ori_ori_n280_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n158_), .B(ori_ori_n126_), .Y(ori_ori_n299_));
  NA3        o277(.A(ori_ori_n299_), .B(ori_ori_n298_), .C(ori_ori_n161_), .Y(ori_ori_n300_));
  OAI210     o278(.A0(ori_ori_n300_), .A1(ori_ori_n297_), .B0(x05), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n296_), .B(x05), .Y(ori_ori_n302_));
  AOI210     o280(.A0(ori_ori_n114_), .A1(ori_ori_n171_), .B0(ori_ori_n302_), .Y(ori_ori_n303_));
  AOI210     o281(.A0(ori_ori_n184_), .A1(ori_ori_n74_), .B0(ori_ori_n101_), .Y(ori_ori_n304_));
  OAI220     o282(.A0(ori_ori_n304_), .A1(ori_ori_n55_), .B0(ori_ori_n253_), .B1(ori_ori_n247_), .Y(ori_ori_n305_));
  OAI210     o283(.A0(ori_ori_n305_), .A1(ori_ori_n303_), .B0(ori_ori_n91_), .Y(ori_ori_n306_));
  AOI210     o284(.A0(ori_ori_n121_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n307_));
  NO2        o285(.A(ori_ori_n142_), .B(ori_ori_n109_), .Y(ori_ori_n308_));
  OAI220     o286(.A0(ori_ori_n308_), .A1(ori_ori_n37_), .B0(ori_ori_n124_), .B1(x13), .Y(ori_ori_n309_));
  OAI210     o287(.A0(ori_ori_n309_), .A1(ori_ori_n307_), .B0(x04), .Y(ori_ori_n310_));
  NO3        o288(.A(ori_ori_n272_), .B(ori_ori_n77_), .C(ori_ori_n55_), .Y(ori_ori_n311_));
  AOI210     o289(.A0(ori_ori_n148_), .A1(ori_ori_n91_), .B0(ori_ori_n121_), .Y(ori_ori_n312_));
  OA210      o290(.A0(ori_ori_n137_), .A1(x12), .B0(ori_ori_n109_), .Y(ori_ori_n313_));
  NO3        o291(.A(ori_ori_n313_), .B(ori_ori_n312_), .C(ori_ori_n311_), .Y(ori_ori_n314_));
  NA4        o292(.A(ori_ori_n314_), .B(ori_ori_n310_), .C(ori_ori_n306_), .D(ori_ori_n301_), .Y(ori04));
  NO2        o293(.A(ori_ori_n81_), .B(ori_ori_n39_), .Y(ori_ori_n316_));
  XO2        o294(.A(ori_ori_n316_), .B(ori_ori_n203_), .Y(ori05));
  AOI210     o295(.A0(ori_ori_n68_), .A1(ori_ori_n51_), .B0(ori_ori_n168_), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n318_), .A1(ori_ori_n252_), .B0(ori_ori_n25_), .Y(ori_ori_n319_));
  AOI210     o297(.A0(x06), .A1(x03), .B0(ori_ori_n24_), .Y(ori_ori_n320_));
  OAI210     o298(.A0(ori_ori_n320_), .A1(ori_ori_n319_), .B0(ori_ori_n91_), .Y(ori_ori_n321_));
  NA2        o299(.A(x11), .B(ori_ori_n31_), .Y(ori_ori_n322_));
  NA2        o300(.A(ori_ori_n23_), .B(ori_ori_n28_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n208_), .B(x03), .Y(ori_ori_n324_));
  OAI220     o302(.A0(ori_ori_n324_), .A1(ori_ori_n323_), .B0(ori_ori_n322_), .B1(ori_ori_n362_), .Y(ori_ori_n325_));
  OAI210     o303(.A0(ori_ori_n26_), .A1(ori_ori_n91_), .B0(x07), .Y(ori_ori_n326_));
  AOI210     o304(.A0(ori_ori_n325_), .A1(x06), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n23_), .B(x00), .Y(ori_ori_n328_));
  BUFFER     o306(.A(ori_ori_n194_), .Y(ori_ori_n329_));
  INV        o307(.A(ori_ori_n329_), .Y(ori_ori_n330_));
  OAI210     o308(.A0(ori_ori_n330_), .A1(ori_ori_n328_), .B0(ori_ori_n91_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n33_), .B(ori_ori_n91_), .Y(ori_ori_n332_));
  AOI210     o310(.A0(ori_ori_n332_), .A1(ori_ori_n83_), .B0(x07), .Y(ori_ori_n333_));
  AOI220     o311(.A0(ori_ori_n333_), .A1(ori_ori_n331_), .B0(ori_ori_n327_), .B1(ori_ori_n321_), .Y(ori_ori_n334_));
  AOI210     o312(.A0(ori_ori_n280_), .A1(ori_ori_n97_), .B0(ori_ori_n215_), .Y(ori_ori_n335_));
  NOi21      o313(.An(ori_ori_n262_), .B(ori_ori_n109_), .Y(ori_ori_n336_));
  NO2        o314(.A(ori_ori_n336_), .B(ori_ori_n216_), .Y(ori_ori_n337_));
  OAI210     o315(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n338_));
  AOI210     o316(.A0(ori_ori_n203_), .A1(ori_ori_n47_), .B0(ori_ori_n338_), .Y(ori_ori_n339_));
  NO4        o317(.A(ori_ori_n339_), .B(ori_ori_n337_), .C(ori_ori_n335_), .D(x08), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n106_), .B(ori_ori_n28_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n220_), .Y(ori_ori_n342_));
  NA3        o320(.A(ori_ori_n275_), .B(ori_ori_n102_), .C(x12), .Y(ori_ori_n343_));
  AO210      o321(.A0(ori_ori_n275_), .A1(ori_ori_n102_), .B0(ori_ori_n203_), .Y(ori_ori_n344_));
  NA3        o322(.A(ori_ori_n344_), .B(ori_ori_n343_), .C(x08), .Y(ori_ori_n345_));
  INV        o323(.A(ori_ori_n345_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n340_), .B(ori_ori_n346_), .Y(ori_ori_n347_));
  NA3        o325(.A(ori_ori_n342_), .B(ori_ori_n336_), .C(ori_ori_n271_), .Y(ori_ori_n348_));
  INV        o326(.A(x14), .Y(ori_ori_n349_));
  NO3        o327(.A(ori_ori_n136_), .B(ori_ori_n71_), .C(ori_ori_n53_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n350_), .B(ori_ori_n349_), .Y(ori_ori_n351_));
  NA2        o329(.A(ori_ori_n351_), .B(ori_ori_n348_), .Y(ori_ori_n352_));
  NA2        o330(.A(ori_ori_n332_), .B(ori_ori_n57_), .Y(ori_ori_n353_));
  NOi21      o331(.An(ori_ori_n223_), .B(ori_ori_n124_), .Y(ori_ori_n354_));
  NO2        o332(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n355_));
  OAI210     o333(.A0(ori_ori_n355_), .A1(ori_ori_n354_), .B0(ori_ori_n91_), .Y(ori_ori_n356_));
  OAI210     o334(.A0(ori_ori_n353_), .A1(ori_ori_n82_), .B0(ori_ori_n356_), .Y(ori_ori_n357_));
  NO4        o335(.A(ori_ori_n357_), .B(ori_ori_n352_), .C(ori_ori_n347_), .D(ori_ori_n334_), .Y(ori06));
  INV        o336(.A(ori_ori_n84_), .Y(ori_ori_n361_));
  INV        o337(.A(x02), .Y(ori_ori_n362_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  INV        m039(.A(mai_mai_n59_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n63_), .B(mai_mai_n24_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(mai_mai_n62_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n66_));
  OAI210     m044(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  AOI220     m045(.A0(mai_mai_n67_), .A1(mai_mai_n59_), .B0(mai_mai_n65_), .B1(mai_mai_n31_), .Y(mai_mai_n68_));
  AOI210     m046(.A0(mai_mai_n68_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x09), .B(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x10), .B(x06), .Y(mai_mai_n71_));
  NA3        m049(.A(mai_mai_n71_), .B(mai_mai_n70_), .C(mai_mai_n28_), .Y(mai_mai_n72_));
  OAI210     m050(.A0(mai_mai_n72_), .A1(x11), .B0(x03), .Y(mai_mai_n73_));
  NOi31      m051(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n411_), .B(mai_mai_n24_), .Y(mai_mai_n75_));
  NO2        m053(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n76_), .B(mai_mai_n36_), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n76_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n48_), .B(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n80_));
  NO2        m058(.A(x08), .B(x01), .Y(mai_mai_n81_));
  OAI210     m059(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n35_), .Y(mai_mai_n82_));
  NA2        m060(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n83_));
  NO3        m061(.A(mai_mai_n82_), .B(mai_mai_n79_), .C(mai_mai_n75_), .Y(mai_mai_n84_));
  AN2        m062(.A(mai_mai_n84_), .B(mai_mai_n73_), .Y(mai_mai_n85_));
  INV        m063(.A(mai_mai_n82_), .Y(mai_mai_n86_));
  NO2        m064(.A(x06), .B(x05), .Y(mai_mai_n87_));
  NA2        m065(.A(x11), .B(x00), .Y(mai_mai_n88_));
  NO2        m066(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n89_));
  NOi21      m067(.An(mai_mai_n88_), .B(mai_mai_n89_), .Y(mai_mai_n90_));
  AOI210     m068(.A0(mai_mai_n87_), .A1(mai_mai_n86_), .B0(mai_mai_n90_), .Y(mai_mai_n91_));
  NOi21      m069(.An(x01), .B(x10), .Y(mai_mai_n92_));
  NO2        m070(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n93_));
  NO3        m071(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(x06), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n94_), .B(mai_mai_n27_), .Y(mai_mai_n95_));
  OAI210     m073(.A0(mai_mai_n91_), .A1(x07), .B0(mai_mai_n95_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n85_), .C(mai_mai_n69_), .Y(mai01));
  INV        m075(.A(x12), .Y(mai_mai_n98_));
  INV        m076(.A(x13), .Y(mai_mai_n99_));
  NA2        m077(.A(x08), .B(x04), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n57_), .Y(mai_mai_n101_));
  NA2        m079(.A(mai_mai_n101_), .B(mai_mai_n87_), .Y(mai_mai_n102_));
  NA2        m080(.A(mai_mai_n92_), .B(mai_mai_n28_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n70_), .Y(mai_mai_n104_));
  NO2        m082(.A(x10), .B(x01), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n106_), .B(mai_mai_n105_), .Y(mai_mai_n107_));
  NA2        m085(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n108_));
  NO3        m086(.A(mai_mai_n108_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n109_));
  AOI210     m087(.A0(mai_mai_n109_), .A1(mai_mai_n107_), .B0(mai_mai_n104_), .Y(mai_mai_n110_));
  AOI210     m088(.A0(mai_mai_n110_), .A1(mai_mai_n102_), .B0(mai_mai_n99_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n112_));
  NOi21      m090(.An(mai_mai_n112_), .B(mai_mai_n58_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n114_));
  NA3        m092(.A(x13), .B(mai_mai_n114_), .C(x06), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n115_), .B(mai_mai_n113_), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n81_), .B(x13), .Y(mai_mai_n117_));
  NA2        m095(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n118_));
  NA2        m096(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n119_), .B(x05), .Y(mai_mai_n120_));
  NA2        m098(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n121_));
  AOI210     m099(.A0(mai_mai_n35_), .A1(mai_mai_n77_), .B0(mai_mai_n113_), .Y(mai_mai_n122_));
  AOI210     m100(.A0(mai_mai_n122_), .A1(mai_mai_n117_), .B0(mai_mai_n71_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n124_));
  NA2        m102(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(mai_mai_n124_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n127_));
  NO2        m105(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n128_));
  NO3        m106(.A(x00), .B(x06), .C(x03), .Y(mai_mai_n129_));
  NO4        m107(.A(mai_mai_n129_), .B(mai_mai_n123_), .C(mai_mai_n116_), .D(mai_mai_n111_), .Y(mai_mai_n130_));
  NA2        m108(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n131_));
  OAI210     m109(.A0(mai_mai_n81_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n132_), .B(mai_mai_n131_), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n134_));
  NA2        m112(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n135_));
  AOI210     m113(.A0(mai_mai_n135_), .A1(mai_mai_n49_), .B0(mai_mai_n134_), .Y(mai_mai_n136_));
  AN2        m114(.A(mai_mai_n136_), .B(mai_mai_n133_), .Y(mai_mai_n137_));
  NO2        m115(.A(x09), .B(x05), .Y(mai_mai_n138_));
  NA2        m116(.A(mai_mai_n138_), .B(mai_mai_n47_), .Y(mai_mai_n139_));
  AOI210     m117(.A0(mai_mai_n139_), .A1(mai_mai_n107_), .B0(mai_mai_n49_), .Y(mai_mai_n140_));
  NA2        m118(.A(x09), .B(x00), .Y(mai_mai_n141_));
  NA2        m119(.A(mai_mai_n112_), .B(mai_mai_n141_), .Y(mai_mai_n142_));
  NA2        m120(.A(mai_mai_n74_), .B(mai_mai_n51_), .Y(mai_mai_n143_));
  AOI210     m121(.A0(mai_mai_n143_), .A1(mai_mai_n142_), .B0(mai_mai_n135_), .Y(mai_mai_n144_));
  NO3        m122(.A(mai_mai_n144_), .B(mai_mai_n140_), .C(mai_mai_n137_), .Y(mai_mai_n145_));
  NO2        m123(.A(x03), .B(x02), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n82_), .B(mai_mai_n99_), .Y(mai_mai_n147_));
  OAI210     m125(.A0(mai_mai_n147_), .A1(mai_mai_n113_), .B0(mai_mai_n146_), .Y(mai_mai_n148_));
  OA210      m126(.A0(mai_mai_n145_), .A1(x11), .B0(mai_mai_n148_), .Y(mai_mai_n149_));
  OAI210     m127(.A0(mai_mai_n130_), .A1(mai_mai_n23_), .B0(mai_mai_n149_), .Y(mai_mai_n150_));
  NAi21      m128(.An(x06), .B(x10), .Y(mai_mai_n151_));
  NOi21      m129(.An(x01), .B(x13), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n99_), .B(x01), .Y(mai_mai_n154_));
  NO2        m132(.A(mai_mai_n154_), .B(x08), .Y(mai_mai_n155_));
  AOI210     m133(.A0(x09), .A1(mai_mai_n153_), .B0(mai_mai_n48_), .Y(mai_mai_n156_));
  AOI210     m134(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n157_));
  OAI210     m135(.A0(mai_mai_n156_), .A1(mai_mai_n152_), .B0(mai_mai_n157_), .Y(mai_mai_n158_));
  NA2        m136(.A(x04), .B(x02), .Y(mai_mai_n159_));
  NA2        m137(.A(x10), .B(x05), .Y(mai_mai_n160_));
  NO2        m138(.A(x09), .B(x01), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n105_), .B(mai_mai_n31_), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n162_), .B(x00), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n112_), .B(x08), .Y(mai_mai_n164_));
  OAI210     m142(.A0(mai_mai_n413_), .A1(x11), .B0(mai_mai_n163_), .Y(mai_mai_n165_));
  NAi21      m143(.An(mai_mai_n159_), .B(mai_mai_n165_), .Y(mai_mai_n166_));
  INV        m144(.A(mai_mai_n25_), .Y(mai_mai_n167_));
  NAi21      m145(.An(x13), .B(x00), .Y(mai_mai_n168_));
  AOI210     m146(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n168_), .Y(mai_mai_n169_));
  AN2        m147(.A(x04), .B(mai_mai_n169_), .Y(mai_mai_n170_));
  BUFFER     m148(.A(mai_mai_n70_), .Y(mai_mai_n171_));
  NO2        m149(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n168_), .B(mai_mai_n36_), .Y(mai_mai_n173_));
  INV        m151(.A(mai_mai_n173_), .Y(mai_mai_n174_));
  OAI210     m152(.A0(mai_mai_n172_), .A1(mai_mai_n171_), .B0(mai_mai_n174_), .Y(mai_mai_n175_));
  OAI210     m153(.A0(mai_mai_n175_), .A1(mai_mai_n170_), .B0(mai_mai_n167_), .Y(mai_mai_n176_));
  NOi21      m154(.An(x09), .B(x00), .Y(mai_mai_n177_));
  NO3        m155(.A(mai_mai_n80_), .B(mai_mai_n177_), .C(mai_mai_n47_), .Y(mai_mai_n178_));
  NA2        m156(.A(x06), .B(x05), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n99_), .B(x12), .Y(mai_mai_n180_));
  NA2        m158(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n181_));
  NA2        m159(.A(mai_mai_n92_), .B(mai_mai_n51_), .Y(mai_mai_n182_));
  NO2        m160(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n183_));
  NA2        m161(.A(mai_mai_n183_), .B(x02), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n184_), .B(mai_mai_n182_), .Y(mai_mai_n185_));
  AOI210     m163(.A0(mai_mai_n181_), .A1(x12), .B0(mai_mai_n185_), .Y(mai_mai_n186_));
  NA4        m164(.A(mai_mai_n186_), .B(mai_mai_n176_), .C(mai_mai_n166_), .D(mai_mai_n158_), .Y(mai_mai_n187_));
  AOI210     m165(.A0(mai_mai_n150_), .A1(mai_mai_n98_), .B0(mai_mai_n187_), .Y(mai_mai_n188_));
  INV        m166(.A(mai_mai_n72_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(mai_mai_n133_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n191_));
  NA2        m169(.A(mai_mai_n191_), .B(mai_mai_n132_), .Y(mai_mai_n192_));
  AOI210     m170(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n124_), .B(x06), .Y(mai_mai_n194_));
  AOI210     m172(.A0(mai_mai_n193_), .A1(mai_mai_n192_), .B0(mai_mai_n194_), .Y(mai_mai_n195_));
  AOI210     m173(.A0(mai_mai_n195_), .A1(mai_mai_n190_), .B0(x12), .Y(mai_mai_n196_));
  INV        m174(.A(mai_mai_n74_), .Y(mai_mai_n197_));
  NO2        m175(.A(mai_mai_n92_), .B(x06), .Y(mai_mai_n198_));
  AOI210     m176(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n199_));
  NO3        m177(.A(mai_mai_n199_), .B(mai_mai_n198_), .C(mai_mai_n41_), .Y(mai_mai_n200_));
  NA4        m178(.A(mai_mai_n151_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n201_));
  NA2        m179(.A(mai_mai_n201_), .B(mai_mai_n135_), .Y(mai_mai_n202_));
  OAI210     m180(.A0(mai_mai_n202_), .A1(mai_mai_n200_), .B0(x02), .Y(mai_mai_n203_));
  AOI210     m181(.A0(mai_mai_n203_), .A1(mai_mai_n57_), .B0(mai_mai_n23_), .Y(mai_mai_n204_));
  OAI210     m182(.A0(mai_mai_n196_), .A1(mai_mai_n57_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  INV        m183(.A(mai_mai_n135_), .Y(mai_mai_n206_));
  NO2        m184(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n207_));
  OAI210     m185(.A0(mai_mai_n76_), .A1(mai_mai_n36_), .B0(mai_mai_n118_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n99_), .B(x03), .Y(mai_mai_n209_));
  NA2        m187(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n210_));
  INV        m188(.A(mai_mai_n151_), .Y(mai_mai_n211_));
  NOi21      m189(.An(x13), .B(x04), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n212_), .B(mai_mai_n177_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n213_), .B(x05), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n211_), .B(mai_mai_n57_), .Y(mai_mai_n215_));
  OAI210     m193(.A0(mai_mai_n210_), .A1(mai_mai_n206_), .B0(mai_mai_n215_), .Y(mai_mai_n216_));
  INV        m194(.A(mai_mai_n89_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n217_), .B(x12), .Y(mai_mai_n218_));
  NA2        m196(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n220_));
  INV        m198(.A(mai_mai_n169_), .Y(mai_mai_n221_));
  AOI210     m199(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n222_));
  NO2        m200(.A(x06), .B(x00), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n224_), .B(x03), .Y(mai_mai_n225_));
  OA210      m203(.A0(mai_mai_n225_), .A1(mai_mai_n223_), .B0(mai_mai_n221_), .Y(mai_mai_n226_));
  NA2        m204(.A(x13), .B(mai_mai_n98_), .Y(mai_mai_n227_));
  NA3        m205(.A(mai_mai_n227_), .B(x12), .C(mai_mai_n90_), .Y(mai_mai_n228_));
  OAI210     m206(.A0(mai_mai_n226_), .A1(mai_mai_n219_), .B0(mai_mai_n228_), .Y(mai_mai_n229_));
  AOI210     m207(.A0(mai_mai_n218_), .A1(mai_mai_n216_), .B0(mai_mai_n229_), .Y(mai_mai_n230_));
  AOI210     m208(.A0(mai_mai_n230_), .A1(mai_mai_n205_), .B0(x07), .Y(mai_mai_n231_));
  NA2        m209(.A(mai_mai_n70_), .B(mai_mai_n29_), .Y(mai_mai_n232_));
  NO2        m210(.A(mai_mai_n212_), .B(mai_mai_n177_), .Y(mai_mai_n233_));
  AOI210     m211(.A0(mai_mai_n233_), .A1(mai_mai_n143_), .B0(mai_mai_n232_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n99_), .B(x06), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n235_), .Y(mai_mai_n236_));
  NO2        m214(.A(x08), .B(x05), .Y(mai_mai_n237_));
  NO2        m215(.A(mai_mai_n237_), .B(mai_mai_n222_), .Y(mai_mai_n238_));
  NA2        m216(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n239_));
  OAI210     m217(.A0(mai_mai_n238_), .A1(mai_mai_n236_), .B0(mai_mai_n239_), .Y(mai_mai_n240_));
  NO2        m218(.A(x12), .B(x02), .Y(mai_mai_n241_));
  INV        m219(.A(mai_mai_n241_), .Y(mai_mai_n242_));
  NO2        m220(.A(mai_mai_n242_), .B(mai_mai_n217_), .Y(mai_mai_n243_));
  OA210      m221(.A0(mai_mai_n240_), .A1(mai_mai_n234_), .B0(mai_mai_n243_), .Y(mai_mai_n244_));
  NA2        m222(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n245_), .B(x01), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n235_), .B(mai_mai_n208_), .Y(mai_mai_n247_));
  NA2        m225(.A(mai_mai_n99_), .B(x04), .Y(mai_mai_n248_));
  OAI210     m226(.A0(x02), .A1(mai_mai_n117_), .B0(mai_mai_n247_), .Y(mai_mai_n249_));
  NO3        m227(.A(mai_mai_n88_), .B(x12), .C(x03), .Y(mai_mai_n250_));
  OAI210     m228(.A0(mai_mai_n249_), .A1(mai_mai_n81_), .B0(mai_mai_n250_), .Y(mai_mai_n251_));
  AOI210     m229(.A0(mai_mai_n182_), .A1(mai_mai_n179_), .B0(mai_mai_n100_), .Y(mai_mai_n252_));
  NOi21      m230(.An(mai_mai_n232_), .B(mai_mai_n198_), .Y(mai_mai_n253_));
  NO2        m231(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n254_));
  OAI210     m232(.A0(mai_mai_n253_), .A1(mai_mai_n252_), .B0(mai_mai_n254_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n256_));
  NO3        m234(.A(mai_mai_n256_), .B(mai_mai_n199_), .C(mai_mai_n172_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n219_), .B(mai_mai_n28_), .Y(mai_mai_n258_));
  OAI210     m236(.A0(mai_mai_n257_), .A1(mai_mai_n206_), .B0(mai_mai_n258_), .Y(mai_mai_n259_));
  NA3        m237(.A(mai_mai_n259_), .B(mai_mai_n255_), .C(mai_mai_n251_), .Y(mai_mai_n260_));
  NO3        m238(.A(mai_mai_n260_), .B(mai_mai_n244_), .C(mai_mai_n231_), .Y(mai_mai_n261_));
  OAI210     m239(.A0(mai_mai_n188_), .A1(mai_mai_n61_), .B0(mai_mai_n261_), .Y(mai02));
  NOi21      m240(.An(mai_mai_n213_), .B(mai_mai_n161_), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n99_), .B(mai_mai_n35_), .Y(mai_mai_n264_));
  NA3        m242(.A(mai_mai_n264_), .B(x10), .C(mai_mai_n56_), .Y(mai_mai_n265_));
  OAI210     m243(.A0(mai_mai_n263_), .A1(mai_mai_n32_), .B0(mai_mai_n265_), .Y(mai_mai_n266_));
  NA2        m244(.A(mai_mai_n266_), .B(mai_mai_n160_), .Y(mai_mai_n267_));
  INV        m245(.A(mai_mai_n160_), .Y(mai_mai_n268_));
  AOI210     m246(.A0(mai_mai_n114_), .A1(mai_mai_n83_), .B0(mai_mai_n199_), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n269_), .B(mai_mai_n99_), .Y(mai_mai_n270_));
  AOI220     m248(.A0(mai_mai_n270_), .A1(mai_mai_n268_), .B0(mai_mai_n147_), .B1(mai_mai_n146_), .Y(mai_mai_n271_));
  AOI210     m249(.A0(mai_mai_n271_), .A1(mai_mai_n267_), .B0(mai_mai_n48_), .Y(mai_mai_n272_));
  NO2        m250(.A(x05), .B(x02), .Y(mai_mai_n273_));
  OAI210     m251(.A0(mai_mai_n192_), .A1(mai_mai_n177_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  AOI220     m252(.A0(mai_mai_n237_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n275_));
  NOi21      m253(.An(mai_mai_n264_), .B(mai_mai_n275_), .Y(mai_mai_n276_));
  AOI210     m254(.A0(mai_mai_n212_), .A1(mai_mai_n76_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  AOI210     m255(.A0(mai_mai_n277_), .A1(mai_mai_n274_), .B0(mai_mai_n135_), .Y(mai_mai_n278_));
  NAi21      m256(.An(mai_mai_n214_), .B(mai_mai_n210_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n224_), .B(mai_mai_n47_), .Y(mai_mai_n280_));
  NA2        m258(.A(mai_mai_n280_), .B(mai_mai_n279_), .Y(mai_mai_n281_));
  AN2        m259(.A(mai_mai_n209_), .B(mai_mai_n208_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n283_));
  NA2        m261(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n284_));
  OA210      m262(.A0(mai_mai_n284_), .A1(x08), .B0(mai_mai_n139_), .Y(mai_mai_n285_));
  AOI210     m263(.A0(mai_mai_n285_), .A1(mai_mai_n132_), .B0(mai_mai_n283_), .Y(mai_mai_n286_));
  OAI210     m264(.A0(mai_mai_n286_), .A1(mai_mai_n282_), .B0(mai_mai_n93_), .Y(mai_mai_n287_));
  NA3        m265(.A(mai_mai_n93_), .B(mai_mai_n81_), .C(mai_mai_n207_), .Y(mai_mai_n288_));
  NA3        m266(.A(mai_mai_n92_), .B(mai_mai_n80_), .C(mai_mai_n42_), .Y(mai_mai_n289_));
  AOI210     m267(.A0(mai_mai_n289_), .A1(mai_mai_n288_), .B0(x04), .Y(mai_mai_n290_));
  NO2        m268(.A(mai_mai_n238_), .B(mai_mai_n103_), .Y(mai_mai_n291_));
  AOI210     m269(.A0(mai_mai_n291_), .A1(x13), .B0(mai_mai_n290_), .Y(mai_mai_n292_));
  NA3        m270(.A(mai_mai_n292_), .B(mai_mai_n287_), .C(mai_mai_n281_), .Y(mai_mai_n293_));
  NO3        m271(.A(mai_mai_n293_), .B(mai_mai_n278_), .C(mai_mai_n272_), .Y(mai_mai_n294_));
  NA2        m272(.A(mai_mai_n134_), .B(x03), .Y(mai_mai_n295_));
  INV        m273(.A(mai_mai_n168_), .Y(mai_mai_n296_));
  AOI220     m274(.A0(x08), .A1(mai_mai_n296_), .B0(mai_mai_n183_), .B1(x08), .Y(mai_mai_n297_));
  OAI210     m275(.A0(mai_mai_n297_), .A1(mai_mai_n256_), .B0(mai_mai_n295_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n298_), .B(mai_mai_n105_), .Y(mai_mai_n299_));
  NA2        m277(.A(mai_mai_n159_), .B(mai_mai_n154_), .Y(mai_mai_n300_));
  AN2        m278(.A(mai_mai_n300_), .B(mai_mai_n164_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n127_), .B(mai_mai_n28_), .Y(mai_mai_n302_));
  OAI210     m280(.A0(mai_mai_n302_), .A1(mai_mai_n301_), .B0(mai_mai_n106_), .Y(mai_mai_n303_));
  NA2        m281(.A(mai_mai_n248_), .B(mai_mai_n98_), .Y(mai_mai_n304_));
  NA2        m282(.A(mai_mai_n98_), .B(mai_mai_n41_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n305_), .B(mai_mai_n304_), .C(mai_mai_n126_), .Y(mai_mai_n306_));
  NA4        m284(.A(mai_mai_n306_), .B(mai_mai_n303_), .C(mai_mai_n299_), .D(mai_mai_n48_), .Y(mai_mai_n307_));
  INV        m285(.A(mai_mai_n183_), .Y(mai_mai_n308_));
  NA2        m286(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n309_));
  OAI220     m287(.A0(mai_mai_n309_), .A1(mai_mai_n412_), .B0(mai_mai_n308_), .B1(mai_mai_n59_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n310_), .B(x02), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n220_), .Y(mai_mai_n312_));
  NA2        m290(.A(mai_mai_n180_), .B(x04), .Y(mai_mai_n313_));
  NO2        m291(.A(mai_mai_n313_), .B(mai_mai_n312_), .Y(mai_mai_n314_));
  NO2        m292(.A(x13), .B(mai_mai_n31_), .Y(mai_mai_n315_));
  OAI210     m293(.A0(mai_mai_n315_), .A1(mai_mai_n314_), .B0(mai_mai_n93_), .Y(mai_mai_n316_));
  NO3        m294(.A(mai_mai_n180_), .B(mai_mai_n153_), .C(mai_mai_n52_), .Y(mai_mai_n317_));
  OAI210     m295(.A0(mai_mai_n141_), .A1(mai_mai_n36_), .B0(mai_mai_n98_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n318_), .A1(mai_mai_n178_), .B0(mai_mai_n317_), .Y(mai_mai_n319_));
  NA4        m297(.A(mai_mai_n319_), .B(mai_mai_n316_), .C(mai_mai_n311_), .D(x06), .Y(mai_mai_n320_));
  NA2        m298(.A(x09), .B(x03), .Y(mai_mai_n321_));
  OAI220     m299(.A0(mai_mai_n321_), .A1(mai_mai_n125_), .B0(mai_mai_n191_), .B1(mai_mai_n63_), .Y(mai_mai_n322_));
  OAI220     m300(.A0(mai_mai_n154_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n323_));
  NO3        m301(.A(mai_mai_n256_), .B(mai_mai_n124_), .C(x08), .Y(mai_mai_n324_));
  AOI210     m302(.A0(mai_mai_n323_), .A1(mai_mai_n206_), .B0(mai_mai_n324_), .Y(mai_mai_n325_));
  NO3        m303(.A(mai_mai_n112_), .B(mai_mai_n125_), .C(mai_mai_n38_), .Y(mai_mai_n326_));
  INV        m304(.A(mai_mai_n326_), .Y(mai_mai_n327_));
  OAI210     m305(.A0(mai_mai_n325_), .A1(mai_mai_n28_), .B0(mai_mai_n327_), .Y(mai_mai_n328_));
  AO220      m306(.A0(mai_mai_n328_), .A1(x04), .B0(mai_mai_n322_), .B1(x05), .Y(mai_mai_n329_));
  AOI210     m307(.A0(mai_mai_n320_), .A1(mai_mai_n307_), .B0(mai_mai_n329_), .Y(mai_mai_n330_));
  OAI210     m308(.A0(mai_mai_n294_), .A1(x12), .B0(mai_mai_n330_), .Y(mai03));
  OR2        m309(.A(mai_mai_n42_), .B(mai_mai_n207_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n147_), .A1(mai_mai_n98_), .B0(mai_mai_n332_), .Y(mai_mai_n333_));
  AO210      m311(.A0(mai_mai_n312_), .A1(mai_mai_n83_), .B0(mai_mai_n313_), .Y(mai_mai_n334_));
  NA2        m312(.A(mai_mai_n180_), .B(mai_mai_n146_), .Y(mai_mai_n335_));
  NA3        m313(.A(mai_mai_n335_), .B(mai_mai_n334_), .C(mai_mai_n184_), .Y(mai_mai_n336_));
  OAI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n333_), .B0(x05), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n332_), .B(x05), .Y(mai_mai_n338_));
  AOI210     m316(.A0(mai_mai_n132_), .A1(mai_mai_n197_), .B0(mai_mai_n338_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n209_), .A1(mai_mai_n77_), .B0(mai_mai_n120_), .Y(mai_mai_n340_));
  OAI220     m318(.A0(mai_mai_n340_), .A1(mai_mai_n59_), .B0(mai_mai_n284_), .B1(mai_mai_n275_), .Y(mai_mai_n341_));
  OAI210     m319(.A0(mai_mai_n341_), .A1(mai_mai_n339_), .B0(mai_mai_n98_), .Y(mai_mai_n342_));
  AOI210     m320(.A0(mai_mai_n139_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n343_));
  NO2        m321(.A(mai_mai_n161_), .B(mai_mai_n128_), .Y(mai_mai_n344_));
  OAI220     m322(.A0(mai_mai_n344_), .A1(mai_mai_n37_), .B0(mai_mai_n142_), .B1(x13), .Y(mai_mai_n345_));
  OAI210     m323(.A0(mai_mai_n345_), .A1(mai_mai_n343_), .B0(x04), .Y(mai_mai_n346_));
  NO3        m324(.A(mai_mai_n305_), .B(mai_mai_n82_), .C(mai_mai_n59_), .Y(mai_mai_n347_));
  AOI210     m325(.A0(mai_mai_n174_), .A1(mai_mai_n98_), .B0(mai_mai_n139_), .Y(mai_mai_n348_));
  OA210      m326(.A0(mai_mai_n155_), .A1(x12), .B0(mai_mai_n128_), .Y(mai_mai_n349_));
  NO3        m327(.A(mai_mai_n349_), .B(mai_mai_n348_), .C(mai_mai_n347_), .Y(mai_mai_n350_));
  NA4        m328(.A(mai_mai_n350_), .B(mai_mai_n346_), .C(mai_mai_n342_), .D(mai_mai_n337_), .Y(mai04));
  NO2        m329(.A(mai_mai_n86_), .B(mai_mai_n39_), .Y(mai_mai_n352_));
  XO2        m330(.A(mai_mai_n352_), .B(mai_mai_n227_), .Y(mai05));
  NO2        m331(.A(mai_mai_n283_), .B(mai_mai_n25_), .Y(mai_mai_n354_));
  NA3        m332(.A(mai_mai_n135_), .B(mai_mai_n127_), .C(mai_mai_n31_), .Y(mai_mai_n355_));
  NO2        m333(.A(mai_mai_n355_), .B(mai_mai_n24_), .Y(mai_mai_n356_));
  OAI210     m334(.A0(mai_mai_n356_), .A1(mai_mai_n354_), .B0(mai_mai_n98_), .Y(mai_mai_n357_));
  OAI210     m335(.A0(mai_mai_n26_), .A1(mai_mai_n98_), .B0(x07), .Y(mai_mai_n358_));
  INV        m336(.A(mai_mai_n358_), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n152_), .B(x05), .Y(mai_mai_n360_));
  NA3        m338(.A(mai_mai_n360_), .B(mai_mai_n223_), .C(mai_mai_n217_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n362_));
  OAI210     m340(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n363_));
  OR3        m341(.A(mai_mai_n363_), .B(mai_mai_n362_), .C(mai_mai_n44_), .Y(mai_mai_n364_));
  NA2        m342(.A(mai_mai_n364_), .B(mai_mai_n361_), .Y(mai_mai_n365_));
  NA2        m343(.A(mai_mai_n365_), .B(mai_mai_n98_), .Y(mai_mai_n366_));
  NA2        m344(.A(mai_mai_n33_), .B(mai_mai_n98_), .Y(mai_mai_n367_));
  AOI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n89_), .B0(x07), .Y(mai_mai_n368_));
  AOI220     m346(.A0(mai_mai_n368_), .A1(mai_mai_n366_), .B0(mai_mai_n359_), .B1(mai_mai_n357_), .Y(mai_mai_n369_));
  OR2        m347(.A(mai_mai_n245_), .B(mai_mai_n242_), .Y(mai_mai_n370_));
  AOI210     m348(.A0(mai_mai_n362_), .A1(x07), .B0(mai_mai_n134_), .Y(mai_mai_n371_));
  OR2        m349(.A(mai_mai_n371_), .B(x03), .Y(mai_mai_n372_));
  NO2        m350(.A(x07), .B(x11), .Y(mai_mai_n373_));
  NO3        m351(.A(mai_mai_n373_), .B(mai_mai_n138_), .C(mai_mai_n28_), .Y(mai_mai_n374_));
  AOI220     m352(.A0(mai_mai_n374_), .A1(mai_mai_n372_), .B0(mai_mai_n370_), .B1(mai_mai_n47_), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n375_), .B(mai_mai_n99_), .Y(mai_mai_n376_));
  AOI210     m354(.A0(mai_mai_n313_), .A1(mai_mai_n108_), .B0(mai_mai_n241_), .Y(mai_mai_n377_));
  NOi21      m355(.An(mai_mai_n295_), .B(mai_mai_n128_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(mai_mai_n242_), .Y(mai_mai_n379_));
  OAI210     m357(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n380_));
  AOI210     m358(.A0(mai_mai_n227_), .A1(mai_mai_n47_), .B0(mai_mai_n380_), .Y(mai_mai_n381_));
  NO4        m359(.A(mai_mai_n381_), .B(mai_mai_n379_), .C(mai_mai_n377_), .D(x08), .Y(mai_mai_n382_));
  NA2        m360(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n383_), .B(x03), .Y(mai_mai_n384_));
  NO2        m362(.A(x13), .B(x12), .Y(mai_mai_n385_));
  NO2        m363(.A(mai_mai_n127_), .B(mai_mai_n28_), .Y(mai_mai_n386_));
  NO2        m364(.A(mai_mai_n386_), .B(mai_mai_n246_), .Y(mai_mai_n387_));
  OR3        m365(.A(mai_mai_n387_), .B(x12), .C(x03), .Y(mai_mai_n388_));
  NA3        m366(.A(mai_mai_n308_), .B(mai_mai_n121_), .C(x12), .Y(mai_mai_n389_));
  AO210      m367(.A0(mai_mai_n308_), .A1(mai_mai_n121_), .B0(mai_mai_n227_), .Y(mai_mai_n390_));
  NA4        m368(.A(mai_mai_n390_), .B(mai_mai_n389_), .C(mai_mai_n388_), .D(x08), .Y(mai_mai_n391_));
  AOI210     m369(.A0(mai_mai_n385_), .A1(mai_mai_n384_), .B0(mai_mai_n391_), .Y(mai_mai_n392_));
  AOI210     m370(.A0(mai_mai_n382_), .A1(mai_mai_n376_), .B0(mai_mai_n392_), .Y(mai_mai_n393_));
  INV        m371(.A(x07), .Y(mai_mai_n394_));
  OAI220     m372(.A0(mai_mai_n394_), .A1(x02), .B0(mai_mai_n138_), .B1(mai_mai_n43_), .Y(mai_mai_n395_));
  OAI210     m373(.A0(mai_mai_n395_), .A1(x11), .B0(mai_mai_n173_), .Y(mai_mai_n396_));
  NA3        m374(.A(mai_mai_n387_), .B(mai_mai_n378_), .C(mai_mai_n304_), .Y(mai_mai_n397_));
  INV        m375(.A(x14), .Y(mai_mai_n398_));
  NO3        m376(.A(mai_mai_n295_), .B(mai_mai_n103_), .C(x11), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n399_), .B(mai_mai_n398_), .Y(mai_mai_n400_));
  NA3        m378(.A(mai_mai_n400_), .B(mai_mai_n397_), .C(mai_mai_n396_), .Y(mai_mai_n401_));
  AOI220     m379(.A0(mai_mai_n367_), .A1(mai_mai_n61_), .B0(mai_mai_n386_), .B1(mai_mai_n153_), .Y(mai_mai_n402_));
  NOi21      m380(.An(mai_mai_n248_), .B(mai_mai_n142_), .Y(mai_mai_n403_));
  NA2        m381(.A(mai_mai_n254_), .B(mai_mai_n211_), .Y(mai_mai_n404_));
  OAI210     m382(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n404_), .Y(mai_mai_n405_));
  OAI210     m383(.A0(mai_mai_n405_), .A1(mai_mai_n403_), .B0(mai_mai_n98_), .Y(mai_mai_n406_));
  OAI210     m384(.A0(mai_mai_n402_), .A1(mai_mai_n88_), .B0(mai_mai_n406_), .Y(mai_mai_n407_));
  NO4        m385(.A(mai_mai_n407_), .B(mai_mai_n401_), .C(mai_mai_n393_), .D(mai_mai_n369_), .Y(mai06));
  INV        m386(.A(x07), .Y(mai_mai_n411_));
  INV        m387(.A(mai_mai_n40_), .Y(mai_mai_n412_));
  INV        m388(.A(x01), .Y(mai_mai_n413_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI210     u039(.A0(x11), .A1(men_men_n48_), .B0(men_men_n61_), .Y(men_men_n62_));
  INV        u040(.A(men_men_n59_), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n29_), .B(x02), .Y(men_men_n64_));
  NA2        u042(.A(men_men_n64_), .B(men_men_n24_), .Y(men_men_n65_));
  OAI220     u043(.A0(men_men_n65_), .A1(men_men_n63_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n66_));
  NA2        u044(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n67_));
  OAI210     u045(.A0(men_men_n30_), .A1(x11), .B0(men_men_n67_), .Y(men_men_n68_));
  AOI220     u046(.A0(men_men_n68_), .A1(men_men_n59_), .B0(men_men_n66_), .B1(men_men_n31_), .Y(men_men_n69_));
  AOI210     u047(.A0(men_men_n69_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n70_));
  NA2        u048(.A(x10), .B(x09), .Y(men_men_n71_));
  NA2        u049(.A(x09), .B(x05), .Y(men_men_n72_));
  NA2        u050(.A(x10), .B(x06), .Y(men_men_n73_));
  NA2        u051(.A(men_men_n73_), .B(men_men_n72_), .Y(men_men_n74_));
  NO2        u052(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n75_));
  OAI210     u053(.A0(men_men_n74_), .A1(x07), .B0(x03), .Y(men_men_n76_));
  NOi31      u054(.An(x08), .B(x04), .C(x00), .Y(men_men_n77_));
  NO2        u055(.A(x10), .B(x09), .Y(men_men_n78_));
  NO2        u056(.A(men_men_n442_), .B(men_men_n24_), .Y(men_men_n79_));
  NO2        u057(.A(x09), .B(men_men_n41_), .Y(men_men_n80_));
  NO2        u058(.A(men_men_n80_), .B(men_men_n36_), .Y(men_men_n81_));
  OAI210     u059(.A0(men_men_n80_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n82_));
  AOI210     u060(.A0(men_men_n81_), .A1(men_men_n48_), .B0(men_men_n82_), .Y(men_men_n83_));
  NO2        u061(.A(men_men_n36_), .B(x00), .Y(men_men_n84_));
  NO2        u062(.A(x08), .B(x01), .Y(men_men_n85_));
  OAI210     u063(.A0(men_men_n85_), .A1(men_men_n84_), .B0(men_men_n35_), .Y(men_men_n86_));
  NO3        u064(.A(men_men_n86_), .B(men_men_n83_), .C(men_men_n79_), .Y(men_men_n87_));
  AN2        u065(.A(men_men_n87_), .B(men_men_n76_), .Y(men_men_n88_));
  INV        u066(.A(men_men_n86_), .Y(men_men_n89_));
  NO2        u067(.A(x06), .B(x05), .Y(men_men_n90_));
  NA2        u068(.A(x11), .B(x00), .Y(men_men_n91_));
  NO2        u069(.A(x11), .B(men_men_n47_), .Y(men_men_n92_));
  NOi21      u070(.An(men_men_n91_), .B(men_men_n92_), .Y(men_men_n93_));
  NOi21      u071(.An(x01), .B(x10), .Y(men_men_n94_));
  NO2        u072(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n95_));
  NO3        u073(.A(men_men_n95_), .B(men_men_n94_), .C(x06), .Y(men_men_n96_));
  NA2        u074(.A(men_men_n96_), .B(men_men_n27_), .Y(men_men_n97_));
  OAI210     u075(.A0(men_men_n443_), .A1(x07), .B0(men_men_n97_), .Y(men_men_n98_));
  NO3        u076(.A(men_men_n98_), .B(men_men_n88_), .C(men_men_n70_), .Y(men01));
  INV        u077(.A(x12), .Y(men_men_n100_));
  INV        u078(.A(x13), .Y(men_men_n101_));
  NA2        u079(.A(men_men_n90_), .B(x01), .Y(men_men_n102_));
  NA2        u080(.A(men_men_n102_), .B(men_men_n71_), .Y(men_men_n103_));
  NA2        u081(.A(x08), .B(x04), .Y(men_men_n104_));
  NA2        u082(.A(x08), .B(men_men_n103_), .Y(men_men_n105_));
  NA2        u083(.A(men_men_n94_), .B(men_men_n28_), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n72_), .Y(men_men_n107_));
  NO2        u085(.A(x10), .B(x01), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n29_), .B(x00), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n108_), .Y(men_men_n110_));
  NA2        u088(.A(x04), .B(men_men_n28_), .Y(men_men_n111_));
  NO3        u089(.A(men_men_n111_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n112_));
  AOI210     u090(.A0(men_men_n112_), .A1(men_men_n110_), .B0(men_men_n107_), .Y(men_men_n113_));
  AOI210     u091(.A0(men_men_n113_), .A1(men_men_n105_), .B0(men_men_n101_), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n56_), .B(x05), .Y(men_men_n115_));
  NOi21      u093(.An(men_men_n115_), .B(men_men_n58_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n101_), .B(men_men_n36_), .Y(men_men_n117_));
  NA3        u095(.A(men_men_n117_), .B(men_men_n444_), .C(x06), .Y(men_men_n118_));
  INV        u096(.A(men_men_n118_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n85_), .B(x13), .Y(men_men_n120_));
  NA2        u098(.A(x09), .B(men_men_n35_), .Y(men_men_n121_));
  NO2        u099(.A(men_men_n121_), .B(men_men_n120_), .Y(men_men_n122_));
  NA2        u100(.A(x13), .B(men_men_n35_), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n123_), .B(x05), .Y(men_men_n124_));
  NO2        u102(.A(men_men_n124_), .B(men_men_n122_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n126_));
  AOI210     u104(.A0(men_men_n57_), .A1(men_men_n81_), .B0(men_men_n116_), .Y(men_men_n127_));
  AOI210     u105(.A0(men_men_n127_), .A1(men_men_n125_), .B0(men_men_n73_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n129_));
  NA2        u107(.A(x10), .B(men_men_n57_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n130_), .B(men_men_n129_), .Y(men_men_n131_));
  NA2        u109(.A(men_men_n51_), .B(x05), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n36_), .B(x04), .Y(men_men_n133_));
  NA3        u111(.A(men_men_n133_), .B(men_men_n132_), .C(x13), .Y(men_men_n134_));
  NO3        u112(.A(men_men_n126_), .B(men_men_n80_), .C(men_men_n36_), .Y(men_men_n135_));
  NO2        u113(.A(men_men_n60_), .B(x05), .Y(men_men_n136_));
  NOi41      u114(.An(men_men_n134_), .B(men_men_n136_), .C(men_men_n135_), .D(men_men_n131_), .Y(men_men_n137_));
  NO3        u115(.A(men_men_n137_), .B(x06), .C(x03), .Y(men_men_n138_));
  NO4        u116(.A(men_men_n138_), .B(men_men_n128_), .C(men_men_n119_), .D(men_men_n114_), .Y(men_men_n139_));
  NA2        u117(.A(x13), .B(men_men_n36_), .Y(men_men_n140_));
  OAI210     u118(.A0(men_men_n85_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n141_));
  INV        u119(.A(men_men_n140_), .Y(men_men_n142_));
  NO2        u120(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n143_));
  OA210      u121(.A0(x00), .A1(men_men_n78_), .B0(men_men_n143_), .Y(men_men_n144_));
  NO2        u122(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n145_));
  NA2        u123(.A(men_men_n29_), .B(x06), .Y(men_men_n146_));
  AN2        u124(.A(men_men_n144_), .B(men_men_n142_), .Y(men_men_n147_));
  NO2        u125(.A(x09), .B(x05), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n148_), .B(men_men_n47_), .Y(men_men_n149_));
  AOI210     u127(.A0(men_men_n149_), .A1(men_men_n110_), .B0(men_men_n49_), .Y(men_men_n150_));
  NA2        u128(.A(x09), .B(x00), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n115_), .B(men_men_n151_), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n77_), .B(men_men_n51_), .Y(men_men_n153_));
  AOI210     u131(.A0(men_men_n153_), .A1(men_men_n152_), .B0(men_men_n146_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n154_), .B(men_men_n150_), .C(men_men_n147_), .Y(men_men_n155_));
  NO2        u133(.A(x03), .B(x02), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n86_), .B(men_men_n101_), .Y(men_men_n157_));
  OAI210     u135(.A0(men_men_n157_), .A1(men_men_n116_), .B0(men_men_n156_), .Y(men_men_n158_));
  OA210      u136(.A0(men_men_n155_), .A1(x11), .B0(men_men_n158_), .Y(men_men_n159_));
  OAI210     u137(.A0(men_men_n139_), .A1(men_men_n23_), .B0(men_men_n159_), .Y(men_men_n160_));
  NA2        u138(.A(men_men_n110_), .B(men_men_n40_), .Y(men_men_n161_));
  NAi21      u139(.An(x06), .B(x10), .Y(men_men_n162_));
  NOi21      u140(.An(x01), .B(x13), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  OR2        u142(.A(men_men_n164_), .B(x08), .Y(men_men_n165_));
  AOI210     u143(.A0(men_men_n165_), .A1(men_men_n161_), .B0(men_men_n41_), .Y(men_men_n166_));
  NO2        u144(.A(men_men_n29_), .B(x03), .Y(men_men_n167_));
  NA2        u145(.A(men_men_n101_), .B(x01), .Y(men_men_n168_));
  NO2        u146(.A(men_men_n168_), .B(x08), .Y(men_men_n169_));
  OAI210     u147(.A0(x05), .A1(men_men_n169_), .B0(men_men_n51_), .Y(men_men_n170_));
  AOI210     u148(.A0(men_men_n170_), .A1(men_men_n167_), .B0(men_men_n48_), .Y(men_men_n171_));
  AOI210     u149(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n172_));
  OAI210     u150(.A0(men_men_n171_), .A1(men_men_n166_), .B0(men_men_n172_), .Y(men_men_n173_));
  NA2        u151(.A(x04), .B(x02), .Y(men_men_n174_));
  NA2        u152(.A(x10), .B(x05), .Y(men_men_n175_));
  NA2        u153(.A(x09), .B(x06), .Y(men_men_n176_));
  NO2        u154(.A(x09), .B(x01), .Y(men_men_n177_));
  NO3        u155(.A(men_men_n177_), .B(men_men_n108_), .C(men_men_n31_), .Y(men_men_n178_));
  NA2        u156(.A(men_men_n178_), .B(x00), .Y(men_men_n179_));
  NO2        u157(.A(men_men_n115_), .B(x08), .Y(men_men_n180_));
  NA3        u158(.A(men_men_n163_), .B(men_men_n162_), .C(men_men_n51_), .Y(men_men_n181_));
  NA2        u159(.A(men_men_n94_), .B(x05), .Y(men_men_n182_));
  OAI210     u160(.A0(men_men_n182_), .A1(men_men_n117_), .B0(men_men_n181_), .Y(men_men_n183_));
  AOI210     u161(.A0(men_men_n180_), .A1(x06), .B0(men_men_n183_), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(x11), .B0(men_men_n179_), .Y(men_men_n185_));
  NAi21      u163(.An(men_men_n174_), .B(men_men_n185_), .Y(men_men_n186_));
  INV        u164(.A(men_men_n25_), .Y(men_men_n187_));
  NAi21      u165(.An(x13), .B(x00), .Y(men_men_n188_));
  AOI210     u166(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n188_), .Y(men_men_n189_));
  AOI220     u167(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n190_));
  OAI210     u168(.A0(men_men_n175_), .A1(men_men_n35_), .B0(men_men_n190_), .Y(men_men_n191_));
  AN2        u169(.A(men_men_n191_), .B(men_men_n189_), .Y(men_men_n192_));
  NO2        u170(.A(men_men_n188_), .B(men_men_n36_), .Y(men_men_n193_));
  INV        u171(.A(men_men_n193_), .Y(men_men_n194_));
  OAI210     u172(.A0(men_men_n194_), .A1(men_men_n176_), .B0(men_men_n73_), .Y(men_men_n195_));
  OAI210     u173(.A0(men_men_n195_), .A1(men_men_n192_), .B0(men_men_n187_), .Y(men_men_n196_));
  NOi21      u174(.An(x09), .B(x00), .Y(men_men_n197_));
  NO3        u175(.A(men_men_n84_), .B(men_men_n197_), .C(men_men_n47_), .Y(men_men_n198_));
  NA2        u176(.A(men_men_n198_), .B(men_men_n130_), .Y(men_men_n199_));
  NA2        u177(.A(x10), .B(x08), .Y(men_men_n200_));
  INV        u178(.A(men_men_n200_), .Y(men_men_n201_));
  NA2        u179(.A(x06), .B(x05), .Y(men_men_n202_));
  OAI210     u180(.A0(men_men_n202_), .A1(men_men_n35_), .B0(men_men_n100_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n201_), .A1(men_men_n58_), .B0(men_men_n203_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n204_), .B(men_men_n199_), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n101_), .B(x12), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n206_), .Y(men_men_n207_));
  NA2        u185(.A(men_men_n94_), .B(men_men_n51_), .Y(men_men_n208_));
  NO2        u186(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n209_), .B(x02), .Y(men_men_n210_));
  NO2        u188(.A(men_men_n210_), .B(men_men_n208_), .Y(men_men_n211_));
  AOI210     u189(.A0(men_men_n207_), .A1(men_men_n205_), .B0(men_men_n211_), .Y(men_men_n212_));
  NA4        u190(.A(men_men_n212_), .B(men_men_n196_), .C(men_men_n186_), .D(men_men_n173_), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n160_), .A1(men_men_n100_), .B0(men_men_n213_), .Y(men_men_n214_));
  NA2        u192(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n215_));
  NA2        u193(.A(men_men_n215_), .B(men_men_n141_), .Y(men_men_n216_));
  AOI210     u194(.A0(men_men_n30_), .A1(x06), .B0(x05), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n129_), .B(x06), .Y(men_men_n218_));
  AOI210     u196(.A0(men_men_n217_), .A1(men_men_n216_), .B0(men_men_n218_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n219_), .B(x12), .Y(men_men_n220_));
  INV        u198(.A(men_men_n77_), .Y(men_men_n221_));
  NA2        u199(.A(men_men_n164_), .B(men_men_n57_), .Y(men_men_n222_));
  INV        u200(.A(men_men_n222_), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n162_), .B(x02), .Y(men_men_n224_));
  AOI210     u202(.A0(men_men_n224_), .A1(men_men_n223_), .B0(men_men_n23_), .Y(men_men_n225_));
  OAI210     u203(.A0(men_men_n220_), .A1(men_men_n57_), .B0(men_men_n225_), .Y(men_men_n226_));
  INV        u204(.A(men_men_n146_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n51_), .B(x03), .Y(men_men_n228_));
  OAI210     u206(.A0(men_men_n80_), .A1(men_men_n36_), .B0(men_men_n121_), .Y(men_men_n229_));
  NO2        u207(.A(men_men_n101_), .B(x03), .Y(men_men_n230_));
  AOI220     u208(.A0(men_men_n230_), .A1(men_men_n229_), .B0(men_men_n77_), .B1(men_men_n228_), .Y(men_men_n231_));
  NA2        u209(.A(men_men_n32_), .B(x06), .Y(men_men_n232_));
  INV        u210(.A(men_men_n162_), .Y(men_men_n233_));
  NOi21      u211(.An(x13), .B(x04), .Y(men_men_n234_));
  NO3        u212(.A(men_men_n234_), .B(men_men_n77_), .C(men_men_n197_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n235_), .B(x05), .Y(men_men_n236_));
  AOI220     u214(.A0(men_men_n236_), .A1(men_men_n232_), .B0(men_men_n233_), .B1(men_men_n57_), .Y(men_men_n237_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n227_), .B0(men_men_n237_), .Y(men_men_n238_));
  INV        u216(.A(men_men_n92_), .Y(men_men_n239_));
  NO2        u217(.A(men_men_n239_), .B(x12), .Y(men_men_n240_));
  NA2        u218(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n241_));
  NO2        u219(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n242_));
  OAI210     u220(.A0(men_men_n242_), .A1(men_men_n191_), .B0(men_men_n189_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n104_), .A1(men_men_n151_), .B0(men_men_n73_), .Y(men_men_n244_));
  INV        u222(.A(men_men_n244_), .Y(men_men_n245_));
  NA2        u223(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n246_));
  INV        u224(.A(x03), .Y(men_men_n247_));
  OA210      u225(.A0(men_men_n247_), .A1(men_men_n245_), .B0(men_men_n243_), .Y(men_men_n248_));
  NA2        u226(.A(x13), .B(men_men_n100_), .Y(men_men_n249_));
  NA3        u227(.A(men_men_n249_), .B(men_men_n203_), .C(men_men_n93_), .Y(men_men_n250_));
  OAI210     u228(.A0(men_men_n248_), .A1(men_men_n241_), .B0(men_men_n250_), .Y(men_men_n251_));
  AOI210     u229(.A0(men_men_n240_), .A1(men_men_n238_), .B0(men_men_n251_), .Y(men_men_n252_));
  AOI210     u230(.A0(men_men_n252_), .A1(men_men_n226_), .B0(x07), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n72_), .B(men_men_n29_), .Y(men_men_n254_));
  AOI210     u232(.A0(men_men_n140_), .A1(men_men_n153_), .B0(men_men_n254_), .Y(men_men_n255_));
  NO2        u233(.A(men_men_n101_), .B(x06), .Y(men_men_n256_));
  INV        u234(.A(men_men_n256_), .Y(men_men_n257_));
  NO2        u235(.A(x08), .B(x05), .Y(men_men_n258_));
  OAI210     u236(.A0(men_men_n77_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n259_));
  NA2        u237(.A(men_men_n257_), .B(men_men_n259_), .Y(men_men_n260_));
  NO2        u238(.A(x12), .B(x02), .Y(men_men_n261_));
  INV        u239(.A(men_men_n261_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n262_), .B(men_men_n239_), .Y(men_men_n263_));
  OA210      u241(.A0(men_men_n260_), .A1(men_men_n255_), .B0(men_men_n263_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n265_), .B(x01), .Y(men_men_n266_));
  NOi21      u244(.An(men_men_n85_), .B(men_men_n121_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n267_), .B(men_men_n266_), .Y(men_men_n268_));
  AOI210     u246(.A0(men_men_n268_), .A1(men_men_n134_), .B0(men_men_n29_), .Y(men_men_n269_));
  NA2        u247(.A(men_men_n256_), .B(men_men_n229_), .Y(men_men_n270_));
  NA2        u248(.A(men_men_n101_), .B(x04), .Y(men_men_n271_));
  NA2        u249(.A(men_men_n271_), .B(men_men_n28_), .Y(men_men_n272_));
  OAI210     u250(.A0(men_men_n272_), .A1(men_men_n120_), .B0(men_men_n270_), .Y(men_men_n273_));
  NO3        u251(.A(men_men_n91_), .B(x12), .C(x03), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n273_), .A1(men_men_n269_), .B0(men_men_n274_), .Y(men_men_n275_));
  AOI210     u253(.A0(men_men_n208_), .A1(men_men_n202_), .B0(men_men_n104_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n25_), .B(x00), .Y(men_men_n277_));
  NA2        u255(.A(men_men_n276_), .B(men_men_n277_), .Y(men_men_n278_));
  NO2        u256(.A(men_men_n241_), .B(men_men_n28_), .Y(men_men_n279_));
  NA2        u257(.A(men_men_n227_), .B(men_men_n279_), .Y(men_men_n280_));
  NA3        u258(.A(men_men_n280_), .B(men_men_n278_), .C(men_men_n275_), .Y(men_men_n281_));
  NO3        u259(.A(men_men_n281_), .B(men_men_n264_), .C(men_men_n253_), .Y(men_men_n282_));
  OAI210     u260(.A0(men_men_n214_), .A1(men_men_n61_), .B0(men_men_n282_), .Y(men02));
  AOI210     u261(.A0(men_men_n140_), .A1(men_men_n86_), .B0(men_men_n132_), .Y(men_men_n284_));
  BUFFER     u262(.A(men_men_n235_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n101_), .B(men_men_n35_), .Y(men_men_n286_));
  NA3        u264(.A(men_men_n286_), .B(men_men_n201_), .C(men_men_n56_), .Y(men_men_n287_));
  OAI210     u265(.A0(men_men_n285_), .A1(men_men_n32_), .B0(men_men_n287_), .Y(men_men_n288_));
  OAI210     u266(.A0(men_men_n288_), .A1(men_men_n284_), .B0(men_men_n175_), .Y(men_men_n289_));
  INV        u267(.A(men_men_n175_), .Y(men_men_n290_));
  NO2        u268(.A(men_men_n86_), .B(men_men_n51_), .Y(men_men_n291_));
  AOI220     u269(.A0(men_men_n291_), .A1(men_men_n290_), .B0(men_men_n157_), .B1(men_men_n156_), .Y(men_men_n292_));
  AOI210     u270(.A0(men_men_n292_), .A1(men_men_n289_), .B0(men_men_n48_), .Y(men_men_n293_));
  NO2        u271(.A(x05), .B(x02), .Y(men_men_n294_));
  OAI210     u272(.A0(men_men_n216_), .A1(men_men_n197_), .B0(men_men_n294_), .Y(men_men_n295_));
  AOI220     u273(.A0(men_men_n258_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n296_));
  NOi21      u274(.An(men_men_n286_), .B(men_men_n296_), .Y(men_men_n297_));
  AOI210     u275(.A0(men_men_n234_), .A1(men_men_n80_), .B0(men_men_n297_), .Y(men_men_n298_));
  AOI210     u276(.A0(men_men_n298_), .A1(men_men_n295_), .B0(men_men_n146_), .Y(men_men_n299_));
  NAi21      u277(.An(men_men_n236_), .B(men_men_n231_), .Y(men_men_n300_));
  NO2        u278(.A(men_men_n246_), .B(men_men_n47_), .Y(men_men_n301_));
  NA2        u279(.A(men_men_n301_), .B(men_men_n300_), .Y(men_men_n302_));
  AN2        u280(.A(men_men_n230_), .B(men_men_n229_), .Y(men_men_n303_));
  OAI210     u281(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n304_));
  NA2        u282(.A(x13), .B(men_men_n28_), .Y(men_men_n305_));
  BUFFER     u283(.A(men_men_n149_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n306_), .A1(men_men_n141_), .B0(men_men_n304_), .Y(men_men_n307_));
  OAI210     u285(.A0(men_men_n307_), .A1(men_men_n303_), .B0(men_men_n95_), .Y(men_men_n308_));
  NA3        u286(.A(men_men_n95_), .B(men_men_n85_), .C(men_men_n228_), .Y(men_men_n309_));
  NA3        u287(.A(men_men_n94_), .B(men_men_n84_), .C(men_men_n42_), .Y(men_men_n310_));
  AOI210     u288(.A0(men_men_n310_), .A1(men_men_n309_), .B0(x04), .Y(men_men_n311_));
  INV        u289(.A(men_men_n156_), .Y(men_men_n312_));
  NO2        u290(.A(men_men_n312_), .B(men_men_n131_), .Y(men_men_n313_));
  AOI210     u291(.A0(men_men_n313_), .A1(x13), .B0(men_men_n311_), .Y(men_men_n314_));
  NA3        u292(.A(men_men_n314_), .B(men_men_n308_), .C(men_men_n302_), .Y(men_men_n315_));
  NO3        u293(.A(men_men_n315_), .B(men_men_n299_), .C(men_men_n293_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n145_), .B(x03), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n188_), .A1(men_men_n51_), .B0(men_men_n317_), .Y(men_men_n318_));
  NA2        u296(.A(men_men_n318_), .B(men_men_n108_), .Y(men_men_n319_));
  INV        u297(.A(men_men_n56_), .Y(men_men_n320_));
  OAI220     u298(.A0(men_men_n271_), .A1(men_men_n320_), .B0(men_men_n132_), .B1(men_men_n28_), .Y(men_men_n321_));
  OAI210     u299(.A0(men_men_n321_), .A1(men_men_n180_), .B0(men_men_n109_), .Y(men_men_n322_));
  NA2        u300(.A(men_men_n271_), .B(men_men_n100_), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n100_), .B(men_men_n41_), .Y(men_men_n324_));
  NA3        u302(.A(men_men_n324_), .B(men_men_n323_), .C(men_men_n131_), .Y(men_men_n325_));
  NA4        u303(.A(men_men_n325_), .B(men_men_n322_), .C(men_men_n319_), .D(men_men_n48_), .Y(men_men_n326_));
  INV        u304(.A(men_men_n209_), .Y(men_men_n327_));
  NO2        u305(.A(men_men_n169_), .B(men_men_n40_), .Y(men_men_n328_));
  NA2        u306(.A(men_men_n32_), .B(x05), .Y(men_men_n329_));
  OAI220     u307(.A0(men_men_n329_), .A1(men_men_n328_), .B0(men_men_n327_), .B1(men_men_n59_), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(x02), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n206_), .B(x04), .Y(men_men_n332_));
  NO2        u310(.A(men_men_n332_), .B(men_men_n36_), .Y(men_men_n333_));
  NO3        u311(.A(men_men_n190_), .B(x13), .C(men_men_n31_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n334_), .A1(men_men_n333_), .B0(men_men_n95_), .Y(men_men_n335_));
  NO3        u313(.A(men_men_n206_), .B(men_men_n167_), .C(men_men_n52_), .Y(men_men_n336_));
  OAI210     u314(.A0(x12), .A1(men_men_n198_), .B0(men_men_n336_), .Y(men_men_n337_));
  NA4        u315(.A(men_men_n337_), .B(men_men_n335_), .C(men_men_n331_), .D(x06), .Y(men_men_n338_));
  NA2        u316(.A(x09), .B(x03), .Y(men_men_n339_));
  OAI220     u317(.A0(men_men_n339_), .A1(men_men_n130_), .B0(men_men_n215_), .B1(men_men_n64_), .Y(men_men_n340_));
  OAI220     u318(.A0(men_men_n168_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n341_), .B(men_men_n227_), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n343_));
  NA2        u321(.A(men_men_n336_), .B(men_men_n343_), .Y(men_men_n344_));
  OAI210     u322(.A0(men_men_n342_), .A1(men_men_n28_), .B0(men_men_n344_), .Y(men_men_n345_));
  AO220      u323(.A0(men_men_n345_), .A1(x04), .B0(men_men_n340_), .B1(x05), .Y(men_men_n346_));
  AOI210     u324(.A0(men_men_n338_), .A1(men_men_n326_), .B0(men_men_n346_), .Y(men_men_n347_));
  OAI210     u325(.A0(men_men_n316_), .A1(x12), .B0(men_men_n347_), .Y(men03));
  OR2        u326(.A(men_men_n42_), .B(men_men_n228_), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n157_), .A1(men_men_n100_), .B0(men_men_n349_), .Y(men_men_n350_));
  NA2        u328(.A(men_men_n206_), .B(men_men_n156_), .Y(men_men_n351_));
  NA2        u329(.A(men_men_n351_), .B(men_men_n210_), .Y(men_men_n352_));
  OAI210     u330(.A0(men_men_n352_), .A1(men_men_n350_), .B0(x05), .Y(men_men_n353_));
  NA2        u331(.A(men_men_n349_), .B(x05), .Y(men_men_n354_));
  AOI210     u332(.A0(men_men_n141_), .A1(men_men_n221_), .B0(men_men_n354_), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n230_), .A1(men_men_n81_), .B0(men_men_n124_), .Y(men_men_n356_));
  OAI220     u334(.A0(men_men_n356_), .A1(men_men_n59_), .B0(men_men_n305_), .B1(men_men_n296_), .Y(men_men_n357_));
  OAI210     u335(.A0(men_men_n357_), .A1(men_men_n355_), .B0(men_men_n100_), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n149_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n359_));
  NO2        u337(.A(men_men_n177_), .B(men_men_n136_), .Y(men_men_n360_));
  OAI220     u338(.A0(men_men_n360_), .A1(men_men_n37_), .B0(men_men_n152_), .B1(x13), .Y(men_men_n361_));
  OAI210     u339(.A0(men_men_n361_), .A1(men_men_n359_), .B0(x04), .Y(men_men_n362_));
  NO3        u340(.A(men_men_n324_), .B(men_men_n86_), .C(men_men_n59_), .Y(men_men_n363_));
  AOI210     u341(.A0(men_men_n194_), .A1(men_men_n100_), .B0(men_men_n149_), .Y(men_men_n364_));
  OA210      u342(.A0(men_men_n169_), .A1(x12), .B0(men_men_n136_), .Y(men_men_n365_));
  NO3        u343(.A(men_men_n365_), .B(men_men_n364_), .C(men_men_n363_), .Y(men_men_n366_));
  NA4        u344(.A(men_men_n366_), .B(men_men_n362_), .C(men_men_n358_), .D(men_men_n353_), .Y(men04));
  NO2        u345(.A(men_men_n89_), .B(men_men_n39_), .Y(men_men_n368_));
  XO2        u346(.A(men_men_n368_), .B(men_men_n249_), .Y(men05));
  AOI210     u347(.A0(men_men_n72_), .A1(men_men_n52_), .B0(men_men_n218_), .Y(men_men_n370_));
  NO2        u348(.A(men_men_n370_), .B(men_men_n25_), .Y(men_men_n371_));
  AOI210     u349(.A0(men_men_n233_), .A1(men_men_n57_), .B0(men_men_n90_), .Y(men_men_n372_));
  NO2        u350(.A(men_men_n372_), .B(men_men_n24_), .Y(men_men_n373_));
  OAI210     u351(.A0(men_men_n373_), .A1(men_men_n371_), .B0(men_men_n100_), .Y(men_men_n374_));
  NA2        u352(.A(x11), .B(men_men_n31_), .Y(men_men_n375_));
  NA2        u353(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n376_));
  NA2        u354(.A(men_men_n254_), .B(x03), .Y(men_men_n377_));
  OAI220     u355(.A0(men_men_n377_), .A1(men_men_n376_), .B0(men_men_n375_), .B1(men_men_n82_), .Y(men_men_n378_));
  OAI210     u356(.A0(men_men_n26_), .A1(men_men_n100_), .B0(x07), .Y(men_men_n379_));
  AOI210     u357(.A0(men_men_n378_), .A1(x06), .B0(men_men_n379_), .Y(men_men_n380_));
  AOI220     u358(.A0(men_men_n82_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n381_));
  NO3        u359(.A(men_men_n381_), .B(men_men_n23_), .C(x00), .Y(men_men_n382_));
  NA2        u360(.A(men_men_n71_), .B(x02), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n383_), .A1(men_men_n377_), .B0(men_men_n256_), .Y(men_men_n384_));
  OR2        u362(.A(men_men_n384_), .B(men_men_n241_), .Y(men_men_n385_));
  NO2        u363(.A(men_men_n23_), .B(x10), .Y(men_men_n386_));
  OAI210     u364(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n387_));
  OR3        u365(.A(men_men_n387_), .B(men_men_n386_), .C(men_men_n44_), .Y(men_men_n388_));
  NA2        u366(.A(men_men_n388_), .B(men_men_n385_), .Y(men_men_n389_));
  OAI210     u367(.A0(men_men_n389_), .A1(men_men_n382_), .B0(men_men_n100_), .Y(men_men_n390_));
  NA2        u368(.A(men_men_n33_), .B(men_men_n100_), .Y(men_men_n391_));
  AOI210     u369(.A0(men_men_n391_), .A1(men_men_n92_), .B0(x07), .Y(men_men_n392_));
  AOI220     u370(.A0(men_men_n392_), .A1(men_men_n390_), .B0(men_men_n380_), .B1(men_men_n374_), .Y(men_men_n393_));
  NA3        u371(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n394_));
  AO210      u372(.A0(men_men_n394_), .A1(men_men_n265_), .B0(men_men_n262_), .Y(men_men_n395_));
  AOI210     u373(.A0(men_men_n386_), .A1(men_men_n75_), .B0(men_men_n145_), .Y(men_men_n396_));
  OR2        u374(.A(men_men_n396_), .B(x03), .Y(men_men_n397_));
  NA2        u375(.A(men_men_n343_), .B(men_men_n61_), .Y(men_men_n398_));
  NO2        u376(.A(men_men_n398_), .B(x11), .Y(men_men_n399_));
  NO3        u377(.A(men_men_n399_), .B(men_men_n148_), .C(men_men_n28_), .Y(men_men_n400_));
  AOI220     u378(.A0(men_men_n400_), .A1(men_men_n397_), .B0(men_men_n395_), .B1(men_men_n47_), .Y(men_men_n401_));
  NO4        u379(.A(men_men_n324_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n402_));
  OAI210     u380(.A0(men_men_n402_), .A1(men_men_n401_), .B0(men_men_n101_), .Y(men_men_n403_));
  AOI210     u381(.A0(men_men_n332_), .A1(men_men_n111_), .B0(men_men_n261_), .Y(men_men_n404_));
  NOi21      u382(.An(men_men_n317_), .B(men_men_n136_), .Y(men_men_n405_));
  OAI210     u383(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n406_));
  AOI210     u384(.A0(men_men_n249_), .A1(men_men_n47_), .B0(men_men_n406_), .Y(men_men_n407_));
  NO3        u385(.A(men_men_n407_), .B(men_men_n404_), .C(x08), .Y(men_men_n408_));
  AOI210     u386(.A0(men_men_n386_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n409_));
  NA2        u387(.A(x09), .B(men_men_n41_), .Y(men_men_n410_));
  OAI220     u388(.A0(men_men_n410_), .A1(men_men_n409_), .B0(men_men_n375_), .B1(men_men_n67_), .Y(men_men_n411_));
  NO2        u389(.A(x13), .B(x12), .Y(men_men_n412_));
  NO2        u390(.A(men_men_n132_), .B(men_men_n28_), .Y(men_men_n413_));
  NO2        u391(.A(men_men_n413_), .B(men_men_n266_), .Y(men_men_n414_));
  OR3        u392(.A(men_men_n414_), .B(x12), .C(x03), .Y(men_men_n415_));
  NA3        u393(.A(men_men_n327_), .B(men_men_n126_), .C(x12), .Y(men_men_n416_));
  AO210      u394(.A0(men_men_n327_), .A1(men_men_n126_), .B0(men_men_n249_), .Y(men_men_n417_));
  NA4        u395(.A(men_men_n417_), .B(men_men_n416_), .C(men_men_n415_), .D(x08), .Y(men_men_n418_));
  AOI210     u396(.A0(men_men_n412_), .A1(men_men_n411_), .B0(men_men_n418_), .Y(men_men_n419_));
  AOI210     u397(.A0(men_men_n408_), .A1(men_men_n403_), .B0(men_men_n419_), .Y(men_men_n420_));
  OAI210     u398(.A0(men_men_n398_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n421_));
  NA2        u399(.A(men_men_n290_), .B(x07), .Y(men_men_n422_));
  OAI220     u400(.A0(men_men_n422_), .A1(men_men_n376_), .B0(men_men_n148_), .B1(men_men_n43_), .Y(men_men_n423_));
  OAI210     u401(.A0(men_men_n423_), .A1(men_men_n421_), .B0(men_men_n193_), .Y(men_men_n424_));
  NA3        u402(.A(men_men_n414_), .B(men_men_n405_), .C(men_men_n323_), .Y(men_men_n425_));
  INV        u403(.A(x14), .Y(men_men_n426_));
  NO3        u404(.A(men_men_n317_), .B(men_men_n106_), .C(x11), .Y(men_men_n427_));
  NO3        u405(.A(men_men_n168_), .B(men_men_n75_), .C(men_men_n57_), .Y(men_men_n428_));
  NO3        u406(.A(men_men_n394_), .B(men_men_n324_), .C(men_men_n188_), .Y(men_men_n429_));
  NO4        u407(.A(men_men_n429_), .B(men_men_n428_), .C(men_men_n427_), .D(men_men_n426_), .Y(men_men_n430_));
  NA3        u408(.A(men_men_n430_), .B(men_men_n425_), .C(men_men_n424_), .Y(men_men_n431_));
  AOI220     u409(.A0(men_men_n391_), .A1(men_men_n61_), .B0(men_men_n413_), .B1(men_men_n167_), .Y(men_men_n432_));
  NOi21      u410(.An(men_men_n271_), .B(men_men_n152_), .Y(men_men_n433_));
  NO3        u411(.A(men_men_n129_), .B(men_men_n24_), .C(x06), .Y(men_men_n434_));
  AOI210     u412(.A0(men_men_n277_), .A1(men_men_n233_), .B0(men_men_n434_), .Y(men_men_n435_));
  OAI210     u413(.A0(men_men_n44_), .A1(x04), .B0(men_men_n435_), .Y(men_men_n436_));
  OAI210     u414(.A0(men_men_n436_), .A1(men_men_n433_), .B0(men_men_n100_), .Y(men_men_n437_));
  OAI210     u415(.A0(men_men_n432_), .A1(men_men_n91_), .B0(men_men_n437_), .Y(men_men_n438_));
  NO4        u416(.A(men_men_n438_), .B(men_men_n431_), .C(men_men_n420_), .D(men_men_n393_), .Y(men06));
  INV        u417(.A(x07), .Y(men_men_n442_));
  INV        u418(.A(men_men_n93_), .Y(men_men_n443_));
  INV        u419(.A(x02), .Y(men_men_n444_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule