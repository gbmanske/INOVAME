//Benchmark atmr_alu4_1266_0.25

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n117_, ori_ori_n118_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n132_, men_men_n133_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  INV        o019(.A(ori_ori_n35_), .Y(ori1));
  INV        o020(.A(i_11_), .Y(ori_ori_n43_));
  NO2        o021(.A(ori_ori_n43_), .B(i_6_), .Y(ori_ori_n44_));
  INV        o022(.A(i_2_), .Y(ori_ori_n45_));
  NA2        o023(.A(i_0_), .B(i_3_), .Y(ori_ori_n46_));
  INV        o024(.A(i_5_), .Y(ori_ori_n47_));
  NO2        o025(.A(i_7_), .B(i_10_), .Y(ori_ori_n48_));
  AOI210     o026(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n48_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_5_), .A1(ori_ori_n46_), .B0(ori_ori_n45_), .Y(ori_ori_n50_));
  NA2        o028(.A(i_0_), .B(i_2_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_7_), .B(i_9_), .Y(ori_ori_n52_));
  NO2        o030(.A(ori_ori_n52_), .B(ori_ori_n51_), .Y(ori_ori_n53_));
  NA2        o031(.A(ori_ori_n50_), .B(ori_ori_n44_), .Y(ori_ori_n54_));
  NA3        o032(.A(i_2_), .B(i_6_), .C(i_8_), .Y(ori_ori_n55_));
  NO2        o033(.A(i_1_), .B(i_6_), .Y(ori_ori_n56_));
  NA2        o034(.A(i_8_), .B(i_7_), .Y(ori_ori_n57_));
  OAI210     o035(.A0(ori_ori_n57_), .A1(ori_ori_n56_), .B0(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n58_), .B(i_12_), .Y(ori_ori_n59_));
  NAi21      o037(.An(i_2_), .B(i_7_), .Y(ori_ori_n60_));
  INV        o038(.A(i_1_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n61_), .B(i_6_), .Y(ori_ori_n62_));
  NA3        o040(.A(ori_ori_n62_), .B(ori_ori_n60_), .C(ori_ori_n31_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_1_), .B(i_10_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(i_6_), .Y(ori_ori_n65_));
  NAi31      o043(.An(ori_ori_n65_), .B(ori_ori_n63_), .C(ori_ori_n59_), .Y(ori_ori_n66_));
  NA2        o044(.A(ori_ori_n49_), .B(i_2_), .Y(ori_ori_n67_));
  AOI210     o045(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n68_));
  NA2        o046(.A(i_1_), .B(i_6_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n69_), .B(ori_ori_n25_), .Y(ori_ori_n70_));
  INV        o048(.A(i_0_), .Y(ori_ori_n71_));
  NAi21      o049(.An(i_5_), .B(i_10_), .Y(ori_ori_n72_));
  NA2        o050(.A(i_5_), .B(i_9_), .Y(ori_ori_n73_));
  AOI210     o051(.A0(ori_ori_n73_), .A1(ori_ori_n72_), .B0(ori_ori_n71_), .Y(ori_ori_n74_));
  NO2        o052(.A(ori_ori_n74_), .B(ori_ori_n70_), .Y(ori_ori_n75_));
  INV        o053(.A(ori_ori_n75_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n76_), .A1(ori_ori_n66_), .B0(i_0_), .Y(ori_ori_n77_));
  NA2        o055(.A(i_12_), .B(i_5_), .Y(ori_ori_n78_));
  NO2        o056(.A(i_3_), .B(i_7_), .Y(ori_ori_n79_));
  INV        o057(.A(i_6_), .Y(ori_ori_n80_));
  NO2        o058(.A(i_2_), .B(i_7_), .Y(ori_ori_n81_));
  INV        o059(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  OAI210     o060(.A0(i_1_), .A1(i_6_), .B0(ori_ori_n82_), .Y(ori_ori_n83_));
  NAi21      o061(.An(i_6_), .B(i_10_), .Y(ori_ori_n84_));
  NA2        o062(.A(i_6_), .B(i_9_), .Y(ori_ori_n85_));
  AOI210     o063(.A0(ori_ori_n85_), .A1(ori_ori_n84_), .B0(ori_ori_n61_), .Y(ori_ori_n86_));
  NA2        o064(.A(i_2_), .B(i_6_), .Y(ori_ori_n87_));
  INV        o065(.A(ori_ori_n86_), .Y(ori_ori_n88_));
  AOI210     o066(.A0(ori_ori_n88_), .A1(ori_ori_n83_), .B0(ori_ori_n78_), .Y(ori_ori_n89_));
  AN3        o067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n90_));
  NAi21      o068(.An(i_6_), .B(i_11_), .Y(ori_ori_n91_));
  INV        o069(.A(i_7_), .Y(ori_ori_n92_));
  NO2        o070(.A(i_0_), .B(i_5_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(ori_ori_n80_), .Y(ori_ori_n94_));
  NA2        o072(.A(i_12_), .B(i_3_), .Y(ori_ori_n95_));
  NAi21      o073(.An(i_7_), .B(i_11_), .Y(ori_ori_n96_));
  NO3        o074(.A(ori_ori_n96_), .B(ori_ori_n84_), .C(ori_ori_n51_), .Y(ori_ori_n97_));
  AN2        o075(.A(i_2_), .B(i_10_), .Y(ori_ori_n98_));
  NA2        o076(.A(i_12_), .B(i_7_), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n61_), .B(ori_ori_n26_), .Y(ori_ori_n100_));
  NA2        o078(.A(i_11_), .B(i_12_), .Y(ori_ori_n101_));
  NAi21      o079(.An(ori_ori_n97_), .B(ori_ori_n101_), .Y(ori_ori_n102_));
  NOi21      o080(.An(i_1_), .B(i_5_), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n103_), .B(i_11_), .Y(ori_ori_n104_));
  NA2        o082(.A(ori_ori_n92_), .B(ori_ori_n37_), .Y(ori_ori_n105_));
  NA2        o083(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n106_), .B(ori_ori_n105_), .Y(ori_ori_n107_));
  NO2        o085(.A(ori_ori_n107_), .B(ori_ori_n45_), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n109_));
  NO2        o087(.A(i_1_), .B(ori_ori_n80_), .Y(ori_ori_n110_));
  NO2        o088(.A(i_6_), .B(i_5_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n111_), .B(i_3_), .Y(ori_ori_n112_));
  AO210      o090(.A0(ori_ori_n112_), .A1(ori_ori_n46_), .B0(ori_ori_n110_), .Y(ori_ori_n113_));
  OAI210     o091(.A0(ori_ori_n113_), .A1(ori_ori_n96_), .B0(ori_ori_n104_), .Y(ori_ori_n114_));
  NO3        o092(.A(ori_ori_n114_), .B(ori_ori_n102_), .C(ori_ori_n89_), .Y(ori_ori_n115_));
  NA3        o093(.A(ori_ori_n115_), .B(ori_ori_n77_), .C(ori_ori_n54_), .Y(ori2));
  NO2        o094(.A(ori_ori_n61_), .B(ori_ori_n37_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n576_), .B(ori_ori_n117_), .Y(ori_ori_n118_));
  NA4        o096(.A(ori_ori_n118_), .B(ori_ori_n75_), .C(ori_ori_n67_), .D(ori_ori_n30_), .Y(ori0));
  NAi21      o097(.An(i_5_), .B(i_11_), .Y(ori_ori_n120_));
  NO2        o098(.A(i_0_), .B(i_1_), .Y(ori_ori_n121_));
  NA2        o099(.A(i_1_), .B(i_5_), .Y(ori_ori_n122_));
  NOi21      o100(.An(i_4_), .B(i_10_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(ori_ori_n40_), .Y(ori_ori_n124_));
  NOi21      o102(.An(i_4_), .B(i_9_), .Y(ori_ori_n125_));
  NOi21      o103(.An(i_11_), .B(i_13_), .Y(ori_ori_n126_));
  NA2        o104(.A(ori_ori_n126_), .B(ori_ori_n125_), .Y(ori_ori_n127_));
  NAi21      o105(.An(i_12_), .B(i_11_), .Y(ori_ori_n128_));
  NO2        o106(.A(ori_ori_n71_), .B(i_5_), .Y(ori_ori_n129_));
  NO2        o107(.A(i_2_), .B(i_1_), .Y(ori_ori_n130_));
  NAi21      o108(.An(i_4_), .B(i_12_), .Y(ori_ori_n131_));
  INV        o109(.A(i_8_), .Y(ori_ori_n132_));
  NO3        o110(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n133_));
  NO2        o111(.A(i_3_), .B(i_8_), .Y(ori_ori_n134_));
  NO3        o112(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n93_), .B(ori_ori_n56_), .Y(ori_ori_n136_));
  NO2        o114(.A(i_13_), .B(i_9_), .Y(ori_ori_n137_));
  NAi21      o115(.An(i_12_), .B(i_3_), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n43_), .B(i_5_), .Y(ori_ori_n139_));
  NA3        o117(.A(i_13_), .B(ori_ori_n132_), .C(i_10_), .Y(ori_ori_n140_));
  NA2        o118(.A(i_0_), .B(i_5_), .Y(ori_ori_n141_));
  NAi31      o119(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n142_));
  NO2        o120(.A(ori_ori_n71_), .B(ori_ori_n26_), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n45_), .B(ori_ori_n61_), .Y(ori_ori_n144_));
  INV        o122(.A(i_13_), .Y(ori_ori_n145_));
  NO2        o123(.A(i_12_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NO2        o124(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n147_));
  INV        o125(.A(i_12_), .Y(ori_ori_n148_));
  NO3        o126(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n149_));
  NA2        o127(.A(i_2_), .B(i_1_), .Y(ori_ori_n150_));
  NO3        o128(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n151_));
  NAi21      o129(.An(i_4_), .B(i_3_), .Y(ori_ori_n152_));
  NO2        o130(.A(i_0_), .B(i_6_), .Y(ori_ori_n153_));
  NOi41      o131(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n154_));
  NO2        o132(.A(i_11_), .B(ori_ori_n145_), .Y(ori_ori_n155_));
  NOi21      o133(.An(i_1_), .B(i_6_), .Y(ori_ori_n156_));
  NAi21      o134(.An(i_3_), .B(i_7_), .Y(ori_ori_n157_));
  NA2        o135(.A(ori_ori_n148_), .B(i_9_), .Y(ori_ori_n158_));
  OR4        o136(.A(ori_ori_n158_), .B(ori_ori_n157_), .C(ori_ori_n156_), .D(ori_ori_n129_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n71_), .B(i_5_), .Y(ori_ori_n160_));
  NA2        o138(.A(i_3_), .B(i_9_), .Y(ori_ori_n161_));
  NAi21      o139(.An(i_7_), .B(i_10_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n162_), .B(ori_ori_n161_), .Y(ori_ori_n163_));
  NA3        o141(.A(ori_ori_n163_), .B(ori_ori_n160_), .C(ori_ori_n62_), .Y(ori_ori_n164_));
  NA2        o142(.A(ori_ori_n164_), .B(ori_ori_n159_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n165_), .B(ori_ori_n155_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n152_), .B(i_2_), .Y(ori_ori_n167_));
  NA2        o145(.A(ori_ori_n155_), .B(i_9_), .Y(ori_ori_n168_));
  NO3        o146(.A(i_11_), .B(ori_ori_n145_), .C(ori_ori_n25_), .Y(ori_ori_n169_));
  NO3        o147(.A(i_12_), .B(ori_ori_n145_), .C(ori_ori_n37_), .Y(ori_ori_n170_));
  AN2        o148(.A(i_3_), .B(i_10_), .Y(ori_ori_n171_));
  NO2        o149(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n172_));
  NO3        o150(.A(ori_ori_n43_), .B(i_13_), .C(i_9_), .Y(ori_ori_n173_));
  NO2        o151(.A(i_2_), .B(i_3_), .Y(ori_ori_n174_));
  OR2        o152(.A(i_0_), .B(i_5_), .Y(ori_ori_n175_));
  NO2        o153(.A(i_12_), .B(i_10_), .Y(ori_ori_n176_));
  NOi21      o154(.An(i_5_), .B(i_0_), .Y(ori_ori_n177_));
  NO2        o155(.A(i_1_), .B(i_7_), .Y(ori_ori_n178_));
  NOi21      o156(.An(ori_ori_n122_), .B(ori_ori_n94_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n179_), .B(ori_ori_n106_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n180_), .B(i_3_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n132_), .B(i_9_), .Y(ori_ori_n182_));
  NA2        o160(.A(ori_ori_n182_), .B(ori_ori_n136_), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n183_), .B(ori_ori_n45_), .Y(ori_ori_n184_));
  INV        o162(.A(ori_ori_n184_), .Y(ori_ori_n185_));
  AOI210     o163(.A0(ori_ori_n185_), .A1(ori_ori_n181_), .B0(ori_ori_n124_), .Y(ori_ori_n186_));
  INV        o164(.A(ori_ori_n186_), .Y(ori_ori_n187_));
  NOi32      o165(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n188_));
  INV        o166(.A(ori_ori_n188_), .Y(ori_ori_n189_));
  NOi32      o167(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n190_));
  NAi21      o168(.An(i_6_), .B(i_1_), .Y(ori_ori_n191_));
  NA3        o169(.A(ori_ori_n191_), .B(ori_ori_n190_), .C(ori_ori_n45_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n192_), .B(i_0_), .Y(ori_ori_n193_));
  NO2        o171(.A(i_1_), .B(ori_ori_n92_), .Y(ori_ori_n194_));
  NAi21      o172(.An(i_3_), .B(i_4_), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n195_), .B(i_9_), .Y(ori_ori_n196_));
  AN2        o174(.A(i_6_), .B(i_7_), .Y(ori_ori_n197_));
  OAI210     o175(.A0(ori_ori_n197_), .A1(ori_ori_n194_), .B0(ori_ori_n196_), .Y(ori_ori_n198_));
  NA2        o176(.A(i_2_), .B(i_7_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n195_), .B(i_10_), .Y(ori_ori_n200_));
  NA3        o178(.A(ori_ori_n200_), .B(ori_ori_n199_), .C(ori_ori_n153_), .Y(ori_ori_n201_));
  AOI210     o179(.A0(ori_ori_n201_), .A1(ori_ori_n198_), .B0(ori_ori_n129_), .Y(ori_ori_n202_));
  AOI210     o180(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n203_));
  OAI210     o181(.A0(ori_ori_n203_), .A1(ori_ori_n130_), .B0(ori_ori_n200_), .Y(ori_ori_n204_));
  AOI220     o182(.A0(ori_ori_n200_), .A1(ori_ori_n178_), .B0(ori_ori_n149_), .B1(ori_ori_n130_), .Y(ori_ori_n205_));
  AOI210     o183(.A0(ori_ori_n205_), .A1(ori_ori_n204_), .B0(i_5_), .Y(ori_ori_n206_));
  NO3        o184(.A(ori_ori_n206_), .B(ori_ori_n202_), .C(ori_ori_n193_), .Y(ori_ori_n207_));
  NO2        o185(.A(ori_ori_n207_), .B(ori_ori_n189_), .Y(ori_ori_n208_));
  AN2        o186(.A(i_12_), .B(i_5_), .Y(ori_ori_n209_));
  INV        o187(.A(ori_ori_n209_), .Y(ori_ori_n210_));
  NO2        o188(.A(i_11_), .B(i_6_), .Y(ori_ori_n211_));
  NO2        o189(.A(i_5_), .B(i_10_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_11_), .B(i_12_), .Y(ori_ori_n213_));
  NAi21      o191(.An(i_13_), .B(i_0_), .Y(ori_ori_n214_));
  NO3        o192(.A(i_1_), .B(i_12_), .C(ori_ori_n80_), .Y(ori_ori_n215_));
  NO2        o193(.A(i_0_), .B(i_11_), .Y(ori_ori_n216_));
  AN2        o194(.A(i_1_), .B(i_6_), .Y(ori_ori_n217_));
  NOi21      o195(.An(i_2_), .B(i_12_), .Y(ori_ori_n218_));
  NAi21      o196(.An(i_9_), .B(i_4_), .Y(ori_ori_n219_));
  OR2        o197(.A(i_13_), .B(i_10_), .Y(ori_ori_n220_));
  NO3        o198(.A(ori_ori_n220_), .B(ori_ori_n101_), .C(ori_ori_n219_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n127_), .B(ori_ori_n105_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n92_), .B(ori_ori_n25_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n170_), .B(ori_ori_n223_), .Y(ori_ori_n224_));
  NO2        o202(.A(ori_ori_n224_), .B(ori_ori_n179_), .Y(ori_ori_n225_));
  NA2        o203(.A(ori_ori_n132_), .B(i_10_), .Y(ori_ori_n226_));
  NA3        o204(.A(ori_ori_n160_), .B(ori_ori_n62_), .C(i_2_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  INV        o206(.A(ori_ori_n228_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n229_), .B(ori_ori_n168_), .Y(ori_ori_n230_));
  NO3        o208(.A(ori_ori_n230_), .B(ori_ori_n225_), .C(ori_ori_n208_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n71_), .B(i_13_), .Y(ori_ori_n232_));
  NO2        o210(.A(i_10_), .B(i_9_), .Y(ori_ori_n233_));
  INV        o211(.A(ori_ori_n91_), .Y(ori_ori_n234_));
  NA2        o212(.A(i_8_), .B(i_9_), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n170_), .B(ori_ori_n136_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n235_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n155_), .B(ori_ori_n172_), .Y(ori_ori_n238_));
  NO3        o216(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n239_));
  INV        o217(.A(ori_ori_n239_), .Y(ori_ori_n240_));
  NA3        o218(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n241_));
  NA4        o219(.A(ori_ori_n120_), .B(ori_ori_n100_), .C(ori_ori_n78_), .D(ori_ori_n23_), .Y(ori_ori_n242_));
  OAI220     o220(.A0(ori_ori_n242_), .A1(ori_ori_n241_), .B0(ori_ori_n240_), .B1(ori_ori_n238_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n243_), .B(ori_ori_n237_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n90_), .B(i_13_), .Y(ori_ori_n245_));
  NO3        o223(.A(i_4_), .B(ori_ori_n47_), .C(i_8_), .Y(ori_ori_n246_));
  NO2        o224(.A(i_6_), .B(i_7_), .Y(ori_ori_n247_));
  NO2        o225(.A(i_11_), .B(i_1_), .Y(ori_ori_n248_));
  NOi21      o226(.An(i_2_), .B(i_7_), .Y(ori_ori_n249_));
  NO2        o227(.A(i_6_), .B(i_10_), .Y(ori_ori_n250_));
  NA3        o228(.A(ori_ori_n154_), .B(ori_ori_n126_), .C(ori_ori_n111_), .Y(ori_ori_n251_));
  NA2        o229(.A(ori_ori_n45_), .B(ori_ori_n43_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n239_), .B(ori_ori_n212_), .Y(ori_ori_n253_));
  NAi21      o231(.An(ori_ori_n140_), .B(ori_ori_n213_), .Y(ori_ori_n254_));
  NA2        o232(.A(ori_ori_n178_), .B(ori_ori_n141_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n255_), .B(ori_ori_n254_), .Y(ori_ori_n256_));
  NA2        o234(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n257_));
  NA2        o235(.A(ori_ori_n173_), .B(ori_ori_n149_), .Y(ori_ori_n258_));
  OAI220     o236(.A0(ori_ori_n258_), .A1(ori_ori_n227_), .B0(ori_ori_n257_), .B1(ori_ori_n245_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n259_), .B(ori_ori_n256_), .Y(ori_ori_n260_));
  NA3        o238(.A(ori_ori_n260_), .B(ori_ori_n251_), .C(ori_ori_n244_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n209_), .B(ori_ori_n145_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n197_), .B(ori_ori_n190_), .Y(ori_ori_n263_));
  OR2        o241(.A(ori_ori_n262_), .B(ori_ori_n263_), .Y(ori_ori_n264_));
  AOI210     o242(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n221_), .Y(ori_ori_n265_));
  NA2        o243(.A(ori_ori_n265_), .B(ori_ori_n264_), .Y(ori_ori_n266_));
  INV        o244(.A(ori_ori_n266_), .Y(ori_ori_n267_));
  NA2        o245(.A(ori_ori_n160_), .B(ori_ori_n62_), .Y(ori_ori_n268_));
  OAI210     o246(.A0(i_8_), .A1(ori_ori_n268_), .B0(ori_ori_n113_), .Y(ori_ori_n269_));
  NA2        o247(.A(ori_ori_n269_), .B(ori_ori_n222_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(ori_ori_n267_), .Y(ori_ori_n271_));
  NO2        o249(.A(i_12_), .B(ori_ori_n132_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n43_), .B(i_10_), .Y(ori_ori_n273_));
  NO2        o251(.A(ori_ori_n273_), .B(i_6_), .Y(ori_ori_n274_));
  NO2        o252(.A(i_0_), .B(i_5_), .Y(ori_ori_n275_));
  NA2        o253(.A(ori_ori_n170_), .B(ori_ori_n79_), .Y(ori_ori_n276_));
  NO2        o254(.A(i_11_), .B(ori_ori_n276_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n144_), .B(ori_ori_n143_), .Y(ori_ori_n278_));
  NA2        o256(.A(ori_ori_n233_), .B(i_4_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n278_), .B(ori_ori_n279_), .Y(ori_ori_n280_));
  AOI210     o258(.A0(ori_ori_n191_), .A1(ori_ori_n45_), .B0(ori_ori_n194_), .Y(ori_ori_n281_));
  NA2        o259(.A(i_0_), .B(ori_ori_n47_), .Y(ori_ori_n282_));
  NA3        o260(.A(ori_ori_n272_), .B(ori_ori_n169_), .C(ori_ori_n282_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n281_), .B(ori_ori_n283_), .Y(ori_ori_n284_));
  NO3        o262(.A(ori_ori_n284_), .B(ori_ori_n280_), .C(ori_ori_n277_), .Y(ori_ori_n285_));
  NOi21      o263(.An(i_10_), .B(i_6_), .Y(ori_ori_n286_));
  NO2        o264(.A(ori_ori_n80_), .B(ori_ori_n25_), .Y(ori_ori_n287_));
  INV        o265(.A(ori_ori_n174_), .Y(ori_ori_n288_));
  NO2        o266(.A(i_12_), .B(ori_ori_n80_), .Y(ori_ori_n289_));
  NA3        o267(.A(ori_ori_n289_), .B(ori_ori_n169_), .C(ori_ori_n282_), .Y(ori_ori_n290_));
  NA3        o268(.A(ori_ori_n211_), .B(ori_ori_n170_), .C(ori_ori_n141_), .Y(ori_ori_n291_));
  AOI210     o269(.A0(ori_ori_n291_), .A1(ori_ori_n290_), .B0(ori_ori_n288_), .Y(ori_ori_n292_));
  OR2        o270(.A(i_2_), .B(i_5_), .Y(ori_ori_n293_));
  OR2        o271(.A(ori_ori_n293_), .B(ori_ori_n217_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n199_), .B(ori_ori_n153_), .Y(ori_ori_n295_));
  AOI210     o273(.A0(ori_ori_n295_), .A1(ori_ori_n294_), .B0(ori_ori_n254_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n296_), .B(ori_ori_n292_), .Y(ori_ori_n297_));
  NA2        o275(.A(ori_ori_n297_), .B(ori_ori_n285_), .Y(ori_ori_n298_));
  NO3        o276(.A(ori_ori_n298_), .B(ori_ori_n271_), .C(ori_ori_n261_), .Y(ori_ori_n299_));
  NA4        o277(.A(ori_ori_n299_), .B(ori_ori_n231_), .C(ori_ori_n187_), .D(ori_ori_n166_), .Y(ori7));
  NO2        o278(.A(ori_ori_n87_), .B(ori_ori_n52_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n250_), .B(ori_ori_n79_), .Y(ori_ori_n302_));
  NA2        o280(.A(i_11_), .B(ori_ori_n132_), .Y(ori_ori_n303_));
  NO2        o281(.A(i_13_), .B(ori_ori_n302_), .Y(ori_ori_n304_));
  NA3        o282(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n148_), .B(i_4_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n306_), .B(i_8_), .Y(ori_ori_n307_));
  NO2        o285(.A(ori_ori_n95_), .B(ori_ori_n305_), .Y(ori_ori_n308_));
  NA2        o286(.A(i_2_), .B(ori_ori_n80_), .Y(ori_ori_n309_));
  OAI210     o287(.A0(ori_ori_n81_), .A1(ori_ori_n134_), .B0(ori_ori_n135_), .Y(ori_ori_n310_));
  NO2        o288(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n311_));
  NA2        o289(.A(i_4_), .B(i_8_), .Y(ori_ori_n312_));
  AOI210     o290(.A0(ori_ori_n312_), .A1(ori_ori_n171_), .B0(ori_ori_n311_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n313_), .B(ori_ori_n309_), .Y(ori_ori_n314_));
  NO4        o292(.A(ori_ori_n314_), .B(ori_ori_n308_), .C(ori_ori_n304_), .D(ori_ori_n301_), .Y(ori_ori_n315_));
  OR2        o293(.A(i_6_), .B(i_10_), .Y(ori_ori_n316_));
  NO2        o294(.A(ori_ori_n316_), .B(ori_ori_n23_), .Y(ori_ori_n317_));
  OR3        o295(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n318_));
  INV        o296(.A(ori_ori_n133_), .Y(ori_ori_n319_));
  INV        o297(.A(ori_ori_n317_), .Y(ori_ori_n320_));
  OR2        o298(.A(ori_ori_n320_), .B(ori_ori_n288_), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n321_), .A1(ori_ori_n315_), .B0(ori_ori_n61_), .Y(ori_ori_n322_));
  NOi21      o300(.An(i_11_), .B(i_7_), .Y(ori_ori_n323_));
  AO210      o301(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n324_));
  NO2        o302(.A(ori_ori_n324_), .B(ori_ori_n323_), .Y(ori_ori_n325_));
  NA2        o303(.A(ori_ori_n325_), .B(ori_ori_n137_), .Y(ori_ori_n326_));
  NA3        o304(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n326_), .B(ori_ori_n61_), .Y(ori_ori_n328_));
  NO3        o306(.A(ori_ori_n162_), .B(ori_ori_n138_), .C(ori_ori_n303_), .Y(ori_ori_n329_));
  OAI210     o307(.A0(ori_ori_n329_), .A1(ori_ori_n146_), .B0(ori_ori_n61_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n218_), .B(ori_ori_n31_), .Y(ori_ori_n331_));
  OR2        o309(.A(ori_ori_n138_), .B(ori_ori_n96_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n332_), .B(ori_ori_n331_), .Y(ori_ori_n333_));
  NO2        o311(.A(i_1_), .B(i_4_), .Y(ori_ori_n334_));
  NA2        o312(.A(ori_ori_n334_), .B(ori_ori_n333_), .Y(ori_ori_n335_));
  NO2        o313(.A(i_1_), .B(i_12_), .Y(ori_ori_n336_));
  NA3        o314(.A(ori_ori_n336_), .B(ori_ori_n98_), .C(ori_ori_n24_), .Y(ori_ori_n337_));
  BUFFER     o315(.A(ori_ori_n337_), .Y(ori_ori_n338_));
  NA3        o316(.A(ori_ori_n338_), .B(ori_ori_n335_), .C(ori_ori_n330_), .Y(ori_ori_n339_));
  OAI210     o317(.A0(ori_ori_n339_), .A1(ori_ori_n328_), .B0(i_6_), .Y(ori_ori_n340_));
  NO2        o318(.A(ori_ori_n327_), .B(ori_ori_n96_), .Y(ori_ori_n341_));
  NA2        o319(.A(ori_ori_n341_), .B(ori_ori_n289_), .Y(ori_ori_n342_));
  NO2        o320(.A(i_6_), .B(i_11_), .Y(ori_ori_n343_));
  INV        o321(.A(ori_ori_n342_), .Y(ori_ori_n344_));
  NO3        o322(.A(ori_ori_n316_), .B(i_8_), .C(ori_ori_n23_), .Y(ori_ori_n345_));
  AOI210     o323(.A0(i_1_), .A1(ori_ori_n163_), .B0(ori_ori_n345_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n346_), .B(ori_ori_n43_), .Y(ori_ori_n347_));
  NA3        o325(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n348_));
  NA2        o326(.A(i_2_), .B(ori_ori_n43_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n349_), .B(ori_ori_n348_), .Y(ori_ori_n350_));
  AOI210     o328(.A0(ori_ori_n248_), .A1(ori_ori_n223_), .B0(ori_ori_n151_), .Y(ori_ori_n351_));
  NO2        o329(.A(ori_ori_n351_), .B(ori_ori_n309_), .Y(ori_ori_n352_));
  OR2        o330(.A(ori_ori_n352_), .B(ori_ori_n350_), .Y(ori_ori_n353_));
  NO3        o331(.A(ori_ori_n353_), .B(ori_ori_n347_), .C(ori_ori_n344_), .Y(ori_ori_n354_));
  NO2        o332(.A(ori_ori_n148_), .B(ori_ori_n92_), .Y(ori_ori_n355_));
  NO2        o333(.A(ori_ori_n355_), .B(ori_ori_n323_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(i_1_), .Y(ori_ori_n357_));
  NO2        o335(.A(ori_ori_n357_), .B(ori_ori_n318_), .Y(ori_ori_n358_));
  NO2        o336(.A(ori_ori_n219_), .B(ori_ori_n80_), .Y(ori_ori_n359_));
  NA2        o337(.A(ori_ori_n358_), .B(ori_ori_n45_), .Y(ori_ori_n360_));
  NA2        o338(.A(i_3_), .B(ori_ori_n132_), .Y(ori_ori_n361_));
  NO2        o339(.A(ori_ori_n361_), .B(ori_ori_n99_), .Y(ori_ori_n362_));
  AN2        o340(.A(ori_ori_n362_), .B(ori_ori_n274_), .Y(ori_ori_n363_));
  NO2        o341(.A(i_8_), .B(ori_ori_n43_), .Y(ori_ori_n364_));
  NA2        o342(.A(i_1_), .B(i_3_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n235_), .B(ori_ori_n87_), .Y(ori_ori_n366_));
  AOI210     o344(.A0(ori_ori_n364_), .A1(ori_ori_n286_), .B0(ori_ori_n366_), .Y(ori_ori_n367_));
  NO2        o345(.A(ori_ori_n367_), .B(ori_ori_n365_), .Y(ori_ori_n368_));
  NO2        o346(.A(ori_ori_n368_), .B(ori_ori_n363_), .Y(ori_ori_n369_));
  NA4        o347(.A(ori_ori_n369_), .B(ori_ori_n360_), .C(ori_ori_n354_), .D(ori_ori_n340_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n197_), .B(ori_ori_n196_), .Y(ori_ori_n371_));
  NO3        o349(.A(ori_ori_n249_), .B(ori_ori_n312_), .C(ori_ori_n80_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n372_), .B(ori_ori_n25_), .Y(ori_ori_n373_));
  NA2        o351(.A(ori_ori_n373_), .B(ori_ori_n371_), .Y(ori_ori_n374_));
  NA2        o352(.A(ori_ori_n374_), .B(i_1_), .Y(ori_ori_n375_));
  INV        o353(.A(i_1_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n375_), .B(i_13_), .Y(ori_ori_n377_));
  OR2        o355(.A(i_11_), .B(i_7_), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n52_), .B(i_12_), .Y(ori_ori_n379_));
  INV        o357(.A(ori_ori_n379_), .Y(ori_ori_n380_));
  NO2        o358(.A(ori_ori_n249_), .B(ori_ori_n24_), .Y(ori_ori_n381_));
  AOI220     o359(.A0(ori_ori_n381_), .A1(ori_ori_n359_), .B0(ori_ori_n154_), .B1(ori_ori_n110_), .Y(ori_ori_n382_));
  OAI220     o360(.A0(ori_ori_n382_), .A1(ori_ori_n41_), .B0(ori_ori_n380_), .B1(ori_ori_n87_), .Y(ori_ori_n383_));
  INV        o361(.A(ori_ori_n383_), .Y(ori_ori_n384_));
  NOi31      o362(.An(ori_ori_n577_), .B(ori_ori_n302_), .C(ori_ori_n43_), .Y(ori_ori_n385_));
  NA2        o363(.A(ori_ori_n109_), .B(i_13_), .Y(ori_ori_n386_));
  NO2        o364(.A(ori_ori_n348_), .B(ori_ori_n99_), .Y(ori_ori_n387_));
  INV        o365(.A(ori_ori_n387_), .Y(ori_ori_n388_));
  OAI220     o366(.A0(ori_ori_n388_), .A1(ori_ori_n69_), .B0(ori_ori_n386_), .B1(ori_ori_n376_), .Y(ori_ori_n389_));
  NO3        o367(.A(ori_ori_n69_), .B(ori_ori_n32_), .C(ori_ori_n92_), .Y(ori_ori_n390_));
  INV        o368(.A(ori_ori_n390_), .Y(ori_ori_n391_));
  AOI210     o369(.A0(ori_ori_n211_), .A1(i_2_), .B0(ori_ori_n86_), .Y(ori_ori_n392_));
  OAI220     o370(.A0(ori_ori_n392_), .A1(ori_ori_n307_), .B0(ori_ori_n391_), .B1(ori_ori_n319_), .Y(ori_ori_n393_));
  NO3        o371(.A(ori_ori_n393_), .B(ori_ori_n389_), .C(ori_ori_n385_), .Y(ori_ori_n394_));
  OR2        o372(.A(i_11_), .B(i_6_), .Y(ori_ori_n395_));
  NA3        o373(.A(ori_ori_n218_), .B(ori_ori_n311_), .C(ori_ori_n91_), .Y(ori_ori_n396_));
  NA2        o374(.A(ori_ori_n343_), .B(i_13_), .Y(ori_ori_n397_));
  NAi21      o375(.An(i_11_), .B(i_12_), .Y(ori_ori_n398_));
  NO3        o376(.A(ori_ori_n398_), .B(i_13_), .C(ori_ori_n80_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n289_), .B(ori_ori_n312_), .Y(ori_ori_n400_));
  AOI210     o378(.A0(ori_ori_n400_), .A1(ori_ori_n173_), .B0(ori_ori_n399_), .Y(ori_ori_n401_));
  NA3        o379(.A(ori_ori_n401_), .B(ori_ori_n397_), .C(ori_ori_n396_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n402_), .B(ori_ori_n61_), .Y(ori_ori_n403_));
  NO2        o381(.A(i_2_), .B(i_12_), .Y(ori_ori_n404_));
  NA3        o382(.A(ori_ori_n403_), .B(ori_ori_n394_), .C(ori_ori_n384_), .Y(ori_ori_n405_));
  OR4        o383(.A(ori_ori_n405_), .B(ori_ori_n377_), .C(ori_ori_n370_), .D(ori_ori_n322_), .Y(ori5));
  NA2        o384(.A(ori_ori_n356_), .B(ori_ori_n167_), .Y(ori_ori_n407_));
  NA3        o385(.A(ori_ori_n24_), .B(ori_ori_n404_), .C(ori_ori_n96_), .Y(ori_ori_n408_));
  NO2        o386(.A(ori_ori_n307_), .B(i_11_), .Y(ori_ori_n409_));
  NA2        o387(.A(ori_ori_n81_), .B(ori_ori_n409_), .Y(ori_ori_n410_));
  NA3        o388(.A(ori_ori_n410_), .B(ori_ori_n408_), .C(ori_ori_n407_), .Y(ori_ori_n411_));
  NO3        o389(.A(i_11_), .B(ori_ori_n148_), .C(i_13_), .Y(ori_ori_n412_));
  NO2        o390(.A(ori_ori_n106_), .B(ori_ori_n23_), .Y(ori_ori_n413_));
  NA2        o391(.A(i_12_), .B(i_8_), .Y(ori_ori_n414_));
  OAI210     o392(.A0(ori_ori_n45_), .A1(i_3_), .B0(ori_ori_n414_), .Y(ori_ori_n415_));
  INV        o393(.A(ori_ori_n233_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n415_), .B(ori_ori_n413_), .Y(ori_ori_n417_));
  INV        o395(.A(ori_ori_n417_), .Y(ori_ori_n418_));
  NO2        o396(.A(ori_ori_n418_), .B(ori_ori_n411_), .Y(ori_ori_n419_));
  INV        o397(.A(ori_ori_n126_), .Y(ori_ori_n420_));
  INV        o398(.A(ori_ori_n154_), .Y(ori_ori_n421_));
  NO2        o399(.A(ori_ori_n421_), .B(ori_ori_n420_), .Y(ori_ori_n422_));
  NO2        o400(.A(ori_ori_n235_), .B(ori_ori_n26_), .Y(ori_ori_n423_));
  NO2        o401(.A(ori_ori_n423_), .B(ori_ori_n223_), .Y(ori_ori_n424_));
  NA2        o402(.A(ori_ori_n424_), .B(i_2_), .Y(ori_ori_n425_));
  INV        o403(.A(ori_ori_n425_), .Y(ori_ori_n426_));
  AOI210     o404(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n220_), .Y(ori_ori_n427_));
  AOI210     o405(.A0(ori_ori_n427_), .A1(ori_ori_n426_), .B0(ori_ori_n422_), .Y(ori_ori_n428_));
  NO2        o406(.A(ori_ori_n131_), .B(ori_ori_n107_), .Y(ori_ori_n429_));
  OAI210     o407(.A0(ori_ori_n429_), .A1(ori_ori_n413_), .B0(i_2_), .Y(ori_ori_n430_));
  INV        o408(.A(ori_ori_n127_), .Y(ori_ori_n431_));
  NO3        o409(.A(ori_ori_n324_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n432_));
  AOI210     o410(.A0(ori_ori_n431_), .A1(ori_ori_n81_), .B0(ori_ori_n432_), .Y(ori_ori_n433_));
  AOI210     o411(.A0(ori_ori_n433_), .A1(ori_ori_n430_), .B0(ori_ori_n132_), .Y(ori_ori_n434_));
  OA210      o412(.A0(ori_ori_n325_), .A1(ori_ori_n108_), .B0(i_13_), .Y(ori_ori_n435_));
  NA2        o413(.A(ori_ori_n133_), .B(ori_ori_n134_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n436_), .B(ori_ori_n199_), .Y(ori_ori_n437_));
  INV        o415(.A(ori_ori_n138_), .Y(ori_ori_n438_));
  NA2        o416(.A(ori_ori_n438_), .B(ori_ori_n223_), .Y(ori_ori_n439_));
  NA3        o417(.A(i_2_), .B(ori_ori_n171_), .C(ori_ori_n106_), .Y(ori_ori_n440_));
  NA2        o418(.A(ori_ori_n440_), .B(ori_ori_n439_), .Y(ori_ori_n441_));
  NO4        o419(.A(ori_ori_n441_), .B(ori_ori_n437_), .C(ori_ori_n435_), .D(ori_ori_n434_), .Y(ori_ori_n442_));
  NO2        o420(.A(ori_ori_n60_), .B(i_12_), .Y(ori_ori_n443_));
  NO2        o421(.A(ori_ori_n443_), .B(ori_ori_n108_), .Y(ori_ori_n444_));
  NO2        o422(.A(ori_ori_n444_), .B(ori_ori_n303_), .Y(ori_ori_n445_));
  NA2        o423(.A(ori_ori_n445_), .B(ori_ori_n36_), .Y(ori_ori_n446_));
  NA4        o424(.A(ori_ori_n446_), .B(ori_ori_n442_), .C(ori_ori_n428_), .D(ori_ori_n419_), .Y(ori6));
  NO2        o425(.A(ori_ori_n142_), .B(ori_ori_n252_), .Y(ori_ori_n448_));
  INV        o426(.A(ori_ori_n177_), .Y(ori_ori_n449_));
  OR2        o427(.A(ori_ori_n449_), .B(i_12_), .Y(ori_ori_n450_));
  INV        o428(.A(ori_ori_n176_), .Y(ori_ori_n451_));
  NA2        o429(.A(ori_ori_n73_), .B(ori_ori_n110_), .Y(ori_ori_n452_));
  NO2        o430(.A(ori_ori_n452_), .B(ori_ori_n451_), .Y(ori_ori_n453_));
  NO2        o431(.A(ori_ori_n156_), .B(i_9_), .Y(ori_ori_n454_));
  NA2        o432(.A(ori_ori_n454_), .B(ori_ori_n443_), .Y(ori_ori_n455_));
  AOI210     o433(.A0(ori_ori_n455_), .A1(ori_ori_n263_), .B0(ori_ori_n129_), .Y(ori_ori_n456_));
  NO2        o434(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n457_));
  NAi32      o435(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n458_));
  NO2        o436(.A(ori_ori_n395_), .B(ori_ori_n458_), .Y(ori_ori_n459_));
  OR3        o437(.A(ori_ori_n459_), .B(ori_ori_n456_), .C(ori_ori_n453_), .Y(ori_ori_n460_));
  NO2        o438(.A(ori_ori_n378_), .B(i_2_), .Y(ori_ori_n461_));
  NA2        o439(.A(ori_ori_n47_), .B(ori_ori_n37_), .Y(ori_ori_n462_));
  INV        o440(.A(ori_ori_n462_), .Y(ori_ori_n463_));
  NA2        o441(.A(ori_ori_n463_), .B(ori_ori_n461_), .Y(ori_ori_n464_));
  BUFFER     o442(.A(ori_ori_n325_), .Y(ori_ori_n465_));
  NA2        o443(.A(ori_ori_n465_), .B(ori_ori_n121_), .Y(ori_ori_n466_));
  AO210      o444(.A0(ori_ori_n253_), .A1(ori_ori_n416_), .B0(ori_ori_n36_), .Y(ori_ori_n467_));
  NA3        o445(.A(ori_ori_n467_), .B(ori_ori_n466_), .C(ori_ori_n464_), .Y(ori_ori_n468_));
  INV        o446(.A(ori_ori_n448_), .Y(ori_ori_n469_));
  NA3        o447(.A(ori_ori_n199_), .B(ori_ori_n149_), .C(ori_ori_n121_), .Y(ori_ori_n470_));
  NA3        o448(.A(ori_ori_n470_), .B(ori_ori_n469_), .C(ori_ori_n310_), .Y(ori_ori_n471_));
  NO2        o449(.A(ori_ori_n316_), .B(i_2_), .Y(ori_ori_n472_));
  OAI210     o450(.A0(ori_ori_n472_), .A1(ori_ori_n78_), .B0(ori_ori_n216_), .Y(ori_ori_n473_));
  INV        o451(.A(ori_ori_n294_), .Y(ori_ori_n474_));
  NA2        o452(.A(ori_ori_n474_), .B(ori_ori_n176_), .Y(ori_ori_n475_));
  NA2        o453(.A(ori_ori_n475_), .B(ori_ori_n473_), .Y(ori_ori_n476_));
  NO4        o454(.A(ori_ori_n476_), .B(ori_ori_n471_), .C(ori_ori_n468_), .D(ori_ori_n460_), .Y(ori_ori_n477_));
  NA3        o455(.A(ori_ori_n477_), .B(ori_ori_n450_), .C(ori_ori_n207_), .Y(ori3));
  NA2        o456(.A(i_12_), .B(i_10_), .Y(ori_ori_n479_));
  NO2        o457(.A(i_11_), .B(ori_ori_n148_), .Y(ori_ori_n480_));
  NA3        o458(.A(ori_ori_n470_), .B(ori_ori_n310_), .C(ori_ori_n198_), .Y(ori_ori_n481_));
  NA2        o459(.A(ori_ori_n481_), .B(ori_ori_n40_), .Y(ori_ori_n482_));
  NOi21      o460(.An(ori_ori_n90_), .B(ori_ori_n424_), .Y(ori_ori_n483_));
  NO3        o461(.A(ori_ori_n332_), .B(ori_ori_n235_), .C(ori_ori_n110_), .Y(ori_ori_n484_));
  NA2        o462(.A(ori_ori_n218_), .B(ori_ori_n44_), .Y(ori_ori_n485_));
  AN2        o463(.A(ori_ori_n234_), .B(ori_ori_n53_), .Y(ori_ori_n486_));
  NO3        o464(.A(ori_ori_n486_), .B(ori_ori_n484_), .C(ori_ori_n483_), .Y(ori_ori_n487_));
  AOI210     o465(.A0(ori_ori_n487_), .A1(ori_ori_n482_), .B0(ori_ori_n47_), .Y(ori_ori_n488_));
  NO4        o466(.A(ori_ori_n203_), .B(ori_ori_n209_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n489_));
  NA2        o467(.A(ori_ori_n129_), .B(ori_ori_n286_), .Y(ori_ori_n490_));
  NOi21      o468(.An(ori_ori_n490_), .B(ori_ori_n489_), .Y(ori_ori_n491_));
  NO2        o469(.A(ori_ori_n491_), .B(ori_ori_n61_), .Y(ori_ori_n492_));
  NOi21      o470(.An(i_5_), .B(i_9_), .Y(ori_ori_n493_));
  NA2        o471(.A(ori_ori_n493_), .B(ori_ori_n232_), .Y(ori_ori_n494_));
  AOI210     o472(.A0(ori_ori_n578_), .A1(ori_ori_n248_), .B0(ori_ori_n372_), .Y(ori_ori_n495_));
  NO2        o473(.A(ori_ori_n495_), .B(ori_ori_n494_), .Y(ori_ori_n496_));
  NO3        o474(.A(ori_ori_n496_), .B(ori_ori_n492_), .C(ori_ori_n488_), .Y(ori_ori_n497_));
  BUFFER     o475(.A(i_0_), .Y(ori_ori_n498_));
  NA2        o476(.A(ori_ori_n287_), .B(i_0_), .Y(ori_ori_n499_));
  NO3        o477(.A(ori_ori_n499_), .B(ori_ori_n210_), .C(ori_ori_n81_), .Y(ori_ori_n500_));
  NO4        o478(.A(ori_ori_n293_), .B(i_12_), .C(ori_ori_n220_), .D(ori_ori_n217_), .Y(ori_ori_n501_));
  AOI210     o479(.A0(ori_ori_n501_), .A1(i_11_), .B0(ori_ori_n500_), .Y(ori_ori_n502_));
  NA2        o480(.A(ori_ori_n412_), .B(ori_ori_n177_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n81_), .B(ori_ori_n56_), .Y(ori_ori_n504_));
  NO2        o482(.A(ori_ori_n504_), .B(ori_ori_n503_), .Y(ori_ori_n505_));
  NO2        o483(.A(ori_ori_n158_), .B(ori_ori_n122_), .Y(ori_ori_n506_));
  NO4        o484(.A(ori_ori_n99_), .B(ori_ori_n56_), .C(ori_ori_n361_), .D(i_5_), .Y(ori_ori_n507_));
  AO220      o485(.A0(ori_ori_n507_), .A1(i_10_), .B0(ori_ori_n506_), .B1(i_6_), .Y(ori_ori_n508_));
  NO2        o486(.A(ori_ori_n508_), .B(ori_ori_n505_), .Y(ori_ori_n509_));
  NA2        o487(.A(ori_ori_n509_), .B(ori_ori_n502_), .Y(ori_ori_n510_));
  NO2        o488(.A(ori_ori_n93_), .B(ori_ori_n37_), .Y(ori_ori_n511_));
  NA2        o489(.A(i_11_), .B(i_9_), .Y(ori_ori_n512_));
  NO3        o490(.A(i_12_), .B(ori_ori_n512_), .C(ori_ori_n309_), .Y(ori_ori_n513_));
  AN2        o491(.A(ori_ori_n513_), .B(ori_ori_n511_), .Y(ori_ori_n514_));
  NO2        o492(.A(ori_ori_n512_), .B(ori_ori_n71_), .Y(ori_ori_n515_));
  INV        o493(.A(ori_ori_n215_), .Y(ori_ori_n516_));
  NO2        o494(.A(ori_ori_n516_), .B(ori_ori_n494_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n517_), .B(ori_ori_n514_), .Y(ori_ori_n518_));
  INV        o496(.A(ori_ori_n175_), .Y(ori_ori_n519_));
  INV        o497(.A(ori_ori_n518_), .Y(ori_ori_n520_));
  INV        o498(.A(ori_ori_n479_), .Y(ori_ori_n521_));
  OA210      o499(.A0(ori_ori_n247_), .A1(ori_ori_n144_), .B0(ori_ori_n246_), .Y(ori_ori_n522_));
  NA2        o500(.A(ori_ori_n521_), .B(ori_ori_n515_), .Y(ori_ori_n523_));
  NA2        o501(.A(ori_ori_n381_), .B(ori_ori_n275_), .Y(ori_ori_n524_));
  NAi21      o502(.An(i_9_), .B(i_5_), .Y(ori_ori_n525_));
  NO2        o503(.A(ori_ori_n525_), .B(ori_ori_n214_), .Y(ori_ori_n526_));
  NA2        o504(.A(ori_ori_n526_), .B(ori_ori_n325_), .Y(ori_ori_n527_));
  OAI220     o505(.A0(ori_ori_n527_), .A1(ori_ori_n80_), .B0(ori_ori_n524_), .B1(ori_ori_n127_), .Y(ori_ori_n528_));
  NO2        o506(.A(ori_ori_n528_), .B(ori_ori_n266_), .Y(ori_ori_n529_));
  NA2        o507(.A(ori_ori_n529_), .B(ori_ori_n523_), .Y(ori_ori_n530_));
  NO3        o508(.A(ori_ori_n530_), .B(ori_ori_n520_), .C(ori_ori_n510_), .Y(ori_ori_n531_));
  NO2        o509(.A(ori_ori_n498_), .B(ori_ori_n398_), .Y(ori_ori_n532_));
  NA2        o510(.A(ori_ori_n153_), .B(ori_ori_n147_), .Y(ori_ori_n533_));
  AOI210     o511(.A0(ori_ori_n533_), .A1(ori_ori_n499_), .B0(ori_ori_n122_), .Y(ori_ori_n534_));
  NO3        o512(.A(ori_ori_n139_), .B(ori_ori_n209_), .C(i_0_), .Y(ori_ori_n535_));
  OAI210     o513(.A0(ori_ori_n535_), .A1(ori_ori_n74_), .B0(i_13_), .Y(ori_ori_n536_));
  INV        o514(.A(ori_ori_n536_), .Y(ori_ori_n537_));
  NO2        o515(.A(ori_ori_n152_), .B(ori_ori_n87_), .Y(ori_ori_n538_));
  AOI210     o516(.A0(ori_ori_n538_), .A1(ori_ori_n532_), .B0(ori_ori_n97_), .Y(ori_ori_n539_));
  OR2        o517(.A(ori_ori_n539_), .B(i_5_), .Y(ori_ori_n540_));
  AOI210     o518(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n128_), .Y(ori_ori_n541_));
  NA2        o519(.A(ori_ori_n541_), .B(ori_ori_n522_), .Y(ori_ori_n542_));
  NO3        o520(.A(ori_ori_n485_), .B(ori_ori_n52_), .C(ori_ori_n47_), .Y(ori_ori_n543_));
  INV        o521(.A(ori_ori_n251_), .Y(ori_ori_n544_));
  NO2        o522(.A(ori_ori_n544_), .B(ori_ori_n543_), .Y(ori_ori_n545_));
  NA3        o523(.A(ori_ori_n212_), .B(ori_ori_n126_), .C(ori_ori_n125_), .Y(ori_ori_n546_));
  INV        o524(.A(ori_ori_n546_), .Y(ori_ori_n547_));
  NO3        o525(.A(ori_ori_n512_), .B(ori_ori_n141_), .C(ori_ori_n131_), .Y(ori_ori_n548_));
  NO2        o526(.A(ori_ori_n548_), .B(ori_ori_n547_), .Y(ori_ori_n549_));
  NA4        o527(.A(ori_ori_n549_), .B(ori_ori_n545_), .C(ori_ori_n542_), .D(ori_ori_n540_), .Y(ori_ori_n550_));
  NO2        o528(.A(ori_ori_n80_), .B(i_5_), .Y(ori_ori_n551_));
  NA3        o529(.A(ori_ori_n480_), .B(ori_ori_n98_), .C(ori_ori_n106_), .Y(ori_ori_n552_));
  INV        o530(.A(ori_ori_n552_), .Y(ori_ori_n553_));
  NA2        o531(.A(ori_ori_n553_), .B(ori_ori_n551_), .Y(ori_ori_n554_));
  NAi21      o532(.An(ori_ori_n151_), .B(ori_ori_n152_), .Y(ori_ori_n555_));
  NO4        o533(.A(ori_ori_n150_), .B(ori_ori_n139_), .C(i_0_), .D(i_12_), .Y(ori_ori_n556_));
  NA2        o534(.A(ori_ori_n556_), .B(ori_ori_n555_), .Y(ori_ori_n557_));
  NA2        o535(.A(ori_ori_n557_), .B(ori_ori_n554_), .Y(ori_ori_n558_));
  NO4        o536(.A(ori_ori_n558_), .B(ori_ori_n550_), .C(ori_ori_n537_), .D(ori_ori_n534_), .Y(ori_ori_n559_));
  OAI210     o537(.A0(ori_ori_n461_), .A1(ori_ori_n457_), .B0(ori_ori_n37_), .Y(ori_ori_n560_));
  INV        o538(.A(ori_ori_n560_), .Y(ori_ori_n561_));
  NA2        o539(.A(ori_ori_n561_), .B(ori_ori_n137_), .Y(ori_ori_n562_));
  NAi31      o540(.An(i_7_), .B(i_2_), .C(i_10_), .Y(ori_ori_n563_));
  NO2        o541(.A(ori_ori_n68_), .B(ori_ori_n563_), .Y(ori_ori_n564_));
  AOI210     o542(.A0(ori_ori_n564_), .A1(ori_ori_n47_), .B0(ori_ori_n501_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n565_), .A1(ori_ori_n562_), .B0(ori_ori_n71_), .Y(ori_ori_n566_));
  INV        o544(.A(ori_ori_n206_), .Y(ori_ori_n567_));
  NO2        o545(.A(ori_ori_n567_), .B(ori_ori_n420_), .Y(ori_ori_n568_));
  NO3        o546(.A(ori_ori_n57_), .B(ori_ori_n56_), .C(i_4_), .Y(ori_ori_n569_));
  OAI210     o547(.A0(ori_ori_n519_), .A1(ori_ori_n172_), .B0(ori_ori_n569_), .Y(ori_ori_n570_));
  NO2        o548(.A(ori_ori_n570_), .B(ori_ori_n398_), .Y(ori_ori_n571_));
  NO3        o549(.A(ori_ori_n571_), .B(ori_ori_n568_), .C(ori_ori_n566_), .Y(ori_ori_n572_));
  NA4        o550(.A(ori_ori_n572_), .B(ori_ori_n559_), .C(ori_ori_n531_), .D(ori_ori_n497_), .Y(ori4));
  INV        o551(.A(i_6_), .Y(ori_ori_n576_));
  INV        o552(.A(i_13_), .Y(ori_ori_n577_));
  INV        o553(.A(i_6_), .Y(ori_ori_n578_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  OAI210     m028(.A0(mai_mai_n50_), .A1(i_3_), .B0(mai_mai_n48_), .Y(mai_mai_n51_));
  AOI210     m029(.A0(mai_mai_n51_), .A1(mai_mai_n47_), .B0(mai_mai_n46_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_0_), .B(i_2_), .Y(mai_mai_n53_));
  NA2        m031(.A(i_7_), .B(i_9_), .Y(mai_mai_n54_));
  NA2        m032(.A(mai_mai_n52_), .B(mai_mai_n45_), .Y(mai_mai_n55_));
  NO2        m033(.A(i_1_), .B(i_6_), .Y(mai_mai_n56_));
  NA2        m034(.A(i_8_), .B(i_7_), .Y(mai_mai_n57_));
  NAi21      m035(.An(i_2_), .B(i_7_), .Y(mai_mai_n58_));
  INV        m036(.A(i_1_), .Y(mai_mai_n59_));
  NA2        m037(.A(mai_mai_n59_), .B(i_6_), .Y(mai_mai_n60_));
  NA2        m038(.A(i_1_), .B(i_10_), .Y(mai_mai_n61_));
  NO2        m039(.A(mai_mai_n61_), .B(i_6_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n63_));
  AOI210     m041(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n64_));
  NA2        m042(.A(i_1_), .B(i_6_), .Y(mai_mai_n65_));
  NO2        m043(.A(mai_mai_n65_), .B(mai_mai_n25_), .Y(mai_mai_n66_));
  INV        m044(.A(i_0_), .Y(mai_mai_n67_));
  NAi21      m045(.An(i_5_), .B(i_10_), .Y(mai_mai_n68_));
  NA2        m046(.A(i_5_), .B(i_9_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n68_), .B0(mai_mai_n67_), .Y(mai_mai_n70_));
  NO2        m048(.A(mai_mai_n70_), .B(mai_mai_n66_), .Y(mai_mai_n71_));
  OAI210     m049(.A0(mai_mai_n64_), .A1(mai_mai_n63_), .B0(mai_mai_n71_), .Y(mai_mai_n72_));
  OAI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n62_), .B0(i_0_), .Y(mai_mai_n73_));
  NA2        m051(.A(i_12_), .B(i_5_), .Y(mai_mai_n74_));
  NA2        m052(.A(i_2_), .B(i_8_), .Y(mai_mai_n75_));
  NO2        m053(.A(i_3_), .B(i_9_), .Y(mai_mai_n76_));
  NO2        m054(.A(i_3_), .B(i_7_), .Y(mai_mai_n77_));
  NO3        m055(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(mai_mai_n59_), .Y(mai_mai_n78_));
  INV        m056(.A(i_6_), .Y(mai_mai_n79_));
  OR4        m057(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n80_));
  INV        m058(.A(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m059(.A(i_2_), .B(i_7_), .Y(mai_mai_n82_));
  NA2        m060(.A(mai_mai_n78_), .B(mai_mai_n80_), .Y(mai_mai_n83_));
  NAi21      m061(.An(i_6_), .B(i_10_), .Y(mai_mai_n84_));
  NA2        m062(.A(i_6_), .B(i_9_), .Y(mai_mai_n85_));
  AOI210     m063(.A0(mai_mai_n85_), .A1(mai_mai_n84_), .B0(mai_mai_n59_), .Y(mai_mai_n86_));
  NA2        m064(.A(i_2_), .B(i_6_), .Y(mai_mai_n87_));
  NO2        m065(.A(mai_mai_n83_), .B(mai_mai_n74_), .Y(mai_mai_n88_));
  AN3        m066(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n89_));
  NAi21      m067(.An(i_6_), .B(i_11_), .Y(mai_mai_n90_));
  NO2        m068(.A(i_5_), .B(i_8_), .Y(mai_mai_n91_));
  NOi21      m069(.An(mai_mai_n91_), .B(mai_mai_n90_), .Y(mai_mai_n92_));
  AOI220     m070(.A0(mai_mai_n92_), .A1(mai_mai_n58_), .B0(mai_mai_n89_), .B1(mai_mai_n32_), .Y(mai_mai_n93_));
  INV        m071(.A(i_7_), .Y(mai_mai_n94_));
  NA2        m072(.A(mai_mai_n46_), .B(mai_mai_n94_), .Y(mai_mai_n95_));
  NO2        m073(.A(i_0_), .B(i_5_), .Y(mai_mai_n96_));
  NO2        m074(.A(mai_mai_n96_), .B(mai_mai_n79_), .Y(mai_mai_n97_));
  NA2        m075(.A(i_12_), .B(i_3_), .Y(mai_mai_n98_));
  INV        m076(.A(mai_mai_n98_), .Y(mai_mai_n99_));
  NA2        m077(.A(mai_mai_n99_), .B(mai_mai_n97_), .Y(mai_mai_n100_));
  NAi21      m078(.An(i_7_), .B(i_11_), .Y(mai_mai_n101_));
  AN2        m079(.A(i_2_), .B(i_10_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(i_7_), .Y(mai_mai_n103_));
  OR2        m081(.A(mai_mai_n74_), .B(mai_mai_n56_), .Y(mai_mai_n104_));
  NO2        m082(.A(i_8_), .B(mai_mai_n94_), .Y(mai_mai_n105_));
  NO3        m083(.A(mai_mai_n105_), .B(mai_mai_n104_), .C(mai_mai_n103_), .Y(mai_mai_n106_));
  NA2        m084(.A(i_12_), .B(i_7_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n59_), .B(mai_mai_n26_), .Y(mai_mai_n108_));
  NA2        m086(.A(mai_mai_n108_), .B(i_0_), .Y(mai_mai_n109_));
  NA2        m087(.A(i_11_), .B(i_12_), .Y(mai_mai_n110_));
  OAI210     m088(.A0(mai_mai_n109_), .A1(mai_mai_n107_), .B0(mai_mai_n110_), .Y(mai_mai_n111_));
  NO2        m089(.A(mai_mai_n111_), .B(mai_mai_n106_), .Y(mai_mai_n112_));
  NA3        m090(.A(mai_mai_n112_), .B(mai_mai_n100_), .C(mai_mai_n93_), .Y(mai_mai_n113_));
  NOi21      m091(.An(i_1_), .B(i_5_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n114_), .B(i_11_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n94_), .B(mai_mai_n37_), .Y(mai_mai_n116_));
  NA2        m094(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(mai_mai_n116_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n118_), .B(mai_mai_n46_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n85_), .B(mai_mai_n84_), .Y(mai_mai_n120_));
  NAi21      m098(.An(i_3_), .B(i_8_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n121_), .B(mai_mai_n58_), .Y(mai_mai_n122_));
  NO2        m100(.A(i_6_), .B(i_5_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(i_3_), .Y(mai_mai_n124_));
  NO2        m102(.A(mai_mai_n122_), .B(mai_mai_n115_), .Y(mai_mai_n125_));
  NO3        m103(.A(mai_mai_n125_), .B(mai_mai_n113_), .C(mai_mai_n88_), .Y(mai_mai_n126_));
  NA3        m104(.A(mai_mai_n126_), .B(mai_mai_n73_), .C(mai_mai_n55_), .Y(mai2));
  NO2        m105(.A(mai_mai_n59_), .B(mai_mai_n37_), .Y(mai_mai_n128_));
  NA2        m106(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n129_), .B(mai_mai_n128_), .Y(mai_mai_n130_));
  NA4        m108(.A(mai_mai_n130_), .B(mai_mai_n71_), .C(mai_mai_n63_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m109(.A(i_8_), .B(i_7_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n132_), .B(i_6_), .Y(mai_mai_n133_));
  NO2        m111(.A(i_12_), .B(i_13_), .Y(mai_mai_n134_));
  NAi21      m112(.An(i_5_), .B(i_11_), .Y(mai_mai_n135_));
  NOi21      m113(.An(mai_mai_n134_), .B(mai_mai_n135_), .Y(mai_mai_n136_));
  NO2        m114(.A(i_0_), .B(i_1_), .Y(mai_mai_n137_));
  NA2        m115(.A(i_2_), .B(i_3_), .Y(mai_mai_n138_));
  NO2        m116(.A(mai_mai_n138_), .B(i_4_), .Y(mai_mai_n139_));
  NA3        m117(.A(mai_mai_n139_), .B(mai_mai_n137_), .C(mai_mai_n136_), .Y(mai_mai_n140_));
  AN2        m118(.A(mai_mai_n134_), .B(mai_mai_n76_), .Y(mai_mai_n141_));
  NA2        m119(.A(i_1_), .B(i_5_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n67_), .B(mai_mai_n46_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(mai_mai_n36_), .Y(mai_mai_n144_));
  NO3        m122(.A(mai_mai_n144_), .B(mai_mai_n142_), .C(i_13_), .Y(mai_mai_n145_));
  OR2        m123(.A(i_0_), .B(i_1_), .Y(mai_mai_n146_));
  NO3        m124(.A(mai_mai_n146_), .B(mai_mai_n74_), .C(i_13_), .Y(mai_mai_n147_));
  NAi32      m125(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n148_));
  NAi21      m126(.An(mai_mai_n148_), .B(mai_mai_n147_), .Y(mai_mai_n149_));
  NOi21      m127(.An(i_4_), .B(i_10_), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n150_), .B(mai_mai_n40_), .Y(mai_mai_n151_));
  NO2        m129(.A(i_3_), .B(i_5_), .Y(mai_mai_n152_));
  NO3        m130(.A(mai_mai_n67_), .B(i_2_), .C(i_1_), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  OAI210     m132(.A0(mai_mai_n154_), .A1(mai_mai_n151_), .B0(mai_mai_n149_), .Y(mai_mai_n155_));
  NO2        m133(.A(mai_mai_n155_), .B(mai_mai_n145_), .Y(mai_mai_n156_));
  AOI210     m134(.A0(mai_mai_n156_), .A1(mai_mai_n140_), .B0(mai_mai_n133_), .Y(mai_mai_n157_));
  NA2        m135(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n158_));
  NOi21      m136(.An(i_4_), .B(i_9_), .Y(mai_mai_n159_));
  NOi21      m137(.An(i_11_), .B(i_13_), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n160_), .B(mai_mai_n159_), .Y(mai_mai_n161_));
  OR2        m139(.A(mai_mai_n161_), .B(mai_mai_n158_), .Y(mai_mai_n162_));
  NO2        m140(.A(i_4_), .B(i_5_), .Y(mai_mai_n163_));
  NAi21      m141(.An(i_12_), .B(i_11_), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n164_), .B(i_13_), .Y(mai_mai_n165_));
  NA3        m143(.A(mai_mai_n165_), .B(mai_mai_n163_), .C(mai_mai_n76_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n166_), .B(mai_mai_n162_), .Y(mai_mai_n167_));
  NO2        m145(.A(mai_mai_n67_), .B(mai_mai_n59_), .Y(mai_mai_n168_));
  NA2        m146(.A(mai_mai_n168_), .B(mai_mai_n46_), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n170_));
  NAi31      m148(.An(mai_mai_n170_), .B(mai_mai_n141_), .C(i_11_), .Y(mai_mai_n171_));
  NA2        m149(.A(i_3_), .B(i_5_), .Y(mai_mai_n172_));
  AOI210     m150(.A0(mai_mai_n161_), .A1(mai_mai_n171_), .B0(mai_mai_n169_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n67_), .B(i_5_), .Y(mai_mai_n174_));
  NO2        m152(.A(i_13_), .B(i_10_), .Y(mai_mai_n175_));
  NA3        m153(.A(mai_mai_n175_), .B(mai_mai_n174_), .C(mai_mai_n44_), .Y(mai_mai_n176_));
  NO2        m154(.A(i_2_), .B(i_1_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n177_), .B(i_3_), .Y(mai_mai_n178_));
  NAi21      m156(.An(i_4_), .B(i_12_), .Y(mai_mai_n179_));
  NO3        m157(.A(mai_mai_n179_), .B(mai_mai_n178_), .C(mai_mai_n176_), .Y(mai_mai_n180_));
  NO3        m158(.A(mai_mai_n180_), .B(mai_mai_n173_), .C(mai_mai_n167_), .Y(mai_mai_n181_));
  INV        m159(.A(i_8_), .Y(mai_mai_n182_));
  INV        m160(.A(i_6_), .Y(mai_mai_n183_));
  NO3        m161(.A(i_3_), .B(mai_mai_n79_), .C(mai_mai_n48_), .Y(mai_mai_n184_));
  NA2        m162(.A(mai_mai_n184_), .B(mai_mai_n105_), .Y(mai_mai_n185_));
  NO3        m163(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n186_));
  NA3        m164(.A(mai_mai_n186_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n188_));
  INV        m166(.A(mai_mai_n188_), .Y(mai_mai_n189_));
  AOI210     m167(.A0(mai_mai_n189_), .A1(mai_mai_n187_), .B0(mai_mai_n185_), .Y(mai_mai_n190_));
  NO2        m168(.A(i_3_), .B(i_8_), .Y(mai_mai_n191_));
  NO3        m169(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n192_));
  NA3        m170(.A(mai_mai_n192_), .B(mai_mai_n191_), .C(mai_mai_n40_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n96_), .B(mai_mai_n56_), .Y(mai_mai_n194_));
  NO2        m172(.A(i_13_), .B(i_9_), .Y(mai_mai_n195_));
  NA3        m173(.A(mai_mai_n195_), .B(i_6_), .C(mai_mai_n182_), .Y(mai_mai_n196_));
  BUFFER     m174(.A(mai_mai_n196_), .Y(mai_mai_n197_));
  NO2        m175(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n198_));
  NO3        m176(.A(i_0_), .B(i_2_), .C(mai_mai_n59_), .Y(mai_mai_n199_));
  NA3        m177(.A(mai_mai_n199_), .B(mai_mai_n198_), .C(i_10_), .Y(mai_mai_n200_));
  OAI210     m178(.A0(mai_mai_n200_), .A1(mai_mai_n197_), .B0(mai_mai_n193_), .Y(mai_mai_n201_));
  AOI210     m179(.A0(mai_mai_n201_), .A1(i_7_), .B0(mai_mai_n190_), .Y(mai_mai_n202_));
  OAI220     m180(.A0(mai_mai_n202_), .A1(i_4_), .B0(mai_mai_n183_), .B1(mai_mai_n181_), .Y(mai_mai_n203_));
  NA3        m181(.A(i_13_), .B(mai_mai_n182_), .C(i_10_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n204_), .B(i_12_), .Y(mai_mai_n205_));
  NA2        m183(.A(i_0_), .B(i_5_), .Y(mai_mai_n206_));
  OAI220     m184(.A0(mai_mai_n79_), .A1(mai_mai_n178_), .B0(mai_mai_n169_), .B1(mai_mai_n124_), .Y(mai_mai_n207_));
  NAi31      m185(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n209_));
  NO2        m187(.A(mai_mai_n46_), .B(mai_mai_n59_), .Y(mai_mai_n210_));
  NA3        m188(.A(mai_mai_n210_), .B(i_3_), .C(mai_mai_n209_), .Y(mai_mai_n211_));
  INV        m189(.A(i_13_), .Y(mai_mai_n212_));
  NO2        m190(.A(i_12_), .B(mai_mai_n212_), .Y(mai_mai_n213_));
  NA3        m191(.A(mai_mai_n213_), .B(mai_mai_n186_), .C(mai_mai_n184_), .Y(mai_mai_n214_));
  OAI210     m192(.A0(mai_mai_n211_), .A1(mai_mai_n208_), .B0(mai_mai_n214_), .Y(mai_mai_n215_));
  AOI220     m193(.A0(mai_mai_n215_), .A1(mai_mai_n132_), .B0(mai_mai_n207_), .B1(mai_mai_n205_), .Y(mai_mai_n216_));
  NO2        m194(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n217_));
  NO2        m195(.A(mai_mai_n172_), .B(i_4_), .Y(mai_mai_n218_));
  NA2        m196(.A(mai_mai_n218_), .B(mai_mai_n217_), .Y(mai_mai_n219_));
  OR2        m197(.A(i_8_), .B(i_7_), .Y(mai_mai_n220_));
  NO2        m198(.A(mai_mai_n220_), .B(mai_mai_n79_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n53_), .B(i_1_), .Y(mai_mai_n222_));
  NA2        m200(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n223_));
  INV        m201(.A(i_12_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n44_), .B(mai_mai_n224_), .Y(mai_mai_n225_));
  NO3        m203(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n226_));
  NA2        m204(.A(i_2_), .B(i_1_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n223_), .B(mai_mai_n219_), .Y(mai_mai_n228_));
  NAi21      m206(.An(i_4_), .B(i_3_), .Y(mai_mai_n229_));
  INV        m207(.A(mai_mai_n69_), .Y(mai_mai_n230_));
  NO2        m208(.A(i_0_), .B(i_6_), .Y(mai_mai_n231_));
  NOi41      m209(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n232_));
  NA2        m210(.A(mai_mai_n232_), .B(mai_mai_n231_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n227_), .B(mai_mai_n172_), .Y(mai_mai_n234_));
  NAi21      m212(.An(mai_mai_n233_), .B(mai_mai_n234_), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n235_), .Y(mai_mai_n236_));
  AOI210     m214(.A0(mai_mai_n236_), .A1(mai_mai_n40_), .B0(mai_mai_n228_), .Y(mai_mai_n237_));
  NO2        m215(.A(i_11_), .B(mai_mai_n212_), .Y(mai_mai_n238_));
  NOi21      m216(.An(i_1_), .B(i_6_), .Y(mai_mai_n239_));
  NAi21      m217(.An(i_3_), .B(i_7_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n224_), .B(i_9_), .Y(mai_mai_n241_));
  NO2        m219(.A(i_12_), .B(i_3_), .Y(mai_mai_n242_));
  NA3        m220(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n243_));
  INV        m221(.A(mai_mai_n133_), .Y(mai_mai_n244_));
  NA2        m222(.A(mai_mai_n224_), .B(i_13_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n245_), .B(mai_mai_n69_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n246_), .B(mai_mai_n244_), .Y(mai_mai_n247_));
  NO2        m225(.A(mai_mai_n220_), .B(mai_mai_n37_), .Y(mai_mai_n248_));
  NA2        m226(.A(i_12_), .B(i_6_), .Y(mai_mai_n249_));
  OR2        m227(.A(i_13_), .B(i_9_), .Y(mai_mai_n250_));
  NO3        m228(.A(mai_mai_n250_), .B(mai_mai_n249_), .C(mai_mai_n48_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n229_), .B(i_2_), .Y(mai_mai_n252_));
  NA3        m230(.A(mai_mai_n252_), .B(mai_mai_n251_), .C(mai_mai_n44_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n238_), .B(i_9_), .Y(mai_mai_n254_));
  OAI210     m232(.A0(mai_mai_n59_), .A1(mai_mai_n254_), .B0(mai_mai_n253_), .Y(mai_mai_n255_));
  NA2        m233(.A(mai_mai_n143_), .B(mai_mai_n59_), .Y(mai_mai_n256_));
  NO3        m234(.A(i_11_), .B(mai_mai_n212_), .C(mai_mai_n25_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n240_), .B(i_8_), .Y(mai_mai_n258_));
  NO2        m236(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n259_));
  NA3        m237(.A(mai_mai_n259_), .B(mai_mai_n258_), .C(mai_mai_n257_), .Y(mai_mai_n260_));
  NA3        m238(.A(i_3_), .B(mai_mai_n248_), .C(mai_mai_n213_), .Y(mai_mai_n261_));
  AOI210     m239(.A0(mai_mai_n261_), .A1(mai_mai_n260_), .B0(mai_mai_n256_), .Y(mai_mai_n262_));
  AOI210     m240(.A0(mai_mai_n255_), .A1(mai_mai_n248_), .B0(mai_mai_n262_), .Y(mai_mai_n263_));
  NA4        m241(.A(mai_mai_n263_), .B(mai_mai_n247_), .C(mai_mai_n237_), .D(mai_mai_n216_), .Y(mai_mai_n264_));
  NO3        m242(.A(i_12_), .B(mai_mai_n212_), .C(mai_mai_n37_), .Y(mai_mai_n265_));
  INV        m243(.A(mai_mai_n265_), .Y(mai_mai_n266_));
  NA2        m244(.A(i_8_), .B(mai_mai_n94_), .Y(mai_mai_n267_));
  NO3        m245(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n268_));
  AOI220     m246(.A0(mai_mai_n268_), .A1(mai_mai_n184_), .B0(mai_mai_n152_), .B1(mai_mai_n222_), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n269_), .B(mai_mai_n267_), .Y(mai_mai_n270_));
  NO3        m248(.A(i_0_), .B(i_2_), .C(mai_mai_n59_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n227_), .B(i_0_), .Y(mai_mai_n272_));
  AOI220     m250(.A0(mai_mai_n272_), .A1(mai_mai_n946_), .B0(mai_mai_n271_), .B1(mai_mai_n132_), .Y(mai_mai_n273_));
  NA2        m251(.A(mai_mai_n259_), .B(mai_mai_n26_), .Y(mai_mai_n274_));
  NO2        m252(.A(mai_mai_n274_), .B(mai_mai_n273_), .Y(mai_mai_n275_));
  NA2        m253(.A(i_0_), .B(i_1_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(i_2_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n57_), .B(i_6_), .Y(mai_mai_n278_));
  NA3        m256(.A(mai_mai_n278_), .B(mai_mai_n277_), .C(mai_mai_n152_), .Y(mai_mai_n279_));
  OAI210     m257(.A0(mai_mai_n154_), .A1(mai_mai_n133_), .B0(mai_mai_n279_), .Y(mai_mai_n280_));
  NO3        m258(.A(mai_mai_n280_), .B(mai_mai_n275_), .C(mai_mai_n270_), .Y(mai_mai_n281_));
  NO2        m259(.A(i_3_), .B(i_10_), .Y(mai_mai_n282_));
  NA3        m260(.A(mai_mai_n282_), .B(mai_mai_n40_), .C(mai_mai_n44_), .Y(mai_mai_n283_));
  NO2        m261(.A(i_2_), .B(mai_mai_n94_), .Y(mai_mai_n284_));
  NA2        m262(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n285_), .B(i_8_), .Y(mai_mai_n286_));
  INV        m264(.A(mai_mai_n286_), .Y(mai_mai_n287_));
  AN2        m265(.A(i_3_), .B(i_10_), .Y(mai_mai_n288_));
  NA3        m266(.A(mai_mai_n186_), .B(mai_mai_n165_), .C(mai_mai_n163_), .Y(mai_mai_n289_));
  NO2        m267(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n290_));
  NO2        m268(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n291_));
  OR2        m269(.A(mai_mai_n287_), .B(mai_mai_n283_), .Y(mai_mai_n292_));
  OAI220     m270(.A0(mai_mai_n292_), .A1(i_6_), .B0(mai_mai_n281_), .B1(mai_mai_n266_), .Y(mai_mai_n293_));
  NO4        m271(.A(mai_mai_n293_), .B(mai_mai_n264_), .C(mai_mai_n203_), .D(mai_mai_n157_), .Y(mai_mai_n294_));
  NO3        m272(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n295_));
  NO3        m273(.A(i_6_), .B(mai_mai_n182_), .C(i_7_), .Y(mai_mai_n296_));
  AOI210     m274(.A0(i_1_), .A1(mai_mai_n227_), .B0(mai_mai_n158_), .Y(mai_mai_n297_));
  NO2        m275(.A(i_2_), .B(i_3_), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n206_), .B(i_5_), .Y(mai_mai_n299_));
  NA4        m277(.A(mai_mai_n299_), .B(mai_mai_n221_), .C(mai_mai_n298_), .D(i_1_), .Y(mai_mai_n300_));
  NA3        m278(.A(mai_mai_n272_), .B(mai_mai_n152_), .C(mai_mai_n105_), .Y(mai_mai_n301_));
  NAi21      m279(.An(i_8_), .B(i_7_), .Y(mai_mai_n302_));
  NO2        m280(.A(mai_mai_n302_), .B(i_6_), .Y(mai_mai_n303_));
  NA3        m281(.A(i_2_), .B(mai_mai_n303_), .C(mai_mai_n152_), .Y(mai_mai_n304_));
  NA3        m282(.A(mai_mai_n304_), .B(mai_mai_n301_), .C(mai_mai_n300_), .Y(mai_mai_n305_));
  OAI210     m283(.A0(mai_mai_n305_), .A1(mai_mai_n297_), .B0(i_4_), .Y(mai_mai_n306_));
  NO2        m284(.A(i_12_), .B(i_10_), .Y(mai_mai_n307_));
  NOi21      m285(.An(i_5_), .B(i_0_), .Y(mai_mai_n308_));
  NO3        m286(.A(mai_mai_n285_), .B(mai_mai_n308_), .C(mai_mai_n121_), .Y(mai_mai_n309_));
  NA4        m287(.A(mai_mai_n77_), .B(mai_mai_n36_), .C(mai_mai_n79_), .D(i_8_), .Y(mai_mai_n310_));
  NA2        m288(.A(mai_mai_n309_), .B(mai_mai_n307_), .Y(mai_mai_n311_));
  NO2        m289(.A(i_6_), .B(i_8_), .Y(mai_mai_n312_));
  NOi21      m290(.An(i_0_), .B(i_2_), .Y(mai_mai_n313_));
  AN2        m291(.A(mai_mai_n313_), .B(mai_mai_n312_), .Y(mai_mai_n314_));
  NO2        m292(.A(i_1_), .B(i_7_), .Y(mai_mai_n315_));
  AO220      m293(.A0(mai_mai_n315_), .A1(mai_mai_n314_), .B0(mai_mai_n303_), .B1(mai_mai_n222_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n316_), .B(i_4_), .Y(mai_mai_n317_));
  NA3        m295(.A(mai_mai_n317_), .B(mai_mai_n311_), .C(mai_mai_n306_), .Y(mai_mai_n318_));
  NO3        m296(.A(mai_mai_n220_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n319_));
  NO3        m297(.A(mai_mai_n302_), .B(i_2_), .C(i_1_), .Y(mai_mai_n320_));
  OAI210     m298(.A0(mai_mai_n320_), .A1(mai_mai_n319_), .B0(i_6_), .Y(mai_mai_n321_));
  NA2        m299(.A(mai_mai_n239_), .B(mai_mai_n284_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n322_), .B(mai_mai_n321_), .Y(mai_mai_n323_));
  NA2        m301(.A(mai_mai_n323_), .B(i_3_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n276_), .B(mai_mai_n75_), .Y(mai_mai_n325_));
  NA2        m303(.A(mai_mai_n325_), .B(mai_mai_n123_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n87_), .B(mai_mai_n182_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n87_), .A1(mai_mai_n326_), .B0(i_3_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n182_), .B(i_9_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(mai_mai_n194_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n328_), .B(mai_mai_n275_), .Y(mai_mai_n331_));
  AOI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n324_), .B0(mai_mai_n151_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n318_), .A1(mai_mai_n295_), .B0(mai_mai_n332_), .Y(mai_mai_n333_));
  NOi32      m311(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n334_));
  INV        m312(.A(mai_mai_n334_), .Y(mai_mai_n335_));
  NAi21      m313(.An(i_0_), .B(i_6_), .Y(mai_mai_n336_));
  NAi21      m314(.An(i_1_), .B(i_5_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n337_), .B(mai_mai_n336_), .Y(mai_mai_n338_));
  NA2        m316(.A(mai_mai_n338_), .B(mai_mai_n25_), .Y(mai_mai_n339_));
  OAI210     m317(.A0(mai_mai_n339_), .A1(mai_mai_n148_), .B0(mai_mai_n233_), .Y(mai_mai_n340_));
  NAi41      m318(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n341_));
  OAI220     m319(.A0(mai_mai_n341_), .A1(mai_mai_n337_), .B0(mai_mai_n208_), .B1(mai_mai_n148_), .Y(mai_mai_n342_));
  AOI210     m320(.A0(mai_mai_n341_), .A1(mai_mai_n148_), .B0(mai_mai_n146_), .Y(mai_mai_n343_));
  OR2        m321(.A(mai_mai_n343_), .B(mai_mai_n342_), .Y(mai_mai_n344_));
  NO2        m322(.A(i_1_), .B(mai_mai_n94_), .Y(mai_mai_n345_));
  NAi21      m323(.An(i_3_), .B(i_4_), .Y(mai_mai_n346_));
  NO2        m324(.A(mai_mai_n346_), .B(i_9_), .Y(mai_mai_n347_));
  OAI210     m325(.A0(i_6_), .A1(mai_mai_n345_), .B0(mai_mai_n347_), .Y(mai_mai_n348_));
  NA2        m326(.A(i_2_), .B(i_7_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n346_), .B(i_10_), .Y(mai_mai_n350_));
  NA3        m328(.A(mai_mai_n350_), .B(mai_mai_n349_), .C(mai_mai_n231_), .Y(mai_mai_n351_));
  AOI210     m329(.A0(mai_mai_n351_), .A1(mai_mai_n348_), .B0(mai_mai_n174_), .Y(mai_mai_n352_));
  AOI210     m330(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n177_), .B0(mai_mai_n350_), .Y(mai_mai_n354_));
  AOI220     m332(.A0(mai_mai_n350_), .A1(mai_mai_n315_), .B0(mai_mai_n226_), .B1(mai_mai_n177_), .Y(mai_mai_n355_));
  AOI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n354_), .B0(i_5_), .Y(mai_mai_n356_));
  NO4        m334(.A(mai_mai_n356_), .B(mai_mai_n352_), .C(mai_mai_n344_), .D(mai_mai_n340_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n357_), .B(mai_mai_n335_), .Y(mai_mai_n358_));
  NO2        m336(.A(mai_mai_n57_), .B(mai_mai_n25_), .Y(mai_mai_n359_));
  AN2        m337(.A(i_12_), .B(i_5_), .Y(mai_mai_n360_));
  NO2        m338(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n361_));
  NA2        m339(.A(mai_mai_n361_), .B(mai_mai_n360_), .Y(mai_mai_n362_));
  NO2        m340(.A(i_11_), .B(i_6_), .Y(mai_mai_n363_));
  NA3        m341(.A(mai_mai_n363_), .B(i_2_), .C(mai_mai_n212_), .Y(mai_mai_n364_));
  NO2        m342(.A(mai_mai_n364_), .B(mai_mai_n362_), .Y(mai_mai_n365_));
  INV        m343(.A(i_5_), .Y(mai_mai_n366_));
  NO2        m344(.A(i_5_), .B(i_10_), .Y(mai_mai_n367_));
  AOI220     m345(.A0(mai_mai_n367_), .A1(mai_mai_n252_), .B0(mai_mai_n366_), .B1(mai_mai_n186_), .Y(mai_mai_n368_));
  NA2        m346(.A(mai_mai_n134_), .B(mai_mai_n45_), .Y(mai_mai_n369_));
  NO2        m347(.A(mai_mai_n369_), .B(mai_mai_n368_), .Y(mai_mai_n370_));
  OAI210     m348(.A0(mai_mai_n370_), .A1(mai_mai_n365_), .B0(mai_mai_n359_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n372_));
  NO2        m350(.A(mai_mai_n140_), .B(mai_mai_n79_), .Y(mai_mai_n373_));
  OAI210     m351(.A0(mai_mai_n373_), .A1(mai_mai_n365_), .B0(mai_mai_n372_), .Y(mai_mai_n374_));
  NO3        m352(.A(mai_mai_n79_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n367_), .B(mai_mai_n224_), .Y(mai_mai_n376_));
  OAI210     m354(.A0(mai_mai_n376_), .A1(mai_mai_n310_), .B0(mai_mai_n208_), .Y(mai_mai_n377_));
  NAi21      m355(.An(i_13_), .B(i_0_), .Y(mai_mai_n378_));
  NO2        m356(.A(mai_mai_n378_), .B(mai_mai_n227_), .Y(mai_mai_n379_));
  NA2        m357(.A(mai_mai_n377_), .B(mai_mai_n379_), .Y(mai_mai_n380_));
  NA3        m358(.A(mai_mai_n380_), .B(mai_mai_n374_), .C(mai_mai_n371_), .Y(mai_mai_n381_));
  NA2        m359(.A(mai_mai_n44_), .B(mai_mai_n212_), .Y(mai_mai_n382_));
  NO2        m360(.A(i_0_), .B(i_11_), .Y(mai_mai_n383_));
  INV        m361(.A(i_5_), .Y(mai_mai_n384_));
  AN2        m362(.A(i_1_), .B(i_6_), .Y(mai_mai_n385_));
  NOi21      m363(.An(i_2_), .B(i_12_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n386_), .B(mai_mai_n385_), .Y(mai_mai_n387_));
  NO2        m365(.A(mai_mai_n387_), .B(mai_mai_n384_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n132_), .B(i_9_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n389_), .B(i_4_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n388_), .B(mai_mai_n390_), .Y(mai_mai_n391_));
  NAi21      m369(.An(i_9_), .B(i_4_), .Y(mai_mai_n392_));
  OR2        m370(.A(i_13_), .B(i_10_), .Y(mai_mai_n393_));
  NO3        m371(.A(mai_mai_n393_), .B(mai_mai_n110_), .C(mai_mai_n392_), .Y(mai_mai_n394_));
  BUFFER     m372(.A(mai_mai_n204_), .Y(mai_mai_n395_));
  NO2        m373(.A(mai_mai_n94_), .B(mai_mai_n25_), .Y(mai_mai_n396_));
  NA2        m374(.A(mai_mai_n259_), .B(mai_mai_n199_), .Y(mai_mai_n397_));
  NO2        m375(.A(mai_mai_n397_), .B(mai_mai_n395_), .Y(mai_mai_n398_));
  INV        m376(.A(mai_mai_n398_), .Y(mai_mai_n399_));
  AOI210     m377(.A0(mai_mai_n399_), .A1(mai_mai_n391_), .B0(mai_mai_n26_), .Y(mai_mai_n400_));
  NA2        m378(.A(mai_mai_n301_), .B(mai_mai_n300_), .Y(mai_mai_n401_));
  AOI220     m379(.A0(mai_mai_n278_), .A1(mai_mai_n268_), .B0(mai_mai_n272_), .B1(i_6_), .Y(mai_mai_n402_));
  NO2        m380(.A(mai_mai_n402_), .B(mai_mai_n158_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n172_), .B(mai_mai_n79_), .Y(mai_mai_n404_));
  AOI220     m382(.A0(mai_mai_n404_), .A1(mai_mai_n277_), .B0(i_3_), .B1(mai_mai_n199_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n405_), .B(mai_mai_n267_), .Y(mai_mai_n406_));
  NO3        m384(.A(mai_mai_n406_), .B(mai_mai_n403_), .C(mai_mai_n401_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n184_), .B(mai_mai_n89_), .Y(mai_mai_n408_));
  NA3        m386(.A(i_2_), .B(mai_mai_n152_), .C(mai_mai_n79_), .Y(mai_mai_n409_));
  AOI210     m387(.A0(mai_mai_n409_), .A1(mai_mai_n408_), .B0(mai_mai_n302_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n278_), .B(mai_mai_n222_), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n411_), .B(mai_mai_n172_), .Y(mai_mai_n412_));
  NA3        m390(.A(mai_mai_n315_), .B(mai_mai_n314_), .C(i_5_), .Y(mai_mai_n413_));
  INV        m391(.A(mai_mai_n296_), .Y(mai_mai_n414_));
  OAI210     m392(.A0(mai_mai_n414_), .A1(mai_mai_n178_), .B0(mai_mai_n413_), .Y(mai_mai_n415_));
  NO3        m393(.A(mai_mai_n415_), .B(mai_mai_n412_), .C(mai_mai_n410_), .Y(mai_mai_n416_));
  AOI210     m394(.A0(mai_mai_n416_), .A1(mai_mai_n407_), .B0(mai_mai_n254_), .Y(mai_mai_n417_));
  NO4        m395(.A(mai_mai_n417_), .B(mai_mai_n400_), .C(mai_mai_n381_), .D(mai_mai_n358_), .Y(mai_mai_n418_));
  NO2        m396(.A(mai_mai_n67_), .B(i_13_), .Y(mai_mai_n419_));
  NA2        m397(.A(mai_mai_n419_), .B(i_2_), .Y(mai_mai_n420_));
  NO2        m398(.A(i_10_), .B(i_9_), .Y(mai_mai_n421_));
  NAi21      m399(.An(i_12_), .B(i_8_), .Y(mai_mai_n422_));
  NO2        m400(.A(mai_mai_n422_), .B(i_3_), .Y(mai_mai_n423_));
  NA2        m401(.A(mai_mai_n423_), .B(mai_mai_n421_), .Y(mai_mai_n424_));
  NA2        m402(.A(i_2_), .B(mai_mai_n97_), .Y(mai_mai_n425_));
  OAI220     m403(.A0(mai_mai_n425_), .A1(mai_mai_n193_), .B0(mai_mai_n424_), .B1(mai_mai_n420_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n291_), .B(i_0_), .Y(mai_mai_n427_));
  NO3        m405(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n428_));
  NA2        m406(.A(mai_mai_n249_), .B(mai_mai_n90_), .Y(mai_mai_n429_));
  NA2        m407(.A(mai_mai_n429_), .B(mai_mai_n428_), .Y(mai_mai_n430_));
  NA2        m408(.A(i_8_), .B(i_9_), .Y(mai_mai_n431_));
  NO2        m409(.A(i_7_), .B(i_2_), .Y(mai_mai_n432_));
  OR2        m410(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  NA2        m411(.A(mai_mai_n265_), .B(mai_mai_n194_), .Y(mai_mai_n434_));
  NO2        m412(.A(mai_mai_n434_), .B(mai_mai_n433_), .Y(mai_mai_n435_));
  NA2        m413(.A(mai_mai_n238_), .B(mai_mai_n290_), .Y(mai_mai_n436_));
  NO3        m414(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n437_));
  INV        m415(.A(mai_mai_n437_), .Y(mai_mai_n438_));
  NA3        m416(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n439_));
  NA3        m417(.A(mai_mai_n135_), .B(mai_mai_n108_), .C(mai_mai_n23_), .Y(mai_mai_n440_));
  OAI220     m418(.A0(mai_mai_n440_), .A1(mai_mai_n439_), .B0(mai_mai_n438_), .B1(mai_mai_n436_), .Y(mai_mai_n441_));
  NO3        m419(.A(mai_mai_n441_), .B(mai_mai_n435_), .C(mai_mai_n426_), .Y(mai_mai_n442_));
  OR2        m420(.A(mai_mai_n276_), .B(mai_mai_n196_), .Y(mai_mai_n443_));
  OA210      m421(.A0(mai_mai_n330_), .A1(mai_mai_n94_), .B0(mai_mai_n279_), .Y(mai_mai_n444_));
  OA220      m422(.A0(mai_mai_n444_), .A1(mai_mai_n151_), .B0(mai_mai_n443_), .B1(mai_mai_n219_), .Y(mai_mai_n445_));
  NA2        m423(.A(mai_mai_n89_), .B(i_13_), .Y(mai_mai_n446_));
  NA2        m424(.A(mai_mai_n404_), .B(mai_mai_n359_), .Y(mai_mai_n447_));
  NO2        m425(.A(i_2_), .B(i_13_), .Y(mai_mai_n448_));
  NA3        m426(.A(mai_mai_n448_), .B(mai_mai_n150_), .C(mai_mai_n92_), .Y(mai_mai_n449_));
  NO2        m427(.A(mai_mai_n447_), .B(mai_mai_n446_), .Y(mai_mai_n450_));
  NO3        m428(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n451_));
  NO2        m429(.A(i_6_), .B(i_7_), .Y(mai_mai_n452_));
  OR2        m430(.A(i_11_), .B(i_8_), .Y(mai_mai_n453_));
  NOi21      m431(.An(i_2_), .B(i_7_), .Y(mai_mai_n454_));
  NAi31      m432(.An(mai_mai_n453_), .B(mai_mai_n454_), .C(mai_mai_n945_), .Y(mai_mai_n455_));
  NO2        m433(.A(mai_mai_n393_), .B(i_6_), .Y(mai_mai_n456_));
  NA2        m434(.A(mai_mai_n456_), .B(mai_mai_n950_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n457_), .B(mai_mai_n455_), .Y(mai_mai_n458_));
  NO2        m436(.A(i_3_), .B(mai_mai_n182_), .Y(mai_mai_n459_));
  NO2        m437(.A(i_6_), .B(i_10_), .Y(mai_mai_n460_));
  NA2        m438(.A(mai_mai_n46_), .B(mai_mai_n44_), .Y(mai_mai_n461_));
  NO2        m439(.A(mai_mai_n146_), .B(i_3_), .Y(mai_mai_n462_));
  NAi31      m440(.An(mai_mai_n461_), .B(mai_mai_n462_), .C(mai_mai_n213_), .Y(mai_mai_n463_));
  NA3        m441(.A(mai_mai_n372_), .B(mai_mai_n168_), .C(mai_mai_n139_), .Y(mai_mai_n464_));
  NA2        m442(.A(mai_mai_n464_), .B(mai_mai_n463_), .Y(mai_mai_n465_));
  NO3        m443(.A(mai_mai_n465_), .B(mai_mai_n458_), .C(mai_mai_n450_), .Y(mai_mai_n466_));
  NA2        m444(.A(mai_mai_n428_), .B(mai_mai_n360_), .Y(mai_mai_n467_));
  NA2        m445(.A(mai_mai_n437_), .B(mai_mai_n367_), .Y(mai_mai_n468_));
  NO2        m446(.A(mai_mai_n468_), .B(mai_mai_n211_), .Y(mai_mai_n469_));
  NO2        m447(.A(i_0_), .B(mai_mai_n79_), .Y(mai_mai_n470_));
  NA3        m448(.A(mai_mai_n470_), .B(i_3_), .C(mai_mai_n132_), .Y(mai_mai_n471_));
  OR3        m449(.A(mai_mai_n285_), .B(mai_mai_n38_), .C(mai_mai_n46_), .Y(mai_mai_n472_));
  NO2        m450(.A(mai_mai_n472_), .B(mai_mai_n471_), .Y(mai_mai_n473_));
  NA2        m451(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n474_));
  NO2        m452(.A(mai_mai_n474_), .B(mai_mai_n446_), .Y(mai_mai_n475_));
  NO3        m453(.A(mai_mai_n475_), .B(mai_mai_n473_), .C(mai_mai_n469_), .Y(mai_mai_n476_));
  NA4        m454(.A(mai_mai_n476_), .B(mai_mai_n466_), .C(mai_mai_n445_), .D(mai_mai_n442_), .Y(mai_mai_n477_));
  NA3        m455(.A(mai_mai_n288_), .B(mai_mai_n165_), .C(mai_mai_n163_), .Y(mai_mai_n478_));
  INV        m456(.A(mai_mai_n478_), .Y(mai_mai_n479_));
  BUFFER     m457(.A(mai_mai_n221_), .Y(mai_mai_n480_));
  NA2        m458(.A(mai_mai_n480_), .B(mai_mai_n479_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n115_), .B(mai_mai_n104_), .Y(mai_mai_n482_));
  AN2        m460(.A(mai_mai_n482_), .B(mai_mai_n428_), .Y(mai_mai_n483_));
  NA2        m461(.A(mai_mai_n295_), .B(mai_mai_n153_), .Y(mai_mai_n484_));
  OAI210     m462(.A0(mai_mai_n484_), .A1(mai_mai_n219_), .B0(mai_mai_n289_), .Y(mai_mai_n485_));
  AOI220     m463(.A0(mai_mai_n485_), .A1(mai_mai_n303_), .B0(mai_mai_n483_), .B1(mai_mai_n291_), .Y(mai_mai_n486_));
  NA4        m464(.A(mai_mai_n419_), .B(mai_mai_n950_), .C(mai_mai_n191_), .D(i_2_), .Y(mai_mai_n487_));
  INV        m465(.A(mai_mai_n487_), .Y(mai_mai_n488_));
  NA2        m466(.A(mai_mai_n334_), .B(mai_mai_n67_), .Y(mai_mai_n489_));
  NO2        m467(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n490_));
  AOI210     m468(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n394_), .Y(mai_mai_n491_));
  INV        m469(.A(mai_mai_n491_), .Y(mai_mai_n492_));
  AOI210     m470(.A0(mai_mai_n488_), .A1(mai_mai_n192_), .B0(mai_mai_n492_), .Y(mai_mai_n493_));
  NO2        m471(.A(i_7_), .B(mai_mai_n187_), .Y(mai_mai_n494_));
  OR2        m472(.A(mai_mai_n172_), .B(i_4_), .Y(mai_mai_n495_));
  INV        m473(.A(mai_mai_n495_), .Y(mai_mai_n496_));
  NA2        m474(.A(mai_mai_n496_), .B(mai_mai_n494_), .Y(mai_mai_n497_));
  NA4        m475(.A(mai_mai_n497_), .B(mai_mai_n493_), .C(mai_mai_n486_), .D(mai_mai_n481_), .Y(mai_mai_n498_));
  NA2        m476(.A(mai_mai_n366_), .B(mai_mai_n277_), .Y(mai_mai_n499_));
  NA2        m477(.A(mai_mai_n362_), .B(mai_mai_n499_), .Y(mai_mai_n500_));
  NO2        m478(.A(i_12_), .B(mai_mai_n182_), .Y(mai_mai_n501_));
  NA2        m479(.A(mai_mai_n501_), .B(mai_mai_n212_), .Y(mai_mai_n502_));
  NA2        m480(.A(mai_mai_n460_), .B(mai_mai_n27_), .Y(mai_mai_n503_));
  NO2        m481(.A(mai_mai_n503_), .B(mai_mai_n502_), .Y(mai_mai_n504_));
  NOi21      m482(.An(mai_mai_n296_), .B(mai_mai_n38_), .Y(mai_mai_n505_));
  OAI210     m483(.A0(mai_mai_n505_), .A1(mai_mai_n504_), .B0(mai_mai_n500_), .Y(mai_mai_n506_));
  NO2        m484(.A(i_8_), .B(i_7_), .Y(mai_mai_n507_));
  INV        m485(.A(mai_mai_n210_), .Y(mai_mai_n508_));
  OAI220     m486(.A0(mai_mai_n46_), .A1(mai_mai_n495_), .B0(mai_mai_n508_), .B1(mai_mai_n229_), .Y(mai_mai_n509_));
  NO2        m487(.A(mai_mai_n949_), .B(i_6_), .Y(mai_mai_n510_));
  NA3        m488(.A(mai_mai_n510_), .B(mai_mai_n509_), .C(mai_mai_n507_), .Y(mai_mai_n511_));
  AOI220     m489(.A0(mai_mai_n404_), .A1(i_2_), .B0(mai_mai_n234_), .B1(mai_mai_n231_), .Y(mai_mai_n512_));
  OAI220     m490(.A0(mai_mai_n512_), .A1(mai_mai_n245_), .B0(mai_mai_n446_), .B1(mai_mai_n124_), .Y(mai_mai_n513_));
  NA2        m491(.A(mai_mai_n513_), .B(mai_mai_n248_), .Y(mai_mai_n514_));
  NA3        m492(.A(mai_mai_n288_), .B(mai_mai_n163_), .C(mai_mai_n89_), .Y(mai_mai_n515_));
  NO2        m493(.A(mai_mai_n209_), .B(mai_mai_n44_), .Y(mai_mai_n516_));
  NO2        m494(.A(mai_mai_n146_), .B(i_5_), .Y(mai_mai_n517_));
  NA2        m495(.A(mai_mai_n517_), .B(mai_mai_n382_), .Y(mai_mai_n518_));
  NO2        m496(.A(mai_mai_n518_), .B(mai_mai_n516_), .Y(mai_mai_n519_));
  NA2        m497(.A(mai_mai_n519_), .B(mai_mai_n437_), .Y(mai_mai_n520_));
  NA4        m498(.A(mai_mai_n520_), .B(mai_mai_n514_), .C(mai_mai_n511_), .D(mai_mai_n506_), .Y(mai_mai_n521_));
  NA3        m499(.A(mai_mai_n206_), .B(mai_mai_n65_), .C(mai_mai_n44_), .Y(mai_mai_n522_));
  NA2        m500(.A(mai_mai_n265_), .B(mai_mai_n77_), .Y(mai_mai_n523_));
  AOI210     m501(.A0(mai_mai_n522_), .A1(mai_mai_n326_), .B0(mai_mai_n523_), .Y(mai_mai_n524_));
  AOI210     m502(.A0(i_6_), .A1(mai_mai_n46_), .B0(mai_mai_n345_), .Y(mai_mai_n525_));
  NA2        m503(.A(mai_mai_n501_), .B(mai_mai_n257_), .Y(mai_mai_n526_));
  NO2        m504(.A(mai_mai_n525_), .B(mai_mai_n526_), .Y(mai_mai_n527_));
  NO2        m505(.A(mai_mai_n527_), .B(mai_mai_n524_), .Y(mai_mai_n528_));
  NO4        m506(.A(mai_mai_n239_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n529_));
  NO3        m507(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n530_));
  NO2        m508(.A(mai_mai_n220_), .B(mai_mai_n36_), .Y(mai_mai_n531_));
  AN2        m509(.A(mai_mai_n531_), .B(mai_mai_n530_), .Y(mai_mai_n532_));
  OA210      m510(.A0(mai_mai_n532_), .A1(mai_mai_n529_), .B0(mai_mai_n334_), .Y(mai_mai_n533_));
  NO2        m511(.A(mai_mai_n393_), .B(i_1_), .Y(mai_mai_n534_));
  NOi31      m512(.An(mai_mai_n534_), .B(mai_mai_n429_), .C(mai_mai_n67_), .Y(mai_mai_n535_));
  AN3        m513(.A(mai_mai_n535_), .B(mai_mai_n390_), .C(i_2_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n402_), .B(mai_mai_n166_), .Y(mai_mai_n537_));
  NO3        m515(.A(mai_mai_n537_), .B(mai_mai_n536_), .C(mai_mai_n533_), .Y(mai_mai_n538_));
  NOi21      m516(.An(i_10_), .B(i_6_), .Y(mai_mai_n539_));
  NA2        m517(.A(mai_mai_n257_), .B(mai_mai_n539_), .Y(mai_mai_n540_));
  NO2        m518(.A(mai_mai_n540_), .B(mai_mai_n427_), .Y(mai_mai_n541_));
  NO2        m519(.A(mai_mai_n107_), .B(mai_mai_n23_), .Y(mai_mai_n542_));
  NA2        m520(.A(mai_mai_n296_), .B(mai_mai_n153_), .Y(mai_mai_n543_));
  AOI220     m521(.A0(mai_mai_n543_), .A1(mai_mai_n411_), .B0(mai_mai_n161_), .B1(mai_mai_n171_), .Y(mai_mai_n544_));
  NO2        m522(.A(mai_mai_n186_), .B(mai_mai_n37_), .Y(mai_mai_n545_));
  NOi31      m523(.An(mai_mai_n136_), .B(mai_mai_n545_), .C(mai_mai_n310_), .Y(mai_mai_n546_));
  NO3        m524(.A(mai_mai_n546_), .B(mai_mai_n544_), .C(mai_mai_n541_), .Y(mai_mai_n547_));
  NO2        m525(.A(mai_mai_n489_), .B(mai_mai_n355_), .Y(mai_mai_n548_));
  NO2        m526(.A(i_12_), .B(mai_mai_n79_), .Y(mai_mai_n549_));
  NO3        m527(.A(i_4_), .B(mai_mai_n321_), .C(mai_mai_n283_), .Y(mai_mai_n550_));
  BUFFER     m528(.A(i_5_), .Y(mai_mai_n551_));
  NO2        m529(.A(mai_mai_n550_), .B(mai_mai_n548_), .Y(mai_mai_n552_));
  NA4        m530(.A(mai_mai_n552_), .B(mai_mai_n547_), .C(mai_mai_n538_), .D(mai_mai_n528_), .Y(mai_mai_n553_));
  NO4        m531(.A(mai_mai_n553_), .B(mai_mai_n521_), .C(mai_mai_n498_), .D(mai_mai_n477_), .Y(mai_mai_n554_));
  NA4        m532(.A(mai_mai_n554_), .B(mai_mai_n418_), .C(mai_mai_n333_), .D(mai_mai_n294_), .Y(mai7));
  NO2        m533(.A(mai_mai_n101_), .B(mai_mai_n84_), .Y(mai_mai_n556_));
  NA2        m534(.A(mai_mai_n460_), .B(mai_mai_n77_), .Y(mai_mai_n557_));
  NA3        m535(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n558_));
  NO2        m536(.A(mai_mai_n224_), .B(i_4_), .Y(mai_mai_n559_));
  NA2        m537(.A(mai_mai_n559_), .B(i_8_), .Y(mai_mai_n560_));
  NO2        m538(.A(mai_mai_n98_), .B(mai_mai_n558_), .Y(mai_mai_n561_));
  OAI210     m539(.A0(mai_mai_n82_), .A1(mai_mai_n191_), .B0(mai_mai_n192_), .Y(mai_mai_n562_));
  NO2        m540(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n563_));
  NO2        m541(.A(mai_mai_n562_), .B(i_13_), .Y(mai_mai_n564_));
  NO3        m542(.A(mai_mai_n564_), .B(mai_mai_n561_), .C(mai_mai_n556_), .Y(mai_mai_n565_));
  AOI210     m543(.A0(mai_mai_n121_), .A1(mai_mai_n58_), .B0(i_10_), .Y(mai_mai_n566_));
  AOI210     m544(.A0(mai_mai_n566_), .A1(mai_mai_n224_), .B0(mai_mai_n150_), .Y(mai_mai_n567_));
  NO2        m545(.A(i_10_), .B(mai_mai_n23_), .Y(mai_mai_n568_));
  OR3        m546(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n569_));
  NO3        m547(.A(mai_mai_n569_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n570_));
  INV        m548(.A(mai_mai_n188_), .Y(mai_mai_n571_));
  NO2        m549(.A(mai_mai_n570_), .B(mai_mai_n568_), .Y(mai_mai_n572_));
  OA220      m550(.A0(mai_mai_n572_), .A1(i_2_), .B0(mai_mai_n567_), .B1(mai_mai_n250_), .Y(mai_mai_n573_));
  AOI210     m551(.A0(mai_mai_n573_), .A1(mai_mai_n565_), .B0(mai_mai_n59_), .Y(mai_mai_n574_));
  NOi21      m552(.An(i_11_), .B(i_7_), .Y(mai_mai_n575_));
  AO210      m553(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n576_));
  NO2        m554(.A(mai_mai_n576_), .B(mai_mai_n575_), .Y(mai_mai_n577_));
  NA2        m555(.A(mai_mai_n577_), .B(mai_mai_n195_), .Y(mai_mai_n578_));
  NA3        m556(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n579_));
  NO2        m557(.A(mai_mai_n578_), .B(mai_mai_n59_), .Y(mai_mai_n580_));
  AO210      m558(.A0(mai_mai_n80_), .A1(mai_mai_n355_), .B0(mai_mai_n41_), .Y(mai_mai_n581_));
  NA2        m559(.A(mai_mai_n213_), .B(mai_mai_n59_), .Y(mai_mai_n582_));
  NO2        m560(.A(mai_mai_n59_), .B(i_9_), .Y(mai_mai_n583_));
  NO2        m561(.A(i_1_), .B(i_12_), .Y(mai_mai_n584_));
  NA2        m562(.A(mai_mai_n582_), .B(mai_mai_n581_), .Y(mai_mai_n585_));
  OAI210     m563(.A0(mai_mai_n585_), .A1(mai_mai_n580_), .B0(i_6_), .Y(mai_mai_n586_));
  NO2        m564(.A(mai_mai_n579_), .B(mai_mai_n101_), .Y(mai_mai_n587_));
  NA2        m565(.A(mai_mai_n587_), .B(mai_mai_n549_), .Y(mai_mai_n588_));
  NO2        m566(.A(i_6_), .B(i_11_), .Y(mai_mai_n589_));
  NA2        m567(.A(mai_mai_n588_), .B(mai_mai_n430_), .Y(mai_mai_n590_));
  NO4        m568(.A(i_12_), .B(mai_mai_n121_), .C(i_13_), .D(mai_mai_n79_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n591_), .B(mai_mai_n583_), .Y(mai_mai_n592_));
  NO3        m570(.A(i_10_), .B(mai_mai_n220_), .C(mai_mai_n23_), .Y(mai_mai_n593_));
  INV        m571(.A(mai_mai_n592_), .Y(mai_mai_n594_));
  NA3        m572(.A(mai_mai_n507_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n595_));
  NA2        m573(.A(mai_mai_n128_), .B(i_9_), .Y(mai_mai_n596_));
  NA2        m574(.A(i_3_), .B(i_9_), .Y(mai_mai_n597_));
  NO2        m575(.A(mai_mai_n596_), .B(mai_mai_n944_), .Y(mai_mai_n598_));
  NA3        m576(.A(mai_mai_n583_), .B(mai_mai_n298_), .C(i_6_), .Y(mai_mai_n599_));
  NO2        m577(.A(mai_mai_n599_), .B(mai_mai_n23_), .Y(mai_mai_n600_));
  NO2        m578(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n601_));
  NA2        m579(.A(mai_mai_n601_), .B(mai_mai_n24_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n602_), .B(i_6_), .Y(mai_mai_n603_));
  OR3        m581(.A(mai_mai_n603_), .B(mai_mai_n600_), .C(mai_mai_n598_), .Y(mai_mai_n604_));
  NO3        m582(.A(mai_mai_n604_), .B(mai_mai_n594_), .C(mai_mai_n590_), .Y(mai_mai_n605_));
  NO2        m583(.A(mai_mai_n392_), .B(mai_mai_n79_), .Y(mai_mai_n606_));
  NO2        m584(.A(mai_mai_n220_), .B(mai_mai_n44_), .Y(mai_mai_n607_));
  NO3        m585(.A(mai_mai_n607_), .B(mai_mai_n291_), .C(mai_mai_n225_), .Y(mai_mai_n608_));
  NO2        m586(.A(mai_mai_n110_), .B(mai_mai_n37_), .Y(mai_mai_n609_));
  NO2        m587(.A(mai_mai_n609_), .B(i_6_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n79_), .B(i_9_), .Y(mai_mai_n611_));
  NO2        m589(.A(mai_mai_n611_), .B(mai_mai_n59_), .Y(mai_mai_n612_));
  NO2        m590(.A(mai_mai_n612_), .B(mai_mai_n584_), .Y(mai_mai_n613_));
  NO4        m591(.A(mai_mai_n613_), .B(mai_mai_n610_), .C(mai_mai_n608_), .D(i_4_), .Y(mai_mai_n614_));
  NA2        m592(.A(i_1_), .B(i_3_), .Y(mai_mai_n615_));
  INV        m593(.A(mai_mai_n614_), .Y(mai_mai_n616_));
  NA3        m594(.A(mai_mai_n616_), .B(mai_mai_n605_), .C(mai_mai_n586_), .Y(mai_mai_n617_));
  NO3        m595(.A(mai_mai_n453_), .B(i_3_), .C(i_7_), .Y(mai_mai_n618_));
  OA210      m596(.A0(mai_mai_n618_), .A1(mai_mai_n232_), .B0(mai_mai_n79_), .Y(mai_mai_n619_));
  NA3        m597(.A(mai_mai_n150_), .B(mai_mai_n77_), .C(mai_mai_n79_), .Y(mai_mai_n620_));
  INV        m598(.A(mai_mai_n620_), .Y(mai_mai_n621_));
  OAI210     m599(.A0(mai_mai_n621_), .A1(mai_mai_n619_), .B0(i_1_), .Y(mai_mai_n622_));
  AOI210     m600(.A0(mai_mai_n249_), .A1(mai_mai_n90_), .B0(i_1_), .Y(mai_mai_n623_));
  NO2        m601(.A(mai_mai_n346_), .B(i_2_), .Y(mai_mai_n624_));
  NA2        m602(.A(mai_mai_n624_), .B(mai_mai_n623_), .Y(mai_mai_n625_));
  AOI210     m603(.A0(mai_mai_n625_), .A1(mai_mai_n622_), .B0(i_13_), .Y(mai_mai_n626_));
  OR2        m604(.A(i_11_), .B(i_7_), .Y(mai_mai_n627_));
  NA2        m605(.A(mai_mai_n99_), .B(mai_mai_n128_), .Y(mai_mai_n628_));
  AOI220     m606(.A0(mai_mai_n448_), .A1(mai_mai_n150_), .B0(i_2_), .B1(mai_mai_n128_), .Y(mai_mai_n629_));
  NA2        m607(.A(mai_mai_n629_), .B(mai_mai_n628_), .Y(mai_mai_n630_));
  NO2        m608(.A(mai_mai_n54_), .B(i_12_), .Y(mai_mai_n631_));
  INV        m609(.A(mai_mai_n631_), .Y(mai_mai_n632_));
  NO2        m610(.A(mai_mai_n454_), .B(mai_mai_n24_), .Y(mai_mai_n633_));
  NA2        m611(.A(mai_mai_n633_), .B(mai_mai_n606_), .Y(mai_mai_n634_));
  OAI220     m612(.A0(mai_mai_n634_), .A1(mai_mai_n41_), .B0(mai_mai_n632_), .B1(mai_mai_n87_), .Y(mai_mai_n635_));
  AOI210     m613(.A0(mai_mai_n630_), .A1(mai_mai_n312_), .B0(mai_mai_n635_), .Y(mai_mai_n636_));
  INV        m614(.A(mai_mai_n107_), .Y(mai_mai_n637_));
  AOI220     m615(.A0(mai_mai_n637_), .A1(mai_mai_n66_), .B0(mai_mai_n363_), .B1(mai_mai_n951_), .Y(mai_mai_n638_));
  NO2        m616(.A(mai_mai_n638_), .B(mai_mai_n229_), .Y(mai_mai_n639_));
  AOI210     m617(.A0(mai_mai_n422_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n640_));
  NOi21      m618(.An(mai_mai_n640_), .B(mai_mai_n557_), .Y(mai_mai_n641_));
  NA2        m619(.A(mai_mai_n120_), .B(i_13_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n597_), .B(mai_mai_n107_), .Y(mai_mai_n643_));
  NO2        m621(.A(mai_mai_n642_), .B(mai_mai_n623_), .Y(mai_mai_n644_));
  AOI220     m622(.A0(mai_mai_n363_), .A1(mai_mai_n951_), .B0(mai_mai_n86_), .B1(mai_mai_n95_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n645_), .B(mai_mai_n560_), .Y(mai_mai_n646_));
  NO4        m624(.A(mai_mai_n646_), .B(mai_mai_n644_), .C(mai_mai_n641_), .D(mai_mai_n639_), .Y(mai_mai_n647_));
  OR2        m625(.A(i_11_), .B(i_6_), .Y(mai_mai_n648_));
  NO2        m626(.A(mai_mai_n597_), .B(mai_mai_n648_), .Y(mai_mai_n649_));
  NA3        m627(.A(mai_mai_n386_), .B(mai_mai_n563_), .C(mai_mai_n90_), .Y(mai_mai_n650_));
  NA2        m628(.A(mai_mai_n589_), .B(i_13_), .Y(mai_mai_n651_));
  NAi21      m629(.An(i_11_), .B(i_12_), .Y(mai_mai_n652_));
  NA2        m630(.A(mai_mai_n651_), .B(mai_mai_n650_), .Y(mai_mai_n653_));
  OAI210     m631(.A0(mai_mai_n653_), .A1(mai_mai_n649_), .B0(mai_mai_n59_), .Y(mai_mai_n654_));
  NO2        m632(.A(i_2_), .B(i_12_), .Y(mai_mai_n655_));
  NA2        m633(.A(mai_mai_n345_), .B(mai_mai_n655_), .Y(mai_mai_n656_));
  NO3        m634(.A(i_9_), .B(mai_mai_n361_), .C(mai_mai_n559_), .Y(mai_mai_n657_));
  NA2        m635(.A(mai_mai_n657_), .B(mai_mai_n345_), .Y(mai_mai_n658_));
  NO2        m636(.A(mai_mai_n121_), .B(i_2_), .Y(mai_mai_n659_));
  NA2        m637(.A(mai_mai_n659_), .B(mai_mai_n584_), .Y(mai_mai_n660_));
  NA3        m638(.A(mai_mai_n660_), .B(mai_mai_n658_), .C(mai_mai_n656_), .Y(mai_mai_n661_));
  NA3        m639(.A(mai_mai_n661_), .B(mai_mai_n45_), .C(mai_mai_n212_), .Y(mai_mai_n662_));
  NA4        m640(.A(mai_mai_n662_), .B(mai_mai_n654_), .C(mai_mai_n647_), .D(mai_mai_n636_), .Y(mai_mai_n663_));
  OR4        m641(.A(mai_mai_n663_), .B(mai_mai_n626_), .C(mai_mai_n617_), .D(mai_mai_n574_), .Y(mai5));
  AN2        m642(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n665_));
  NA3        m643(.A(mai_mai_n665_), .B(mai_mai_n655_), .C(mai_mai_n101_), .Y(mai_mai_n666_));
  INV        m644(.A(mai_mai_n666_), .Y(mai_mai_n667_));
  NO3        m645(.A(i_11_), .B(mai_mai_n224_), .C(i_13_), .Y(mai_mai_n668_));
  NO2        m646(.A(mai_mai_n117_), .B(mai_mai_n23_), .Y(mai_mai_n669_));
  NA2        m647(.A(i_12_), .B(i_8_), .Y(mai_mai_n670_));
  INV        m648(.A(mai_mai_n421_), .Y(mai_mai_n671_));
  NA2        m649(.A(i_2_), .B(mai_mai_n669_), .Y(mai_mai_n672_));
  INV        m650(.A(mai_mai_n672_), .Y(mai_mai_n673_));
  NO2        m651(.A(mai_mai_n673_), .B(mai_mai_n667_), .Y(mai_mai_n674_));
  INV        m652(.A(mai_mai_n160_), .Y(mai_mai_n675_));
  INV        m653(.A(mai_mai_n232_), .Y(mai_mai_n676_));
  OAI210     m654(.A0(mai_mai_n624_), .A1(mai_mai_n423_), .B0(mai_mai_n103_), .Y(mai_mai_n677_));
  AOI210     m655(.A0(mai_mai_n677_), .A1(mai_mai_n676_), .B0(mai_mai_n675_), .Y(mai_mai_n678_));
  NO2        m656(.A(mai_mai_n431_), .B(mai_mai_n26_), .Y(mai_mai_n679_));
  INV        m657(.A(mai_mai_n678_), .Y(mai_mai_n680_));
  INV        m658(.A(mai_mai_n161_), .Y(mai_mai_n681_));
  NO3        m659(.A(mai_mai_n576_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n682_));
  AOI210     m660(.A0(mai_mai_n681_), .A1(mai_mai_n82_), .B0(mai_mai_n682_), .Y(mai_mai_n683_));
  NO2        m661(.A(mai_mai_n683_), .B(mai_mai_n182_), .Y(mai_mai_n684_));
  OA210      m662(.A0(mai_mai_n577_), .A1(mai_mai_n119_), .B0(i_13_), .Y(mai_mai_n685_));
  INV        m663(.A(mai_mai_n141_), .Y(mai_mai_n686_));
  NO2        m664(.A(mai_mai_n686_), .B(mai_mai_n349_), .Y(mai_mai_n687_));
  NO2        m665(.A(mai_mai_n138_), .B(mai_mai_n490_), .Y(mai_mai_n688_));
  NA2        m666(.A(mai_mai_n688_), .B(mai_mai_n396_), .Y(mai_mai_n689_));
  NO2        m667(.A(mai_mai_n95_), .B(mai_mai_n44_), .Y(mai_mai_n690_));
  INV        m668(.A(mai_mai_n284_), .Y(mai_mai_n691_));
  NA4        m669(.A(mai_mai_n691_), .B(mai_mai_n288_), .C(mai_mai_n117_), .D(mai_mai_n42_), .Y(mai_mai_n692_));
  OAI210     m670(.A0(mai_mai_n692_), .A1(mai_mai_n690_), .B0(mai_mai_n689_), .Y(mai_mai_n693_));
  NO4        m671(.A(mai_mai_n693_), .B(mai_mai_n687_), .C(mai_mai_n685_), .D(mai_mai_n684_), .Y(mai_mai_n694_));
  INV        m672(.A(mai_mai_n542_), .Y(mai_mai_n695_));
  NA2        m673(.A(mai_mai_n668_), .B(mai_mai_n258_), .Y(mai_mai_n696_));
  NA2        m674(.A(mai_mai_n696_), .B(mai_mai_n695_), .Y(mai_mai_n697_));
  NO2        m675(.A(mai_mai_n58_), .B(i_12_), .Y(mai_mai_n698_));
  AOI220     m676(.A0(mai_mai_n698_), .A1(mai_mai_n36_), .B0(mai_mai_n697_), .B1(mai_mai_n46_), .Y(mai_mai_n699_));
  NA4        m677(.A(mai_mai_n699_), .B(mai_mai_n694_), .C(mai_mai_n680_), .D(mai_mai_n674_), .Y(mai6));
  NO3        m678(.A(i_9_), .B(mai_mai_n290_), .C(i_1_), .Y(mai_mai_n701_));
  NO2        m679(.A(mai_mai_n174_), .B(mai_mai_n129_), .Y(mai_mai_n702_));
  OAI210     m680(.A0(mai_mai_n702_), .A1(mai_mai_n701_), .B0(mai_mai_n659_), .Y(mai_mai_n703_));
  NA4        m681(.A(mai_mai_n367_), .B(mai_mai_n459_), .C(mai_mai_n65_), .D(mai_mai_n94_), .Y(mai_mai_n704_));
  INV        m682(.A(mai_mai_n704_), .Y(mai_mai_n705_));
  NO2        m683(.A(i_11_), .B(i_9_), .Y(mai_mai_n706_));
  NO2        m684(.A(mai_mai_n705_), .B(mai_mai_n308_), .Y(mai_mai_n707_));
  AO210      m685(.A0(mai_mai_n707_), .A1(mai_mai_n703_), .B0(i_12_), .Y(mai_mai_n708_));
  NA2        m686(.A(mai_mai_n350_), .B(mai_mai_n315_), .Y(mai_mai_n709_));
  NA2        m687(.A(mai_mai_n549_), .B(mai_mai_n59_), .Y(mai_mai_n710_));
  NA2        m688(.A(mai_mai_n618_), .B(mai_mai_n65_), .Y(mai_mai_n711_));
  BUFFER     m689(.A(mai_mai_n80_), .Y(mai_mai_n712_));
  NA4        m690(.A(mai_mai_n712_), .B(mai_mai_n711_), .C(mai_mai_n710_), .D(mai_mai_n709_), .Y(mai_mai_n713_));
  INV        m691(.A(mai_mai_n185_), .Y(mai_mai_n714_));
  AOI220     m692(.A0(mai_mai_n714_), .A1(mai_mai_n706_), .B0(mai_mai_n713_), .B1(mai_mai_n67_), .Y(mai_mai_n715_));
  INV        m693(.A(mai_mai_n307_), .Y(mai_mai_n716_));
  INV        m694(.A(mai_mai_n117_), .Y(mai_mai_n717_));
  NA2        m695(.A(mai_mai_n717_), .B(mai_mai_n46_), .Y(mai_mai_n718_));
  NO2        m696(.A(mai_mai_n718_), .B(mai_mai_n716_), .Y(mai_mai_n719_));
  NO2        m697(.A(mai_mai_n239_), .B(i_9_), .Y(mai_mai_n720_));
  NA2        m698(.A(mai_mai_n720_), .B(mai_mai_n698_), .Y(mai_mai_n721_));
  NO2        m699(.A(mai_mai_n721_), .B(mai_mai_n174_), .Y(mai_mai_n722_));
  NO2        m700(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n723_));
  NA3        m701(.A(mai_mai_n723_), .B(mai_mai_n452_), .C(mai_mai_n367_), .Y(mai_mai_n724_));
  OAI210     m702(.A0(mai_mai_n618_), .A1(mai_mai_n531_), .B0(mai_mai_n530_), .Y(mai_mai_n725_));
  NA2        m703(.A(mai_mai_n725_), .B(mai_mai_n724_), .Y(mai_mai_n726_));
  OR3        m704(.A(mai_mai_n726_), .B(mai_mai_n722_), .C(mai_mai_n719_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n627_), .B(i_2_), .Y(mai_mai_n728_));
  NA2        m706(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n729_));
  OAI210     m707(.A0(mai_mai_n729_), .A1(mai_mai_n385_), .B0(mai_mai_n339_), .Y(mai_mai_n730_));
  NA2        m708(.A(mai_mai_n730_), .B(mai_mai_n728_), .Y(mai_mai_n731_));
  AO220      m709(.A0(mai_mai_n338_), .A1(mai_mai_n329_), .B0(mai_mai_n375_), .B1(i_8_), .Y(mai_mai_n732_));
  NA3        m710(.A(mai_mai_n732_), .B(mai_mai_n242_), .C(i_7_), .Y(mai_mai_n733_));
  BUFFER     m711(.A(mai_mai_n423_), .Y(mai_mai_n734_));
  NA3        m712(.A(mai_mai_n734_), .B(mai_mai_n137_), .C(mai_mai_n63_), .Y(mai_mai_n735_));
  AO210      m713(.A0(mai_mai_n468_), .A1(mai_mai_n671_), .B0(mai_mai_n36_), .Y(mai_mai_n736_));
  NA4        m714(.A(mai_mai_n736_), .B(mai_mai_n735_), .C(mai_mai_n733_), .D(mai_mai_n731_), .Y(mai_mai_n737_));
  OAI210     m715(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n80_), .Y(mai_mai_n738_));
  NA2        m716(.A(mai_mai_n738_), .B(mai_mai_n530_), .Y(mai_mai_n739_));
  OAI210     m717(.A0(mai_mai_n375_), .A1(mai_mai_n192_), .B0(mai_mai_n64_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n740_), .B(mai_mai_n739_), .Y(mai_mai_n741_));
  AO210      m719(.A0(mai_mai_n490_), .A1(mai_mai_n46_), .B0(mai_mai_n81_), .Y(mai_mai_n742_));
  NA3        m720(.A(mai_mai_n742_), .B(mai_mai_n460_), .C(mai_mai_n206_), .Y(mai_mai_n743_));
  AOI210     m721(.A0(mai_mai_n423_), .A1(mai_mai_n421_), .B0(mai_mai_n529_), .Y(mai_mai_n744_));
  NA2        m722(.A(mai_mai_n104_), .B(mai_mai_n383_), .Y(mai_mai_n745_));
  NA2        m723(.A(mai_mai_n231_), .B(mai_mai_n46_), .Y(mai_mai_n746_));
  NA3        m724(.A(mai_mai_n745_), .B(mai_mai_n744_), .C(mai_mai_n743_), .Y(mai_mai_n747_));
  NO4        m725(.A(mai_mai_n747_), .B(mai_mai_n741_), .C(mai_mai_n737_), .D(mai_mai_n727_), .Y(mai_mai_n748_));
  NA4        m726(.A(mai_mai_n748_), .B(mai_mai_n715_), .C(mai_mai_n708_), .D(mai_mai_n357_), .Y(mai3));
  NA2        m727(.A(i_6_), .B(i_7_), .Y(mai_mai_n750_));
  NO2        m728(.A(mai_mai_n750_), .B(i_0_), .Y(mai_mai_n751_));
  NO2        m729(.A(i_11_), .B(mai_mai_n224_), .Y(mai_mai_n752_));
  OAI210     m730(.A0(mai_mai_n751_), .A1(mai_mai_n272_), .B0(mai_mai_n752_), .Y(mai_mai_n753_));
  INV        m731(.A(mai_mai_n753_), .Y(mai_mai_n754_));
  NO3        m732(.A(mai_mai_n427_), .B(mai_mai_n84_), .C(mai_mai_n44_), .Y(mai_mai_n755_));
  OA210      m733(.A0(mai_mai_n755_), .A1(mai_mai_n754_), .B0(mai_mai_n163_), .Y(mai_mai_n756_));
  NA2        m734(.A(mai_mai_n386_), .B(mai_mai_n45_), .Y(mai_mai_n757_));
  NO4        m735(.A(mai_mai_n353_), .B(mai_mai_n360_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n758_));
  NA2        m736(.A(mai_mai_n174_), .B(mai_mai_n539_), .Y(mai_mai_n759_));
  NOi21      m737(.An(mai_mai_n759_), .B(mai_mai_n758_), .Y(mai_mai_n760_));
  NA2        m738(.A(mai_mai_n640_), .B(mai_mai_n611_), .Y(mai_mai_n761_));
  NA2        m739(.A(mai_mai_n313_), .B(i_5_), .Y(mai_mai_n762_));
  OAI220     m740(.A0(mai_mai_n762_), .A1(mai_mai_n761_), .B0(mai_mai_n760_), .B1(mai_mai_n59_), .Y(mai_mai_n763_));
  NOi21      m741(.An(i_5_), .B(i_9_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n764_), .B(mai_mai_n419_), .Y(mai_mai_n765_));
  NO2        m743(.A(mai_mai_n164_), .B(mai_mai_n138_), .Y(mai_mai_n766_));
  NA2        m744(.A(mai_mai_n766_), .B(mai_mai_n231_), .Y(mai_mai_n767_));
  NO2        m745(.A(mai_mai_n767_), .B(mai_mai_n170_), .Y(mai_mai_n768_));
  NO3        m746(.A(mai_mai_n768_), .B(mai_mai_n763_), .C(mai_mai_n756_), .Y(mai_mai_n769_));
  NA2        m747(.A(mai_mai_n174_), .B(mai_mai_n24_), .Y(mai_mai_n770_));
  NO2        m748(.A(mai_mai_n609_), .B(mai_mai_n556_), .Y(mai_mai_n771_));
  NO2        m749(.A(mai_mai_n771_), .B(mai_mai_n770_), .Y(mai_mai_n772_));
  NA2        m750(.A(mai_mai_n295_), .B(mai_mai_n122_), .Y(mai_mai_n773_));
  NAi21      m751(.An(mai_mai_n151_), .B(i_5_), .Y(mai_mai_n774_));
  OAI220     m752(.A0(mai_mai_n774_), .A1(mai_mai_n746_), .B0(mai_mai_n773_), .B1(mai_mai_n376_), .Y(mai_mai_n775_));
  NO2        m753(.A(mai_mai_n775_), .B(mai_mai_n772_), .Y(mai_mai_n776_));
  NO2        m754(.A(mai_mai_n367_), .B(mai_mai_n276_), .Y(mai_mai_n777_));
  NA2        m755(.A(mai_mai_n777_), .B(mai_mai_n643_), .Y(mai_mai_n778_));
  INV        m756(.A(mai_mai_n452_), .Y(mai_mai_n779_));
  AN2        m757(.A(mai_mai_n89_), .B(mai_mai_n230_), .Y(mai_mai_n780_));
  NA2        m758(.A(mai_mai_n668_), .B(mai_mai_n308_), .Y(mai_mai_n781_));
  NO2        m759(.A(mai_mai_n602_), .B(mai_mai_n508_), .Y(mai_mai_n782_));
  NO2        m760(.A(mai_mai_n241_), .B(mai_mai_n142_), .Y(mai_mai_n783_));
  NA2        m761(.A(i_0_), .B(i_10_), .Y(mai_mai_n784_));
  AN2        m762(.A(mai_mai_n783_), .B(i_6_), .Y(mai_mai_n785_));
  NA2        m763(.A(mai_mai_n174_), .B(mai_mai_n77_), .Y(mai_mai_n786_));
  NA2        m764(.A(mai_mai_n534_), .B(i_4_), .Y(mai_mai_n787_));
  NA2        m765(.A(mai_mai_n177_), .B(mai_mai_n191_), .Y(mai_mai_n788_));
  OAI220     m766(.A0(mai_mai_n788_), .A1(mai_mai_n781_), .B0(mai_mai_n787_), .B1(mai_mai_n786_), .Y(mai_mai_n789_));
  NO4        m767(.A(mai_mai_n789_), .B(mai_mai_n785_), .C(mai_mai_n782_), .D(mai_mai_n780_), .Y(mai_mai_n790_));
  NA3        m768(.A(mai_mai_n790_), .B(mai_mai_n778_), .C(mai_mai_n776_), .Y(mai_mai_n791_));
  NA2        m769(.A(i_11_), .B(i_9_), .Y(mai_mai_n792_));
  NO2        m770(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n793_));
  NA2        m771(.A(mai_mai_n372_), .B(mai_mai_n168_), .Y(mai_mai_n794_));
  NA2        m772(.A(mai_mai_n794_), .B(mai_mai_n149_), .Y(mai_mai_n795_));
  NO2        m773(.A(mai_mai_n792_), .B(mai_mai_n67_), .Y(mai_mai_n796_));
  NO2        m774(.A(mai_mai_n164_), .B(i_0_), .Y(mai_mai_n797_));
  NA2        m775(.A(mai_mai_n452_), .B(mai_mai_n218_), .Y(mai_mai_n798_));
  NA2        m776(.A(i_6_), .B(i_4_), .Y(mai_mai_n799_));
  OAI220     m777(.A0(mai_mai_n799_), .A1(mai_mai_n765_), .B0(mai_mai_n798_), .B1(mai_mai_n164_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n800_), .B(mai_mai_n795_), .Y(mai_mai_n801_));
  NA2        m779(.A(mai_mai_n601_), .B(mai_mai_n114_), .Y(mai_mai_n802_));
  NO2        m780(.A(i_6_), .B(mai_mai_n802_), .Y(mai_mai_n803_));
  AOI210     m781(.A0(mai_mai_n422_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n804_));
  NA2        m782(.A(mai_mai_n160_), .B(mai_mai_n96_), .Y(mai_mai_n805_));
  NOi32      m783(.An(mai_mai_n804_), .Bn(mai_mai_n177_), .C(mai_mai_n805_), .Y(mai_mai_n806_));
  NA2        m784(.A(mai_mai_n563_), .B(mai_mai_n308_), .Y(mai_mai_n807_));
  NO2        m785(.A(mai_mai_n807_), .B(mai_mai_n757_), .Y(mai_mai_n808_));
  NO3        m786(.A(mai_mai_n808_), .B(mai_mai_n806_), .C(mai_mai_n803_), .Y(mai_mai_n809_));
  NOi21      m787(.An(i_7_), .B(i_5_), .Y(mai_mai_n810_));
  NOi31      m788(.An(mai_mai_n810_), .B(i_0_), .C(mai_mai_n652_), .Y(mai_mai_n811_));
  NO3        m789(.A(mai_mai_n378_), .B(mai_mai_n341_), .C(mai_mai_n337_), .Y(mai_mai_n812_));
  NO2        m790(.A(mai_mai_n243_), .B(i_5_), .Y(mai_mai_n813_));
  INV        m791(.A(mai_mai_n652_), .Y(mai_mai_n814_));
  AOI210     m792(.A0(mai_mai_n814_), .A1(mai_mai_n813_), .B0(mai_mai_n812_), .Y(mai_mai_n815_));
  NA3        m793(.A(mai_mai_n815_), .B(mai_mai_n809_), .C(mai_mai_n801_), .Y(mai_mai_n816_));
  NO2        m794(.A(mai_mai_n770_), .B(mai_mai_n227_), .Y(mai_mai_n817_));
  AN2        m795(.A(mai_mai_n312_), .B(mai_mai_n308_), .Y(mai_mai_n818_));
  AN2        m796(.A(mai_mai_n818_), .B(mai_mai_n766_), .Y(mai_mai_n819_));
  OAI210     m797(.A0(mai_mai_n819_), .A1(mai_mai_n817_), .B0(i_10_), .Y(mai_mai_n820_));
  NA3        m798(.A(mai_mai_n451_), .B(mai_mai_n386_), .C(mai_mai_n45_), .Y(mai_mai_n821_));
  OAI210     m799(.A0(mai_mai_n774_), .A1(mai_mai_n779_), .B0(mai_mai_n821_), .Y(mai_mai_n822_));
  NO2        m800(.A(mai_mai_n242_), .B(mai_mai_n46_), .Y(mai_mai_n823_));
  NA2        m801(.A(mai_mai_n796_), .B(mai_mai_n288_), .Y(mai_mai_n824_));
  OAI210     m802(.A0(mai_mai_n823_), .A1(mai_mai_n176_), .B0(mai_mai_n824_), .Y(mai_mai_n825_));
  AOI220     m803(.A0(mai_mai_n825_), .A1(mai_mai_n452_), .B0(mai_mai_n822_), .B1(mai_mai_n67_), .Y(mai_mai_n826_));
  NA3        m804(.A(mai_mai_n729_), .B(mai_mai_n359_), .C(i_6_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n87_), .B(mai_mai_n44_), .Y(mai_mai_n828_));
  NO2        m806(.A(mai_mai_n69_), .B(mai_mai_n670_), .Y(mai_mai_n829_));
  AOI220     m807(.A0(mai_mai_n829_), .A1(mai_mai_n828_), .B0(mai_mai_n163_), .B1(mai_mai_n556_), .Y(mai_mai_n830_));
  AOI210     m808(.A0(mai_mai_n830_), .A1(mai_mai_n827_), .B0(mai_mai_n47_), .Y(mai_mai_n831_));
  NO3        m809(.A(mai_mai_n551_), .B(mai_mai_n336_), .C(mai_mai_n24_), .Y(mai_mai_n832_));
  AOI210     m810(.A0(mai_mai_n633_), .A1(mai_mai_n517_), .B0(mai_mai_n832_), .Y(mai_mai_n833_));
  NO2        m811(.A(mai_mai_n558_), .B(mai_mai_n98_), .Y(mai_mai_n834_));
  NA2        m812(.A(mai_mai_n834_), .B(i_0_), .Y(mai_mai_n835_));
  OAI220     m813(.A0(mai_mai_n835_), .A1(mai_mai_n79_), .B0(mai_mai_n833_), .B1(mai_mai_n161_), .Y(mai_mai_n836_));
  NO3        m814(.A(mai_mai_n836_), .B(mai_mai_n831_), .C(mai_mai_n492_), .Y(mai_mai_n837_));
  NA3        m815(.A(mai_mai_n837_), .B(mai_mai_n826_), .C(mai_mai_n820_), .Y(mai_mai_n838_));
  NO3        m816(.A(mai_mai_n838_), .B(mai_mai_n816_), .C(mai_mai_n791_), .Y(mai_mai_n839_));
  NO2        m817(.A(i_0_), .B(mai_mai_n652_), .Y(mai_mai_n840_));
  NO3        m818(.A(mai_mai_n98_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n841_));
  AO220      m819(.A0(mai_mai_n841_), .A1(mai_mai_n44_), .B0(mai_mai_n840_), .B1(mai_mai_n163_), .Y(mai_mai_n842_));
  NO2        m820(.A(mai_mai_n710_), .B(mai_mai_n805_), .Y(mai_mai_n843_));
  AOI210     m821(.A0(mai_mai_n842_), .A1(mai_mai_n327_), .B0(mai_mai_n843_), .Y(mai_mai_n844_));
  NA3        m822(.A(mai_mai_n136_), .B(mai_mai_n611_), .C(mai_mai_n67_), .Y(mai_mai_n845_));
  NO2        m823(.A(mai_mai_n725_), .B(mai_mai_n378_), .Y(mai_mai_n846_));
  NA3        m824(.A(mai_mai_n751_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n847_));
  NA2        m825(.A(mai_mai_n752_), .B(i_9_), .Y(mai_mai_n848_));
  AOI210     m826(.A0(mai_mai_n847_), .A1(mai_mai_n471_), .B0(mai_mai_n848_), .Y(mai_mai_n849_));
  NO2        m827(.A(mai_mai_n849_), .B(mai_mai_n846_), .Y(mai_mai_n850_));
  NA3        m828(.A(mai_mai_n850_), .B(mai_mai_n845_), .C(mai_mai_n844_), .Y(mai_mai_n851_));
  NA2        m829(.A(mai_mai_n818_), .B(mai_mai_n349_), .Y(mai_mai_n852_));
  AOI210     m830(.A0(mai_mai_n283_), .A1(mai_mai_n151_), .B0(mai_mai_n852_), .Y(mai_mai_n853_));
  NA2        m831(.A(mai_mai_n40_), .B(mai_mai_n44_), .Y(mai_mai_n854_));
  NA2        m832(.A(mai_mai_n793_), .B(mai_mai_n462_), .Y(mai_mai_n855_));
  AOI210     m833(.A0(mai_mai_n854_), .A1(mai_mai_n151_), .B0(mai_mai_n855_), .Y(mai_mai_n856_));
  NO2        m834(.A(mai_mai_n856_), .B(mai_mai_n853_), .Y(mai_mai_n857_));
  NO3        m835(.A(mai_mai_n784_), .B(mai_mai_n764_), .C(mai_mai_n179_), .Y(mai_mai_n858_));
  AOI220     m836(.A0(mai_mai_n858_), .A1(i_11_), .B0(mai_mai_n535_), .B1(mai_mai_n69_), .Y(mai_mai_n859_));
  NO3        m837(.A(mai_mai_n198_), .B(mai_mai_n360_), .C(i_0_), .Y(mai_mai_n860_));
  OAI210     m838(.A0(mai_mai_n860_), .A1(mai_mai_n70_), .B0(i_13_), .Y(mai_mai_n861_));
  INV        m839(.A(mai_mai_n206_), .Y(mai_mai_n862_));
  OAI220     m840(.A0(mai_mai_n502_), .A1(mai_mai_n129_), .B0(mai_mai_n947_), .B1(mai_mai_n571_), .Y(mai_mai_n863_));
  NA2        m841(.A(mai_mai_n863_), .B(mai_mai_n862_), .Y(mai_mai_n864_));
  NA4        m842(.A(mai_mai_n864_), .B(mai_mai_n861_), .C(mai_mai_n859_), .D(mai_mai_n857_), .Y(mai_mai_n865_));
  NA2        m843(.A(mai_mai_n810_), .B(mai_mai_n462_), .Y(mai_mai_n866_));
  INV        m844(.A(mai_mai_n165_), .Y(mai_mai_n867_));
  OR2        m845(.A(mai_mai_n867_), .B(mai_mai_n866_), .Y(mai_mai_n868_));
  AOI210     m846(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n164_), .Y(mai_mai_n869_));
  NA3        m847(.A(mai_mai_n568_), .B(mai_mai_n174_), .C(mai_mai_n77_), .Y(mai_mai_n870_));
  NA2        m848(.A(mai_mai_n870_), .B(mai_mai_n515_), .Y(mai_mai_n871_));
  NO3        m849(.A(mai_mai_n757_), .B(mai_mai_n54_), .C(mai_mai_n48_), .Y(mai_mai_n872_));
  NA2        m850(.A(mai_mai_n467_), .B(mai_mai_n449_), .Y(mai_mai_n873_));
  NO3        m851(.A(mai_mai_n873_), .B(mai_mai_n872_), .C(mai_mai_n871_), .Y(mai_mai_n874_));
  NA3        m852(.A(mai_mai_n793_), .B(mai_mai_n272_), .C(mai_mai_n217_), .Y(mai_mai_n875_));
  INV        m853(.A(mai_mai_n875_), .Y(mai_mai_n876_));
  NA3        m854(.A(mai_mai_n367_), .B(mai_mai_n314_), .C(mai_mai_n209_), .Y(mai_mai_n877_));
  INV        m855(.A(mai_mai_n877_), .Y(mai_mai_n878_));
  NO3        m856(.A(mai_mai_n792_), .B(mai_mai_n206_), .C(mai_mai_n179_), .Y(mai_mai_n879_));
  NO3        m857(.A(mai_mai_n879_), .B(mai_mai_n878_), .C(mai_mai_n876_), .Y(mai_mai_n880_));
  NA3        m858(.A(mai_mai_n880_), .B(mai_mai_n874_), .C(mai_mai_n868_), .Y(mai_mai_n881_));
  INV        m859(.A(mai_mai_n570_), .Y(mai_mai_n882_));
  NO3        m860(.A(mai_mai_n882_), .B(mai_mai_n948_), .C(i_3_), .Y(mai_mai_n883_));
  INV        m861(.A(mai_mai_n883_), .Y(mai_mai_n884_));
  NA3        m862(.A(mai_mai_n288_), .B(i_5_), .C(mai_mai_n182_), .Y(mai_mai_n885_));
  NA2        m863(.A(mai_mai_n885_), .B(mai_mai_n229_), .Y(mai_mai_n886_));
  NO4        m864(.A(mai_mai_n227_), .B(mai_mai_n198_), .C(i_0_), .D(i_12_), .Y(mai_mai_n887_));
  AOI220     m865(.A0(mai_mai_n887_), .A1(mai_mai_n886_), .B0(mai_mai_n705_), .B1(mai_mai_n165_), .Y(mai_mai_n888_));
  AN2        m866(.A(mai_mai_n784_), .B(mai_mai_n142_), .Y(mai_mai_n889_));
  NO3        m867(.A(mai_mai_n889_), .B(i_12_), .C(mai_mai_n595_), .Y(mai_mai_n890_));
  NA2        m868(.A(mai_mai_n890_), .B(mai_mai_n206_), .Y(mai_mai_n891_));
  NA3        m869(.A(mai_mai_n91_), .B(mai_mai_n539_), .C(i_11_), .Y(mai_mai_n892_));
  NO2        m870(.A(mai_mai_n892_), .B(mai_mai_n144_), .Y(mai_mai_n893_));
  NA2        m871(.A(mai_mai_n810_), .B(mai_mai_n448_), .Y(mai_mai_n894_));
  NA2        m872(.A(mai_mai_n60_), .B(mai_mai_n94_), .Y(mai_mai_n895_));
  OAI220     m873(.A0(mai_mai_n895_), .A1(mai_mai_n885_), .B0(mai_mai_n894_), .B1(mai_mai_n612_), .Y(mai_mai_n896_));
  AOI210     m874(.A0(mai_mai_n896_), .A1(mai_mai_n797_), .B0(mai_mai_n893_), .Y(mai_mai_n897_));
  NA4        m875(.A(mai_mai_n897_), .B(mai_mai_n891_), .C(mai_mai_n888_), .D(mai_mai_n884_), .Y(mai_mai_n898_));
  NO4        m876(.A(mai_mai_n898_), .B(mai_mai_n881_), .C(mai_mai_n865_), .D(mai_mai_n851_), .Y(mai_mai_n899_));
  OAI210     m877(.A0(mai_mai_n728_), .A1(mai_mai_n723_), .B0(mai_mai_n37_), .Y(mai_mai_n900_));
  NA3        m878(.A(mai_mai_n804_), .B(mai_mai_n345_), .C(i_5_), .Y(mai_mai_n901_));
  NA3        m879(.A(mai_mai_n901_), .B(mai_mai_n900_), .C(mai_mai_n567_), .Y(mai_mai_n902_));
  NA2        m880(.A(mai_mai_n902_), .B(mai_mai_n195_), .Y(mai_mai_n903_));
  NA2        m881(.A(mai_mai_n175_), .B(mai_mai_n177_), .Y(mai_mai_n904_));
  AO210      m882(.A0(i_11_), .A1(mai_mai_n33_), .B0(mai_mai_n904_), .Y(mai_mai_n905_));
  NAi31      m883(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n906_));
  NO2        m884(.A(mai_mai_n64_), .B(mai_mai_n906_), .Y(mai_mai_n907_));
  NO2        m885(.A(mai_mai_n907_), .B(mai_mai_n593_), .Y(mai_mai_n908_));
  NA2        m886(.A(mai_mai_n908_), .B(mai_mai_n905_), .Y(mai_mai_n909_));
  NO2        m887(.A(mai_mai_n439_), .B(mai_mai_n249_), .Y(mai_mai_n910_));
  NO4        m888(.A(mai_mai_n220_), .B(mai_mai_n135_), .C(mai_mai_n615_), .D(mai_mai_n37_), .Y(mai_mai_n911_));
  NO2        m889(.A(mai_mai_n911_), .B(mai_mai_n910_), .Y(mai_mai_n912_));
  OAI210     m890(.A0(mai_mai_n892_), .A1(mai_mai_n138_), .B0(mai_mai_n912_), .Y(mai_mai_n913_));
  AOI210     m891(.A0(mai_mai_n909_), .A1(mai_mai_n48_), .B0(mai_mai_n913_), .Y(mai_mai_n914_));
  AOI210     m892(.A0(mai_mai_n914_), .A1(mai_mai_n903_), .B0(mai_mai_n67_), .Y(mai_mai_n915_));
  NO2        m893(.A(mai_mai_n532_), .B(mai_mai_n356_), .Y(mai_mai_n916_));
  NO2        m894(.A(mai_mai_n916_), .B(mai_mai_n675_), .Y(mai_mai_n917_));
  INV        m895(.A(mai_mai_n101_), .Y(mai_mai_n918_));
  NA2        m896(.A(mai_mai_n918_), .B(mai_mai_n70_), .Y(mai_mai_n919_));
  AOI210     m897(.A0(mai_mai_n869_), .A1(mai_mai_n793_), .B0(mai_mai_n811_), .Y(mai_mai_n920_));
  AOI210     m898(.A0(mai_mai_n920_), .A1(mai_mai_n919_), .B0(mai_mai_n615_), .Y(mai_mai_n921_));
  INV        m899(.A(mai_mai_n243_), .Y(mai_mai_n922_));
  NA2        m900(.A(mai_mai_n922_), .B(mai_mai_n70_), .Y(mai_mai_n923_));
  NO2        m901(.A(mai_mai_n923_), .B(mai_mai_n224_), .Y(mai_mai_n924_));
  NA3        m902(.A(mai_mai_n89_), .B(mai_mai_n290_), .C(mai_mai_n31_), .Y(mai_mai_n925_));
  INV        m903(.A(mai_mai_n925_), .Y(mai_mai_n926_));
  NO3        m904(.A(mai_mai_n926_), .B(mai_mai_n924_), .C(mai_mai_n921_), .Y(mai_mai_n927_));
  OAI210     m905(.A0(mai_mai_n251_), .A1(mai_mai_n147_), .B0(mai_mai_n82_), .Y(mai_mai_n928_));
  NA2        m906(.A(mai_mai_n679_), .B(mai_mai_n272_), .Y(mai_mai_n929_));
  AOI210     m907(.A0(mai_mai_n929_), .A1(mai_mai_n928_), .B0(i_11_), .Y(mai_mai_n930_));
  INV        m908(.A(mai_mai_n195_), .Y(mai_mai_n931_));
  NA2        m909(.A(mai_mai_n153_), .B(i_5_), .Y(mai_mai_n932_));
  NO2        m910(.A(mai_mai_n931_), .B(mai_mai_n932_), .Y(mai_mai_n933_));
  NO3        m911(.A(i_9_), .B(mai_mai_n453_), .C(mai_mai_n240_), .Y(mai_mai_n934_));
  NO2        m912(.A(mai_mai_n934_), .B(mai_mai_n529_), .Y(mai_mai_n935_));
  INV        m913(.A(mai_mai_n342_), .Y(mai_mai_n936_));
  AOI210     m914(.A0(mai_mai_n936_), .A1(mai_mai_n935_), .B0(mai_mai_n41_), .Y(mai_mai_n937_));
  NO3        m915(.A(mai_mai_n937_), .B(mai_mai_n933_), .C(mai_mai_n930_), .Y(mai_mai_n938_));
  OAI210     m916(.A0(mai_mai_n927_), .A1(i_4_), .B0(mai_mai_n938_), .Y(mai_mai_n939_));
  NO3        m917(.A(mai_mai_n939_), .B(mai_mai_n917_), .C(mai_mai_n915_), .Y(mai_mai_n940_));
  NA4        m918(.A(mai_mai_n940_), .B(mai_mai_n899_), .C(mai_mai_n839_), .D(mai_mai_n769_), .Y(mai4));
  INV        m919(.A(i_2_), .Y(mai_mai_n944_));
  INV        m920(.A(i_3_), .Y(mai_mai_n945_));
  INV        m921(.A(i_7_), .Y(mai_mai_n946_));
  INV        m922(.A(i_6_), .Y(mai_mai_n947_));
  INV        m923(.A(i_0_), .Y(mai_mai_n948_));
  INV        m924(.A(i_10_), .Y(mai_mai_n949_));
  INV        m925(.A(i_4_), .Y(mai_mai_n950_));
  INV        m926(.A(i_1_), .Y(mai_mai_n951_));
  NAi21      u000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u002(.A(i_9_), .Y(men_men_n25_));
  INV        u003(.A(i_3_), .Y(men_men_n26_));
  NO2        u004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u013(.A(i_4_), .Y(men_men_n36_));
  INV        u014(.A(i_10_), .Y(men_men_n37_));
  BUFFER     u015(.A(i_11_), .Y(men_men_n38_));
  NOi21      u016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u017(.A(men_men_n39_), .Y(men_men_n40_));
  NO2        u018(.A(men_men_n36_), .B(i_3_), .Y(men_men_n41_));
  NAi31      u019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u020(.A(men_men_n35_), .Y(men1));
  INV        u021(.A(i_11_), .Y(men_men_n44_));
  NO2        u022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u023(.A(i_2_), .Y(men_men_n46_));
  NA2        u024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u025(.A(i_5_), .Y(men_men_n48_));
  NO2        u026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  NA2        u028(.A(i_0_), .B(i_2_), .Y(men_men_n51_));
  NA2        u029(.A(i_7_), .B(i_9_), .Y(men_men_n52_));
  NO2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NA3        u031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n54_));
  NO2        u032(.A(i_1_), .B(i_6_), .Y(men_men_n55_));
  NA2        u033(.A(i_8_), .B(i_7_), .Y(men_men_n56_));
  OAI210     u034(.A0(men_men_n56_), .A1(men_men_n55_), .B0(men_men_n54_), .Y(men_men_n57_));
  NA2        u035(.A(men_men_n57_), .B(i_12_), .Y(men_men_n58_));
  NAi21      u036(.An(i_2_), .B(i_7_), .Y(men_men_n59_));
  INV        u037(.A(i_1_), .Y(men_men_n60_));
  NA2        u038(.A(men_men_n60_), .B(i_6_), .Y(men_men_n61_));
  NA3        u039(.A(men_men_n61_), .B(men_men_n59_), .C(men_men_n31_), .Y(men_men_n62_));
  NA2        u040(.A(men_men_n62_), .B(men_men_n58_), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n50_), .B(i_2_), .Y(men_men_n64_));
  AOI210     u042(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n65_));
  NA2        u043(.A(i_1_), .B(i_6_), .Y(men_men_n66_));
  NO2        u044(.A(men_men_n66_), .B(men_men_n25_), .Y(men_men_n67_));
  INV        u045(.A(i_0_), .Y(men_men_n68_));
  NAi21      u046(.An(i_5_), .B(i_10_), .Y(men_men_n69_));
  NA2        u047(.A(i_5_), .B(i_9_), .Y(men_men_n70_));
  AOI210     u048(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n68_), .Y(men_men_n71_));
  NO2        u049(.A(men_men_n71_), .B(men_men_n67_), .Y(men_men_n72_));
  OAI210     u050(.A0(men_men_n65_), .A1(men_men_n64_), .B0(men_men_n72_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n73_), .A1(men_men_n63_), .B0(i_0_), .Y(men_men_n74_));
  NA2        u052(.A(i_12_), .B(i_5_), .Y(men_men_n75_));
  NA2        u053(.A(i_2_), .B(i_8_), .Y(men_men_n76_));
  NO2        u054(.A(i_3_), .B(i_9_), .Y(men_men_n77_));
  NO2        u055(.A(i_3_), .B(i_7_), .Y(men_men_n78_));
  INV        u056(.A(i_6_), .Y(men_men_n79_));
  OR4        u057(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n80_));
  INV        u058(.A(men_men_n80_), .Y(men_men_n81_));
  NO2        u059(.A(i_2_), .B(i_7_), .Y(men_men_n82_));
  NAi21      u060(.An(i_6_), .B(i_10_), .Y(men_men_n83_));
  NA2        u061(.A(i_6_), .B(i_9_), .Y(men_men_n84_));
  AOI210     u062(.A0(men_men_n84_), .A1(men_men_n83_), .B0(men_men_n60_), .Y(men_men_n85_));
  NA2        u063(.A(i_2_), .B(i_6_), .Y(men_men_n86_));
  NO3        u064(.A(men_men_n86_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n87_));
  NO2        u065(.A(men_men_n87_), .B(men_men_n85_), .Y(men_men_n88_));
  AOI210     u066(.A0(men_men_n88_), .A1(men_men_n76_), .B0(men_men_n75_), .Y(men_men_n89_));
  AN3        u067(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n90_));
  NAi21      u068(.An(i_6_), .B(i_11_), .Y(men_men_n91_));
  NO2        u069(.A(i_5_), .B(i_8_), .Y(men_men_n92_));
  NOi21      u070(.An(men_men_n92_), .B(men_men_n91_), .Y(men_men_n93_));
  AOI220     u071(.A0(men_men_n93_), .A1(men_men_n59_), .B0(men_men_n90_), .B1(men_men_n32_), .Y(men_men_n94_));
  INV        u072(.A(i_7_), .Y(men_men_n95_));
  NA2        u073(.A(men_men_n46_), .B(men_men_n95_), .Y(men_men_n96_));
  NO2        u074(.A(i_0_), .B(i_5_), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n97_), .B(men_men_n79_), .Y(men_men_n98_));
  NA2        u076(.A(i_12_), .B(i_3_), .Y(men_men_n99_));
  INV        u077(.A(men_men_n99_), .Y(men_men_n100_));
  NA3        u078(.A(men_men_n100_), .B(men_men_n98_), .C(men_men_n96_), .Y(men_men_n101_));
  NAi21      u079(.An(i_7_), .B(i_11_), .Y(men_men_n102_));
  NO3        u080(.A(men_men_n102_), .B(men_men_n83_), .C(men_men_n51_), .Y(men_men_n103_));
  AN2        u081(.A(i_2_), .B(i_10_), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(i_7_), .Y(men_men_n105_));
  OR2        u083(.A(men_men_n75_), .B(men_men_n55_), .Y(men_men_n106_));
  NO2        u084(.A(i_8_), .B(men_men_n95_), .Y(men_men_n107_));
  NO3        u085(.A(men_men_n107_), .B(men_men_n106_), .C(men_men_n105_), .Y(men_men_n108_));
  NA2        u086(.A(i_12_), .B(i_7_), .Y(men_men_n109_));
  NA2        u087(.A(i_3_), .B(i_0_), .Y(men_men_n110_));
  NA2        u088(.A(i_11_), .B(i_12_), .Y(men_men_n111_));
  OAI210     u089(.A0(men_men_n110_), .A1(men_men_n109_), .B0(men_men_n111_), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n112_), .B(men_men_n108_), .Y(men_men_n113_));
  NAi41      u091(.An(men_men_n103_), .B(men_men_n113_), .C(men_men_n101_), .D(men_men_n94_), .Y(men_men_n114_));
  NOi21      u092(.An(i_1_), .B(i_5_), .Y(men_men_n115_));
  NA2        u093(.A(men_men_n115_), .B(i_11_), .Y(men_men_n116_));
  NA2        u094(.A(men_men_n95_), .B(men_men_n37_), .Y(men_men_n117_));
  NA2        u095(.A(i_7_), .B(men_men_n25_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n118_), .B(men_men_n117_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(men_men_n46_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n84_), .B(men_men_n83_), .Y(men_men_n121_));
  NAi21      u099(.An(i_3_), .B(i_8_), .Y(men_men_n122_));
  NA2        u100(.A(men_men_n122_), .B(men_men_n59_), .Y(men_men_n123_));
  NOi31      u101(.An(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .Y(men_men_n124_));
  NO2        u102(.A(i_1_), .B(men_men_n79_), .Y(men_men_n125_));
  NO2        u103(.A(i_6_), .B(i_5_), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n126_), .B(i_3_), .Y(men_men_n127_));
  AO210      u105(.A0(men_men_n127_), .A1(men_men_n47_), .B0(men_men_n125_), .Y(men_men_n128_));
  OAI220     u106(.A0(men_men_n128_), .A1(men_men_n102_), .B0(men_men_n124_), .B1(men_men_n116_), .Y(men_men_n129_));
  NO3        u107(.A(men_men_n129_), .B(men_men_n114_), .C(men_men_n89_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n130_), .B(men_men_n74_), .Y(men2));
  NO2        u109(.A(men_men_n60_), .B(men_men_n37_), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n982_), .B(men_men_n132_), .Y(men_men_n133_));
  NA4        u111(.A(men_men_n133_), .B(men_men_n72_), .C(men_men_n64_), .D(men_men_n30_), .Y(men0));
  AN2        u112(.A(i_8_), .B(i_7_), .Y(men_men_n135_));
  NA2        u113(.A(men_men_n135_), .B(i_6_), .Y(men_men_n136_));
  NO2        u114(.A(i_12_), .B(i_13_), .Y(men_men_n137_));
  NAi21      u115(.An(i_5_), .B(i_11_), .Y(men_men_n138_));
  NOi21      u116(.An(men_men_n137_), .B(men_men_n138_), .Y(men_men_n139_));
  NO2        u117(.A(i_0_), .B(i_1_), .Y(men_men_n140_));
  NA2        u118(.A(i_2_), .B(i_3_), .Y(men_men_n141_));
  NO2        u119(.A(men_men_n141_), .B(i_4_), .Y(men_men_n142_));
  NA3        u120(.A(men_men_n142_), .B(men_men_n140_), .C(men_men_n139_), .Y(men_men_n143_));
  OR2        u121(.A(men_men_n143_), .B(men_men_n25_), .Y(men_men_n144_));
  AN2        u122(.A(men_men_n137_), .B(men_men_n77_), .Y(men_men_n145_));
  NO2        u123(.A(men_men_n145_), .B(men_men_n27_), .Y(men_men_n146_));
  NA2        u124(.A(i_1_), .B(i_5_), .Y(men_men_n147_));
  NO2        u125(.A(men_men_n68_), .B(men_men_n46_), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n148_), .B(men_men_n36_), .Y(men_men_n149_));
  NO3        u127(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n150_));
  OR2        u128(.A(i_0_), .B(i_1_), .Y(men_men_n151_));
  NO3        u129(.A(men_men_n151_), .B(men_men_n75_), .C(i_13_), .Y(men_men_n152_));
  NAi32      u130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n153_));
  NAi21      u131(.An(men_men_n153_), .B(men_men_n152_), .Y(men_men_n154_));
  NOi21      u132(.An(i_4_), .B(i_10_), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n155_), .B(men_men_n39_), .Y(men_men_n156_));
  NO2        u134(.A(i_3_), .B(i_5_), .Y(men_men_n157_));
  NO3        u135(.A(men_men_n68_), .B(i_2_), .C(i_1_), .Y(men_men_n158_));
  OAI210     u136(.A0(i_2_), .A1(men_men_n156_), .B0(men_men_n154_), .Y(men_men_n159_));
  NO2        u137(.A(men_men_n159_), .B(men_men_n150_), .Y(men_men_n160_));
  AOI210     u138(.A0(men_men_n160_), .A1(men_men_n144_), .B0(men_men_n136_), .Y(men_men_n161_));
  NA3        u139(.A(men_men_n68_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n162_));
  NOi21      u140(.An(i_4_), .B(i_9_), .Y(men_men_n163_));
  NOi21      u141(.An(i_11_), .B(i_13_), .Y(men_men_n164_));
  NA2        u142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  NO2        u143(.A(i_4_), .B(i_5_), .Y(men_men_n166_));
  NAi21      u144(.An(i_12_), .B(i_11_), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n167_), .B(i_13_), .Y(men_men_n168_));
  NA2        u146(.A(men_men_n168_), .B(men_men_n166_), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n169_), .A1(men_men_n165_), .B0(men_men_n162_), .Y(men_men_n170_));
  NO2        u148(.A(men_men_n68_), .B(men_men_n60_), .Y(men_men_n171_));
  NA2        u149(.A(men_men_n36_), .B(i_5_), .Y(men_men_n172_));
  NAi31      u150(.An(men_men_n172_), .B(men_men_n145_), .C(i_11_), .Y(men_men_n173_));
  NA2        u151(.A(i_3_), .B(i_5_), .Y(men_men_n174_));
  OR2        u152(.A(men_men_n174_), .B(men_men_n165_), .Y(men_men_n175_));
  AOI210     u153(.A0(men_men_n175_), .A1(men_men_n173_), .B0(i_2_), .Y(men_men_n176_));
  NO2        u154(.A(men_men_n68_), .B(i_5_), .Y(men_men_n177_));
  NO2        u155(.A(i_13_), .B(i_10_), .Y(men_men_n178_));
  NA3        u156(.A(men_men_n178_), .B(men_men_n177_), .C(men_men_n44_), .Y(men_men_n179_));
  NO2        u157(.A(i_2_), .B(i_1_), .Y(men_men_n180_));
  NA2        u158(.A(men_men_n180_), .B(i_3_), .Y(men_men_n181_));
  NAi21      u159(.An(i_4_), .B(i_12_), .Y(men_men_n182_));
  NO3        u160(.A(men_men_n182_), .B(men_men_n181_), .C(men_men_n25_), .Y(men_men_n183_));
  NO3        u161(.A(men_men_n183_), .B(men_men_n176_), .C(men_men_n170_), .Y(men_men_n184_));
  INV        u162(.A(i_8_), .Y(men_men_n185_));
  NO2        u163(.A(men_men_n185_), .B(i_7_), .Y(men_men_n186_));
  NA2        u164(.A(men_men_n186_), .B(i_6_), .Y(men_men_n187_));
  NO3        u165(.A(i_3_), .B(men_men_n79_), .C(men_men_n48_), .Y(men_men_n188_));
  NA2        u166(.A(men_men_n188_), .B(men_men_n107_), .Y(men_men_n189_));
  NO3        u167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n190_));
  NA3        u168(.A(men_men_n190_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n191_));
  NO3        u169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n192_));
  OAI210     u170(.A0(men_men_n90_), .A1(i_12_), .B0(men_men_n192_), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n193_), .A1(men_men_n191_), .B0(men_men_n189_), .Y(men_men_n194_));
  NO2        u172(.A(i_3_), .B(i_8_), .Y(men_men_n195_));
  NO3        u173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n196_));
  NA3        u174(.A(men_men_n196_), .B(men_men_n195_), .C(men_men_n39_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n97_), .B(men_men_n55_), .Y(men_men_n198_));
  INV        u176(.A(men_men_n198_), .Y(men_men_n199_));
  NO2        u177(.A(i_13_), .B(i_9_), .Y(men_men_n200_));
  NAi21      u178(.An(i_12_), .B(i_3_), .Y(men_men_n201_));
  NO2        u179(.A(men_men_n44_), .B(i_5_), .Y(men_men_n202_));
  NO3        u180(.A(i_0_), .B(i_2_), .C(men_men_n60_), .Y(men_men_n203_));
  NA2        u181(.A(men_men_n203_), .B(i_10_), .Y(men_men_n204_));
  OAI220     u182(.A0(men_men_n204_), .A1(men_men_n201_), .B0(men_men_n199_), .B1(men_men_n197_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n205_), .A1(i_7_), .B0(men_men_n194_), .Y(men_men_n206_));
  OAI220     u184(.A0(men_men_n206_), .A1(i_4_), .B0(men_men_n187_), .B1(men_men_n184_), .Y(men_men_n207_));
  NAi21      u185(.An(i_12_), .B(i_7_), .Y(men_men_n208_));
  NA3        u186(.A(i_13_), .B(men_men_n185_), .C(i_10_), .Y(men_men_n209_));
  NO2        u187(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  NA2        u188(.A(i_0_), .B(i_5_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n211_), .B(men_men_n98_), .Y(men_men_n212_));
  OAI220     u190(.A0(men_men_n212_), .A1(men_men_n181_), .B0(i_2_), .B1(men_men_n127_), .Y(men_men_n213_));
  NAi31      u191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n36_), .B(i_13_), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n68_), .B(men_men_n26_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n46_), .B(men_men_n60_), .Y(men_men_n217_));
  NA3        u195(.A(men_men_n217_), .B(men_men_n216_), .C(men_men_n215_), .Y(men_men_n218_));
  INV        u196(.A(i_13_), .Y(men_men_n219_));
  NO2        u197(.A(i_12_), .B(men_men_n219_), .Y(men_men_n220_));
  NA3        u198(.A(men_men_n220_), .B(men_men_n190_), .C(men_men_n188_), .Y(men_men_n221_));
  OAI210     u199(.A0(men_men_n218_), .A1(men_men_n214_), .B0(men_men_n221_), .Y(men_men_n222_));
  AOI220     u200(.A0(men_men_n222_), .A1(men_men_n135_), .B0(men_men_n213_), .B1(men_men_n210_), .Y(men_men_n223_));
  NO2        u201(.A(i_12_), .B(men_men_n37_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n174_), .B(i_4_), .Y(men_men_n225_));
  NA2        u203(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  OR2        u204(.A(i_8_), .B(i_7_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n227_), .B(men_men_n79_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n51_), .B(i_1_), .Y(men_men_n229_));
  NA2        u207(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  INV        u208(.A(i_12_), .Y(men_men_n231_));
  NO3        u209(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n232_));
  NA2        u210(.A(i_2_), .B(i_1_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n230_), .B(men_men_n226_), .Y(men_men_n234_));
  NO3        u212(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n235_));
  NAi21      u213(.An(i_4_), .B(i_3_), .Y(men_men_n236_));
  NO2        u214(.A(i_0_), .B(i_6_), .Y(men_men_n237_));
  NOi41      u215(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n238_));
  NA2        u216(.A(men_men_n238_), .B(men_men_n237_), .Y(men_men_n239_));
  NO2        u217(.A(men_men_n233_), .B(men_men_n174_), .Y(men_men_n240_));
  NAi21      u218(.An(men_men_n239_), .B(men_men_n240_), .Y(men_men_n241_));
  INV        u219(.A(men_men_n241_), .Y(men_men_n242_));
  AOI220     u220(.A0(men_men_n242_), .A1(men_men_n39_), .B0(men_men_n234_), .B1(men_men_n200_), .Y(men_men_n243_));
  NO2        u221(.A(i_11_), .B(men_men_n219_), .Y(men_men_n244_));
  NOi21      u222(.An(i_1_), .B(i_6_), .Y(men_men_n245_));
  NAi21      u223(.An(i_3_), .B(i_7_), .Y(men_men_n246_));
  OR4        u224(.A(i_12_), .B(men_men_n246_), .C(men_men_n245_), .D(men_men_n177_), .Y(men_men_n247_));
  NO2        u225(.A(i_12_), .B(i_3_), .Y(men_men_n248_));
  NA2        u226(.A(men_men_n68_), .B(i_5_), .Y(men_men_n249_));
  NA2        u227(.A(i_3_), .B(i_9_), .Y(men_men_n250_));
  NAi21      u228(.An(i_7_), .B(i_10_), .Y(men_men_n251_));
  NO2        u229(.A(men_men_n251_), .B(men_men_n250_), .Y(men_men_n252_));
  NA2        u230(.A(men_men_n252_), .B(men_men_n249_), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n253_), .B(men_men_n247_), .Y(men_men_n254_));
  INV        u232(.A(men_men_n136_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n231_), .B(i_13_), .Y(men_men_n256_));
  NO2        u234(.A(men_men_n256_), .B(men_men_n70_), .Y(men_men_n257_));
  AOI220     u235(.A0(men_men_n257_), .A1(men_men_n255_), .B0(men_men_n254_), .B1(men_men_n244_), .Y(men_men_n258_));
  NO2        u236(.A(men_men_n227_), .B(men_men_n37_), .Y(men_men_n259_));
  NA2        u237(.A(i_12_), .B(i_6_), .Y(men_men_n260_));
  OR2        u238(.A(i_13_), .B(i_9_), .Y(men_men_n261_));
  NO3        u239(.A(men_men_n261_), .B(men_men_n260_), .C(men_men_n48_), .Y(men_men_n262_));
  NO2        u240(.A(men_men_n236_), .B(i_2_), .Y(men_men_n263_));
  NA3        u241(.A(men_men_n263_), .B(men_men_n262_), .C(men_men_n44_), .Y(men_men_n264_));
  NA2        u242(.A(men_men_n244_), .B(i_9_), .Y(men_men_n265_));
  OAI210     u243(.A0(men_men_n68_), .A1(men_men_n265_), .B0(men_men_n264_), .Y(men_men_n266_));
  NO3        u244(.A(i_11_), .B(men_men_n219_), .C(men_men_n25_), .Y(men_men_n267_));
  NO2        u245(.A(men_men_n246_), .B(i_8_), .Y(men_men_n268_));
  NO2        u246(.A(i_6_), .B(men_men_n48_), .Y(men_men_n269_));
  NA3        u247(.A(men_men_n269_), .B(men_men_n268_), .C(men_men_n267_), .Y(men_men_n270_));
  NO3        u248(.A(men_men_n26_), .B(men_men_n79_), .C(i_5_), .Y(men_men_n271_));
  NA3        u249(.A(men_men_n271_), .B(men_men_n259_), .C(men_men_n220_), .Y(men_men_n272_));
  AOI210     u250(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n46_), .Y(men_men_n273_));
  AOI210     u251(.A0(men_men_n266_), .A1(men_men_n259_), .B0(men_men_n273_), .Y(men_men_n274_));
  NA4        u252(.A(men_men_n274_), .B(men_men_n258_), .C(men_men_n243_), .D(men_men_n223_), .Y(men_men_n275_));
  NO3        u253(.A(i_12_), .B(men_men_n219_), .C(men_men_n37_), .Y(men_men_n276_));
  INV        u254(.A(men_men_n276_), .Y(men_men_n277_));
  NOi21      u255(.An(men_men_n157_), .B(men_men_n79_), .Y(men_men_n278_));
  NO3        u256(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n279_));
  AOI220     u257(.A0(men_men_n279_), .A1(men_men_n188_), .B0(men_men_n278_), .B1(men_men_n229_), .Y(men_men_n280_));
  NO2        u258(.A(men_men_n280_), .B(i_7_), .Y(men_men_n281_));
  NO2        u259(.A(men_men_n233_), .B(i_0_), .Y(men_men_n282_));
  AOI220     u260(.A0(men_men_n282_), .A1(men_men_n186_), .B0(i_1_), .B1(men_men_n135_), .Y(men_men_n283_));
  NA2        u261(.A(men_men_n269_), .B(men_men_n26_), .Y(men_men_n284_));
  NO2        u262(.A(men_men_n284_), .B(men_men_n283_), .Y(men_men_n285_));
  NA2        u263(.A(i_0_), .B(i_1_), .Y(men_men_n286_));
  NO2        u264(.A(men_men_n286_), .B(i_2_), .Y(men_men_n287_));
  NO2        u265(.A(men_men_n56_), .B(i_6_), .Y(men_men_n288_));
  NO3        u266(.A(men_men_n135_), .B(men_men_n285_), .C(men_men_n281_), .Y(men_men_n289_));
  NO2        u267(.A(i_3_), .B(i_10_), .Y(men_men_n290_));
  NA3        u268(.A(men_men_n290_), .B(men_men_n39_), .C(men_men_n44_), .Y(men_men_n291_));
  NO2        u269(.A(i_2_), .B(men_men_n95_), .Y(men_men_n292_));
  NA2        u270(.A(i_1_), .B(men_men_n36_), .Y(men_men_n293_));
  NOi21      u271(.An(men_men_n211_), .B(men_men_n97_), .Y(men_men_n294_));
  NA3        u272(.A(men_men_n294_), .B(i_1_), .C(men_men_n292_), .Y(men_men_n295_));
  AN2        u273(.A(i_3_), .B(i_10_), .Y(men_men_n296_));
  NA3        u274(.A(men_men_n296_), .B(men_men_n168_), .C(men_men_n166_), .Y(men_men_n297_));
  NO2        u275(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n298_));
  OR2        u276(.A(men_men_n295_), .B(men_men_n291_), .Y(men_men_n299_));
  OAI220     u277(.A0(men_men_n299_), .A1(i_6_), .B0(men_men_n289_), .B1(men_men_n277_), .Y(men_men_n300_));
  NO4        u278(.A(men_men_n300_), .B(men_men_n275_), .C(men_men_n207_), .D(men_men_n161_), .Y(men_men_n301_));
  NO3        u279(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n302_));
  NO2        u280(.A(men_men_n56_), .B(men_men_n79_), .Y(men_men_n303_));
  NA2        u281(.A(men_men_n282_), .B(men_men_n303_), .Y(men_men_n304_));
  NO3        u282(.A(i_6_), .B(men_men_n185_), .C(i_7_), .Y(men_men_n305_));
  NA2        u283(.A(men_men_n305_), .B(men_men_n190_), .Y(men_men_n306_));
  AOI210     u284(.A0(men_men_n306_), .A1(men_men_n304_), .B0(i_5_), .Y(men_men_n307_));
  NO2        u285(.A(i_2_), .B(i_3_), .Y(men_men_n308_));
  OR2        u286(.A(i_0_), .B(i_5_), .Y(men_men_n309_));
  NA2        u287(.A(men_men_n211_), .B(men_men_n309_), .Y(men_men_n310_));
  NA4        u288(.A(men_men_n310_), .B(men_men_n228_), .C(men_men_n308_), .D(i_1_), .Y(men_men_n311_));
  NA3        u289(.A(men_men_n282_), .B(men_men_n278_), .C(men_men_n107_), .Y(men_men_n312_));
  NAi21      u290(.An(i_8_), .B(i_7_), .Y(men_men_n313_));
  NO2        u291(.A(men_men_n313_), .B(i_6_), .Y(men_men_n314_));
  NO2        u292(.A(men_men_n151_), .B(men_men_n46_), .Y(men_men_n315_));
  NA3        u293(.A(men_men_n315_), .B(men_men_n314_), .C(men_men_n157_), .Y(men_men_n316_));
  NA3        u294(.A(men_men_n316_), .B(men_men_n312_), .C(men_men_n311_), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n317_), .A1(men_men_n307_), .B0(i_4_), .Y(men_men_n318_));
  NO2        u296(.A(i_12_), .B(i_10_), .Y(men_men_n319_));
  NOi21      u297(.An(i_5_), .B(i_0_), .Y(men_men_n320_));
  AOI210     u298(.A0(i_2_), .A1(men_men_n48_), .B0(men_men_n95_), .Y(men_men_n321_));
  NO3        u299(.A(men_men_n321_), .B(men_men_n293_), .C(men_men_n122_), .Y(men_men_n322_));
  NA4        u300(.A(men_men_n78_), .B(men_men_n36_), .C(men_men_n79_), .D(i_8_), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n322_), .B(men_men_n319_), .Y(men_men_n324_));
  NO2        u302(.A(i_6_), .B(i_8_), .Y(men_men_n325_));
  NOi21      u303(.An(i_0_), .B(i_2_), .Y(men_men_n326_));
  AN2        u304(.A(men_men_n326_), .B(men_men_n325_), .Y(men_men_n327_));
  NO2        u305(.A(i_1_), .B(i_7_), .Y(men_men_n328_));
  NA3        u306(.A(men_men_n325_), .B(men_men_n41_), .C(i_5_), .Y(men_men_n329_));
  NA3        u307(.A(men_men_n329_), .B(men_men_n324_), .C(men_men_n318_), .Y(men_men_n330_));
  NO2        u308(.A(i_8_), .B(men_men_n310_), .Y(men_men_n331_));
  NO2        u309(.A(men_men_n97_), .B(men_men_n118_), .Y(men_men_n332_));
  OAI210     u310(.A0(men_men_n332_), .A1(men_men_n331_), .B0(i_3_), .Y(men_men_n333_));
  NO2        u311(.A(men_men_n286_), .B(men_men_n76_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n334_), .B(men_men_n126_), .Y(men_men_n335_));
  NA3        u313(.A(men_men_n294_), .B(i_8_), .C(men_men_n60_), .Y(men_men_n336_));
  AOI210     u314(.A0(men_men_n336_), .A1(men_men_n335_), .B0(i_7_), .Y(men_men_n337_));
  NO2        u315(.A(men_men_n185_), .B(i_9_), .Y(men_men_n338_));
  NA2        u316(.A(men_men_n338_), .B(men_men_n198_), .Y(men_men_n339_));
  NO2        u317(.A(men_men_n337_), .B(men_men_n285_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n340_), .A1(men_men_n333_), .B0(men_men_n156_), .Y(men_men_n341_));
  AOI210     u319(.A0(men_men_n330_), .A1(men_men_n302_), .B0(men_men_n341_), .Y(men_men_n342_));
  NOi32      u320(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n343_));
  INV        u321(.A(men_men_n343_), .Y(men_men_n344_));
  NAi21      u322(.An(i_0_), .B(i_6_), .Y(men_men_n345_));
  NAi21      u323(.An(i_1_), .B(i_5_), .Y(men_men_n346_));
  NA2        u324(.A(men_men_n346_), .B(men_men_n345_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n347_), .B(men_men_n25_), .Y(men_men_n348_));
  OAI210     u326(.A0(men_men_n348_), .A1(men_men_n153_), .B0(men_men_n239_), .Y(men_men_n349_));
  NAi41      u327(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n350_), .A1(men_men_n346_), .B0(men_men_n214_), .B1(men_men_n153_), .Y(men_men_n351_));
  AOI210     u329(.A0(men_men_n350_), .A1(men_men_n153_), .B0(men_men_n151_), .Y(men_men_n352_));
  NOi32      u330(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n353_));
  NA2        u331(.A(men_men_n353_), .B(men_men_n46_), .Y(men_men_n354_));
  NO2        u332(.A(men_men_n354_), .B(i_0_), .Y(men_men_n355_));
  OR3        u333(.A(men_men_n355_), .B(men_men_n352_), .C(men_men_n351_), .Y(men_men_n356_));
  NO2        u334(.A(i_1_), .B(men_men_n95_), .Y(men_men_n357_));
  NAi21      u335(.An(i_3_), .B(i_4_), .Y(men_men_n358_));
  NO2        u336(.A(men_men_n358_), .B(i_9_), .Y(men_men_n359_));
  AN2        u337(.A(i_6_), .B(i_7_), .Y(men_men_n360_));
  OAI210     u338(.A0(men_men_n360_), .A1(men_men_n357_), .B0(men_men_n359_), .Y(men_men_n361_));
  NA2        u339(.A(i_2_), .B(i_7_), .Y(men_men_n362_));
  NO2        u340(.A(men_men_n358_), .B(i_10_), .Y(men_men_n363_));
  AOI220     u341(.A0(men_men_n363_), .A1(men_men_n328_), .B0(men_men_n232_), .B1(men_men_n180_), .Y(men_men_n364_));
  NO2        u342(.A(men_men_n356_), .B(men_men_n349_), .Y(men_men_n365_));
  NO2        u343(.A(men_men_n365_), .B(men_men_n344_), .Y(men_men_n366_));
  NO2        u344(.A(men_men_n56_), .B(men_men_n25_), .Y(men_men_n367_));
  AN2        u345(.A(i_12_), .B(i_5_), .Y(men_men_n368_));
  NO2        u346(.A(i_4_), .B(men_men_n26_), .Y(men_men_n369_));
  NA2        u347(.A(men_men_n369_), .B(men_men_n368_), .Y(men_men_n370_));
  NO2        u348(.A(i_11_), .B(i_6_), .Y(men_men_n371_));
  NA3        u349(.A(men_men_n371_), .B(men_men_n315_), .C(men_men_n219_), .Y(men_men_n372_));
  NO2        u350(.A(men_men_n372_), .B(men_men_n370_), .Y(men_men_n373_));
  NO2        u351(.A(men_men_n236_), .B(i_5_), .Y(men_men_n374_));
  NO2        u352(.A(i_5_), .B(i_10_), .Y(men_men_n375_));
  NA2        u353(.A(men_men_n137_), .B(men_men_n45_), .Y(men_men_n376_));
  NO2        u354(.A(men_men_n376_), .B(men_men_n236_), .Y(men_men_n377_));
  OAI210     u355(.A0(men_men_n377_), .A1(men_men_n373_), .B0(men_men_n367_), .Y(men_men_n378_));
  NO2        u356(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n379_));
  INV        u357(.A(men_men_n143_), .Y(men_men_n380_));
  OAI210     u358(.A0(men_men_n380_), .A1(men_men_n373_), .B0(men_men_n379_), .Y(men_men_n381_));
  NO3        u359(.A(men_men_n79_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n382_));
  NO2        u360(.A(i_3_), .B(men_men_n95_), .Y(men_men_n383_));
  NA2        u361(.A(men_men_n290_), .B(men_men_n70_), .Y(men_men_n384_));
  NO2        u362(.A(i_11_), .B(i_12_), .Y(men_men_n385_));
  NA2        u363(.A(men_men_n385_), .B(men_men_n36_), .Y(men_men_n386_));
  NO2        u364(.A(men_men_n384_), .B(men_men_n386_), .Y(men_men_n387_));
  NA2        u365(.A(men_men_n375_), .B(men_men_n231_), .Y(men_men_n388_));
  NA3        u366(.A(men_men_n107_), .B(men_men_n41_), .C(i_11_), .Y(men_men_n389_));
  NO2        u367(.A(men_men_n389_), .B(men_men_n214_), .Y(men_men_n390_));
  NAi21      u368(.An(i_13_), .B(i_0_), .Y(men_men_n391_));
  NO2        u369(.A(men_men_n391_), .B(men_men_n233_), .Y(men_men_n392_));
  OAI210     u370(.A0(men_men_n390_), .A1(men_men_n387_), .B0(men_men_n392_), .Y(men_men_n393_));
  NA3        u371(.A(men_men_n393_), .B(men_men_n381_), .C(men_men_n378_), .Y(men_men_n394_));
  NO3        u372(.A(i_1_), .B(i_12_), .C(men_men_n79_), .Y(men_men_n395_));
  NO2        u373(.A(i_0_), .B(i_11_), .Y(men_men_n396_));
  AN2        u374(.A(i_1_), .B(i_6_), .Y(men_men_n397_));
  NOi21      u375(.An(i_2_), .B(i_12_), .Y(men_men_n398_));
  NA2        u376(.A(men_men_n398_), .B(men_men_n397_), .Y(men_men_n399_));
  INV        u377(.A(men_men_n399_), .Y(men_men_n400_));
  NA2        u378(.A(men_men_n135_), .B(i_9_), .Y(men_men_n401_));
  NO2        u379(.A(men_men_n401_), .B(i_4_), .Y(men_men_n402_));
  NA2        u380(.A(men_men_n400_), .B(men_men_n402_), .Y(men_men_n403_));
  OR2        u381(.A(i_13_), .B(i_10_), .Y(men_men_n404_));
  NO2        u382(.A(men_men_n165_), .B(men_men_n117_), .Y(men_men_n405_));
  OR2        u383(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n406_));
  NO2        u384(.A(men_men_n95_), .B(men_men_n25_), .Y(men_men_n407_));
  NA2        u385(.A(men_men_n276_), .B(men_men_n407_), .Y(men_men_n408_));
  OAI220     u386(.A0(men_men_n60_), .A1(men_men_n406_), .B0(men_men_n408_), .B1(men_men_n97_), .Y(men_men_n409_));
  INV        u387(.A(men_men_n409_), .Y(men_men_n410_));
  AOI210     u388(.A0(men_men_n410_), .A1(men_men_n403_), .B0(men_men_n26_), .Y(men_men_n411_));
  NA2        u389(.A(men_men_n312_), .B(men_men_n311_), .Y(men_men_n412_));
  AOI220     u390(.A0(men_men_n288_), .A1(men_men_n279_), .B0(men_men_n282_), .B1(men_men_n303_), .Y(men_men_n413_));
  NO2        u391(.A(men_men_n413_), .B(i_5_), .Y(men_men_n414_));
  NO2        u392(.A(men_men_n174_), .B(men_men_n79_), .Y(men_men_n415_));
  AOI220     u393(.A0(men_men_n415_), .A1(men_men_n287_), .B0(men_men_n271_), .B1(men_men_n203_), .Y(men_men_n416_));
  NO2        u394(.A(men_men_n416_), .B(i_7_), .Y(men_men_n417_));
  NO3        u395(.A(men_men_n417_), .B(men_men_n414_), .C(men_men_n412_), .Y(men_men_n418_));
  NA2        u396(.A(men_men_n188_), .B(men_men_n90_), .Y(men_men_n419_));
  AOI210     u397(.A0(men_men_n151_), .A1(men_men_n419_), .B0(men_men_n313_), .Y(men_men_n420_));
  NA3        u398(.A(men_men_n249_), .B(men_men_n61_), .C(i_2_), .Y(men_men_n421_));
  NA2        u399(.A(men_men_n288_), .B(men_men_n229_), .Y(men_men_n422_));
  OAI220     u400(.A0(men_men_n422_), .A1(men_men_n174_), .B0(men_men_n421_), .B1(men_men_n978_), .Y(men_men_n423_));
  NO2        u401(.A(i_3_), .B(men_men_n48_), .Y(men_men_n424_));
  NA2        u402(.A(men_men_n327_), .B(men_men_n424_), .Y(men_men_n425_));
  NA2        u403(.A(men_men_n305_), .B(men_men_n310_), .Y(men_men_n426_));
  OAI210     u404(.A0(men_men_n426_), .A1(men_men_n181_), .B0(men_men_n425_), .Y(men_men_n427_));
  NO3        u405(.A(men_men_n427_), .B(men_men_n423_), .C(men_men_n420_), .Y(men_men_n428_));
  AOI210     u406(.A0(men_men_n428_), .A1(men_men_n418_), .B0(men_men_n265_), .Y(men_men_n429_));
  NO4        u407(.A(men_men_n429_), .B(men_men_n411_), .C(men_men_n394_), .D(men_men_n366_), .Y(men_men_n430_));
  NO2        u408(.A(men_men_n68_), .B(i_13_), .Y(men_men_n431_));
  NO2        u409(.A(i_10_), .B(i_9_), .Y(men_men_n432_));
  NAi21      u410(.An(i_12_), .B(i_8_), .Y(men_men_n433_));
  NO2        u411(.A(men_men_n433_), .B(i_3_), .Y(men_men_n434_));
  NO2        u412(.A(men_men_n46_), .B(i_4_), .Y(men_men_n435_));
  NA2        u413(.A(men_men_n435_), .B(men_men_n98_), .Y(men_men_n436_));
  NO2        u414(.A(men_men_n436_), .B(men_men_n197_), .Y(men_men_n437_));
  NA2        u415(.A(men_men_n298_), .B(i_0_), .Y(men_men_n438_));
  NO3        u416(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n439_));
  NA2        u417(.A(men_men_n260_), .B(men_men_n91_), .Y(men_men_n440_));
  NA2        u418(.A(men_men_n440_), .B(men_men_n439_), .Y(men_men_n441_));
  NA2        u419(.A(i_8_), .B(i_9_), .Y(men_men_n442_));
  NO2        u420(.A(men_men_n441_), .B(men_men_n438_), .Y(men_men_n443_));
  NO3        u421(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n444_));
  NA3        u422(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n445_));
  NO2        u423(.A(men_men_n443_), .B(men_men_n437_), .Y(men_men_n446_));
  NA2        u424(.A(men_men_n287_), .B(men_men_n102_), .Y(men_men_n447_));
  OA220      u425(.A0(men_men_n339_), .A1(men_men_n156_), .B0(men_men_n447_), .B1(men_men_n226_), .Y(men_men_n448_));
  NA2        u426(.A(men_men_n90_), .B(i_13_), .Y(men_men_n449_));
  NA2        u427(.A(men_men_n415_), .B(men_men_n367_), .Y(men_men_n450_));
  NO2        u428(.A(i_2_), .B(i_13_), .Y(men_men_n451_));
  NA3        u429(.A(men_men_n451_), .B(men_men_n155_), .C(men_men_n93_), .Y(men_men_n452_));
  OAI220     u430(.A0(men_men_n452_), .A1(men_men_n231_), .B0(men_men_n450_), .B1(men_men_n449_), .Y(men_men_n453_));
  NO3        u431(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n454_));
  NO2        u432(.A(i_6_), .B(i_7_), .Y(men_men_n455_));
  NA2        u433(.A(men_men_n455_), .B(men_men_n454_), .Y(men_men_n456_));
  NO2        u434(.A(i_11_), .B(i_1_), .Y(men_men_n457_));
  OR2        u435(.A(i_11_), .B(i_8_), .Y(men_men_n458_));
  NOi21      u436(.An(i_2_), .B(i_7_), .Y(men_men_n459_));
  NAi31      u437(.An(men_men_n458_), .B(men_men_n459_), .C(i_0_), .Y(men_men_n460_));
  NO2        u438(.A(men_men_n404_), .B(i_6_), .Y(men_men_n461_));
  NA3        u439(.A(men_men_n461_), .B(i_1_), .C(men_men_n70_), .Y(men_men_n462_));
  NO2        u440(.A(men_men_n462_), .B(men_men_n460_), .Y(men_men_n463_));
  NO2        u441(.A(i_3_), .B(men_men_n185_), .Y(men_men_n464_));
  NO2        u442(.A(i_6_), .B(i_10_), .Y(men_men_n465_));
  NA4        u443(.A(men_men_n465_), .B(men_men_n302_), .C(men_men_n464_), .D(men_men_n231_), .Y(men_men_n466_));
  NO2        u444(.A(men_men_n466_), .B(men_men_n149_), .Y(men_men_n467_));
  NA3        u445(.A(men_men_n238_), .B(men_men_n164_), .C(men_men_n126_), .Y(men_men_n468_));
  NA2        u446(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n469_));
  NO2        u447(.A(men_men_n151_), .B(i_3_), .Y(men_men_n470_));
  NAi31      u448(.An(men_men_n469_), .B(men_men_n470_), .C(men_men_n220_), .Y(men_men_n471_));
  NA3        u449(.A(men_men_n379_), .B(men_men_n171_), .C(men_men_n142_), .Y(men_men_n472_));
  NA3        u450(.A(men_men_n472_), .B(men_men_n471_), .C(men_men_n468_), .Y(men_men_n473_));
  NO4        u451(.A(men_men_n473_), .B(men_men_n467_), .C(men_men_n463_), .D(men_men_n453_), .Y(men_men_n474_));
  NA2        u452(.A(men_men_n439_), .B(men_men_n368_), .Y(men_men_n475_));
  NAi21      u453(.An(men_men_n209_), .B(men_men_n385_), .Y(men_men_n476_));
  NO2        u454(.A(men_men_n26_), .B(i_5_), .Y(men_men_n477_));
  NO2        u455(.A(i_0_), .B(men_men_n79_), .Y(men_men_n478_));
  NA3        u456(.A(men_men_n478_), .B(men_men_n477_), .C(men_men_n135_), .Y(men_men_n479_));
  NO2        u457(.A(men_men_n38_), .B(men_men_n479_), .Y(men_men_n480_));
  NA2        u458(.A(men_men_n302_), .B(men_men_n232_), .Y(men_men_n481_));
  NO2        u459(.A(men_men_n481_), .B(men_men_n421_), .Y(men_men_n482_));
  NA4        u460(.A(men_men_n296_), .B(men_men_n217_), .C(men_men_n68_), .D(men_men_n231_), .Y(men_men_n483_));
  NO2        u461(.A(men_men_n483_), .B(men_men_n456_), .Y(men_men_n484_));
  NO3        u462(.A(men_men_n484_), .B(men_men_n482_), .C(men_men_n480_), .Y(men_men_n485_));
  NA4        u463(.A(men_men_n485_), .B(men_men_n474_), .C(men_men_n448_), .D(men_men_n446_), .Y(men_men_n486_));
  NA3        u464(.A(men_men_n296_), .B(men_men_n168_), .C(men_men_n166_), .Y(men_men_n487_));
  OAI210     u465(.A0(men_men_n291_), .A1(men_men_n172_), .B0(men_men_n487_), .Y(men_men_n488_));
  AN2        u466(.A(men_men_n279_), .B(men_men_n228_), .Y(men_men_n489_));
  NA2        u467(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n490_));
  NA2        u468(.A(men_men_n116_), .B(men_men_n106_), .Y(men_men_n491_));
  AN2        u469(.A(men_men_n491_), .B(men_men_n439_), .Y(men_men_n492_));
  OAI210     u470(.A0(i_2_), .A1(men_men_n226_), .B0(men_men_n297_), .Y(men_men_n493_));
  AOI220     u471(.A0(men_men_n493_), .A1(men_men_n314_), .B0(men_men_n492_), .B1(men_men_n298_), .Y(men_men_n494_));
  NA2        u472(.A(men_men_n368_), .B(men_men_n219_), .Y(men_men_n495_));
  NA2        u473(.A(men_men_n343_), .B(men_men_n68_), .Y(men_men_n496_));
  NA2        u474(.A(men_men_n360_), .B(men_men_n353_), .Y(men_men_n497_));
  OR2        u475(.A(men_men_n495_), .B(men_men_n497_), .Y(men_men_n498_));
  NO2        u476(.A(men_men_n36_), .B(i_8_), .Y(men_men_n499_));
  INV        u477(.A(men_men_n498_), .Y(men_men_n500_));
  OAI210     u478(.A0(i_8_), .A1(men_men_n60_), .B0(men_men_n128_), .Y(men_men_n501_));
  INV        u479(.A(men_men_n259_), .Y(men_men_n502_));
  NO2        u480(.A(men_men_n502_), .B(men_men_n191_), .Y(men_men_n503_));
  AOI220     u481(.A0(i_6_), .A1(men_men_n503_), .B0(men_men_n501_), .B1(men_men_n405_), .Y(men_men_n504_));
  NA4        u482(.A(men_men_n504_), .B(men_men_n498_), .C(men_men_n494_), .D(men_men_n490_), .Y(men_men_n505_));
  NA2        u483(.A(men_men_n374_), .B(men_men_n287_), .Y(men_men_n506_));
  OAI210     u484(.A0(men_men_n370_), .A1(men_men_n162_), .B0(men_men_n506_), .Y(men_men_n507_));
  NO2        u485(.A(i_12_), .B(men_men_n185_), .Y(men_men_n508_));
  NA2        u486(.A(men_men_n508_), .B(men_men_n219_), .Y(men_men_n509_));
  NO2        u487(.A(men_men_n404_), .B(men_men_n38_), .Y(men_men_n510_));
  NA2        u488(.A(men_men_n510_), .B(men_men_n507_), .Y(men_men_n511_));
  NO2        u489(.A(i_8_), .B(i_7_), .Y(men_men_n512_));
  AOI220     u490(.A0(men_men_n315_), .A1(men_men_n39_), .B0(men_men_n229_), .B1(men_men_n200_), .Y(men_men_n513_));
  OAI220     u491(.A0(men_men_n513_), .A1(men_men_n174_), .B0(i_5_), .B1(men_men_n236_), .Y(men_men_n514_));
  NA2        u492(.A(men_men_n44_), .B(i_10_), .Y(men_men_n515_));
  NO2        u493(.A(men_men_n515_), .B(i_6_), .Y(men_men_n516_));
  NA3        u494(.A(men_men_n516_), .B(men_men_n514_), .C(men_men_n512_), .Y(men_men_n517_));
  AOI220     u495(.A0(men_men_n415_), .A1(men_men_n315_), .B0(men_men_n240_), .B1(men_men_n237_), .Y(men_men_n518_));
  OAI220     u496(.A0(men_men_n518_), .A1(men_men_n256_), .B0(men_men_n449_), .B1(men_men_n127_), .Y(men_men_n519_));
  NA2        u497(.A(men_men_n519_), .B(men_men_n259_), .Y(men_men_n520_));
  NOi31      u498(.An(men_men_n282_), .B(men_men_n291_), .C(men_men_n172_), .Y(men_men_n521_));
  NA3        u499(.A(men_men_n296_), .B(men_men_n166_), .C(men_men_n90_), .Y(men_men_n522_));
  NO2        u500(.A(men_men_n151_), .B(i_5_), .Y(men_men_n523_));
  NA2        u501(.A(men_men_n523_), .B(men_men_n308_), .Y(men_men_n524_));
  NA2        u502(.A(men_men_n524_), .B(men_men_n522_), .Y(men_men_n525_));
  OAI210     u503(.A0(men_men_n525_), .A1(men_men_n521_), .B0(men_men_n444_), .Y(men_men_n526_));
  NA4        u504(.A(men_men_n526_), .B(men_men_n520_), .C(men_men_n517_), .D(men_men_n511_), .Y(men_men_n527_));
  NA2        u505(.A(men_men_n276_), .B(men_men_n78_), .Y(men_men_n528_));
  NO2        u506(.A(men_men_n335_), .B(men_men_n528_), .Y(men_men_n529_));
  NA2        u507(.A(men_men_n288_), .B(men_men_n279_), .Y(men_men_n530_));
  NO2        u508(.A(men_men_n530_), .B(men_men_n165_), .Y(men_men_n531_));
  NA2        u509(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n532_));
  NA2        u510(.A(men_men_n432_), .B(men_men_n215_), .Y(men_men_n533_));
  NO2        u511(.A(men_men_n532_), .B(men_men_n533_), .Y(men_men_n534_));
  NA3        u512(.A(men_men_n508_), .B(men_men_n267_), .C(i_5_), .Y(men_men_n535_));
  NO2        u513(.A(i_1_), .B(men_men_n535_), .Y(men_men_n536_));
  NO4        u514(.A(men_men_n536_), .B(men_men_n534_), .C(men_men_n531_), .D(men_men_n529_), .Y(men_men_n537_));
  NO4        u515(.A(men_men_n245_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n538_));
  NO3        u516(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n539_));
  NO2        u517(.A(men_men_n227_), .B(men_men_n36_), .Y(men_men_n540_));
  AN2        u518(.A(men_men_n540_), .B(men_men_n539_), .Y(men_men_n541_));
  OA210      u519(.A0(men_men_n541_), .A1(men_men_n538_), .B0(men_men_n343_), .Y(men_men_n542_));
  NO2        u520(.A(men_men_n404_), .B(i_1_), .Y(men_men_n543_));
  NOi31      u521(.An(men_men_n543_), .B(men_men_n440_), .C(men_men_n68_), .Y(men_men_n544_));
  AN3        u522(.A(men_men_n544_), .B(men_men_n402_), .C(men_men_n477_), .Y(men_men_n545_));
  NO2        u523(.A(men_men_n413_), .B(men_men_n169_), .Y(men_men_n546_));
  NO3        u524(.A(men_men_n546_), .B(men_men_n545_), .C(men_men_n542_), .Y(men_men_n547_));
  NO2        u525(.A(men_men_n79_), .B(men_men_n25_), .Y(men_men_n548_));
  NA2        u526(.A(men_men_n276_), .B(men_men_n548_), .Y(men_men_n549_));
  NO2        u527(.A(men_men_n549_), .B(men_men_n438_), .Y(men_men_n550_));
  NO2        u528(.A(men_men_n109_), .B(men_men_n23_), .Y(men_men_n551_));
  INV        u529(.A(men_men_n305_), .Y(men_men_n552_));
  AOI220     u530(.A0(men_men_n552_), .A1(men_men_n422_), .B0(men_men_n175_), .B1(men_men_n173_), .Y(men_men_n553_));
  NOi21      u531(.An(men_men_n139_), .B(men_men_n323_), .Y(men_men_n554_));
  NO3        u532(.A(men_men_n554_), .B(men_men_n553_), .C(men_men_n550_), .Y(men_men_n555_));
  NO2        u533(.A(men_men_n496_), .B(men_men_n364_), .Y(men_men_n556_));
  NO2        u534(.A(i_12_), .B(men_men_n79_), .Y(men_men_n557_));
  NA3        u535(.A(men_men_n557_), .B(men_men_n267_), .C(i_5_), .Y(men_men_n558_));
  NO2        u536(.A(men_men_n558_), .B(i_3_), .Y(men_men_n559_));
  NA2        u537(.A(men_men_n166_), .B(i_0_), .Y(men_men_n560_));
  NO3        u538(.A(men_men_n560_), .B(men_men_n977_), .C(men_men_n291_), .Y(men_men_n561_));
  OR2        u539(.A(i_2_), .B(i_5_), .Y(men_men_n562_));
  OR2        u540(.A(men_men_n562_), .B(men_men_n397_), .Y(men_men_n563_));
  AOI210     u541(.A0(men_men_n362_), .A1(men_men_n237_), .B0(men_men_n190_), .Y(men_men_n564_));
  AOI210     u542(.A0(men_men_n564_), .A1(men_men_n563_), .B0(men_men_n476_), .Y(men_men_n565_));
  NO4        u543(.A(men_men_n565_), .B(men_men_n561_), .C(men_men_n559_), .D(men_men_n556_), .Y(men_men_n566_));
  NA4        u544(.A(men_men_n566_), .B(men_men_n555_), .C(men_men_n547_), .D(men_men_n537_), .Y(men_men_n567_));
  NO4        u545(.A(men_men_n567_), .B(men_men_n527_), .C(men_men_n505_), .D(men_men_n486_), .Y(men_men_n568_));
  NA4        u546(.A(men_men_n568_), .B(men_men_n430_), .C(men_men_n342_), .D(men_men_n301_), .Y(men7));
  NO2        u547(.A(men_men_n86_), .B(men_men_n52_), .Y(men_men_n570_));
  NO2        u548(.A(men_men_n102_), .B(men_men_n83_), .Y(men_men_n571_));
  NA2        u549(.A(men_men_n369_), .B(men_men_n571_), .Y(men_men_n572_));
  NA2        u550(.A(men_men_n465_), .B(men_men_n78_), .Y(men_men_n573_));
  NA2        u551(.A(men_men_n137_), .B(i_8_), .Y(men_men_n574_));
  OAI210     u552(.A0(men_men_n574_), .A1(men_men_n573_), .B0(men_men_n572_), .Y(men_men_n575_));
  NA3        u553(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n576_));
  NO2        u554(.A(men_men_n231_), .B(i_4_), .Y(men_men_n577_));
  NA2        u555(.A(men_men_n577_), .B(i_8_), .Y(men_men_n578_));
  NA2        u556(.A(i_2_), .B(men_men_n79_), .Y(men_men_n579_));
  OAI210     u557(.A0(men_men_n82_), .A1(men_men_n195_), .B0(men_men_n196_), .Y(men_men_n580_));
  NA2        u558(.A(i_4_), .B(i_8_), .Y(men_men_n581_));
  NA2        u559(.A(men_men_n581_), .B(men_men_n296_), .Y(men_men_n582_));
  OAI220     u560(.A0(men_men_n582_), .A1(men_men_n579_), .B0(men_men_n580_), .B1(i_13_), .Y(men_men_n583_));
  NO3        u561(.A(men_men_n583_), .B(men_men_n575_), .C(men_men_n570_), .Y(men_men_n584_));
  AOI210     u562(.A0(men_men_n122_), .A1(men_men_n59_), .B0(i_10_), .Y(men_men_n585_));
  AOI210     u563(.A0(men_men_n585_), .A1(men_men_n231_), .B0(men_men_n155_), .Y(men_men_n586_));
  OR2        u564(.A(i_6_), .B(i_10_), .Y(men_men_n587_));
  NO2        u565(.A(men_men_n587_), .B(men_men_n23_), .Y(men_men_n588_));
  OR3        u566(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n589_));
  NO3        u567(.A(men_men_n589_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n590_));
  INV        u568(.A(men_men_n192_), .Y(men_men_n591_));
  INV        u569(.A(men_men_n590_), .Y(men_men_n592_));
  OA220      u570(.A0(men_men_n592_), .A1(i_3_), .B0(men_men_n586_), .B1(men_men_n261_), .Y(men_men_n593_));
  AOI210     u571(.A0(men_men_n593_), .A1(men_men_n584_), .B0(men_men_n60_), .Y(men_men_n594_));
  NOi21      u572(.An(i_11_), .B(i_7_), .Y(men_men_n595_));
  AO210      u573(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n596_));
  NO2        u574(.A(men_men_n596_), .B(men_men_n595_), .Y(men_men_n597_));
  NA3        u575(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n598_));
  NAi31      u576(.An(men_men_n598_), .B(men_men_n208_), .C(i_11_), .Y(men_men_n599_));
  NO2        u577(.A(men_men_n599_), .B(men_men_n60_), .Y(men_men_n600_));
  NA2        u578(.A(men_men_n81_), .B(men_men_n60_), .Y(men_men_n601_));
  AO210      u579(.A0(men_men_n601_), .A1(men_men_n364_), .B0(men_men_n40_), .Y(men_men_n602_));
  NO2        u580(.A(men_men_n60_), .B(i_9_), .Y(men_men_n603_));
  NA2        u581(.A(men_men_n60_), .B(men_men_n985_), .Y(men_men_n604_));
  NO2        u582(.A(i_1_), .B(i_12_), .Y(men_men_n605_));
  NA2        u583(.A(men_men_n604_), .B(men_men_n602_), .Y(men_men_n606_));
  OAI210     u584(.A0(men_men_n606_), .A1(men_men_n600_), .B0(i_6_), .Y(men_men_n607_));
  NO2        u585(.A(i_6_), .B(i_11_), .Y(men_men_n608_));
  INV        u586(.A(men_men_n441_), .Y(men_men_n609_));
  NO4        u587(.A(men_men_n208_), .B(men_men_n122_), .C(i_13_), .D(men_men_n79_), .Y(men_men_n610_));
  NA2        u588(.A(men_men_n610_), .B(men_men_n603_), .Y(men_men_n611_));
  NO3        u589(.A(men_men_n587_), .B(men_men_n227_), .C(men_men_n23_), .Y(men_men_n612_));
  AOI210     u590(.A0(i_1_), .A1(men_men_n252_), .B0(men_men_n612_), .Y(men_men_n613_));
  OAI210     u591(.A0(men_men_n613_), .A1(men_men_n44_), .B0(men_men_n611_), .Y(men_men_n614_));
  NA3        u592(.A(men_men_n512_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n615_));
  NA2        u593(.A(men_men_n132_), .B(i_9_), .Y(men_men_n616_));
  NA3        u594(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n617_));
  NO2        u595(.A(men_men_n46_), .B(i_1_), .Y(men_men_n618_));
  NA3        u596(.A(men_men_n618_), .B(men_men_n260_), .C(men_men_n44_), .Y(men_men_n619_));
  OAI220     u597(.A0(men_men_n619_), .A1(men_men_n617_), .B0(men_men_n616_), .B1(men_men_n974_), .Y(men_men_n620_));
  NA3        u598(.A(men_men_n603_), .B(men_men_n308_), .C(i_6_), .Y(men_men_n621_));
  NO2        u599(.A(men_men_n621_), .B(men_men_n23_), .Y(men_men_n622_));
  AOI210     u600(.A0(men_men_n457_), .A1(men_men_n407_), .B0(men_men_n235_), .Y(men_men_n623_));
  NO2        u601(.A(men_men_n623_), .B(men_men_n579_), .Y(men_men_n624_));
  NAi21      u602(.An(men_men_n615_), .B(men_men_n85_), .Y(men_men_n625_));
  NA2        u603(.A(men_men_n618_), .B(men_men_n260_), .Y(men_men_n626_));
  NO2        u604(.A(i_11_), .B(men_men_n37_), .Y(men_men_n627_));
  NA2        u605(.A(men_men_n627_), .B(men_men_n24_), .Y(men_men_n628_));
  OAI210     u606(.A0(men_men_n628_), .A1(men_men_n626_), .B0(men_men_n625_), .Y(men_men_n629_));
  OR4        u607(.A(men_men_n629_), .B(men_men_n624_), .C(men_men_n622_), .D(men_men_n620_), .Y(men_men_n630_));
  NO3        u608(.A(men_men_n630_), .B(men_men_n614_), .C(men_men_n609_), .Y(men_men_n631_));
  NO2        u609(.A(men_men_n231_), .B(men_men_n95_), .Y(men_men_n632_));
  NO2        u610(.A(men_men_n632_), .B(men_men_n595_), .Y(men_men_n633_));
  NA2        u611(.A(men_men_n633_), .B(i_1_), .Y(men_men_n634_));
  NO2        u612(.A(men_men_n634_), .B(men_men_n589_), .Y(men_men_n635_));
  NA2        u613(.A(men_men_n635_), .B(men_men_n46_), .Y(men_men_n636_));
  NO2        u614(.A(men_men_n980_), .B(men_men_n109_), .Y(men_men_n637_));
  AN2        u615(.A(men_men_n637_), .B(men_men_n516_), .Y(men_men_n638_));
  NO2        u616(.A(men_men_n227_), .B(men_men_n44_), .Y(men_men_n639_));
  NO3        u617(.A(men_men_n639_), .B(men_men_n298_), .C(i_11_), .Y(men_men_n640_));
  NO2        u618(.A(men_men_n111_), .B(men_men_n37_), .Y(men_men_n641_));
  NO2        u619(.A(men_men_n641_), .B(i_6_), .Y(men_men_n642_));
  NO2        u620(.A(men_men_n79_), .B(i_9_), .Y(men_men_n643_));
  NO2        u621(.A(men_men_n643_), .B(men_men_n60_), .Y(men_men_n644_));
  NO2        u622(.A(men_men_n644_), .B(men_men_n605_), .Y(men_men_n645_));
  NO4        u623(.A(men_men_n645_), .B(men_men_n642_), .C(men_men_n640_), .D(i_4_), .Y(men_men_n646_));
  NA2        u624(.A(i_1_), .B(i_3_), .Y(men_men_n647_));
  NO2        u625(.A(men_men_n442_), .B(men_men_n86_), .Y(men_men_n648_));
  AOI210     u626(.A0(men_men_n639_), .A1(i_10_), .B0(men_men_n648_), .Y(men_men_n649_));
  NO2        u627(.A(men_men_n649_), .B(men_men_n647_), .Y(men_men_n650_));
  NO3        u628(.A(men_men_n650_), .B(men_men_n646_), .C(men_men_n638_), .Y(men_men_n651_));
  NA4        u629(.A(men_men_n651_), .B(men_men_n636_), .C(men_men_n631_), .D(men_men_n607_), .Y(men_men_n652_));
  NO3        u630(.A(men_men_n458_), .B(i_3_), .C(i_7_), .Y(men_men_n653_));
  NOi21      u631(.An(men_men_n653_), .B(i_10_), .Y(men_men_n654_));
  AN2        u632(.A(men_men_n238_), .B(men_men_n79_), .Y(men_men_n655_));
  NA2        u633(.A(men_men_n360_), .B(men_men_n359_), .Y(men_men_n656_));
  NA3        u634(.A(men_men_n465_), .B(men_men_n499_), .C(men_men_n46_), .Y(men_men_n657_));
  NO3        u635(.A(men_men_n459_), .B(men_men_n581_), .C(men_men_n79_), .Y(men_men_n658_));
  NA2        u636(.A(men_men_n658_), .B(men_men_n25_), .Y(men_men_n659_));
  NA3        u637(.A(men_men_n155_), .B(men_men_n78_), .C(men_men_n79_), .Y(men_men_n660_));
  NA4        u638(.A(men_men_n660_), .B(men_men_n659_), .C(men_men_n657_), .D(men_men_n656_), .Y(men_men_n661_));
  OAI210     u639(.A0(men_men_n661_), .A1(men_men_n655_), .B0(i_1_), .Y(men_men_n662_));
  AOI210     u640(.A0(men_men_n260_), .A1(men_men_n91_), .B0(i_1_), .Y(men_men_n663_));
  NO2        u641(.A(men_men_n358_), .B(i_2_), .Y(men_men_n664_));
  NA2        u642(.A(men_men_n664_), .B(men_men_n663_), .Y(men_men_n665_));
  OAI210     u643(.A0(men_men_n621_), .A1(men_men_n433_), .B0(men_men_n665_), .Y(men_men_n666_));
  INV        u644(.A(men_men_n666_), .Y(men_men_n667_));
  AOI210     u645(.A0(men_men_n667_), .A1(men_men_n662_), .B0(i_13_), .Y(men_men_n668_));
  OR2        u646(.A(i_11_), .B(i_7_), .Y(men_men_n669_));
  NA3        u647(.A(men_men_n669_), .B(men_men_n100_), .C(men_men_n132_), .Y(men_men_n670_));
  AOI220     u648(.A0(men_men_n451_), .A1(men_men_n155_), .B0(men_men_n435_), .B1(men_men_n132_), .Y(men_men_n671_));
  OAI210     u649(.A0(men_men_n671_), .A1(men_men_n44_), .B0(men_men_n670_), .Y(men_men_n672_));
  NA2        u650(.A(men_men_n238_), .B(men_men_n125_), .Y(men_men_n673_));
  NO2        u651(.A(men_men_n673_), .B(men_men_n40_), .Y(men_men_n674_));
  AOI210     u652(.A0(men_men_n672_), .A1(men_men_n325_), .B0(men_men_n674_), .Y(men_men_n675_));
  AOI220     u653(.A0(i_7_), .A1(men_men_n67_), .B0(men_men_n371_), .B1(men_men_n618_), .Y(men_men_n676_));
  NO2        u654(.A(men_men_n676_), .B(men_men_n236_), .Y(men_men_n677_));
  NA2        u655(.A(men_men_n121_), .B(i_13_), .Y(men_men_n678_));
  NO2        u656(.A(men_men_n617_), .B(men_men_n109_), .Y(men_men_n679_));
  INV        u657(.A(men_men_n679_), .Y(men_men_n680_));
  OAI220     u658(.A0(men_men_n680_), .A1(men_men_n66_), .B0(men_men_n678_), .B1(men_men_n663_), .Y(men_men_n681_));
  NO3        u659(.A(men_men_n66_), .B(men_men_n32_), .C(men_men_n95_), .Y(men_men_n682_));
  NA2        u660(.A(men_men_n26_), .B(men_men_n185_), .Y(men_men_n683_));
  NA2        u661(.A(men_men_n683_), .B(i_7_), .Y(men_men_n684_));
  NO3        u662(.A(men_men_n459_), .B(men_men_n231_), .C(men_men_n79_), .Y(men_men_n685_));
  AOI210     u663(.A0(men_men_n685_), .A1(men_men_n684_), .B0(men_men_n682_), .Y(men_men_n686_));
  NO2        u664(.A(men_men_n686_), .B(men_men_n591_), .Y(men_men_n687_));
  NO3        u665(.A(men_men_n687_), .B(men_men_n681_), .C(men_men_n677_), .Y(men_men_n688_));
  OR2        u666(.A(i_11_), .B(i_6_), .Y(men_men_n689_));
  NA3        u667(.A(men_men_n577_), .B(men_men_n683_), .C(i_7_), .Y(men_men_n690_));
  AOI210     u668(.A0(men_men_n690_), .A1(men_men_n680_), .B0(men_men_n689_), .Y(men_men_n691_));
  NA2        u669(.A(men_men_n608_), .B(i_13_), .Y(men_men_n692_));
  NA2        u670(.A(men_men_n96_), .B(men_men_n683_), .Y(men_men_n693_));
  NAi21      u671(.An(i_11_), .B(i_12_), .Y(men_men_n694_));
  NOi41      u672(.An(men_men_n105_), .B(men_men_n694_), .C(i_13_), .D(men_men_n79_), .Y(men_men_n695_));
  NO2        u673(.A(men_men_n459_), .B(men_men_n581_), .Y(men_men_n696_));
  AOI220     u674(.A0(men_men_n696_), .A1(men_men_n302_), .B0(men_men_n695_), .B1(men_men_n693_), .Y(men_men_n697_));
  NA2        u675(.A(men_men_n697_), .B(men_men_n692_), .Y(men_men_n698_));
  OAI210     u676(.A0(men_men_n698_), .A1(men_men_n691_), .B0(men_men_n60_), .Y(men_men_n699_));
  NO2        u677(.A(i_2_), .B(i_12_), .Y(men_men_n700_));
  NA2        u678(.A(men_men_n357_), .B(men_men_n700_), .Y(men_men_n701_));
  OAI210     u679(.A0(i_8_), .A1(men_men_n359_), .B0(men_men_n357_), .Y(men_men_n702_));
  NO2        u680(.A(men_men_n122_), .B(i_2_), .Y(men_men_n703_));
  NA2        u681(.A(men_men_n703_), .B(men_men_n605_), .Y(men_men_n704_));
  NA3        u682(.A(men_men_n704_), .B(men_men_n702_), .C(men_men_n701_), .Y(men_men_n705_));
  NA3        u683(.A(men_men_n705_), .B(men_men_n45_), .C(men_men_n219_), .Y(men_men_n706_));
  NA4        u684(.A(men_men_n706_), .B(men_men_n699_), .C(men_men_n688_), .D(men_men_n675_), .Y(men_men_n707_));
  OR4        u685(.A(men_men_n707_), .B(men_men_n668_), .C(men_men_n652_), .D(men_men_n594_), .Y(men5));
  AOI210     u686(.A0(men_men_n633_), .A1(men_men_n263_), .B0(men_men_n405_), .Y(men_men_n709_));
  NO2        u687(.A(men_men_n578_), .B(i_11_), .Y(men_men_n710_));
  NA2        u688(.A(men_men_n82_), .B(men_men_n710_), .Y(men_men_n711_));
  NA2        u689(.A(men_men_n711_), .B(men_men_n709_), .Y(men_men_n712_));
  NO3        u690(.A(i_11_), .B(men_men_n231_), .C(i_13_), .Y(men_men_n713_));
  NO2        u691(.A(men_men_n118_), .B(men_men_n23_), .Y(men_men_n714_));
  NA2        u692(.A(i_12_), .B(i_8_), .Y(men_men_n715_));
  INV        u693(.A(men_men_n715_), .Y(men_men_n716_));
  INV        u694(.A(men_men_n432_), .Y(men_men_n717_));
  AOI220     u695(.A0(men_men_n308_), .A1(men_men_n551_), .B0(men_men_n716_), .B1(men_men_n714_), .Y(men_men_n718_));
  INV        u696(.A(men_men_n718_), .Y(men_men_n719_));
  NO2        u697(.A(men_men_n719_), .B(men_men_n712_), .Y(men_men_n720_));
  INV        u698(.A(men_men_n164_), .Y(men_men_n721_));
  OAI210     u699(.A0(men_men_n664_), .A1(men_men_n434_), .B0(men_men_n105_), .Y(men_men_n722_));
  NO2        u700(.A(men_men_n722_), .B(men_men_n721_), .Y(men_men_n723_));
  NO2        u701(.A(men_men_n442_), .B(men_men_n26_), .Y(men_men_n724_));
  NO2        u702(.A(men_men_n724_), .B(men_men_n407_), .Y(men_men_n725_));
  NA2        u703(.A(men_men_n725_), .B(i_2_), .Y(men_men_n726_));
  INV        u704(.A(men_men_n726_), .Y(men_men_n727_));
  AOI210     u705(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n404_), .Y(men_men_n728_));
  AOI210     u706(.A0(men_men_n728_), .A1(men_men_n727_), .B0(men_men_n723_), .Y(men_men_n729_));
  OA210      u707(.A0(men_men_n597_), .A1(men_men_n120_), .B0(i_13_), .Y(men_men_n730_));
  NA2        u708(.A(men_men_n192_), .B(men_men_n195_), .Y(men_men_n731_));
  NA2        u709(.A(men_men_n145_), .B(i_8_), .Y(men_men_n732_));
  AOI210     u710(.A0(men_men_n732_), .A1(men_men_n731_), .B0(men_men_n362_), .Y(men_men_n733_));
  AOI210     u711(.A0(men_men_n201_), .A1(men_men_n141_), .B0(men_men_n499_), .Y(men_men_n734_));
  NA2        u712(.A(men_men_n734_), .B(men_men_n407_), .Y(men_men_n735_));
  NO2        u713(.A(men_men_n96_), .B(men_men_n44_), .Y(men_men_n736_));
  INV        u714(.A(men_men_n292_), .Y(men_men_n737_));
  NA4        u715(.A(men_men_n737_), .B(men_men_n296_), .C(men_men_n118_), .D(men_men_n42_), .Y(men_men_n738_));
  OAI210     u716(.A0(men_men_n738_), .A1(men_men_n736_), .B0(men_men_n735_), .Y(men_men_n739_));
  NO3        u717(.A(men_men_n739_), .B(men_men_n733_), .C(men_men_n730_), .Y(men_men_n740_));
  NA2        u718(.A(men_men_n551_), .B(men_men_n28_), .Y(men_men_n741_));
  NA2        u719(.A(men_men_n713_), .B(men_men_n268_), .Y(men_men_n742_));
  NA2        u720(.A(men_men_n742_), .B(men_men_n741_), .Y(men_men_n743_));
  AOI220     u721(.A0(men_men_n120_), .A1(men_men_n36_), .B0(men_men_n743_), .B1(men_men_n46_), .Y(men_men_n744_));
  NA4        u722(.A(men_men_n744_), .B(men_men_n740_), .C(men_men_n729_), .D(men_men_n720_), .Y(men6));
  NA2        u723(.A(men_men_n981_), .B(men_men_n703_), .Y(men_men_n746_));
  NA4        u724(.A(men_men_n375_), .B(men_men_n464_), .C(men_men_n66_), .D(men_men_n95_), .Y(men_men_n747_));
  INV        u725(.A(men_men_n747_), .Y(men_men_n748_));
  NO2        u726(.A(men_men_n214_), .B(men_men_n469_), .Y(men_men_n749_));
  INV        u727(.A(i_9_), .Y(men_men_n750_));
  NO2        u728(.A(men_men_n748_), .B(men_men_n320_), .Y(men_men_n751_));
  AO210      u729(.A0(men_men_n751_), .A1(men_men_n746_), .B0(i_12_), .Y(men_men_n752_));
  NA2        u730(.A(men_men_n363_), .B(men_men_n328_), .Y(men_men_n753_));
  NA2        u731(.A(men_men_n557_), .B(men_men_n60_), .Y(men_men_n754_));
  NA2        u732(.A(men_men_n654_), .B(men_men_n66_), .Y(men_men_n755_));
  NA4        u733(.A(men_men_n601_), .B(men_men_n755_), .C(men_men_n754_), .D(men_men_n753_), .Y(men_men_n756_));
  INV        u734(.A(men_men_n189_), .Y(men_men_n757_));
  AOI220     u735(.A0(men_men_n757_), .A1(men_men_n750_), .B0(men_men_n756_), .B1(men_men_n68_), .Y(men_men_n758_));
  INV        u736(.A(men_men_n319_), .Y(men_men_n759_));
  NA2        u737(.A(men_men_n70_), .B(men_men_n125_), .Y(men_men_n760_));
  AOI210     u738(.A0(men_men_n118_), .A1(men_men_n760_), .B0(men_men_n759_), .Y(men_men_n761_));
  NO2        u739(.A(men_men_n497_), .B(men_men_n177_), .Y(men_men_n762_));
  INV        u740(.A(i_11_), .Y(men_men_n763_));
  NA3        u741(.A(men_men_n763_), .B(men_men_n455_), .C(men_men_n375_), .Y(men_men_n764_));
  NAi32      u742(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n765_));
  NO2        u743(.A(men_men_n689_), .B(men_men_n765_), .Y(men_men_n766_));
  OAI210     u744(.A0(men_men_n653_), .A1(men_men_n540_), .B0(men_men_n539_), .Y(men_men_n767_));
  NAi31      u745(.An(men_men_n766_), .B(men_men_n767_), .C(men_men_n764_), .Y(men_men_n768_));
  OR3        u746(.A(men_men_n768_), .B(men_men_n762_), .C(men_men_n761_), .Y(men_men_n769_));
  NA3        u747(.A(men_men_n338_), .B(men_men_n248_), .C(i_7_), .Y(men_men_n770_));
  OR2        u748(.A(men_men_n597_), .B(men_men_n434_), .Y(men_men_n771_));
  NA2        u749(.A(men_men_n771_), .B(men_men_n140_), .Y(men_men_n772_));
  OR2        u750(.A(men_men_n717_), .B(men_men_n36_), .Y(men_men_n773_));
  NA3        u751(.A(men_men_n773_), .B(men_men_n772_), .C(men_men_n770_), .Y(men_men_n774_));
  AOI220     u752(.A0(men_men_n979_), .A1(men_men_n539_), .B0(men_men_n749_), .B1(men_men_n684_), .Y(men_men_n775_));
  NA3        u753(.A(men_men_n362_), .B(men_men_n232_), .C(men_men_n140_), .Y(men_men_n776_));
  NA2        u754(.A(men_men_n382_), .B(men_men_n65_), .Y(men_men_n777_));
  NA4        u755(.A(men_men_n777_), .B(men_men_n776_), .C(men_men_n775_), .D(men_men_n580_), .Y(men_men_n778_));
  AO210      u756(.A0(men_men_n499_), .A1(men_men_n46_), .B0(men_men_n81_), .Y(men_men_n779_));
  NA3        u757(.A(men_men_n779_), .B(men_men_n465_), .C(men_men_n211_), .Y(men_men_n780_));
  AOI210     u758(.A0(men_men_n434_), .A1(men_men_n432_), .B0(men_men_n538_), .Y(men_men_n781_));
  NO2        u759(.A(men_men_n587_), .B(men_men_n96_), .Y(men_men_n782_));
  OAI210     u760(.A0(men_men_n782_), .A1(men_men_n106_), .B0(men_men_n396_), .Y(men_men_n783_));
  NA2        u761(.A(men_men_n237_), .B(men_men_n46_), .Y(men_men_n784_));
  INV        u762(.A(men_men_n563_), .Y(men_men_n785_));
  NA3        u763(.A(men_men_n785_), .B(men_men_n319_), .C(i_7_), .Y(men_men_n786_));
  NA4        u764(.A(men_men_n786_), .B(men_men_n783_), .C(men_men_n781_), .D(men_men_n780_), .Y(men_men_n787_));
  NO4        u765(.A(men_men_n787_), .B(men_men_n778_), .C(men_men_n774_), .D(men_men_n769_), .Y(men_men_n788_));
  NA4        u766(.A(men_men_n788_), .B(men_men_n758_), .C(men_men_n752_), .D(men_men_n365_), .Y(men3));
  NA2        u767(.A(i_12_), .B(i_10_), .Y(men_men_n790_));
  NA2        u768(.A(i_6_), .B(i_7_), .Y(men_men_n791_));
  NO2        u769(.A(men_men_n791_), .B(i_0_), .Y(men_men_n792_));
  NO2        u770(.A(i_11_), .B(men_men_n231_), .Y(men_men_n793_));
  NO3        u771(.A(men_men_n438_), .B(men_men_n83_), .C(men_men_n44_), .Y(men_men_n794_));
  AN2        u772(.A(men_men_n794_), .B(men_men_n166_), .Y(men_men_n795_));
  NA3        u773(.A(men_men_n776_), .B(men_men_n580_), .C(men_men_n361_), .Y(men_men_n796_));
  NA2        u774(.A(men_men_n796_), .B(men_men_n39_), .Y(men_men_n797_));
  NO3        u775(.A(men_men_n201_), .B(men_men_n442_), .C(men_men_n125_), .Y(men_men_n798_));
  NA2        u776(.A(men_men_n398_), .B(men_men_n45_), .Y(men_men_n799_));
  AN2        u777(.A(men_men_n440_), .B(men_men_n53_), .Y(men_men_n800_));
  NO2        u778(.A(men_men_n800_), .B(men_men_n798_), .Y(men_men_n801_));
  AOI210     u779(.A0(men_men_n801_), .A1(men_men_n797_), .B0(men_men_n48_), .Y(men_men_n802_));
  NA2        u780(.A(men_men_n984_), .B(men_men_n643_), .Y(men_men_n803_));
  NA2        u781(.A(men_men_n326_), .B(men_men_n424_), .Y(men_men_n804_));
  NO2        u782(.A(men_men_n804_), .B(men_men_n803_), .Y(men_men_n805_));
  NOi21      u783(.An(i_5_), .B(i_9_), .Y(men_men_n806_));
  NA2        u784(.A(men_men_n806_), .B(men_men_n431_), .Y(men_men_n807_));
  AOI210     u785(.A0(men_men_n260_), .A1(men_men_n457_), .B0(men_men_n658_), .Y(men_men_n808_));
  NO2        u786(.A(men_men_n808_), .B(men_men_n807_), .Y(men_men_n809_));
  NO4        u787(.A(men_men_n809_), .B(men_men_n805_), .C(men_men_n802_), .D(men_men_n795_), .Y(men_men_n810_));
  NA2        u788(.A(men_men_n177_), .B(men_men_n24_), .Y(men_men_n811_));
  INV        u789(.A(men_men_n641_), .Y(men_men_n812_));
  NO2        u790(.A(men_men_n812_), .B(men_men_n811_), .Y(men_men_n813_));
  NA2        u791(.A(men_men_n302_), .B(men_men_n123_), .Y(men_men_n814_));
  NAi21      u792(.An(men_men_n156_), .B(men_men_n424_), .Y(men_men_n815_));
  OAI220     u793(.A0(men_men_n815_), .A1(men_men_n784_), .B0(men_men_n814_), .B1(men_men_n388_), .Y(men_men_n816_));
  NO2        u794(.A(men_men_n816_), .B(men_men_n813_), .Y(men_men_n817_));
  NA2        u795(.A(men_men_n548_), .B(i_0_), .Y(men_men_n818_));
  NO3        u796(.A(men_men_n818_), .B(men_men_n370_), .C(men_men_n82_), .Y(men_men_n819_));
  NO4        u797(.A(men_men_n562_), .B(men_men_n208_), .C(men_men_n404_), .D(men_men_n397_), .Y(men_men_n820_));
  AOI210     u798(.A0(men_men_n820_), .A1(i_11_), .B0(men_men_n819_), .Y(men_men_n821_));
  NA2        u799(.A(men_men_n713_), .B(men_men_n320_), .Y(men_men_n822_));
  AOI210     u800(.A0(men_men_n465_), .A1(men_men_n82_), .B0(men_men_n55_), .Y(men_men_n823_));
  OAI220     u801(.A0(men_men_n823_), .A1(men_men_n822_), .B0(men_men_n628_), .B1(i_5_), .Y(men_men_n824_));
  NA2        u802(.A(i_0_), .B(i_10_), .Y(men_men_n825_));
  AOI220     u803(.A0(men_men_n326_), .A1(men_men_n92_), .B0(men_men_n177_), .B1(men_men_n78_), .Y(men_men_n826_));
  NA2        u804(.A(men_men_n543_), .B(i_4_), .Y(men_men_n827_));
  NA2        u805(.A(men_men_n180_), .B(men_men_n195_), .Y(men_men_n828_));
  OAI220     u806(.A0(men_men_n828_), .A1(men_men_n822_), .B0(men_men_n827_), .B1(men_men_n826_), .Y(men_men_n829_));
  NO2        u807(.A(men_men_n829_), .B(men_men_n824_), .Y(men_men_n830_));
  NA3        u808(.A(men_men_n830_), .B(men_men_n821_), .C(men_men_n817_), .Y(men_men_n831_));
  NO2        u809(.A(men_men_n97_), .B(men_men_n37_), .Y(men_men_n832_));
  NA2        u810(.A(i_11_), .B(i_9_), .Y(men_men_n833_));
  NO3        u811(.A(i_12_), .B(men_men_n833_), .C(men_men_n579_), .Y(men_men_n834_));
  AN2        u812(.A(men_men_n834_), .B(men_men_n832_), .Y(men_men_n835_));
  NA2        u813(.A(men_men_n379_), .B(men_men_n171_), .Y(men_men_n836_));
  NA2        u814(.A(men_men_n836_), .B(men_men_n154_), .Y(men_men_n837_));
  NO2        u815(.A(men_men_n833_), .B(men_men_n68_), .Y(men_men_n838_));
  NO2        u816(.A(men_men_n167_), .B(i_0_), .Y(men_men_n839_));
  AOI210     u817(.A0(men_men_n360_), .A1(men_men_n41_), .B0(men_men_n395_), .Y(men_men_n840_));
  NO2        u818(.A(men_men_n840_), .B(men_men_n807_), .Y(men_men_n841_));
  NO3        u819(.A(men_men_n841_), .B(men_men_n837_), .C(men_men_n835_), .Y(men_men_n842_));
  NA2        u820(.A(men_men_n627_), .B(men_men_n115_), .Y(men_men_n843_));
  NO2        u821(.A(i_6_), .B(men_men_n843_), .Y(men_men_n844_));
  AOI210     u822(.A0(men_men_n433_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n845_));
  NA2        u823(.A(men_men_n164_), .B(men_men_n97_), .Y(men_men_n846_));
  NOi32      u824(.An(men_men_n845_), .Bn(men_men_n180_), .C(men_men_n846_), .Y(men_men_n847_));
  NO2        u825(.A(men_men_n976_), .B(men_men_n799_), .Y(men_men_n848_));
  NO3        u826(.A(men_men_n848_), .B(men_men_n847_), .C(men_men_n844_), .Y(men_men_n849_));
  NOi21      u827(.An(i_7_), .B(i_5_), .Y(men_men_n850_));
  NOi31      u828(.An(men_men_n850_), .B(i_0_), .C(men_men_n694_), .Y(men_men_n851_));
  NA3        u829(.A(men_men_n851_), .B(men_men_n369_), .C(i_6_), .Y(men_men_n852_));
  OA210      u830(.A0(men_men_n846_), .A1(men_men_n497_), .B0(men_men_n852_), .Y(men_men_n853_));
  NO3        u831(.A(men_men_n391_), .B(men_men_n350_), .C(men_men_n346_), .Y(men_men_n854_));
  INV        u832(.A(men_men_n309_), .Y(men_men_n855_));
  NO2        u833(.A(men_men_n694_), .B(men_men_n250_), .Y(men_men_n856_));
  AOI210     u834(.A0(men_men_n856_), .A1(men_men_n855_), .B0(men_men_n854_), .Y(men_men_n857_));
  NA4        u835(.A(men_men_n857_), .B(men_men_n853_), .C(men_men_n849_), .D(men_men_n842_), .Y(men_men_n858_));
  AN2        u836(.A(men_men_n325_), .B(men_men_n320_), .Y(men_men_n859_));
  NO2        u837(.A(men_men_n790_), .B(men_men_n308_), .Y(men_men_n860_));
  BUFFER     u838(.A(men_men_n454_), .Y(men_men_n861_));
  NA2        u839(.A(men_men_n860_), .B(men_men_n838_), .Y(men_men_n862_));
  NO2        u840(.A(men_men_n815_), .B(i_6_), .Y(men_men_n863_));
  NA2        u841(.A(men_men_n838_), .B(men_men_n296_), .Y(men_men_n864_));
  NA2        u842(.A(men_men_n179_), .B(men_men_n864_), .Y(men_men_n865_));
  AOI220     u843(.A0(men_men_n865_), .A1(men_men_n455_), .B0(men_men_n863_), .B1(men_men_n68_), .Y(men_men_n866_));
  NO2        u844(.A(men_men_n70_), .B(men_men_n715_), .Y(men_men_n867_));
  INV        u845(.A(men_men_n867_), .Y(men_men_n868_));
  NO2        u846(.A(men_men_n868_), .B(men_men_n47_), .Y(men_men_n869_));
  NO3        u847(.A(men_men_n562_), .B(men_men_n345_), .C(men_men_n24_), .Y(men_men_n870_));
  INV        u848(.A(men_men_n870_), .Y(men_men_n871_));
  NAi21      u849(.An(i_9_), .B(i_5_), .Y(men_men_n872_));
  NO2        u850(.A(men_men_n872_), .B(men_men_n391_), .Y(men_men_n873_));
  NO2        u851(.A(men_men_n576_), .B(men_men_n99_), .Y(men_men_n874_));
  AOI220     u852(.A0(men_men_n874_), .A1(i_0_), .B0(men_men_n873_), .B1(men_men_n597_), .Y(men_men_n875_));
  OAI220     u853(.A0(men_men_n875_), .A1(men_men_n79_), .B0(men_men_n871_), .B1(men_men_n165_), .Y(men_men_n876_));
  NO3        u854(.A(men_men_n876_), .B(men_men_n869_), .C(men_men_n500_), .Y(men_men_n877_));
  NA3        u855(.A(men_men_n877_), .B(men_men_n866_), .C(men_men_n862_), .Y(men_men_n878_));
  NO3        u856(.A(men_men_n878_), .B(men_men_n858_), .C(men_men_n831_), .Y(men_men_n879_));
  NO2        u857(.A(i_0_), .B(men_men_n694_), .Y(men_men_n880_));
  NA2        u858(.A(men_men_n68_), .B(men_men_n44_), .Y(men_men_n881_));
  AN2        u859(.A(men_men_n880_), .B(men_men_n166_), .Y(men_men_n882_));
  NO2        u860(.A(men_men_n754_), .B(men_men_n846_), .Y(men_men_n883_));
  AOI210     u861(.A0(men_men_n882_), .A1(i_8_), .B0(men_men_n883_), .Y(men_men_n884_));
  NA2        u862(.A(men_men_n703_), .B(men_men_n139_), .Y(men_men_n885_));
  INV        u863(.A(men_men_n885_), .Y(men_men_n886_));
  NA2        u864(.A(men_men_n886_), .B(men_men_n643_), .Y(men_men_n887_));
  NO2        u865(.A(men_men_n767_), .B(men_men_n391_), .Y(men_men_n888_));
  NA3        u866(.A(men_men_n792_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n889_));
  NA2        u867(.A(men_men_n793_), .B(i_9_), .Y(men_men_n890_));
  AOI210     u868(.A0(men_men_n889_), .A1(men_men_n479_), .B0(men_men_n890_), .Y(men_men_n891_));
  OAI210     u869(.A0(men_men_n237_), .A1(i_9_), .B0(men_men_n224_), .Y(men_men_n892_));
  AOI210     u870(.A0(men_men_n892_), .A1(men_men_n818_), .B0(men_men_n147_), .Y(men_men_n893_));
  NO3        u871(.A(men_men_n893_), .B(men_men_n891_), .C(men_men_n888_), .Y(men_men_n894_));
  NA3        u872(.A(men_men_n894_), .B(men_men_n887_), .C(men_men_n884_), .Y(men_men_n895_));
  INV        u873(.A(men_men_n859_), .Y(men_men_n896_));
  AOI210     u874(.A0(men_men_n291_), .A1(men_men_n156_), .B0(men_men_n896_), .Y(men_men_n897_));
  NA3        u875(.A(men_men_n39_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n898_));
  NA2        u876(.A(i_5_), .B(men_men_n470_), .Y(men_men_n899_));
  AOI210     u877(.A0(men_men_n898_), .A1(men_men_n156_), .B0(men_men_n899_), .Y(men_men_n900_));
  NO2        u878(.A(men_men_n900_), .B(men_men_n897_), .Y(men_men_n901_));
  NO3        u879(.A(men_men_n825_), .B(men_men_n806_), .C(men_men_n182_), .Y(men_men_n902_));
  AOI220     u880(.A0(men_men_n902_), .A1(i_11_), .B0(men_men_n544_), .B1(men_men_n70_), .Y(men_men_n903_));
  NO3        u881(.A(men_men_n202_), .B(men_men_n368_), .C(i_0_), .Y(men_men_n904_));
  OAI210     u882(.A0(men_men_n904_), .A1(men_men_n71_), .B0(i_13_), .Y(men_men_n905_));
  OAI220     u883(.A0(men_men_n509_), .A1(men_men_n982_), .B0(i_12_), .B1(men_men_n591_), .Y(men_men_n906_));
  NA3        u884(.A(men_men_n906_), .B(men_men_n383_), .C(i_0_), .Y(men_men_n907_));
  NA4        u885(.A(men_men_n907_), .B(men_men_n905_), .C(men_men_n903_), .D(men_men_n901_), .Y(men_men_n908_));
  NO2        u886(.A(men_men_n236_), .B(men_men_n86_), .Y(men_men_n909_));
  AOI210     u887(.A0(men_men_n909_), .A1(men_men_n880_), .B0(men_men_n103_), .Y(men_men_n910_));
  AOI210     u888(.A0(men_men_n792_), .A1(men_men_n157_), .B0(men_men_n470_), .Y(men_men_n911_));
  NA2        u889(.A(men_men_n338_), .B(men_men_n168_), .Y(men_men_n912_));
  OA220      u890(.A0(men_men_n912_), .A1(men_men_n911_), .B0(men_men_n910_), .B1(i_5_), .Y(men_men_n913_));
  AOI210     u891(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n167_), .Y(men_men_n914_));
  NA2        u892(.A(men_men_n914_), .B(men_men_n861_), .Y(men_men_n915_));
  NA3        u893(.A(men_men_n475_), .B(men_men_n468_), .C(men_men_n452_), .Y(men_men_n916_));
  INV        u894(.A(men_men_n916_), .Y(men_men_n917_));
  NA3        u895(.A(men_men_n375_), .B(men_men_n164_), .C(men_men_n163_), .Y(men_men_n918_));
  NA3        u896(.A(men_men_n375_), .B(men_men_n327_), .C(men_men_n215_), .Y(men_men_n919_));
  INV        u897(.A(men_men_n919_), .Y(men_men_n920_));
  NOi31      u898(.An(men_men_n374_), .B(men_men_n881_), .C(men_men_n233_), .Y(men_men_n921_));
  NO3        u899(.A(men_men_n921_), .B(men_men_n920_), .C(men_men_n975_), .Y(men_men_n922_));
  NA4        u900(.A(men_men_n922_), .B(men_men_n917_), .C(men_men_n915_), .D(men_men_n913_), .Y(men_men_n923_));
  INV        u901(.A(i_5_), .Y(men_men_n924_));
  NA3        u902(.A(men_men_n793_), .B(men_men_n104_), .C(men_men_n118_), .Y(men_men_n925_));
  INV        u903(.A(men_men_n925_), .Y(men_men_n926_));
  NA2        u904(.A(men_men_n926_), .B(men_men_n924_), .Y(men_men_n927_));
  NO4        u905(.A(men_men_n233_), .B(men_men_n202_), .C(i_0_), .D(i_12_), .Y(men_men_n928_));
  AOI220     u906(.A0(men_men_n928_), .A1(i_10_), .B0(men_men_n748_), .B1(men_men_n168_), .Y(men_men_n929_));
  BUFFER     u907(.A(men_men_n825_), .Y(men_men_n930_));
  NO3        u908(.A(men_men_n930_), .B(i_12_), .C(men_men_n125_), .Y(men_men_n931_));
  NA2        u909(.A(men_men_n931_), .B(men_men_n211_), .Y(men_men_n932_));
  NA2        u910(.A(men_men_n850_), .B(men_men_n451_), .Y(men_men_n933_));
  OAI220     u911(.A0(i_7_), .A1(men_men_n983_), .B0(men_men_n933_), .B1(men_men_n644_), .Y(men_men_n934_));
  NA2        u912(.A(men_men_n934_), .B(men_men_n839_), .Y(men_men_n935_));
  NA4        u913(.A(men_men_n935_), .B(men_men_n932_), .C(men_men_n929_), .D(men_men_n927_), .Y(men_men_n936_));
  NO4        u914(.A(men_men_n936_), .B(men_men_n923_), .C(men_men_n908_), .D(men_men_n895_), .Y(men_men_n937_));
  NA3        u915(.A(men_men_n845_), .B(men_men_n357_), .C(i_5_), .Y(men_men_n938_));
  NA2        u916(.A(men_men_n938_), .B(men_men_n586_), .Y(men_men_n939_));
  NA2        u917(.A(men_men_n939_), .B(men_men_n200_), .Y(men_men_n940_));
  AN2        u918(.A(men_men_n669_), .B(men_men_n358_), .Y(men_men_n941_));
  NA2        u919(.A(men_men_n178_), .B(men_men_n180_), .Y(men_men_n942_));
  AO210      u920(.A0(men_men_n941_), .A1(men_men_n33_), .B0(men_men_n942_), .Y(men_men_n943_));
  OAI210     u921(.A0(men_men_n590_), .A1(men_men_n588_), .B0(men_men_n308_), .Y(men_men_n944_));
  NA2        u922(.A(men_men_n944_), .B(men_men_n943_), .Y(men_men_n945_));
  NO2        u923(.A(men_men_n445_), .B(men_men_n260_), .Y(men_men_n946_));
  NO2        u924(.A(men_men_n946_), .B(men_men_n820_), .Y(men_men_n947_));
  INV        u925(.A(men_men_n947_), .Y(men_men_n948_));
  AOI210     u926(.A0(men_men_n945_), .A1(men_men_n48_), .B0(men_men_n948_), .Y(men_men_n949_));
  AOI210     u927(.A0(men_men_n949_), .A1(men_men_n940_), .B0(men_men_n68_), .Y(men_men_n950_));
  INV        u928(.A(men_men_n71_), .Y(men_men_n951_));
  INV        u929(.A(men_men_n851_), .Y(men_men_n952_));
  AOI210     u930(.A0(men_men_n952_), .A1(men_men_n951_), .B0(men_men_n647_), .Y(men_men_n953_));
  NA2        u931(.A(i_8_), .B(men_men_n71_), .Y(men_men_n954_));
  NO2        u932(.A(men_men_n954_), .B(men_men_n231_), .Y(men_men_n955_));
  NO2        u933(.A(men_men_n955_), .B(men_men_n953_), .Y(men_men_n956_));
  OAI210     u934(.A0(men_men_n262_), .A1(men_men_n152_), .B0(men_men_n82_), .Y(men_men_n957_));
  NA3        u935(.A(men_men_n724_), .B(men_men_n282_), .C(men_men_n75_), .Y(men_men_n958_));
  AOI210     u936(.A0(men_men_n958_), .A1(men_men_n957_), .B0(i_11_), .Y(men_men_n959_));
  NA2        u937(.A(men_men_n581_), .B(men_men_n208_), .Y(men_men_n960_));
  OAI210     u938(.A0(men_men_n960_), .A1(men_men_n845_), .B0(men_men_n200_), .Y(men_men_n961_));
  NA2        u939(.A(men_men_n158_), .B(i_5_), .Y(men_men_n962_));
  AOI210     u940(.A0(men_men_n961_), .A1(men_men_n731_), .B0(men_men_n962_), .Y(men_men_n963_));
  NO4        u941(.A(men_men_n872_), .B(men_men_n458_), .C(men_men_n246_), .D(men_men_n245_), .Y(men_men_n964_));
  NO2        u942(.A(men_men_n964_), .B(men_men_n538_), .Y(men_men_n965_));
  INV        u943(.A(men_men_n351_), .Y(men_men_n966_));
  AOI210     u944(.A0(men_men_n966_), .A1(men_men_n965_), .B0(men_men_n40_), .Y(men_men_n967_));
  NO3        u945(.A(men_men_n967_), .B(men_men_n963_), .C(men_men_n959_), .Y(men_men_n968_));
  OAI210     u946(.A0(men_men_n956_), .A1(i_4_), .B0(men_men_n968_), .Y(men_men_n969_));
  NO3        u947(.A(men_men_n969_), .B(men_men_n541_), .C(men_men_n950_), .Y(men_men_n970_));
  NA4        u948(.A(men_men_n970_), .B(men_men_n937_), .C(men_men_n879_), .D(men_men_n810_), .Y(men4));
  INV        u949(.A(i_2_), .Y(men_men_n974_));
  INV        u950(.A(men_men_n918_), .Y(men_men_n975_));
  INV        u951(.A(men_men_n320_), .Y(men_men_n976_));
  INV        u952(.A(i_6_), .Y(men_men_n977_));
  INV        u953(.A(i_10_), .Y(men_men_n978_));
  INV        u954(.A(i_11_), .Y(men_men_n979_));
  INV        u955(.A(i_3_), .Y(men_men_n980_));
  INV        u956(.A(i_9_), .Y(men_men_n981_));
  INV        u957(.A(i_6_), .Y(men_men_n982_));
  INV        u958(.A(i_5_), .Y(men_men_n983_));
  INV        u959(.A(i_12_), .Y(men_men_n984_));
  INV        u960(.A(men_men_n201_), .Y(men_men_n985_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule