//Benchmark atmr_9sym_175_0.0625

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n152_, ori_ori_n153_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n150_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n153_, men_men_n154_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  INV        o002(.A(i_5_), .Y(ori_ori_n13_));
  NOi21      o003(.An(i_3_), .B(i_7_), .Y(ori_ori_n14_));
  NA3        o004(.A(ori_ori_n14_), .B(i_0_), .C(ori_ori_n13_), .Y(ori_ori_n15_));
  INV        o005(.A(i_0_), .Y(ori_ori_n16_));
  NOi21      o006(.An(i_1_), .B(i_3_), .Y(ori_ori_n17_));
  NA3        o007(.A(ori_ori_n17_), .B(ori_ori_n16_), .C(i_2_), .Y(ori_ori_n18_));
  AOI210     o008(.A0(ori_ori_n18_), .A1(ori_ori_n15_), .B0(ori_ori_n153_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA3        o012(.A(i_6_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  NA2        o014(.A(ori_ori_n24_), .B(i_5_), .Y(ori_ori_n25_));
  AOI210     o015(.A0(ori_ori_n25_), .A1(ori_ori_n23_), .B0(ori_ori_n21_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n27_));
  NA2        o017(.A(ori_ori_n16_), .B(i_5_), .Y(ori_ori_n28_));
  INV        o018(.A(i_2_), .Y(ori_ori_n29_));
  NOi21      o019(.An(i_6_), .B(i_8_), .Y(ori_ori_n30_));
  NOi21      o020(.An(i_7_), .B(i_1_), .Y(ori_ori_n31_));
  NOi21      o021(.An(i_5_), .B(i_6_), .Y(ori_ori_n32_));
  AOI220     o022(.A0(ori_ori_n32_), .A1(ori_ori_n31_), .B0(ori_ori_n30_), .B1(i_5_), .Y(ori_ori_n33_));
  NO3        o023(.A(ori_ori_n33_), .B(ori_ori_n29_), .C(i_4_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_0_), .B(i_4_), .Y(ori_ori_n35_));
  INV        o025(.A(i_1_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_3_), .B(i_0_), .Y(ori_ori_n37_));
  NA2        o027(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o028(.A(ori_ori_n23_), .B(ori_ori_n38_), .Y(ori_ori_n39_));
  NO2        o029(.A(ori_ori_n39_), .B(ori_ori_n34_), .Y(ori_ori_n40_));
  NOi21      o030(.An(i_4_), .B(i_0_), .Y(ori_ori_n41_));
  NO2        o031(.A(ori_ori_n24_), .B(ori_ori_n14_), .Y(ori_ori_n42_));
  NA2        o032(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n43_));
  NOi21      o033(.An(i_2_), .B(i_8_), .Y(ori_ori_n44_));
  NO2        o034(.A(ori_ori_n41_), .B(ori_ori_n35_), .Y(ori_ori_n45_));
  NO3        o035(.A(ori_ori_n45_), .B(ori_ori_n43_), .C(ori_ori_n42_), .Y(ori_ori_n46_));
  INV        o036(.A(ori_ori_n46_), .Y(ori_ori_n47_));
  NOi31      o037(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n48_));
  NA2        o038(.A(ori_ori_n48_), .B(i_0_), .Y(ori_ori_n49_));
  NOi21      o039(.An(i_4_), .B(i_3_), .Y(ori_ori_n50_));
  NOi21      o040(.An(i_1_), .B(i_4_), .Y(ori_ori_n51_));
  OAI210     o041(.A0(ori_ori_n51_), .A1(ori_ori_n50_), .B0(ori_ori_n44_), .Y(ori_ori_n52_));
  NA2        o042(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  AN2        o043(.A(i_8_), .B(i_7_), .Y(ori_ori_n54_));
  INV        o044(.A(ori_ori_n54_), .Y(ori_ori_n55_));
  NOi21      o045(.An(i_8_), .B(i_7_), .Y(ori_ori_n56_));
  NA3        o046(.A(ori_ori_n56_), .B(ori_ori_n50_), .C(i_6_), .Y(ori_ori_n57_));
  OAI210     o047(.A0(ori_ori_n55_), .A1(ori_ori_n43_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  AOI220     o048(.A0(ori_ori_n58_), .A1(ori_ori_n29_), .B0(ori_ori_n53_), .B1(ori_ori_n32_), .Y(ori_ori_n59_));
  NA4        o049(.A(ori_ori_n59_), .B(ori_ori_n47_), .C(ori_ori_n40_), .D(ori_ori_n27_), .Y(ori_ori_n60_));
  NA2        o050(.A(i_8_), .B(i_7_), .Y(ori_ori_n61_));
  NO3        o051(.A(ori_ori_n61_), .B(ori_ori_n153_), .C(i_1_), .Y(ori_ori_n62_));
  NA2        o052(.A(i_8_), .B(ori_ori_n22_), .Y(ori_ori_n63_));
  NOi21      o053(.An(i_1_), .B(i_2_), .Y(ori_ori_n64_));
  NO2        o054(.A(ori_ori_n152_), .B(ori_ori_n63_), .Y(ori_ori_n65_));
  OAI210     o055(.A0(ori_ori_n65_), .A1(ori_ori_n62_), .B0(ori_ori_n13_), .Y(ori_ori_n66_));
  NA3        o056(.A(ori_ori_n56_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n67_));
  INV        o057(.A(ori_ori_n67_), .Y(ori_ori_n68_));
  NA2        o058(.A(ori_ori_n17_), .B(i_6_), .Y(ori_ori_n69_));
  INV        o059(.A(ori_ori_n69_), .Y(ori_ori_n70_));
  INV        o060(.A(i_0_), .Y(ori_ori_n71_));
  AOI220     o061(.A0(ori_ori_n71_), .A1(ori_ori_n70_), .B0(ori_ori_n68_), .B1(ori_ori_n50_), .Y(ori_ori_n72_));
  NA2        o062(.A(ori_ori_n72_), .B(ori_ori_n66_), .Y(ori_ori_n73_));
  NOi21      o063(.An(i_7_), .B(i_8_), .Y(ori_ori_n74_));
  NOi21      o064(.An(i_6_), .B(i_5_), .Y(ori_ori_n75_));
  NA2        o065(.A(ori_ori_n75_), .B(ori_ori_n64_), .Y(ori_ori_n76_));
  NA3        o066(.A(ori_ori_n24_), .B(i_2_), .C(ori_ori_n13_), .Y(ori_ori_n77_));
  NO2        o067(.A(i_3_), .B(ori_ori_n77_), .Y(ori_ori_n78_));
  AOI220     o068(.A0(ori_ori_n37_), .A1(ori_ori_n36_), .B0(ori_ori_n17_), .B1(ori_ori_n29_), .Y(ori_ori_n79_));
  NA2        o069(.A(ori_ori_n20_), .B(i_7_), .Y(ori_ori_n80_));
  NO2        o070(.A(ori_ori_n80_), .B(ori_ori_n79_), .Y(ori_ori_n81_));
  NO2        o071(.A(ori_ori_n81_), .B(ori_ori_n78_), .Y(ori_ori_n82_));
  NA3        o072(.A(ori_ori_n56_), .B(ori_ori_n29_), .C(i_3_), .Y(ori_ori_n83_));
  NA2        o073(.A(ori_ori_n36_), .B(i_6_), .Y(ori_ori_n84_));
  AOI210     o074(.A0(ori_ori_n84_), .A1(ori_ori_n21_), .B0(ori_ori_n83_), .Y(ori_ori_n85_));
  NOi21      o075(.An(i_2_), .B(i_1_), .Y(ori_ori_n86_));
  AN3        o076(.A(ori_ori_n74_), .B(ori_ori_n86_), .C(ori_ori_n41_), .Y(ori_ori_n87_));
  NAi21      o077(.An(i_6_), .B(i_0_), .Y(ori_ori_n88_));
  NA3        o078(.A(ori_ori_n51_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n89_));
  NOi21      o079(.An(i_4_), .B(i_6_), .Y(ori_ori_n90_));
  NA3        o080(.A(i_5_), .B(ori_ori_n64_), .C(ori_ori_n90_), .Y(ori_ori_n91_));
  OAI210     o081(.A0(ori_ori_n89_), .A1(ori_ori_n88_), .B0(ori_ori_n91_), .Y(ori_ori_n92_));
  NA2        o082(.A(ori_ori_n64_), .B(ori_ori_n30_), .Y(ori_ori_n93_));
  NO3        o083(.A(ori_ori_n92_), .B(ori_ori_n87_), .C(ori_ori_n85_), .Y(ori_ori_n94_));
  NA2        o084(.A(ori_ori_n56_), .B(ori_ori_n12_), .Y(ori_ori_n95_));
  NA2        o085(.A(ori_ori_n30_), .B(ori_ori_n13_), .Y(ori_ori_n96_));
  NOi21      o086(.An(i_3_), .B(i_1_), .Y(ori_ori_n97_));
  NA2        o087(.A(ori_ori_n97_), .B(i_4_), .Y(ori_ori_n98_));
  AOI210     o088(.A0(ori_ori_n96_), .A1(ori_ori_n95_), .B0(ori_ori_n98_), .Y(ori_ori_n99_));
  INV        o089(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NA4        o090(.A(ori_ori_n100_), .B(ori_ori_n94_), .C(ori_ori_n82_), .D(ori_ori_n76_), .Y(ori_ori_n101_));
  NA2        o091(.A(ori_ori_n44_), .B(ori_ori_n14_), .Y(ori_ori_n102_));
  NOi31      o092(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n103_));
  NOi31      o093(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n104_));
  OAI210     o094(.A0(ori_ori_n104_), .A1(ori_ori_n103_), .B0(i_7_), .Y(ori_ori_n105_));
  NA3        o095(.A(ori_ori_n30_), .B(i_2_), .C(ori_ori_n13_), .Y(ori_ori_n106_));
  NA3        o096(.A(ori_ori_n106_), .B(ori_ori_n105_), .C(ori_ori_n93_), .Y(ori_ori_n107_));
  NA2        o097(.A(ori_ori_n107_), .B(ori_ori_n35_), .Y(ori_ori_n108_));
  NA2        o098(.A(ori_ori_n50_), .B(ori_ori_n31_), .Y(ori_ori_n109_));
  AOI210     o099(.A0(ori_ori_n109_), .A1(ori_ori_n67_), .B0(ori_ori_n28_), .Y(ori_ori_n110_));
  NA4        o100(.A(ori_ori_n54_), .B(ori_ori_n86_), .C(ori_ori_n16_), .D(ori_ori_n12_), .Y(ori_ori_n111_));
  NAi31      o101(.An(ori_ori_n88_), .B(ori_ori_n74_), .C(ori_ori_n86_), .Y(ori_ori_n112_));
  NA3        o102(.A(ori_ori_n56_), .B(ori_ori_n48_), .C(i_6_), .Y(ori_ori_n113_));
  NA3        o103(.A(ori_ori_n113_), .B(ori_ori_n112_), .C(ori_ori_n111_), .Y(ori_ori_n114_));
  NOi21      o104(.An(i_0_), .B(i_2_), .Y(ori_ori_n115_));
  NA3        o105(.A(ori_ori_n115_), .B(ori_ori_n31_), .C(ori_ori_n90_), .Y(ori_ori_n116_));
  NOi32      o106(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n117_));
  NA2        o107(.A(ori_ori_n117_), .B(ori_ori_n103_), .Y(ori_ori_n118_));
  NA3        o108(.A(ori_ori_n115_), .B(ori_ori_n50_), .C(ori_ori_n30_), .Y(ori_ori_n119_));
  NA3        o109(.A(ori_ori_n119_), .B(ori_ori_n118_), .C(ori_ori_n116_), .Y(ori_ori_n120_));
  NA4        o110(.A(ori_ori_n48_), .B(i_6_), .C(ori_ori_n13_), .D(i_7_), .Y(ori_ori_n121_));
  NA4        o111(.A(ori_ori_n51_), .B(ori_ori_n32_), .C(ori_ori_n16_), .D(i_8_), .Y(ori_ori_n122_));
  NA2        o112(.A(ori_ori_n51_), .B(ori_ori_n37_), .Y(ori_ori_n123_));
  NA3        o113(.A(ori_ori_n123_), .B(ori_ori_n122_), .C(ori_ori_n121_), .Y(ori_ori_n124_));
  NO4        o114(.A(ori_ori_n124_), .B(ori_ori_n120_), .C(ori_ori_n114_), .D(ori_ori_n110_), .Y(ori_ori_n125_));
  NOi21      o115(.An(i_5_), .B(i_2_), .Y(ori_ori_n126_));
  NA2        o116(.A(ori_ori_n126_), .B(ori_ori_n74_), .Y(ori_ori_n127_));
  AOI210     o117(.A0(ori_ori_n127_), .A1(ori_ori_n102_), .B0(ori_ori_n84_), .Y(ori_ori_n128_));
  NO3        o118(.A(ori_ori_n20_), .B(ori_ori_n11_), .C(ori_ori_n13_), .Y(ori_ori_n129_));
  NA2        o119(.A(i_2_), .B(i_4_), .Y(ori_ori_n130_));
  INV        o120(.A(ori_ori_n130_), .Y(ori_ori_n131_));
  NO2        o121(.A(i_8_), .B(i_7_), .Y(ori_ori_n132_));
  OA210      o122(.A0(ori_ori_n131_), .A1(ori_ori_n129_), .B0(ori_ori_n132_), .Y(ori_ori_n133_));
  NA2        o123(.A(ori_ori_n97_), .B(i_0_), .Y(ori_ori_n134_));
  NO2        o124(.A(ori_ori_n134_), .B(i_4_), .Y(ori_ori_n135_));
  NO3        o125(.A(ori_ori_n135_), .B(ori_ori_n133_), .C(ori_ori_n128_), .Y(ori_ori_n136_));
  NA2        o126(.A(ori_ori_n74_), .B(ori_ori_n12_), .Y(ori_ori_n137_));
  NA2        o127(.A(i_1_), .B(ori_ori_n13_), .Y(ori_ori_n138_));
  NA2        o128(.A(ori_ori_n41_), .B(i_3_), .Y(ori_ori_n139_));
  AOI210     o129(.A0(ori_ori_n139_), .A1(ori_ori_n138_), .B0(ori_ori_n137_), .Y(ori_ori_n140_));
  NA3        o130(.A(ori_ori_n115_), .B(ori_ori_n56_), .C(ori_ori_n90_), .Y(ori_ori_n141_));
  OAI210     o131(.A0(ori_ori_n83_), .A1(ori_ori_n28_), .B0(ori_ori_n141_), .Y(ori_ori_n142_));
  NA4        o132(.A(i_5_), .B(ori_ori_n54_), .C(ori_ori_n36_), .D(ori_ori_n20_), .Y(ori_ori_n143_));
  NOi31      o133(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n144_));
  NA2        o134(.A(ori_ori_n117_), .B(ori_ori_n144_), .Y(ori_ori_n145_));
  NA2        o135(.A(ori_ori_n145_), .B(ori_ori_n143_), .Y(ori_ori_n146_));
  NO3        o136(.A(ori_ori_n146_), .B(ori_ori_n142_), .C(ori_ori_n140_), .Y(ori_ori_n147_));
  NA4        o137(.A(ori_ori_n147_), .B(ori_ori_n136_), .C(ori_ori_n125_), .D(ori_ori_n108_), .Y(ori_ori_n148_));
  OR4        o138(.A(ori_ori_n148_), .B(ori_ori_n101_), .C(ori_ori_n73_), .D(ori_ori_n60_), .Y(ori00));
  INV        o139(.A(i_2_), .Y(ori_ori_n152_));
  INV        o140(.A(i_4_), .Y(ori_ori_n153_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  INV        m002(.A(i_5_), .Y(mai_mai_n13_));
  NOi21      m003(.An(i_3_), .B(i_7_), .Y(mai_mai_n14_));
  INV        m004(.A(i_0_), .Y(mai_mai_n15_));
  NOi21      m005(.An(i_1_), .B(i_3_), .Y(mai_mai_n16_));
  INV        m006(.A(i_4_), .Y(mai_mai_n17_));
  NA2        m007(.A(i_0_), .B(mai_mai_n17_), .Y(mai_mai_n18_));
  INV        m008(.A(i_7_), .Y(mai_mai_n19_));
  NA3        m009(.A(i_6_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n20_));
  NOi21      m010(.An(i_8_), .B(i_6_), .Y(mai_mai_n21_));
  NOi21      m011(.An(i_1_), .B(i_8_), .Y(mai_mai_n22_));
  AOI220     m012(.A0(mai_mai_n22_), .A1(i_2_), .B0(mai_mai_n21_), .B1(i_5_), .Y(mai_mai_n23_));
  AOI210     m013(.A0(mai_mai_n23_), .A1(mai_mai_n20_), .B0(mai_mai_n18_), .Y(mai_mai_n24_));
  NA2        m014(.A(mai_mai_n24_), .B(mai_mai_n11_), .Y(mai_mai_n25_));
  NA2        m015(.A(mai_mai_n15_), .B(i_5_), .Y(mai_mai_n26_));
  NO2        m016(.A(i_2_), .B(i_4_), .Y(mai_mai_n27_));
  NA3        m017(.A(mai_mai_n27_), .B(i_6_), .C(i_8_), .Y(mai_mai_n28_));
  INV        m018(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  INV        m019(.A(i_2_), .Y(mai_mai_n30_));
  NOi21      m020(.An(i_5_), .B(i_0_), .Y(mai_mai_n31_));
  NOi21      m021(.An(i_6_), .B(i_8_), .Y(mai_mai_n32_));
  NOi21      m022(.An(i_7_), .B(i_1_), .Y(mai_mai_n33_));
  NOi21      m023(.An(i_5_), .B(i_6_), .Y(mai_mai_n34_));
  AOI220     m024(.A0(mai_mai_n34_), .A1(mai_mai_n33_), .B0(mai_mai_n32_), .B1(mai_mai_n31_), .Y(mai_mai_n35_));
  NO3        m025(.A(mai_mai_n35_), .B(mai_mai_n30_), .C(i_4_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_0_), .B(i_4_), .Y(mai_mai_n37_));
  XO2        m027(.A(i_1_), .B(i_3_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_7_), .B(i_5_), .Y(mai_mai_n39_));
  AN3        m029(.A(mai_mai_n39_), .B(mai_mai_n38_), .C(mai_mai_n37_), .Y(mai_mai_n40_));
  INV        m030(.A(i_1_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_3_), .B(i_0_), .Y(mai_mai_n42_));
  NA2        m032(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA3        m033(.A(i_6_), .B(mai_mai_n13_), .C(i_7_), .Y(mai_mai_n44_));
  AOI210     m034(.A0(mai_mai_n44_), .A1(mai_mai_n20_), .B0(mai_mai_n43_), .Y(mai_mai_n45_));
  NO4        m035(.A(mai_mai_n45_), .B(mai_mai_n40_), .C(mai_mai_n36_), .D(mai_mai_n29_), .Y(mai_mai_n46_));
  INV        m036(.A(i_8_), .Y(mai_mai_n47_));
  NA2        m037(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n48_));
  NO3        m038(.A(mai_mai_n48_), .B(i_2_), .C(mai_mai_n47_), .Y(mai_mai_n49_));
  NOi21      m039(.An(i_4_), .B(i_0_), .Y(mai_mai_n50_));
  AOI210     m040(.A0(mai_mai_n50_), .A1(mai_mai_n21_), .B0(mai_mai_n14_), .Y(mai_mai_n51_));
  NA2        m041(.A(i_1_), .B(mai_mai_n13_), .Y(mai_mai_n52_));
  NOi21      m042(.An(i_2_), .B(i_8_), .Y(mai_mai_n53_));
  NO3        m043(.A(mai_mai_n53_), .B(mai_mai_n50_), .C(mai_mai_n37_), .Y(mai_mai_n54_));
  NO3        m044(.A(mai_mai_n54_), .B(mai_mai_n52_), .C(mai_mai_n51_), .Y(mai_mai_n55_));
  NO2        m045(.A(mai_mai_n55_), .B(mai_mai_n49_), .Y(mai_mai_n56_));
  NOi31      m046(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n57_));
  NA2        m047(.A(mai_mai_n57_), .B(i_0_), .Y(mai_mai_n58_));
  NOi21      m048(.An(i_4_), .B(i_3_), .Y(mai_mai_n59_));
  NOi21      m049(.An(i_1_), .B(i_4_), .Y(mai_mai_n60_));
  OAI210     m050(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n53_), .Y(mai_mai_n61_));
  NA2        m051(.A(mai_mai_n61_), .B(mai_mai_n58_), .Y(mai_mai_n62_));
  NA2        m052(.A(i_8_), .B(mai_mai_n12_), .Y(mai_mai_n63_));
  NOi21      m053(.An(i_8_), .B(i_7_), .Y(mai_mai_n64_));
  NO2        m054(.A(mai_mai_n63_), .B(mai_mai_n52_), .Y(mai_mai_n65_));
  AOI220     m055(.A0(mai_mai_n65_), .A1(mai_mai_n30_), .B0(mai_mai_n62_), .B1(mai_mai_n34_), .Y(mai_mai_n66_));
  NA4        m056(.A(mai_mai_n66_), .B(mai_mai_n56_), .C(mai_mai_n46_), .D(mai_mai_n25_), .Y(mai_mai_n67_));
  NA2        m057(.A(i_8_), .B(i_7_), .Y(mai_mai_n68_));
  NO3        m058(.A(mai_mai_n68_), .B(i_6_), .C(i_1_), .Y(mai_mai_n69_));
  NA2        m059(.A(i_8_), .B(mai_mai_n19_), .Y(mai_mai_n70_));
  AOI220     m060(.A0(mai_mai_n42_), .A1(i_1_), .B0(mai_mai_n38_), .B1(i_2_), .Y(mai_mai_n71_));
  NOi21      m061(.An(i_1_), .B(i_2_), .Y(mai_mai_n72_));
  NO2        m062(.A(mai_mai_n71_), .B(mai_mai_n70_), .Y(mai_mai_n73_));
  OAI210     m063(.A0(mai_mai_n73_), .A1(mai_mai_n69_), .B0(mai_mai_n13_), .Y(mai_mai_n74_));
  NA3        m064(.A(mai_mai_n64_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n75_));
  NA3        m065(.A(mai_mai_n16_), .B(i_2_), .C(i_6_), .Y(mai_mai_n76_));
  INV        m066(.A(mai_mai_n76_), .Y(mai_mai_n77_));
  NO2        m067(.A(i_0_), .B(i_4_), .Y(mai_mai_n78_));
  AOI220     m068(.A0(mai_mai_n78_), .A1(mai_mai_n77_), .B0(mai_mai_n22_), .B1(mai_mai_n59_), .Y(mai_mai_n79_));
  NA2        m069(.A(mai_mai_n79_), .B(mai_mai_n74_), .Y(mai_mai_n80_));
  NA2        m070(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n81_));
  NOi21      m071(.An(i_7_), .B(i_8_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n82_), .B(mai_mai_n12_), .Y(mai_mai_n83_));
  OAI210     m073(.A0(mai_mai_n83_), .A1(mai_mai_n11_), .B0(mai_mai_n81_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n84_), .B(mai_mai_n72_), .Y(mai_mai_n85_));
  NA3        m075(.A(mai_mai_n21_), .B(i_2_), .C(mai_mai_n13_), .Y(mai_mai_n86_));
  AOI210     m076(.A0(mai_mai_n18_), .A1(mai_mai_n48_), .B0(mai_mai_n86_), .Y(mai_mai_n87_));
  AOI220     m077(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n16_), .B1(mai_mai_n30_), .Y(mai_mai_n88_));
  NA3        m078(.A(mai_mai_n17_), .B(i_5_), .C(i_7_), .Y(mai_mai_n89_));
  NA2        m079(.A(i_4_), .B(i_5_), .Y(mai_mai_n90_));
  NA3        m080(.A(mai_mai_n68_), .B(mai_mai_n16_), .C(mai_mai_n15_), .Y(mai_mai_n91_));
  OAI220     m081(.A0(mai_mai_n91_), .A1(mai_mai_n90_), .B0(mai_mai_n89_), .B1(mai_mai_n88_), .Y(mai_mai_n92_));
  NO2        m082(.A(mai_mai_n92_), .B(mai_mai_n87_), .Y(mai_mai_n93_));
  NA2        m083(.A(mai_mai_n41_), .B(i_6_), .Y(mai_mai_n94_));
  NAi21      m084(.An(i_6_), .B(i_0_), .Y(mai_mai_n95_));
  NA3        m085(.A(mai_mai_n60_), .B(i_5_), .C(mai_mai_n19_), .Y(mai_mai_n96_));
  NOi21      m086(.An(i_4_), .B(i_6_), .Y(mai_mai_n97_));
  NO2        m087(.A(mai_mai_n96_), .B(mai_mai_n95_), .Y(mai_mai_n98_));
  NA2        m088(.A(mai_mai_n72_), .B(mai_mai_n32_), .Y(mai_mai_n99_));
  NOi21      m089(.An(mai_mai_n39_), .B(mai_mai_n99_), .Y(mai_mai_n100_));
  NO2        m090(.A(mai_mai_n100_), .B(mai_mai_n98_), .Y(mai_mai_n101_));
  NOi31      m091(.An(mai_mai_n50_), .B(mai_mai_n150_), .C(i_2_), .Y(mai_mai_n102_));
  NOi21      m092(.An(i_3_), .B(i_1_), .Y(mai_mai_n103_));
  NA2        m093(.A(mai_mai_n103_), .B(i_4_), .Y(mai_mai_n104_));
  NO2        m094(.A(i_8_), .B(mai_mai_n104_), .Y(mai_mai_n105_));
  NA2        m095(.A(mai_mai_n82_), .B(mai_mai_n13_), .Y(mai_mai_n106_));
  NOi31      m096(.An(mai_mai_n42_), .B(mai_mai_n106_), .C(mai_mai_n30_), .Y(mai_mai_n107_));
  NO3        m097(.A(mai_mai_n107_), .B(mai_mai_n105_), .C(mai_mai_n102_), .Y(mai_mai_n108_));
  NA4        m098(.A(mai_mai_n108_), .B(mai_mai_n101_), .C(mai_mai_n93_), .D(mai_mai_n85_), .Y(mai_mai_n109_));
  NA2        m099(.A(mai_mai_n53_), .B(mai_mai_n14_), .Y(mai_mai_n110_));
  NOi31      m100(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n111_));
  NA2        m101(.A(mai_mai_n111_), .B(i_7_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n32_), .B(mai_mai_n13_), .Y(mai_mai_n113_));
  NA4        m103(.A(mai_mai_n113_), .B(mai_mai_n112_), .C(mai_mai_n110_), .D(mai_mai_n99_), .Y(mai_mai_n114_));
  NA2        m104(.A(mai_mai_n114_), .B(mai_mai_n37_), .Y(mai_mai_n115_));
  NA2        m105(.A(mai_mai_n59_), .B(mai_mai_n33_), .Y(mai_mai_n116_));
  AOI210     m106(.A0(mai_mai_n116_), .A1(mai_mai_n75_), .B0(mai_mai_n26_), .Y(mai_mai_n117_));
  NA3        m107(.A(mai_mai_n64_), .B(mai_mai_n57_), .C(i_6_), .Y(mai_mai_n118_));
  INV        m108(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  NA2        m109(.A(mai_mai_n59_), .B(mai_mai_n32_), .Y(mai_mai_n120_));
  INV        m110(.A(mai_mai_n120_), .Y(mai_mai_n121_));
  NA4        m111(.A(mai_mai_n57_), .B(i_6_), .C(mai_mai_n13_), .D(i_7_), .Y(mai_mai_n122_));
  NA4        m112(.A(mai_mai_n60_), .B(mai_mai_n34_), .C(mai_mai_n15_), .D(i_8_), .Y(mai_mai_n123_));
  NA4        m113(.A(mai_mai_n60_), .B(mai_mai_n42_), .C(i_5_), .D(mai_mai_n19_), .Y(mai_mai_n124_));
  NA3        m114(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n122_), .Y(mai_mai_n125_));
  NO4        m115(.A(mai_mai_n125_), .B(mai_mai_n121_), .C(mai_mai_n119_), .D(mai_mai_n117_), .Y(mai_mai_n126_));
  BUFFER     m116(.A(i_5_), .Y(mai_mai_n127_));
  NA2        m117(.A(mai_mai_n127_), .B(mai_mai_n82_), .Y(mai_mai_n128_));
  AOI210     m118(.A0(mai_mai_n128_), .A1(mai_mai_n110_), .B0(mai_mai_n94_), .Y(mai_mai_n129_));
  NO3        m119(.A(i_2_), .B(mai_mai_n17_), .C(mai_mai_n11_), .Y(mai_mai_n130_));
  NO2        m120(.A(i_8_), .B(i_7_), .Y(mai_mai_n131_));
  AN2        m121(.A(mai_mai_n130_), .B(mai_mai_n131_), .Y(mai_mai_n132_));
  NA4        m122(.A(mai_mai_n103_), .B(i_0_), .C(i_5_), .D(mai_mai_n19_), .Y(mai_mai_n133_));
  NO2        m123(.A(mai_mai_n133_), .B(i_4_), .Y(mai_mai_n134_));
  NO3        m124(.A(mai_mai_n134_), .B(mai_mai_n132_), .C(mai_mai_n129_), .Y(mai_mai_n135_));
  NA2        m125(.A(mai_mai_n82_), .B(mai_mai_n12_), .Y(mai_mai_n136_));
  NA2        m126(.A(i_2_), .B(mai_mai_n13_), .Y(mai_mai_n137_));
  NO2        m127(.A(mai_mai_n137_), .B(mai_mai_n136_), .Y(mai_mai_n138_));
  NA2        m128(.A(mai_mai_n64_), .B(mai_mai_n97_), .Y(mai_mai_n139_));
  INV        m129(.A(mai_mai_n139_), .Y(mai_mai_n140_));
  NA3        m130(.A(mai_mai_n53_), .B(mai_mai_n31_), .C(mai_mai_n14_), .Y(mai_mai_n141_));
  NOi31      m131(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n142_));
  NA2        m132(.A(i_4_), .B(mai_mai_n142_), .Y(mai_mai_n143_));
  NA2        m133(.A(mai_mai_n143_), .B(mai_mai_n141_), .Y(mai_mai_n144_));
  NO3        m134(.A(mai_mai_n144_), .B(mai_mai_n140_), .C(mai_mai_n138_), .Y(mai_mai_n145_));
  NA4        m135(.A(mai_mai_n145_), .B(mai_mai_n135_), .C(mai_mai_n126_), .D(mai_mai_n115_), .Y(mai_mai_n146_));
  OR4        m136(.A(mai_mai_n146_), .B(mai_mai_n109_), .C(mai_mai_n80_), .D(mai_mai_n67_), .Y(mai00));
  INV        m137(.A(i_8_), .Y(mai_mai_n150_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NO2        u013(.A(men_men_n153_), .B(men_men_n22_), .Y(men_men_n24_));
  AOI210     u014(.A0(men_men_n24_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n25_));
  NA2        u015(.A(i_0_), .B(men_men_n14_), .Y(men_men_n26_));
  NA2        u016(.A(men_men_n17_), .B(i_5_), .Y(men_men_n27_));
  NO2        u017(.A(i_2_), .B(i_4_), .Y(men_men_n28_));
  NA3        u018(.A(men_men_n28_), .B(i_6_), .C(i_8_), .Y(men_men_n29_));
  AOI210     u019(.A0(men_men_n27_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n30_));
  INV        u020(.A(i_2_), .Y(men_men_n31_));
  NOi21      u021(.An(i_6_), .B(i_8_), .Y(men_men_n32_));
  NOi21      u022(.An(i_7_), .B(i_1_), .Y(men_men_n33_));
  NOi21      u023(.An(i_5_), .B(i_6_), .Y(men_men_n34_));
  NOi21      u024(.An(i_0_), .B(i_4_), .Y(men_men_n35_));
  XO2        u025(.A(i_1_), .B(i_3_), .Y(men_men_n36_));
  NOi21      u026(.An(i_7_), .B(i_5_), .Y(men_men_n37_));
  AN3        u027(.A(men_men_n37_), .B(men_men_n36_), .C(men_men_n35_), .Y(men_men_n38_));
  INV        u028(.A(i_1_), .Y(men_men_n39_));
  NOi21      u029(.An(i_3_), .B(i_0_), .Y(men_men_n40_));
  NA2        u030(.A(men_men_n40_), .B(men_men_n39_), .Y(men_men_n41_));
  NA3        u031(.A(i_6_), .B(men_men_n14_), .C(i_7_), .Y(men_men_n42_));
  AOI210     u032(.A0(men_men_n42_), .A1(men_men_n154_), .B0(men_men_n41_), .Y(men_men_n43_));
  NO3        u033(.A(men_men_n43_), .B(men_men_n38_), .C(men_men_n30_), .Y(men_men_n44_));
  INV        u034(.A(i_8_), .Y(men_men_n45_));
  NOi21      u035(.An(i_4_), .B(i_0_), .Y(men_men_n46_));
  INV        u036(.A(men_men_n15_), .Y(men_men_n47_));
  NA2        u037(.A(i_1_), .B(men_men_n14_), .Y(men_men_n48_));
  NO2        u038(.A(men_men_n46_), .B(men_men_n35_), .Y(men_men_n49_));
  NO3        u039(.A(men_men_n49_), .B(men_men_n48_), .C(men_men_n47_), .Y(men_men_n50_));
  INV        u040(.A(men_men_n50_), .Y(men_men_n51_));
  NOi31      u041(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n52_));
  NOi21      u042(.An(i_4_), .B(i_3_), .Y(men_men_n53_));
  AN2        u043(.A(i_8_), .B(i_7_), .Y(men_men_n54_));
  NA2        u044(.A(men_men_n54_), .B(men_men_n12_), .Y(men_men_n55_));
  NOi21      u045(.An(i_8_), .B(i_7_), .Y(men_men_n56_));
  NA3        u046(.A(men_men_n56_), .B(men_men_n53_), .C(i_6_), .Y(men_men_n57_));
  OAI210     u047(.A0(men_men_n55_), .A1(men_men_n48_), .B0(men_men_n57_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(men_men_n31_), .Y(men_men_n59_));
  NA4        u049(.A(men_men_n59_), .B(men_men_n51_), .C(men_men_n44_), .D(men_men_n25_), .Y(men_men_n60_));
  NA2        u050(.A(i_8_), .B(i_7_), .Y(men_men_n61_));
  NO3        u051(.A(men_men_n61_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n62_));
  NA2        u052(.A(i_8_), .B(men_men_n23_), .Y(men_men_n63_));
  AOI220     u053(.A0(men_men_n40_), .A1(i_1_), .B0(men_men_n36_), .B1(i_2_), .Y(men_men_n64_));
  NOi21      u054(.An(i_1_), .B(i_2_), .Y(men_men_n65_));
  NA3        u055(.A(men_men_n65_), .B(men_men_n46_), .C(i_6_), .Y(men_men_n66_));
  OAI210     u056(.A0(men_men_n64_), .A1(men_men_n63_), .B0(men_men_n66_), .Y(men_men_n67_));
  OAI210     u057(.A0(men_men_n67_), .A1(men_men_n62_), .B0(men_men_n14_), .Y(men_men_n68_));
  NA3        u058(.A(men_men_n56_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n69_));
  NA3        u059(.A(i_1_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n70_));
  NA2        u060(.A(men_men_n70_), .B(men_men_n69_), .Y(men_men_n71_));
  NOi32      u061(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n72_));
  NA2        u062(.A(men_men_n72_), .B(i_3_), .Y(men_men_n73_));
  NA3        u063(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n74_));
  NA2        u064(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n75_));
  NO2        u065(.A(i_0_), .B(i_4_), .Y(men_men_n76_));
  AOI220     u066(.A0(men_men_n76_), .A1(men_men_n75_), .B0(men_men_n71_), .B1(men_men_n53_), .Y(men_men_n77_));
  NA2        u067(.A(men_men_n77_), .B(men_men_n68_), .Y(men_men_n78_));
  NAi21      u068(.An(i_3_), .B(i_6_), .Y(men_men_n79_));
  NO3        u069(.A(men_men_n79_), .B(i_0_), .C(men_men_n45_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n32_), .B(i_5_), .Y(men_men_n81_));
  NOi21      u071(.An(i_7_), .B(i_8_), .Y(men_men_n82_));
  NOi31      u072(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n83_));
  AOI210     u073(.A0(men_men_n82_), .A1(men_men_n12_), .B0(men_men_n83_), .Y(men_men_n84_));
  OAI210     u074(.A0(men_men_n84_), .A1(men_men_n11_), .B0(men_men_n81_), .Y(men_men_n85_));
  OAI210     u075(.A0(men_men_n85_), .A1(men_men_n80_), .B0(men_men_n65_), .Y(men_men_n86_));
  INV        u076(.A(i_5_), .Y(men_men_n87_));
  NA3        u077(.A(men_men_n61_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n88_));
  NO2        u078(.A(men_men_n88_), .B(men_men_n87_), .Y(men_men_n89_));
  INV        u079(.A(men_men_n89_), .Y(men_men_n90_));
  NA3        u080(.A(men_men_n56_), .B(men_men_n31_), .C(i_3_), .Y(men_men_n91_));
  NA2        u081(.A(men_men_n39_), .B(i_6_), .Y(men_men_n92_));
  AOI210     u082(.A0(men_men_n92_), .A1(men_men_n22_), .B0(men_men_n91_), .Y(men_men_n93_));
  NAi21      u083(.An(i_6_), .B(i_0_), .Y(men_men_n94_));
  NOi21      u084(.An(i_4_), .B(i_6_), .Y(men_men_n95_));
  NOi21      u085(.An(i_5_), .B(i_3_), .Y(men_men_n96_));
  NA3        u086(.A(men_men_n96_), .B(men_men_n65_), .C(men_men_n95_), .Y(men_men_n97_));
  INV        u087(.A(men_men_n97_), .Y(men_men_n98_));
  NA2        u088(.A(men_men_n65_), .B(men_men_n32_), .Y(men_men_n99_));
  NOi21      u089(.An(men_men_n37_), .B(men_men_n99_), .Y(men_men_n100_));
  NO3        u090(.A(men_men_n100_), .B(men_men_n98_), .C(men_men_n93_), .Y(men_men_n101_));
  INV        u091(.A(i_1_), .Y(men_men_n102_));
  NA2        u092(.A(men_men_n102_), .B(i_7_), .Y(men_men_n103_));
  NOi21      u093(.An(men_men_n46_), .B(men_men_n103_), .Y(men_men_n104_));
  NA2        u094(.A(men_men_n56_), .B(men_men_n12_), .Y(men_men_n105_));
  NA2        u095(.A(men_men_n32_), .B(men_men_n14_), .Y(men_men_n106_));
  NOi21      u096(.An(i_3_), .B(i_1_), .Y(men_men_n107_));
  NA2        u097(.A(men_men_n107_), .B(i_4_), .Y(men_men_n108_));
  AOI210     u098(.A0(men_men_n106_), .A1(men_men_n105_), .B0(men_men_n108_), .Y(men_men_n109_));
  NOi31      u099(.An(men_men_n40_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n110_));
  NO3        u100(.A(men_men_n110_), .B(men_men_n109_), .C(men_men_n104_), .Y(men_men_n111_));
  NA4        u101(.A(men_men_n111_), .B(men_men_n101_), .C(men_men_n90_), .D(men_men_n86_), .Y(men_men_n112_));
  NOi31      u102(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n113_));
  NOi31      u103(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n114_));
  OAI210     u104(.A0(men_men_n114_), .A1(men_men_n113_), .B0(i_7_), .Y(men_men_n115_));
  NA3        u105(.A(men_men_n32_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NA2        u107(.A(men_men_n117_), .B(men_men_n35_), .Y(men_men_n118_));
  NA4        u108(.A(men_men_n54_), .B(i_2_), .C(men_men_n17_), .D(men_men_n12_), .Y(men_men_n119_));
  NAi31      u109(.An(men_men_n94_), .B(men_men_n82_), .C(i_2_), .Y(men_men_n120_));
  NA3        u110(.A(men_men_n56_), .B(men_men_n52_), .C(i_6_), .Y(men_men_n121_));
  NA3        u111(.A(men_men_n121_), .B(men_men_n120_), .C(men_men_n119_), .Y(men_men_n122_));
  NOi21      u112(.An(i_0_), .B(i_2_), .Y(men_men_n123_));
  NA3        u113(.A(men_men_n123_), .B(men_men_n33_), .C(men_men_n95_), .Y(men_men_n124_));
  NA3        u114(.A(men_men_n46_), .B(men_men_n37_), .C(men_men_n18_), .Y(men_men_n125_));
  NA3        u115(.A(men_men_n123_), .B(men_men_n53_), .C(men_men_n32_), .Y(men_men_n126_));
  NA3        u116(.A(men_men_n126_), .B(men_men_n125_), .C(men_men_n124_), .Y(men_men_n127_));
  NA4        u117(.A(men_men_n52_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n128_));
  NA3        u118(.A(men_men_n34_), .B(men_men_n17_), .C(i_8_), .Y(men_men_n129_));
  NA2        u119(.A(men_men_n129_), .B(men_men_n128_), .Y(men_men_n130_));
  NO3        u120(.A(men_men_n130_), .B(men_men_n127_), .C(men_men_n122_), .Y(men_men_n131_));
  NA2        u121(.A(men_men_n54_), .B(men_men_n28_), .Y(men_men_n132_));
  NO2        u122(.A(men_men_n132_), .B(men_men_n92_), .Y(men_men_n133_));
  NO3        u123(.A(i_2_), .B(men_men_n11_), .C(men_men_n14_), .Y(men_men_n134_));
  NA2        u124(.A(i_2_), .B(i_4_), .Y(men_men_n135_));
  AOI210     u125(.A0(men_men_n94_), .A1(men_men_n79_), .B0(men_men_n135_), .Y(men_men_n136_));
  NO2        u126(.A(i_8_), .B(i_7_), .Y(men_men_n137_));
  OA210      u127(.A0(men_men_n136_), .A1(men_men_n134_), .B0(men_men_n137_), .Y(men_men_n138_));
  NA2        u128(.A(i_5_), .B(men_men_n23_), .Y(men_men_n139_));
  NO2        u129(.A(men_men_n139_), .B(i_4_), .Y(men_men_n140_));
  NO3        u130(.A(men_men_n140_), .B(men_men_n138_), .C(men_men_n133_), .Y(men_men_n141_));
  NA3        u131(.A(men_men_n123_), .B(men_men_n56_), .C(men_men_n95_), .Y(men_men_n142_));
  OAI210     u132(.A0(men_men_n91_), .A1(men_men_n27_), .B0(men_men_n142_), .Y(men_men_n143_));
  NA2        u133(.A(men_men_n96_), .B(men_men_n39_), .Y(men_men_n144_));
  NOi31      u134(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n145_));
  NA2        u135(.A(men_men_n72_), .B(men_men_n145_), .Y(men_men_n146_));
  NA2        u136(.A(men_men_n146_), .B(men_men_n144_), .Y(men_men_n147_));
  NO2        u137(.A(men_men_n147_), .B(men_men_n143_), .Y(men_men_n148_));
  NA4        u138(.A(men_men_n148_), .B(men_men_n141_), .C(men_men_n131_), .D(men_men_n118_), .Y(men_men_n149_));
  OR4        u139(.A(men_men_n149_), .B(men_men_n112_), .C(men_men_n78_), .D(men_men_n60_), .Y(men00));
  INV        u140(.A(i_1_), .Y(men_men_n153_));
  INV        u141(.A(i_5_), .Y(men_men_n154_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule