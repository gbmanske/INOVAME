//Benchmark atmr_max1024_476_0.25

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n383_, mai_mai_n384_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n404_, men_men_n405_, men_men_n406_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO3        o012(.A(ori_ori_n27_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  NA3        o021(.A(x7), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n38_));
  NA2        o022(.A(x4), .B(x3), .Y(ori_ori_n39_));
  AOI210     o023(.A0(ori_ori_n38_), .A1(ori_ori_n23_), .B0(ori_ori_n39_), .Y(ori_ori_n40_));
  NO2        o024(.A(x2), .B(x0), .Y(ori_ori_n41_));
  INV        o025(.A(x3), .Y(ori_ori_n42_));
  NO2        o026(.A(ori_ori_n42_), .B(ori_ori_n18_), .Y(ori_ori_n43_));
  INV        o027(.A(ori_ori_n43_), .Y(ori_ori_n44_));
  NO2        o028(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n45_));
  OAI210     o029(.A0(ori_ori_n45_), .A1(ori_ori_n44_), .B0(ori_ori_n41_), .Y(ori_ori_n46_));
  INV        o030(.A(x4), .Y(ori_ori_n47_));
  NO2        o031(.A(ori_ori_n47_), .B(ori_ori_n17_), .Y(ori_ori_n48_));
  NA2        o032(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n49_));
  OAI210     o033(.A0(ori_ori_n49_), .A1(ori_ori_n20_), .B0(ori_ori_n46_), .Y(ori_ori_n50_));
  NA2        o034(.A(x7), .B(ori_ori_n37_), .Y(ori_ori_n51_));
  AOI220     o035(.A0(ori_ori_n51_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n52_));
  INV        o036(.A(x2), .Y(ori_ori_n53_));
  NO2        o037(.A(ori_ori_n53_), .B(ori_ori_n17_), .Y(ori_ori_n54_));
  NA2        o038(.A(ori_ori_n42_), .B(ori_ori_n18_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n55_), .B(ori_ori_n54_), .Y(ori_ori_n56_));
  OAI210     o040(.A0(ori_ori_n52_), .A1(ori_ori_n32_), .B0(ori_ori_n56_), .Y(ori_ori_n57_));
  NO3        o041(.A(ori_ori_n57_), .B(ori_ori_n50_), .C(ori_ori_n40_), .Y(ori01));
  NA2        o042(.A(ori_ori_n42_), .B(x1), .Y(ori_ori_n59_));
  INV        o043(.A(x9), .Y(ori_ori_n60_));
  NO2        o044(.A(x7), .B(x6), .Y(ori_ori_n61_));
  NO2        o045(.A(ori_ori_n59_), .B(x5), .Y(ori_ori_n62_));
  NO2        o046(.A(x2), .B(x1), .Y(ori_ori_n63_));
  OA210      o047(.A0(ori_ori_n63_), .A1(ori_ori_n62_), .B0(ori_ori_n61_), .Y(ori_ori_n64_));
  OAI210     o048(.A0(ori_ori_n43_), .A1(ori_ori_n25_), .B0(ori_ori_n53_), .Y(ori_ori_n65_));
  OAI210     o049(.A0(ori_ori_n55_), .A1(ori_ori_n20_), .B0(ori_ori_n65_), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n66_), .B(ori_ori_n64_), .Y(ori_ori_n67_));
  NA2        o051(.A(ori_ori_n67_), .B(x4), .Y(ori_ori_n68_));
  NA2        o052(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n69_));
  OAI210     o053(.A0(ori_ori_n69_), .A1(ori_ori_n55_), .B0(x0), .Y(ori_ori_n70_));
  NA2        o054(.A(x5), .B(x3), .Y(ori_ori_n71_));
  NO2        o055(.A(x8), .B(x6), .Y(ori_ori_n72_));
  NAi21      o056(.An(x4), .B(x3), .Y(ori_ori_n73_));
  INV        o057(.A(ori_ori_n73_), .Y(ori_ori_n74_));
  NO2        o058(.A(ori_ori_n74_), .B(ori_ori_n22_), .Y(ori_ori_n75_));
  NO2        o059(.A(x4), .B(x2), .Y(ori_ori_n76_));
  NO2        o060(.A(ori_ori_n76_), .B(x3), .Y(ori_ori_n77_));
  NO3        o061(.A(ori_ori_n77_), .B(ori_ori_n75_), .C(ori_ori_n18_), .Y(ori_ori_n78_));
  NO2        o062(.A(ori_ori_n78_), .B(ori_ori_n70_), .Y(ori_ori_n79_));
  NA2        o063(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n80_));
  INV        o064(.A(x8), .Y(ori_ori_n81_));
  NA2        o065(.A(x2), .B(x1), .Y(ori_ori_n82_));
  AOI210     o066(.A0(ori_ori_n55_), .A1(ori_ori_n25_), .B0(ori_ori_n53_), .Y(ori_ori_n83_));
  OAI210     o067(.A0(ori_ori_n44_), .A1(ori_ori_n37_), .B0(ori_ori_n47_), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n84_), .B(ori_ori_n83_), .Y(ori_ori_n85_));
  NA2        o069(.A(x4), .B(ori_ori_n42_), .Y(ori_ori_n86_));
  NO2        o070(.A(ori_ori_n47_), .B(ori_ori_n53_), .Y(ori_ori_n87_));
  AOI210     o071(.A0(ori_ori_n86_), .A1(ori_ori_n51_), .B0(x1), .Y(ori_ori_n88_));
  NO2        o072(.A(x3), .B(x2), .Y(ori_ori_n89_));
  NA3        o073(.A(ori_ori_n89_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n90_));
  AOI210     o074(.A0(x8), .A1(x6), .B0(ori_ori_n90_), .Y(ori_ori_n91_));
  NA2        o075(.A(ori_ori_n53_), .B(x1), .Y(ori_ori_n92_));
  OAI210     o076(.A0(ori_ori_n92_), .A1(ori_ori_n39_), .B0(ori_ori_n17_), .Y(ori_ori_n93_));
  NO4        o077(.A(ori_ori_n93_), .B(ori_ori_n91_), .C(ori_ori_n88_), .D(ori_ori_n85_), .Y(ori_ori_n94_));
  AO210      o078(.A0(ori_ori_n79_), .A1(ori_ori_n68_), .B0(ori_ori_n94_), .Y(ori02));
  NO2        o079(.A(x3), .B(ori_ori_n53_), .Y(ori_ori_n96_));
  NA2        o080(.A(ori_ori_n53_), .B(ori_ori_n17_), .Y(ori_ori_n97_));
  NA2        o081(.A(ori_ori_n42_), .B(x0), .Y(ori_ori_n98_));
  INV        o082(.A(ori_ori_n98_), .Y(ori_ori_n99_));
  NA2        o083(.A(ori_ori_n99_), .B(x1), .Y(ori_ori_n100_));
  NO3        o084(.A(ori_ori_n100_), .B(x7), .C(x5), .Y(ori_ori_n101_));
  INV        o085(.A(x8), .Y(ori_ori_n102_));
  NO2        o086(.A(x4), .B(x1), .Y(ori_ori_n103_));
  NA2        o087(.A(ori_ori_n103_), .B(x2), .Y(ori_ori_n104_));
  NOi21      o088(.An(x0), .B(x4), .Y(ori_ori_n105_));
  AOI210     o089(.A0(ori_ori_n354_), .A1(ori_ori_n104_), .B0(ori_ori_n71_), .Y(ori_ori_n106_));
  NO2        o090(.A(x5), .B(ori_ori_n47_), .Y(ori_ori_n107_));
  NA2        o091(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n108_));
  AOI210     o092(.A0(ori_ori_n108_), .A1(ori_ori_n92_), .B0(ori_ori_n98_), .Y(ori_ori_n109_));
  OAI210     o093(.A0(ori_ori_n109_), .A1(ori_ori_n35_), .B0(ori_ori_n107_), .Y(ori_ori_n110_));
  NO2        o094(.A(x7), .B(x0), .Y(ori_ori_n111_));
  NO2        o095(.A(ori_ori_n76_), .B(ori_ori_n87_), .Y(ori_ori_n112_));
  NO2        o096(.A(ori_ori_n112_), .B(x3), .Y(ori_ori_n113_));
  NA2        o097(.A(ori_ori_n111_), .B(ori_ori_n113_), .Y(ori_ori_n114_));
  NO2        o098(.A(ori_ori_n21_), .B(ori_ori_n42_), .Y(ori_ori_n115_));
  NO2        o099(.A(ori_ori_n47_), .B(x2), .Y(ori_ori_n116_));
  NA2        o100(.A(ori_ori_n116_), .B(ori_ori_n115_), .Y(ori_ori_n117_));
  NA4        o101(.A(ori_ori_n117_), .B(ori_ori_n114_), .C(ori_ori_n110_), .D(ori_ori_n36_), .Y(ori_ori_n118_));
  NO3        o102(.A(ori_ori_n118_), .B(ori_ori_n106_), .C(ori_ori_n101_), .Y(ori_ori_n119_));
  NO3        o103(.A(ori_ori_n71_), .B(ori_ori_n69_), .C(ori_ori_n24_), .Y(ori_ori_n120_));
  NO2        o104(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n121_));
  NA2        o105(.A(x7), .B(x3), .Y(ori_ori_n122_));
  NO2        o106(.A(ori_ori_n86_), .B(x5), .Y(ori_ori_n123_));
  NO2        o107(.A(x9), .B(x7), .Y(ori_ori_n124_));
  NOi21      o108(.An(x8), .B(x0), .Y(ori_ori_n125_));
  OA210      o109(.A0(ori_ori_n124_), .A1(x1), .B0(ori_ori_n125_), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n42_), .B(x2), .Y(ori_ori_n127_));
  INV        o111(.A(x7), .Y(ori_ori_n128_));
  NA2        o112(.A(ori_ori_n128_), .B(ori_ori_n18_), .Y(ori_ori_n129_));
  AOI220     o113(.A0(ori_ori_n129_), .A1(ori_ori_n127_), .B0(ori_ori_n96_), .B1(x7), .Y(ori_ori_n130_));
  NO2        o114(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n131_));
  NO2        o115(.A(ori_ori_n131_), .B(ori_ori_n105_), .Y(ori_ori_n132_));
  NO2        o116(.A(ori_ori_n132_), .B(ori_ori_n130_), .Y(ori_ori_n133_));
  AOI210     o117(.A0(ori_ori_n126_), .A1(ori_ori_n123_), .B0(ori_ori_n133_), .Y(ori_ori_n134_));
  OAI210     o118(.A0(ori_ori_n122_), .A1(ori_ori_n49_), .B0(ori_ori_n134_), .Y(ori_ori_n135_));
  NA2        o119(.A(x5), .B(x1), .Y(ori_ori_n136_));
  INV        o120(.A(ori_ori_n136_), .Y(ori_ori_n137_));
  AOI210     o121(.A0(ori_ori_n137_), .A1(ori_ori_n105_), .B0(ori_ori_n36_), .Y(ori_ori_n138_));
  NAi21      o122(.An(x2), .B(x7), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n139_), .B(ori_ori_n47_), .Y(ori_ori_n140_));
  NA2        o124(.A(ori_ori_n140_), .B(ori_ori_n62_), .Y(ori_ori_n141_));
  NAi31      o125(.An(ori_ori_n71_), .B(x7), .C(ori_ori_n35_), .Y(ori_ori_n142_));
  NA3        o126(.A(ori_ori_n142_), .B(ori_ori_n141_), .C(ori_ori_n138_), .Y(ori_ori_n143_));
  NO3        o127(.A(ori_ori_n143_), .B(ori_ori_n135_), .C(ori_ori_n120_), .Y(ori_ori_n144_));
  NO2        o128(.A(ori_ori_n144_), .B(ori_ori_n119_), .Y(ori_ori_n145_));
  NA2        o129(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n146_));
  NA2        o130(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n147_));
  NA3        o131(.A(ori_ori_n147_), .B(ori_ori_n146_), .C(ori_ori_n24_), .Y(ori_ori_n148_));
  AN2        o132(.A(ori_ori_n148_), .B(ori_ori_n116_), .Y(ori_ori_n149_));
  NA2        o133(.A(x8), .B(x0), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n128_), .B(ori_ori_n25_), .Y(ori_ori_n151_));
  NA2        o135(.A(x2), .B(x0), .Y(ori_ori_n152_));
  NA2        o136(.A(x4), .B(x1), .Y(ori_ori_n153_));
  NAi21      o137(.An(ori_ori_n103_), .B(ori_ori_n153_), .Y(ori_ori_n154_));
  NOi21      o138(.An(ori_ori_n154_), .B(ori_ori_n152_), .Y(ori_ori_n155_));
  NO2        o139(.A(ori_ori_n155_), .B(ori_ori_n149_), .Y(ori_ori_n156_));
  NO2        o140(.A(ori_ori_n156_), .B(ori_ori_n42_), .Y(ori_ori_n157_));
  NO2        o141(.A(ori_ori_n148_), .B(ori_ori_n69_), .Y(ori_ori_n158_));
  INV        o142(.A(ori_ori_n107_), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n92_), .B(ori_ori_n17_), .Y(ori_ori_n160_));
  AOI210     o144(.A0(ori_ori_n35_), .A1(ori_ori_n81_), .B0(ori_ori_n160_), .Y(ori_ori_n161_));
  NO3        o145(.A(ori_ori_n161_), .B(ori_ori_n159_), .C(x7), .Y(ori_ori_n162_));
  NA3        o146(.A(ori_ori_n154_), .B(ori_ori_n159_), .C(ori_ori_n41_), .Y(ori_ori_n163_));
  OAI210     o147(.A0(ori_ori_n147_), .A1(ori_ori_n112_), .B0(ori_ori_n163_), .Y(ori_ori_n164_));
  NO3        o148(.A(ori_ori_n164_), .B(ori_ori_n162_), .C(ori_ori_n158_), .Y(ori_ori_n165_));
  NO2        o149(.A(ori_ori_n165_), .B(x3), .Y(ori_ori_n166_));
  NO3        o150(.A(ori_ori_n166_), .B(ori_ori_n157_), .C(ori_ori_n145_), .Y(ori03));
  NO2        o151(.A(ori_ori_n47_), .B(x3), .Y(ori_ori_n168_));
  NO2        o152(.A(ori_ori_n71_), .B(x6), .Y(ori_ori_n169_));
  NA2        o153(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n170_));
  NO2        o154(.A(ori_ori_n170_), .B(x4), .Y(ori_ori_n171_));
  NO2        o155(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n172_));
  INV        o156(.A(ori_ori_n169_), .Y(ori_ori_n173_));
  NA2        o157(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n174_), .B(ori_ori_n170_), .Y(ori_ori_n175_));
  NA2        o159(.A(x9), .B(ori_ori_n53_), .Y(ori_ori_n176_));
  INV        o160(.A(ori_ori_n175_), .Y(ori_ori_n177_));
  NO3        o161(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n178_));
  NO2        o162(.A(x5), .B(x1), .Y(ori_ori_n179_));
  NO2        o163(.A(ori_ori_n174_), .B(ori_ori_n146_), .Y(ori_ori_n180_));
  NO3        o164(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n181_));
  AOI220     o165(.A0(ori_ori_n181_), .A1(ori_ori_n47_), .B0(ori_ori_n178_), .B1(ori_ori_n107_), .Y(ori_ori_n182_));
  NA3        o166(.A(ori_ori_n182_), .B(ori_ori_n177_), .C(ori_ori_n173_), .Y(ori_ori_n183_));
  NO2        o167(.A(ori_ori_n47_), .B(ori_ori_n42_), .Y(ori_ori_n184_));
  NA2        o168(.A(ori_ori_n184_), .B(ori_ori_n19_), .Y(ori_ori_n185_));
  NO2        o169(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n186_));
  NO2        o170(.A(ori_ori_n186_), .B(x6), .Y(ori_ori_n187_));
  NOi21      o171(.An(ori_ori_n76_), .B(ori_ori_n187_), .Y(ori_ori_n188_));
  NA2        o172(.A(ori_ori_n186_), .B(x6), .Y(ori_ori_n189_));
  AOI210     o173(.A0(ori_ori_n189_), .A1(ori_ori_n188_), .B0(ori_ori_n128_), .Y(ori_ori_n190_));
  AO210      o174(.A0(ori_ori_n190_), .A1(ori_ori_n185_), .B0(ori_ori_n151_), .Y(ori_ori_n191_));
  NA2        o175(.A(ori_ori_n42_), .B(ori_ori_n53_), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n153_), .B(x6), .Y(ori_ori_n193_));
  NA2        o177(.A(ori_ori_n193_), .B(x5), .Y(ori_ori_n194_));
  NA2        o178(.A(x6), .B(ori_ori_n47_), .Y(ori_ori_n195_));
  NO2        o179(.A(ori_ori_n136_), .B(ori_ori_n42_), .Y(ori_ori_n196_));
  OAI210     o180(.A0(ori_ori_n196_), .A1(ori_ori_n180_), .B0(ori_ori_n352_), .Y(ori_ori_n197_));
  NA2        o181(.A(ori_ori_n107_), .B(x6), .Y(ori_ori_n198_));
  INV        o182(.A(ori_ori_n62_), .Y(ori_ori_n199_));
  NA3        o183(.A(ori_ori_n199_), .B(ori_ori_n198_), .C(ori_ori_n197_), .Y(ori_ori_n200_));
  NA2        o184(.A(ori_ori_n200_), .B(x2), .Y(ori_ori_n201_));
  NA3        o185(.A(ori_ori_n201_), .B(ori_ori_n194_), .C(ori_ori_n191_), .Y(ori_ori_n202_));
  AOI210     o186(.A0(ori_ori_n183_), .A1(x8), .B0(ori_ori_n202_), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n81_), .B(x3), .Y(ori_ori_n204_));
  NA2        o188(.A(ori_ori_n204_), .B(ori_ori_n171_), .Y(ori_ori_n205_));
  NO3        o189(.A(ori_ori_n80_), .B(ori_ori_n72_), .C(ori_ori_n25_), .Y(ori_ori_n206_));
  AOI210     o190(.A0(ori_ori_n187_), .A1(ori_ori_n131_), .B0(ori_ori_n206_), .Y(ori_ori_n207_));
  AOI210     o191(.A0(ori_ori_n207_), .A1(ori_ori_n205_), .B0(x2), .Y(ori_ori_n208_));
  NO2        o192(.A(x4), .B(ori_ori_n53_), .Y(ori_ori_n209_));
  AOI220     o193(.A0(ori_ori_n171_), .A1(ori_ori_n160_), .B0(ori_ori_n209_), .B1(ori_ori_n62_), .Y(ori_ori_n210_));
  NA2        o194(.A(ori_ori_n60_), .B(x6), .Y(ori_ori_n211_));
  NA2        o195(.A(ori_ori_n42_), .B(ori_ori_n17_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n174_), .B(x6), .Y(ori_ori_n213_));
  NO2        o197(.A(ori_ori_n174_), .B(x6), .Y(ori_ori_n214_));
  INV        o198(.A(ori_ori_n214_), .Y(ori_ori_n215_));
  NA3        o199(.A(ori_ori_n215_), .B(ori_ori_n213_), .C(ori_ori_n121_), .Y(ori_ori_n216_));
  NA3        o200(.A(ori_ori_n216_), .B(ori_ori_n210_), .C(ori_ori_n128_), .Y(ori_ori_n217_));
  NA2        o201(.A(ori_ori_n60_), .B(x2), .Y(ori_ori_n218_));
  NA2        o202(.A(x6), .B(x2), .Y(ori_ori_n219_));
  NA2        o203(.A(x9), .B(ori_ori_n42_), .Y(ori_ori_n220_));
  NO2        o204(.A(ori_ori_n220_), .B(ori_ori_n170_), .Y(ori_ori_n221_));
  OR3        o205(.A(ori_ori_n221_), .B(ori_ori_n169_), .C(ori_ori_n123_), .Y(ori_ori_n222_));
  NA2        o206(.A(x4), .B(x0), .Y(ori_ori_n223_));
  NA2        o207(.A(ori_ori_n222_), .B(ori_ori_n41_), .Y(ori_ori_n224_));
  NO2        o208(.A(ori_ori_n224_), .B(x8), .Y(ori_ori_n225_));
  INV        o209(.A(ori_ori_n211_), .Y(ori_ori_n226_));
  OAI210     o210(.A0(x0), .A1(ori_ori_n179_), .B0(ori_ori_n226_), .Y(ori_ori_n227_));
  INV        o211(.A(ori_ori_n150_), .Y(ori_ori_n228_));
  OAI210     o212(.A0(ori_ori_n228_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n229_));
  AOI210     o213(.A0(ori_ori_n229_), .A1(ori_ori_n227_), .B0(ori_ori_n192_), .Y(ori_ori_n230_));
  NO4        o214(.A(ori_ori_n230_), .B(ori_ori_n225_), .C(ori_ori_n217_), .D(ori_ori_n208_), .Y(ori_ori_n231_));
  NA2        o215(.A(ori_ori_n214_), .B(x2), .Y(ori_ori_n232_));
  OAI210     o216(.A0(ori_ori_n228_), .A1(x6), .B0(ori_ori_n43_), .Y(ori_ori_n233_));
  AOI210     o217(.A0(ori_ori_n233_), .A1(ori_ori_n232_), .B0(ori_ori_n159_), .Y(ori_ori_n234_));
  NOi21      o218(.An(ori_ori_n219_), .B(ori_ori_n17_), .Y(ori_ori_n235_));
  NA3        o219(.A(ori_ori_n235_), .B(ori_ori_n179_), .C(ori_ori_n39_), .Y(ori_ori_n236_));
  AOI210     o220(.A0(ori_ori_n36_), .A1(ori_ori_n53_), .B0(x0), .Y(ori_ori_n237_));
  NA3        o221(.A(ori_ori_n237_), .B(ori_ori_n137_), .C(ori_ori_n32_), .Y(ori_ori_n238_));
  NA2        o222(.A(x3), .B(x2), .Y(ori_ori_n239_));
  AOI220     o223(.A0(ori_ori_n239_), .A1(ori_ori_n192_), .B0(ori_ori_n238_), .B1(ori_ori_n236_), .Y(ori_ori_n240_));
  NAi21      o224(.An(x4), .B(x0), .Y(ori_ori_n241_));
  NO3        o225(.A(ori_ori_n241_), .B(ori_ori_n43_), .C(x2), .Y(ori_ori_n242_));
  OAI210     o226(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n242_), .Y(ori_ori_n243_));
  NO2        o227(.A(ori_ori_n237_), .B(ori_ori_n235_), .Y(ori_ori_n244_));
  AOI220     o228(.A0(ori_ori_n244_), .A1(ori_ori_n74_), .B0(ori_ori_n18_), .B1(ori_ori_n31_), .Y(ori_ori_n245_));
  AOI210     o229(.A0(ori_ori_n245_), .A1(ori_ori_n243_), .B0(ori_ori_n25_), .Y(ori_ori_n246_));
  NA3        o230(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n247_));
  OAI210     o231(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(ori_ori_n247_), .Y(ori_ori_n248_));
  INV        o232(.A(ori_ori_n180_), .Y(ori_ori_n249_));
  NA2        o233(.A(ori_ori_n36_), .B(ori_ori_n42_), .Y(ori_ori_n250_));
  OR2        o234(.A(ori_ori_n250_), .B(ori_ori_n223_), .Y(ori_ori_n251_));
  OAI220     o235(.A0(ori_ori_n251_), .A1(ori_ori_n136_), .B0(ori_ori_n195_), .B1(ori_ori_n249_), .Y(ori_ori_n252_));
  AO210      o236(.A0(ori_ori_n248_), .A1(ori_ori_n123_), .B0(ori_ori_n252_), .Y(ori_ori_n253_));
  NO4        o237(.A(ori_ori_n253_), .B(ori_ori_n246_), .C(ori_ori_n240_), .D(ori_ori_n234_), .Y(ori_ori_n254_));
  OAI210     o238(.A0(ori_ori_n231_), .A1(ori_ori_n203_), .B0(ori_ori_n254_), .Y(ori04));
  NO2        o239(.A(x2), .B(x1), .Y(ori_ori_n256_));
  OAI210     o240(.A0(ori_ori_n212_), .A1(ori_ori_n256_), .B0(ori_ori_n36_), .Y(ori_ori_n257_));
  NO2        o241(.A(ori_ori_n256_), .B(ori_ori_n241_), .Y(ori_ori_n258_));
  AOI210     o242(.A0(ori_ori_n60_), .A1(x4), .B0(ori_ori_n97_), .Y(ori_ori_n259_));
  OAI210     o243(.A0(ori_ori_n259_), .A1(ori_ori_n258_), .B0(ori_ori_n204_), .Y(ori_ori_n260_));
  NO2        o244(.A(ori_ori_n239_), .B(ori_ori_n172_), .Y(ori_ori_n261_));
  NA2        o245(.A(x9), .B(x0), .Y(ori_ori_n262_));
  AOI210     o246(.A0(ori_ori_n80_), .A1(ori_ori_n69_), .B0(ori_ori_n262_), .Y(ori_ori_n263_));
  OAI210     o247(.A0(ori_ori_n263_), .A1(ori_ori_n261_), .B0(ori_ori_n81_), .Y(ori_ori_n264_));
  NA3        o248(.A(ori_ori_n264_), .B(x6), .C(ori_ori_n260_), .Y(ori_ori_n265_));
  NA2        o249(.A(ori_ori_n265_), .B(ori_ori_n257_), .Y(ori_ori_n266_));
  NO2        o250(.A(ori_ori_n176_), .B(ori_ori_n98_), .Y(ori_ori_n267_));
  NO3        o251(.A(ori_ori_n211_), .B(x2), .C(ori_ori_n18_), .Y(ori_ori_n268_));
  NO2        o252(.A(ori_ori_n268_), .B(ori_ori_n267_), .Y(ori_ori_n269_));
  OAI210     o253(.A0(x8), .A1(ori_ori_n92_), .B0(ori_ori_n150_), .Y(ori_ori_n270_));
  NA3        o254(.A(ori_ori_n270_), .B(x6), .C(x3), .Y(ori_ori_n271_));
  NOi21      o255(.An(ori_ori_n125_), .B(ori_ori_n108_), .Y(ori_ori_n272_));
  AOI210     o256(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n273_));
  OAI220     o257(.A0(ori_ori_n273_), .A1(ori_ori_n250_), .B0(ori_ori_n218_), .B1(ori_ori_n247_), .Y(ori_ori_n274_));
  AOI210     o258(.A0(ori_ori_n272_), .A1(x6), .B0(ori_ori_n274_), .Y(ori_ori_n275_));
  NA2        o259(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n276_));
  OAI210     o260(.A0(ori_ori_n92_), .A1(ori_ori_n17_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  NA2        o261(.A(ori_ori_n277_), .B(ori_ori_n72_), .Y(ori_ori_n278_));
  NA4        o262(.A(ori_ori_n278_), .B(ori_ori_n275_), .C(ori_ori_n271_), .D(ori_ori_n269_), .Y(ori_ori_n279_));
  OAI210     o263(.A0(x1), .A1(x3), .B0(ori_ori_n242_), .Y(ori_ori_n280_));
  NA2        o264(.A(ori_ori_n178_), .B(ori_ori_n76_), .Y(ori_ori_n281_));
  NA3        o265(.A(ori_ori_n281_), .B(ori_ori_n280_), .C(ori_ori_n128_), .Y(ori_ori_n282_));
  AOI210     o266(.A0(ori_ori_n279_), .A1(x4), .B0(ori_ori_n282_), .Y(ori_ori_n283_));
  NA3        o267(.A(ori_ori_n258_), .B(ori_ori_n176_), .C(ori_ori_n81_), .Y(ori_ori_n284_));
  NA2        o268(.A(x4), .B(ori_ori_n82_), .Y(ori_ori_n285_));
  AOI210     o269(.A0(ori_ori_n285_), .A1(ori_ori_n284_), .B0(x3), .Y(ori_ori_n286_));
  INV        o270(.A(ori_ori_n82_), .Y(ori_ori_n287_));
  NO2        o271(.A(ori_ori_n81_), .B(x4), .Y(ori_ori_n288_));
  AOI220     o272(.A0(ori_ori_n288_), .A1(ori_ori_n43_), .B0(ori_ori_n105_), .B1(ori_ori_n287_), .Y(ori_ori_n289_));
  NA3        o273(.A(ori_ori_n289_), .B(ori_ori_n185_), .C(x6), .Y(ori_ori_n290_));
  NO2        o274(.A(ori_ori_n125_), .B(ori_ori_n73_), .Y(ori_ori_n291_));
  NO2        o275(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n292_));
  NOi21      o276(.An(ori_ori_n103_), .B(ori_ori_n27_), .Y(ori_ori_n293_));
  AOI210     o277(.A0(ori_ori_n292_), .A1(ori_ori_n291_), .B0(ori_ori_n293_), .Y(ori_ori_n294_));
  OAI210     o278(.A0(ori_ori_n152_), .A1(ori_ori_n60_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  OAI220     o279(.A0(ori_ori_n295_), .A1(x6), .B0(ori_ori_n290_), .B1(ori_ori_n286_), .Y(ori_ori_n296_));
  OAI210     o280(.A0(x6), .A1(ori_ori_n47_), .B0(ori_ori_n41_), .Y(ori_ori_n297_));
  OAI210     o281(.A0(ori_ori_n297_), .A1(ori_ori_n81_), .B0(ori_ori_n251_), .Y(ori_ori_n298_));
  AOI210     o282(.A0(ori_ori_n298_), .A1(ori_ori_n18_), .B0(ori_ori_n128_), .Y(ori_ori_n299_));
  AO220      o283(.A0(ori_ori_n299_), .A1(ori_ori_n296_), .B0(ori_ori_n283_), .B1(ori_ori_n266_), .Y(ori_ori_n300_));
  NA2        o284(.A(ori_ori_n292_), .B(x6), .Y(ori_ori_n301_));
  AOI210     o285(.A0(x6), .A1(x1), .B0(ori_ori_n127_), .Y(ori_ori_n302_));
  NA2        o286(.A(ori_ori_n288_), .B(x0), .Y(ori_ori_n303_));
  NA2        o287(.A(ori_ori_n76_), .B(x6), .Y(ori_ori_n304_));
  OAI210     o288(.A0(ori_ori_n303_), .A1(ori_ori_n302_), .B0(ori_ori_n304_), .Y(ori_ori_n305_));
  AOI220     o289(.A0(ori_ori_n305_), .A1(ori_ori_n301_), .B0(ori_ori_n181_), .B1(ori_ori_n48_), .Y(ori_ori_n306_));
  NA2        o290(.A(ori_ori_n306_), .B(ori_ori_n300_), .Y(ori_ori_n307_));
  NA2        o291(.A(ori_ori_n168_), .B(ori_ori_n128_), .Y(ori_ori_n308_));
  OAI210     o292(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n192_), .Y(ori_ori_n309_));
  AO220      o293(.A0(ori_ori_n309_), .A1(ori_ori_n124_), .B0(ori_ori_n96_), .B1(x4), .Y(ori_ori_n310_));
  NA3        o294(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n311_));
  NA2        o295(.A(ori_ori_n184_), .B(x0), .Y(ori_ori_n312_));
  OAI220     o296(.A0(ori_ori_n312_), .A1(ori_ori_n176_), .B0(ori_ori_n311_), .B1(ori_ori_n287_), .Y(ori_ori_n313_));
  AOI210     o297(.A0(ori_ori_n310_), .A1(ori_ori_n102_), .B0(ori_ori_n313_), .Y(ori_ori_n314_));
  AOI210     o298(.A0(ori_ori_n314_), .A1(ori_ori_n308_), .B0(ori_ori_n25_), .Y(ori_ori_n315_));
  NA2        o299(.A(ori_ori_n315_), .B(x6), .Y(ori_ori_n316_));
  NO2        o300(.A(x0), .B(ori_ori_n32_), .Y(ori_ori_n317_));
  NO2        o301(.A(ori_ori_n128_), .B(x0), .Y(ori_ori_n318_));
  AOI220     o302(.A0(ori_ori_n318_), .A1(ori_ori_n184_), .B0(ori_ori_n168_), .B1(ori_ori_n128_), .Y(ori_ori_n319_));
  AOI210     o303(.A0(x7), .A1(ori_ori_n209_), .B0(x1), .Y(ori_ori_n320_));
  OAI210     o304(.A0(ori_ori_n319_), .A1(x8), .B0(ori_ori_n320_), .Y(ori_ori_n321_));
  NAi31      o305(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n322_));
  OAI210     o306(.A0(ori_ori_n322_), .A1(x4), .B0(ori_ori_n139_), .Y(ori_ori_n323_));
  NA3        o307(.A(ori_ori_n323_), .B(ori_ori_n122_), .C(x9), .Y(ori_ori_n324_));
  NA2        o308(.A(ori_ori_n291_), .B(ori_ori_n128_), .Y(ori_ori_n325_));
  NA4        o309(.A(ori_ori_n325_), .B(x1), .C(ori_ori_n324_), .D(ori_ori_n49_), .Y(ori_ori_n326_));
  OAI210     o310(.A0(ori_ori_n321_), .A1(ori_ori_n317_), .B0(ori_ori_n326_), .Y(ori_ori_n327_));
  NOi31      o311(.An(ori_ori_n318_), .B(ori_ori_n32_), .C(x8), .Y(ori_ori_n328_));
  NA2        o312(.A(ori_ori_n353_), .B(ori_ori_n128_), .Y(ori_ori_n329_));
  NO2        o313(.A(ori_ori_n329_), .B(ori_ori_n53_), .Y(ori_ori_n330_));
  NO2        o314(.A(ori_ori_n330_), .B(ori_ori_n328_), .Y(ori_ori_n331_));
  AOI210     o315(.A0(ori_ori_n331_), .A1(ori_ori_n327_), .B0(ori_ori_n25_), .Y(ori_ori_n332_));
  NA4        o316(.A(ori_ori_n31_), .B(ori_ori_n81_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n333_));
  NO3        o317(.A(ori_ori_n218_), .B(ori_ori_n150_), .C(ori_ori_n39_), .Y(ori_ori_n334_));
  NA2        o318(.A(ori_ori_n334_), .B(x7), .Y(ori_ori_n335_));
  NA2        o319(.A(ori_ori_n335_), .B(ori_ori_n333_), .Y(ori_ori_n336_));
  OAI210     o320(.A0(ori_ori_n336_), .A1(ori_ori_n332_), .B0(ori_ori_n36_), .Y(ori_ori_n337_));
  NA2        o321(.A(ori_ori_n212_), .B(ori_ori_n21_), .Y(ori_ori_n338_));
  NO2        o322(.A(ori_ori_n136_), .B(ori_ori_n111_), .Y(ori_ori_n339_));
  NA2        o323(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  AOI210     o324(.A0(ori_ori_n340_), .A1(ori_ori_n142_), .B0(ori_ori_n28_), .Y(ori_ori_n341_));
  NA2        o325(.A(ori_ori_n53_), .B(ori_ori_n322_), .Y(ori_ori_n342_));
  NA2        o326(.A(ori_ori_n342_), .B(ori_ori_n151_), .Y(ori_ori_n343_));
  OAI220     o327(.A0(ori_ori_n220_), .A1(x2), .B0(ori_ori_n136_), .B1(ori_ori_n42_), .Y(ori_ori_n344_));
  NA2        o328(.A(ori_ori_n344_), .B(ori_ori_n111_), .Y(ori_ori_n345_));
  AOI210     o329(.A0(ori_ori_n345_), .A1(ori_ori_n343_), .B0(ori_ori_n195_), .Y(ori_ori_n346_));
  NO2        o330(.A(ori_ori_n346_), .B(ori_ori_n341_), .Y(ori_ori_n347_));
  NA3        o331(.A(ori_ori_n347_), .B(ori_ori_n337_), .C(ori_ori_n316_), .Y(ori_ori_n348_));
  AOI210     o332(.A0(ori_ori_n307_), .A1(ori_ori_n25_), .B0(ori_ori_n348_), .Y(ori05));
  INV        o333(.A(x6), .Y(ori_ori_n352_));
  INV        o334(.A(x4), .Y(ori_ori_n353_));
  INV        o335(.A(x0), .Y(ori_ori_n354_));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  NAi21      m004(.An(mai_mai_n20_), .B(mai_mai_n19_), .Y(mai_mai_n21_));
  NA2        m005(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n22_));
  INV        m006(.A(x5), .Y(mai_mai_n23_));
  NA2        m007(.A(x7), .B(x6), .Y(mai_mai_n24_));
  NA2        m008(.A(x8), .B(x3), .Y(mai_mai_n25_));
  NA2        m009(.A(x4), .B(x2), .Y(mai_mai_n26_));
  INV        m010(.A(mai_mai_n22_), .Y(mai_mai_n27_));
  NO2        m011(.A(x4), .B(x3), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OA210      m013(.A0(mai_mai_n29_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n30_));
  NOi31      m014(.An(mai_mai_n21_), .B(mai_mai_n30_), .C(mai_mai_n27_), .Y(mai00));
  NO2        m015(.A(x1), .B(x0), .Y(mai_mai_n32_));
  INV        m016(.A(x6), .Y(mai_mai_n33_));
  NO2        m017(.A(mai_mai_n33_), .B(mai_mai_n23_), .Y(mai_mai_n34_));
  NA2        m018(.A(x4), .B(x3), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n21_), .B(mai_mai_n35_), .Y(mai_mai_n36_));
  NO2        m020(.A(x2), .B(x0), .Y(mai_mai_n37_));
  INV        m021(.A(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n39_));
  INV        m023(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m024(.A(mai_mai_n34_), .B(x4), .Y(mai_mai_n41_));
  OAI210     m025(.A0(mai_mai_n41_), .A1(mai_mai_n40_), .B0(mai_mai_n37_), .Y(mai_mai_n42_));
  INV        m026(.A(x4), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n43_), .B(mai_mai_n17_), .Y(mai_mai_n44_));
  NA2        m028(.A(mai_mai_n44_), .B(x2), .Y(mai_mai_n45_));
  NA2        m029(.A(mai_mai_n45_), .B(mai_mai_n42_), .Y(mai_mai_n46_));
  AOI210     m030(.A0(mai_mai_n20_), .A1(mai_mai_n19_), .B0(mai_mai_n32_), .Y(mai_mai_n47_));
  INV        m031(.A(x2), .Y(mai_mai_n48_));
  NO2        m032(.A(mai_mai_n48_), .B(mai_mai_n17_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n38_), .B(mai_mai_n18_), .Y(mai_mai_n50_));
  NA2        m034(.A(mai_mai_n50_), .B(mai_mai_n49_), .Y(mai_mai_n51_));
  OAI210     m035(.A0(mai_mai_n47_), .A1(mai_mai_n29_), .B0(mai_mai_n51_), .Y(mai_mai_n52_));
  NO3        m036(.A(mai_mai_n52_), .B(mai_mai_n46_), .C(mai_mai_n36_), .Y(mai01));
  NA2        m037(.A(x8), .B(x7), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n38_), .B(x1), .Y(mai_mai_n55_));
  INV        m039(.A(x9), .Y(mai_mai_n56_));
  NO2        m040(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n57_));
  NO2        m041(.A(mai_mai_n55_), .B(x5), .Y(mai_mai_n58_));
  NO2        m042(.A(x8), .B(x2), .Y(mai_mai_n59_));
  OAI210     m043(.A0(mai_mai_n39_), .A1(mai_mai_n23_), .B0(mai_mai_n48_), .Y(mai_mai_n60_));
  OAI210     m044(.A0(mai_mai_n50_), .A1(mai_mai_n20_), .B0(mai_mai_n60_), .Y(mai_mai_n61_));
  NAi31      m045(.An(x1), .B(x9), .C(x5), .Y(mai_mai_n62_));
  INV        m046(.A(mai_mai_n61_), .Y(mai_mai_n63_));
  OAI210     m047(.A0(mai_mai_n63_), .A1(mai_mai_n57_), .B0(x4), .Y(mai_mai_n64_));
  NA2        m048(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n65_));
  OAI210     m049(.A0(mai_mai_n65_), .A1(mai_mai_n50_), .B0(x0), .Y(mai_mai_n66_));
  NA2        m050(.A(x5), .B(x3), .Y(mai_mai_n67_));
  NO2        m051(.A(x8), .B(x6), .Y(mai_mai_n68_));
  NO2        m052(.A(mai_mai_n67_), .B(mai_mai_n48_), .Y(mai_mai_n69_));
  NAi21      m053(.An(x4), .B(x3), .Y(mai_mai_n70_));
  INV        m054(.A(mai_mai_n70_), .Y(mai_mai_n71_));
  NO2        m055(.A(mai_mai_n71_), .B(mai_mai_n20_), .Y(mai_mai_n72_));
  NO2        m056(.A(x4), .B(x2), .Y(mai_mai_n73_));
  NO2        m057(.A(mai_mai_n73_), .B(x3), .Y(mai_mai_n74_));
  NO3        m058(.A(mai_mai_n74_), .B(mai_mai_n72_), .C(mai_mai_n18_), .Y(mai_mai_n75_));
  NO3        m059(.A(mai_mai_n75_), .B(mai_mai_n69_), .C(mai_mai_n66_), .Y(mai_mai_n76_));
  NO4        m060(.A(x7), .B(x6), .C(mai_mai_n38_), .D(x1), .Y(mai_mai_n77_));
  NA2        m061(.A(mai_mai_n56_), .B(mai_mai_n43_), .Y(mai_mai_n78_));
  INV        m062(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m063(.A0(mai_mai_n77_), .A1(mai_mai_n58_), .B0(mai_mai_n79_), .Y(mai_mai_n80_));
  NA2        m064(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n81_));
  NO2        m065(.A(mai_mai_n81_), .B(mai_mai_n23_), .Y(mai_mai_n82_));
  INV        m066(.A(x8), .Y(mai_mai_n83_));
  NO2        m067(.A(x2), .B(mai_mai_n82_), .Y(mai_mai_n84_));
  NO2        m068(.A(mai_mai_n84_), .B(mai_mai_n24_), .Y(mai_mai_n85_));
  AOI210     m069(.A0(mai_mai_n50_), .A1(mai_mai_n23_), .B0(mai_mai_n48_), .Y(mai_mai_n86_));
  NA2        m070(.A(mai_mai_n40_), .B(mai_mai_n43_), .Y(mai_mai_n87_));
  NO3        m071(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(mai_mai_n85_), .Y(mai_mai_n88_));
  NA2        m072(.A(x4), .B(mai_mai_n38_), .Y(mai_mai_n89_));
  NO2        m073(.A(mai_mai_n43_), .B(mai_mai_n48_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n89_), .B(x1), .Y(mai_mai_n91_));
  NO2        m075(.A(x3), .B(x2), .Y(mai_mai_n92_));
  NA2        m076(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n93_));
  OAI210     m077(.A0(mai_mai_n93_), .A1(mai_mai_n35_), .B0(mai_mai_n17_), .Y(mai_mai_n94_));
  NO3        m078(.A(mai_mai_n94_), .B(mai_mai_n91_), .C(mai_mai_n88_), .Y(mai_mai_n95_));
  AO220      m079(.A0(mai_mai_n95_), .A1(mai_mai_n80_), .B0(mai_mai_n76_), .B1(mai_mai_n64_), .Y(mai02));
  NO2        m080(.A(x3), .B(mai_mai_n48_), .Y(mai_mai_n97_));
  NO2        m081(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n98_));
  OAI210     m082(.A0(mai_mai_n78_), .A1(x2), .B0(x3), .Y(mai_mai_n99_));
  AOI220     m083(.A0(mai_mai_n99_), .A1(mai_mai_n98_), .B0(mai_mai_n97_), .B1(x4), .Y(mai_mai_n100_));
  NO3        m084(.A(mai_mai_n100_), .B(x7), .C(x5), .Y(mai_mai_n101_));
  OR2        m085(.A(x8), .B(x0), .Y(mai_mai_n102_));
  INV        m086(.A(mai_mai_n102_), .Y(mai_mai_n103_));
  NAi21      m087(.An(x2), .B(x8), .Y(mai_mai_n104_));
  INV        m088(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NO2        m089(.A(x4), .B(x1), .Y(mai_mai_n106_));
  NOi21      m090(.An(x0), .B(x1), .Y(mai_mai_n107_));
  NO3        m091(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n108_));
  NOi21      m092(.An(x0), .B(x4), .Y(mai_mai_n109_));
  NO2        m093(.A(x5), .B(mai_mai_n43_), .Y(mai_mai_n110_));
  NA2        m094(.A(mai_mai_n32_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  NAi21      m095(.An(x0), .B(x4), .Y(mai_mai_n112_));
  NO2        m096(.A(mai_mai_n112_), .B(x1), .Y(mai_mai_n113_));
  NO2        m097(.A(x7), .B(x0), .Y(mai_mai_n114_));
  NO2        m098(.A(mai_mai_n73_), .B(mai_mai_n90_), .Y(mai_mai_n115_));
  NO2        m099(.A(mai_mai_n115_), .B(x3), .Y(mai_mai_n116_));
  OAI210     m100(.A0(mai_mai_n114_), .A1(mai_mai_n113_), .B0(mai_mai_n116_), .Y(mai_mai_n117_));
  NA2        m101(.A(x5), .B(x0), .Y(mai_mai_n118_));
  NO2        m102(.A(mai_mai_n43_), .B(x2), .Y(mai_mai_n119_));
  NA3        m103(.A(mai_mai_n119_), .B(mai_mai_n118_), .C(x3), .Y(mai_mai_n120_));
  NA4        m104(.A(mai_mai_n120_), .B(mai_mai_n117_), .C(mai_mai_n111_), .D(mai_mai_n33_), .Y(mai_mai_n121_));
  NO2        m105(.A(mai_mai_n121_), .B(mai_mai_n101_), .Y(mai_mai_n122_));
  NO3        m106(.A(mai_mai_n67_), .B(mai_mai_n65_), .C(mai_mai_n22_), .Y(mai_mai_n123_));
  NO2        m107(.A(mai_mai_n26_), .B(mai_mai_n23_), .Y(mai_mai_n124_));
  AOI220     m108(.A0(mai_mai_n107_), .A1(mai_mai_n124_), .B0(mai_mai_n58_), .B1(mai_mai_n17_), .Y(mai_mai_n125_));
  NO3        m109(.A(mai_mai_n125_), .B(mai_mai_n54_), .C(mai_mai_n56_), .Y(mai_mai_n126_));
  NA2        m110(.A(x7), .B(x3), .Y(mai_mai_n127_));
  NO2        m111(.A(mai_mai_n89_), .B(x5), .Y(mai_mai_n128_));
  NO2        m112(.A(x9), .B(x7), .Y(mai_mai_n129_));
  NOi21      m113(.An(x8), .B(x0), .Y(mai_mai_n130_));
  NO2        m114(.A(mai_mai_n38_), .B(x2), .Y(mai_mai_n131_));
  INV        m115(.A(x7), .Y(mai_mai_n132_));
  NA2        m116(.A(mai_mai_n132_), .B(mai_mai_n18_), .Y(mai_mai_n133_));
  NO2        m117(.A(mai_mai_n23_), .B(x4), .Y(mai_mai_n134_));
  NA2        m118(.A(mai_mai_n130_), .B(mai_mai_n128_), .Y(mai_mai_n135_));
  OAI210     m119(.A0(mai_mai_n127_), .A1(mai_mai_n45_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NA2        m120(.A(x5), .B(x1), .Y(mai_mai_n137_));
  INV        m121(.A(mai_mai_n137_), .Y(mai_mai_n138_));
  AOI210     m122(.A0(mai_mai_n138_), .A1(mai_mai_n109_), .B0(mai_mai_n33_), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n56_), .B(mai_mai_n83_), .Y(mai_mai_n140_));
  NO2        m124(.A(x2), .B(mai_mai_n140_), .Y(mai_mai_n141_));
  NA2        m125(.A(mai_mai_n141_), .B(mai_mai_n58_), .Y(mai_mai_n142_));
  NA2        m126(.A(mai_mai_n142_), .B(mai_mai_n139_), .Y(mai_mai_n143_));
  NO4        m127(.A(mai_mai_n143_), .B(mai_mai_n136_), .C(mai_mai_n126_), .D(mai_mai_n123_), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n144_), .B(mai_mai_n122_), .Y(mai_mai_n145_));
  NO2        m129(.A(mai_mai_n118_), .B(mai_mai_n115_), .Y(mai_mai_n146_));
  NA2        m130(.A(mai_mai_n23_), .B(mai_mai_n18_), .Y(mai_mai_n147_));
  NA2        m131(.A(mai_mai_n23_), .B(mai_mai_n17_), .Y(mai_mai_n148_));
  NA3        m132(.A(mai_mai_n148_), .B(mai_mai_n147_), .C(mai_mai_n22_), .Y(mai_mai_n149_));
  AN2        m133(.A(mai_mai_n149_), .B(mai_mai_n119_), .Y(mai_mai_n150_));
  NA2        m134(.A(x8), .B(x0), .Y(mai_mai_n151_));
  NO2        m135(.A(mai_mai_n132_), .B(mai_mai_n23_), .Y(mai_mai_n152_));
  NO2        m136(.A(mai_mai_n107_), .B(x4), .Y(mai_mai_n153_));
  NA2        m137(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  AOI210     m138(.A0(mai_mai_n151_), .A1(x1), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  NA2        m139(.A(x2), .B(x0), .Y(mai_mai_n156_));
  NA2        m140(.A(x4), .B(x1), .Y(mai_mai_n157_));
  NAi21      m141(.An(mai_mai_n106_), .B(mai_mai_n157_), .Y(mai_mai_n158_));
  NOi31      m142(.An(mai_mai_n158_), .B(mai_mai_n134_), .C(mai_mai_n156_), .Y(mai_mai_n159_));
  NO4        m143(.A(mai_mai_n159_), .B(mai_mai_n155_), .C(mai_mai_n150_), .D(mai_mai_n146_), .Y(mai_mai_n160_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n38_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n149_), .B(mai_mai_n65_), .Y(mai_mai_n162_));
  INV        m146(.A(mai_mai_n110_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n93_), .B(mai_mai_n17_), .Y(mai_mai_n164_));
  NA2        m148(.A(mai_mai_n158_), .B(mai_mai_n37_), .Y(mai_mai_n165_));
  OAI210     m149(.A0(mai_mai_n148_), .A1(mai_mai_n115_), .B0(mai_mai_n165_), .Y(mai_mai_n166_));
  NO2        m150(.A(mai_mai_n166_), .B(mai_mai_n162_), .Y(mai_mai_n167_));
  NO2        m151(.A(mai_mai_n167_), .B(x3), .Y(mai_mai_n168_));
  NO3        m152(.A(mai_mai_n168_), .B(mai_mai_n161_), .C(mai_mai_n145_), .Y(mai03));
  NO2        m153(.A(mai_mai_n43_), .B(x3), .Y(mai_mai_n170_));
  NO2        m154(.A(x6), .B(mai_mai_n23_), .Y(mai_mai_n171_));
  NO2        m155(.A(mai_mai_n48_), .B(x1), .Y(mai_mai_n172_));
  OAI210     m156(.A0(mai_mai_n172_), .A1(mai_mai_n23_), .B0(x6), .Y(mai_mai_n173_));
  NO2        m157(.A(mai_mai_n173_), .B(mai_mai_n17_), .Y(mai_mai_n174_));
  NA2        m158(.A(mai_mai_n174_), .B(mai_mai_n170_), .Y(mai_mai_n175_));
  NO2        m159(.A(mai_mai_n67_), .B(x6), .Y(mai_mai_n176_));
  NA2        m160(.A(x6), .B(mai_mai_n23_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n177_), .B(x4), .Y(mai_mai_n178_));
  NO2        m162(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n179_));
  AO220      m163(.A0(mai_mai_n179_), .A1(mai_mai_n178_), .B0(mai_mai_n176_), .B1(mai_mai_n49_), .Y(mai_mai_n180_));
  NA2        m164(.A(mai_mai_n180_), .B(mai_mai_n56_), .Y(mai_mai_n181_));
  NA2        m165(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n182_));
  AOI210     m166(.A0(mai_mai_n23_), .A1(x3), .B0(mai_mai_n156_), .Y(mai_mai_n183_));
  NA2        m167(.A(mai_mai_n183_), .B(mai_mai_n23_), .Y(mai_mai_n184_));
  NO3        m168(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n185_));
  NO2        m169(.A(x5), .B(x1), .Y(mai_mai_n186_));
  NA2        m170(.A(mai_mai_n186_), .B(mai_mai_n17_), .Y(mai_mai_n187_));
  NO3        m171(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n188_));
  NA2        m172(.A(mai_mai_n383_), .B(mai_mai_n43_), .Y(mai_mai_n189_));
  NA4        m173(.A(mai_mai_n189_), .B(mai_mai_n184_), .C(mai_mai_n181_), .D(mai_mai_n175_), .Y(mai_mai_n190_));
  NO2        m174(.A(mai_mai_n43_), .B(mai_mai_n38_), .Y(mai_mai_n191_));
  NA2        m175(.A(mai_mai_n191_), .B(mai_mai_n19_), .Y(mai_mai_n192_));
  NO2        m176(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n193_));
  INV        m177(.A(x6), .Y(mai_mai_n194_));
  NOi21      m178(.An(mai_mai_n73_), .B(mai_mai_n194_), .Y(mai_mai_n195_));
  NA2        m179(.A(mai_mai_n56_), .B(mai_mai_n83_), .Y(mai_mai_n196_));
  NO2        m180(.A(mai_mai_n195_), .B(mai_mai_n132_), .Y(mai_mai_n197_));
  NA2        m181(.A(mai_mai_n38_), .B(mai_mai_n48_), .Y(mai_mai_n198_));
  OAI210     m182(.A0(mai_mai_n198_), .A1(mai_mai_n23_), .B0(mai_mai_n148_), .Y(mai_mai_n199_));
  NO3        m183(.A(mai_mai_n157_), .B(mai_mai_n56_), .C(x6), .Y(mai_mai_n200_));
  AOI220     m184(.A0(mai_mai_n200_), .A1(mai_mai_n199_), .B0(mai_mai_n119_), .B1(mai_mai_n82_), .Y(mai_mai_n201_));
  NA2        m185(.A(x6), .B(mai_mai_n43_), .Y(mai_mai_n202_));
  OAI210     m186(.A0(mai_mai_n103_), .A1(mai_mai_n68_), .B0(x4), .Y(mai_mai_n203_));
  AOI210     m187(.A0(mai_mai_n203_), .A1(mai_mai_n202_), .B0(mai_mai_n67_), .Y(mai_mai_n204_));
  NA2        m188(.A(mai_mai_n171_), .B(mai_mai_n113_), .Y(mai_mai_n205_));
  NA3        m189(.A(mai_mai_n182_), .B(mai_mai_n110_), .C(x6), .Y(mai_mai_n206_));
  OAI210     m190(.A0(mai_mai_n83_), .A1(mai_mai_n33_), .B0(mai_mai_n58_), .Y(mai_mai_n207_));
  NA3        m191(.A(mai_mai_n207_), .B(mai_mai_n206_), .C(mai_mai_n205_), .Y(mai_mai_n208_));
  OAI210     m192(.A0(mai_mai_n208_), .A1(mai_mai_n204_), .B0(x2), .Y(mai_mai_n209_));
  NA3        m193(.A(mai_mai_n209_), .B(mai_mai_n201_), .C(mai_mai_n197_), .Y(mai_mai_n210_));
  AOI210     m194(.A0(mai_mai_n190_), .A1(x8), .B0(mai_mai_n210_), .Y(mai_mai_n211_));
  NO2        m195(.A(mai_mai_n81_), .B(mai_mai_n23_), .Y(mai_mai_n212_));
  AOI210     m196(.A0(mai_mai_n194_), .A1(mai_mai_n134_), .B0(mai_mai_n212_), .Y(mai_mai_n213_));
  NO2        m197(.A(mai_mai_n213_), .B(x2), .Y(mai_mai_n214_));
  AOI220     m198(.A0(mai_mai_n178_), .A1(mai_mai_n164_), .B0(x2), .B1(mai_mai_n58_), .Y(mai_mai_n215_));
  NA3        m199(.A(mai_mai_n23_), .B(x3), .C(x2), .Y(mai_mai_n216_));
  AOI210     m200(.A0(mai_mai_n216_), .A1(mai_mai_n118_), .B0(x9), .Y(mai_mai_n217_));
  NA2        m201(.A(mai_mai_n38_), .B(mai_mai_n17_), .Y(mai_mai_n218_));
  NO2        m202(.A(mai_mai_n218_), .B(mai_mai_n23_), .Y(mai_mai_n219_));
  OAI210     m203(.A0(mai_mai_n219_), .A1(mai_mai_n217_), .B0(mai_mai_n106_), .Y(mai_mai_n220_));
  NA2        m204(.A(mai_mai_n182_), .B(x6), .Y(mai_mai_n221_));
  NO2        m205(.A(mai_mai_n182_), .B(x6), .Y(mai_mai_n222_));
  NAi21      m206(.An(mai_mai_n140_), .B(mai_mai_n222_), .Y(mai_mai_n223_));
  NA3        m207(.A(mai_mai_n223_), .B(mai_mai_n221_), .C(mai_mai_n124_), .Y(mai_mai_n224_));
  NA4        m208(.A(mai_mai_n224_), .B(mai_mai_n220_), .C(mai_mai_n215_), .D(mai_mai_n132_), .Y(mai_mai_n225_));
  NA2        m209(.A(mai_mai_n171_), .B(mai_mai_n193_), .Y(mai_mai_n226_));
  NO2        m210(.A(x9), .B(x6), .Y(mai_mai_n227_));
  NO2        m211(.A(mai_mai_n118_), .B(mai_mai_n18_), .Y(mai_mai_n228_));
  NAi21      m212(.An(mai_mai_n228_), .B(mai_mai_n216_), .Y(mai_mai_n229_));
  NAi21      m213(.An(x1), .B(x4), .Y(mai_mai_n230_));
  AOI210     m214(.A0(x3), .A1(x2), .B0(mai_mai_n43_), .Y(mai_mai_n231_));
  OAI210     m215(.A0(mai_mai_n118_), .A1(x3), .B0(mai_mai_n231_), .Y(mai_mai_n232_));
  AOI220     m216(.A0(mai_mai_n232_), .A1(mai_mai_n230_), .B0(mai_mai_n229_), .B1(mai_mai_n227_), .Y(mai_mai_n233_));
  NA2        m217(.A(mai_mai_n233_), .B(mai_mai_n226_), .Y(mai_mai_n234_));
  NA2        m218(.A(mai_mai_n56_), .B(x2), .Y(mai_mai_n235_));
  NO2        m219(.A(mai_mai_n235_), .B(mai_mai_n226_), .Y(mai_mai_n236_));
  NO3        m220(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n237_));
  NA2        m221(.A(x6), .B(x2), .Y(mai_mai_n238_));
  NO2        m222(.A(mai_mai_n238_), .B(mai_mai_n147_), .Y(mai_mai_n239_));
  NO2        m223(.A(mai_mai_n237_), .B(mai_mai_n239_), .Y(mai_mai_n240_));
  OAI220     m224(.A0(mai_mai_n240_), .A1(mai_mai_n38_), .B0(mai_mai_n153_), .B1(mai_mai_n41_), .Y(mai_mai_n241_));
  OAI210     m225(.A0(mai_mai_n241_), .A1(mai_mai_n236_), .B0(mai_mai_n234_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n176_), .B(mai_mai_n37_), .Y(mai_mai_n243_));
  AOI210     m227(.A0(mai_mai_n243_), .A1(mai_mai_n242_), .B0(x8), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n228_), .A1(mai_mai_n186_), .B0(x6), .Y(mai_mai_n245_));
  NO2        m229(.A(mai_mai_n245_), .B(mai_mai_n198_), .Y(mai_mai_n246_));
  NO4        m230(.A(mai_mai_n246_), .B(mai_mai_n244_), .C(mai_mai_n225_), .D(mai_mai_n214_), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n140_), .B(x1), .Y(mai_mai_n248_));
  NO3        m232(.A(mai_mai_n248_), .B(x3), .C(mai_mai_n33_), .Y(mai_mai_n249_));
  OAI210     m233(.A0(mai_mai_n249_), .A1(mai_mai_n222_), .B0(x2), .Y(mai_mai_n250_));
  OAI210     m234(.A0(x8), .A1(x6), .B0(mai_mai_n39_), .Y(mai_mai_n251_));
  AOI210     m235(.A0(mai_mai_n251_), .A1(mai_mai_n250_), .B0(mai_mai_n163_), .Y(mai_mai_n252_));
  NOi21      m236(.An(mai_mai_n238_), .B(mai_mai_n17_), .Y(mai_mai_n253_));
  NA3        m237(.A(mai_mai_n253_), .B(mai_mai_n186_), .C(mai_mai_n35_), .Y(mai_mai_n254_));
  AOI210     m238(.A0(mai_mai_n33_), .A1(mai_mai_n48_), .B0(x0), .Y(mai_mai_n255_));
  NA3        m239(.A(mai_mai_n255_), .B(mai_mai_n138_), .C(mai_mai_n29_), .Y(mai_mai_n256_));
  NA2        m240(.A(x3), .B(x2), .Y(mai_mai_n257_));
  AOI220     m241(.A0(mai_mai_n257_), .A1(mai_mai_n198_), .B0(mai_mai_n256_), .B1(mai_mai_n254_), .Y(mai_mai_n258_));
  NAi21      m242(.An(x4), .B(x0), .Y(mai_mai_n259_));
  NO3        m243(.A(mai_mai_n259_), .B(mai_mai_n39_), .C(x2), .Y(mai_mai_n260_));
  OAI210     m244(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n260_), .Y(mai_mai_n261_));
  NO2        m245(.A(x9), .B(x8), .Y(mai_mai_n262_));
  NA3        m246(.A(mai_mai_n262_), .B(mai_mai_n33_), .C(mai_mai_n48_), .Y(mai_mai_n263_));
  OAI210     m247(.A0(mai_mai_n255_), .A1(mai_mai_n253_), .B0(mai_mai_n263_), .Y(mai_mai_n264_));
  NA2        m248(.A(mai_mai_n264_), .B(mai_mai_n71_), .Y(mai_mai_n265_));
  AOI210     m249(.A0(mai_mai_n265_), .A1(mai_mai_n261_), .B0(mai_mai_n23_), .Y(mai_mai_n266_));
  NO2        m250(.A(mai_mai_n255_), .B(mai_mai_n253_), .Y(mai_mai_n267_));
  AN2        m251(.A(mai_mai_n267_), .B(mai_mai_n128_), .Y(mai_mai_n268_));
  NO4        m252(.A(mai_mai_n268_), .B(mai_mai_n266_), .C(mai_mai_n258_), .D(mai_mai_n252_), .Y(mai_mai_n269_));
  OAI210     m253(.A0(mai_mai_n247_), .A1(mai_mai_n211_), .B0(mai_mai_n269_), .Y(mai04));
  OAI210     m254(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n271_));
  NA3        m255(.A(mai_mai_n271_), .B(mai_mai_n237_), .C(mai_mai_n74_), .Y(mai_mai_n272_));
  NO2        m256(.A(x2), .B(x1), .Y(mai_mai_n273_));
  OAI210     m257(.A0(mai_mai_n218_), .A1(mai_mai_n273_), .B0(mai_mai_n33_), .Y(mai_mai_n274_));
  NO2        m258(.A(mai_mai_n273_), .B(mai_mai_n259_), .Y(mai_mai_n275_));
  NO2        m259(.A(mai_mai_n235_), .B(mai_mai_n81_), .Y(mai_mai_n276_));
  NO2        m260(.A(mai_mai_n276_), .B(mai_mai_n33_), .Y(mai_mai_n277_));
  NO2        m261(.A(mai_mai_n257_), .B(mai_mai_n179_), .Y(mai_mai_n278_));
  NA2        m262(.A(mai_mai_n278_), .B(mai_mai_n83_), .Y(mai_mai_n279_));
  NA2        m263(.A(mai_mai_n279_), .B(mai_mai_n277_), .Y(mai_mai_n280_));
  NA2        m264(.A(mai_mai_n280_), .B(mai_mai_n274_), .Y(mai_mai_n281_));
  NO3        m265(.A(x9), .B(mai_mai_n104_), .C(mai_mai_n18_), .Y(mai_mai_n282_));
  INV        m266(.A(mai_mai_n282_), .Y(mai_mai_n283_));
  OAI210     m267(.A0(mai_mai_n102_), .A1(mai_mai_n93_), .B0(mai_mai_n151_), .Y(mai_mai_n284_));
  NA3        m268(.A(mai_mai_n284_), .B(x6), .C(x3), .Y(mai_mai_n285_));
  NA2        m269(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n286_));
  OAI210     m270(.A0(mai_mai_n93_), .A1(mai_mai_n17_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  AOI220     m271(.A0(mai_mai_n287_), .A1(mai_mai_n68_), .B0(mai_mai_n276_), .B1(mai_mai_n83_), .Y(mai_mai_n288_));
  NA3        m272(.A(mai_mai_n288_), .B(mai_mai_n285_), .C(mai_mai_n283_), .Y(mai_mai_n289_));
  OAI210     m273(.A0(mai_mai_n98_), .A1(x3), .B0(mai_mai_n260_), .Y(mai_mai_n290_));
  NA3        m274(.A(mai_mai_n196_), .B(mai_mai_n185_), .C(mai_mai_n73_), .Y(mai_mai_n291_));
  NA3        m275(.A(mai_mai_n291_), .B(mai_mai_n290_), .C(mai_mai_n132_), .Y(mai_mai_n292_));
  AOI210     m276(.A0(mai_mai_n289_), .A1(x4), .B0(mai_mai_n292_), .Y(mai_mai_n293_));
  NA2        m277(.A(mai_mai_n275_), .B(mai_mai_n83_), .Y(mai_mai_n294_));
  NOi21      m278(.An(x4), .B(x0), .Y(mai_mai_n295_));
  XO2        m279(.A(x4), .B(x0), .Y(mai_mai_n296_));
  AOI210     m280(.A0(x2), .A1(x8), .B0(mai_mai_n295_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n297_), .A1(mai_mai_n294_), .B0(x3), .Y(mai_mai_n298_));
  NO3        m282(.A(mai_mai_n296_), .B(mai_mai_n140_), .C(x2), .Y(mai_mai_n299_));
  NO3        m283(.A(mai_mai_n196_), .B(mai_mai_n26_), .C(mai_mai_n22_), .Y(mai_mai_n300_));
  NO2        m284(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n301_));
  NA3        m285(.A(mai_mai_n301_), .B(mai_mai_n192_), .C(x6), .Y(mai_mai_n302_));
  NO2        m286(.A(mai_mai_n38_), .B(x0), .Y(mai_mai_n303_));
  NO2        m287(.A(mai_mai_n130_), .B(mai_mai_n70_), .Y(mai_mai_n304_));
  NOi21      m288(.An(mai_mai_n106_), .B(mai_mai_n25_), .Y(mai_mai_n305_));
  AOI210     m289(.A0(mai_mai_n384_), .A1(mai_mai_n304_), .B0(mai_mai_n305_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n93_), .A1(mai_mai_n56_), .B0(mai_mai_n306_), .Y(mai_mai_n307_));
  OAI220     m291(.A0(mai_mai_n307_), .A1(x6), .B0(mai_mai_n302_), .B1(mai_mai_n298_), .Y(mai_mai_n308_));
  AO220      m292(.A0(x7), .A1(mai_mai_n308_), .B0(mai_mai_n293_), .B1(mai_mai_n281_), .Y(mai_mai_n309_));
  NA2        m293(.A(mai_mai_n188_), .B(mai_mai_n44_), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n309_), .C(mai_mai_n272_), .Y(mai_mai_n311_));
  AOI210     m295(.A0(mai_mai_n172_), .A1(x8), .B0(mai_mai_n98_), .Y(mai_mai_n312_));
  NA2        m296(.A(mai_mai_n312_), .B(mai_mai_n286_), .Y(mai_mai_n313_));
  NA3        m297(.A(mai_mai_n313_), .B(mai_mai_n170_), .C(mai_mai_n132_), .Y(mai_mai_n314_));
  AO220      m298(.A0(x4), .A1(mai_mai_n129_), .B0(mai_mai_n97_), .B1(x4), .Y(mai_mai_n315_));
  NA3        m299(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n316_));
  NO2        m300(.A(mai_mai_n316_), .B(x2), .Y(mai_mai_n317_));
  AOI210     m301(.A0(mai_mai_n315_), .A1(mai_mai_n103_), .B0(mai_mai_n317_), .Y(mai_mai_n318_));
  AOI210     m302(.A0(mai_mai_n318_), .A1(mai_mai_n314_), .B0(mai_mai_n23_), .Y(mai_mai_n319_));
  NA3        m303(.A(mai_mai_n105_), .B(mai_mai_n191_), .C(x0), .Y(mai_mai_n320_));
  NA2        m304(.A(mai_mai_n170_), .B(mai_mai_n179_), .Y(mai_mai_n321_));
  NO2        m305(.A(mai_mai_n321_), .B(mai_mai_n23_), .Y(mai_mai_n322_));
  AOI210     m306(.A0(mai_mai_n104_), .A1(mai_mai_n102_), .B0(mai_mai_n37_), .Y(mai_mai_n323_));
  NOi21      m307(.An(mai_mai_n323_), .B(mai_mai_n157_), .Y(mai_mai_n324_));
  OAI210     m308(.A0(mai_mai_n324_), .A1(mai_mai_n322_), .B0(mai_mai_n129_), .Y(mai_mai_n325_));
  NAi31      m309(.An(mai_mai_n45_), .B(mai_mai_n248_), .C(mai_mai_n152_), .Y(mai_mai_n326_));
  NA3        m310(.A(mai_mai_n326_), .B(mai_mai_n325_), .C(mai_mai_n320_), .Y(mai_mai_n327_));
  OAI210     m311(.A0(mai_mai_n327_), .A1(mai_mai_n319_), .B0(x6), .Y(mai_mai_n328_));
  OAI210     m312(.A0(mai_mai_n140_), .A1(mai_mai_n43_), .B0(mai_mai_n114_), .Y(mai_mai_n329_));
  AOI210     m313(.A0(mai_mai_n35_), .A1(mai_mai_n29_), .B0(mai_mai_n329_), .Y(mai_mai_n330_));
  NO2        m314(.A(mai_mai_n132_), .B(x0), .Y(mai_mai_n331_));
  AOI220     m315(.A0(mai_mai_n331_), .A1(mai_mai_n191_), .B0(mai_mai_n170_), .B1(mai_mai_n132_), .Y(mai_mai_n332_));
  INV        m316(.A(x1), .Y(mai_mai_n333_));
  OAI210     m317(.A0(mai_mai_n332_), .A1(x8), .B0(mai_mai_n333_), .Y(mai_mai_n334_));
  NO4        m318(.A(x8), .B(mai_mai_n259_), .C(x9), .D(x2), .Y(mai_mai_n335_));
  NOi21      m319(.An(mai_mai_n108_), .B(mai_mai_n156_), .Y(mai_mai_n336_));
  NO3        m320(.A(mai_mai_n336_), .B(mai_mai_n335_), .C(mai_mai_n18_), .Y(mai_mai_n337_));
  NO3        m321(.A(x9), .B(mai_mai_n132_), .C(x0), .Y(mai_mai_n338_));
  AOI220     m322(.A0(mai_mai_n338_), .A1(x8), .B0(mai_mai_n304_), .B1(mai_mai_n132_), .Y(mai_mai_n339_));
  NA2        m323(.A(mai_mai_n339_), .B(mai_mai_n337_), .Y(mai_mai_n340_));
  OAI210     m324(.A0(mai_mai_n334_), .A1(mai_mai_n330_), .B0(mai_mai_n340_), .Y(mai_mai_n341_));
  NOi31      m325(.An(mai_mai_n331_), .B(mai_mai_n29_), .C(x8), .Y(mai_mai_n342_));
  INV        m326(.A(mai_mai_n112_), .Y(mai_mai_n343_));
  NO3        m327(.A(mai_mai_n343_), .B(mai_mai_n108_), .C(mai_mai_n38_), .Y(mai_mai_n344_));
  NOi31      m328(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n345_));
  AOI220     m329(.A0(mai_mai_n345_), .A1(mai_mai_n295_), .B0(mai_mai_n109_), .B1(x3), .Y(mai_mai_n346_));
  AOI210     m330(.A0(mai_mai_n230_), .A1(mai_mai_n54_), .B0(mai_mai_n107_), .Y(mai_mai_n347_));
  OAI210     m331(.A0(mai_mai_n347_), .A1(x3), .B0(mai_mai_n346_), .Y(mai_mai_n348_));
  NO3        m332(.A(mai_mai_n348_), .B(mai_mai_n344_), .C(x2), .Y(mai_mai_n349_));
  NO2        m333(.A(mai_mai_n296_), .B(mai_mai_n262_), .Y(mai_mai_n350_));
  INV        m334(.A(mai_mai_n316_), .Y(mai_mai_n351_));
  AOI220     m335(.A0(mai_mai_n351_), .A1(mai_mai_n83_), .B0(mai_mai_n350_), .B1(mai_mai_n132_), .Y(mai_mai_n352_));
  NO2        m336(.A(mai_mai_n352_), .B(mai_mai_n48_), .Y(mai_mai_n353_));
  NO3        m337(.A(mai_mai_n353_), .B(mai_mai_n349_), .C(mai_mai_n342_), .Y(mai_mai_n354_));
  AOI210     m338(.A0(mai_mai_n354_), .A1(mai_mai_n341_), .B0(mai_mai_n23_), .Y(mai_mai_n355_));
  NO3        m339(.A(mai_mai_n56_), .B(x4), .C(x1), .Y(mai_mai_n356_));
  NO3        m340(.A(mai_mai_n59_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n357_));
  AOI220     m341(.A0(mai_mai_n357_), .A1(mai_mai_n231_), .B0(mai_mai_n356_), .B1(mai_mai_n323_), .Y(mai_mai_n358_));
  NO2        m342(.A(mai_mai_n358_), .B(mai_mai_n92_), .Y(mai_mai_n359_));
  NO3        m343(.A(mai_mai_n235_), .B(mai_mai_n151_), .C(mai_mai_n35_), .Y(mai_mai_n360_));
  OAI210     m344(.A0(mai_mai_n360_), .A1(mai_mai_n359_), .B0(x7), .Y(mai_mai_n361_));
  NA2        m345(.A(mai_mai_n131_), .B(mai_mai_n113_), .Y(mai_mai_n362_));
  NA2        m346(.A(mai_mai_n362_), .B(mai_mai_n361_), .Y(mai_mai_n363_));
  OAI210     m347(.A0(mai_mai_n363_), .A1(mai_mai_n355_), .B0(mai_mai_n33_), .Y(mai_mai_n364_));
  NO2        m348(.A(mai_mai_n338_), .B(mai_mai_n179_), .Y(mai_mai_n365_));
  NO4        m349(.A(mai_mai_n365_), .B(mai_mai_n67_), .C(x4), .D(mai_mai_n48_), .Y(mai_mai_n366_));
  NA2        m350(.A(mai_mai_n303_), .B(mai_mai_n152_), .Y(mai_mai_n367_));
  NA2        m351(.A(x3), .B(mai_mai_n48_), .Y(mai_mai_n368_));
  AOI210     m352(.A0(x2), .A1(mai_mai_n25_), .B0(mai_mai_n62_), .Y(mai_mai_n369_));
  OAI210     m353(.A0(mai_mai_n129_), .A1(mai_mai_n18_), .B0(x7), .Y(mai_mai_n370_));
  NO3        m354(.A(mai_mai_n345_), .B(x3), .C(mai_mai_n48_), .Y(mai_mai_n371_));
  AOI210     m355(.A0(mai_mai_n371_), .A1(mai_mai_n370_), .B0(mai_mai_n369_), .Y(mai_mai_n372_));
  OAI210     m356(.A0(mai_mai_n133_), .A1(mai_mai_n368_), .B0(mai_mai_n372_), .Y(mai_mai_n373_));
  NA2        m357(.A(mai_mai_n373_), .B(x0), .Y(mai_mai_n374_));
  AOI210     m358(.A0(mai_mai_n374_), .A1(mai_mai_n367_), .B0(mai_mai_n202_), .Y(mai_mai_n375_));
  INV        m359(.A(x5), .Y(mai_mai_n376_));
  NO4        m360(.A(mai_mai_n93_), .B(mai_mai_n376_), .C(mai_mai_n54_), .D(mai_mai_n29_), .Y(mai_mai_n377_));
  NO3        m361(.A(mai_mai_n377_), .B(mai_mai_n375_), .C(mai_mai_n366_), .Y(mai_mai_n378_));
  NA3        m362(.A(mai_mai_n378_), .B(mai_mai_n364_), .C(mai_mai_n328_), .Y(mai_mai_n379_));
  AOI210     m363(.A0(mai_mai_n311_), .A1(mai_mai_n23_), .B0(mai_mai_n379_), .Y(mai05));
  INV        m364(.A(mai_mai_n187_), .Y(mai_mai_n383_));
  INV        m365(.A(x2), .Y(mai_mai_n384_));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  INV        u005(.A(men_men_n19_), .Y(men_men_n22_));
  NA2        u006(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n23_));
  INV        u007(.A(x5), .Y(men_men_n24_));
  NA2        u008(.A(x7), .B(x6), .Y(men_men_n25_));
  NA2        u009(.A(x8), .B(x3), .Y(men_men_n26_));
  NA2        u010(.A(x4), .B(x2), .Y(men_men_n27_));
  NO4        u011(.A(men_men_n27_), .B(men_men_n26_), .C(men_men_n25_), .D(men_men_n24_), .Y(men_men_n28_));
  NO2        u012(.A(men_men_n28_), .B(men_men_n23_), .Y(men_men_n29_));
  NO2        u013(.A(x4), .B(x3), .Y(men_men_n30_));
  INV        u014(.A(men_men_n30_), .Y(men_men_n31_));
  NOi21      u015(.An(men_men_n22_), .B(men_men_n29_), .Y(men00));
  NO2        u016(.A(x1), .B(x0), .Y(men_men_n33_));
  INV        u017(.A(x6), .Y(men_men_n34_));
  NO2        u018(.A(men_men_n34_), .B(men_men_n24_), .Y(men_men_n35_));
  AN2        u019(.A(x8), .B(x7), .Y(men_men_n36_));
  NA3        u020(.A(men_men_n36_), .B(men_men_n35_), .C(men_men_n33_), .Y(men_men_n37_));
  NA2        u021(.A(x4), .B(x3), .Y(men_men_n38_));
  AOI210     u022(.A0(men_men_n37_), .A1(men_men_n22_), .B0(men_men_n38_), .Y(men_men_n39_));
  NO2        u023(.A(x2), .B(x0), .Y(men_men_n40_));
  INV        u024(.A(x3), .Y(men_men_n41_));
  NO2        u025(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n42_));
  INV        u026(.A(men_men_n42_), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n35_), .B(x4), .Y(men_men_n44_));
  OAI210     u028(.A0(men_men_n44_), .A1(men_men_n43_), .B0(men_men_n40_), .Y(men_men_n45_));
  INV        u029(.A(x4), .Y(men_men_n46_));
  NO2        u030(.A(men_men_n46_), .B(men_men_n17_), .Y(men_men_n47_));
  NA2        u031(.A(men_men_n47_), .B(x2), .Y(men_men_n48_));
  OAI210     u032(.A0(men_men_n48_), .A1(men_men_n20_), .B0(men_men_n45_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n36_), .B(men_men_n35_), .Y(men_men_n50_));
  NA2        u034(.A(men_men_n50_), .B(men_men_n33_), .Y(men_men_n51_));
  INV        u035(.A(x2), .Y(men_men_n52_));
  NO2        u036(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n53_));
  NA2        u037(.A(men_men_n41_), .B(men_men_n18_), .Y(men_men_n54_));
  NA2        u038(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  OAI210     u039(.A0(men_men_n51_), .A1(men_men_n31_), .B0(men_men_n55_), .Y(men_men_n56_));
  NO3        u040(.A(men_men_n56_), .B(men_men_n49_), .C(men_men_n39_), .Y(men01));
  NA2        u041(.A(x8), .B(x7), .Y(men_men_n58_));
  NA2        u042(.A(men_men_n41_), .B(x1), .Y(men_men_n59_));
  INV        u043(.A(x9), .Y(men_men_n60_));
  NO2        u044(.A(men_men_n60_), .B(men_men_n34_), .Y(men_men_n61_));
  INV        u045(.A(men_men_n61_), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n59_), .Y(men_men_n63_));
  NO2        u047(.A(x7), .B(x6), .Y(men_men_n64_));
  NO2        u048(.A(men_men_n59_), .B(x5), .Y(men_men_n65_));
  NO2        u049(.A(x8), .B(x2), .Y(men_men_n66_));
  INV        u050(.A(men_men_n66_), .Y(men_men_n67_));
  OA210      u051(.A0(men_men_n66_), .A1(men_men_n65_), .B0(men_men_n64_), .Y(men_men_n68_));
  OAI210     u052(.A0(men_men_n42_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n69_));
  OAI210     u053(.A0(men_men_n54_), .A1(men_men_n20_), .B0(men_men_n69_), .Y(men_men_n70_));
  NAi31      u054(.An(x1), .B(x9), .C(x5), .Y(men_men_n71_));
  OAI220     u055(.A0(men_men_n71_), .A1(men_men_n41_), .B0(men_men_n70_), .B1(men_men_n68_), .Y(men_men_n72_));
  OAI210     u056(.A0(men_men_n72_), .A1(men_men_n63_), .B0(x4), .Y(men_men_n73_));
  NA2        u057(.A(men_men_n46_), .B(x2), .Y(men_men_n74_));
  OAI210     u058(.A0(men_men_n74_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n75_));
  NA2        u059(.A(x5), .B(x3), .Y(men_men_n76_));
  NO2        u060(.A(x8), .B(x6), .Y(men_men_n77_));
  NO4        u061(.A(men_men_n77_), .B(men_men_n76_), .C(men_men_n64_), .D(men_men_n52_), .Y(men_men_n78_));
  NAi21      u062(.An(x4), .B(x3), .Y(men_men_n79_));
  INV        u063(.A(men_men_n79_), .Y(men_men_n80_));
  NO2        u064(.A(x4), .B(x2), .Y(men_men_n81_));
  NO2        u065(.A(men_men_n81_), .B(x3), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n79_), .B(men_men_n18_), .Y(men_men_n83_));
  NO3        u067(.A(men_men_n83_), .B(men_men_n78_), .C(men_men_n75_), .Y(men_men_n84_));
  NO3        u068(.A(men_men_n21_), .B(men_men_n41_), .C(x1), .Y(men_men_n85_));
  INV        u069(.A(x4), .Y(men_men_n86_));
  NA2        u070(.A(men_men_n85_), .B(men_men_n86_), .Y(men_men_n87_));
  NA2        u071(.A(x3), .B(men_men_n18_), .Y(men_men_n88_));
  NO2        u072(.A(men_men_n88_), .B(men_men_n24_), .Y(men_men_n89_));
  INV        u073(.A(x8), .Y(men_men_n90_));
  NA2        u074(.A(x2), .B(x1), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n90_), .Y(men_men_n92_));
  NO2        u076(.A(men_men_n92_), .B(men_men_n89_), .Y(men_men_n93_));
  NO2        u077(.A(men_men_n93_), .B(men_men_n25_), .Y(men_men_n94_));
  AOI210     u078(.A0(men_men_n54_), .A1(men_men_n24_), .B0(men_men_n52_), .Y(men_men_n95_));
  OAI210     u079(.A0(men_men_n43_), .A1(men_men_n35_), .B0(men_men_n46_), .Y(men_men_n96_));
  NO3        u080(.A(men_men_n96_), .B(men_men_n95_), .C(men_men_n94_), .Y(men_men_n97_));
  NA2        u081(.A(x4), .B(men_men_n41_), .Y(men_men_n98_));
  NO2        u082(.A(men_men_n46_), .B(men_men_n52_), .Y(men_men_n99_));
  OAI210     u083(.A0(men_men_n99_), .A1(men_men_n41_), .B0(men_men_n18_), .Y(men_men_n100_));
  AOI210     u084(.A0(men_men_n98_), .A1(men_men_n50_), .B0(men_men_n100_), .Y(men_men_n101_));
  NO2        u085(.A(x3), .B(x2), .Y(men_men_n102_));
  NA2        u086(.A(men_men_n102_), .B(men_men_n24_), .Y(men_men_n103_));
  INV        u087(.A(men_men_n103_), .Y(men_men_n104_));
  NA2        u088(.A(men_men_n52_), .B(x1), .Y(men_men_n105_));
  OAI210     u089(.A0(men_men_n105_), .A1(men_men_n38_), .B0(men_men_n17_), .Y(men_men_n106_));
  NO4        u090(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n101_), .D(men_men_n97_), .Y(men_men_n107_));
  AO220      u091(.A0(men_men_n107_), .A1(men_men_n87_), .B0(men_men_n84_), .B1(men_men_n73_), .Y(men02));
  NO2        u092(.A(x3), .B(men_men_n52_), .Y(men_men_n109_));
  NA2        u093(.A(men_men_n52_), .B(men_men_n17_), .Y(men_men_n110_));
  NA2        u094(.A(men_men_n41_), .B(x0), .Y(men_men_n111_));
  NO2        u095(.A(x4), .B(men_men_n110_), .Y(men_men_n112_));
  AOI220     u096(.A0(men_men_n112_), .A1(x1), .B0(men_men_n109_), .B1(x4), .Y(men_men_n113_));
  NO3        u097(.A(men_men_n113_), .B(x7), .C(x5), .Y(men_men_n114_));
  NA2        u098(.A(x9), .B(x2), .Y(men_men_n115_));
  OR2        u099(.A(x8), .B(x0), .Y(men_men_n116_));
  INV        u100(.A(men_men_n116_), .Y(men_men_n117_));
  NAi21      u101(.An(x2), .B(x8), .Y(men_men_n118_));
  INV        u102(.A(men_men_n118_), .Y(men_men_n119_));
  OAI220     u103(.A0(men_men_n119_), .A1(men_men_n117_), .B0(men_men_n115_), .B1(x7), .Y(men_men_n120_));
  NO2        u104(.A(x4), .B(x1), .Y(men_men_n121_));
  NA3        u105(.A(men_men_n121_), .B(men_men_n120_), .C(men_men_n58_), .Y(men_men_n122_));
  NOi21      u106(.An(x0), .B(x1), .Y(men_men_n123_));
  NO3        u107(.A(x9), .B(x8), .C(x7), .Y(men_men_n124_));
  NOi21      u108(.An(x0), .B(x4), .Y(men_men_n125_));
  NAi21      u109(.An(x8), .B(x7), .Y(men_men_n126_));
  NO2        u110(.A(men_men_n126_), .B(men_men_n60_), .Y(men_men_n127_));
  AOI220     u111(.A0(men_men_n127_), .A1(men_men_n125_), .B0(men_men_n124_), .B1(men_men_n123_), .Y(men_men_n128_));
  AOI210     u112(.A0(men_men_n128_), .A1(men_men_n122_), .B0(men_men_n76_), .Y(men_men_n129_));
  NO2        u113(.A(x5), .B(men_men_n46_), .Y(men_men_n130_));
  NA2        u114(.A(x2), .B(men_men_n18_), .Y(men_men_n131_));
  AOI210     u115(.A0(men_men_n131_), .A1(men_men_n105_), .B0(men_men_n111_), .Y(men_men_n132_));
  OAI210     u116(.A0(men_men_n132_), .A1(men_men_n33_), .B0(men_men_n130_), .Y(men_men_n133_));
  NAi21      u117(.An(x0), .B(x4), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x1), .Y(men_men_n135_));
  NO2        u119(.A(x7), .B(x0), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n81_), .B(men_men_n99_), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x3), .Y(men_men_n138_));
  OAI210     u122(.A0(men_men_n136_), .A1(men_men_n135_), .B0(men_men_n138_), .Y(men_men_n139_));
  NA2        u123(.A(x5), .B(x0), .Y(men_men_n140_));
  NO2        u124(.A(men_men_n46_), .B(x2), .Y(men_men_n141_));
  NA3        u125(.A(men_men_n139_), .B(men_men_n133_), .C(men_men_n34_), .Y(men_men_n142_));
  NO3        u126(.A(men_men_n142_), .B(men_men_n129_), .C(men_men_n114_), .Y(men_men_n143_));
  NO2        u127(.A(men_men_n27_), .B(men_men_n24_), .Y(men_men_n144_));
  AOI220     u128(.A0(men_men_n123_), .A1(men_men_n144_), .B0(men_men_n65_), .B1(men_men_n17_), .Y(men_men_n145_));
  NO2        u129(.A(men_men_n145_), .B(men_men_n58_), .Y(men_men_n146_));
  NO2        u130(.A(x9), .B(x7), .Y(men_men_n147_));
  NOi21      u131(.An(x8), .B(x0), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n41_), .B(x2), .Y(men_men_n149_));
  INV        u133(.A(x7), .Y(men_men_n150_));
  NA2        u134(.A(men_men_n150_), .B(men_men_n18_), .Y(men_men_n151_));
  AOI220     u135(.A0(men_men_n151_), .A1(men_men_n149_), .B0(men_men_n109_), .B1(men_men_n36_), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n24_), .B(x4), .Y(men_men_n153_));
  NO2        u137(.A(men_men_n153_), .B(men_men_n125_), .Y(men_men_n154_));
  NO2        u138(.A(men_men_n154_), .B(men_men_n152_), .Y(men_men_n155_));
  NA2        u139(.A(x5), .B(x1), .Y(men_men_n156_));
  INV        u140(.A(men_men_n156_), .Y(men_men_n157_));
  AOI210     u141(.A0(men_men_n157_), .A1(men_men_n125_), .B0(men_men_n34_), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n60_), .B(men_men_n90_), .Y(men_men_n159_));
  NAi21      u143(.An(x2), .B(x7), .Y(men_men_n160_));
  NAi31      u144(.An(men_men_n76_), .B(men_men_n36_), .C(men_men_n33_), .Y(men_men_n161_));
  NA2        u145(.A(men_men_n161_), .B(men_men_n158_), .Y(men_men_n162_));
  NO3        u146(.A(men_men_n162_), .B(men_men_n155_), .C(men_men_n146_), .Y(men_men_n163_));
  NO2        u147(.A(men_men_n163_), .B(men_men_n143_), .Y(men_men_n164_));
  NO2        u148(.A(men_men_n140_), .B(men_men_n137_), .Y(men_men_n165_));
  NA2        u149(.A(men_men_n24_), .B(men_men_n18_), .Y(men_men_n166_));
  NA2        u150(.A(men_men_n24_), .B(men_men_n17_), .Y(men_men_n167_));
  NA3        u151(.A(men_men_n167_), .B(men_men_n166_), .C(men_men_n23_), .Y(men_men_n168_));
  AN2        u152(.A(men_men_n168_), .B(men_men_n141_), .Y(men_men_n169_));
  NA2        u153(.A(x8), .B(x0), .Y(men_men_n170_));
  NO2        u154(.A(men_men_n150_), .B(men_men_n24_), .Y(men_men_n171_));
  NO2        u155(.A(men_men_n123_), .B(x4), .Y(men_men_n172_));
  NA2        u156(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  AOI210     u157(.A0(men_men_n170_), .A1(men_men_n131_), .B0(men_men_n173_), .Y(men_men_n174_));
  NA2        u158(.A(x2), .B(x0), .Y(men_men_n175_));
  NA2        u159(.A(x4), .B(x1), .Y(men_men_n176_));
  NAi21      u160(.An(men_men_n121_), .B(men_men_n176_), .Y(men_men_n177_));
  NO3        u161(.A(men_men_n174_), .B(men_men_n169_), .C(men_men_n165_), .Y(men_men_n178_));
  NO2        u162(.A(men_men_n178_), .B(men_men_n41_), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n168_), .B(men_men_n74_), .Y(men_men_n180_));
  INV        u164(.A(men_men_n130_), .Y(men_men_n181_));
  NO2        u165(.A(men_men_n105_), .B(men_men_n17_), .Y(men_men_n182_));
  AOI210     u166(.A0(men_men_n33_), .A1(men_men_n90_), .B0(men_men_n182_), .Y(men_men_n183_));
  NO3        u167(.A(men_men_n183_), .B(men_men_n181_), .C(x7), .Y(men_men_n184_));
  NA3        u168(.A(men_men_n177_), .B(men_men_n181_), .C(men_men_n40_), .Y(men_men_n185_));
  OAI210     u169(.A0(men_men_n167_), .A1(men_men_n137_), .B0(men_men_n185_), .Y(men_men_n186_));
  NO3        u170(.A(men_men_n186_), .B(men_men_n184_), .C(men_men_n180_), .Y(men_men_n187_));
  NO2        u171(.A(men_men_n187_), .B(x3), .Y(men_men_n188_));
  NO3        u172(.A(men_men_n188_), .B(men_men_n179_), .C(men_men_n164_), .Y(men03));
  NO2        u173(.A(men_men_n46_), .B(x3), .Y(men_men_n190_));
  NO2        u174(.A(x6), .B(men_men_n24_), .Y(men_men_n191_));
  NO2        u175(.A(men_men_n52_), .B(x1), .Y(men_men_n192_));
  INV        u176(.A(men_men_n61_), .Y(men_men_n193_));
  OAI220     u177(.A0(men_men_n193_), .A1(men_men_n17_), .B0(men_men_n24_), .B1(men_men_n105_), .Y(men_men_n194_));
  NA2        u178(.A(men_men_n194_), .B(men_men_n190_), .Y(men_men_n195_));
  NA2        u179(.A(x6), .B(men_men_n24_), .Y(men_men_n196_));
  NO2        u180(.A(men_men_n18_), .B(x0), .Y(men_men_n197_));
  NA2        u181(.A(x3), .B(men_men_n17_), .Y(men_men_n198_));
  NO2        u182(.A(men_men_n198_), .B(men_men_n196_), .Y(men_men_n199_));
  NA2        u183(.A(x9), .B(men_men_n52_), .Y(men_men_n200_));
  NA2        u184(.A(men_men_n200_), .B(x4), .Y(men_men_n201_));
  NA2        u185(.A(men_men_n196_), .B(men_men_n79_), .Y(men_men_n202_));
  AOI210     u186(.A0(men_men_n24_), .A1(x3), .B0(men_men_n175_), .Y(men_men_n203_));
  AOI220     u187(.A0(men_men_n203_), .A1(men_men_n202_), .B0(men_men_n201_), .B1(men_men_n199_), .Y(men_men_n204_));
  NO2        u188(.A(x5), .B(x1), .Y(men_men_n205_));
  AOI220     u189(.A0(men_men_n205_), .A1(men_men_n17_), .B0(men_men_n102_), .B1(x5), .Y(men_men_n206_));
  NO2        u190(.A(men_men_n198_), .B(men_men_n166_), .Y(men_men_n207_));
  INV        u191(.A(men_men_n207_), .Y(men_men_n208_));
  OAI210     u192(.A0(men_men_n206_), .A1(men_men_n62_), .B0(men_men_n208_), .Y(men_men_n209_));
  NA2        u193(.A(men_men_n209_), .B(men_men_n46_), .Y(men_men_n210_));
  NA3        u194(.A(men_men_n210_), .B(men_men_n204_), .C(men_men_n195_), .Y(men_men_n211_));
  NO2        u195(.A(x3), .B(men_men_n17_), .Y(men_men_n212_));
  NO2        u196(.A(men_men_n212_), .B(x6), .Y(men_men_n213_));
  NOi21      u197(.An(men_men_n81_), .B(men_men_n213_), .Y(men_men_n214_));
  NA2        u198(.A(men_men_n60_), .B(men_men_n90_), .Y(men_men_n215_));
  NA3        u199(.A(men_men_n215_), .B(men_men_n212_), .C(x6), .Y(men_men_n216_));
  AOI210     u200(.A0(men_men_n216_), .A1(men_men_n214_), .B0(men_men_n150_), .Y(men_men_n217_));
  OR2        u201(.A(men_men_n217_), .B(men_men_n171_), .Y(men_men_n218_));
  NA2        u202(.A(men_men_n41_), .B(men_men_n52_), .Y(men_men_n219_));
  INV        u203(.A(men_men_n167_), .Y(men_men_n220_));
  NO2        u204(.A(men_men_n176_), .B(x6), .Y(men_men_n221_));
  AOI220     u205(.A0(men_men_n221_), .A1(men_men_n220_), .B0(men_men_n141_), .B1(men_men_n89_), .Y(men_men_n222_));
  NA2        u206(.A(x6), .B(men_men_n46_), .Y(men_men_n223_));
  OAI210     u207(.A0(men_men_n117_), .A1(men_men_n77_), .B0(x4), .Y(men_men_n224_));
  AOI210     u208(.A0(men_men_n224_), .A1(men_men_n223_), .B0(men_men_n76_), .Y(men_men_n225_));
  NO2        u209(.A(men_men_n60_), .B(x6), .Y(men_men_n226_));
  NO2        u210(.A(men_men_n156_), .B(men_men_n41_), .Y(men_men_n227_));
  OAI210     u211(.A0(men_men_n227_), .A1(men_men_n207_), .B0(men_men_n226_), .Y(men_men_n228_));
  NA2        u212(.A(men_men_n191_), .B(men_men_n135_), .Y(men_men_n229_));
  OAI210     u213(.A0(men_men_n90_), .A1(men_men_n34_), .B0(men_men_n65_), .Y(men_men_n230_));
  NA3        u214(.A(men_men_n230_), .B(men_men_n229_), .C(men_men_n228_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n225_), .B0(x2), .Y(men_men_n232_));
  NA3        u216(.A(men_men_n232_), .B(men_men_n222_), .C(men_men_n218_), .Y(men_men_n233_));
  AOI210     u217(.A0(men_men_n211_), .A1(x8), .B0(men_men_n233_), .Y(men_men_n234_));
  NO2        u218(.A(men_men_n90_), .B(x3), .Y(men_men_n235_));
  NA2        u219(.A(men_men_n405_), .B(men_men_n65_), .Y(men_men_n236_));
  NA2        u220(.A(men_men_n60_), .B(x6), .Y(men_men_n237_));
  NA3        u221(.A(men_men_n24_), .B(x3), .C(x2), .Y(men_men_n238_));
  INV        u222(.A(men_men_n237_), .Y(men_men_n239_));
  NA2        u223(.A(men_men_n41_), .B(men_men_n17_), .Y(men_men_n240_));
  NA2        u224(.A(men_men_n239_), .B(men_men_n121_), .Y(men_men_n241_));
  NA2        u225(.A(men_men_n198_), .B(x6), .Y(men_men_n242_));
  NA2        u226(.A(men_men_n242_), .B(men_men_n144_), .Y(men_men_n243_));
  NA4        u227(.A(men_men_n243_), .B(men_men_n241_), .C(men_men_n236_), .D(men_men_n150_), .Y(men_men_n244_));
  NA2        u228(.A(men_men_n191_), .B(men_men_n212_), .Y(men_men_n245_));
  INV        u229(.A(x6), .Y(men_men_n246_));
  NO2        u230(.A(men_men_n140_), .B(men_men_n18_), .Y(men_men_n247_));
  NAi21      u231(.An(men_men_n247_), .B(men_men_n238_), .Y(men_men_n248_));
  NAi21      u232(.An(x1), .B(x4), .Y(men_men_n249_));
  AOI210     u233(.A0(x3), .A1(x2), .B0(men_men_n46_), .Y(men_men_n250_));
  OAI210     u234(.A0(men_men_n140_), .A1(x3), .B0(men_men_n250_), .Y(men_men_n251_));
  AOI220     u235(.A0(men_men_n251_), .A1(men_men_n249_), .B0(men_men_n248_), .B1(men_men_n246_), .Y(men_men_n252_));
  NA2        u236(.A(men_men_n252_), .B(men_men_n245_), .Y(men_men_n253_));
  NO2        u237(.A(men_men_n404_), .B(men_men_n245_), .Y(men_men_n254_));
  NO3        u238(.A(x9), .B(x6), .C(x0), .Y(men_men_n255_));
  NA2        u239(.A(men_men_n105_), .B(men_men_n24_), .Y(men_men_n256_));
  NA2        u240(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  OAI220     u241(.A0(men_men_n257_), .A1(men_men_n41_), .B0(men_men_n172_), .B1(men_men_n44_), .Y(men_men_n258_));
  OAI210     u242(.A0(men_men_n258_), .A1(men_men_n254_), .B0(men_men_n253_), .Y(men_men_n259_));
  NO2        u243(.A(x3), .B(men_men_n196_), .Y(men_men_n260_));
  NA2        u244(.A(x4), .B(x0), .Y(men_men_n261_));
  NO2        u245(.A(men_men_n71_), .B(x6), .Y(men_men_n262_));
  AOI210     u246(.A0(men_men_n260_), .A1(men_men_n40_), .B0(men_men_n262_), .Y(men_men_n263_));
  AOI210     u247(.A0(men_men_n263_), .A1(men_men_n259_), .B0(x8), .Y(men_men_n264_));
  NA2        u248(.A(x0), .B(men_men_n20_), .Y(men_men_n265_));
  NO2        u249(.A(men_men_n265_), .B(men_men_n219_), .Y(men_men_n266_));
  NO3        u250(.A(men_men_n266_), .B(men_men_n264_), .C(men_men_n244_), .Y(men_men_n267_));
  NO2        u251(.A(men_men_n159_), .B(x1), .Y(men_men_n268_));
  NO3        u252(.A(men_men_n268_), .B(x3), .C(men_men_n34_), .Y(men_men_n269_));
  NA2        u253(.A(men_men_n269_), .B(x2), .Y(men_men_n270_));
  OAI210     u254(.A0(x0), .A1(x6), .B0(men_men_n42_), .Y(men_men_n271_));
  AOI210     u255(.A0(men_men_n271_), .A1(men_men_n270_), .B0(men_men_n181_), .Y(men_men_n272_));
  NA3        u256(.A(x0), .B(men_men_n205_), .C(men_men_n38_), .Y(men_men_n273_));
  AOI210     u257(.A0(men_men_n34_), .A1(men_men_n52_), .B0(x0), .Y(men_men_n274_));
  NA3        u258(.A(men_men_n274_), .B(men_men_n157_), .C(men_men_n31_), .Y(men_men_n275_));
  NA2        u259(.A(x3), .B(x2), .Y(men_men_n276_));
  AOI220     u260(.A0(men_men_n276_), .A1(men_men_n219_), .B0(men_men_n275_), .B1(men_men_n273_), .Y(men_men_n277_));
  NAi21      u261(.An(x4), .B(x0), .Y(men_men_n278_));
  NO3        u262(.A(men_men_n278_), .B(men_men_n42_), .C(x2), .Y(men_men_n279_));
  OAI210     u263(.A0(x6), .A1(men_men_n18_), .B0(men_men_n279_), .Y(men_men_n280_));
  OAI220     u264(.A0(men_men_n23_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n281_));
  NO2        u265(.A(x9), .B(x8), .Y(men_men_n282_));
  NA3        u266(.A(men_men_n282_), .B(men_men_n34_), .C(men_men_n52_), .Y(men_men_n283_));
  OAI210     u267(.A0(men_men_n274_), .A1(x0), .B0(men_men_n283_), .Y(men_men_n284_));
  AOI220     u268(.A0(men_men_n284_), .A1(men_men_n80_), .B0(men_men_n281_), .B1(men_men_n30_), .Y(men_men_n285_));
  AOI210     u269(.A0(men_men_n285_), .A1(men_men_n280_), .B0(men_men_n24_), .Y(men_men_n286_));
  INV        u270(.A(men_men_n207_), .Y(men_men_n287_));
  NA2        u271(.A(men_men_n34_), .B(men_men_n41_), .Y(men_men_n288_));
  OR2        u272(.A(men_men_n288_), .B(men_men_n261_), .Y(men_men_n289_));
  OAI220     u273(.A0(men_men_n289_), .A1(men_men_n156_), .B0(men_men_n223_), .B1(men_men_n287_), .Y(men_men_n290_));
  NO4        u274(.A(men_men_n290_), .B(men_men_n286_), .C(men_men_n277_), .D(men_men_n272_), .Y(men_men_n291_));
  OAI210     u275(.A0(men_men_n267_), .A1(men_men_n234_), .B0(men_men_n291_), .Y(men04));
  NA2        u276(.A(men_men_n255_), .B(men_men_n82_), .Y(men_men_n293_));
  NA2        u277(.A(men_men_n52_), .B(men_men_n235_), .Y(men_men_n294_));
  NA3        u278(.A(men_men_n88_), .B(x6), .C(men_men_n294_), .Y(men_men_n295_));
  NA2        u279(.A(men_men_n295_), .B(x6), .Y(men_men_n296_));
  NO2        u280(.A(men_men_n200_), .B(men_men_n111_), .Y(men_men_n297_));
  INV        u281(.A(men_men_n297_), .Y(men_men_n298_));
  OAI210     u282(.A0(men_men_n404_), .A1(x6), .B0(men_men_n288_), .Y(men_men_n299_));
  AOI210     u283(.A0(men_men_n148_), .A1(men_men_n61_), .B0(men_men_n299_), .Y(men_men_n300_));
  NA2        u284(.A(men_men_n300_), .B(men_men_n298_), .Y(men_men_n301_));
  AOI210     u285(.A0(men_men_n301_), .A1(x4), .B0(x7), .Y(men_men_n302_));
  XO2        u286(.A(x4), .B(x0), .Y(men_men_n303_));
  OAI210     u287(.A0(men_men_n303_), .A1(men_men_n115_), .B0(men_men_n249_), .Y(men_men_n304_));
  NA2        u288(.A(men_men_n304_), .B(x8), .Y(men_men_n305_));
  NO2        u289(.A(men_men_n305_), .B(x3), .Y(men_men_n306_));
  INV        u290(.A(men_men_n91_), .Y(men_men_n307_));
  NO2        u291(.A(men_men_n90_), .B(x4), .Y(men_men_n308_));
  AOI220     u292(.A0(men_men_n308_), .A1(men_men_n42_), .B0(men_men_n125_), .B1(men_men_n307_), .Y(men_men_n309_));
  NO3        u293(.A(men_men_n303_), .B(men_men_n159_), .C(x2), .Y(men_men_n310_));
  NO3        u294(.A(men_men_n215_), .B(men_men_n27_), .C(men_men_n23_), .Y(men_men_n311_));
  NO2        u295(.A(men_men_n311_), .B(men_men_n310_), .Y(men_men_n312_));
  NA3        u296(.A(men_men_n312_), .B(men_men_n309_), .C(x6), .Y(men_men_n313_));
  OAI220     u297(.A0(men_men_n278_), .A1(men_men_n88_), .B0(men_men_n175_), .B1(men_men_n90_), .Y(men_men_n314_));
  NO2        u298(.A(men_men_n41_), .B(x0), .Y(men_men_n315_));
  OR2        u299(.A(men_men_n308_), .B(men_men_n315_), .Y(men_men_n316_));
  NO2        u300(.A(men_men_n148_), .B(men_men_n105_), .Y(men_men_n317_));
  AOI220     u301(.A0(men_men_n317_), .A1(men_men_n316_), .B0(men_men_n314_), .B1(men_men_n59_), .Y(men_men_n318_));
  INV        u302(.A(men_men_n318_), .Y(men_men_n319_));
  OAI220     u303(.A0(men_men_n319_), .A1(x6), .B0(men_men_n313_), .B1(men_men_n306_), .Y(men_men_n320_));
  OAI210     u304(.A0(men_men_n61_), .A1(men_men_n46_), .B0(men_men_n40_), .Y(men_men_n321_));
  OAI210     u305(.A0(men_men_n321_), .A1(men_men_n90_), .B0(men_men_n289_), .Y(men_men_n322_));
  AOI210     u306(.A0(men_men_n322_), .A1(men_men_n18_), .B0(men_men_n150_), .Y(men_men_n323_));
  AO220      u307(.A0(men_men_n323_), .A1(men_men_n320_), .B0(men_men_n302_), .B1(men_men_n296_), .Y(men_men_n324_));
  NA2        u308(.A(men_men_n308_), .B(x0), .Y(men_men_n325_));
  NO2        u309(.A(men_men_n325_), .B(men_men_n41_), .Y(men_men_n326_));
  INV        u310(.A(men_men_n326_), .Y(men_men_n327_));
  NA3        u311(.A(men_men_n327_), .B(men_men_n324_), .C(men_men_n293_), .Y(men_men_n328_));
  NA3        u312(.A(x7), .B(x3), .C(x0), .Y(men_men_n329_));
  NA2        u313(.A(x3), .B(x0), .Y(men_men_n330_));
  OAI220     u314(.A0(men_men_n330_), .A1(men_men_n200_), .B0(men_men_n329_), .B1(men_men_n307_), .Y(men_men_n331_));
  INV        u315(.A(men_men_n331_), .Y(men_men_n332_));
  NO2        u316(.A(men_men_n332_), .B(men_men_n24_), .Y(men_men_n333_));
  NA3        u317(.A(men_men_n119_), .B(x3), .C(x0), .Y(men_men_n334_));
  OAI210     u318(.A0(men_men_n190_), .A1(men_men_n66_), .B0(men_men_n197_), .Y(men_men_n335_));
  NA3        u319(.A(men_men_n192_), .B(men_men_n212_), .C(x8), .Y(men_men_n336_));
  AOI210     u320(.A0(men_men_n336_), .A1(men_men_n335_), .B0(men_men_n24_), .Y(men_men_n337_));
  AOI210     u321(.A0(men_men_n118_), .A1(men_men_n116_), .B0(men_men_n40_), .Y(men_men_n338_));
  NOi31      u322(.An(men_men_n338_), .B(men_men_n315_), .C(men_men_n176_), .Y(men_men_n339_));
  OAI210     u323(.A0(men_men_n339_), .A1(men_men_n337_), .B0(men_men_n147_), .Y(men_men_n340_));
  NAi31      u324(.An(men_men_n48_), .B(men_men_n268_), .C(men_men_n171_), .Y(men_men_n341_));
  NA3        u325(.A(men_men_n341_), .B(men_men_n340_), .C(men_men_n334_), .Y(men_men_n342_));
  OAI210     u326(.A0(men_men_n342_), .A1(men_men_n333_), .B0(x6), .Y(men_men_n343_));
  INV        u327(.A(men_men_n136_), .Y(men_men_n344_));
  NA3        u328(.A(men_men_n53_), .B(men_men_n36_), .C(men_men_n30_), .Y(men_men_n345_));
  AOI220     u329(.A0(men_men_n345_), .A1(men_men_n344_), .B0(men_men_n38_), .B1(men_men_n31_), .Y(men_men_n346_));
  AOI210     u330(.A0(men_men_n127_), .A1(men_men_n405_), .B0(x1), .Y(men_men_n347_));
  INV        u331(.A(men_men_n347_), .Y(men_men_n348_));
  NAi31      u332(.An(x2), .B(x8), .C(x0), .Y(men_men_n349_));
  NA2        u333(.A(men_men_n406_), .B(x9), .Y(men_men_n350_));
  NO4        u334(.A(men_men_n126_), .B(men_men_n278_), .C(x9), .D(x2), .Y(men_men_n351_));
  NOi21      u335(.An(men_men_n124_), .B(men_men_n175_), .Y(men_men_n352_));
  NO3        u336(.A(men_men_n352_), .B(men_men_n351_), .C(men_men_n18_), .Y(men_men_n353_));
  NO3        u337(.A(x9), .B(men_men_n150_), .C(x0), .Y(men_men_n354_));
  NA2        u338(.A(men_men_n354_), .B(men_men_n235_), .Y(men_men_n355_));
  NA4        u339(.A(men_men_n355_), .B(men_men_n353_), .C(men_men_n350_), .D(men_men_n48_), .Y(men_men_n356_));
  OAI210     u340(.A0(men_men_n348_), .A1(men_men_n346_), .B0(men_men_n356_), .Y(men_men_n357_));
  AOI210     u341(.A0(men_men_n36_), .A1(x9), .B0(men_men_n134_), .Y(men_men_n358_));
  NO3        u342(.A(men_men_n358_), .B(men_men_n124_), .C(men_men_n41_), .Y(men_men_n359_));
  AOI210     u343(.A0(men_men_n249_), .A1(men_men_n58_), .B0(men_men_n123_), .Y(men_men_n360_));
  NO2        u344(.A(men_men_n360_), .B(x3), .Y(men_men_n361_));
  NO3        u345(.A(men_men_n361_), .B(men_men_n359_), .C(x2), .Y(men_men_n362_));
  OAI220     u346(.A0(men_men_n303_), .A1(men_men_n282_), .B0(men_men_n278_), .B1(men_men_n41_), .Y(men_men_n363_));
  AOI210     u347(.A0(x9), .A1(men_men_n46_), .B0(men_men_n329_), .Y(men_men_n364_));
  AOI220     u348(.A0(men_men_n364_), .A1(men_men_n90_), .B0(men_men_n363_), .B1(men_men_n150_), .Y(men_men_n365_));
  NO2        u349(.A(men_men_n365_), .B(men_men_n52_), .Y(men_men_n366_));
  NO2        u350(.A(men_men_n366_), .B(men_men_n362_), .Y(men_men_n367_));
  AOI210     u351(.A0(men_men_n367_), .A1(men_men_n357_), .B0(men_men_n24_), .Y(men_men_n368_));
  NA4        u352(.A(men_men_n30_), .B(men_men_n90_), .C(x2), .D(men_men_n17_), .Y(men_men_n369_));
  NO3        u353(.A(men_men_n60_), .B(x4), .C(x1), .Y(men_men_n370_));
  NO3        u354(.A(men_men_n66_), .B(men_men_n18_), .C(x0), .Y(men_men_n371_));
  AOI220     u355(.A0(men_men_n371_), .A1(men_men_n250_), .B0(men_men_n370_), .B1(men_men_n338_), .Y(men_men_n372_));
  NO2        u356(.A(men_men_n372_), .B(men_men_n102_), .Y(men_men_n373_));
  NA2        u357(.A(men_men_n373_), .B(x7), .Y(men_men_n374_));
  NA2        u358(.A(men_men_n215_), .B(x7), .Y(men_men_n375_));
  NA3        u359(.A(men_men_n375_), .B(men_men_n149_), .C(men_men_n135_), .Y(men_men_n376_));
  NA3        u360(.A(men_men_n376_), .B(men_men_n374_), .C(men_men_n369_), .Y(men_men_n377_));
  OAI210     u361(.A0(men_men_n377_), .A1(men_men_n368_), .B0(men_men_n34_), .Y(men_men_n378_));
  NO2        u362(.A(men_men_n354_), .B(men_men_n197_), .Y(men_men_n379_));
  NO4        u363(.A(men_men_n379_), .B(men_men_n76_), .C(x4), .D(men_men_n52_), .Y(men_men_n380_));
  NA2        u364(.A(men_men_n240_), .B(men_men_n21_), .Y(men_men_n381_));
  NO2        u365(.A(men_men_n156_), .B(men_men_n136_), .Y(men_men_n382_));
  NA2        u366(.A(men_men_n382_), .B(men_men_n381_), .Y(men_men_n383_));
  AOI210     u367(.A0(men_men_n383_), .A1(men_men_n161_), .B0(men_men_n27_), .Y(men_men_n384_));
  AOI220     u368(.A0(men_men_n315_), .A1(men_men_n90_), .B0(men_men_n148_), .B1(men_men_n192_), .Y(men_men_n385_));
  NA3        u369(.A(men_men_n385_), .B(men_men_n349_), .C(men_men_n88_), .Y(men_men_n386_));
  NA2        u370(.A(men_men_n386_), .B(men_men_n171_), .Y(men_men_n387_));
  OAI220     u371(.A0(x3), .A1(men_men_n67_), .B0(men_men_n156_), .B1(men_men_n41_), .Y(men_men_n388_));
  NA2        u372(.A(x3), .B(men_men_n52_), .Y(men_men_n389_));
  AOI210     u373(.A0(men_men_n160_), .A1(men_men_n26_), .B0(men_men_n71_), .Y(men_men_n390_));
  OAI210     u374(.A0(men_men_n147_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n391_));
  NO2        u375(.A(x3), .B(men_men_n52_), .Y(men_men_n392_));
  AOI210     u376(.A0(men_men_n392_), .A1(men_men_n391_), .B0(men_men_n390_), .Y(men_men_n393_));
  OAI210     u377(.A0(men_men_n151_), .A1(men_men_n389_), .B0(men_men_n393_), .Y(men_men_n394_));
  AOI220     u378(.A0(men_men_n394_), .A1(x0), .B0(men_men_n388_), .B1(men_men_n136_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n395_), .A1(men_men_n387_), .B0(men_men_n223_), .Y(men_men_n396_));
  NA2        u380(.A(x9), .B(x5), .Y(men_men_n397_));
  NO4        u381(.A(men_men_n105_), .B(men_men_n397_), .C(men_men_n58_), .D(men_men_n31_), .Y(men_men_n398_));
  NO4        u382(.A(men_men_n398_), .B(men_men_n396_), .C(men_men_n384_), .D(men_men_n380_), .Y(men_men_n399_));
  NA3        u383(.A(men_men_n399_), .B(men_men_n378_), .C(men_men_n343_), .Y(men_men_n400_));
  AOI210     u384(.A0(men_men_n328_), .A1(men_men_n24_), .B0(men_men_n400_), .Y(men05));
  INV        u385(.A(x2), .Y(men_men_n404_));
  INV        u386(.A(x4), .Y(men_men_n405_));
  INV        u387(.A(x2), .Y(men_men_n406_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule