//Benchmark atmr_9sym_175_0.0313

module atmr_9sym(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, z0);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;
 output z0;
 wire ori_ori_n11_, ori_ori_n12_, ori_ori_n13_, ori_ori_n14_, ori_ori_n15_, ori_ori_n16_, ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n167_, mai_mai_n11_, mai_mai_n12_, mai_mai_n13_, mai_mai_n14_, mai_mai_n15_, mai_mai_n16_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n174_, men_men_n11_, men_men_n12_, men_men_n13_, men_men_n14_, men_men_n15_, men_men_n16_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n172_, men_men_n173_, men_men_n174_, ori00, mai00, men00;
  INV        o000(.A(i_3_), .Y(ori_ori_n11_));
  INV        o001(.A(i_6_), .Y(ori_ori_n12_));
  NA2        o002(.A(i_4_), .B(ori_ori_n12_), .Y(ori_ori_n13_));
  INV        o003(.A(i_5_), .Y(ori_ori_n14_));
  NOi21      o004(.An(i_3_), .B(i_7_), .Y(ori_ori_n15_));
  NA3        o005(.A(ori_ori_n15_), .B(i_0_), .C(ori_ori_n14_), .Y(ori_ori_n16_));
  INV        o006(.A(i_0_), .Y(ori_ori_n17_));
  NOi21      o007(.An(i_1_), .B(i_3_), .Y(ori_ori_n18_));
  NO2        o008(.A(ori_ori_n16_), .B(ori_ori_n13_), .Y(ori_ori_n19_));
  INV        o009(.A(i_4_), .Y(ori_ori_n20_));
  NA2        o010(.A(i_0_), .B(ori_ori_n20_), .Y(ori_ori_n21_));
  INV        o011(.A(i_7_), .Y(ori_ori_n22_));
  NA3        o012(.A(i_6_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n23_));
  NOi21      o013(.An(i_8_), .B(i_6_), .Y(ori_ori_n24_));
  NOi21      o014(.An(i_1_), .B(i_8_), .Y(ori_ori_n25_));
  AOI220     o015(.A0(ori_ori_n25_), .A1(i_2_), .B0(ori_ori_n24_), .B1(i_5_), .Y(ori_ori_n26_));
  AOI210     o016(.A0(ori_ori_n26_), .A1(ori_ori_n23_), .B0(ori_ori_n21_), .Y(ori_ori_n27_));
  AOI210     o017(.A0(ori_ori_n27_), .A1(ori_ori_n11_), .B0(ori_ori_n19_), .Y(ori_ori_n28_));
  NA2        o018(.A(i_0_), .B(ori_ori_n14_), .Y(ori_ori_n29_));
  NA2        o019(.A(ori_ori_n17_), .B(i_5_), .Y(ori_ori_n30_));
  NO2        o020(.A(i_2_), .B(i_4_), .Y(ori_ori_n31_));
  NA3        o021(.A(ori_ori_n31_), .B(i_6_), .C(i_8_), .Y(ori_ori_n32_));
  AOI210     o022(.A0(ori_ori_n30_), .A1(ori_ori_n29_), .B0(ori_ori_n32_), .Y(ori_ori_n33_));
  INV        o023(.A(i_2_), .Y(ori_ori_n34_));
  NOi21      o024(.An(i_5_), .B(i_0_), .Y(ori_ori_n35_));
  NOi21      o025(.An(i_6_), .B(i_8_), .Y(ori_ori_n36_));
  NOi21      o026(.An(i_7_), .B(i_1_), .Y(ori_ori_n37_));
  NOi21      o027(.An(i_5_), .B(i_6_), .Y(ori_ori_n38_));
  AOI220     o028(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n36_), .B1(ori_ori_n35_), .Y(ori_ori_n39_));
  NO3        o029(.A(ori_ori_n39_), .B(ori_ori_n34_), .C(i_4_), .Y(ori_ori_n40_));
  NOi21      o030(.An(i_0_), .B(i_4_), .Y(ori_ori_n41_));
  XO2        o031(.A(i_1_), .B(i_3_), .Y(ori_ori_n42_));
  NOi21      o032(.An(i_7_), .B(i_5_), .Y(ori_ori_n43_));
  AN3        o033(.A(ori_ori_n43_), .B(ori_ori_n42_), .C(ori_ori_n41_), .Y(ori_ori_n44_));
  INV        o034(.A(i_1_), .Y(ori_ori_n45_));
  NOi21      o035(.An(i_3_), .B(i_0_), .Y(ori_ori_n46_));
  NA2        o036(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o037(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n48_));
  NO4        o038(.A(ori_ori_n48_), .B(ori_ori_n44_), .C(ori_ori_n40_), .D(ori_ori_n33_), .Y(ori_ori_n49_));
  NA2        o039(.A(i_1_), .B(ori_ori_n11_), .Y(ori_ori_n50_));
  NOi21      o040(.An(i_4_), .B(i_0_), .Y(ori_ori_n51_));
  NO2        o041(.A(ori_ori_n24_), .B(ori_ori_n15_), .Y(ori_ori_n52_));
  NA2        o042(.A(i_1_), .B(ori_ori_n14_), .Y(ori_ori_n53_));
  NOi21      o043(.An(i_2_), .B(i_8_), .Y(ori_ori_n54_));
  NO3        o044(.A(ori_ori_n54_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori_ori_n55_));
  NO3        o045(.A(ori_ori_n55_), .B(ori_ori_n53_), .C(ori_ori_n52_), .Y(ori_ori_n56_));
  INV        o046(.A(ori_ori_n56_), .Y(ori_ori_n57_));
  NOi31      o047(.An(i_2_), .B(i_1_), .C(i_3_), .Y(ori_ori_n58_));
  NOi21      o048(.An(i_4_), .B(i_3_), .Y(ori_ori_n59_));
  NOi21      o049(.An(i_1_), .B(i_4_), .Y(ori_ori_n60_));
  AN2        o050(.A(i_8_), .B(i_7_), .Y(ori_ori_n61_));
  INV        o051(.A(ori_ori_n61_), .Y(ori_ori_n62_));
  NOi21      o052(.An(i_8_), .B(i_7_), .Y(ori_ori_n63_));
  NA3        o053(.A(ori_ori_n63_), .B(ori_ori_n59_), .C(i_6_), .Y(ori_ori_n64_));
  OAI210     o054(.A0(ori_ori_n62_), .A1(ori_ori_n53_), .B0(ori_ori_n64_), .Y(ori_ori_n65_));
  AOI220     o055(.A0(ori_ori_n65_), .A1(ori_ori_n34_), .B0(ori_ori_n54_), .B1(ori_ori_n38_), .Y(ori_ori_n66_));
  NA4        o056(.A(ori_ori_n66_), .B(ori_ori_n57_), .C(ori_ori_n49_), .D(ori_ori_n28_), .Y(ori_ori_n67_));
  NA2        o057(.A(i_8_), .B(ori_ori_n22_), .Y(ori_ori_n68_));
  AOI220     o058(.A0(ori_ori_n46_), .A1(i_1_), .B0(ori_ori_n42_), .B1(i_2_), .Y(ori_ori_n69_));
  NOi21      o059(.An(i_1_), .B(i_2_), .Y(ori_ori_n70_));
  NO2        o060(.A(ori_ori_n69_), .B(ori_ori_n68_), .Y(ori_ori_n71_));
  NA2        o061(.A(ori_ori_n71_), .B(ori_ori_n14_), .Y(ori_ori_n72_));
  NA3        o062(.A(ori_ori_n63_), .B(i_2_), .C(ori_ori_n12_), .Y(ori_ori_n73_));
  NA2        o063(.A(ori_ori_n25_), .B(ori_ori_n14_), .Y(ori_ori_n74_));
  NA2        o064(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  NOi32      o065(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(ori_ori_n76_));
  NA2        o066(.A(ori_ori_n76_), .B(i_3_), .Y(ori_ori_n77_));
  NA2        o067(.A(ori_ori_n18_), .B(i_6_), .Y(ori_ori_n78_));
  NA2        o068(.A(ori_ori_n78_), .B(ori_ori_n77_), .Y(ori_ori_n79_));
  INV        o069(.A(i_0_), .Y(ori_ori_n80_));
  AOI220     o070(.A0(ori_ori_n80_), .A1(ori_ori_n79_), .B0(ori_ori_n75_), .B1(ori_ori_n59_), .Y(ori_ori_n81_));
  NA2        o071(.A(ori_ori_n81_), .B(ori_ori_n72_), .Y(ori_ori_n82_));
  NA2        o072(.A(ori_ori_n36_), .B(ori_ori_n35_), .Y(ori_ori_n83_));
  NOi21      o073(.An(i_7_), .B(i_8_), .Y(ori_ori_n84_));
  NOi21      o074(.An(i_6_), .B(i_5_), .Y(ori_ori_n85_));
  AOI210     o075(.A0(ori_ori_n84_), .A1(ori_ori_n12_), .B0(ori_ori_n85_), .Y(ori_ori_n86_));
  OAI210     o076(.A0(ori_ori_n86_), .A1(ori_ori_n11_), .B0(ori_ori_n83_), .Y(ori_ori_n87_));
  NA2        o077(.A(ori_ori_n87_), .B(ori_ori_n70_), .Y(ori_ori_n88_));
  NA3        o078(.A(ori_ori_n24_), .B(i_2_), .C(ori_ori_n14_), .Y(ori_ori_n89_));
  AOI210     o079(.A0(ori_ori_n21_), .A1(ori_ori_n50_), .B0(ori_ori_n89_), .Y(ori_ori_n90_));
  AOI220     o080(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n18_), .B1(ori_ori_n34_), .Y(ori_ori_n91_));
  NA3        o081(.A(ori_ori_n20_), .B(i_5_), .C(i_7_), .Y(ori_ori_n92_));
  NO2        o082(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NO2        o083(.A(ori_ori_n93_), .B(ori_ori_n90_), .Y(ori_ori_n94_));
  NA3        o084(.A(ori_ori_n63_), .B(ori_ori_n34_), .C(i_3_), .Y(ori_ori_n95_));
  NA2        o085(.A(ori_ori_n45_), .B(i_6_), .Y(ori_ori_n96_));
  AOI210     o086(.A0(ori_ori_n96_), .A1(ori_ori_n21_), .B0(ori_ori_n95_), .Y(ori_ori_n97_));
  NOi21      o087(.An(i_2_), .B(i_1_), .Y(ori_ori_n98_));
  AN3        o088(.A(ori_ori_n84_), .B(ori_ori_n98_), .C(ori_ori_n51_), .Y(ori_ori_n99_));
  NAi21      o089(.An(i_6_), .B(i_0_), .Y(ori_ori_n100_));
  NA3        o090(.A(ori_ori_n60_), .B(i_5_), .C(ori_ori_n22_), .Y(ori_ori_n101_));
  NOi21      o091(.An(i_4_), .B(i_6_), .Y(ori_ori_n102_));
  NOi21      o092(.An(i_5_), .B(i_3_), .Y(ori_ori_n103_));
  NA3        o093(.A(ori_ori_n103_), .B(ori_ori_n70_), .C(ori_ori_n102_), .Y(ori_ori_n104_));
  OAI210     o094(.A0(ori_ori_n101_), .A1(ori_ori_n100_), .B0(ori_ori_n104_), .Y(ori_ori_n105_));
  NA2        o095(.A(ori_ori_n70_), .B(ori_ori_n36_), .Y(ori_ori_n106_));
  NO3        o096(.A(ori_ori_n105_), .B(ori_ori_n99_), .C(ori_ori_n97_), .Y(ori_ori_n107_));
  NOi31      o097(.An(ori_ori_n51_), .B(ori_ori_n167_), .C(i_2_), .Y(ori_ori_n108_));
  NA2        o098(.A(ori_ori_n63_), .B(ori_ori_n12_), .Y(ori_ori_n109_));
  NA2        o099(.A(ori_ori_n36_), .B(ori_ori_n14_), .Y(ori_ori_n110_));
  NOi21      o100(.An(i_3_), .B(i_1_), .Y(ori_ori_n111_));
  NA2        o101(.A(ori_ori_n111_), .B(i_4_), .Y(ori_ori_n112_));
  AOI210     o102(.A0(ori_ori_n110_), .A1(ori_ori_n109_), .B0(ori_ori_n112_), .Y(ori_ori_n113_));
  NOi31      o103(.An(ori_ori_n46_), .B(i_5_), .C(ori_ori_n34_), .Y(ori_ori_n114_));
  NO3        o104(.A(ori_ori_n114_), .B(ori_ori_n113_), .C(ori_ori_n108_), .Y(ori_ori_n115_));
  NA4        o105(.A(ori_ori_n115_), .B(ori_ori_n107_), .C(ori_ori_n94_), .D(ori_ori_n88_), .Y(ori_ori_n116_));
  NA2        o106(.A(ori_ori_n54_), .B(ori_ori_n15_), .Y(ori_ori_n117_));
  NOi31      o107(.An(i_6_), .B(i_1_), .C(i_8_), .Y(ori_ori_n118_));
  NOi31      o108(.An(i_5_), .B(i_2_), .C(i_6_), .Y(ori_ori_n119_));
  OAI210     o109(.A0(ori_ori_n119_), .A1(ori_ori_n118_), .B0(i_7_), .Y(ori_ori_n120_));
  NA2        o110(.A(ori_ori_n36_), .B(ori_ori_n14_), .Y(ori_ori_n121_));
  NA4        o111(.A(ori_ori_n121_), .B(ori_ori_n120_), .C(ori_ori_n117_), .D(ori_ori_n106_), .Y(ori_ori_n122_));
  NA2        o112(.A(ori_ori_n122_), .B(ori_ori_n41_), .Y(ori_ori_n123_));
  NA2        o113(.A(ori_ori_n59_), .B(ori_ori_n37_), .Y(ori_ori_n124_));
  AOI210     o114(.A0(ori_ori_n124_), .A1(ori_ori_n73_), .B0(ori_ori_n30_), .Y(ori_ori_n125_));
  NA3        o115(.A(ori_ori_n61_), .B(ori_ori_n98_), .C(ori_ori_n12_), .Y(ori_ori_n126_));
  NAi31      o116(.An(ori_ori_n100_), .B(ori_ori_n84_), .C(ori_ori_n98_), .Y(ori_ori_n127_));
  NA3        o117(.A(ori_ori_n63_), .B(ori_ori_n58_), .C(i_6_), .Y(ori_ori_n128_));
  NA3        o118(.A(ori_ori_n128_), .B(ori_ori_n127_), .C(ori_ori_n126_), .Y(ori_ori_n129_));
  NOi21      o119(.An(i_0_), .B(i_2_), .Y(ori_ori_n130_));
  NA3        o120(.A(ori_ori_n130_), .B(ori_ori_n37_), .C(ori_ori_n102_), .Y(ori_ori_n131_));
  NOi32      o121(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(ori_ori_n132_));
  NA2        o122(.A(ori_ori_n132_), .B(ori_ori_n118_), .Y(ori_ori_n133_));
  NA3        o123(.A(ori_ori_n130_), .B(ori_ori_n59_), .C(ori_ori_n36_), .Y(ori_ori_n134_));
  NA3        o124(.A(ori_ori_n134_), .B(ori_ori_n133_), .C(ori_ori_n131_), .Y(ori_ori_n135_));
  NA4        o125(.A(ori_ori_n58_), .B(i_6_), .C(ori_ori_n14_), .D(i_7_), .Y(ori_ori_n136_));
  NA4        o126(.A(ori_ori_n60_), .B(ori_ori_n38_), .C(ori_ori_n17_), .D(i_8_), .Y(ori_ori_n137_));
  NA4        o127(.A(ori_ori_n60_), .B(ori_ori_n46_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n138_));
  NA3        o128(.A(ori_ori_n138_), .B(ori_ori_n137_), .C(ori_ori_n136_), .Y(ori_ori_n139_));
  NO4        o129(.A(ori_ori_n139_), .B(ori_ori_n135_), .C(ori_ori_n129_), .D(ori_ori_n125_), .Y(ori_ori_n140_));
  INV        o130(.A(i_2_), .Y(ori_ori_n141_));
  AOI220     o131(.A0(ori_ori_n141_), .A1(ori_ori_n84_), .B0(ori_ori_n61_), .B1(ori_ori_n31_), .Y(ori_ori_n142_));
  NO2        o132(.A(ori_ori_n142_), .B(ori_ori_n96_), .Y(ori_ori_n143_));
  NO4        o133(.A(i_2_), .B(ori_ori_n20_), .C(ori_ori_n11_), .D(ori_ori_n14_), .Y(ori_ori_n144_));
  NA2        o134(.A(i_2_), .B(i_4_), .Y(ori_ori_n145_));
  INV        o135(.A(ori_ori_n145_), .Y(ori_ori_n146_));
  NO2        o136(.A(i_8_), .B(i_7_), .Y(ori_ori_n147_));
  OA210      o137(.A0(ori_ori_n146_), .A1(ori_ori_n144_), .B0(ori_ori_n147_), .Y(ori_ori_n148_));
  NA4        o138(.A(ori_ori_n111_), .B(i_0_), .C(i_5_), .D(ori_ori_n22_), .Y(ori_ori_n149_));
  NO2        o139(.A(ori_ori_n149_), .B(i_4_), .Y(ori_ori_n150_));
  NO3        o140(.A(ori_ori_n150_), .B(ori_ori_n148_), .C(ori_ori_n143_), .Y(ori_ori_n151_));
  NA2        o141(.A(ori_ori_n84_), .B(ori_ori_n12_), .Y(ori_ori_n152_));
  NA3        o142(.A(i_2_), .B(i_1_), .C(ori_ori_n14_), .Y(ori_ori_n153_));
  NA2        o143(.A(ori_ori_n51_), .B(i_3_), .Y(ori_ori_n154_));
  AOI210     o144(.A0(ori_ori_n154_), .A1(ori_ori_n153_), .B0(ori_ori_n152_), .Y(ori_ori_n155_));
  NA3        o145(.A(ori_ori_n130_), .B(ori_ori_n63_), .C(ori_ori_n102_), .Y(ori_ori_n156_));
  OAI210     o146(.A0(ori_ori_n95_), .A1(ori_ori_n30_), .B0(ori_ori_n156_), .Y(ori_ori_n157_));
  NA4        o147(.A(ori_ori_n103_), .B(ori_ori_n61_), .C(ori_ori_n45_), .D(ori_ori_n20_), .Y(ori_ori_n158_));
  NOi31      o148(.An(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n159_));
  OAI210     o149(.A0(ori_ori_n132_), .A1(ori_ori_n76_), .B0(ori_ori_n159_), .Y(ori_ori_n160_));
  NA2        o150(.A(ori_ori_n160_), .B(ori_ori_n158_), .Y(ori_ori_n161_));
  NO3        o151(.A(ori_ori_n161_), .B(ori_ori_n157_), .C(ori_ori_n155_), .Y(ori_ori_n162_));
  NA4        o152(.A(ori_ori_n162_), .B(ori_ori_n151_), .C(ori_ori_n140_), .D(ori_ori_n123_), .Y(ori_ori_n163_));
  OR4        o153(.A(ori_ori_n163_), .B(ori_ori_n116_), .C(ori_ori_n82_), .D(ori_ori_n67_), .Y(ori00));
  INV        o154(.A(i_8_), .Y(ori_ori_n167_));
  INV        m000(.A(i_3_), .Y(mai_mai_n11_));
  INV        m001(.A(i_6_), .Y(mai_mai_n12_));
  NA2        m002(.A(i_4_), .B(mai_mai_n12_), .Y(mai_mai_n13_));
  INV        m003(.A(i_5_), .Y(mai_mai_n14_));
  NOi21      m004(.An(i_3_), .B(i_7_), .Y(mai_mai_n15_));
  NA3        m005(.A(mai_mai_n15_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n16_));
  INV        m006(.A(i_0_), .Y(mai_mai_n17_));
  NOi21      m007(.An(i_1_), .B(i_3_), .Y(mai_mai_n18_));
  NA3        m008(.A(mai_mai_n18_), .B(mai_mai_n17_), .C(i_2_), .Y(mai_mai_n19_));
  AOI210     m009(.A0(mai_mai_n19_), .A1(mai_mai_n16_), .B0(mai_mai_n13_), .Y(mai_mai_n20_));
  INV        m010(.A(i_4_), .Y(mai_mai_n21_));
  NA2        m011(.A(i_0_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  INV        m012(.A(i_7_), .Y(mai_mai_n23_));
  NA3        m013(.A(i_6_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n24_));
  NOi21      m014(.An(i_8_), .B(i_6_), .Y(mai_mai_n25_));
  NOi21      m015(.An(i_1_), .B(i_8_), .Y(mai_mai_n26_));
  AOI220     m016(.A0(mai_mai_n26_), .A1(i_2_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n27_));
  AOI210     m017(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n22_), .Y(mai_mai_n28_));
  AOI210     m018(.A0(mai_mai_n28_), .A1(mai_mai_n11_), .B0(mai_mai_n20_), .Y(mai_mai_n29_));
  NA2        m019(.A(i_0_), .B(mai_mai_n14_), .Y(mai_mai_n30_));
  NA2        m020(.A(mai_mai_n17_), .B(i_5_), .Y(mai_mai_n31_));
  NO2        m021(.A(i_2_), .B(i_4_), .Y(mai_mai_n32_));
  NA3        m022(.A(mai_mai_n32_), .B(i_6_), .C(i_8_), .Y(mai_mai_n33_));
  AOI210     m023(.A0(mai_mai_n31_), .A1(mai_mai_n30_), .B0(mai_mai_n33_), .Y(mai_mai_n34_));
  INV        m024(.A(i_2_), .Y(mai_mai_n35_));
  NOi21      m025(.An(i_5_), .B(i_0_), .Y(mai_mai_n36_));
  NOi21      m026(.An(i_6_), .B(i_8_), .Y(mai_mai_n37_));
  NOi21      m027(.An(i_7_), .B(i_1_), .Y(mai_mai_n38_));
  NOi21      m028(.An(i_5_), .B(i_6_), .Y(mai_mai_n39_));
  AOI220     m029(.A0(mai_mai_n39_), .A1(mai_mai_n38_), .B0(mai_mai_n37_), .B1(mai_mai_n36_), .Y(mai_mai_n40_));
  NO3        m030(.A(mai_mai_n40_), .B(mai_mai_n35_), .C(i_4_), .Y(mai_mai_n41_));
  NOi21      m031(.An(i_0_), .B(i_4_), .Y(mai_mai_n42_));
  NOi21      m032(.An(i_7_), .B(i_5_), .Y(mai_mai_n43_));
  AN2        m033(.A(mai_mai_n43_), .B(mai_mai_n42_), .Y(mai_mai_n44_));
  INV        m034(.A(i_1_), .Y(mai_mai_n45_));
  NOi21      m035(.An(i_3_), .B(i_0_), .Y(mai_mai_n46_));
  NA2        m036(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NA3        m037(.A(i_6_), .B(mai_mai_n14_), .C(i_7_), .Y(mai_mai_n48_));
  AOI210     m038(.A0(mai_mai_n48_), .A1(mai_mai_n24_), .B0(mai_mai_n47_), .Y(mai_mai_n49_));
  NO4        m039(.A(mai_mai_n49_), .B(mai_mai_n44_), .C(mai_mai_n41_), .D(mai_mai_n34_), .Y(mai_mai_n50_));
  INV        m040(.A(i_8_), .Y(mai_mai_n51_));
  NA2        m041(.A(i_1_), .B(mai_mai_n11_), .Y(mai_mai_n52_));
  NO4        m042(.A(mai_mai_n52_), .B(mai_mai_n30_), .C(i_2_), .D(mai_mai_n51_), .Y(mai_mai_n53_));
  NOi21      m043(.An(i_4_), .B(i_0_), .Y(mai_mai_n54_));
  AOI210     m044(.A0(mai_mai_n54_), .A1(mai_mai_n25_), .B0(mai_mai_n15_), .Y(mai_mai_n55_));
  NA2        m045(.A(i_1_), .B(mai_mai_n14_), .Y(mai_mai_n56_));
  NOi21      m046(.An(i_2_), .B(i_8_), .Y(mai_mai_n57_));
  NO2        m047(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n58_));
  NO2        m048(.A(mai_mai_n58_), .B(mai_mai_n53_), .Y(mai_mai_n59_));
  NOi31      m049(.An(i_2_), .B(i_1_), .C(i_3_), .Y(mai_mai_n60_));
  NOi21      m050(.An(i_4_), .B(i_3_), .Y(mai_mai_n61_));
  NOi21      m051(.An(i_1_), .B(i_4_), .Y(mai_mai_n62_));
  OAI210     m052(.A0(mai_mai_n62_), .A1(mai_mai_n61_), .B0(mai_mai_n57_), .Y(mai_mai_n63_));
  INV        m053(.A(mai_mai_n63_), .Y(mai_mai_n64_));
  AN2        m054(.A(i_8_), .B(i_7_), .Y(mai_mai_n65_));
  NA2        m055(.A(mai_mai_n65_), .B(mai_mai_n12_), .Y(mai_mai_n66_));
  NOi21      m056(.An(i_8_), .B(i_7_), .Y(mai_mai_n67_));
  NA3        m057(.A(mai_mai_n67_), .B(mai_mai_n61_), .C(i_6_), .Y(mai_mai_n68_));
  OAI210     m058(.A0(mai_mai_n66_), .A1(mai_mai_n56_), .B0(mai_mai_n68_), .Y(mai_mai_n69_));
  AOI220     m059(.A0(mai_mai_n69_), .A1(mai_mai_n35_), .B0(mai_mai_n64_), .B1(mai_mai_n39_), .Y(mai_mai_n70_));
  NA4        m060(.A(mai_mai_n70_), .B(mai_mai_n59_), .C(mai_mai_n50_), .D(mai_mai_n29_), .Y(mai_mai_n71_));
  NA2        m061(.A(i_8_), .B(i_7_), .Y(mai_mai_n72_));
  NO3        m062(.A(mai_mai_n72_), .B(mai_mai_n13_), .C(i_1_), .Y(mai_mai_n73_));
  NA2        m063(.A(i_8_), .B(mai_mai_n23_), .Y(mai_mai_n74_));
  NOi21      m064(.An(i_1_), .B(i_2_), .Y(mai_mai_n75_));
  NA3        m065(.A(mai_mai_n75_), .B(mai_mai_n54_), .C(i_6_), .Y(mai_mai_n76_));
  OAI210     m066(.A0(mai_mai_n174_), .A1(mai_mai_n74_), .B0(mai_mai_n76_), .Y(mai_mai_n77_));
  OAI210     m067(.A0(mai_mai_n77_), .A1(mai_mai_n73_), .B0(mai_mai_n14_), .Y(mai_mai_n78_));
  NA3        m068(.A(mai_mai_n67_), .B(i_2_), .C(mai_mai_n12_), .Y(mai_mai_n79_));
  NA3        m069(.A(mai_mai_n26_), .B(i_0_), .C(mai_mai_n14_), .Y(mai_mai_n80_));
  NA2        m070(.A(mai_mai_n80_), .B(mai_mai_n79_), .Y(mai_mai_n81_));
  NOi32      m071(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(mai_mai_n82_));
  NA2        m072(.A(mai_mai_n82_), .B(i_3_), .Y(mai_mai_n83_));
  NA3        m073(.A(mai_mai_n18_), .B(i_2_), .C(i_6_), .Y(mai_mai_n84_));
  NA2        m074(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  NO2        m075(.A(i_0_), .B(i_4_), .Y(mai_mai_n86_));
  AOI220     m076(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n81_), .B1(mai_mai_n61_), .Y(mai_mai_n87_));
  NA2        m077(.A(mai_mai_n87_), .B(mai_mai_n78_), .Y(mai_mai_n88_));
  NAi21      m078(.An(i_3_), .B(i_6_), .Y(mai_mai_n89_));
  NO3        m079(.A(mai_mai_n89_), .B(i_0_), .C(mai_mai_n51_), .Y(mai_mai_n90_));
  NA2        m080(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n91_));
  NOi21      m081(.An(i_7_), .B(i_8_), .Y(mai_mai_n92_));
  NOi31      m082(.An(i_6_), .B(i_5_), .C(i_7_), .Y(mai_mai_n93_));
  AOI210     m083(.A0(mai_mai_n92_), .A1(mai_mai_n12_), .B0(mai_mai_n93_), .Y(mai_mai_n94_));
  OAI210     m084(.A0(mai_mai_n94_), .A1(mai_mai_n11_), .B0(mai_mai_n91_), .Y(mai_mai_n95_));
  OAI210     m085(.A0(mai_mai_n95_), .A1(mai_mai_n90_), .B0(mai_mai_n75_), .Y(mai_mai_n96_));
  NA3        m086(.A(mai_mai_n25_), .B(i_2_), .C(mai_mai_n14_), .Y(mai_mai_n97_));
  AOI210     m087(.A0(mai_mai_n22_), .A1(mai_mai_n52_), .B0(mai_mai_n97_), .Y(mai_mai_n98_));
  AOI220     m088(.A0(mai_mai_n46_), .A1(mai_mai_n45_), .B0(mai_mai_n18_), .B1(mai_mai_n35_), .Y(mai_mai_n99_));
  NA3        m089(.A(mai_mai_n21_), .B(i_5_), .C(i_7_), .Y(mai_mai_n100_));
  NO2        m090(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NO2        m091(.A(mai_mai_n101_), .B(mai_mai_n98_), .Y(mai_mai_n102_));
  NA3        m092(.A(mai_mai_n67_), .B(mai_mai_n35_), .C(i_3_), .Y(mai_mai_n103_));
  NA2        m093(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n104_));
  AOI210     m094(.A0(mai_mai_n104_), .A1(mai_mai_n22_), .B0(mai_mai_n103_), .Y(mai_mai_n105_));
  NOi21      m095(.An(i_2_), .B(i_1_), .Y(mai_mai_n106_));
  NAi21      m096(.An(i_6_), .B(i_0_), .Y(mai_mai_n107_));
  NA3        m097(.A(mai_mai_n62_), .B(i_5_), .C(mai_mai_n23_), .Y(mai_mai_n108_));
  NOi21      m098(.An(i_4_), .B(i_6_), .Y(mai_mai_n109_));
  NOi21      m099(.An(i_5_), .B(i_3_), .Y(mai_mai_n110_));
  NA3        m100(.A(mai_mai_n110_), .B(mai_mai_n75_), .C(mai_mai_n109_), .Y(mai_mai_n111_));
  OAI210     m101(.A0(mai_mai_n108_), .A1(mai_mai_n107_), .B0(mai_mai_n111_), .Y(mai_mai_n112_));
  NA2        m102(.A(mai_mai_n75_), .B(mai_mai_n37_), .Y(mai_mai_n113_));
  NOi21      m103(.An(mai_mai_n43_), .B(mai_mai_n113_), .Y(mai_mai_n114_));
  NO3        m104(.A(mai_mai_n114_), .B(mai_mai_n112_), .C(mai_mai_n105_), .Y(mai_mai_n115_));
  NOi21      m105(.An(i_6_), .B(i_1_), .Y(mai_mai_n116_));
  AOI220     m106(.A0(mai_mai_n116_), .A1(i_7_), .B0(mai_mai_n25_), .B1(i_5_), .Y(mai_mai_n117_));
  NOi31      m107(.An(mai_mai_n54_), .B(mai_mai_n117_), .C(i_2_), .Y(mai_mai_n118_));
  NA2        m108(.A(mai_mai_n67_), .B(mai_mai_n12_), .Y(mai_mai_n119_));
  NA2        m109(.A(mai_mai_n37_), .B(mai_mai_n14_), .Y(mai_mai_n120_));
  NOi21      m110(.An(i_3_), .B(i_1_), .Y(mai_mai_n121_));
  NA2        m111(.A(mai_mai_n121_), .B(i_4_), .Y(mai_mai_n122_));
  AOI210     m112(.A0(mai_mai_n120_), .A1(mai_mai_n119_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  AOI220     m113(.A0(mai_mai_n92_), .A1(mai_mai_n14_), .B0(mai_mai_n109_), .B1(mai_mai_n23_), .Y(mai_mai_n124_));
  NOi31      m114(.An(mai_mai_n46_), .B(mai_mai_n124_), .C(mai_mai_n35_), .Y(mai_mai_n125_));
  NO3        m115(.A(mai_mai_n125_), .B(mai_mai_n123_), .C(mai_mai_n118_), .Y(mai_mai_n126_));
  NA4        m116(.A(mai_mai_n126_), .B(mai_mai_n115_), .C(mai_mai_n102_), .D(mai_mai_n96_), .Y(mai_mai_n127_));
  NA2        m117(.A(mai_mai_n57_), .B(mai_mai_n15_), .Y(mai_mai_n128_));
  NOi31      m118(.An(i_5_), .B(i_2_), .C(i_6_), .Y(mai_mai_n129_));
  NA2        m119(.A(mai_mai_n129_), .B(i_7_), .Y(mai_mai_n130_));
  NA3        m120(.A(mai_mai_n130_), .B(mai_mai_n128_), .C(mai_mai_n113_), .Y(mai_mai_n131_));
  NA2        m121(.A(mai_mai_n131_), .B(mai_mai_n42_), .Y(mai_mai_n132_));
  NO2        m122(.A(mai_mai_n79_), .B(mai_mai_n31_), .Y(mai_mai_n133_));
  NA4        m123(.A(mai_mai_n65_), .B(mai_mai_n106_), .C(mai_mai_n17_), .D(mai_mai_n12_), .Y(mai_mai_n134_));
  NAi31      m124(.An(mai_mai_n107_), .B(mai_mai_n92_), .C(mai_mai_n106_), .Y(mai_mai_n135_));
  NA3        m125(.A(mai_mai_n67_), .B(mai_mai_n60_), .C(i_6_), .Y(mai_mai_n136_));
  NA3        m126(.A(mai_mai_n136_), .B(mai_mai_n135_), .C(mai_mai_n134_), .Y(mai_mai_n137_));
  NOi21      m127(.An(i_0_), .B(i_2_), .Y(mai_mai_n138_));
  NA3        m128(.A(mai_mai_n138_), .B(mai_mai_n38_), .C(mai_mai_n109_), .Y(mai_mai_n139_));
  NA3        m129(.A(mai_mai_n54_), .B(mai_mai_n43_), .C(mai_mai_n18_), .Y(mai_mai_n140_));
  NA3        m130(.A(mai_mai_n138_), .B(mai_mai_n61_), .C(mai_mai_n37_), .Y(mai_mai_n141_));
  NA3        m131(.A(mai_mai_n141_), .B(mai_mai_n140_), .C(mai_mai_n139_), .Y(mai_mai_n142_));
  NA4        m132(.A(mai_mai_n60_), .B(i_6_), .C(mai_mai_n14_), .D(i_7_), .Y(mai_mai_n143_));
  NA4        m133(.A(mai_mai_n62_), .B(mai_mai_n39_), .C(mai_mai_n17_), .D(i_8_), .Y(mai_mai_n144_));
  NA4        m134(.A(mai_mai_n62_), .B(mai_mai_n46_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n145_));
  NA3        m135(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(mai_mai_n143_), .Y(mai_mai_n146_));
  NO4        m136(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n137_), .D(mai_mai_n133_), .Y(mai_mai_n147_));
  AOI220     m137(.A0(i_5_), .A1(mai_mai_n92_), .B0(mai_mai_n65_), .B1(mai_mai_n32_), .Y(mai_mai_n148_));
  AOI210     m138(.A0(mai_mai_n148_), .A1(mai_mai_n128_), .B0(mai_mai_n104_), .Y(mai_mai_n149_));
  NO4        m139(.A(i_2_), .B(mai_mai_n21_), .C(mai_mai_n11_), .D(mai_mai_n14_), .Y(mai_mai_n150_));
  NA2        m140(.A(i_2_), .B(i_4_), .Y(mai_mai_n151_));
  AOI210     m141(.A0(mai_mai_n107_), .A1(mai_mai_n89_), .B0(mai_mai_n151_), .Y(mai_mai_n152_));
  NO2        m142(.A(i_8_), .B(i_7_), .Y(mai_mai_n153_));
  OA210      m143(.A0(mai_mai_n152_), .A1(mai_mai_n150_), .B0(mai_mai_n153_), .Y(mai_mai_n154_));
  NA4        m144(.A(mai_mai_n121_), .B(i_0_), .C(i_5_), .D(mai_mai_n23_), .Y(mai_mai_n155_));
  NO2        m145(.A(mai_mai_n155_), .B(i_4_), .Y(mai_mai_n156_));
  NO3        m146(.A(mai_mai_n156_), .B(mai_mai_n154_), .C(mai_mai_n149_), .Y(mai_mai_n157_));
  NA2        m147(.A(mai_mai_n92_), .B(mai_mai_n12_), .Y(mai_mai_n158_));
  NA3        m148(.A(i_2_), .B(i_1_), .C(mai_mai_n14_), .Y(mai_mai_n159_));
  NA2        m149(.A(mai_mai_n54_), .B(i_3_), .Y(mai_mai_n160_));
  AOI210     m150(.A0(mai_mai_n160_), .A1(mai_mai_n159_), .B0(mai_mai_n158_), .Y(mai_mai_n161_));
  NA3        m151(.A(mai_mai_n138_), .B(mai_mai_n67_), .C(mai_mai_n109_), .Y(mai_mai_n162_));
  OAI210     m152(.A0(mai_mai_n103_), .A1(mai_mai_n31_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  NA3        m153(.A(mai_mai_n110_), .B(mai_mai_n65_), .C(mai_mai_n45_), .Y(mai_mai_n164_));
  NA3        m154(.A(mai_mai_n57_), .B(mai_mai_n36_), .C(mai_mai_n15_), .Y(mai_mai_n165_));
  NOi31      m155(.An(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n166_));
  NA2        m156(.A(mai_mai_n82_), .B(mai_mai_n166_), .Y(mai_mai_n167_));
  NA3        m157(.A(mai_mai_n167_), .B(mai_mai_n165_), .C(mai_mai_n164_), .Y(mai_mai_n168_));
  NO3        m158(.A(mai_mai_n168_), .B(mai_mai_n163_), .C(mai_mai_n161_), .Y(mai_mai_n169_));
  NA4        m159(.A(mai_mai_n169_), .B(mai_mai_n157_), .C(mai_mai_n147_), .D(mai_mai_n132_), .Y(mai_mai_n170_));
  OR4        m160(.A(mai_mai_n170_), .B(mai_mai_n127_), .C(mai_mai_n88_), .D(mai_mai_n71_), .Y(mai00));
  INV        m161(.A(i_2_), .Y(mai_mai_n174_));
  INV        u000(.A(i_3_), .Y(men_men_n11_));
  INV        u001(.A(i_6_), .Y(men_men_n12_));
  NA2        u002(.A(i_4_), .B(men_men_n12_), .Y(men_men_n13_));
  INV        u003(.A(i_5_), .Y(men_men_n14_));
  NOi21      u004(.An(i_3_), .B(i_7_), .Y(men_men_n15_));
  NA3        u005(.A(men_men_n15_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n16_));
  INV        u006(.A(i_0_), .Y(men_men_n17_));
  NOi21      u007(.An(i_1_), .B(i_3_), .Y(men_men_n18_));
  NA3        u008(.A(men_men_n18_), .B(men_men_n17_), .C(i_2_), .Y(men_men_n19_));
  AOI210     u009(.A0(men_men_n19_), .A1(men_men_n16_), .B0(men_men_n13_), .Y(men_men_n20_));
  INV        u010(.A(i_4_), .Y(men_men_n21_));
  NA2        u011(.A(i_0_), .B(men_men_n21_), .Y(men_men_n22_));
  INV        u012(.A(i_7_), .Y(men_men_n23_));
  NOi21      u013(.An(i_8_), .B(i_6_), .Y(men_men_n24_));
  AOI210     u014(.A0(men_men_n172_), .A1(men_men_n173_), .B0(men_men_n22_), .Y(men_men_n25_));
  AOI210     u015(.A0(men_men_n25_), .A1(men_men_n11_), .B0(men_men_n20_), .Y(men_men_n26_));
  NA2        u016(.A(i_0_), .B(men_men_n14_), .Y(men_men_n27_));
  NA2        u017(.A(men_men_n17_), .B(i_5_), .Y(men_men_n28_));
  NO2        u018(.A(i_2_), .B(i_4_), .Y(men_men_n29_));
  NA3        u019(.A(men_men_n29_), .B(i_6_), .C(i_8_), .Y(men_men_n30_));
  AOI210     u020(.A0(men_men_n28_), .A1(men_men_n27_), .B0(men_men_n30_), .Y(men_men_n31_));
  INV        u021(.A(i_2_), .Y(men_men_n32_));
  NOi21      u022(.An(i_5_), .B(i_0_), .Y(men_men_n33_));
  NOi21      u023(.An(i_6_), .B(i_8_), .Y(men_men_n34_));
  NOi21      u024(.An(i_7_), .B(i_1_), .Y(men_men_n35_));
  NOi21      u025(.An(i_5_), .B(i_6_), .Y(men_men_n36_));
  AOI220     u026(.A0(men_men_n36_), .A1(men_men_n35_), .B0(men_men_n34_), .B1(men_men_n33_), .Y(men_men_n37_));
  NO3        u027(.A(men_men_n37_), .B(men_men_n32_), .C(i_4_), .Y(men_men_n38_));
  NOi21      u028(.An(i_0_), .B(i_4_), .Y(men_men_n39_));
  XO2        u029(.A(i_1_), .B(i_3_), .Y(men_men_n40_));
  NOi21      u030(.An(i_7_), .B(i_5_), .Y(men_men_n41_));
  AN3        u031(.A(men_men_n41_), .B(men_men_n40_), .C(men_men_n39_), .Y(men_men_n42_));
  INV        u032(.A(i_1_), .Y(men_men_n43_));
  NOi21      u033(.An(i_3_), .B(i_0_), .Y(men_men_n44_));
  NO3        u034(.A(men_men_n42_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n45_));
  INV        u035(.A(i_8_), .Y(men_men_n46_));
  NOi21      u036(.An(i_4_), .B(i_0_), .Y(men_men_n47_));
  AOI210     u037(.A0(men_men_n47_), .A1(men_men_n24_), .B0(men_men_n15_), .Y(men_men_n48_));
  NA2        u038(.A(i_1_), .B(men_men_n14_), .Y(men_men_n49_));
  NOi21      u039(.An(i_2_), .B(i_8_), .Y(men_men_n50_));
  NO3        u040(.A(men_men_n50_), .B(men_men_n47_), .C(men_men_n39_), .Y(men_men_n51_));
  NO3        u041(.A(men_men_n51_), .B(men_men_n49_), .C(men_men_n48_), .Y(men_men_n52_));
  INV        u042(.A(men_men_n52_), .Y(men_men_n53_));
  NOi31      u043(.An(i_2_), .B(i_1_), .C(i_3_), .Y(men_men_n54_));
  NA2        u044(.A(men_men_n54_), .B(i_0_), .Y(men_men_n55_));
  NOi21      u045(.An(i_4_), .B(i_3_), .Y(men_men_n56_));
  NOi21      u046(.An(i_1_), .B(i_4_), .Y(men_men_n57_));
  OAI210     u047(.A0(men_men_n57_), .A1(men_men_n56_), .B0(men_men_n50_), .Y(men_men_n58_));
  NA2        u048(.A(men_men_n58_), .B(men_men_n55_), .Y(men_men_n59_));
  AN2        u049(.A(i_8_), .B(i_7_), .Y(men_men_n60_));
  NA2        u050(.A(men_men_n60_), .B(men_men_n12_), .Y(men_men_n61_));
  NOi21      u051(.An(i_8_), .B(i_7_), .Y(men_men_n62_));
  NA3        u052(.A(men_men_n62_), .B(men_men_n56_), .C(i_6_), .Y(men_men_n63_));
  OAI210     u053(.A0(men_men_n61_), .A1(men_men_n49_), .B0(men_men_n63_), .Y(men_men_n64_));
  AOI220     u054(.A0(men_men_n64_), .A1(men_men_n32_), .B0(men_men_n59_), .B1(men_men_n36_), .Y(men_men_n65_));
  NA4        u055(.A(men_men_n65_), .B(men_men_n53_), .C(men_men_n45_), .D(men_men_n26_), .Y(men_men_n66_));
  NA2        u056(.A(i_8_), .B(i_7_), .Y(men_men_n67_));
  NO3        u057(.A(men_men_n67_), .B(men_men_n13_), .C(i_1_), .Y(men_men_n68_));
  NA2        u058(.A(i_8_), .B(men_men_n23_), .Y(men_men_n69_));
  AOI220     u059(.A0(men_men_n44_), .A1(i_1_), .B0(men_men_n40_), .B1(i_2_), .Y(men_men_n70_));
  NOi21      u060(.An(i_1_), .B(i_2_), .Y(men_men_n71_));
  NA3        u061(.A(men_men_n71_), .B(men_men_n47_), .C(i_6_), .Y(men_men_n72_));
  OAI210     u062(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n72_), .Y(men_men_n73_));
  OAI210     u063(.A0(men_men_n73_), .A1(men_men_n68_), .B0(men_men_n14_), .Y(men_men_n74_));
  NA3        u064(.A(men_men_n62_), .B(i_2_), .C(men_men_n12_), .Y(men_men_n75_));
  NA3        u065(.A(i_1_), .B(i_0_), .C(men_men_n14_), .Y(men_men_n76_));
  NA2        u066(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  NOi32      u067(.An(i_8_), .Bn(i_7_), .C(i_5_), .Y(men_men_n78_));
  NA2        u068(.A(men_men_n78_), .B(i_3_), .Y(men_men_n79_));
  NA3        u069(.A(men_men_n18_), .B(i_2_), .C(i_6_), .Y(men_men_n80_));
  NA2        u070(.A(men_men_n80_), .B(men_men_n79_), .Y(men_men_n81_));
  NO2        u071(.A(i_0_), .B(i_4_), .Y(men_men_n82_));
  AOI220     u072(.A0(men_men_n82_), .A1(men_men_n81_), .B0(men_men_n77_), .B1(men_men_n56_), .Y(men_men_n83_));
  NA2        u073(.A(men_men_n83_), .B(men_men_n74_), .Y(men_men_n84_));
  NAi21      u074(.An(i_3_), .B(i_6_), .Y(men_men_n85_));
  NO3        u075(.A(men_men_n85_), .B(i_0_), .C(men_men_n46_), .Y(men_men_n86_));
  NA2        u076(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n87_));
  NOi21      u077(.An(i_7_), .B(i_8_), .Y(men_men_n88_));
  NOi31      u078(.An(i_6_), .B(i_5_), .C(i_7_), .Y(men_men_n89_));
  AOI210     u079(.A0(men_men_n88_), .A1(men_men_n12_), .B0(men_men_n89_), .Y(men_men_n90_));
  OAI210     u080(.A0(men_men_n90_), .A1(men_men_n11_), .B0(men_men_n87_), .Y(men_men_n91_));
  OAI210     u081(.A0(men_men_n91_), .A1(men_men_n86_), .B0(men_men_n71_), .Y(men_men_n92_));
  NA3        u082(.A(men_men_n24_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n93_));
  NO2        u083(.A(men_men_n22_), .B(men_men_n93_), .Y(men_men_n94_));
  NA2        u084(.A(men_men_n44_), .B(men_men_n43_), .Y(men_men_n95_));
  OAI210     u085(.A0(i_4_), .A1(i_7_), .B0(i_5_), .Y(men_men_n96_));
  NA3        u086(.A(men_men_n67_), .B(men_men_n18_), .C(men_men_n17_), .Y(men_men_n97_));
  OAI220     u087(.A0(men_men_n97_), .A1(men_men_n96_), .B0(men_men_n174_), .B1(men_men_n95_), .Y(men_men_n98_));
  NO2        u088(.A(men_men_n98_), .B(men_men_n94_), .Y(men_men_n99_));
  NA3        u089(.A(men_men_n62_), .B(men_men_n32_), .C(i_3_), .Y(men_men_n100_));
  NA2        u090(.A(men_men_n43_), .B(i_6_), .Y(men_men_n101_));
  AOI210     u091(.A0(men_men_n101_), .A1(men_men_n22_), .B0(men_men_n100_), .Y(men_men_n102_));
  NOi21      u092(.An(i_2_), .B(i_1_), .Y(men_men_n103_));
  AN3        u093(.A(men_men_n88_), .B(men_men_n103_), .C(men_men_n47_), .Y(men_men_n104_));
  NAi21      u094(.An(i_6_), .B(i_0_), .Y(men_men_n105_));
  NOi21      u095(.An(i_4_), .B(i_6_), .Y(men_men_n106_));
  NOi21      u096(.An(i_5_), .B(i_3_), .Y(men_men_n107_));
  NA3        u097(.A(men_men_n107_), .B(men_men_n71_), .C(men_men_n106_), .Y(men_men_n108_));
  INV        u098(.A(men_men_n108_), .Y(men_men_n109_));
  NA2        u099(.A(men_men_n71_), .B(men_men_n34_), .Y(men_men_n110_));
  NOi21      u100(.An(men_men_n41_), .B(men_men_n110_), .Y(men_men_n111_));
  NO4        u101(.A(men_men_n111_), .B(men_men_n109_), .C(men_men_n104_), .D(men_men_n102_), .Y(men_men_n112_));
  NOi21      u102(.An(i_6_), .B(i_1_), .Y(men_men_n113_));
  AOI220     u103(.A0(men_men_n113_), .A1(i_7_), .B0(men_men_n24_), .B1(i_5_), .Y(men_men_n114_));
  NOi31      u104(.An(men_men_n47_), .B(men_men_n114_), .C(i_2_), .Y(men_men_n115_));
  NA2        u105(.A(men_men_n62_), .B(men_men_n12_), .Y(men_men_n116_));
  NA2        u106(.A(men_men_n34_), .B(men_men_n14_), .Y(men_men_n117_));
  NOi21      u107(.An(i_3_), .B(i_1_), .Y(men_men_n118_));
  NA2        u108(.A(men_men_n118_), .B(i_4_), .Y(men_men_n119_));
  AOI210     u109(.A0(men_men_n117_), .A1(men_men_n116_), .B0(men_men_n119_), .Y(men_men_n120_));
  AOI220     u110(.A0(men_men_n88_), .A1(men_men_n14_), .B0(men_men_n106_), .B1(men_men_n23_), .Y(men_men_n121_));
  NOi31      u111(.An(men_men_n44_), .B(men_men_n121_), .C(men_men_n32_), .Y(men_men_n122_));
  NO3        u112(.A(men_men_n122_), .B(men_men_n120_), .C(men_men_n115_), .Y(men_men_n123_));
  NA4        u113(.A(men_men_n123_), .B(men_men_n112_), .C(men_men_n99_), .D(men_men_n92_), .Y(men_men_n124_));
  NA2        u114(.A(men_men_n50_), .B(men_men_n15_), .Y(men_men_n125_));
  NOi31      u115(.An(i_6_), .B(i_1_), .C(i_8_), .Y(men_men_n126_));
  NOi31      u116(.An(i_5_), .B(i_2_), .C(i_6_), .Y(men_men_n127_));
  OAI210     u117(.A0(men_men_n127_), .A1(men_men_n126_), .B0(i_7_), .Y(men_men_n128_));
  NA3        u118(.A(men_men_n34_), .B(i_2_), .C(men_men_n14_), .Y(men_men_n129_));
  NA4        u119(.A(men_men_n129_), .B(men_men_n128_), .C(men_men_n125_), .D(men_men_n110_), .Y(men_men_n130_));
  NA2        u120(.A(men_men_n130_), .B(men_men_n39_), .Y(men_men_n131_));
  NA2        u121(.A(men_men_n56_), .B(men_men_n35_), .Y(men_men_n132_));
  AOI210     u122(.A0(men_men_n132_), .A1(men_men_n75_), .B0(men_men_n28_), .Y(men_men_n133_));
  NAi31      u123(.An(men_men_n105_), .B(men_men_n88_), .C(men_men_n103_), .Y(men_men_n134_));
  NA3        u124(.A(men_men_n62_), .B(men_men_n54_), .C(i_6_), .Y(men_men_n135_));
  NA2        u125(.A(men_men_n135_), .B(men_men_n134_), .Y(men_men_n136_));
  NOi21      u126(.An(i_0_), .B(i_2_), .Y(men_men_n137_));
  NA3        u127(.A(men_men_n137_), .B(men_men_n35_), .C(men_men_n106_), .Y(men_men_n138_));
  NA3        u128(.A(men_men_n47_), .B(men_men_n41_), .C(men_men_n18_), .Y(men_men_n139_));
  NOi32      u129(.An(i_4_), .Bn(i_5_), .C(i_3_), .Y(men_men_n140_));
  NA2        u130(.A(men_men_n140_), .B(men_men_n126_), .Y(men_men_n141_));
  NA3        u131(.A(men_men_n137_), .B(men_men_n56_), .C(men_men_n34_), .Y(men_men_n142_));
  NA4        u132(.A(men_men_n142_), .B(men_men_n141_), .C(men_men_n139_), .D(men_men_n138_), .Y(men_men_n143_));
  NA4        u133(.A(men_men_n54_), .B(i_6_), .C(men_men_n14_), .D(i_7_), .Y(men_men_n144_));
  NA4        u134(.A(men_men_n57_), .B(men_men_n36_), .C(men_men_n17_), .D(i_8_), .Y(men_men_n145_));
  NA2        u135(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n146_));
  NO4        u136(.A(men_men_n146_), .B(men_men_n143_), .C(men_men_n136_), .D(men_men_n133_), .Y(men_men_n147_));
  NA2        u137(.A(men_men_n60_), .B(men_men_n29_), .Y(men_men_n148_));
  AOI210     u138(.A0(men_men_n148_), .A1(men_men_n125_), .B0(men_men_n101_), .Y(men_men_n149_));
  NO3        u139(.A(i_2_), .B(men_men_n11_), .C(men_men_n14_), .Y(men_men_n150_));
  NA2        u140(.A(i_2_), .B(i_4_), .Y(men_men_n151_));
  AOI210     u141(.A0(men_men_n105_), .A1(men_men_n85_), .B0(men_men_n151_), .Y(men_men_n152_));
  NO2        u142(.A(i_8_), .B(i_7_), .Y(men_men_n153_));
  OA210      u143(.A0(men_men_n152_), .A1(men_men_n150_), .B0(men_men_n153_), .Y(men_men_n154_));
  NO2        u144(.A(men_men_n154_), .B(men_men_n149_), .Y(men_men_n155_));
  NA2        u145(.A(men_men_n88_), .B(men_men_n12_), .Y(men_men_n156_));
  NA3        u146(.A(i_2_), .B(i_1_), .C(men_men_n14_), .Y(men_men_n157_));
  NO2        u147(.A(men_men_n157_), .B(men_men_n156_), .Y(men_men_n158_));
  NA3        u148(.A(men_men_n137_), .B(men_men_n62_), .C(men_men_n106_), .Y(men_men_n159_));
  INV        u149(.A(men_men_n159_), .Y(men_men_n160_));
  NA4        u150(.A(men_men_n107_), .B(men_men_n60_), .C(men_men_n43_), .D(men_men_n21_), .Y(men_men_n161_));
  NA3        u151(.A(men_men_n89_), .B(men_men_n118_), .C(i_0_), .Y(men_men_n162_));
  NA2        u152(.A(men_men_n33_), .B(men_men_n15_), .Y(men_men_n163_));
  NOi31      u153(.An(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n164_));
  OAI210     u154(.A0(men_men_n140_), .A1(men_men_n78_), .B0(men_men_n164_), .Y(men_men_n165_));
  NA4        u155(.A(men_men_n165_), .B(men_men_n163_), .C(men_men_n162_), .D(men_men_n161_), .Y(men_men_n166_));
  NO3        u156(.A(men_men_n166_), .B(men_men_n160_), .C(men_men_n158_), .Y(men_men_n167_));
  NA4        u157(.A(men_men_n167_), .B(men_men_n155_), .C(men_men_n147_), .D(men_men_n131_), .Y(men_men_n168_));
  OR4        u158(.A(men_men_n168_), .B(men_men_n124_), .C(men_men_n84_), .D(men_men_n66_), .Y(men00));
  INV        u159(.A(i_1_), .Y(men_men_n172_));
  INV        u160(.A(i_5_), .Y(men_men_n173_));
  INV        u161(.A(i_7_), .Y(men_men_n174_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
endmodule