//Benchmark atmr_alu4_1266_0.0625

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n133_, ori_ori_n134_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n987_, mai_mai_n988_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NA2        o032(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n55_));
  NO2        o033(.A(i_1_), .B(i_6_), .Y(ori_ori_n56_));
  NA2        o034(.A(i_8_), .B(i_7_), .Y(ori_ori_n57_));
  NAi21      o035(.An(i_2_), .B(i_7_), .Y(ori_ori_n58_));
  INV        o036(.A(i_1_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(i_6_), .Y(ori_ori_n60_));
  NA3        o038(.A(ori_ori_n60_), .B(ori_ori_n58_), .C(ori_ori_n31_), .Y(ori_ori_n61_));
  NA2        o039(.A(i_1_), .B(i_10_), .Y(ori_ori_n62_));
  NO2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NAi21      o041(.An(ori_ori_n63_), .B(ori_ori_n61_), .Y(ori_ori_n64_));
  NA2        o042(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n65_));
  AOI210     o043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n66_));
  NA2        o044(.A(i_1_), .B(i_6_), .Y(ori_ori_n67_));
  NO2        o045(.A(ori_ori_n67_), .B(ori_ori_n25_), .Y(ori_ori_n68_));
  INV        o046(.A(i_0_), .Y(ori_ori_n69_));
  NAi21      o047(.An(i_5_), .B(i_10_), .Y(ori_ori_n70_));
  NA2        o048(.A(i_5_), .B(i_9_), .Y(ori_ori_n71_));
  AOI210     o049(.A0(ori_ori_n71_), .A1(ori_ori_n70_), .B0(ori_ori_n69_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n72_), .B(ori_ori_n68_), .Y(ori_ori_n73_));
  OAI210     o051(.A0(ori_ori_n66_), .A1(ori_ori_n65_), .B0(ori_ori_n73_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n64_), .B0(i_0_), .Y(ori_ori_n75_));
  NA2        o053(.A(i_12_), .B(i_5_), .Y(ori_ori_n76_));
  NA2        o054(.A(i_2_), .B(i_8_), .Y(ori_ori_n77_));
  NO2        o055(.A(ori_ori_n77_), .B(ori_ori_n56_), .Y(ori_ori_n78_));
  NO2        o056(.A(i_3_), .B(i_7_), .Y(ori_ori_n79_));
  INV        o057(.A(i_6_), .Y(ori_ori_n80_));
  OR4        o058(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(ori_ori_n81_));
  INV        o059(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_2_), .B(i_7_), .Y(ori_ori_n83_));
  INV        o061(.A(ori_ori_n78_), .Y(ori_ori_n84_));
  NAi21      o062(.An(i_6_), .B(i_10_), .Y(ori_ori_n85_));
  NA2        o063(.A(i_6_), .B(i_9_), .Y(ori_ori_n86_));
  AOI210     o064(.A0(ori_ori_n86_), .A1(ori_ori_n85_), .B0(ori_ori_n59_), .Y(ori_ori_n87_));
  NA2        o065(.A(i_2_), .B(i_6_), .Y(ori_ori_n88_));
  NO2        o066(.A(ori_ori_n88_), .B(ori_ori_n25_), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n89_), .B(ori_ori_n87_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n84_), .B0(ori_ori_n76_), .Y(ori_ori_n91_));
  AN3        o069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n92_));
  NAi21      o070(.An(i_6_), .B(i_11_), .Y(ori_ori_n93_));
  NA2        o071(.A(ori_ori_n92_), .B(ori_ori_n32_), .Y(ori_ori_n94_));
  INV        o072(.A(i_7_), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n46_), .B(ori_ori_n95_), .Y(ori_ori_n96_));
  NO2        o074(.A(i_0_), .B(i_5_), .Y(ori_ori_n97_));
  NO2        o075(.A(ori_ori_n97_), .B(ori_ori_n80_), .Y(ori_ori_n98_));
  NA2        o076(.A(i_12_), .B(i_3_), .Y(ori_ori_n99_));
  INV        o077(.A(ori_ori_n99_), .Y(ori_ori_n100_));
  NA3        o078(.A(ori_ori_n100_), .B(ori_ori_n98_), .C(ori_ori_n96_), .Y(ori_ori_n101_));
  NAi21      o079(.An(i_7_), .B(i_11_), .Y(ori_ori_n102_));
  NO3        o080(.A(ori_ori_n102_), .B(ori_ori_n85_), .C(ori_ori_n53_), .Y(ori_ori_n103_));
  AN2        o081(.A(i_2_), .B(i_10_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n104_), .B(i_7_), .Y(ori_ori_n105_));
  OR2        o083(.A(ori_ori_n76_), .B(ori_ori_n56_), .Y(ori_ori_n106_));
  NO2        o084(.A(i_8_), .B(ori_ori_n95_), .Y(ori_ori_n107_));
  NO3        o085(.A(ori_ori_n107_), .B(ori_ori_n106_), .C(ori_ori_n105_), .Y(ori_ori_n108_));
  NA2        o086(.A(i_12_), .B(i_7_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n59_), .B(ori_ori_n26_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n110_), .B(i_0_), .Y(ori_ori_n111_));
  NA2        o089(.A(i_11_), .B(i_12_), .Y(ori_ori_n112_));
  OAI210     o090(.A0(ori_ori_n111_), .A1(ori_ori_n109_), .B0(ori_ori_n112_), .Y(ori_ori_n113_));
  NO2        o091(.A(ori_ori_n113_), .B(ori_ori_n108_), .Y(ori_ori_n114_));
  NAi41      o092(.An(ori_ori_n103_), .B(ori_ori_n114_), .C(ori_ori_n101_), .D(ori_ori_n94_), .Y(ori_ori_n115_));
  NOi21      o093(.An(i_1_), .B(i_5_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n116_), .B(i_11_), .Y(ori_ori_n117_));
  NA2        o095(.A(ori_ori_n95_), .B(ori_ori_n37_), .Y(ori_ori_n118_));
  NA2        o096(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n119_));
  NA2        o097(.A(ori_ori_n119_), .B(ori_ori_n118_), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n120_), .B(ori_ori_n46_), .Y(ori_ori_n121_));
  NA2        o099(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n122_));
  NAi21      o100(.An(i_3_), .B(i_8_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n123_), .B(ori_ori_n58_), .Y(ori_ori_n124_));
  NOi31      o102(.An(ori_ori_n124_), .B(ori_ori_n122_), .C(ori_ori_n121_), .Y(ori_ori_n125_));
  NO2        o103(.A(i_1_), .B(ori_ori_n80_), .Y(ori_ori_n126_));
  NO2        o104(.A(i_6_), .B(i_5_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(i_3_), .Y(ori_ori_n128_));
  AO210      o106(.A0(ori_ori_n128_), .A1(ori_ori_n47_), .B0(ori_ori_n126_), .Y(ori_ori_n129_));
  OAI220     o107(.A0(ori_ori_n129_), .A1(ori_ori_n102_), .B0(ori_ori_n125_), .B1(ori_ori_n117_), .Y(ori_ori_n130_));
  NO3        o108(.A(ori_ori_n130_), .B(ori_ori_n115_), .C(ori_ori_n91_), .Y(ori_ori_n131_));
  NA3        o109(.A(ori_ori_n131_), .B(ori_ori_n75_), .C(ori_ori_n55_), .Y(ori2));
  NO2        o110(.A(ori_ori_n59_), .B(ori_ori_n37_), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n828_), .B(ori_ori_n133_), .Y(ori_ori_n134_));
  NA4        o112(.A(ori_ori_n134_), .B(ori_ori_n73_), .C(ori_ori_n65_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o113(.A(i_8_), .B(i_7_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(i_6_), .Y(ori_ori_n137_));
  NO2        o115(.A(i_12_), .B(i_13_), .Y(ori_ori_n138_));
  NAi21      o116(.An(i_5_), .B(i_11_), .Y(ori_ori_n139_));
  NOi21      o117(.An(ori_ori_n138_), .B(ori_ori_n139_), .Y(ori_ori_n140_));
  NO2        o118(.A(i_0_), .B(i_1_), .Y(ori_ori_n141_));
  NA2        o119(.A(i_2_), .B(i_3_), .Y(ori_ori_n142_));
  NO2        o120(.A(ori_ori_n142_), .B(i_4_), .Y(ori_ori_n143_));
  NA3        o121(.A(ori_ori_n143_), .B(ori_ori_n141_), .C(ori_ori_n140_), .Y(ori_ori_n144_));
  NA2        o122(.A(i_1_), .B(i_5_), .Y(ori_ori_n145_));
  OR2        o123(.A(i_0_), .B(i_1_), .Y(ori_ori_n146_));
  NAi32      o124(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n147_));
  NOi21      o125(.An(i_4_), .B(i_10_), .Y(ori_ori_n148_));
  NA2        o126(.A(ori_ori_n148_), .B(ori_ori_n40_), .Y(ori_ori_n149_));
  NO3        o127(.A(ori_ori_n69_), .B(i_2_), .C(i_1_), .Y(ori_ori_n150_));
  INV        o128(.A(ori_ori_n150_), .Y(ori_ori_n151_));
  NOi21      o129(.An(i_4_), .B(i_9_), .Y(ori_ori_n152_));
  NOi21      o130(.An(i_11_), .B(i_13_), .Y(ori_ori_n153_));
  NA2        o131(.A(ori_ori_n153_), .B(ori_ori_n152_), .Y(ori_ori_n154_));
  NO2        o132(.A(i_4_), .B(i_5_), .Y(ori_ori_n155_));
  NAi21      o133(.An(i_12_), .B(i_11_), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n156_), .B(i_13_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n69_), .B(ori_ori_n59_), .Y(ori_ori_n158_));
  NA2        o136(.A(i_3_), .B(i_5_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n69_), .B(i_5_), .Y(ori_ori_n160_));
  NO2        o138(.A(i_13_), .B(i_10_), .Y(ori_ori_n161_));
  NA3        o139(.A(ori_ori_n161_), .B(ori_ori_n160_), .C(ori_ori_n44_), .Y(ori_ori_n162_));
  NO2        o140(.A(i_2_), .B(i_1_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n163_), .B(i_3_), .Y(ori_ori_n164_));
  NAi21      o142(.An(i_4_), .B(i_12_), .Y(ori_ori_n165_));
  INV        o143(.A(i_8_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n166_), .B(i_7_), .Y(ori_ori_n167_));
  NO3        o145(.A(i_3_), .B(ori_ori_n80_), .C(ori_ori_n48_), .Y(ori_ori_n168_));
  NA2        o146(.A(ori_ori_n168_), .B(ori_ori_n107_), .Y(ori_ori_n169_));
  NO3        o147(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n170_));
  NO3        o148(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n171_));
  NO2        o149(.A(i_3_), .B(i_8_), .Y(ori_ori_n172_));
  NO3        o150(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n173_));
  NA3        o151(.A(ori_ori_n173_), .B(ori_ori_n172_), .C(ori_ori_n40_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n97_), .B(ori_ori_n56_), .Y(ori_ori_n175_));
  INV        o153(.A(ori_ori_n175_), .Y(ori_ori_n176_));
  NO2        o154(.A(i_13_), .B(i_9_), .Y(ori_ori_n177_));
  NAi21      o155(.An(i_12_), .B(i_3_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n176_), .B(ori_ori_n174_), .Y(ori_ori_n180_));
  NA2        o158(.A(ori_ori_n180_), .B(i_7_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n181_), .B(i_4_), .Y(ori_ori_n182_));
  NAi21      o160(.An(i_12_), .B(i_7_), .Y(ori_ori_n183_));
  NA3        o161(.A(i_13_), .B(ori_ori_n166_), .C(i_10_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n184_), .B(ori_ori_n183_), .Y(ori_ori_n185_));
  NA2        o163(.A(i_0_), .B(i_5_), .Y(ori_ori_n186_));
  OAI220     o164(.A0(ori_ori_n80_), .A1(ori_ori_n164_), .B0(i_2_), .B1(ori_ori_n128_), .Y(ori_ori_n187_));
  NAi31      o165(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n46_), .B(ori_ori_n59_), .Y(ori_ori_n190_));
  NA3        o168(.A(ori_ori_n190_), .B(i_3_), .C(ori_ori_n189_), .Y(ori_ori_n191_));
  INV        o169(.A(i_13_), .Y(ori_ori_n192_));
  NO2        o170(.A(i_12_), .B(ori_ori_n192_), .Y(ori_ori_n193_));
  NA3        o171(.A(ori_ori_n193_), .B(ori_ori_n170_), .C(ori_ori_n168_), .Y(ori_ori_n194_));
  OAI210     o172(.A0(ori_ori_n191_), .A1(ori_ori_n188_), .B0(ori_ori_n194_), .Y(ori_ori_n195_));
  AOI220     o173(.A0(ori_ori_n195_), .A1(ori_ori_n136_), .B0(ori_ori_n187_), .B1(ori_ori_n185_), .Y(ori_ori_n196_));
  NO2        o174(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n197_));
  OR2        o175(.A(i_8_), .B(i_7_), .Y(ori_ori_n198_));
  INV        o176(.A(i_12_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n44_), .B(ori_ori_n199_), .Y(ori_ori_n200_));
  NO3        o178(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n201_));
  NA2        o179(.A(i_2_), .B(i_1_), .Y(ori_ori_n202_));
  NO3        o180(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n203_));
  NAi21      o181(.An(i_4_), .B(i_3_), .Y(ori_ori_n204_));
  NO2        o182(.A(i_0_), .B(i_6_), .Y(ori_ori_n205_));
  NOi41      o183(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n202_), .B(ori_ori_n159_), .Y(ori_ori_n207_));
  NO2        o185(.A(i_11_), .B(ori_ori_n192_), .Y(ori_ori_n208_));
  NOi21      o186(.An(i_1_), .B(i_6_), .Y(ori_ori_n209_));
  NAi21      o187(.An(i_3_), .B(i_7_), .Y(ori_ori_n210_));
  NA2        o188(.A(ori_ori_n199_), .B(i_9_), .Y(ori_ori_n211_));
  OR4        o189(.A(ori_ori_n211_), .B(ori_ori_n210_), .C(ori_ori_n209_), .D(ori_ori_n160_), .Y(ori_ori_n212_));
  NO2        o190(.A(i_12_), .B(i_3_), .Y(ori_ori_n213_));
  NA2        o191(.A(ori_ori_n69_), .B(i_5_), .Y(ori_ori_n214_));
  NA2        o192(.A(i_3_), .B(i_9_), .Y(ori_ori_n215_));
  NAi21      o193(.An(i_7_), .B(i_10_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n216_), .B(ori_ori_n215_), .Y(ori_ori_n217_));
  NA3        o195(.A(ori_ori_n217_), .B(ori_ori_n214_), .C(ori_ori_n60_), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n218_), .B(ori_ori_n212_), .Y(ori_ori_n219_));
  INV        o197(.A(ori_ori_n137_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n199_), .B(i_13_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n221_), .B(ori_ori_n71_), .Y(ori_ori_n222_));
  AOI220     o200(.A0(ori_ori_n222_), .A1(ori_ori_n220_), .B0(ori_ori_n219_), .B1(ori_ori_n208_), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n198_), .B(ori_ori_n37_), .Y(ori_ori_n224_));
  NA2        o202(.A(i_12_), .B(i_6_), .Y(ori_ori_n225_));
  OR2        o203(.A(i_13_), .B(i_9_), .Y(ori_ori_n226_));
  NO3        o204(.A(ori_ori_n226_), .B(ori_ori_n225_), .C(ori_ori_n48_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n204_), .B(i_2_), .Y(ori_ori_n228_));
  NA3        o206(.A(ori_ori_n228_), .B(ori_ori_n227_), .C(ori_ori_n44_), .Y(ori_ori_n229_));
  NA2        o207(.A(ori_ori_n208_), .B(i_9_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n214_), .B(ori_ori_n60_), .Y(ori_ori_n231_));
  OAI210     o209(.A0(ori_ori_n231_), .A1(ori_ori_n230_), .B0(ori_ori_n229_), .Y(ori_ori_n232_));
  NO3        o210(.A(i_11_), .B(ori_ori_n192_), .C(ori_ori_n25_), .Y(ori_ori_n233_));
  NO2        o211(.A(ori_ori_n210_), .B(i_8_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n232_), .B(ori_ori_n224_), .Y(ori_ori_n235_));
  NA3        o213(.A(ori_ori_n235_), .B(ori_ori_n223_), .C(ori_ori_n196_), .Y(ori_ori_n236_));
  NO3        o214(.A(i_12_), .B(ori_ori_n192_), .C(ori_ori_n37_), .Y(ori_ori_n237_));
  INV        o215(.A(ori_ori_n237_), .Y(ori_ori_n238_));
  NO3        o216(.A(i_0_), .B(i_2_), .C(ori_ori_n59_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n202_), .B(i_0_), .Y(ori_ori_n240_));
  AOI220     o218(.A0(ori_ori_n240_), .A1(ori_ori_n167_), .B0(ori_ori_n239_), .B1(ori_ori_n136_), .Y(ori_ori_n241_));
  NA2        o219(.A(i_5_), .B(ori_ori_n26_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n242_), .B(ori_ori_n241_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n151_), .B(ori_ori_n137_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n244_), .B(ori_ori_n243_), .Y(ori_ori_n245_));
  NO2        o223(.A(i_3_), .B(i_10_), .Y(ori_ori_n246_));
  NO2        o224(.A(i_2_), .B(ori_ori_n95_), .Y(ori_ori_n247_));
  AN2        o225(.A(i_3_), .B(i_10_), .Y(ori_ori_n248_));
  NO2        o226(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n249_));
  NO2        o227(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n245_), .B(ori_ori_n238_), .Y(ori_ori_n251_));
  NO3        o229(.A(ori_ori_n251_), .B(ori_ori_n236_), .C(ori_ori_n182_), .Y(ori_ori_n252_));
  NO3        o230(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n253_));
  NO3        o231(.A(i_6_), .B(ori_ori_n166_), .C(i_7_), .Y(ori_ori_n254_));
  NO2        o232(.A(i_2_), .B(i_3_), .Y(ori_ori_n255_));
  OR2        o233(.A(i_0_), .B(i_5_), .Y(ori_ori_n256_));
  NO2        o234(.A(ori_ori_n146_), .B(ori_ori_n46_), .Y(ori_ori_n257_));
  NO2        o235(.A(i_12_), .B(i_10_), .Y(ori_ori_n258_));
  NOi21      o236(.An(i_5_), .B(i_0_), .Y(ori_ori_n259_));
  NO2        o237(.A(i_2_), .B(ori_ori_n95_), .Y(ori_ori_n260_));
  NO4        o238(.A(ori_ori_n260_), .B(i_4_), .C(ori_ori_n259_), .D(ori_ori_n123_), .Y(ori_ori_n261_));
  NA4        o239(.A(ori_ori_n79_), .B(ori_ori_n36_), .C(ori_ori_n80_), .D(i_8_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n261_), .B(ori_ori_n258_), .Y(ori_ori_n263_));
  NO2        o241(.A(i_6_), .B(i_8_), .Y(ori_ori_n264_));
  NOi21      o242(.An(i_0_), .B(i_2_), .Y(ori_ori_n265_));
  AN2        o243(.A(ori_ori_n265_), .B(ori_ori_n264_), .Y(ori_ori_n266_));
  NO2        o244(.A(i_1_), .B(i_7_), .Y(ori_ori_n267_));
  INV        o245(.A(ori_ori_n263_), .Y(ori_ori_n268_));
  NA3        o246(.A(ori_ori_n209_), .B(ori_ori_n247_), .C(ori_ori_n166_), .Y(ori_ori_n269_));
  NO2        o247(.A(ori_ori_n166_), .B(i_9_), .Y(ori_ori_n270_));
  NA2        o248(.A(ori_ori_n270_), .B(ori_ori_n175_), .Y(ori_ori_n271_));
  INV        o249(.A(ori_ori_n243_), .Y(ori_ori_n272_));
  AOI210     o250(.A0(ori_ori_n272_), .A1(ori_ori_n269_), .B0(ori_ori_n149_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n268_), .A1(ori_ori_n253_), .B0(ori_ori_n273_), .Y(ori_ori_n274_));
  NOi32      o252(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n275_));
  INV        o253(.A(ori_ori_n275_), .Y(ori_ori_n276_));
  NAi21      o254(.An(i_0_), .B(i_6_), .Y(ori_ori_n277_));
  NAi21      o255(.An(i_1_), .B(i_5_), .Y(ori_ori_n278_));
  NA2        o256(.A(ori_ori_n278_), .B(ori_ori_n277_), .Y(ori_ori_n279_));
  NA2        o257(.A(ori_ori_n279_), .B(ori_ori_n25_), .Y(ori_ori_n280_));
  NO2        o258(.A(ori_ori_n280_), .B(ori_ori_n147_), .Y(ori_ori_n281_));
  NAi41      o259(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n282_));
  OAI220     o260(.A0(ori_ori_n282_), .A1(ori_ori_n278_), .B0(ori_ori_n188_), .B1(ori_ori_n147_), .Y(ori_ori_n283_));
  AOI210     o261(.A0(ori_ori_n282_), .A1(ori_ori_n147_), .B0(ori_ori_n146_), .Y(ori_ori_n284_));
  NOi32      o262(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n285_));
  NAi21      o263(.An(i_6_), .B(i_1_), .Y(ori_ori_n286_));
  NA3        o264(.A(ori_ori_n286_), .B(ori_ori_n285_), .C(ori_ori_n46_), .Y(ori_ori_n287_));
  NO2        o265(.A(ori_ori_n287_), .B(i_0_), .Y(ori_ori_n288_));
  OR3        o266(.A(ori_ori_n288_), .B(ori_ori_n284_), .C(ori_ori_n283_), .Y(ori_ori_n289_));
  NO2        o267(.A(i_1_), .B(ori_ori_n95_), .Y(ori_ori_n290_));
  NAi21      o268(.An(i_3_), .B(i_4_), .Y(ori_ori_n291_));
  NO2        o269(.A(ori_ori_n291_), .B(i_9_), .Y(ori_ori_n292_));
  AN2        o270(.A(i_6_), .B(i_7_), .Y(ori_ori_n293_));
  OAI210     o271(.A0(ori_ori_n293_), .A1(ori_ori_n290_), .B0(ori_ori_n292_), .Y(ori_ori_n294_));
  NA2        o272(.A(i_2_), .B(i_7_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n291_), .B(i_10_), .Y(ori_ori_n296_));
  NA3        o274(.A(ori_ori_n296_), .B(ori_ori_n295_), .C(ori_ori_n205_), .Y(ori_ori_n297_));
  AOI210     o275(.A0(ori_ori_n297_), .A1(ori_ori_n294_), .B0(ori_ori_n160_), .Y(ori_ori_n298_));
  AOI210     o276(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n299_));
  OAI210     o277(.A0(ori_ori_n299_), .A1(ori_ori_n163_), .B0(ori_ori_n296_), .Y(ori_ori_n300_));
  AOI220     o278(.A0(ori_ori_n296_), .A1(ori_ori_n267_), .B0(ori_ori_n201_), .B1(ori_ori_n163_), .Y(ori_ori_n301_));
  AOI210     o279(.A0(ori_ori_n301_), .A1(ori_ori_n300_), .B0(i_5_), .Y(ori_ori_n302_));
  NO4        o280(.A(ori_ori_n302_), .B(ori_ori_n298_), .C(ori_ori_n289_), .D(ori_ori_n281_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n303_), .B(ori_ori_n276_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n57_), .B(ori_ori_n25_), .Y(ori_ori_n305_));
  AN2        o283(.A(i_12_), .B(i_5_), .Y(ori_ori_n306_));
  NA2        o284(.A(ori_ori_n829_), .B(ori_ori_n306_), .Y(ori_ori_n307_));
  NO2        o285(.A(i_11_), .B(i_6_), .Y(ori_ori_n308_));
  NA3        o286(.A(ori_ori_n308_), .B(ori_ori_n257_), .C(ori_ori_n192_), .Y(ori_ori_n309_));
  NO2        o287(.A(ori_ori_n309_), .B(ori_ori_n307_), .Y(ori_ori_n310_));
  NO2        o288(.A(i_5_), .B(i_10_), .Y(ori_ori_n311_));
  NA2        o289(.A(ori_ori_n311_), .B(ori_ori_n228_), .Y(ori_ori_n312_));
  NA2        o290(.A(ori_ori_n138_), .B(ori_ori_n45_), .Y(ori_ori_n313_));
  NO2        o291(.A(ori_ori_n313_), .B(ori_ori_n312_), .Y(ori_ori_n314_));
  OAI210     o292(.A0(ori_ori_n314_), .A1(ori_ori_n310_), .B0(ori_ori_n305_), .Y(ori_ori_n315_));
  NO2        o293(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n316_));
  NO2        o294(.A(ori_ori_n144_), .B(ori_ori_n80_), .Y(ori_ori_n317_));
  OAI210     o295(.A0(ori_ori_n317_), .A1(ori_ori_n310_), .B0(ori_ori_n316_), .Y(ori_ori_n318_));
  NO3        o296(.A(ori_ori_n80_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n319_));
  NA3        o297(.A(ori_ori_n246_), .B(ori_ori_n71_), .C(ori_ori_n54_), .Y(ori_ori_n320_));
  NO2        o298(.A(i_11_), .B(i_12_), .Y(ori_ori_n321_));
  NA2        o299(.A(ori_ori_n321_), .B(ori_ori_n36_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n320_), .B(ori_ori_n322_), .Y(ori_ori_n323_));
  NA2        o301(.A(ori_ori_n311_), .B(ori_ori_n199_), .Y(ori_ori_n324_));
  NAi21      o302(.An(i_13_), .B(i_0_), .Y(ori_ori_n325_));
  NO2        o303(.A(ori_ori_n325_), .B(ori_ori_n202_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n323_), .B(ori_ori_n326_), .Y(ori_ori_n327_));
  NA3        o305(.A(ori_ori_n327_), .B(ori_ori_n318_), .C(ori_ori_n315_), .Y(ori_ori_n328_));
  NA2        o306(.A(ori_ori_n44_), .B(ori_ori_n192_), .Y(ori_ori_n329_));
  NO3        o307(.A(i_1_), .B(i_12_), .C(ori_ori_n80_), .Y(ori_ori_n330_));
  NO2        o308(.A(i_0_), .B(i_11_), .Y(ori_ori_n331_));
  NOi21      o309(.An(i_2_), .B(i_12_), .Y(ori_ori_n332_));
  OR2        o310(.A(i_13_), .B(i_10_), .Y(ori_ori_n333_));
  NO2        o311(.A(ori_ori_n154_), .B(ori_ori_n118_), .Y(ori_ori_n334_));
  NO2        o312(.A(ori_ori_n95_), .B(ori_ori_n25_), .Y(ori_ori_n335_));
  NO2        o313(.A(ori_ori_n159_), .B(ori_ori_n80_), .Y(ori_ori_n336_));
  NA2        o314(.A(ori_ori_n166_), .B(i_10_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n214_), .B(ori_ori_n60_), .C(i_2_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n338_), .B(ori_ori_n337_), .Y(ori_ori_n339_));
  NO2        o317(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n340_));
  NA3        o318(.A(ori_ori_n267_), .B(ori_ori_n266_), .C(ori_ori_n340_), .Y(ori_ori_n341_));
  INV        o319(.A(ori_ori_n254_), .Y(ori_ori_n342_));
  OAI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n164_), .B0(ori_ori_n341_), .Y(ori_ori_n343_));
  NO2        o321(.A(ori_ori_n343_), .B(ori_ori_n339_), .Y(ori_ori_n344_));
  NO2        o322(.A(ori_ori_n344_), .B(ori_ori_n230_), .Y(ori_ori_n345_));
  NO3        o323(.A(ori_ori_n345_), .B(ori_ori_n328_), .C(ori_ori_n304_), .Y(ori_ori_n346_));
  NO2        o324(.A(ori_ori_n69_), .B(i_13_), .Y(ori_ori_n347_));
  NO2        o325(.A(i_10_), .B(i_9_), .Y(ori_ori_n348_));
  NAi21      o326(.An(i_12_), .B(i_8_), .Y(ori_ori_n349_));
  NO2        o327(.A(ori_ori_n349_), .B(i_3_), .Y(ori_ori_n350_));
  NO2        o328(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n351_));
  NA2        o329(.A(ori_ori_n351_), .B(ori_ori_n98_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n174_), .Y(ori_ori_n353_));
  NA2        o331(.A(ori_ori_n250_), .B(i_0_), .Y(ori_ori_n354_));
  NO3        o332(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n355_));
  NA2        o333(.A(ori_ori_n225_), .B(ori_ori_n93_), .Y(ori_ori_n356_));
  NA2        o334(.A(ori_ori_n356_), .B(ori_ori_n355_), .Y(ori_ori_n357_));
  NA2        o335(.A(i_8_), .B(i_9_), .Y(ori_ori_n358_));
  AOI210     o336(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n359_));
  OR2        o337(.A(ori_ori_n359_), .B(ori_ori_n358_), .Y(ori_ori_n360_));
  NA2        o338(.A(ori_ori_n237_), .B(ori_ori_n175_), .Y(ori_ori_n361_));
  OAI220     o339(.A0(ori_ori_n361_), .A1(ori_ori_n360_), .B0(ori_ori_n357_), .B1(ori_ori_n354_), .Y(ori_ori_n362_));
  NA2        o340(.A(ori_ori_n208_), .B(ori_ori_n249_), .Y(ori_ori_n363_));
  NO3        o341(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n364_));
  INV        o342(.A(ori_ori_n364_), .Y(ori_ori_n365_));
  NA3        o343(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n366_));
  NA4        o344(.A(ori_ori_n139_), .B(ori_ori_n110_), .C(ori_ori_n76_), .D(ori_ori_n23_), .Y(ori_ori_n367_));
  OAI220     o345(.A0(ori_ori_n367_), .A1(ori_ori_n366_), .B0(ori_ori_n365_), .B1(ori_ori_n363_), .Y(ori_ori_n368_));
  NO3        o346(.A(ori_ori_n368_), .B(ori_ori_n362_), .C(ori_ori_n353_), .Y(ori_ori_n369_));
  OR2        o347(.A(ori_ori_n271_), .B(ori_ori_n149_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n92_), .B(i_13_), .Y(ori_ori_n371_));
  NA2        o349(.A(ori_ori_n336_), .B(ori_ori_n305_), .Y(ori_ori_n372_));
  NO2        o350(.A(i_2_), .B(i_13_), .Y(ori_ori_n373_));
  NO2        o351(.A(ori_ori_n372_), .B(ori_ori_n371_), .Y(ori_ori_n374_));
  NO3        o352(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n375_));
  NO2        o353(.A(i_6_), .B(i_7_), .Y(ori_ori_n376_));
  NO2        o354(.A(i_11_), .B(i_1_), .Y(ori_ori_n377_));
  OR2        o355(.A(i_11_), .B(i_8_), .Y(ori_ori_n378_));
  NOi21      o356(.An(i_2_), .B(i_7_), .Y(ori_ori_n379_));
  NO2        o357(.A(i_3_), .B(ori_ori_n166_), .Y(ori_ori_n380_));
  NO2        o358(.A(i_6_), .B(i_10_), .Y(ori_ori_n381_));
  NA3        o359(.A(ori_ori_n206_), .B(ori_ori_n153_), .C(ori_ori_n127_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n383_));
  NO2        o361(.A(ori_ori_n146_), .B(i_3_), .Y(ori_ori_n384_));
  NAi31      o362(.An(ori_ori_n383_), .B(ori_ori_n384_), .C(ori_ori_n193_), .Y(ori_ori_n385_));
  NA3        o363(.A(ori_ori_n316_), .B(ori_ori_n158_), .C(ori_ori_n143_), .Y(ori_ori_n386_));
  NA3        o364(.A(ori_ori_n386_), .B(ori_ori_n385_), .C(ori_ori_n382_), .Y(ori_ori_n387_));
  NO2        o365(.A(ori_ori_n387_), .B(ori_ori_n374_), .Y(ori_ori_n388_));
  NA2        o366(.A(ori_ori_n355_), .B(ori_ori_n306_), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n364_), .B(ori_ori_n311_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n390_), .B(ori_ori_n191_), .Y(ori_ori_n391_));
  NAi21      o369(.An(ori_ori_n184_), .B(ori_ori_n321_), .Y(ori_ori_n392_));
  NA2        o370(.A(ori_ori_n267_), .B(ori_ori_n186_), .Y(ori_ori_n393_));
  NO2        o371(.A(ori_ori_n393_), .B(ori_ori_n392_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n253_), .B(ori_ori_n201_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n395_), .B(ori_ori_n338_), .Y(ori_ori_n396_));
  NO3        o374(.A(ori_ori_n396_), .B(ori_ori_n394_), .C(ori_ori_n391_), .Y(ori_ori_n397_));
  NA4        o375(.A(ori_ori_n397_), .B(ori_ori_n388_), .C(ori_ori_n370_), .D(ori_ori_n369_), .Y(ori_ori_n398_));
  NA2        o376(.A(ori_ori_n117_), .B(ori_ori_n106_), .Y(ori_ori_n399_));
  AN2        o377(.A(ori_ori_n399_), .B(ori_ori_n355_), .Y(ori_ori_n400_));
  NA2        o378(.A(ori_ori_n400_), .B(ori_ori_n250_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n275_), .B(ori_ori_n69_), .Y(ori_ori_n402_));
  NO2        o380(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n403_));
  NA2        o381(.A(ori_ori_n39_), .B(i_13_), .Y(ori_ori_n404_));
  OAI210     o382(.A0(i_8_), .A1(ori_ori_n59_), .B0(ori_ori_n129_), .Y(ori_ori_n405_));
  NA2        o383(.A(ori_ori_n405_), .B(ori_ori_n334_), .Y(ori_ori_n406_));
  NA3        o384(.A(ori_ori_n406_), .B(ori_ori_n404_), .C(ori_ori_n401_), .Y(ori_ori_n407_));
  NO2        o385(.A(i_12_), .B(ori_ori_n166_), .Y(ori_ori_n408_));
  NO2        o386(.A(i_8_), .B(i_7_), .Y(ori_ori_n409_));
  AOI220     o387(.A0(ori_ori_n336_), .A1(ori_ori_n257_), .B0(ori_ori_n207_), .B1(ori_ori_n205_), .Y(ori_ori_n410_));
  OAI220     o388(.A0(ori_ori_n410_), .A1(ori_ori_n221_), .B0(ori_ori_n371_), .B1(ori_ori_n128_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n411_), .B(ori_ori_n224_), .Y(ori_ori_n412_));
  NA3        o390(.A(ori_ori_n248_), .B(ori_ori_n155_), .C(ori_ori_n92_), .Y(ori_ori_n413_));
  NO2        o391(.A(ori_ori_n146_), .B(i_5_), .Y(ori_ori_n414_));
  NA3        o392(.A(ori_ori_n414_), .B(ori_ori_n329_), .C(ori_ori_n255_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(ori_ori_n413_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n416_), .B(ori_ori_n364_), .Y(ori_ori_n417_));
  NA2        o395(.A(ori_ori_n417_), .B(ori_ori_n412_), .Y(ori_ori_n418_));
  AOI210     o396(.A0(ori_ori_n286_), .A1(ori_ori_n46_), .B0(ori_ori_n290_), .Y(ori_ori_n419_));
  NA2        o397(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n420_));
  NA3        o398(.A(ori_ori_n408_), .B(ori_ori_n233_), .C(ori_ori_n420_), .Y(ori_ori_n421_));
  NO2        o399(.A(ori_ori_n419_), .B(ori_ori_n421_), .Y(ori_ori_n422_));
  INV        o400(.A(ori_ori_n422_), .Y(ori_ori_n423_));
  NO4        o401(.A(ori_ori_n209_), .B(ori_ori_n42_), .C(i_2_), .D(ori_ori_n48_), .Y(ori_ori_n424_));
  NO3        o402(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n198_), .B(ori_ori_n36_), .Y(ori_ori_n426_));
  NO2        o404(.A(ori_ori_n333_), .B(i_1_), .Y(ori_ori_n427_));
  NOi31      o405(.An(ori_ori_n427_), .B(ori_ori_n356_), .C(ori_ori_n69_), .Y(ori_ori_n428_));
  NOi21      o406(.An(i_10_), .B(i_6_), .Y(ori_ori_n429_));
  NO2        o407(.A(ori_ori_n80_), .B(ori_ori_n25_), .Y(ori_ori_n430_));
  AOI220     o408(.A0(ori_ori_n237_), .A1(ori_ori_n430_), .B0(ori_ori_n233_), .B1(ori_ori_n429_), .Y(ori_ori_n431_));
  NO2        o409(.A(ori_ori_n431_), .B(ori_ori_n354_), .Y(ori_ori_n432_));
  NO2        o410(.A(ori_ori_n109_), .B(ori_ori_n23_), .Y(ori_ori_n433_));
  NOi21      o411(.An(ori_ori_n140_), .B(ori_ori_n262_), .Y(ori_ori_n434_));
  NO2        o412(.A(ori_ori_n434_), .B(ori_ori_n432_), .Y(ori_ori_n435_));
  NO2        o413(.A(ori_ori_n402_), .B(ori_ori_n301_), .Y(ori_ori_n436_));
  INV        o414(.A(ori_ori_n255_), .Y(ori_ori_n437_));
  NO2        o415(.A(i_12_), .B(ori_ori_n80_), .Y(ori_ori_n438_));
  NA3        o416(.A(ori_ori_n438_), .B(ori_ori_n233_), .C(ori_ori_n420_), .Y(ori_ori_n439_));
  NA3        o417(.A(ori_ori_n308_), .B(ori_ori_n237_), .C(ori_ori_n186_), .Y(ori_ori_n440_));
  AOI210     o418(.A0(ori_ori_n440_), .A1(ori_ori_n439_), .B0(ori_ori_n437_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n295_), .B(ori_ori_n205_), .Y(ori_ori_n442_));
  NO2        o420(.A(ori_ori_n442_), .B(ori_ori_n392_), .Y(ori_ori_n443_));
  NO3        o421(.A(ori_ori_n443_), .B(ori_ori_n441_), .C(ori_ori_n436_), .Y(ori_ori_n444_));
  NA3        o422(.A(ori_ori_n444_), .B(ori_ori_n435_), .C(ori_ori_n423_), .Y(ori_ori_n445_));
  NO4        o423(.A(ori_ori_n445_), .B(ori_ori_n418_), .C(ori_ori_n407_), .D(ori_ori_n398_), .Y(ori_ori_n446_));
  NA4        o424(.A(ori_ori_n446_), .B(ori_ori_n346_), .C(ori_ori_n274_), .D(ori_ori_n252_), .Y(ori7));
  NO2        o425(.A(ori_ori_n88_), .B(ori_ori_n54_), .Y(ori_ori_n448_));
  NO2        o426(.A(ori_ori_n102_), .B(ori_ori_n85_), .Y(ori_ori_n449_));
  NA2        o427(.A(ori_ori_n829_), .B(ori_ori_n449_), .Y(ori_ori_n450_));
  NA2        o428(.A(ori_ori_n381_), .B(ori_ori_n79_), .Y(ori_ori_n451_));
  NA2        o429(.A(i_11_), .B(ori_ori_n166_), .Y(ori_ori_n452_));
  NA2        o430(.A(ori_ori_n138_), .B(ori_ori_n452_), .Y(ori_ori_n453_));
  OAI210     o431(.A0(ori_ori_n453_), .A1(ori_ori_n451_), .B0(ori_ori_n450_), .Y(ori_ori_n454_));
  NO2        o432(.A(ori_ori_n199_), .B(i_4_), .Y(ori_ori_n455_));
  NA2        o433(.A(ori_ori_n455_), .B(i_8_), .Y(ori_ori_n456_));
  NA2        o434(.A(i_2_), .B(ori_ori_n80_), .Y(ori_ori_n457_));
  OAI210     o435(.A0(ori_ori_n83_), .A1(ori_ori_n172_), .B0(ori_ori_n173_), .Y(ori_ori_n458_));
  NO2        o436(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n459_));
  NA2        o437(.A(i_4_), .B(i_8_), .Y(ori_ori_n460_));
  AOI210     o438(.A0(ori_ori_n460_), .A1(ori_ori_n248_), .B0(ori_ori_n459_), .Y(ori_ori_n461_));
  OAI220     o439(.A0(ori_ori_n461_), .A1(ori_ori_n457_), .B0(ori_ori_n458_), .B1(i_13_), .Y(ori_ori_n462_));
  NO3        o440(.A(ori_ori_n462_), .B(ori_ori_n454_), .C(ori_ori_n448_), .Y(ori_ori_n463_));
  AOI210     o441(.A0(ori_ori_n123_), .A1(ori_ori_n58_), .B0(i_10_), .Y(ori_ori_n464_));
  AOI210     o442(.A0(ori_ori_n464_), .A1(ori_ori_n199_), .B0(ori_ori_n148_), .Y(ori_ori_n465_));
  OR2        o443(.A(i_6_), .B(i_10_), .Y(ori_ori_n466_));
  INV        o444(.A(ori_ori_n171_), .Y(ori_ori_n467_));
  OR2        o445(.A(ori_ori_n465_), .B(ori_ori_n226_), .Y(ori_ori_n468_));
  AOI210     o446(.A0(ori_ori_n468_), .A1(ori_ori_n463_), .B0(ori_ori_n59_), .Y(ori_ori_n469_));
  NOi21      o447(.An(i_11_), .B(i_7_), .Y(ori_ori_n470_));
  AO210      o448(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n471_));
  NO2        o449(.A(ori_ori_n471_), .B(ori_ori_n470_), .Y(ori_ori_n472_));
  NA2        o450(.A(ori_ori_n472_), .B(ori_ori_n177_), .Y(ori_ori_n473_));
  NA3        o451(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n474_));
  NAi31      o452(.An(ori_ori_n474_), .B(ori_ori_n183_), .C(i_11_), .Y(ori_ori_n475_));
  AOI210     o453(.A0(ori_ori_n475_), .A1(ori_ori_n473_), .B0(ori_ori_n59_), .Y(ori_ori_n476_));
  NA2        o454(.A(ori_ori_n82_), .B(ori_ori_n59_), .Y(ori_ori_n477_));
  AO210      o455(.A0(ori_ori_n477_), .A1(ori_ori_n301_), .B0(ori_ori_n41_), .Y(ori_ori_n478_));
  NO3        o456(.A(ori_ori_n216_), .B(ori_ori_n178_), .C(ori_ori_n452_), .Y(ori_ori_n479_));
  OAI210     o457(.A0(ori_ori_n479_), .A1(ori_ori_n193_), .B0(ori_ori_n59_), .Y(ori_ori_n480_));
  NA2        o458(.A(ori_ori_n332_), .B(ori_ori_n31_), .Y(ori_ori_n481_));
  OR2        o459(.A(ori_ori_n178_), .B(ori_ori_n102_), .Y(ori_ori_n482_));
  NA2        o460(.A(ori_ori_n482_), .B(ori_ori_n481_), .Y(ori_ori_n483_));
  NO2        o461(.A(ori_ori_n59_), .B(i_9_), .Y(ori_ori_n484_));
  NO2        o462(.A(ori_ori_n484_), .B(i_4_), .Y(ori_ori_n485_));
  NA2        o463(.A(ori_ori_n485_), .B(ori_ori_n483_), .Y(ori_ori_n486_));
  NO2        o464(.A(i_1_), .B(i_12_), .Y(ori_ori_n487_));
  NA3        o465(.A(ori_ori_n487_), .B(ori_ori_n104_), .C(ori_ori_n24_), .Y(ori_ori_n488_));
  BUFFER     o466(.A(ori_ori_n488_), .Y(ori_ori_n489_));
  NA4        o467(.A(ori_ori_n489_), .B(ori_ori_n486_), .C(ori_ori_n480_), .D(ori_ori_n478_), .Y(ori_ori_n490_));
  OAI210     o468(.A0(ori_ori_n490_), .A1(ori_ori_n476_), .B0(i_6_), .Y(ori_ori_n491_));
  NO2        o469(.A(ori_ori_n474_), .B(ori_ori_n102_), .Y(ori_ori_n492_));
  NA2        o470(.A(ori_ori_n492_), .B(ori_ori_n438_), .Y(ori_ori_n493_));
  NO2        o471(.A(ori_ori_n199_), .B(ori_ori_n80_), .Y(ori_ori_n494_));
  NO2        o472(.A(ori_ori_n494_), .B(i_11_), .Y(ori_ori_n495_));
  NA2        o473(.A(ori_ori_n493_), .B(ori_ori_n357_), .Y(ori_ori_n496_));
  NO3        o474(.A(ori_ori_n466_), .B(ori_ori_n198_), .C(ori_ori_n23_), .Y(ori_ori_n497_));
  AOI210     o475(.A0(i_1_), .A1(ori_ori_n217_), .B0(ori_ori_n497_), .Y(ori_ori_n498_));
  NO2        o476(.A(ori_ori_n498_), .B(ori_ori_n44_), .Y(ori_ori_n499_));
  NA3        o477(.A(ori_ori_n409_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n500_));
  INV        o478(.A(i_2_), .Y(ori_ori_n501_));
  NA2        o479(.A(ori_ori_n133_), .B(i_9_), .Y(ori_ori_n502_));
  NA3        o480(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n504_));
  NA3        o482(.A(ori_ori_n504_), .B(ori_ori_n225_), .C(ori_ori_n44_), .Y(ori_ori_n505_));
  OAI220     o483(.A0(ori_ori_n505_), .A1(ori_ori_n503_), .B0(ori_ori_n502_), .B1(ori_ori_n501_), .Y(ori_ori_n506_));
  NA3        o484(.A(ori_ori_n484_), .B(ori_ori_n255_), .C(i_6_), .Y(ori_ori_n507_));
  NO2        o485(.A(ori_ori_n507_), .B(ori_ori_n23_), .Y(ori_ori_n508_));
  AOI210     o486(.A0(ori_ori_n377_), .A1(ori_ori_n335_), .B0(ori_ori_n203_), .Y(ori_ori_n509_));
  NO2        o487(.A(ori_ori_n509_), .B(ori_ori_n457_), .Y(ori_ori_n510_));
  NO2        o488(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n511_));
  OR3        o489(.A(ori_ori_n510_), .B(ori_ori_n508_), .C(ori_ori_n506_), .Y(ori_ori_n512_));
  NO3        o490(.A(ori_ori_n512_), .B(ori_ori_n499_), .C(ori_ori_n496_), .Y(ori_ori_n513_));
  NO2        o491(.A(ori_ori_n199_), .B(ori_ori_n95_), .Y(ori_ori_n514_));
  NO2        o492(.A(ori_ori_n514_), .B(ori_ori_n470_), .Y(ori_ori_n515_));
  NO2        o493(.A(ori_ori_n198_), .B(ori_ori_n44_), .Y(ori_ori_n516_));
  NO3        o494(.A(ori_ori_n516_), .B(ori_ori_n250_), .C(ori_ori_n200_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n112_), .B(ori_ori_n37_), .Y(ori_ori_n518_));
  NO2        o496(.A(ori_ori_n518_), .B(i_6_), .Y(ori_ori_n519_));
  NO2        o497(.A(ori_ori_n80_), .B(i_9_), .Y(ori_ori_n520_));
  NO2        o498(.A(ori_ori_n520_), .B(ori_ori_n59_), .Y(ori_ori_n521_));
  NO2        o499(.A(ori_ori_n521_), .B(ori_ori_n487_), .Y(ori_ori_n522_));
  NO4        o500(.A(ori_ori_n522_), .B(ori_ori_n519_), .C(ori_ori_n517_), .D(i_4_), .Y(ori_ori_n523_));
  NA2        o501(.A(i_1_), .B(i_3_), .Y(ori_ori_n524_));
  INV        o502(.A(ori_ori_n523_), .Y(ori_ori_n525_));
  NA3        o503(.A(ori_ori_n525_), .B(ori_ori_n513_), .C(ori_ori_n491_), .Y(ori_ori_n526_));
  NO3        o504(.A(ori_ori_n378_), .B(i_3_), .C(i_7_), .Y(ori_ori_n527_));
  NOi21      o505(.An(ori_ori_n527_), .B(i_10_), .Y(ori_ori_n528_));
  OA210      o506(.A0(ori_ori_n528_), .A1(ori_ori_n206_), .B0(ori_ori_n80_), .Y(ori_ori_n529_));
  NA3        o507(.A(ori_ori_n381_), .B(ori_ori_n403_), .C(ori_ori_n46_), .Y(ori_ori_n530_));
  NO3        o508(.A(ori_ori_n379_), .B(ori_ori_n460_), .C(ori_ori_n80_), .Y(ori_ori_n531_));
  NA2        o509(.A(ori_ori_n531_), .B(ori_ori_n25_), .Y(ori_ori_n532_));
  NA3        o510(.A(ori_ori_n148_), .B(ori_ori_n79_), .C(ori_ori_n80_), .Y(ori_ori_n533_));
  NA3        o511(.A(ori_ori_n533_), .B(ori_ori_n532_), .C(ori_ori_n530_), .Y(ori_ori_n534_));
  OAI210     o512(.A0(ori_ori_n534_), .A1(ori_ori_n529_), .B0(i_1_), .Y(ori_ori_n535_));
  AOI210     o513(.A0(ori_ori_n225_), .A1(ori_ori_n93_), .B0(i_1_), .Y(ori_ori_n536_));
  NO2        o514(.A(ori_ori_n291_), .B(i_2_), .Y(ori_ori_n537_));
  NA2        o515(.A(ori_ori_n537_), .B(ori_ori_n536_), .Y(ori_ori_n538_));
  OAI210     o516(.A0(ori_ori_n507_), .A1(ori_ori_n349_), .B0(ori_ori_n538_), .Y(ori_ori_n539_));
  INV        o517(.A(ori_ori_n539_), .Y(ori_ori_n540_));
  AOI210     o518(.A0(ori_ori_n540_), .A1(ori_ori_n535_), .B0(i_13_), .Y(ori_ori_n541_));
  NA2        o519(.A(ori_ori_n100_), .B(ori_ori_n133_), .Y(ori_ori_n542_));
  AOI220     o520(.A0(ori_ori_n373_), .A1(ori_ori_n148_), .B0(ori_ori_n351_), .B1(ori_ori_n133_), .Y(ori_ori_n543_));
  OAI210     o521(.A0(ori_ori_n543_), .A1(ori_ori_n44_), .B0(ori_ori_n542_), .Y(ori_ori_n544_));
  NO2        o522(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n545_));
  NO2        o523(.A(ori_ori_n379_), .B(ori_ori_n24_), .Y(ori_ori_n546_));
  NO2        o524(.A(ori_ori_n827_), .B(ori_ori_n88_), .Y(ori_ori_n547_));
  AOI210     o525(.A0(ori_ori_n544_), .A1(ori_ori_n264_), .B0(ori_ori_n547_), .Y(ori_ori_n548_));
  INV        o526(.A(ori_ori_n109_), .Y(ori_ori_n549_));
  AOI220     o527(.A0(ori_ori_n549_), .A1(ori_ori_n68_), .B0(ori_ori_n308_), .B1(ori_ori_n504_), .Y(ori_ori_n550_));
  NO2        o528(.A(ori_ori_n550_), .B(ori_ori_n204_), .Y(ori_ori_n551_));
  AOI210     o529(.A0(ori_ori_n349_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n552_));
  NOi31      o530(.An(ori_ori_n552_), .B(ori_ori_n451_), .C(ori_ori_n44_), .Y(ori_ori_n553_));
  NA2        o531(.A(ori_ori_n122_), .B(i_13_), .Y(ori_ori_n554_));
  NO2        o532(.A(ori_ori_n503_), .B(ori_ori_n109_), .Y(ori_ori_n555_));
  INV        o533(.A(ori_ori_n555_), .Y(ori_ori_n556_));
  OAI220     o534(.A0(ori_ori_n556_), .A1(ori_ori_n67_), .B0(ori_ori_n554_), .B1(ori_ori_n536_), .Y(ori_ori_n557_));
  NO3        o535(.A(ori_ori_n67_), .B(ori_ori_n32_), .C(ori_ori_n95_), .Y(ori_ori_n558_));
  NA2        o536(.A(ori_ori_n26_), .B(ori_ori_n166_), .Y(ori_ori_n559_));
  INV        o537(.A(i_7_), .Y(ori_ori_n560_));
  INV        o538(.A(ori_ori_n558_), .Y(ori_ori_n561_));
  AOI220     o539(.A0(ori_ori_n308_), .A1(ori_ori_n504_), .B0(ori_ori_n87_), .B1(ori_ori_n96_), .Y(ori_ori_n562_));
  OAI220     o540(.A0(ori_ori_n562_), .A1(ori_ori_n456_), .B0(ori_ori_n561_), .B1(ori_ori_n467_), .Y(ori_ori_n563_));
  NO4        o541(.A(ori_ori_n563_), .B(ori_ori_n557_), .C(ori_ori_n553_), .D(ori_ori_n551_), .Y(ori_ori_n564_));
  OR2        o542(.A(i_11_), .B(i_6_), .Y(ori_ori_n565_));
  NA3        o543(.A(ori_ori_n455_), .B(ori_ori_n559_), .C(i_7_), .Y(ori_ori_n566_));
  AOI210     o544(.A0(ori_ori_n566_), .A1(ori_ori_n556_), .B0(ori_ori_n565_), .Y(ori_ori_n567_));
  NA3        o545(.A(ori_ori_n332_), .B(ori_ori_n459_), .C(ori_ori_n93_), .Y(ori_ori_n568_));
  NA2        o546(.A(ori_ori_n495_), .B(i_13_), .Y(ori_ori_n569_));
  NA2        o547(.A(ori_ori_n96_), .B(ori_ori_n559_), .Y(ori_ori_n570_));
  NAi21      o548(.An(i_11_), .B(i_12_), .Y(ori_ori_n571_));
  NOi41      o549(.An(ori_ori_n105_), .B(ori_ori_n571_), .C(i_13_), .D(ori_ori_n80_), .Y(ori_ori_n572_));
  NO3        o550(.A(ori_ori_n379_), .B(ori_ori_n438_), .C(ori_ori_n460_), .Y(ori_ori_n573_));
  AOI220     o551(.A0(ori_ori_n573_), .A1(ori_ori_n253_), .B0(ori_ori_n572_), .B1(ori_ori_n570_), .Y(ori_ori_n574_));
  NA3        o552(.A(ori_ori_n574_), .B(ori_ori_n569_), .C(ori_ori_n568_), .Y(ori_ori_n575_));
  OAI210     o553(.A0(ori_ori_n575_), .A1(ori_ori_n567_), .B0(ori_ori_n59_), .Y(ori_ori_n576_));
  NO2        o554(.A(i_2_), .B(i_12_), .Y(ori_ori_n577_));
  NA2        o555(.A(ori_ori_n290_), .B(ori_ori_n577_), .Y(ori_ori_n578_));
  INV        o556(.A(ori_ori_n578_), .Y(ori_ori_n579_));
  NA3        o557(.A(ori_ori_n579_), .B(ori_ori_n45_), .C(ori_ori_n192_), .Y(ori_ori_n580_));
  NA4        o558(.A(ori_ori_n580_), .B(ori_ori_n576_), .C(ori_ori_n564_), .D(ori_ori_n548_), .Y(ori_ori_n581_));
  OR4        o559(.A(ori_ori_n581_), .B(ori_ori_n541_), .C(ori_ori_n526_), .D(ori_ori_n469_), .Y(ori5));
  NA2        o560(.A(ori_ori_n515_), .B(ori_ori_n228_), .Y(ori_ori_n583_));
  AN2        o561(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n584_));
  NA3        o562(.A(ori_ori_n584_), .B(ori_ori_n577_), .C(ori_ori_n102_), .Y(ori_ori_n585_));
  NO2        o563(.A(ori_ori_n456_), .B(i_11_), .Y(ori_ori_n586_));
  NA2        o564(.A(ori_ori_n83_), .B(ori_ori_n586_), .Y(ori_ori_n587_));
  NA3        o565(.A(ori_ori_n587_), .B(ori_ori_n585_), .C(ori_ori_n583_), .Y(ori_ori_n588_));
  NO3        o566(.A(i_11_), .B(ori_ori_n199_), .C(i_13_), .Y(ori_ori_n589_));
  NO2        o567(.A(ori_ori_n119_), .B(ori_ori_n23_), .Y(ori_ori_n590_));
  NA2        o568(.A(i_12_), .B(i_8_), .Y(ori_ori_n591_));
  OAI210     o569(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n591_), .Y(ori_ori_n592_));
  INV        o570(.A(ori_ori_n348_), .Y(ori_ori_n593_));
  AOI220     o571(.A0(ori_ori_n255_), .A1(ori_ori_n433_), .B0(ori_ori_n592_), .B1(ori_ori_n590_), .Y(ori_ori_n594_));
  INV        o572(.A(ori_ori_n594_), .Y(ori_ori_n595_));
  NO2        o573(.A(ori_ori_n595_), .B(ori_ori_n588_), .Y(ori_ori_n596_));
  INV        o574(.A(ori_ori_n153_), .Y(ori_ori_n597_));
  INV        o575(.A(ori_ori_n206_), .Y(ori_ori_n598_));
  OAI210     o576(.A0(ori_ori_n537_), .A1(ori_ori_n350_), .B0(ori_ori_n105_), .Y(ori_ori_n599_));
  AOI210     o577(.A0(ori_ori_n599_), .A1(ori_ori_n598_), .B0(ori_ori_n597_), .Y(ori_ori_n600_));
  NO2        o578(.A(ori_ori_n358_), .B(ori_ori_n26_), .Y(ori_ori_n601_));
  NO2        o579(.A(ori_ori_n601_), .B(ori_ori_n335_), .Y(ori_ori_n602_));
  NA2        o580(.A(ori_ori_n602_), .B(i_2_), .Y(ori_ori_n603_));
  INV        o581(.A(ori_ori_n603_), .Y(ori_ori_n604_));
  AOI210     o582(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n333_), .Y(ori_ori_n605_));
  AOI210     o583(.A0(ori_ori_n605_), .A1(ori_ori_n604_), .B0(ori_ori_n600_), .Y(ori_ori_n606_));
  NO2        o584(.A(ori_ori_n165_), .B(ori_ori_n120_), .Y(ori_ori_n607_));
  OAI210     o585(.A0(ori_ori_n607_), .A1(ori_ori_n590_), .B0(i_2_), .Y(ori_ori_n608_));
  INV        o586(.A(ori_ori_n154_), .Y(ori_ori_n609_));
  NO3        o587(.A(ori_ori_n471_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n610_));
  AOI210     o588(.A0(ori_ori_n609_), .A1(ori_ori_n83_), .B0(ori_ori_n610_), .Y(ori_ori_n611_));
  AOI210     o589(.A0(ori_ori_n611_), .A1(ori_ori_n608_), .B0(ori_ori_n166_), .Y(ori_ori_n612_));
  OA210      o590(.A0(ori_ori_n472_), .A1(ori_ori_n121_), .B0(i_13_), .Y(ori_ori_n613_));
  AOI210     o591(.A0(ori_ori_n178_), .A1(ori_ori_n142_), .B0(ori_ori_n403_), .Y(ori_ori_n614_));
  NA2        o592(.A(ori_ori_n614_), .B(ori_ori_n335_), .Y(ori_ori_n615_));
  NO2        o593(.A(ori_ori_n96_), .B(ori_ori_n44_), .Y(ori_ori_n616_));
  INV        o594(.A(ori_ori_n247_), .Y(ori_ori_n617_));
  NA4        o595(.A(ori_ori_n617_), .B(ori_ori_n248_), .C(ori_ori_n119_), .D(ori_ori_n42_), .Y(ori_ori_n618_));
  OAI210     o596(.A0(ori_ori_n618_), .A1(ori_ori_n616_), .B0(ori_ori_n615_), .Y(ori_ori_n619_));
  NO3        o597(.A(ori_ori_n619_), .B(ori_ori_n613_), .C(ori_ori_n612_), .Y(ori_ori_n620_));
  NA2        o598(.A(ori_ori_n433_), .B(ori_ori_n28_), .Y(ori_ori_n621_));
  NA2        o599(.A(ori_ori_n589_), .B(ori_ori_n234_), .Y(ori_ori_n622_));
  NA2        o600(.A(ori_ori_n622_), .B(ori_ori_n621_), .Y(ori_ori_n623_));
  NO2        o601(.A(ori_ori_n58_), .B(i_12_), .Y(ori_ori_n624_));
  NO2        o602(.A(ori_ori_n624_), .B(ori_ori_n121_), .Y(ori_ori_n625_));
  NO2        o603(.A(ori_ori_n625_), .B(ori_ori_n452_), .Y(ori_ori_n626_));
  AOI220     o604(.A0(ori_ori_n626_), .A1(ori_ori_n36_), .B0(ori_ori_n623_), .B1(ori_ori_n46_), .Y(ori_ori_n627_));
  NA4        o605(.A(ori_ori_n627_), .B(ori_ori_n620_), .C(ori_ori_n606_), .D(ori_ori_n596_), .Y(ori6));
  NA4        o606(.A(ori_ori_n311_), .B(ori_ori_n380_), .C(ori_ori_n67_), .D(ori_ori_n95_), .Y(ori_ori_n629_));
  INV        o607(.A(ori_ori_n629_), .Y(ori_ori_n630_));
  NO2        o608(.A(ori_ori_n188_), .B(ori_ori_n383_), .Y(ori_ori_n631_));
  NO2        o609(.A(i_11_), .B(i_9_), .Y(ori_ori_n632_));
  NO2        o610(.A(ori_ori_n630_), .B(ori_ori_n259_), .Y(ori_ori_n633_));
  OR2        o611(.A(ori_ori_n633_), .B(i_12_), .Y(ori_ori_n634_));
  NA2        o612(.A(ori_ori_n296_), .B(ori_ori_n267_), .Y(ori_ori_n635_));
  NA2        o613(.A(ori_ori_n438_), .B(ori_ori_n59_), .Y(ori_ori_n636_));
  NA2        o614(.A(ori_ori_n528_), .B(ori_ori_n67_), .Y(ori_ori_n637_));
  BUFFER     o615(.A(ori_ori_n477_), .Y(ori_ori_n638_));
  NA4        o616(.A(ori_ori_n638_), .B(ori_ori_n637_), .C(ori_ori_n636_), .D(ori_ori_n635_), .Y(ori_ori_n639_));
  INV        o617(.A(ori_ori_n169_), .Y(ori_ori_n640_));
  AOI220     o618(.A0(ori_ori_n640_), .A1(ori_ori_n632_), .B0(ori_ori_n639_), .B1(ori_ori_n69_), .Y(ori_ori_n641_));
  INV        o619(.A(ori_ori_n258_), .Y(ori_ori_n642_));
  NA2        o620(.A(ori_ori_n71_), .B(ori_ori_n126_), .Y(ori_ori_n643_));
  INV        o621(.A(ori_ori_n119_), .Y(ori_ori_n644_));
  NA2        o622(.A(ori_ori_n644_), .B(ori_ori_n46_), .Y(ori_ori_n645_));
  AOI210     o623(.A0(ori_ori_n645_), .A1(ori_ori_n643_), .B0(ori_ori_n642_), .Y(ori_ori_n646_));
  NO2        o624(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n647_));
  NA3        o625(.A(ori_ori_n647_), .B(ori_ori_n376_), .C(ori_ori_n311_), .Y(ori_ori_n648_));
  NAi32      o626(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n649_));
  NO2        o627(.A(ori_ori_n565_), .B(ori_ori_n649_), .Y(ori_ori_n650_));
  OAI210     o628(.A0(ori_ori_n527_), .A1(ori_ori_n426_), .B0(ori_ori_n425_), .Y(ori_ori_n651_));
  NAi31      o629(.An(ori_ori_n650_), .B(ori_ori_n651_), .C(ori_ori_n648_), .Y(ori_ori_n652_));
  OR2        o630(.A(ori_ori_n652_), .B(ori_ori_n646_), .Y(ori_ori_n653_));
  AO220      o631(.A0(ori_ori_n279_), .A1(ori_ori_n270_), .B0(ori_ori_n319_), .B1(ori_ori_n452_), .Y(ori_ori_n654_));
  NA3        o632(.A(ori_ori_n654_), .B(ori_ori_n213_), .C(i_7_), .Y(ori_ori_n655_));
  BUFFER     o633(.A(ori_ori_n472_), .Y(ori_ori_n656_));
  NA3        o634(.A(ori_ori_n656_), .B(ori_ori_n141_), .C(ori_ori_n65_), .Y(ori_ori_n657_));
  AO210      o635(.A0(ori_ori_n390_), .A1(ori_ori_n593_), .B0(ori_ori_n36_), .Y(ori_ori_n658_));
  NA3        o636(.A(ori_ori_n658_), .B(ori_ori_n657_), .C(ori_ori_n655_), .Y(ori_ori_n659_));
  OAI210     o637(.A0(ori_ori_n494_), .A1(i_11_), .B0(ori_ori_n81_), .Y(ori_ori_n660_));
  AOI220     o638(.A0(ori_ori_n660_), .A1(ori_ori_n425_), .B0(ori_ori_n631_), .B1(ori_ori_n560_), .Y(ori_ori_n661_));
  NA3        o639(.A(ori_ori_n295_), .B(ori_ori_n201_), .C(ori_ori_n141_), .Y(ori_ori_n662_));
  NA2        o640(.A(ori_ori_n319_), .B(ori_ori_n66_), .Y(ori_ori_n663_));
  NA4        o641(.A(ori_ori_n663_), .B(ori_ori_n662_), .C(ori_ori_n661_), .D(ori_ori_n458_), .Y(ori_ori_n664_));
  AO210      o642(.A0(ori_ori_n403_), .A1(ori_ori_n46_), .B0(ori_ori_n82_), .Y(ori_ori_n665_));
  NA3        o643(.A(ori_ori_n665_), .B(ori_ori_n381_), .C(ori_ori_n186_), .Y(ori_ori_n666_));
  AOI210     o644(.A0(ori_ori_n350_), .A1(ori_ori_n348_), .B0(ori_ori_n424_), .Y(ori_ori_n667_));
  NO2        o645(.A(ori_ori_n466_), .B(ori_ori_n96_), .Y(ori_ori_n668_));
  OAI210     o646(.A0(ori_ori_n668_), .A1(ori_ori_n106_), .B0(ori_ori_n331_), .Y(ori_ori_n669_));
  NA2        o647(.A(ori_ori_n205_), .B(ori_ori_n46_), .Y(ori_ori_n670_));
  NA3        o648(.A(ori_ori_n669_), .B(ori_ori_n667_), .C(ori_ori_n666_), .Y(ori_ori_n671_));
  NO4        o649(.A(ori_ori_n671_), .B(ori_ori_n664_), .C(ori_ori_n659_), .D(ori_ori_n653_), .Y(ori_ori_n672_));
  NA4        o650(.A(ori_ori_n672_), .B(ori_ori_n641_), .C(ori_ori_n634_), .D(ori_ori_n303_), .Y(ori3));
  NA2        o651(.A(i_12_), .B(i_10_), .Y(ori_ori_n674_));
  NO2        o652(.A(i_11_), .B(ori_ori_n199_), .Y(ori_ori_n675_));
  NA3        o653(.A(ori_ori_n662_), .B(ori_ori_n458_), .C(ori_ori_n294_), .Y(ori_ori_n676_));
  NA2        o654(.A(ori_ori_n676_), .B(ori_ori_n40_), .Y(ori_ori_n677_));
  NOi21      o655(.An(ori_ori_n92_), .B(ori_ori_n602_), .Y(ori_ori_n678_));
  NO3        o656(.A(ori_ori_n482_), .B(ori_ori_n358_), .C(ori_ori_n126_), .Y(ori_ori_n679_));
  NA2        o657(.A(ori_ori_n332_), .B(ori_ori_n45_), .Y(ori_ori_n680_));
  NO2        o658(.A(ori_ori_n679_), .B(ori_ori_n678_), .Y(ori_ori_n681_));
  AOI210     o659(.A0(ori_ori_n681_), .A1(ori_ori_n677_), .B0(ori_ori_n48_), .Y(ori_ori_n682_));
  NO4        o660(.A(ori_ori_n299_), .B(ori_ori_n306_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n683_));
  NA2        o661(.A(ori_ori_n160_), .B(ori_ori_n429_), .Y(ori_ori_n684_));
  NOi21      o662(.An(ori_ori_n684_), .B(ori_ori_n683_), .Y(ori_ori_n685_));
  NO2        o663(.A(ori_ori_n685_), .B(ori_ori_n59_), .Y(ori_ori_n686_));
  NOi21      o664(.An(i_5_), .B(i_9_), .Y(ori_ori_n687_));
  NA2        o665(.A(ori_ori_n687_), .B(ori_ori_n347_), .Y(ori_ori_n688_));
  BUFFER     o666(.A(ori_ori_n225_), .Y(ori_ori_n689_));
  AOI210     o667(.A0(ori_ori_n689_), .A1(ori_ori_n377_), .B0(ori_ori_n531_), .Y(ori_ori_n690_));
  NO2        o668(.A(ori_ori_n690_), .B(ori_ori_n688_), .Y(ori_ori_n691_));
  NO3        o669(.A(ori_ori_n691_), .B(ori_ori_n686_), .C(ori_ori_n682_), .Y(ori_ori_n692_));
  NA2        o670(.A(ori_ori_n160_), .B(ori_ori_n24_), .Y(ori_ori_n693_));
  NO2        o671(.A(ori_ori_n518_), .B(ori_ori_n449_), .Y(ori_ori_n694_));
  NO2        o672(.A(ori_ori_n694_), .B(ori_ori_n693_), .Y(ori_ori_n695_));
  NA2        o673(.A(ori_ori_n253_), .B(ori_ori_n124_), .Y(ori_ori_n696_));
  NAi21      o674(.An(ori_ori_n149_), .B(ori_ori_n340_), .Y(ori_ori_n697_));
  OAI220     o675(.A0(ori_ori_n697_), .A1(ori_ori_n670_), .B0(ori_ori_n696_), .B1(ori_ori_n324_), .Y(ori_ori_n698_));
  NO2        o676(.A(ori_ori_n698_), .B(ori_ori_n695_), .Y(ori_ori_n699_));
  NA2        o677(.A(ori_ori_n430_), .B(i_0_), .Y(ori_ori_n700_));
  NO3        o678(.A(ori_ori_n700_), .B(ori_ori_n307_), .C(ori_ori_n83_), .Y(ori_ori_n701_));
  INV        o679(.A(ori_ori_n701_), .Y(ori_ori_n702_));
  NA2        o680(.A(ori_ori_n589_), .B(ori_ori_n259_), .Y(ori_ori_n703_));
  AOI210     o681(.A0(ori_ori_n381_), .A1(ori_ori_n83_), .B0(ori_ori_n56_), .Y(ori_ori_n704_));
  NO2        o682(.A(ori_ori_n704_), .B(ori_ori_n703_), .Y(ori_ori_n705_));
  NA2        o683(.A(i_0_), .B(i_10_), .Y(ori_ori_n706_));
  INV        o684(.A(ori_ori_n705_), .Y(ori_ori_n707_));
  NA3        o685(.A(ori_ori_n707_), .B(ori_ori_n702_), .C(ori_ori_n699_), .Y(ori_ori_n708_));
  NO2        o686(.A(ori_ori_n97_), .B(ori_ori_n37_), .Y(ori_ori_n709_));
  NA2        o687(.A(i_11_), .B(i_9_), .Y(ori_ori_n710_));
  NO3        o688(.A(i_12_), .B(ori_ori_n710_), .C(ori_ori_n457_), .Y(ori_ori_n711_));
  AN2        o689(.A(ori_ori_n711_), .B(ori_ori_n709_), .Y(ori_ori_n712_));
  NA2        o690(.A(ori_ori_n316_), .B(ori_ori_n158_), .Y(ori_ori_n713_));
  INV        o691(.A(ori_ori_n713_), .Y(ori_ori_n714_));
  NO2        o692(.A(ori_ori_n710_), .B(ori_ori_n69_), .Y(ori_ori_n715_));
  NO2        o693(.A(ori_ori_n156_), .B(i_0_), .Y(ori_ori_n716_));
  INV        o694(.A(ori_ori_n330_), .Y(ori_ori_n717_));
  NO2        o695(.A(ori_ori_n717_), .B(ori_ori_n688_), .Y(ori_ori_n718_));
  NO3        o696(.A(ori_ori_n718_), .B(ori_ori_n714_), .C(ori_ori_n712_), .Y(ori_ori_n719_));
  NA2        o697(.A(ori_ori_n511_), .B(ori_ori_n116_), .Y(ori_ori_n720_));
  NO2        o698(.A(i_6_), .B(ori_ori_n720_), .Y(ori_ori_n721_));
  NA2        o699(.A(ori_ori_n153_), .B(ori_ori_n97_), .Y(ori_ori_n722_));
  NA2        o700(.A(ori_ori_n459_), .B(ori_ori_n259_), .Y(ori_ori_n723_));
  NO2        o701(.A(ori_ori_n723_), .B(ori_ori_n680_), .Y(ori_ori_n724_));
  NO2        o702(.A(ori_ori_n724_), .B(ori_ori_n721_), .Y(ori_ori_n725_));
  NOi21      o703(.An(i_7_), .B(i_5_), .Y(ori_ori_n726_));
  NOi31      o704(.An(ori_ori_n726_), .B(i_0_), .C(ori_ori_n571_), .Y(ori_ori_n727_));
  NA3        o705(.A(ori_ori_n727_), .B(ori_ori_n829_), .C(i_6_), .Y(ori_ori_n728_));
  BUFFER     o706(.A(ori_ori_n728_), .Y(ori_ori_n729_));
  INV        o707(.A(ori_ori_n256_), .Y(ori_ori_n730_));
  NA3        o708(.A(ori_ori_n729_), .B(ori_ori_n725_), .C(ori_ori_n719_), .Y(ori_ori_n731_));
  NO2        o709(.A(ori_ori_n674_), .B(ori_ori_n255_), .Y(ori_ori_n732_));
  OA210      o710(.A0(ori_ori_n376_), .A1(ori_ori_n190_), .B0(ori_ori_n375_), .Y(ori_ori_n733_));
  NA2        o711(.A(ori_ori_n732_), .B(ori_ori_n715_), .Y(ori_ori_n734_));
  NA3        o712(.A(ori_ori_n375_), .B(ori_ori_n332_), .C(ori_ori_n45_), .Y(ori_ori_n735_));
  OAI210     o713(.A0(ori_ori_n697_), .A1(i_7_), .B0(ori_ori_n735_), .Y(ori_ori_n736_));
  NA2        o714(.A(ori_ori_n715_), .B(ori_ori_n248_), .Y(ori_ori_n737_));
  OAI210     o715(.A0(i_3_), .A1(ori_ori_n162_), .B0(ori_ori_n737_), .Y(ori_ori_n738_));
  AOI220     o716(.A0(ori_ori_n738_), .A1(ori_ori_n376_), .B0(ori_ori_n736_), .B1(ori_ori_n69_), .Y(ori_ori_n739_));
  NA3        o717(.A(i_5_), .B(ori_ori_n305_), .C(ori_ori_n494_), .Y(ori_ori_n740_));
  NA2        o718(.A(ori_ori_n88_), .B(ori_ori_n44_), .Y(ori_ori_n741_));
  NO2        o719(.A(ori_ori_n71_), .B(ori_ori_n591_), .Y(ori_ori_n742_));
  AOI220     o720(.A0(ori_ori_n742_), .A1(ori_ori_n741_), .B0(ori_ori_n155_), .B1(ori_ori_n449_), .Y(ori_ori_n743_));
  AOI210     o721(.A0(ori_ori_n743_), .A1(ori_ori_n740_), .B0(ori_ori_n47_), .Y(ori_ori_n744_));
  NO3        o722(.A(i_5_), .B(ori_ori_n277_), .C(ori_ori_n24_), .Y(ori_ori_n745_));
  AOI210     o723(.A0(ori_ori_n546_), .A1(ori_ori_n414_), .B0(ori_ori_n745_), .Y(ori_ori_n746_));
  NAi21      o724(.An(i_9_), .B(i_5_), .Y(ori_ori_n747_));
  NO2        o725(.A(ori_ori_n747_), .B(ori_ori_n325_), .Y(ori_ori_n748_));
  NA2        o726(.A(ori_ori_n748_), .B(ori_ori_n472_), .Y(ori_ori_n749_));
  OAI220     o727(.A0(ori_ori_n749_), .A1(ori_ori_n80_), .B0(ori_ori_n746_), .B1(ori_ori_n154_), .Y(ori_ori_n750_));
  NO2        o728(.A(ori_ori_n750_), .B(ori_ori_n744_), .Y(ori_ori_n751_));
  NA3        o729(.A(ori_ori_n751_), .B(ori_ori_n739_), .C(ori_ori_n734_), .Y(ori_ori_n752_));
  NO3        o730(.A(ori_ori_n752_), .B(ori_ori_n731_), .C(ori_ori_n708_), .Y(ori_ori_n753_));
  NO2        o731(.A(i_0_), .B(ori_ori_n571_), .Y(ori_ori_n754_));
  NO2        o732(.A(ori_ori_n636_), .B(ori_ori_n722_), .Y(ori_ori_n755_));
  INV        o733(.A(ori_ori_n755_), .Y(ori_ori_n756_));
  NO2        o734(.A(ori_ori_n651_), .B(ori_ori_n325_), .Y(ori_ori_n757_));
  NA2        o735(.A(ori_ori_n205_), .B(ori_ori_n197_), .Y(ori_ori_n758_));
  AOI210     o736(.A0(ori_ori_n758_), .A1(ori_ori_n700_), .B0(ori_ori_n145_), .Y(ori_ori_n759_));
  NO2        o737(.A(ori_ori_n759_), .B(ori_ori_n757_), .Y(ori_ori_n760_));
  NA2        o738(.A(ori_ori_n760_), .B(ori_ori_n756_), .Y(ori_ori_n761_));
  NO3        o739(.A(ori_ori_n706_), .B(ori_ori_n687_), .C(ori_ori_n165_), .Y(ori_ori_n762_));
  AOI220     o740(.A0(ori_ori_n762_), .A1(i_11_), .B0(ori_ori_n428_), .B1(ori_ori_n71_), .Y(ori_ori_n763_));
  NO3        o741(.A(ori_ori_n179_), .B(ori_ori_n306_), .C(i_0_), .Y(ori_ori_n764_));
  OAI210     o742(.A0(ori_ori_n764_), .A1(ori_ori_n72_), .B0(i_13_), .Y(ori_ori_n765_));
  NA2        o743(.A(ori_ori_n765_), .B(ori_ori_n763_), .Y(ori_ori_n766_));
  NO2        o744(.A(ori_ori_n204_), .B(ori_ori_n88_), .Y(ori_ori_n767_));
  AOI210     o745(.A0(ori_ori_n767_), .A1(ori_ori_n754_), .B0(ori_ori_n103_), .Y(ori_ori_n768_));
  OR2        o746(.A(ori_ori_n768_), .B(i_5_), .Y(ori_ori_n769_));
  AOI210     o747(.A0(i_0_), .A1(ori_ori_n25_), .B0(ori_ori_n156_), .Y(ori_ori_n770_));
  NA2        o748(.A(ori_ori_n770_), .B(ori_ori_n733_), .Y(ori_ori_n771_));
  NO3        o749(.A(ori_ori_n680_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n772_));
  NA2        o750(.A(ori_ori_n389_), .B(ori_ori_n382_), .Y(ori_ori_n773_));
  NO2        o751(.A(ori_ori_n773_), .B(ori_ori_n772_), .Y(ori_ori_n774_));
  NA3        o752(.A(ori_ori_n311_), .B(ori_ori_n153_), .C(ori_ori_n152_), .Y(ori_ori_n775_));
  NA3        o753(.A(i_5_), .B(ori_ori_n240_), .C(ori_ori_n197_), .Y(ori_ori_n776_));
  NA2        o754(.A(ori_ori_n776_), .B(ori_ori_n775_), .Y(ori_ori_n777_));
  NA3        o755(.A(ori_ori_n311_), .B(ori_ori_n266_), .C(ori_ori_n189_), .Y(ori_ori_n778_));
  INV        o756(.A(ori_ori_n778_), .Y(ori_ori_n779_));
  NO3        o757(.A(ori_ori_n710_), .B(ori_ori_n186_), .C(ori_ori_n165_), .Y(ori_ori_n780_));
  NO3        o758(.A(ori_ori_n780_), .B(ori_ori_n779_), .C(ori_ori_n777_), .Y(ori_ori_n781_));
  NA4        o759(.A(ori_ori_n781_), .B(ori_ori_n774_), .C(ori_ori_n771_), .D(ori_ori_n769_), .Y(ori_ori_n782_));
  NO2        o760(.A(ori_ori_n80_), .B(i_5_), .Y(ori_ori_n783_));
  NA3        o761(.A(ori_ori_n675_), .B(ori_ori_n104_), .C(ori_ori_n119_), .Y(ori_ori_n784_));
  INV        o762(.A(ori_ori_n784_), .Y(ori_ori_n785_));
  NA2        o763(.A(ori_ori_n785_), .B(ori_ori_n783_), .Y(ori_ori_n786_));
  NA3        o764(.A(ori_ori_n248_), .B(i_5_), .C(ori_ori_n166_), .Y(ori_ori_n787_));
  NAi31      o765(.An(ori_ori_n203_), .B(ori_ori_n787_), .C(ori_ori_n204_), .Y(ori_ori_n788_));
  NO4        o766(.A(ori_ori_n202_), .B(ori_ori_n179_), .C(i_0_), .D(i_12_), .Y(ori_ori_n789_));
  AOI220     o767(.A0(ori_ori_n789_), .A1(ori_ori_n788_), .B0(ori_ori_n630_), .B1(ori_ori_n157_), .Y(ori_ori_n790_));
  AN2        o768(.A(ori_ori_n706_), .B(ori_ori_n145_), .Y(ori_ori_n791_));
  NO4        o769(.A(ori_ori_n791_), .B(i_12_), .C(ori_ori_n500_), .D(ori_ori_n126_), .Y(ori_ori_n792_));
  NA2        o770(.A(ori_ori_n792_), .B(ori_ori_n186_), .Y(ori_ori_n793_));
  NA2        o771(.A(ori_ori_n726_), .B(ori_ori_n373_), .Y(ori_ori_n794_));
  NA2        o772(.A(ori_ori_n60_), .B(ori_ori_n95_), .Y(ori_ori_n795_));
  OAI220     o773(.A0(ori_ori_n795_), .A1(ori_ori_n787_), .B0(ori_ori_n794_), .B1(ori_ori_n521_), .Y(ori_ori_n796_));
  NA2        o774(.A(ori_ori_n796_), .B(ori_ori_n716_), .Y(ori_ori_n797_));
  NA4        o775(.A(ori_ori_n797_), .B(ori_ori_n793_), .C(ori_ori_n790_), .D(ori_ori_n786_), .Y(ori_ori_n798_));
  NO4        o776(.A(ori_ori_n798_), .B(ori_ori_n782_), .C(ori_ori_n766_), .D(ori_ori_n761_), .Y(ori_ori_n799_));
  NA2        o777(.A(ori_ori_n647_), .B(ori_ori_n37_), .Y(ori_ori_n800_));
  NA2        o778(.A(ori_ori_n800_), .B(ori_ori_n465_), .Y(ori_ori_n801_));
  NA2        o779(.A(ori_ori_n801_), .B(ori_ori_n177_), .Y(ori_ori_n802_));
  NA2        o780(.A(ori_ori_n497_), .B(ori_ori_n48_), .Y(ori_ori_n803_));
  AOI210     o781(.A0(ori_ori_n803_), .A1(ori_ori_n802_), .B0(ori_ori_n69_), .Y(ori_ori_n804_));
  INV        o782(.A(ori_ori_n302_), .Y(ori_ori_n805_));
  NO2        o783(.A(ori_ori_n805_), .B(ori_ori_n597_), .Y(ori_ori_n806_));
  INV        o784(.A(ori_ori_n72_), .Y(ori_ori_n807_));
  AOI210     o785(.A0(ori_ori_n770_), .A1(i_5_), .B0(ori_ori_n727_), .Y(ori_ori_n808_));
  AOI210     o786(.A0(ori_ori_n808_), .A1(ori_ori_n807_), .B0(ori_ori_n524_), .Y(ori_ori_n809_));
  INV        o787(.A(ori_ori_n809_), .Y(ori_ori_n810_));
  NA2        o788(.A(ori_ori_n227_), .B(ori_ori_n83_), .Y(ori_ori_n811_));
  NA3        o789(.A(ori_ori_n601_), .B(ori_ori_n240_), .C(ori_ori_n76_), .Y(ori_ori_n812_));
  AOI210     o790(.A0(ori_ori_n812_), .A1(ori_ori_n811_), .B0(i_11_), .Y(ori_ori_n813_));
  NO3        o791(.A(ori_ori_n57_), .B(ori_ori_n56_), .C(i_4_), .Y(ori_ori_n814_));
  OAI210     o792(.A0(ori_ori_n730_), .A1(ori_ori_n249_), .B0(ori_ori_n814_), .Y(ori_ori_n815_));
  NO2        o793(.A(ori_ori_n815_), .B(ori_ori_n571_), .Y(ori_ori_n816_));
  NO4        o794(.A(ori_ori_n747_), .B(ori_ori_n378_), .C(ori_ori_n210_), .D(ori_ori_n209_), .Y(ori_ori_n817_));
  NO2        o795(.A(ori_ori_n817_), .B(ori_ori_n424_), .Y(ori_ori_n818_));
  INV        o796(.A(ori_ori_n283_), .Y(ori_ori_n819_));
  AOI210     o797(.A0(ori_ori_n819_), .A1(ori_ori_n818_), .B0(ori_ori_n41_), .Y(ori_ori_n820_));
  NO3        o798(.A(ori_ori_n820_), .B(ori_ori_n816_), .C(ori_ori_n813_), .Y(ori_ori_n821_));
  OAI210     o799(.A0(ori_ori_n810_), .A1(i_4_), .B0(ori_ori_n821_), .Y(ori_ori_n822_));
  NO3        o800(.A(ori_ori_n822_), .B(ori_ori_n806_), .C(ori_ori_n804_), .Y(ori_ori_n823_));
  NA4        o801(.A(ori_ori_n823_), .B(ori_ori_n799_), .C(ori_ori_n753_), .D(ori_ori_n692_), .Y(ori4));
  INV        o802(.A(ori_ori_n545_), .Y(ori_ori_n827_));
  INV        o803(.A(i_6_), .Y(ori_ori_n828_));
  INV        o804(.A(i_4_), .Y(ori_ori_n829_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m021(.A(mai_mai_n35_), .Y(mai1));
  INV        m022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m024(.A(i_2_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NO2        m026(.A(i_7_), .B(i_10_), .Y(mai_mai_n49_));
  AOI210     m027(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n49_), .Y(mai_mai_n50_));
  NA2        m028(.A(i_0_), .B(i_2_), .Y(mai_mai_n51_));
  NA2        m029(.A(i_7_), .B(i_9_), .Y(mai_mai_n52_));
  NO2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NA3        m031(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n54_));
  NO2        m032(.A(i_1_), .B(i_6_), .Y(mai_mai_n55_));
  NA2        m033(.A(i_8_), .B(i_7_), .Y(mai_mai_n56_));
  OAI210     m034(.A0(mai_mai_n56_), .A1(mai_mai_n55_), .B0(mai_mai_n54_), .Y(mai_mai_n57_));
  NA2        m035(.A(mai_mai_n57_), .B(i_12_), .Y(mai_mai_n58_));
  NAi21      m036(.An(i_2_), .B(i_7_), .Y(mai_mai_n59_));
  INV        m037(.A(i_1_), .Y(mai_mai_n60_));
  NA2        m038(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n61_));
  NA3        m039(.A(mai_mai_n61_), .B(mai_mai_n59_), .C(mai_mai_n31_), .Y(mai_mai_n62_));
  NA2        m040(.A(i_1_), .B(i_10_), .Y(mai_mai_n63_));
  NO2        m041(.A(mai_mai_n63_), .B(i_6_), .Y(mai_mai_n64_));
  NAi31      m042(.An(mai_mai_n64_), .B(mai_mai_n62_), .C(mai_mai_n58_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n50_), .B(i_2_), .Y(mai_mai_n66_));
  AOI210     m044(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n67_));
  NA2        m045(.A(i_1_), .B(i_6_), .Y(mai_mai_n68_));
  NO2        m046(.A(mai_mai_n68_), .B(mai_mai_n25_), .Y(mai_mai_n69_));
  INV        m047(.A(i_0_), .Y(mai_mai_n70_));
  NAi21      m048(.An(i_5_), .B(i_10_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_5_), .B(i_9_), .Y(mai_mai_n72_));
  AOI210     m050(.A0(mai_mai_n72_), .A1(mai_mai_n71_), .B0(mai_mai_n70_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n69_), .Y(mai_mai_n74_));
  OAI210     m052(.A0(mai_mai_n67_), .A1(mai_mai_n66_), .B0(mai_mai_n74_), .Y(mai_mai_n75_));
  OAI210     m053(.A0(mai_mai_n75_), .A1(mai_mai_n65_), .B0(i_0_), .Y(mai_mai_n76_));
  NA2        m054(.A(i_12_), .B(i_5_), .Y(mai_mai_n77_));
  NA2        m055(.A(i_2_), .B(i_8_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n78_), .B(mai_mai_n55_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_3_), .B(i_9_), .Y(mai_mai_n80_));
  NO2        m058(.A(i_3_), .B(i_7_), .Y(mai_mai_n81_));
  NO2        m059(.A(mai_mai_n80_), .B(mai_mai_n60_), .Y(mai_mai_n82_));
  INV        m060(.A(i_6_), .Y(mai_mai_n83_));
  OR4        m061(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n84_));
  INV        m062(.A(mai_mai_n84_), .Y(mai_mai_n85_));
  NO2        m063(.A(i_2_), .B(i_7_), .Y(mai_mai_n86_));
  NO2        m064(.A(mai_mai_n85_), .B(mai_mai_n86_), .Y(mai_mai_n87_));
  OAI210     m065(.A0(mai_mai_n82_), .A1(mai_mai_n79_), .B0(mai_mai_n87_), .Y(mai_mai_n88_));
  NAi21      m066(.An(i_6_), .B(i_10_), .Y(mai_mai_n89_));
  NA2        m067(.A(i_6_), .B(i_9_), .Y(mai_mai_n90_));
  AOI210     m068(.A0(mai_mai_n90_), .A1(mai_mai_n89_), .B0(mai_mai_n60_), .Y(mai_mai_n91_));
  NA2        m069(.A(i_2_), .B(i_6_), .Y(mai_mai_n92_));
  INV        m070(.A(mai_mai_n91_), .Y(mai_mai_n93_));
  AOI210     m071(.A0(mai_mai_n93_), .A1(mai_mai_n88_), .B0(mai_mai_n77_), .Y(mai_mai_n94_));
  AN3        m072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n95_));
  NAi21      m073(.An(i_6_), .B(i_11_), .Y(mai_mai_n96_));
  NO2        m074(.A(i_5_), .B(i_8_), .Y(mai_mai_n97_));
  NOi21      m075(.An(mai_mai_n97_), .B(mai_mai_n96_), .Y(mai_mai_n98_));
  AOI220     m076(.A0(mai_mai_n98_), .A1(mai_mai_n59_), .B0(mai_mai_n95_), .B1(mai_mai_n32_), .Y(mai_mai_n99_));
  INV        m077(.A(i_7_), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n47_), .B(mai_mai_n100_), .Y(mai_mai_n101_));
  NO2        m079(.A(i_0_), .B(i_5_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(mai_mai_n83_), .Y(mai_mai_n103_));
  NA2        m081(.A(i_12_), .B(i_3_), .Y(mai_mai_n104_));
  INV        m082(.A(mai_mai_n104_), .Y(mai_mai_n105_));
  NA3        m083(.A(mai_mai_n105_), .B(mai_mai_n103_), .C(mai_mai_n101_), .Y(mai_mai_n106_));
  NAi21      m084(.An(i_7_), .B(i_11_), .Y(mai_mai_n107_));
  NO3        m085(.A(mai_mai_n107_), .B(mai_mai_n89_), .C(mai_mai_n51_), .Y(mai_mai_n108_));
  AN2        m086(.A(i_2_), .B(i_10_), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(i_7_), .Y(mai_mai_n110_));
  OR2        m088(.A(mai_mai_n77_), .B(mai_mai_n55_), .Y(mai_mai_n111_));
  NO2        m089(.A(i_8_), .B(mai_mai_n100_), .Y(mai_mai_n112_));
  NA2        m090(.A(i_12_), .B(i_7_), .Y(mai_mai_n113_));
  NA2        m091(.A(i_11_), .B(i_12_), .Y(mai_mai_n114_));
  NAi41      m092(.An(mai_mai_n108_), .B(mai_mai_n114_), .C(mai_mai_n106_), .D(mai_mai_n99_), .Y(mai_mai_n115_));
  NOi21      m093(.An(i_1_), .B(i_5_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(i_11_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n100_), .B(mai_mai_n37_), .Y(mai_mai_n118_));
  NA2        m096(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n118_), .Y(mai_mai_n120_));
  NO2        m098(.A(mai_mai_n120_), .B(mai_mai_n47_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n122_));
  NAi21      m100(.An(i_3_), .B(i_8_), .Y(mai_mai_n123_));
  NA2        m101(.A(mai_mai_n123_), .B(mai_mai_n59_), .Y(mai_mai_n124_));
  NOi31      m102(.An(mai_mai_n124_), .B(mai_mai_n122_), .C(mai_mai_n121_), .Y(mai_mai_n125_));
  NO2        m103(.A(i_1_), .B(mai_mai_n83_), .Y(mai_mai_n126_));
  NO2        m104(.A(i_6_), .B(i_5_), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n127_), .B(i_3_), .Y(mai_mai_n128_));
  OAI220     m106(.A0(mai_mai_n128_), .A1(mai_mai_n107_), .B0(mai_mai_n125_), .B1(mai_mai_n117_), .Y(mai_mai_n129_));
  NO3        m107(.A(mai_mai_n129_), .B(mai_mai_n115_), .C(mai_mai_n94_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n76_), .Y(mai2));
  NO2        m109(.A(mai_mai_n60_), .B(mai_mai_n37_), .Y(mai_mai_n132_));
  NA2        m110(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n133_), .B(mai_mai_n132_), .Y(mai_mai_n134_));
  NA4        m112(.A(mai_mai_n134_), .B(mai_mai_n74_), .C(mai_mai_n66_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m113(.A(i_8_), .B(i_7_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n136_), .B(i_6_), .Y(mai_mai_n137_));
  NO2        m115(.A(i_12_), .B(i_13_), .Y(mai_mai_n138_));
  NAi21      m116(.An(i_5_), .B(i_11_), .Y(mai_mai_n139_));
  NOi21      m117(.An(mai_mai_n138_), .B(mai_mai_n139_), .Y(mai_mai_n140_));
  NO2        m118(.A(i_0_), .B(i_1_), .Y(mai_mai_n141_));
  NA2        m119(.A(i_2_), .B(i_3_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n142_), .B(i_4_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(mai_mai_n140_), .Y(mai_mai_n144_));
  AN2        m122(.A(mai_mai_n138_), .B(mai_mai_n80_), .Y(mai_mai_n145_));
  NO2        m123(.A(mai_mai_n145_), .B(mai_mai_n27_), .Y(mai_mai_n146_));
  NA2        m124(.A(i_1_), .B(i_5_), .Y(mai_mai_n147_));
  NO2        m125(.A(mai_mai_n70_), .B(mai_mai_n47_), .Y(mai_mai_n148_));
  NA2        m126(.A(mai_mai_n148_), .B(mai_mai_n36_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n147_), .C(mai_mai_n146_), .Y(mai_mai_n150_));
  OR2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NO3        m129(.A(mai_mai_n151_), .B(mai_mai_n77_), .C(i_13_), .Y(mai_mai_n152_));
  NAi32      m130(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n153_));
  NAi21      m131(.An(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  NOi21      m132(.An(i_4_), .B(i_10_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n155_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NO2        m134(.A(i_3_), .B(i_5_), .Y(mai_mai_n157_));
  NO3        m135(.A(mai_mai_n70_), .B(i_2_), .C(i_1_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  OAI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n156_), .B0(mai_mai_n154_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n160_), .B(mai_mai_n150_), .Y(mai_mai_n161_));
  AOI210     m139(.A0(mai_mai_n161_), .A1(mai_mai_n144_), .B0(mai_mai_n137_), .Y(mai_mai_n162_));
  NA3        m140(.A(mai_mai_n70_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n163_));
  NA2        m141(.A(i_3_), .B(mai_mai_n48_), .Y(mai_mai_n164_));
  NOi21      m142(.An(i_4_), .B(i_9_), .Y(mai_mai_n165_));
  NOi21      m143(.An(i_11_), .B(i_13_), .Y(mai_mai_n166_));
  NA2        m144(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  NO2        m145(.A(i_4_), .B(i_5_), .Y(mai_mai_n168_));
  NAi21      m146(.An(i_12_), .B(i_11_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(i_13_), .Y(mai_mai_n170_));
  NA3        m148(.A(mai_mai_n170_), .B(mai_mai_n168_), .C(mai_mai_n80_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n167_), .B0(mai_mai_n163_), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n70_), .B(mai_mai_n60_), .Y(mai_mai_n173_));
  INV        m151(.A(mai_mai_n173_), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n175_));
  NAi31      m153(.An(mai_mai_n175_), .B(mai_mai_n145_), .C(i_11_), .Y(mai_mai_n176_));
  NA2        m154(.A(i_3_), .B(i_5_), .Y(mai_mai_n177_));
  OR2        m155(.A(mai_mai_n177_), .B(mai_mai_n167_), .Y(mai_mai_n178_));
  AOI210     m156(.A0(mai_mai_n178_), .A1(mai_mai_n176_), .B0(mai_mai_n174_), .Y(mai_mai_n179_));
  NO2        m157(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n180_));
  NO2        m158(.A(i_13_), .B(i_10_), .Y(mai_mai_n181_));
  NA3        m159(.A(mai_mai_n181_), .B(mai_mai_n180_), .C(mai_mai_n45_), .Y(mai_mai_n182_));
  NO2        m160(.A(i_2_), .B(i_1_), .Y(mai_mai_n183_));
  NA2        m161(.A(mai_mai_n183_), .B(i_3_), .Y(mai_mai_n184_));
  NAi21      m162(.An(i_4_), .B(i_12_), .Y(mai_mai_n185_));
  NO3        m163(.A(mai_mai_n184_), .B(mai_mai_n182_), .C(mai_mai_n25_), .Y(mai_mai_n186_));
  NO3        m164(.A(mai_mai_n186_), .B(mai_mai_n179_), .C(mai_mai_n172_), .Y(mai_mai_n187_));
  INV        m165(.A(i_8_), .Y(mai_mai_n188_));
  NO2        m166(.A(mai_mai_n188_), .B(i_7_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n189_), .B(i_6_), .Y(mai_mai_n190_));
  NO3        m168(.A(i_3_), .B(mai_mai_n83_), .C(mai_mai_n48_), .Y(mai_mai_n191_));
  NA2        m169(.A(mai_mai_n191_), .B(mai_mai_n112_), .Y(mai_mai_n192_));
  NO3        m170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n193_));
  NA3        m171(.A(mai_mai_n193_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n194_));
  NO3        m172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n195_));
  OAI210     m173(.A0(mai_mai_n95_), .A1(i_12_), .B0(mai_mai_n195_), .Y(mai_mai_n196_));
  AOI210     m174(.A0(mai_mai_n196_), .A1(mai_mai_n194_), .B0(mai_mai_n192_), .Y(mai_mai_n197_));
  NO2        m175(.A(i_3_), .B(i_8_), .Y(mai_mai_n198_));
  NO3        m176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n102_), .B(mai_mai_n55_), .Y(mai_mai_n200_));
  NO2        m178(.A(i_13_), .B(i_9_), .Y(mai_mai_n201_));
  NA3        m179(.A(mai_mai_n201_), .B(i_6_), .C(mai_mai_n188_), .Y(mai_mai_n202_));
  NAi21      m180(.An(i_12_), .B(i_3_), .Y(mai_mai_n203_));
  OR2        m181(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n205_));
  NO3        m183(.A(i_0_), .B(i_2_), .C(mai_mai_n60_), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n206_), .B(mai_mai_n205_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n207_), .B(mai_mai_n204_), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n208_), .B(mai_mai_n197_), .Y(mai_mai_n209_));
  OAI220     m187(.A0(mai_mai_n209_), .A1(i_4_), .B0(mai_mai_n190_), .B1(mai_mai_n187_), .Y(mai_mai_n210_));
  NAi21      m188(.An(i_12_), .B(i_7_), .Y(mai_mai_n211_));
  NA3        m189(.A(i_13_), .B(mai_mai_n188_), .C(i_10_), .Y(mai_mai_n212_));
  NA2        m190(.A(i_0_), .B(i_5_), .Y(mai_mai_n213_));
  NAi31      m191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n70_), .B(mai_mai_n26_), .Y(mai_mai_n216_));
  NO2        m194(.A(mai_mai_n47_), .B(mai_mai_n60_), .Y(mai_mai_n217_));
  INV        m195(.A(i_13_), .Y(mai_mai_n218_));
  NO2        m196(.A(i_12_), .B(mai_mai_n218_), .Y(mai_mai_n219_));
  NO2        m197(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n220_));
  NO2        m198(.A(mai_mai_n177_), .B(i_4_), .Y(mai_mai_n221_));
  NA2        m199(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  OR2        m200(.A(i_8_), .B(i_7_), .Y(mai_mai_n223_));
  NO2        m201(.A(mai_mai_n223_), .B(mai_mai_n83_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n51_), .B(i_1_), .Y(mai_mai_n225_));
  NA2        m203(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n226_));
  INV        m204(.A(i_12_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n45_), .B(mai_mai_n227_), .Y(mai_mai_n228_));
  NO3        m206(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n229_));
  NA2        m207(.A(i_2_), .B(i_1_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n226_), .B(mai_mai_n222_), .Y(mai_mai_n231_));
  NO3        m209(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n232_));
  NAi21      m210(.An(i_4_), .B(i_3_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n233_), .B(mai_mai_n72_), .Y(mai_mai_n234_));
  NO2        m212(.A(i_0_), .B(i_6_), .Y(mai_mai_n235_));
  NOi41      m213(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n236_));
  NA2        m214(.A(mai_mai_n236_), .B(mai_mai_n235_), .Y(mai_mai_n237_));
  NO2        m215(.A(mai_mai_n230_), .B(mai_mai_n177_), .Y(mai_mai_n238_));
  NAi21      m216(.An(mai_mai_n237_), .B(mai_mai_n238_), .Y(mai_mai_n239_));
  INV        m217(.A(mai_mai_n239_), .Y(mai_mai_n240_));
  AOI210     m218(.A0(mai_mai_n240_), .A1(mai_mai_n40_), .B0(mai_mai_n231_), .Y(mai_mai_n241_));
  NO2        m219(.A(i_11_), .B(mai_mai_n218_), .Y(mai_mai_n242_));
  NOi21      m220(.An(i_1_), .B(i_6_), .Y(mai_mai_n243_));
  NAi21      m221(.An(i_3_), .B(i_7_), .Y(mai_mai_n244_));
  NA2        m222(.A(mai_mai_n227_), .B(i_9_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n48_), .B(mai_mai_n25_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n70_), .B(i_5_), .Y(mai_mai_n247_));
  NA3        m225(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n223_), .B(mai_mai_n37_), .Y(mai_mai_n249_));
  NA2        m227(.A(i_12_), .B(i_6_), .Y(mai_mai_n250_));
  OR2        m228(.A(i_13_), .B(i_9_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n233_), .B(i_2_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n242_), .B(i_9_), .Y(mai_mai_n253_));
  NA2        m231(.A(mai_mai_n148_), .B(mai_mai_n60_), .Y(mai_mai_n254_));
  NO3        m232(.A(i_11_), .B(mai_mai_n218_), .C(mai_mai_n25_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n244_), .B(i_8_), .Y(mai_mai_n256_));
  NA3        m234(.A(i_5_), .B(mai_mai_n256_), .C(mai_mai_n255_), .Y(mai_mai_n257_));
  NO3        m235(.A(mai_mai_n26_), .B(mai_mai_n83_), .C(i_5_), .Y(mai_mai_n258_));
  NA3        m236(.A(mai_mai_n258_), .B(mai_mai_n249_), .C(mai_mai_n219_), .Y(mai_mai_n259_));
  AOI210     m237(.A0(mai_mai_n259_), .A1(mai_mai_n257_), .B0(mai_mai_n254_), .Y(mai_mai_n260_));
  INV        m238(.A(mai_mai_n260_), .Y(mai_mai_n261_));
  NA2        m239(.A(mai_mai_n261_), .B(mai_mai_n241_), .Y(mai_mai_n262_));
  NO3        m240(.A(i_12_), .B(mai_mai_n218_), .C(mai_mai_n37_), .Y(mai_mai_n263_));
  INV        m241(.A(mai_mai_n263_), .Y(mai_mai_n264_));
  NA2        m242(.A(i_8_), .B(mai_mai_n100_), .Y(mai_mai_n265_));
  NOi21      m243(.An(mai_mai_n157_), .B(mai_mai_n83_), .Y(mai_mai_n266_));
  NO3        m244(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n267_));
  AOI220     m245(.A0(mai_mai_n267_), .A1(mai_mai_n191_), .B0(mai_mai_n266_), .B1(mai_mai_n225_), .Y(mai_mai_n268_));
  NO2        m246(.A(mai_mai_n268_), .B(mai_mai_n265_), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n230_), .B(i_0_), .Y(mai_mai_n270_));
  NA2        m248(.A(i_0_), .B(i_1_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n271_), .B(i_2_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n56_), .B(i_6_), .Y(mai_mai_n273_));
  NA3        m251(.A(mai_mai_n273_), .B(mai_mai_n272_), .C(mai_mai_n157_), .Y(mai_mai_n274_));
  OAI210     m252(.A0(mai_mai_n159_), .A1(mai_mai_n137_), .B0(mai_mai_n274_), .Y(mai_mai_n275_));
  NO2        m253(.A(mai_mai_n275_), .B(mai_mai_n269_), .Y(mai_mai_n276_));
  NO2        m254(.A(i_3_), .B(i_10_), .Y(mai_mai_n277_));
  NA3        m255(.A(mai_mai_n277_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n278_));
  NO2        m256(.A(i_2_), .B(mai_mai_n100_), .Y(mai_mai_n279_));
  NA2        m257(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n280_), .B(i_8_), .Y(mai_mai_n281_));
  NA2        m259(.A(mai_mai_n281_), .B(mai_mai_n279_), .Y(mai_mai_n282_));
  AN2        m260(.A(i_3_), .B(i_10_), .Y(mai_mai_n283_));
  NA4        m261(.A(mai_mai_n283_), .B(mai_mai_n193_), .C(mai_mai_n170_), .D(mai_mai_n168_), .Y(mai_mai_n284_));
  NO2        m262(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n285_));
  NO2        m263(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n286_));
  OR2        m264(.A(mai_mai_n282_), .B(mai_mai_n278_), .Y(mai_mai_n287_));
  OAI220     m265(.A0(mai_mai_n287_), .A1(i_6_), .B0(mai_mai_n276_), .B1(mai_mai_n264_), .Y(mai_mai_n288_));
  NO4        m266(.A(mai_mai_n288_), .B(mai_mai_n262_), .C(mai_mai_n210_), .D(mai_mai_n162_), .Y(mai_mai_n289_));
  NO3        m267(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n290_));
  INV        m268(.A(mai_mai_n56_), .Y(mai_mai_n291_));
  NA2        m269(.A(mai_mai_n270_), .B(mai_mai_n291_), .Y(mai_mai_n292_));
  NO3        m270(.A(i_6_), .B(mai_mai_n188_), .C(i_7_), .Y(mai_mai_n293_));
  INV        m271(.A(mai_mai_n293_), .Y(mai_mai_n294_));
  AOI210     m272(.A0(mai_mai_n294_), .A1(mai_mai_n292_), .B0(mai_mai_n164_), .Y(mai_mai_n295_));
  NO2        m273(.A(i_2_), .B(i_3_), .Y(mai_mai_n296_));
  OR2        m274(.A(i_0_), .B(i_5_), .Y(mai_mai_n297_));
  NA2        m275(.A(mai_mai_n213_), .B(mai_mai_n297_), .Y(mai_mai_n298_));
  NA4        m276(.A(mai_mai_n298_), .B(mai_mai_n224_), .C(mai_mai_n296_), .D(i_1_), .Y(mai_mai_n299_));
  NA3        m277(.A(mai_mai_n270_), .B(mai_mai_n266_), .C(mai_mai_n112_), .Y(mai_mai_n300_));
  NAi21      m278(.An(i_8_), .B(i_7_), .Y(mai_mai_n301_));
  NO2        m279(.A(mai_mai_n301_), .B(i_6_), .Y(mai_mai_n302_));
  NO2        m280(.A(mai_mai_n151_), .B(mai_mai_n47_), .Y(mai_mai_n303_));
  NA3        m281(.A(mai_mai_n303_), .B(mai_mai_n302_), .C(mai_mai_n157_), .Y(mai_mai_n304_));
  NA3        m282(.A(mai_mai_n304_), .B(mai_mai_n300_), .C(mai_mai_n299_), .Y(mai_mai_n305_));
  OAI210     m283(.A0(mai_mai_n305_), .A1(mai_mai_n295_), .B0(i_4_), .Y(mai_mai_n306_));
  NO2        m284(.A(i_12_), .B(i_10_), .Y(mai_mai_n307_));
  NOi21      m285(.An(i_5_), .B(i_0_), .Y(mai_mai_n308_));
  NA4        m286(.A(mai_mai_n81_), .B(mai_mai_n36_), .C(mai_mai_n83_), .D(i_8_), .Y(mai_mai_n309_));
  NO2        m287(.A(i_6_), .B(i_8_), .Y(mai_mai_n310_));
  NOi21      m288(.An(i_0_), .B(i_2_), .Y(mai_mai_n311_));
  AN2        m289(.A(mai_mai_n311_), .B(mai_mai_n310_), .Y(mai_mai_n312_));
  NO2        m290(.A(i_1_), .B(i_7_), .Y(mai_mai_n313_));
  AO220      m291(.A0(mai_mai_n313_), .A1(mai_mai_n312_), .B0(mai_mai_n302_), .B1(mai_mai_n225_), .Y(mai_mai_n314_));
  NA3        m292(.A(mai_mai_n314_), .B(mai_mai_n42_), .C(i_5_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n315_), .B(mai_mai_n306_), .Y(mai_mai_n316_));
  NO3        m294(.A(mai_mai_n223_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n317_));
  NO3        m295(.A(mai_mai_n301_), .B(i_2_), .C(i_1_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n318_), .A1(mai_mai_n317_), .B0(i_6_), .Y(mai_mai_n319_));
  NO2        m297(.A(mai_mai_n319_), .B(mai_mai_n298_), .Y(mai_mai_n320_));
  NOi21      m298(.An(mai_mai_n147_), .B(mai_mai_n103_), .Y(mai_mai_n321_));
  NO2        m299(.A(mai_mai_n321_), .B(mai_mai_n119_), .Y(mai_mai_n322_));
  OAI210     m300(.A0(mai_mai_n322_), .A1(mai_mai_n320_), .B0(i_3_), .Y(mai_mai_n323_));
  INV        m301(.A(mai_mai_n81_), .Y(mai_mai_n324_));
  NO2        m302(.A(mai_mai_n271_), .B(mai_mai_n78_), .Y(mai_mai_n325_));
  NA2        m303(.A(mai_mai_n325_), .B(mai_mai_n127_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n92_), .B(mai_mai_n188_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n327_), .B(mai_mai_n60_), .Y(mai_mai_n328_));
  AOI210     m306(.A0(mai_mai_n328_), .A1(mai_mai_n326_), .B0(mai_mai_n324_), .Y(mai_mai_n329_));
  NO2        m307(.A(mai_mai_n188_), .B(i_9_), .Y(mai_mai_n330_));
  NA2        m308(.A(mai_mai_n330_), .B(mai_mai_n200_), .Y(mai_mai_n331_));
  NO2        m309(.A(mai_mai_n331_), .B(mai_mai_n47_), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n332_), .B(mai_mai_n329_), .Y(mai_mai_n333_));
  AOI210     m311(.A0(mai_mai_n333_), .A1(mai_mai_n323_), .B0(mai_mai_n156_), .Y(mai_mai_n334_));
  AOI210     m312(.A0(mai_mai_n316_), .A1(mai_mai_n290_), .B0(mai_mai_n334_), .Y(mai_mai_n335_));
  NOi32      m313(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n336_));
  INV        m314(.A(mai_mai_n336_), .Y(mai_mai_n337_));
  NAi21      m315(.An(i_1_), .B(i_5_), .Y(mai_mai_n338_));
  NAi41      m316(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n339_));
  OAI220     m317(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n214_), .B1(mai_mai_n153_), .Y(mai_mai_n340_));
  NO2        m318(.A(mai_mai_n153_), .B(mai_mai_n151_), .Y(mai_mai_n341_));
  NOi32      m319(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n342_));
  NAi21      m320(.An(i_6_), .B(i_1_), .Y(mai_mai_n343_));
  NA3        m321(.A(mai_mai_n343_), .B(mai_mai_n342_), .C(mai_mai_n47_), .Y(mai_mai_n344_));
  NO2        m322(.A(mai_mai_n344_), .B(i_0_), .Y(mai_mai_n345_));
  OR3        m323(.A(mai_mai_n345_), .B(mai_mai_n341_), .C(mai_mai_n340_), .Y(mai_mai_n346_));
  NO2        m324(.A(i_1_), .B(mai_mai_n100_), .Y(mai_mai_n347_));
  NAi21      m325(.An(i_3_), .B(i_4_), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(i_9_), .Y(mai_mai_n349_));
  AN2        m327(.A(i_6_), .B(i_7_), .Y(mai_mai_n350_));
  NA2        m328(.A(i_2_), .B(i_7_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n348_), .B(i_10_), .Y(mai_mai_n352_));
  AOI210     m330(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n353_));
  OAI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n183_), .B0(mai_mai_n352_), .Y(mai_mai_n354_));
  AOI220     m332(.A0(mai_mai_n352_), .A1(mai_mai_n313_), .B0(mai_mai_n229_), .B1(mai_mai_n183_), .Y(mai_mai_n355_));
  AOI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n354_), .B0(i_5_), .Y(mai_mai_n356_));
  NO3        m334(.A(mai_mai_n356_), .B(mai_mai_n346_), .C(mai_mai_n987_), .Y(mai_mai_n357_));
  NO2        m335(.A(mai_mai_n357_), .B(mai_mai_n337_), .Y(mai_mai_n358_));
  NO2        m336(.A(mai_mai_n56_), .B(mai_mai_n25_), .Y(mai_mai_n359_));
  AN2        m337(.A(i_12_), .B(i_5_), .Y(mai_mai_n360_));
  NO2        m338(.A(i_11_), .B(i_6_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n233_), .B(i_5_), .Y(mai_mai_n362_));
  NO2        m340(.A(i_5_), .B(i_10_), .Y(mai_mai_n363_));
  AOI220     m341(.A0(mai_mai_n363_), .A1(mai_mai_n252_), .B0(mai_mai_n362_), .B1(mai_mai_n193_), .Y(mai_mai_n364_));
  NA2        m342(.A(mai_mai_n138_), .B(mai_mai_n46_), .Y(mai_mai_n365_));
  NO2        m343(.A(mai_mai_n365_), .B(mai_mai_n364_), .Y(mai_mai_n366_));
  NA2        m344(.A(mai_mai_n366_), .B(mai_mai_n359_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n368_));
  NO3        m346(.A(mai_mai_n83_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n369_));
  NO2        m347(.A(i_3_), .B(mai_mai_n100_), .Y(mai_mai_n370_));
  NO2        m348(.A(i_11_), .B(i_12_), .Y(mai_mai_n371_));
  NA3        m349(.A(mai_mai_n112_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n372_));
  NO2        m350(.A(mai_mai_n372_), .B(mai_mai_n214_), .Y(mai_mai_n373_));
  NAi21      m351(.An(i_13_), .B(i_0_), .Y(mai_mai_n374_));
  INV        m352(.A(mai_mai_n374_), .Y(mai_mai_n375_));
  NA2        m353(.A(mai_mai_n373_), .B(mai_mai_n375_), .Y(mai_mai_n376_));
  NA2        m354(.A(mai_mai_n376_), .B(mai_mai_n367_), .Y(mai_mai_n377_));
  NO3        m355(.A(i_1_), .B(i_12_), .C(mai_mai_n83_), .Y(mai_mai_n378_));
  NO2        m356(.A(i_0_), .B(i_11_), .Y(mai_mai_n379_));
  AN2        m357(.A(i_1_), .B(i_6_), .Y(mai_mai_n380_));
  NOi21      m358(.An(i_2_), .B(i_12_), .Y(mai_mai_n381_));
  NA2        m359(.A(mai_mai_n381_), .B(mai_mai_n380_), .Y(mai_mai_n382_));
  INV        m360(.A(mai_mai_n382_), .Y(mai_mai_n383_));
  NA2        m361(.A(mai_mai_n136_), .B(i_9_), .Y(mai_mai_n384_));
  NO2        m362(.A(mai_mai_n384_), .B(i_4_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n383_), .B(mai_mai_n385_), .Y(mai_mai_n386_));
  NAi21      m364(.An(i_9_), .B(i_4_), .Y(mai_mai_n387_));
  OR2        m365(.A(i_13_), .B(i_10_), .Y(mai_mai_n388_));
  NO3        m366(.A(mai_mai_n388_), .B(mai_mai_n114_), .C(mai_mai_n387_), .Y(mai_mai_n389_));
  OR2        m367(.A(mai_mai_n212_), .B(mai_mai_n211_), .Y(mai_mai_n390_));
  NO2        m368(.A(mai_mai_n100_), .B(mai_mai_n25_), .Y(mai_mai_n391_));
  NA2        m369(.A(mai_mai_n263_), .B(mai_mai_n391_), .Y(mai_mai_n392_));
  NA2        m370(.A(i_5_), .B(mai_mai_n206_), .Y(mai_mai_n393_));
  OAI220     m371(.A0(mai_mai_n393_), .A1(mai_mai_n390_), .B0(mai_mai_n392_), .B1(mai_mai_n321_), .Y(mai_mai_n394_));
  INV        m372(.A(mai_mai_n394_), .Y(mai_mai_n395_));
  AOI210     m373(.A0(mai_mai_n395_), .A1(mai_mai_n386_), .B0(mai_mai_n26_), .Y(mai_mai_n396_));
  NA2        m374(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n397_));
  AOI220     m375(.A0(mai_mai_n273_), .A1(mai_mai_n267_), .B0(mai_mai_n270_), .B1(mai_mai_n291_), .Y(mai_mai_n398_));
  NO2        m376(.A(mai_mai_n398_), .B(mai_mai_n164_), .Y(mai_mai_n399_));
  AOI220     m377(.A0(i_3_), .A1(mai_mai_n272_), .B0(mai_mai_n258_), .B1(mai_mai_n206_), .Y(mai_mai_n400_));
  NO2        m378(.A(mai_mai_n400_), .B(mai_mai_n265_), .Y(mai_mai_n401_));
  NO3        m379(.A(mai_mai_n401_), .B(mai_mai_n399_), .C(mai_mai_n397_), .Y(mai_mai_n402_));
  NA2        m380(.A(mai_mai_n191_), .B(mai_mai_n95_), .Y(mai_mai_n403_));
  NA3        m381(.A(mai_mai_n303_), .B(mai_mai_n157_), .C(mai_mai_n83_), .Y(mai_mai_n404_));
  AOI210     m382(.A0(mai_mai_n404_), .A1(mai_mai_n403_), .B0(mai_mai_n301_), .Y(mai_mai_n405_));
  NA2        m383(.A(mai_mai_n188_), .B(i_10_), .Y(mai_mai_n406_));
  NA3        m384(.A(mai_mai_n247_), .B(mai_mai_n61_), .C(i_2_), .Y(mai_mai_n407_));
  NA2        m385(.A(mai_mai_n273_), .B(mai_mai_n225_), .Y(mai_mai_n408_));
  OAI220     m386(.A0(mai_mai_n408_), .A1(mai_mai_n177_), .B0(mai_mai_n407_), .B1(mai_mai_n406_), .Y(mai_mai_n409_));
  NA3        m387(.A(mai_mai_n313_), .B(mai_mai_n312_), .C(i_5_), .Y(mai_mai_n410_));
  NA2        m388(.A(mai_mai_n293_), .B(mai_mai_n298_), .Y(mai_mai_n411_));
  OAI210     m389(.A0(mai_mai_n411_), .A1(mai_mai_n184_), .B0(mai_mai_n410_), .Y(mai_mai_n412_));
  NO3        m390(.A(mai_mai_n412_), .B(mai_mai_n409_), .C(mai_mai_n405_), .Y(mai_mai_n413_));
  AOI210     m391(.A0(mai_mai_n413_), .A1(mai_mai_n402_), .B0(mai_mai_n253_), .Y(mai_mai_n414_));
  NO4        m392(.A(mai_mai_n414_), .B(mai_mai_n396_), .C(mai_mai_n377_), .D(mai_mai_n358_), .Y(mai_mai_n415_));
  NO2        m393(.A(mai_mai_n70_), .B(i_13_), .Y(mai_mai_n416_));
  NO2        m394(.A(i_10_), .B(i_9_), .Y(mai_mai_n417_));
  NAi21      m395(.An(i_12_), .B(i_8_), .Y(mai_mai_n418_));
  NO2        m396(.A(mai_mai_n418_), .B(i_3_), .Y(mai_mai_n419_));
  INV        m397(.A(i_0_), .Y(mai_mai_n420_));
  NO3        m398(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n421_));
  NA2        m399(.A(mai_mai_n250_), .B(mai_mai_n96_), .Y(mai_mai_n422_));
  NA2        m400(.A(mai_mai_n422_), .B(mai_mai_n421_), .Y(mai_mai_n423_));
  NA2        m401(.A(i_8_), .B(i_9_), .Y(mai_mai_n424_));
  NA2        m402(.A(mai_mai_n263_), .B(mai_mai_n200_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n425_), .B(mai_mai_n424_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n242_), .B(mai_mai_n285_), .Y(mai_mai_n427_));
  NO3        m405(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n428_));
  INV        m406(.A(mai_mai_n428_), .Y(mai_mai_n429_));
  NA3        m407(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n430_));
  NO2        m408(.A(mai_mai_n429_), .B(mai_mai_n427_), .Y(mai_mai_n431_));
  NO2        m409(.A(mai_mai_n431_), .B(mai_mai_n426_), .Y(mai_mai_n432_));
  NA2        m410(.A(mai_mai_n272_), .B(mai_mai_n107_), .Y(mai_mai_n433_));
  OR2        m411(.A(mai_mai_n433_), .B(mai_mai_n202_), .Y(mai_mai_n434_));
  OA210      m412(.A0(mai_mai_n331_), .A1(mai_mai_n100_), .B0(mai_mai_n274_), .Y(mai_mai_n435_));
  OA220      m413(.A0(mai_mai_n435_), .A1(mai_mai_n156_), .B0(mai_mai_n434_), .B1(mai_mai_n222_), .Y(mai_mai_n436_));
  NA2        m414(.A(mai_mai_n95_), .B(i_13_), .Y(mai_mai_n437_));
  NO2        m415(.A(i_2_), .B(i_13_), .Y(mai_mai_n438_));
  NO3        m416(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n439_));
  NO2        m417(.A(i_6_), .B(i_7_), .Y(mai_mai_n440_));
  NA2        m418(.A(mai_mai_n440_), .B(mai_mai_n439_), .Y(mai_mai_n441_));
  NO2        m419(.A(i_11_), .B(i_1_), .Y(mai_mai_n442_));
  OR2        m420(.A(i_11_), .B(i_8_), .Y(mai_mai_n443_));
  NOi21      m421(.An(i_2_), .B(i_7_), .Y(mai_mai_n444_));
  NAi31      m422(.An(mai_mai_n443_), .B(mai_mai_n444_), .C(i_0_), .Y(mai_mai_n445_));
  NO2        m423(.A(mai_mai_n388_), .B(i_6_), .Y(mai_mai_n446_));
  NA3        m424(.A(mai_mai_n446_), .B(i_1_), .C(mai_mai_n72_), .Y(mai_mai_n447_));
  NO2        m425(.A(mai_mai_n447_), .B(mai_mai_n445_), .Y(mai_mai_n448_));
  NO2        m426(.A(i_3_), .B(mai_mai_n188_), .Y(mai_mai_n449_));
  NO2        m427(.A(i_6_), .B(i_10_), .Y(mai_mai_n450_));
  NA4        m428(.A(mai_mai_n450_), .B(mai_mai_n290_), .C(mai_mai_n449_), .D(mai_mai_n227_), .Y(mai_mai_n451_));
  NO2        m429(.A(mai_mai_n451_), .B(mai_mai_n149_), .Y(mai_mai_n452_));
  NA3        m430(.A(mai_mai_n236_), .B(mai_mai_n166_), .C(mai_mai_n127_), .Y(mai_mai_n453_));
  NA2        m431(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n454_));
  NO2        m432(.A(mai_mai_n151_), .B(i_3_), .Y(mai_mai_n455_));
  NAi31      m433(.An(mai_mai_n454_), .B(mai_mai_n455_), .C(mai_mai_n219_), .Y(mai_mai_n456_));
  NA3        m434(.A(mai_mai_n368_), .B(mai_mai_n173_), .C(mai_mai_n143_), .Y(mai_mai_n457_));
  NA3        m435(.A(mai_mai_n457_), .B(mai_mai_n456_), .C(mai_mai_n453_), .Y(mai_mai_n458_));
  NO3        m436(.A(mai_mai_n458_), .B(mai_mai_n452_), .C(mai_mai_n448_), .Y(mai_mai_n459_));
  NA2        m437(.A(mai_mai_n421_), .B(mai_mai_n360_), .Y(mai_mai_n460_));
  NAi21      m438(.An(mai_mai_n212_), .B(mai_mai_n371_), .Y(mai_mai_n461_));
  NO2        m439(.A(mai_mai_n26_), .B(i_5_), .Y(mai_mai_n462_));
  NO2        m440(.A(i_0_), .B(mai_mai_n83_), .Y(mai_mai_n463_));
  NA3        m441(.A(mai_mai_n463_), .B(mai_mai_n462_), .C(mai_mai_n136_), .Y(mai_mai_n464_));
  OR3        m442(.A(mai_mai_n280_), .B(mai_mai_n38_), .C(mai_mai_n47_), .Y(mai_mai_n465_));
  NO2        m443(.A(mai_mai_n465_), .B(mai_mai_n464_), .Y(mai_mai_n466_));
  NA2        m444(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n467_));
  NA2        m445(.A(mai_mai_n290_), .B(mai_mai_n229_), .Y(mai_mai_n468_));
  OAI220     m446(.A0(mai_mai_n468_), .A1(mai_mai_n407_), .B0(mai_mai_n467_), .B1(mai_mai_n437_), .Y(mai_mai_n469_));
  NA4        m447(.A(mai_mai_n283_), .B(mai_mai_n217_), .C(mai_mai_n70_), .D(mai_mai_n227_), .Y(mai_mai_n470_));
  NO2        m448(.A(mai_mai_n470_), .B(mai_mai_n441_), .Y(mai_mai_n471_));
  NO3        m449(.A(mai_mai_n471_), .B(mai_mai_n469_), .C(mai_mai_n466_), .Y(mai_mai_n472_));
  NA4        m450(.A(mai_mai_n472_), .B(mai_mai_n459_), .C(mai_mai_n436_), .D(mai_mai_n432_), .Y(mai_mai_n473_));
  NA3        m451(.A(mai_mai_n283_), .B(mai_mai_n170_), .C(mai_mai_n168_), .Y(mai_mai_n474_));
  OAI210     m452(.A0(mai_mai_n278_), .A1(mai_mai_n175_), .B0(mai_mai_n474_), .Y(mai_mai_n475_));
  AN2        m453(.A(mai_mai_n267_), .B(mai_mai_n224_), .Y(mai_mai_n476_));
  NA2        m454(.A(mai_mai_n476_), .B(mai_mai_n475_), .Y(mai_mai_n477_));
  NA2        m455(.A(mai_mai_n290_), .B(mai_mai_n158_), .Y(mai_mai_n478_));
  OAI210     m456(.A0(mai_mai_n478_), .A1(mai_mai_n222_), .B0(mai_mai_n284_), .Y(mai_mai_n479_));
  NA2        m457(.A(mai_mai_n479_), .B(mai_mai_n302_), .Y(mai_mai_n480_));
  NA2        m458(.A(mai_mai_n360_), .B(mai_mai_n218_), .Y(mai_mai_n481_));
  NA2        m459(.A(mai_mai_n336_), .B(mai_mai_n70_), .Y(mai_mai_n482_));
  NA2        m460(.A(mai_mai_n350_), .B(mai_mai_n342_), .Y(mai_mai_n483_));
  OR2        m461(.A(mai_mai_n481_), .B(mai_mai_n483_), .Y(mai_mai_n484_));
  NO2        m462(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n485_));
  NAi41      m463(.An(mai_mai_n482_), .B(mai_mai_n450_), .C(mai_mai_n485_), .D(mai_mai_n47_), .Y(mai_mai_n486_));
  AOI210     m464(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n389_), .Y(mai_mai_n487_));
  NA3        m465(.A(mai_mai_n487_), .B(mai_mai_n486_), .C(mai_mai_n484_), .Y(mai_mai_n488_));
  INV        m466(.A(mai_mai_n488_), .Y(mai_mai_n489_));
  AOI210     m467(.A0(mai_mai_n189_), .A1(i_9_), .B0(mai_mai_n249_), .Y(mai_mai_n490_));
  NO2        m468(.A(mai_mai_n490_), .B(mai_mai_n194_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n177_), .B(mai_mai_n83_), .Y(mai_mai_n492_));
  NA2        m470(.A(mai_mai_n492_), .B(mai_mai_n491_), .Y(mai_mai_n493_));
  NA4        m471(.A(mai_mai_n493_), .B(mai_mai_n489_), .C(mai_mai_n480_), .D(mai_mai_n477_), .Y(mai_mai_n494_));
  NA2        m472(.A(mai_mai_n362_), .B(mai_mai_n272_), .Y(mai_mai_n495_));
  NA2        m473(.A(mai_mai_n163_), .B(mai_mai_n495_), .Y(mai_mai_n496_));
  NO2        m474(.A(i_12_), .B(mai_mai_n188_), .Y(mai_mai_n497_));
  NA2        m475(.A(mai_mai_n497_), .B(mai_mai_n218_), .Y(mai_mai_n498_));
  NO3        m476(.A(i_6_), .B(mai_mai_n498_), .C(mai_mai_n433_), .Y(mai_mai_n499_));
  NOi31      m477(.An(mai_mai_n293_), .B(mai_mai_n388_), .C(mai_mai_n38_), .Y(mai_mai_n500_));
  OAI210     m478(.A0(mai_mai_n500_), .A1(mai_mai_n499_), .B0(mai_mai_n496_), .Y(mai_mai_n501_));
  NO2        m479(.A(i_8_), .B(i_7_), .Y(mai_mai_n502_));
  INV        m480(.A(i_5_), .Y(mai_mai_n503_));
  NA2        m481(.A(mai_mai_n503_), .B(mai_mai_n217_), .Y(mai_mai_n504_));
  AOI220     m482(.A0(mai_mai_n303_), .A1(mai_mai_n40_), .B0(mai_mai_n225_), .B1(mai_mai_n201_), .Y(mai_mai_n505_));
  OAI220     m483(.A0(mai_mai_n505_), .A1(mai_mai_n177_), .B0(mai_mai_n504_), .B1(mai_mai_n233_), .Y(mai_mai_n506_));
  NA2        m484(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n507_));
  NO2        m485(.A(mai_mai_n507_), .B(i_6_), .Y(mai_mai_n508_));
  NA3        m486(.A(mai_mai_n508_), .B(mai_mai_n506_), .C(mai_mai_n502_), .Y(mai_mai_n509_));
  NO2        m487(.A(mai_mai_n437_), .B(mai_mai_n128_), .Y(mai_mai_n510_));
  NA2        m488(.A(mai_mai_n510_), .B(mai_mai_n249_), .Y(mai_mai_n511_));
  NOi31      m489(.An(mai_mai_n270_), .B(mai_mai_n278_), .C(mai_mai_n175_), .Y(mai_mai_n512_));
  NA2        m490(.A(mai_mai_n512_), .B(mai_mai_n428_), .Y(mai_mai_n513_));
  NA4        m491(.A(mai_mai_n513_), .B(mai_mai_n511_), .C(mai_mai_n509_), .D(mai_mai_n501_), .Y(mai_mai_n514_));
  NA3        m492(.A(mai_mai_n213_), .B(mai_mai_n68_), .C(mai_mai_n45_), .Y(mai_mai_n515_));
  NA2        m493(.A(mai_mai_n263_), .B(mai_mai_n81_), .Y(mai_mai_n516_));
  AOI210     m494(.A0(mai_mai_n515_), .A1(mai_mai_n326_), .B0(mai_mai_n516_), .Y(mai_mai_n517_));
  NA2        m495(.A(mai_mai_n273_), .B(mai_mai_n267_), .Y(mai_mai_n518_));
  NO2        m496(.A(mai_mai_n518_), .B(mai_mai_n167_), .Y(mai_mai_n519_));
  NA2        m497(.A(mai_mai_n217_), .B(mai_mai_n216_), .Y(mai_mai_n520_));
  NA2        m498(.A(mai_mai_n417_), .B(mai_mai_n215_), .Y(mai_mai_n521_));
  NO2        m499(.A(mai_mai_n520_), .B(mai_mai_n521_), .Y(mai_mai_n522_));
  AOI210     m500(.A0(mai_mai_n343_), .A1(mai_mai_n47_), .B0(mai_mai_n347_), .Y(mai_mai_n523_));
  NA2        m501(.A(i_0_), .B(mai_mai_n48_), .Y(mai_mai_n524_));
  NA3        m502(.A(mai_mai_n497_), .B(mai_mai_n255_), .C(mai_mai_n524_), .Y(mai_mai_n525_));
  NO2        m503(.A(mai_mai_n523_), .B(mai_mai_n525_), .Y(mai_mai_n526_));
  NO4        m504(.A(mai_mai_n526_), .B(mai_mai_n522_), .C(mai_mai_n519_), .D(mai_mai_n517_), .Y(mai_mai_n527_));
  NO4        m505(.A(mai_mai_n243_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n528_));
  NO3        m506(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n529_));
  NO2        m507(.A(mai_mai_n223_), .B(mai_mai_n36_), .Y(mai_mai_n530_));
  AN2        m508(.A(mai_mai_n530_), .B(mai_mai_n529_), .Y(mai_mai_n531_));
  OA210      m509(.A0(mai_mai_n531_), .A1(mai_mai_n528_), .B0(mai_mai_n336_), .Y(mai_mai_n532_));
  NO2        m510(.A(mai_mai_n388_), .B(i_1_), .Y(mai_mai_n533_));
  NOi31      m511(.An(mai_mai_n533_), .B(mai_mai_n422_), .C(mai_mai_n70_), .Y(mai_mai_n534_));
  AN4        m512(.A(mai_mai_n534_), .B(mai_mai_n385_), .C(mai_mai_n462_), .D(i_2_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n398_), .B(mai_mai_n171_), .Y(mai_mai_n536_));
  NO3        m514(.A(mai_mai_n536_), .B(mai_mai_n535_), .C(mai_mai_n532_), .Y(mai_mai_n537_));
  NO2        m515(.A(mai_mai_n113_), .B(mai_mai_n23_), .Y(mai_mai_n538_));
  NA2        m516(.A(mai_mai_n293_), .B(mai_mai_n158_), .Y(mai_mai_n539_));
  AOI220     m517(.A0(mai_mai_n539_), .A1(mai_mai_n408_), .B0(mai_mai_n178_), .B1(mai_mai_n176_), .Y(mai_mai_n540_));
  NO2        m518(.A(mai_mai_n193_), .B(mai_mai_n37_), .Y(mai_mai_n541_));
  NOi31      m519(.An(mai_mai_n140_), .B(mai_mai_n541_), .C(mai_mai_n309_), .Y(mai_mai_n542_));
  NO2        m520(.A(mai_mai_n542_), .B(mai_mai_n540_), .Y(mai_mai_n543_));
  INV        m521(.A(mai_mai_n296_), .Y(mai_mai_n544_));
  NO2        m522(.A(i_12_), .B(mai_mai_n83_), .Y(mai_mai_n545_));
  NA3        m523(.A(mai_mai_n545_), .B(mai_mai_n255_), .C(mai_mai_n524_), .Y(mai_mai_n546_));
  NA3        m524(.A(mai_mai_n361_), .B(mai_mai_n263_), .C(mai_mai_n213_), .Y(mai_mai_n547_));
  AOI210     m525(.A0(mai_mai_n547_), .A1(mai_mai_n546_), .B0(mai_mai_n544_), .Y(mai_mai_n548_));
  NA2        m526(.A(mai_mai_n168_), .B(i_0_), .Y(mai_mai_n549_));
  NO3        m527(.A(mai_mai_n549_), .B(mai_mai_n319_), .C(mai_mai_n278_), .Y(mai_mai_n550_));
  OR2        m528(.A(i_2_), .B(i_5_), .Y(mai_mai_n551_));
  OR2        m529(.A(mai_mai_n551_), .B(mai_mai_n380_), .Y(mai_mai_n552_));
  AOI210     m530(.A0(mai_mai_n351_), .A1(mai_mai_n235_), .B0(mai_mai_n193_), .Y(mai_mai_n553_));
  AOI210     m531(.A0(mai_mai_n553_), .A1(mai_mai_n552_), .B0(mai_mai_n461_), .Y(mai_mai_n554_));
  NO3        m532(.A(mai_mai_n554_), .B(mai_mai_n550_), .C(mai_mai_n548_), .Y(mai_mai_n555_));
  NA4        m533(.A(mai_mai_n555_), .B(mai_mai_n543_), .C(mai_mai_n537_), .D(mai_mai_n527_), .Y(mai_mai_n556_));
  NO4        m534(.A(mai_mai_n556_), .B(mai_mai_n514_), .C(mai_mai_n494_), .D(mai_mai_n473_), .Y(mai_mai_n557_));
  NA4        m535(.A(mai_mai_n557_), .B(mai_mai_n415_), .C(mai_mai_n335_), .D(mai_mai_n289_), .Y(mai7));
  NO2        m536(.A(mai_mai_n92_), .B(mai_mai_n52_), .Y(mai_mai_n559_));
  NO2        m537(.A(mai_mai_n107_), .B(mai_mai_n89_), .Y(mai_mai_n560_));
  NA2        m538(.A(i_3_), .B(mai_mai_n560_), .Y(mai_mai_n561_));
  NA2        m539(.A(mai_mai_n450_), .B(mai_mai_n81_), .Y(mai_mai_n562_));
  NA2        m540(.A(i_11_), .B(mai_mai_n188_), .Y(mai_mai_n563_));
  NA2        m541(.A(mai_mai_n138_), .B(mai_mai_n563_), .Y(mai_mai_n564_));
  OAI210     m542(.A0(mai_mai_n564_), .A1(mai_mai_n562_), .B0(mai_mai_n561_), .Y(mai_mai_n565_));
  NA3        m543(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n566_));
  NO2        m544(.A(mai_mai_n227_), .B(i_4_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n567_), .B(i_8_), .Y(mai_mai_n568_));
  NO2        m546(.A(mai_mai_n104_), .B(mai_mai_n566_), .Y(mai_mai_n569_));
  NA2        m547(.A(i_2_), .B(mai_mai_n83_), .Y(mai_mai_n570_));
  OAI210     m548(.A0(mai_mai_n86_), .A1(mai_mai_n198_), .B0(mai_mai_n199_), .Y(mai_mai_n571_));
  NO2        m549(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n572_));
  NA2        m550(.A(i_4_), .B(i_8_), .Y(mai_mai_n573_));
  NO3        m551(.A(mai_mai_n569_), .B(mai_mai_n565_), .C(mai_mai_n559_), .Y(mai_mai_n574_));
  AOI210     m552(.A0(mai_mai_n123_), .A1(mai_mai_n59_), .B0(i_10_), .Y(mai_mai_n575_));
  AOI210     m553(.A0(mai_mai_n575_), .A1(mai_mai_n227_), .B0(mai_mai_n155_), .Y(mai_mai_n576_));
  OR2        m554(.A(i_6_), .B(i_10_), .Y(mai_mai_n577_));
  NO2        m555(.A(mai_mai_n577_), .B(mai_mai_n23_), .Y(mai_mai_n578_));
  OR3        m556(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n579_));
  NO3        m557(.A(mai_mai_n579_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n580_));
  INV        m558(.A(mai_mai_n195_), .Y(mai_mai_n581_));
  NO2        m559(.A(mai_mai_n580_), .B(mai_mai_n578_), .Y(mai_mai_n582_));
  OA220      m560(.A0(mai_mai_n582_), .A1(mai_mai_n544_), .B0(mai_mai_n576_), .B1(mai_mai_n251_), .Y(mai_mai_n583_));
  AOI210     m561(.A0(mai_mai_n583_), .A1(mai_mai_n574_), .B0(mai_mai_n60_), .Y(mai_mai_n584_));
  NOi21      m562(.An(i_11_), .B(i_7_), .Y(mai_mai_n585_));
  AO210      m563(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n586_));
  NO2        m564(.A(mai_mai_n586_), .B(mai_mai_n585_), .Y(mai_mai_n587_));
  NA2        m565(.A(mai_mai_n587_), .B(mai_mai_n201_), .Y(mai_mai_n588_));
  NA3        m566(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n589_));
  NO2        m567(.A(mai_mai_n588_), .B(mai_mai_n60_), .Y(mai_mai_n590_));
  NA2        m568(.A(mai_mai_n85_), .B(mai_mai_n60_), .Y(mai_mai_n591_));
  AO210      m569(.A0(mai_mai_n591_), .A1(mai_mai_n355_), .B0(mai_mai_n41_), .Y(mai_mai_n592_));
  NA2        m570(.A(mai_mai_n219_), .B(mai_mai_n60_), .Y(mai_mai_n593_));
  NO2        m571(.A(mai_mai_n60_), .B(i_9_), .Y(mai_mai_n594_));
  NO2        m572(.A(i_1_), .B(i_12_), .Y(mai_mai_n595_));
  NA3        m573(.A(mai_mai_n595_), .B(mai_mai_n109_), .C(mai_mai_n24_), .Y(mai_mai_n596_));
  BUFFER     m574(.A(mai_mai_n596_), .Y(mai_mai_n597_));
  NA3        m575(.A(mai_mai_n597_), .B(mai_mai_n593_), .C(mai_mai_n592_), .Y(mai_mai_n598_));
  OAI210     m576(.A0(mai_mai_n598_), .A1(mai_mai_n590_), .B0(i_6_), .Y(mai_mai_n599_));
  NO2        m577(.A(mai_mai_n589_), .B(mai_mai_n107_), .Y(mai_mai_n600_));
  NA2        m578(.A(mai_mai_n600_), .B(mai_mai_n545_), .Y(mai_mai_n601_));
  NO2        m579(.A(i_6_), .B(i_11_), .Y(mai_mai_n602_));
  NA2        m580(.A(mai_mai_n601_), .B(mai_mai_n423_), .Y(mai_mai_n603_));
  NO4        m581(.A(mai_mai_n211_), .B(mai_mai_n123_), .C(i_13_), .D(mai_mai_n83_), .Y(mai_mai_n604_));
  NA2        m582(.A(mai_mai_n604_), .B(mai_mai_n594_), .Y(mai_mai_n605_));
  INV        m583(.A(mai_mai_n605_), .Y(mai_mai_n606_));
  NA3        m584(.A(mai_mai_n502_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n607_));
  INV        m585(.A(i_2_), .Y(mai_mai_n608_));
  NA2        m586(.A(mai_mai_n132_), .B(i_9_), .Y(mai_mai_n609_));
  NA3        m587(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n610_));
  NO2        m588(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n611_));
  NA3        m589(.A(mai_mai_n611_), .B(mai_mai_n250_), .C(mai_mai_n45_), .Y(mai_mai_n612_));
  OAI220     m590(.A0(mai_mai_n612_), .A1(mai_mai_n610_), .B0(mai_mai_n609_), .B1(mai_mai_n608_), .Y(mai_mai_n613_));
  NA3        m591(.A(mai_mai_n594_), .B(mai_mai_n296_), .C(i_6_), .Y(mai_mai_n614_));
  NO2        m592(.A(mai_mai_n614_), .B(mai_mai_n23_), .Y(mai_mai_n615_));
  AOI210     m593(.A0(mai_mai_n442_), .A1(mai_mai_n391_), .B0(mai_mai_n232_), .Y(mai_mai_n616_));
  NO2        m594(.A(mai_mai_n616_), .B(mai_mai_n570_), .Y(mai_mai_n617_));
  NAi21      m595(.An(mai_mai_n607_), .B(mai_mai_n91_), .Y(mai_mai_n618_));
  NA2        m596(.A(mai_mai_n611_), .B(mai_mai_n250_), .Y(mai_mai_n619_));
  NO2        m597(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n620_));
  NA2        m598(.A(mai_mai_n620_), .B(mai_mai_n24_), .Y(mai_mai_n621_));
  OAI210     m599(.A0(mai_mai_n621_), .A1(mai_mai_n619_), .B0(mai_mai_n618_), .Y(mai_mai_n622_));
  OR4        m600(.A(mai_mai_n622_), .B(mai_mai_n617_), .C(mai_mai_n615_), .D(mai_mai_n613_), .Y(mai_mai_n623_));
  NO3        m601(.A(mai_mai_n623_), .B(mai_mai_n606_), .C(mai_mai_n603_), .Y(mai_mai_n624_));
  NO2        m602(.A(mai_mai_n227_), .B(mai_mai_n100_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n625_), .B(mai_mai_n585_), .Y(mai_mai_n626_));
  NA2        m604(.A(mai_mai_n626_), .B(i_1_), .Y(mai_mai_n627_));
  NO2        m605(.A(mai_mai_n627_), .B(mai_mai_n579_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n387_), .B(mai_mai_n83_), .Y(mai_mai_n629_));
  NA2        m607(.A(mai_mai_n628_), .B(mai_mai_n47_), .Y(mai_mai_n630_));
  NA2        m608(.A(i_3_), .B(mai_mai_n188_), .Y(mai_mai_n631_));
  NO2        m609(.A(mai_mai_n631_), .B(mai_mai_n113_), .Y(mai_mai_n632_));
  AN2        m610(.A(mai_mai_n632_), .B(mai_mai_n508_), .Y(mai_mai_n633_));
  NO2        m611(.A(mai_mai_n223_), .B(mai_mai_n45_), .Y(mai_mai_n634_));
  NO3        m612(.A(mai_mai_n634_), .B(mai_mai_n286_), .C(mai_mai_n228_), .Y(mai_mai_n635_));
  NO2        m613(.A(mai_mai_n114_), .B(mai_mai_n37_), .Y(mai_mai_n636_));
  NO2        m614(.A(mai_mai_n636_), .B(i_6_), .Y(mai_mai_n637_));
  NO2        m615(.A(mai_mai_n83_), .B(i_9_), .Y(mai_mai_n638_));
  NO2        m616(.A(mai_mai_n638_), .B(mai_mai_n60_), .Y(mai_mai_n639_));
  NO2        m617(.A(mai_mai_n639_), .B(mai_mai_n595_), .Y(mai_mai_n640_));
  NO4        m618(.A(mai_mai_n640_), .B(mai_mai_n637_), .C(mai_mai_n635_), .D(i_4_), .Y(mai_mai_n641_));
  NA2        m619(.A(i_1_), .B(i_3_), .Y(mai_mai_n642_));
  NO2        m620(.A(mai_mai_n424_), .B(mai_mai_n92_), .Y(mai_mai_n643_));
  INV        m621(.A(mai_mai_n643_), .Y(mai_mai_n644_));
  NO2        m622(.A(mai_mai_n644_), .B(mai_mai_n642_), .Y(mai_mai_n645_));
  NO3        m623(.A(mai_mai_n645_), .B(mai_mai_n641_), .C(mai_mai_n633_), .Y(mai_mai_n646_));
  NA4        m624(.A(mai_mai_n646_), .B(mai_mai_n630_), .C(mai_mai_n624_), .D(mai_mai_n599_), .Y(mai_mai_n647_));
  NA2        m625(.A(mai_mai_n350_), .B(mai_mai_n349_), .Y(mai_mai_n648_));
  INV        m626(.A(mai_mai_n648_), .Y(mai_mai_n649_));
  NA2        m627(.A(mai_mai_n649_), .B(i_1_), .Y(mai_mai_n650_));
  AOI210     m628(.A0(mai_mai_n250_), .A1(mai_mai_n96_), .B0(i_1_), .Y(mai_mai_n651_));
  NO2        m629(.A(mai_mai_n348_), .B(i_2_), .Y(mai_mai_n652_));
  NA2        m630(.A(mai_mai_n652_), .B(mai_mai_n651_), .Y(mai_mai_n653_));
  OAI210     m631(.A0(mai_mai_n614_), .A1(mai_mai_n418_), .B0(mai_mai_n653_), .Y(mai_mai_n654_));
  INV        m632(.A(mai_mai_n654_), .Y(mai_mai_n655_));
  AOI210     m633(.A0(mai_mai_n655_), .A1(mai_mai_n650_), .B0(i_13_), .Y(mai_mai_n656_));
  OR2        m634(.A(i_11_), .B(i_7_), .Y(mai_mai_n657_));
  NA3        m635(.A(mai_mai_n657_), .B(mai_mai_n105_), .C(mai_mai_n132_), .Y(mai_mai_n658_));
  AOI220     m636(.A0(mai_mai_n438_), .A1(mai_mai_n155_), .B0(i_2_), .B1(mai_mai_n132_), .Y(mai_mai_n659_));
  OAI210     m637(.A0(mai_mai_n659_), .A1(mai_mai_n45_), .B0(mai_mai_n658_), .Y(mai_mai_n660_));
  NO2        m638(.A(mai_mai_n52_), .B(i_12_), .Y(mai_mai_n661_));
  INV        m639(.A(mai_mai_n661_), .Y(mai_mai_n662_));
  NO2        m640(.A(mai_mai_n444_), .B(mai_mai_n24_), .Y(mai_mai_n663_));
  AOI220     m641(.A0(mai_mai_n663_), .A1(mai_mai_n629_), .B0(mai_mai_n236_), .B1(mai_mai_n126_), .Y(mai_mai_n664_));
  OAI220     m642(.A0(mai_mai_n664_), .A1(mai_mai_n41_), .B0(mai_mai_n662_), .B1(mai_mai_n92_), .Y(mai_mai_n665_));
  AOI210     m643(.A0(mai_mai_n660_), .A1(mai_mai_n310_), .B0(mai_mai_n665_), .Y(mai_mai_n666_));
  INV        m644(.A(mai_mai_n113_), .Y(mai_mai_n667_));
  AOI220     m645(.A0(mai_mai_n667_), .A1(mai_mai_n69_), .B0(mai_mai_n361_), .B1(mai_mai_n611_), .Y(mai_mai_n668_));
  NO2        m646(.A(mai_mai_n668_), .B(mai_mai_n233_), .Y(mai_mai_n669_));
  AOI210     m647(.A0(mai_mai_n418_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n670_));
  NOi31      m648(.An(mai_mai_n670_), .B(mai_mai_n562_), .C(mai_mai_n45_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n122_), .B(i_13_), .Y(mai_mai_n672_));
  NO2        m650(.A(mai_mai_n610_), .B(mai_mai_n113_), .Y(mai_mai_n673_));
  INV        m651(.A(mai_mai_n673_), .Y(mai_mai_n674_));
  OAI220     m652(.A0(mai_mai_n674_), .A1(mai_mai_n68_), .B0(mai_mai_n672_), .B1(mai_mai_n651_), .Y(mai_mai_n675_));
  NO3        m653(.A(mai_mai_n68_), .B(mai_mai_n32_), .C(mai_mai_n100_), .Y(mai_mai_n676_));
  NA2        m654(.A(mai_mai_n26_), .B(mai_mai_n188_), .Y(mai_mai_n677_));
  NA2        m655(.A(mai_mai_n677_), .B(i_7_), .Y(mai_mai_n678_));
  NO3        m656(.A(mai_mai_n444_), .B(mai_mai_n227_), .C(mai_mai_n83_), .Y(mai_mai_n679_));
  AOI210     m657(.A0(mai_mai_n679_), .A1(mai_mai_n678_), .B0(mai_mai_n676_), .Y(mai_mai_n680_));
  NA2        m658(.A(mai_mai_n91_), .B(mai_mai_n101_), .Y(mai_mai_n681_));
  OAI220     m659(.A0(mai_mai_n681_), .A1(mai_mai_n568_), .B0(mai_mai_n680_), .B1(mai_mai_n581_), .Y(mai_mai_n682_));
  NO4        m660(.A(mai_mai_n682_), .B(mai_mai_n675_), .C(mai_mai_n671_), .D(mai_mai_n669_), .Y(mai_mai_n683_));
  OR2        m661(.A(i_11_), .B(i_6_), .Y(mai_mai_n684_));
  NA3        m662(.A(mai_mai_n567_), .B(mai_mai_n677_), .C(i_7_), .Y(mai_mai_n685_));
  AOI210     m663(.A0(mai_mai_n685_), .A1(mai_mai_n674_), .B0(mai_mai_n684_), .Y(mai_mai_n686_));
  NA3        m664(.A(mai_mai_n381_), .B(mai_mai_n572_), .C(mai_mai_n96_), .Y(mai_mai_n687_));
  NA2        m665(.A(mai_mai_n602_), .B(i_13_), .Y(mai_mai_n688_));
  NA2        m666(.A(mai_mai_n101_), .B(mai_mai_n677_), .Y(mai_mai_n689_));
  NAi21      m667(.An(i_11_), .B(i_12_), .Y(mai_mai_n690_));
  NOi41      m668(.An(mai_mai_n110_), .B(mai_mai_n690_), .C(i_13_), .D(mai_mai_n83_), .Y(mai_mai_n691_));
  NO3        m669(.A(mai_mai_n444_), .B(mai_mai_n545_), .C(mai_mai_n573_), .Y(mai_mai_n692_));
  AOI220     m670(.A0(mai_mai_n692_), .A1(mai_mai_n290_), .B0(mai_mai_n691_), .B1(mai_mai_n689_), .Y(mai_mai_n693_));
  NA3        m671(.A(mai_mai_n693_), .B(mai_mai_n688_), .C(mai_mai_n687_), .Y(mai_mai_n694_));
  OAI210     m672(.A0(mai_mai_n694_), .A1(mai_mai_n686_), .B0(mai_mai_n60_), .Y(mai_mai_n695_));
  NO2        m673(.A(i_2_), .B(i_12_), .Y(mai_mai_n696_));
  NA2        m674(.A(mai_mai_n347_), .B(mai_mai_n696_), .Y(mai_mai_n697_));
  NO3        m675(.A(i_9_), .B(i_3_), .C(mai_mai_n567_), .Y(mai_mai_n698_));
  NA2        m676(.A(mai_mai_n698_), .B(mai_mai_n347_), .Y(mai_mai_n699_));
  NO2        m677(.A(mai_mai_n123_), .B(i_2_), .Y(mai_mai_n700_));
  NA2        m678(.A(mai_mai_n700_), .B(mai_mai_n595_), .Y(mai_mai_n701_));
  NA3        m679(.A(mai_mai_n701_), .B(mai_mai_n699_), .C(mai_mai_n697_), .Y(mai_mai_n702_));
  NA3        m680(.A(mai_mai_n702_), .B(mai_mai_n46_), .C(mai_mai_n218_), .Y(mai_mai_n703_));
  NA4        m681(.A(mai_mai_n703_), .B(mai_mai_n695_), .C(mai_mai_n683_), .D(mai_mai_n666_), .Y(mai_mai_n704_));
  OR4        m682(.A(mai_mai_n704_), .B(mai_mai_n656_), .C(mai_mai_n647_), .D(mai_mai_n584_), .Y(mai5));
  NA2        m683(.A(mai_mai_n626_), .B(mai_mai_n252_), .Y(mai_mai_n706_));
  AN2        m684(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n707_));
  NA3        m685(.A(mai_mai_n707_), .B(mai_mai_n696_), .C(mai_mai_n107_), .Y(mai_mai_n708_));
  NO2        m686(.A(mai_mai_n568_), .B(i_11_), .Y(mai_mai_n709_));
  NA2        m687(.A(mai_mai_n86_), .B(mai_mai_n709_), .Y(mai_mai_n710_));
  NA3        m688(.A(mai_mai_n710_), .B(mai_mai_n708_), .C(mai_mai_n706_), .Y(mai_mai_n711_));
  NO3        m689(.A(i_11_), .B(mai_mai_n227_), .C(i_13_), .Y(mai_mai_n712_));
  NO2        m690(.A(mai_mai_n119_), .B(mai_mai_n23_), .Y(mai_mai_n713_));
  NA2        m691(.A(i_12_), .B(i_8_), .Y(mai_mai_n714_));
  OAI210     m692(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n714_), .Y(mai_mai_n715_));
  INV        m693(.A(mai_mai_n417_), .Y(mai_mai_n716_));
  AOI220     m694(.A0(mai_mai_n296_), .A1(mai_mai_n538_), .B0(mai_mai_n715_), .B1(mai_mai_n713_), .Y(mai_mai_n717_));
  INV        m695(.A(mai_mai_n717_), .Y(mai_mai_n718_));
  NO2        m696(.A(mai_mai_n718_), .B(mai_mai_n711_), .Y(mai_mai_n719_));
  INV        m697(.A(mai_mai_n166_), .Y(mai_mai_n720_));
  INV        m698(.A(mai_mai_n236_), .Y(mai_mai_n721_));
  OAI210     m699(.A0(mai_mai_n652_), .A1(mai_mai_n419_), .B0(mai_mai_n110_), .Y(mai_mai_n722_));
  AOI210     m700(.A0(mai_mai_n722_), .A1(mai_mai_n721_), .B0(mai_mai_n720_), .Y(mai_mai_n723_));
  NO2        m701(.A(mai_mai_n424_), .B(mai_mai_n26_), .Y(mai_mai_n724_));
  NO2        m702(.A(mai_mai_n724_), .B(mai_mai_n391_), .Y(mai_mai_n725_));
  NA2        m703(.A(mai_mai_n725_), .B(i_2_), .Y(mai_mai_n726_));
  INV        m704(.A(mai_mai_n726_), .Y(mai_mai_n727_));
  AOI210     m705(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n388_), .Y(mai_mai_n728_));
  AOI210     m706(.A0(mai_mai_n728_), .A1(mai_mai_n727_), .B0(mai_mai_n723_), .Y(mai_mai_n729_));
  NO2        m707(.A(mai_mai_n185_), .B(mai_mai_n120_), .Y(mai_mai_n730_));
  OAI210     m708(.A0(mai_mai_n730_), .A1(mai_mai_n713_), .B0(i_2_), .Y(mai_mai_n731_));
  INV        m709(.A(mai_mai_n167_), .Y(mai_mai_n732_));
  NO3        m710(.A(mai_mai_n586_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n733_));
  AOI210     m711(.A0(mai_mai_n732_), .A1(mai_mai_n86_), .B0(mai_mai_n733_), .Y(mai_mai_n734_));
  AOI210     m712(.A0(mai_mai_n734_), .A1(mai_mai_n731_), .B0(mai_mai_n188_), .Y(mai_mai_n735_));
  OA210      m713(.A0(mai_mai_n587_), .A1(mai_mai_n121_), .B0(i_13_), .Y(mai_mai_n736_));
  NA2        m714(.A(mai_mai_n195_), .B(mai_mai_n198_), .Y(mai_mai_n737_));
  NA2        m715(.A(mai_mai_n145_), .B(mai_mai_n563_), .Y(mai_mai_n738_));
  AOI210     m716(.A0(mai_mai_n738_), .A1(mai_mai_n737_), .B0(mai_mai_n351_), .Y(mai_mai_n739_));
  AOI210     m717(.A0(mai_mai_n203_), .A1(mai_mai_n142_), .B0(mai_mai_n485_), .Y(mai_mai_n740_));
  NA2        m718(.A(mai_mai_n740_), .B(mai_mai_n391_), .Y(mai_mai_n741_));
  NO2        m719(.A(mai_mai_n101_), .B(mai_mai_n45_), .Y(mai_mai_n742_));
  INV        m720(.A(mai_mai_n279_), .Y(mai_mai_n743_));
  NA4        m721(.A(mai_mai_n743_), .B(mai_mai_n283_), .C(mai_mai_n119_), .D(mai_mai_n43_), .Y(mai_mai_n744_));
  OAI210     m722(.A0(mai_mai_n744_), .A1(mai_mai_n742_), .B0(mai_mai_n741_), .Y(mai_mai_n745_));
  NO4        m723(.A(mai_mai_n745_), .B(mai_mai_n739_), .C(mai_mai_n736_), .D(mai_mai_n735_), .Y(mai_mai_n746_));
  NA2        m724(.A(mai_mai_n538_), .B(mai_mai_n28_), .Y(mai_mai_n747_));
  NA2        m725(.A(mai_mai_n712_), .B(mai_mai_n256_), .Y(mai_mai_n748_));
  NA2        m726(.A(mai_mai_n748_), .B(mai_mai_n747_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n59_), .B(i_12_), .Y(mai_mai_n750_));
  NO2        m728(.A(mai_mai_n750_), .B(mai_mai_n121_), .Y(mai_mai_n751_));
  NO2        m729(.A(mai_mai_n751_), .B(mai_mai_n563_), .Y(mai_mai_n752_));
  AOI220     m730(.A0(mai_mai_n752_), .A1(mai_mai_n36_), .B0(mai_mai_n749_), .B1(mai_mai_n47_), .Y(mai_mai_n753_));
  NA4        m731(.A(mai_mai_n753_), .B(mai_mai_n746_), .C(mai_mai_n729_), .D(mai_mai_n719_), .Y(mai6));
  NO3        m732(.A(mai_mai_n246_), .B(mai_mai_n285_), .C(i_1_), .Y(mai_mai_n755_));
  NO2        m733(.A(mai_mai_n180_), .B(mai_mai_n133_), .Y(mai_mai_n756_));
  OAI210     m734(.A0(mai_mai_n756_), .A1(mai_mai_n755_), .B0(mai_mai_n700_), .Y(mai_mai_n757_));
  NA4        m735(.A(mai_mai_n363_), .B(mai_mai_n449_), .C(mai_mai_n68_), .D(mai_mai_n100_), .Y(mai_mai_n758_));
  INV        m736(.A(mai_mai_n758_), .Y(mai_mai_n759_));
  NO2        m737(.A(mai_mai_n214_), .B(mai_mai_n454_), .Y(mai_mai_n760_));
  NO2        m738(.A(i_11_), .B(i_9_), .Y(mai_mai_n761_));
  NO2        m739(.A(mai_mai_n759_), .B(mai_mai_n308_), .Y(mai_mai_n762_));
  AO210      m740(.A0(mai_mai_n762_), .A1(mai_mai_n757_), .B0(i_12_), .Y(mai_mai_n763_));
  NA2        m741(.A(mai_mai_n352_), .B(mai_mai_n313_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n545_), .B(mai_mai_n60_), .Y(mai_mai_n765_));
  BUFFER     m743(.A(mai_mai_n591_), .Y(mai_mai_n766_));
  NA3        m744(.A(mai_mai_n766_), .B(mai_mai_n765_), .C(mai_mai_n764_), .Y(mai_mai_n767_));
  INV        m745(.A(mai_mai_n192_), .Y(mai_mai_n768_));
  AOI220     m746(.A0(mai_mai_n768_), .A1(mai_mai_n761_), .B0(mai_mai_n767_), .B1(mai_mai_n70_), .Y(mai_mai_n769_));
  INV        m747(.A(mai_mai_n307_), .Y(mai_mai_n770_));
  NA2        m748(.A(mai_mai_n72_), .B(mai_mai_n126_), .Y(mai_mai_n771_));
  INV        m749(.A(mai_mai_n119_), .Y(mai_mai_n772_));
  NA2        m750(.A(mai_mai_n772_), .B(mai_mai_n47_), .Y(mai_mai_n773_));
  AOI210     m751(.A0(mai_mai_n773_), .A1(mai_mai_n771_), .B0(mai_mai_n770_), .Y(mai_mai_n774_));
  NO2        m752(.A(mai_mai_n243_), .B(i_9_), .Y(mai_mai_n775_));
  NA2        m753(.A(mai_mai_n775_), .B(mai_mai_n750_), .Y(mai_mai_n776_));
  AOI210     m754(.A0(mai_mai_n776_), .A1(mai_mai_n483_), .B0(mai_mai_n180_), .Y(mai_mai_n777_));
  NAi32      m755(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n778_));
  NO2        m756(.A(mai_mai_n684_), .B(mai_mai_n778_), .Y(mai_mai_n779_));
  OR3        m757(.A(mai_mai_n779_), .B(mai_mai_n777_), .C(mai_mai_n774_), .Y(mai_mai_n780_));
  NO2        m758(.A(mai_mai_n657_), .B(i_2_), .Y(mai_mai_n781_));
  NA2        m759(.A(mai_mai_n48_), .B(mai_mai_n37_), .Y(mai_mai_n782_));
  NO2        m760(.A(mai_mai_n782_), .B(mai_mai_n380_), .Y(mai_mai_n783_));
  NA2        m761(.A(mai_mai_n783_), .B(mai_mai_n781_), .Y(mai_mai_n784_));
  OR2        m762(.A(mai_mai_n587_), .B(mai_mai_n419_), .Y(mai_mai_n785_));
  NA3        m763(.A(mai_mai_n785_), .B(mai_mai_n141_), .C(mai_mai_n66_), .Y(mai_mai_n786_));
  OR2        m764(.A(mai_mai_n716_), .B(mai_mai_n36_), .Y(mai_mai_n787_));
  NA3        m765(.A(mai_mai_n787_), .B(mai_mai_n786_), .C(mai_mai_n784_), .Y(mai_mai_n788_));
  OAI210     m766(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n84_), .Y(mai_mai_n789_));
  AOI220     m767(.A0(mai_mai_n789_), .A1(mai_mai_n529_), .B0(mai_mai_n760_), .B1(mai_mai_n678_), .Y(mai_mai_n790_));
  NA2        m768(.A(mai_mai_n369_), .B(mai_mai_n67_), .Y(mai_mai_n791_));
  NA3        m769(.A(mai_mai_n791_), .B(mai_mai_n790_), .C(mai_mai_n571_), .Y(mai_mai_n792_));
  BUFFER     m770(.A(mai_mai_n85_), .Y(mai_mai_n793_));
  NA3        m771(.A(mai_mai_n793_), .B(mai_mai_n450_), .C(mai_mai_n213_), .Y(mai_mai_n794_));
  AOI210     m772(.A0(mai_mai_n419_), .A1(mai_mai_n417_), .B0(mai_mai_n528_), .Y(mai_mai_n795_));
  NO2        m773(.A(mai_mai_n577_), .B(mai_mai_n101_), .Y(mai_mai_n796_));
  OAI210     m774(.A0(mai_mai_n796_), .A1(mai_mai_n111_), .B0(mai_mai_n379_), .Y(mai_mai_n797_));
  INV        m775(.A(mai_mai_n552_), .Y(mai_mai_n798_));
  NA3        m776(.A(mai_mai_n798_), .B(mai_mai_n307_), .C(i_7_), .Y(mai_mai_n799_));
  NA4        m777(.A(mai_mai_n799_), .B(mai_mai_n797_), .C(mai_mai_n795_), .D(mai_mai_n794_), .Y(mai_mai_n800_));
  NO4        m778(.A(mai_mai_n800_), .B(mai_mai_n792_), .C(mai_mai_n788_), .D(mai_mai_n780_), .Y(mai_mai_n801_));
  NA4        m779(.A(mai_mai_n801_), .B(mai_mai_n769_), .C(mai_mai_n763_), .D(mai_mai_n357_), .Y(mai3));
  NA2        m780(.A(i_6_), .B(i_7_), .Y(mai_mai_n803_));
  NO2        m781(.A(mai_mai_n803_), .B(i_0_), .Y(mai_mai_n804_));
  NO2        m782(.A(i_11_), .B(mai_mai_n227_), .Y(mai_mai_n805_));
  OAI210     m783(.A0(mai_mai_n804_), .A1(mai_mai_n270_), .B0(mai_mai_n805_), .Y(mai_mai_n806_));
  NO2        m784(.A(mai_mai_n806_), .B(mai_mai_n188_), .Y(mai_mai_n807_));
  NO3        m785(.A(mai_mai_n420_), .B(mai_mai_n89_), .C(mai_mai_n45_), .Y(mai_mai_n808_));
  OA210      m786(.A0(mai_mai_n808_), .A1(mai_mai_n807_), .B0(mai_mai_n168_), .Y(mai_mai_n809_));
  NA2        m787(.A(mai_mai_n381_), .B(mai_mai_n46_), .Y(mai_mai_n810_));
  AN2        m788(.A(mai_mai_n422_), .B(mai_mai_n53_), .Y(mai_mai_n811_));
  INV        m789(.A(mai_mai_n811_), .Y(mai_mai_n812_));
  NO2        m790(.A(mai_mai_n812_), .B(mai_mai_n48_), .Y(mai_mai_n813_));
  NO4        m791(.A(mai_mai_n353_), .B(mai_mai_n360_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n814_));
  NA2        m792(.A(mai_mai_n670_), .B(mai_mai_n638_), .Y(mai_mai_n815_));
  NA2        m793(.A(mai_mai_n311_), .B(i_5_), .Y(mai_mai_n816_));
  OAI220     m794(.A0(mai_mai_n816_), .A1(mai_mai_n815_), .B0(mai_mai_n988_), .B1(mai_mai_n60_), .Y(mai_mai_n817_));
  NOi21      m795(.An(i_5_), .B(i_9_), .Y(mai_mai_n818_));
  NA2        m796(.A(mai_mai_n818_), .B(mai_mai_n416_), .Y(mai_mai_n819_));
  BUFFER     m797(.A(mai_mai_n250_), .Y(mai_mai_n820_));
  NA2        m798(.A(mai_mai_n820_), .B(mai_mai_n442_), .Y(mai_mai_n821_));
  NO3        m799(.A(mai_mai_n384_), .B(mai_mai_n250_), .C(mai_mai_n70_), .Y(mai_mai_n822_));
  NO2        m800(.A(mai_mai_n169_), .B(mai_mai_n142_), .Y(mai_mai_n823_));
  AOI210     m801(.A0(mai_mai_n823_), .A1(mai_mai_n235_), .B0(mai_mai_n822_), .Y(mai_mai_n824_));
  OAI220     m802(.A0(mai_mai_n824_), .A1(mai_mai_n175_), .B0(mai_mai_n821_), .B1(mai_mai_n819_), .Y(mai_mai_n825_));
  NO4        m803(.A(mai_mai_n825_), .B(mai_mai_n817_), .C(mai_mai_n813_), .D(mai_mai_n809_), .Y(mai_mai_n826_));
  NA2        m804(.A(mai_mai_n180_), .B(mai_mai_n24_), .Y(mai_mai_n827_));
  NO2        m805(.A(mai_mai_n636_), .B(mai_mai_n560_), .Y(mai_mai_n828_));
  NO2        m806(.A(mai_mai_n828_), .B(mai_mai_n827_), .Y(mai_mai_n829_));
  INV        m807(.A(mai_mai_n829_), .Y(mai_mai_n830_));
  NO2        m808(.A(mai_mai_n363_), .B(mai_mai_n271_), .Y(mai_mai_n831_));
  NA2        m809(.A(mai_mai_n831_), .B(mai_mai_n673_), .Y(mai_mai_n832_));
  NO4        m810(.A(mai_mai_n551_), .B(mai_mai_n211_), .C(mai_mai_n388_), .D(mai_mai_n380_), .Y(mai_mai_n833_));
  NA2        m811(.A(mai_mai_n833_), .B(i_11_), .Y(mai_mai_n834_));
  AN2        m812(.A(mai_mai_n95_), .B(mai_mai_n234_), .Y(mai_mai_n835_));
  NA2        m813(.A(mai_mai_n712_), .B(mai_mai_n308_), .Y(mai_mai_n836_));
  AOI210     m814(.A0(mai_mai_n450_), .A1(mai_mai_n86_), .B0(mai_mai_n55_), .Y(mai_mai_n837_));
  OAI220     m815(.A0(mai_mai_n837_), .A1(mai_mai_n836_), .B0(mai_mai_n621_), .B1(mai_mai_n504_), .Y(mai_mai_n838_));
  NO2        m816(.A(mai_mai_n245_), .B(mai_mai_n147_), .Y(mai_mai_n839_));
  INV        m817(.A(mai_mai_n507_), .Y(mai_mai_n840_));
  NO4        m818(.A(mai_mai_n113_), .B(mai_mai_n55_), .C(mai_mai_n631_), .D(i_5_), .Y(mai_mai_n841_));
  AO220      m819(.A0(mai_mai_n841_), .A1(mai_mai_n840_), .B0(mai_mai_n839_), .B1(i_6_), .Y(mai_mai_n842_));
  AOI220     m820(.A0(mai_mai_n311_), .A1(mai_mai_n97_), .B0(mai_mai_n180_), .B1(mai_mai_n81_), .Y(mai_mai_n843_));
  NA2        m821(.A(mai_mai_n533_), .B(i_4_), .Y(mai_mai_n844_));
  INV        m822(.A(mai_mai_n183_), .Y(mai_mai_n845_));
  OAI220     m823(.A0(mai_mai_n845_), .A1(mai_mai_n836_), .B0(mai_mai_n844_), .B1(mai_mai_n843_), .Y(mai_mai_n846_));
  NO4        m824(.A(mai_mai_n846_), .B(mai_mai_n842_), .C(mai_mai_n838_), .D(mai_mai_n835_), .Y(mai_mai_n847_));
  NA4        m825(.A(mai_mai_n847_), .B(mai_mai_n834_), .C(mai_mai_n832_), .D(mai_mai_n830_), .Y(mai_mai_n848_));
  NA2        m826(.A(i_11_), .B(i_9_), .Y(mai_mai_n849_));
  NO2        m827(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n850_));
  NA2        m828(.A(mai_mai_n368_), .B(mai_mai_n173_), .Y(mai_mai_n851_));
  NA2        m829(.A(mai_mai_n851_), .B(mai_mai_n154_), .Y(mai_mai_n852_));
  NO2        m830(.A(mai_mai_n849_), .B(mai_mai_n70_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n169_), .B(i_0_), .Y(mai_mai_n854_));
  INV        m832(.A(mai_mai_n854_), .Y(mai_mai_n855_));
  NA2        m833(.A(mai_mai_n440_), .B(mai_mai_n221_), .Y(mai_mai_n856_));
  AOI210     m834(.A0(mai_mai_n350_), .A1(mai_mai_n42_), .B0(mai_mai_n378_), .Y(mai_mai_n857_));
  OAI220     m835(.A0(mai_mai_n857_), .A1(mai_mai_n819_), .B0(mai_mai_n856_), .B1(mai_mai_n855_), .Y(mai_mai_n858_));
  NO2        m836(.A(mai_mai_n858_), .B(mai_mai_n852_), .Y(mai_mai_n859_));
  NA2        m837(.A(mai_mai_n620_), .B(mai_mai_n116_), .Y(mai_mai_n860_));
  NO2        m838(.A(i_6_), .B(mai_mai_n860_), .Y(mai_mai_n861_));
  AOI210     m839(.A0(mai_mai_n418_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n862_));
  NA2        m840(.A(mai_mai_n166_), .B(mai_mai_n102_), .Y(mai_mai_n863_));
  NOi32      m841(.An(mai_mai_n862_), .Bn(mai_mai_n183_), .C(mai_mai_n863_), .Y(mai_mai_n864_));
  NA2        m842(.A(mai_mai_n572_), .B(mai_mai_n308_), .Y(mai_mai_n865_));
  NO2        m843(.A(mai_mai_n865_), .B(mai_mai_n810_), .Y(mai_mai_n866_));
  NO3        m844(.A(mai_mai_n866_), .B(mai_mai_n864_), .C(mai_mai_n861_), .Y(mai_mai_n867_));
  NOi21      m845(.An(i_7_), .B(i_5_), .Y(mai_mai_n868_));
  OR2        m846(.A(mai_mai_n863_), .B(mai_mai_n483_), .Y(mai_mai_n869_));
  NO3        m847(.A(mai_mai_n374_), .B(mai_mai_n339_), .C(mai_mai_n338_), .Y(mai_mai_n870_));
  NO2        m848(.A(mai_mai_n248_), .B(mai_mai_n297_), .Y(mai_mai_n871_));
  INV        m849(.A(mai_mai_n690_), .Y(mai_mai_n872_));
  AOI210     m850(.A0(mai_mai_n872_), .A1(mai_mai_n871_), .B0(mai_mai_n870_), .Y(mai_mai_n873_));
  NA4        m851(.A(mai_mai_n873_), .B(mai_mai_n869_), .C(mai_mai_n867_), .D(mai_mai_n859_), .Y(mai_mai_n874_));
  AN2        m852(.A(mai_mai_n310_), .B(mai_mai_n308_), .Y(mai_mai_n875_));
  AN2        m853(.A(mai_mai_n875_), .B(mai_mai_n823_), .Y(mai_mai_n876_));
  INV        m854(.A(mai_mai_n876_), .Y(mai_mai_n877_));
  OA210      m855(.A0(mai_mai_n440_), .A1(mai_mai_n217_), .B0(mai_mai_n439_), .Y(mai_mai_n878_));
  NA2        m856(.A(mai_mai_n853_), .B(mai_mai_n283_), .Y(mai_mai_n879_));
  OAI210     m857(.A0(i_2_), .A1(mai_mai_n182_), .B0(mai_mai_n879_), .Y(mai_mai_n880_));
  NA2        m858(.A(mai_mai_n880_), .B(mai_mai_n440_), .Y(mai_mai_n881_));
  NAi21      m859(.An(i_9_), .B(i_5_), .Y(mai_mai_n882_));
  NO2        m860(.A(mai_mai_n882_), .B(mai_mai_n374_), .Y(mai_mai_n883_));
  NO2        m861(.A(mai_mai_n566_), .B(mai_mai_n104_), .Y(mai_mai_n884_));
  AOI220     m862(.A0(mai_mai_n884_), .A1(i_0_), .B0(mai_mai_n883_), .B1(mai_mai_n587_), .Y(mai_mai_n885_));
  NO2        m863(.A(mai_mai_n885_), .B(mai_mai_n83_), .Y(mai_mai_n886_));
  NO2        m864(.A(mai_mai_n886_), .B(mai_mai_n488_), .Y(mai_mai_n887_));
  NA3        m865(.A(mai_mai_n887_), .B(mai_mai_n881_), .C(mai_mai_n877_), .Y(mai_mai_n888_));
  NO3        m866(.A(mai_mai_n888_), .B(mai_mai_n874_), .C(mai_mai_n848_), .Y(mai_mai_n889_));
  NO2        m867(.A(i_0_), .B(mai_mai_n690_), .Y(mai_mai_n890_));
  NA2        m868(.A(mai_mai_n70_), .B(mai_mai_n45_), .Y(mai_mai_n891_));
  INV        m869(.A(mai_mai_n891_), .Y(mai_mai_n892_));
  NO3        m870(.A(mai_mai_n104_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n893_));
  AO220      m871(.A0(mai_mai_n893_), .A1(mai_mai_n892_), .B0(mai_mai_n890_), .B1(mai_mai_n168_), .Y(mai_mai_n894_));
  AOI210     m872(.A0(mai_mai_n765_), .A1(mai_mai_n648_), .B0(mai_mai_n863_), .Y(mai_mai_n895_));
  AOI210     m873(.A0(mai_mai_n894_), .A1(mai_mai_n327_), .B0(mai_mai_n895_), .Y(mai_mai_n896_));
  NA2        m874(.A(mai_mai_n700_), .B(mai_mai_n140_), .Y(mai_mai_n897_));
  INV        m875(.A(mai_mai_n897_), .Y(mai_mai_n898_));
  NA3        m876(.A(mai_mai_n898_), .B(mai_mai_n638_), .C(mai_mai_n70_), .Y(mai_mai_n899_));
  NA3        m877(.A(mai_mai_n804_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n900_));
  NA2        m878(.A(mai_mai_n805_), .B(i_9_), .Y(mai_mai_n901_));
  AOI210     m879(.A0(mai_mai_n900_), .A1(mai_mai_n464_), .B0(mai_mai_n901_), .Y(mai_mai_n902_));
  NA2        m880(.A(mai_mai_n235_), .B(mai_mai_n220_), .Y(mai_mai_n903_));
  NO2        m881(.A(mai_mai_n903_), .B(mai_mai_n147_), .Y(mai_mai_n904_));
  NO2        m882(.A(mai_mai_n904_), .B(mai_mai_n902_), .Y(mai_mai_n905_));
  NA3        m883(.A(mai_mai_n905_), .B(mai_mai_n899_), .C(mai_mai_n896_), .Y(mai_mai_n906_));
  NA2        m884(.A(mai_mai_n875_), .B(mai_mai_n351_), .Y(mai_mai_n907_));
  AOI210     m885(.A0(mai_mai_n278_), .A1(mai_mai_n156_), .B0(mai_mai_n907_), .Y(mai_mai_n908_));
  NA3        m886(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n909_));
  NA2        m887(.A(mai_mai_n850_), .B(mai_mai_n455_), .Y(mai_mai_n910_));
  AOI210     m888(.A0(mai_mai_n909_), .A1(mai_mai_n156_), .B0(mai_mai_n910_), .Y(mai_mai_n911_));
  NO2        m889(.A(mai_mai_n911_), .B(mai_mai_n908_), .Y(mai_mai_n912_));
  NA2        m890(.A(mai_mai_n534_), .B(mai_mai_n72_), .Y(mai_mai_n913_));
  NO3        m891(.A(mai_mai_n205_), .B(mai_mai_n360_), .C(i_0_), .Y(mai_mai_n914_));
  OAI210     m892(.A0(mai_mai_n914_), .A1(mai_mai_n73_), .B0(i_13_), .Y(mai_mai_n915_));
  INV        m893(.A(mai_mai_n213_), .Y(mai_mai_n916_));
  OAI220     m894(.A0(mai_mai_n498_), .A1(mai_mai_n133_), .B0(i_12_), .B1(mai_mai_n581_), .Y(mai_mai_n917_));
  NA3        m895(.A(mai_mai_n917_), .B(mai_mai_n370_), .C(mai_mai_n916_), .Y(mai_mai_n918_));
  NA4        m896(.A(mai_mai_n918_), .B(mai_mai_n915_), .C(mai_mai_n913_), .D(mai_mai_n912_), .Y(mai_mai_n919_));
  INV        m897(.A(mai_mai_n108_), .Y(mai_mai_n920_));
  AOI220     m898(.A0(mai_mai_n868_), .A1(mai_mai_n455_), .B0(mai_mai_n804_), .B1(mai_mai_n157_), .Y(mai_mai_n921_));
  NA2        m899(.A(mai_mai_n330_), .B(mai_mai_n170_), .Y(mai_mai_n922_));
  OA220      m900(.A0(mai_mai_n922_), .A1(mai_mai_n921_), .B0(mai_mai_n920_), .B1(i_5_), .Y(mai_mai_n923_));
  AOI210     m901(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n169_), .Y(mai_mai_n924_));
  NA2        m902(.A(mai_mai_n924_), .B(mai_mai_n878_), .Y(mai_mai_n925_));
  NA3        m903(.A(mai_mai_n578_), .B(mai_mai_n180_), .C(mai_mai_n81_), .Y(mai_mai_n926_));
  INV        m904(.A(mai_mai_n926_), .Y(mai_mai_n927_));
  NO3        m905(.A(mai_mai_n810_), .B(mai_mai_n52_), .C(mai_mai_n48_), .Y(mai_mai_n928_));
  NA2        m906(.A(mai_mai_n460_), .B(mai_mai_n453_), .Y(mai_mai_n929_));
  NO3        m907(.A(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n927_), .Y(mai_mai_n930_));
  NA3        m908(.A(mai_mai_n363_), .B(mai_mai_n166_), .C(mai_mai_n165_), .Y(mai_mai_n931_));
  NA3        m909(.A(mai_mai_n850_), .B(mai_mai_n270_), .C(mai_mai_n220_), .Y(mai_mai_n932_));
  NA2        m910(.A(mai_mai_n932_), .B(mai_mai_n931_), .Y(mai_mai_n933_));
  NOi31      m911(.An(mai_mai_n362_), .B(mai_mai_n891_), .C(mai_mai_n230_), .Y(mai_mai_n934_));
  NO3        m912(.A(mai_mai_n849_), .B(mai_mai_n213_), .C(mai_mai_n185_), .Y(mai_mai_n935_));
  NO3        m913(.A(mai_mai_n935_), .B(mai_mai_n934_), .C(mai_mai_n933_), .Y(mai_mai_n936_));
  NA4        m914(.A(mai_mai_n936_), .B(mai_mai_n930_), .C(mai_mai_n925_), .D(mai_mai_n923_), .Y(mai_mai_n937_));
  INV        m915(.A(mai_mai_n580_), .Y(mai_mai_n938_));
  NO3        m916(.A(mai_mai_n938_), .B(mai_mai_n524_), .C(mai_mai_n324_), .Y(mai_mai_n939_));
  INV        m917(.A(mai_mai_n939_), .Y(mai_mai_n940_));
  NA2        m918(.A(mai_mai_n759_), .B(mai_mai_n170_), .Y(mai_mai_n941_));
  NA3        m919(.A(mai_mai_n97_), .B(i_10_), .C(i_11_), .Y(mai_mai_n942_));
  NO2        m920(.A(mai_mai_n942_), .B(mai_mai_n149_), .Y(mai_mai_n943_));
  NA2        m921(.A(mai_mai_n868_), .B(mai_mai_n438_), .Y(mai_mai_n944_));
  NO2        m922(.A(mai_mai_n944_), .B(mai_mai_n639_), .Y(mai_mai_n945_));
  AOI210     m923(.A0(mai_mai_n945_), .A1(mai_mai_n854_), .B0(mai_mai_n943_), .Y(mai_mai_n946_));
  NA3        m924(.A(mai_mai_n946_), .B(mai_mai_n941_), .C(mai_mai_n940_), .Y(mai_mai_n947_));
  NO4        m925(.A(mai_mai_n947_), .B(mai_mai_n937_), .C(mai_mai_n919_), .D(mai_mai_n906_), .Y(mai_mai_n948_));
  NA2        m926(.A(mai_mai_n781_), .B(mai_mai_n37_), .Y(mai_mai_n949_));
  NA3        m927(.A(mai_mai_n862_), .B(mai_mai_n347_), .C(i_5_), .Y(mai_mai_n950_));
  NA3        m928(.A(mai_mai_n950_), .B(mai_mai_n949_), .C(mai_mai_n576_), .Y(mai_mai_n951_));
  NA2        m929(.A(mai_mai_n951_), .B(mai_mai_n201_), .Y(mai_mai_n952_));
  AN2        m930(.A(mai_mai_n657_), .B(mai_mai_n348_), .Y(mai_mai_n953_));
  NA2        m931(.A(mai_mai_n181_), .B(mai_mai_n183_), .Y(mai_mai_n954_));
  AO210      m932(.A0(mai_mai_n953_), .A1(mai_mai_n33_), .B0(mai_mai_n954_), .Y(mai_mai_n955_));
  OAI210     m933(.A0(mai_mai_n580_), .A1(mai_mai_n578_), .B0(mai_mai_n296_), .Y(mai_mai_n956_));
  NAi31      m934(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n957_));
  NO2        m935(.A(mai_mai_n67_), .B(mai_mai_n957_), .Y(mai_mai_n958_));
  INV        m936(.A(mai_mai_n958_), .Y(mai_mai_n959_));
  NA3        m937(.A(mai_mai_n959_), .B(mai_mai_n956_), .C(mai_mai_n955_), .Y(mai_mai_n960_));
  NO2        m938(.A(mai_mai_n430_), .B(mai_mai_n250_), .Y(mai_mai_n961_));
  NO4        m939(.A(mai_mai_n223_), .B(mai_mai_n139_), .C(mai_mai_n642_), .D(mai_mai_n37_), .Y(mai_mai_n962_));
  NO3        m940(.A(mai_mai_n962_), .B(mai_mai_n961_), .C(mai_mai_n833_), .Y(mai_mai_n963_));
  OAI210     m941(.A0(mai_mai_n942_), .A1(mai_mai_n142_), .B0(mai_mai_n963_), .Y(mai_mai_n964_));
  AOI210     m942(.A0(mai_mai_n960_), .A1(mai_mai_n48_), .B0(mai_mai_n964_), .Y(mai_mai_n965_));
  AOI210     m943(.A0(mai_mai_n965_), .A1(mai_mai_n952_), .B0(mai_mai_n70_), .Y(mai_mai_n966_));
  NO2        m944(.A(mai_mai_n531_), .B(mai_mai_n356_), .Y(mai_mai_n967_));
  NO2        m945(.A(mai_mai_n967_), .B(mai_mai_n720_), .Y(mai_mai_n968_));
  NA2        m946(.A(mai_mai_n248_), .B(mai_mai_n54_), .Y(mai_mai_n969_));
  AOI220     m947(.A0(mai_mai_n969_), .A1(mai_mai_n73_), .B0(mai_mai_n325_), .B1(mai_mai_n246_), .Y(mai_mai_n970_));
  NO2        m948(.A(mai_mai_n970_), .B(mai_mai_n227_), .Y(mai_mai_n971_));
  INV        m949(.A(mai_mai_n971_), .Y(mai_mai_n972_));
  NA2        m950(.A(mai_mai_n573_), .B(mai_mai_n211_), .Y(mai_mai_n973_));
  OAI210     m951(.A0(mai_mai_n973_), .A1(mai_mai_n862_), .B0(mai_mai_n201_), .Y(mai_mai_n974_));
  NA2        m952(.A(mai_mai_n158_), .B(i_5_), .Y(mai_mai_n975_));
  NO2        m953(.A(mai_mai_n974_), .B(mai_mai_n975_), .Y(mai_mai_n976_));
  NO4        m954(.A(mai_mai_n882_), .B(mai_mai_n443_), .C(mai_mai_n244_), .D(mai_mai_n243_), .Y(mai_mai_n977_));
  NO2        m955(.A(mai_mai_n977_), .B(mai_mai_n528_), .Y(mai_mai_n978_));
  INV        m956(.A(mai_mai_n340_), .Y(mai_mai_n979_));
  AOI210     m957(.A0(mai_mai_n979_), .A1(mai_mai_n978_), .B0(mai_mai_n41_), .Y(mai_mai_n980_));
  NO2        m958(.A(mai_mai_n980_), .B(mai_mai_n976_), .Y(mai_mai_n981_));
  OAI210     m959(.A0(mai_mai_n972_), .A1(i_4_), .B0(mai_mai_n981_), .Y(mai_mai_n982_));
  NO3        m960(.A(mai_mai_n982_), .B(mai_mai_n968_), .C(mai_mai_n966_), .Y(mai_mai_n983_));
  NA4        m961(.A(mai_mai_n983_), .B(mai_mai_n948_), .C(mai_mai_n889_), .D(mai_mai_n826_), .Y(mai4));
  INV        m962(.A(mai_mai_n237_), .Y(mai_mai_n987_));
  INV        m963(.A(mai_mai_n814_), .Y(mai_mai_n988_));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NAi31      u0019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n42_));
  INV        u0020(.A(men_men_n35_), .Y(men1));
  INV        u0021(.A(i_11_), .Y(men_men_n44_));
  NO2        u0022(.A(men_men_n44_), .B(i_6_), .Y(men_men_n45_));
  INV        u0023(.A(i_2_), .Y(men_men_n46_));
  NA2        u0024(.A(i_0_), .B(i_3_), .Y(men_men_n47_));
  INV        u0025(.A(i_5_), .Y(men_men_n48_));
  NO2        u0026(.A(i_7_), .B(i_10_), .Y(men_men_n49_));
  AOI210     u0027(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n49_), .Y(men_men_n50_));
  OAI210     u0028(.A0(men_men_n50_), .A1(i_3_), .B0(men_men_n48_), .Y(men_men_n51_));
  AOI210     u0029(.A0(men_men_n51_), .A1(men_men_n47_), .B0(men_men_n46_), .Y(men_men_n52_));
  NA2        u0030(.A(i_0_), .B(i_2_), .Y(men_men_n53_));
  NA2        u0031(.A(i_7_), .B(i_9_), .Y(men_men_n54_));
  NO2        u0032(.A(men_men_n54_), .B(men_men_n53_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n52_), .B(men_men_n45_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n50_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(i_3_), .B(i_9_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_7_), .Y(men_men_n83_));
  NO3        u0061(.A(men_men_n83_), .B(men_men_n82_), .C(men_men_n63_), .Y(men_men_n84_));
  INV        u0062(.A(i_6_), .Y(men_men_n85_));
  NO2        u0063(.A(i_2_), .B(i_7_), .Y(men_men_n86_));
  INV        u0064(.A(men_men_n86_), .Y(men_men_n87_));
  NA2        u0065(.A(men_men_n84_), .B(men_men_n87_), .Y(men_men_n88_));
  NAi21      u0066(.An(i_6_), .B(i_10_), .Y(men_men_n89_));
  NA2        u0067(.A(i_6_), .B(i_9_), .Y(men_men_n90_));
  AOI210     u0068(.A0(men_men_n90_), .A1(men_men_n89_), .B0(men_men_n63_), .Y(men_men_n91_));
  NA2        u0069(.A(i_2_), .B(i_6_), .Y(men_men_n92_));
  NO3        u0070(.A(men_men_n92_), .B(men_men_n49_), .C(men_men_n25_), .Y(men_men_n93_));
  NO2        u0071(.A(men_men_n93_), .B(men_men_n91_), .Y(men_men_n94_));
  AOI210     u0072(.A0(men_men_n94_), .A1(men_men_n88_), .B0(men_men_n80_), .Y(men_men_n95_));
  AN3        u0073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n96_));
  NAi21      u0074(.An(i_6_), .B(i_11_), .Y(men_men_n97_));
  NO2        u0075(.A(i_5_), .B(i_8_), .Y(men_men_n98_));
  NOi21      u0076(.An(men_men_n98_), .B(men_men_n97_), .Y(men_men_n99_));
  AOI220     u0077(.A0(men_men_n99_), .A1(men_men_n62_), .B0(men_men_n96_), .B1(men_men_n32_), .Y(men_men_n100_));
  INV        u0078(.A(i_7_), .Y(men_men_n101_));
  NA2        u0079(.A(men_men_n46_), .B(men_men_n101_), .Y(men_men_n102_));
  NO2        u0080(.A(i_0_), .B(i_5_), .Y(men_men_n103_));
  NO2        u0081(.A(men_men_n103_), .B(men_men_n85_), .Y(men_men_n104_));
  NA2        u0082(.A(i_12_), .B(i_3_), .Y(men_men_n105_));
  INV        u0083(.A(men_men_n105_), .Y(men_men_n106_));
  NA3        u0084(.A(men_men_n106_), .B(men_men_n104_), .C(men_men_n102_), .Y(men_men_n107_));
  NAi21      u0085(.An(i_7_), .B(i_11_), .Y(men_men_n108_));
  AN2        u0086(.A(i_2_), .B(i_10_), .Y(men_men_n109_));
  NO2        u0087(.A(men_men_n109_), .B(i_7_), .Y(men_men_n110_));
  OR2        u0088(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n111_));
  NO2        u0089(.A(i_8_), .B(men_men_n101_), .Y(men_men_n112_));
  NO3        u0090(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n110_), .Y(men_men_n113_));
  NA2        u0091(.A(i_12_), .B(i_7_), .Y(men_men_n114_));
  NO2        u0092(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n115_));
  NA2        u0093(.A(men_men_n115_), .B(i_0_), .Y(men_men_n116_));
  NA2        u0094(.A(i_11_), .B(i_12_), .Y(men_men_n117_));
  OAI210     u0095(.A0(men_men_n116_), .A1(men_men_n114_), .B0(men_men_n117_), .Y(men_men_n118_));
  NO2        u0096(.A(men_men_n118_), .B(men_men_n113_), .Y(men_men_n119_));
  NA3        u0097(.A(men_men_n119_), .B(men_men_n107_), .C(men_men_n100_), .Y(men_men_n120_));
  NOi21      u0098(.An(i_1_), .B(i_5_), .Y(men_men_n121_));
  NA2        u0099(.A(men_men_n121_), .B(i_11_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n101_), .B(men_men_n37_), .Y(men_men_n123_));
  NA2        u0101(.A(i_7_), .B(men_men_n25_), .Y(men_men_n124_));
  NA2        u0102(.A(men_men_n124_), .B(men_men_n123_), .Y(men_men_n125_));
  NO2        u0103(.A(men_men_n125_), .B(men_men_n46_), .Y(men_men_n126_));
  NA2        u0104(.A(men_men_n90_), .B(men_men_n89_), .Y(men_men_n127_));
  NAi21      u0105(.An(i_3_), .B(i_8_), .Y(men_men_n128_));
  NA2        u0106(.A(men_men_n128_), .B(men_men_n62_), .Y(men_men_n129_));
  NOi31      u0107(.An(men_men_n129_), .B(men_men_n127_), .C(men_men_n126_), .Y(men_men_n130_));
  NO2        u0108(.A(i_1_), .B(men_men_n85_), .Y(men_men_n131_));
  NO2        u0109(.A(i_6_), .B(i_5_), .Y(men_men_n132_));
  NA2        u0110(.A(men_men_n132_), .B(i_3_), .Y(men_men_n133_));
  AO210      u0111(.A0(men_men_n133_), .A1(men_men_n47_), .B0(men_men_n131_), .Y(men_men_n134_));
  OAI220     u0112(.A0(men_men_n134_), .A1(men_men_n108_), .B0(men_men_n130_), .B1(men_men_n122_), .Y(men_men_n135_));
  NO3        u0113(.A(men_men_n135_), .B(men_men_n120_), .C(men_men_n95_), .Y(men_men_n136_));
  NA3        u0114(.A(men_men_n136_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0115(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n138_));
  NA2        u0116(.A(i_6_), .B(men_men_n25_), .Y(men_men_n139_));
  NA2        u0117(.A(men_men_n139_), .B(men_men_n138_), .Y(men_men_n140_));
  NA4        u0118(.A(men_men_n140_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0119(.A(i_8_), .B(i_7_), .Y(men_men_n142_));
  NA2        u0120(.A(men_men_n142_), .B(i_6_), .Y(men_men_n143_));
  NO2        u0121(.A(i_12_), .B(i_13_), .Y(men_men_n144_));
  NAi21      u0122(.An(i_5_), .B(i_11_), .Y(men_men_n145_));
  NOi21      u0123(.An(men_men_n144_), .B(men_men_n145_), .Y(men_men_n146_));
  NO2        u0124(.A(i_0_), .B(i_1_), .Y(men_men_n147_));
  NA2        u0125(.A(i_2_), .B(i_3_), .Y(men_men_n148_));
  NO2        u0126(.A(men_men_n148_), .B(i_4_), .Y(men_men_n149_));
  NA3        u0127(.A(men_men_n149_), .B(men_men_n147_), .C(men_men_n146_), .Y(men_men_n150_));
  OR2        u0128(.A(men_men_n150_), .B(men_men_n25_), .Y(men_men_n151_));
  AN2        u0129(.A(men_men_n144_), .B(men_men_n82_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n152_), .B(men_men_n27_), .Y(men_men_n153_));
  NA2        u0131(.A(i_1_), .B(i_5_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n73_), .B(men_men_n46_), .Y(men_men_n155_));
  NA2        u0133(.A(men_men_n155_), .B(men_men_n36_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n156_), .B(men_men_n154_), .C(men_men_n153_), .Y(men_men_n157_));
  OR2        u0135(.A(i_0_), .B(i_1_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n159_));
  NAi32      u0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n160_));
  NAi21      u0138(.An(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0139(.An(i_4_), .B(i_10_), .Y(men_men_n162_));
  NA2        u0140(.A(men_men_n162_), .B(men_men_n40_), .Y(men_men_n163_));
  NO2        u0141(.A(i_3_), .B(i_5_), .Y(men_men_n164_));
  NO3        u0142(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n165_));
  INV        u0143(.A(men_men_n165_), .Y(men_men_n166_));
  OAI210     u0144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n167_));
  NO2        u0145(.A(men_men_n167_), .B(men_men_n157_), .Y(men_men_n168_));
  AOI210     u0146(.A0(men_men_n168_), .A1(men_men_n151_), .B0(men_men_n143_), .Y(men_men_n169_));
  NA2        u0147(.A(men_men_n46_), .B(i_1_), .Y(men_men_n170_));
  NA2        u0148(.A(i_3_), .B(men_men_n48_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_4_), .B(i_9_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_11_), .B(i_13_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  OR2        u0152(.A(men_men_n174_), .B(men_men_n171_), .Y(men_men_n175_));
  NO2        u0153(.A(i_4_), .B(i_5_), .Y(men_men_n176_));
  NAi21      u0154(.An(i_12_), .B(i_11_), .Y(men_men_n177_));
  NO2        u0155(.A(men_men_n177_), .B(i_13_), .Y(men_men_n178_));
  NA3        u0156(.A(men_men_n178_), .B(men_men_n176_), .C(men_men_n82_), .Y(men_men_n179_));
  AOI210     u0157(.A0(men_men_n179_), .A1(men_men_n175_), .B0(men_men_n170_), .Y(men_men_n180_));
  NO2        u0158(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n181_));
  NA2        u0159(.A(men_men_n181_), .B(men_men_n46_), .Y(men_men_n182_));
  NA2        u0160(.A(men_men_n36_), .B(i_5_), .Y(men_men_n183_));
  NAi31      u0161(.An(men_men_n183_), .B(men_men_n152_), .C(i_11_), .Y(men_men_n184_));
  NA2        u0162(.A(i_3_), .B(i_5_), .Y(men_men_n185_));
  OR2        u0163(.A(men_men_n185_), .B(men_men_n174_), .Y(men_men_n186_));
  AOI210     u0164(.A0(men_men_n186_), .A1(men_men_n184_), .B0(men_men_n182_), .Y(men_men_n187_));
  NO2        u0165(.A(men_men_n73_), .B(i_5_), .Y(men_men_n188_));
  NO2        u0166(.A(i_13_), .B(i_10_), .Y(men_men_n189_));
  NA3        u0167(.A(men_men_n189_), .B(men_men_n188_), .C(men_men_n44_), .Y(men_men_n190_));
  NO2        u0168(.A(i_2_), .B(i_1_), .Y(men_men_n191_));
  NA2        u0169(.A(men_men_n191_), .B(i_3_), .Y(men_men_n192_));
  NAi21      u0170(.An(i_4_), .B(i_12_), .Y(men_men_n193_));
  NO4        u0171(.A(men_men_n193_), .B(men_men_n192_), .C(men_men_n190_), .D(men_men_n25_), .Y(men_men_n194_));
  NO3        u0172(.A(men_men_n194_), .B(men_men_n187_), .C(men_men_n180_), .Y(men_men_n195_));
  INV        u0173(.A(i_8_), .Y(men_men_n196_));
  NA2        u0174(.A(i_8_), .B(i_6_), .Y(men_men_n197_));
  NO3        u0175(.A(i_3_), .B(men_men_n85_), .C(men_men_n48_), .Y(men_men_n198_));
  NA2        u0176(.A(men_men_n198_), .B(men_men_n112_), .Y(men_men_n199_));
  NO3        u0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n200_));
  NA3        u0178(.A(men_men_n200_), .B(men_men_n40_), .C(men_men_n44_), .Y(men_men_n201_));
  NO3        u0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n202_));
  OAI210     u0180(.A0(men_men_n96_), .A1(i_12_), .B0(men_men_n202_), .Y(men_men_n203_));
  AOI210     u0181(.A0(men_men_n203_), .A1(men_men_n201_), .B0(men_men_n199_), .Y(men_men_n204_));
  NO2        u0182(.A(i_3_), .B(i_8_), .Y(men_men_n205_));
  NO3        u0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n206_));
  NA3        u0184(.A(men_men_n206_), .B(men_men_n205_), .C(men_men_n40_), .Y(men_men_n207_));
  NO2        u0185(.A(i_13_), .B(i_9_), .Y(men_men_n208_));
  NA3        u0186(.A(men_men_n208_), .B(i_6_), .C(men_men_n196_), .Y(men_men_n209_));
  NAi21      u0187(.An(i_12_), .B(i_3_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n44_), .B(i_5_), .Y(men_men_n211_));
  NO3        u0189(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n212_));
  NA3        u0190(.A(men_men_n212_), .B(men_men_n211_), .C(i_10_), .Y(men_men_n213_));
  OAI220     u0191(.A0(men_men_n213_), .A1(men_men_n209_), .B0(men_men_n103_), .B1(men_men_n207_), .Y(men_men_n214_));
  AOI210     u0192(.A0(men_men_n214_), .A1(i_7_), .B0(men_men_n204_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(i_4_), .B0(men_men_n197_), .B1(men_men_n195_), .Y(men_men_n216_));
  NAi21      u0194(.An(i_12_), .B(i_7_), .Y(men_men_n217_));
  NA3        u0195(.A(i_13_), .B(men_men_n196_), .C(i_10_), .Y(men_men_n218_));
  NO2        u0196(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n219_));
  NA2        u0197(.A(i_0_), .B(i_5_), .Y(men_men_n220_));
  NA2        u0198(.A(men_men_n220_), .B(men_men_n104_), .Y(men_men_n221_));
  OAI220     u0199(.A0(men_men_n221_), .A1(men_men_n192_), .B0(men_men_n182_), .B1(men_men_n133_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n36_), .B(i_13_), .Y(men_men_n223_));
  NO2        u0201(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n224_));
  NO2        u0202(.A(men_men_n46_), .B(men_men_n63_), .Y(men_men_n225_));
  NA3        u0203(.A(men_men_n225_), .B(men_men_n224_), .C(men_men_n223_), .Y(men_men_n226_));
  INV        u0204(.A(i_13_), .Y(men_men_n227_));
  NO2        u0205(.A(i_12_), .B(men_men_n227_), .Y(men_men_n228_));
  NA3        u0206(.A(men_men_n228_), .B(men_men_n200_), .C(men_men_n198_), .Y(men_men_n229_));
  OAI210     u0207(.A0(men_men_n226_), .A1(i_9_), .B0(men_men_n229_), .Y(men_men_n230_));
  AOI220     u0208(.A0(men_men_n230_), .A1(men_men_n142_), .B0(men_men_n222_), .B1(men_men_n219_), .Y(men_men_n231_));
  NO2        u0209(.A(i_12_), .B(men_men_n37_), .Y(men_men_n232_));
  NO2        u0210(.A(men_men_n185_), .B(i_4_), .Y(men_men_n233_));
  NA2        u0211(.A(men_men_n233_), .B(men_men_n232_), .Y(men_men_n234_));
  OR2        u0212(.A(i_8_), .B(i_7_), .Y(men_men_n235_));
  NO2        u0213(.A(men_men_n235_), .B(men_men_n85_), .Y(men_men_n236_));
  NO2        u0214(.A(men_men_n53_), .B(i_1_), .Y(men_men_n237_));
  NA2        u0215(.A(men_men_n237_), .B(men_men_n236_), .Y(men_men_n238_));
  INV        u0216(.A(i_12_), .Y(men_men_n239_));
  NO2        u0217(.A(men_men_n44_), .B(men_men_n239_), .Y(men_men_n240_));
  NO3        u0218(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n241_));
  NA2        u0219(.A(i_2_), .B(i_1_), .Y(men_men_n242_));
  NO2        u0220(.A(men_men_n238_), .B(men_men_n234_), .Y(men_men_n243_));
  NO3        u0221(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n244_));
  NAi21      u0222(.An(i_4_), .B(i_3_), .Y(men_men_n245_));
  INV        u0223(.A(men_men_n75_), .Y(men_men_n246_));
  NO2        u0224(.A(i_0_), .B(i_6_), .Y(men_men_n247_));
  NOi41      u0225(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n248_));
  NA2        u0226(.A(men_men_n248_), .B(men_men_n247_), .Y(men_men_n249_));
  NO2        u0227(.A(men_men_n242_), .B(men_men_n185_), .Y(men_men_n250_));
  NAi21      u0228(.An(men_men_n249_), .B(men_men_n250_), .Y(men_men_n251_));
  INV        u0229(.A(men_men_n251_), .Y(men_men_n252_));
  AOI220     u0230(.A0(men_men_n252_), .A1(men_men_n40_), .B0(men_men_n243_), .B1(men_men_n208_), .Y(men_men_n253_));
  NO2        u0231(.A(i_11_), .B(men_men_n227_), .Y(men_men_n254_));
  NOi21      u0232(.An(i_1_), .B(i_6_), .Y(men_men_n255_));
  NAi21      u0233(.An(i_3_), .B(i_7_), .Y(men_men_n256_));
  NA2        u0234(.A(men_men_n239_), .B(i_9_), .Y(men_men_n257_));
  OR4        u0235(.A(men_men_n257_), .B(men_men_n256_), .C(men_men_n255_), .D(men_men_n188_), .Y(men_men_n258_));
  NO2        u0236(.A(i_12_), .B(i_3_), .Y(men_men_n259_));
  NA2        u0237(.A(men_men_n73_), .B(i_5_), .Y(men_men_n260_));
  NA2        u0238(.A(i_3_), .B(i_9_), .Y(men_men_n261_));
  NAi21      u0239(.An(i_7_), .B(i_10_), .Y(men_men_n262_));
  NO2        u0240(.A(men_men_n262_), .B(men_men_n261_), .Y(men_men_n263_));
  NA3        u0241(.A(men_men_n263_), .B(men_men_n260_), .C(men_men_n64_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n264_), .B(men_men_n258_), .Y(men_men_n265_));
  NA3        u0243(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n266_));
  INV        u0244(.A(men_men_n143_), .Y(men_men_n267_));
  NA2        u0245(.A(men_men_n239_), .B(i_13_), .Y(men_men_n268_));
  NO2        u0246(.A(men_men_n268_), .B(men_men_n75_), .Y(men_men_n269_));
  AOI220     u0247(.A0(men_men_n269_), .A1(men_men_n267_), .B0(men_men_n265_), .B1(men_men_n254_), .Y(men_men_n270_));
  NO2        u0248(.A(men_men_n235_), .B(men_men_n37_), .Y(men_men_n271_));
  NA2        u0249(.A(i_12_), .B(i_6_), .Y(men_men_n272_));
  OR2        u0250(.A(i_13_), .B(i_9_), .Y(men_men_n273_));
  NO3        u0251(.A(men_men_n273_), .B(men_men_n272_), .C(men_men_n48_), .Y(men_men_n274_));
  NO2        u0252(.A(men_men_n245_), .B(i_2_), .Y(men_men_n275_));
  NA3        u0253(.A(men_men_n275_), .B(men_men_n274_), .C(men_men_n44_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n254_), .B(i_9_), .Y(men_men_n277_));
  NA2        u0255(.A(men_men_n260_), .B(men_men_n64_), .Y(men_men_n278_));
  OAI210     u0256(.A0(men_men_n278_), .A1(men_men_n277_), .B0(men_men_n276_), .Y(men_men_n279_));
  NA2        u0257(.A(men_men_n155_), .B(men_men_n63_), .Y(men_men_n280_));
  NO3        u0258(.A(i_11_), .B(men_men_n227_), .C(men_men_n25_), .Y(men_men_n281_));
  NO2        u0259(.A(men_men_n256_), .B(i_8_), .Y(men_men_n282_));
  NO2        u0260(.A(i_6_), .B(men_men_n48_), .Y(men_men_n283_));
  NA3        u0261(.A(men_men_n283_), .B(men_men_n282_), .C(men_men_n281_), .Y(men_men_n284_));
  NO3        u0262(.A(men_men_n26_), .B(men_men_n85_), .C(i_5_), .Y(men_men_n285_));
  NA3        u0263(.A(men_men_n285_), .B(men_men_n271_), .C(men_men_n228_), .Y(men_men_n286_));
  AOI210     u0264(.A0(men_men_n286_), .A1(men_men_n284_), .B0(men_men_n280_), .Y(men_men_n287_));
  AOI210     u0265(.A0(men_men_n279_), .A1(men_men_n271_), .B0(men_men_n287_), .Y(men_men_n288_));
  NA4        u0266(.A(men_men_n288_), .B(men_men_n270_), .C(men_men_n253_), .D(men_men_n231_), .Y(men_men_n289_));
  NO3        u0267(.A(i_12_), .B(men_men_n227_), .C(men_men_n37_), .Y(men_men_n290_));
  INV        u0268(.A(men_men_n290_), .Y(men_men_n291_));
  NA2        u0269(.A(i_8_), .B(men_men_n101_), .Y(men_men_n292_));
  NO3        u0270(.A(i_0_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n293_));
  AOI220     u0271(.A0(men_men_n293_), .A1(men_men_n198_), .B0(men_men_n164_), .B1(men_men_n237_), .Y(men_men_n294_));
  NO2        u0272(.A(men_men_n294_), .B(men_men_n292_), .Y(men_men_n295_));
  NO2        u0273(.A(men_men_n242_), .B(i_0_), .Y(men_men_n296_));
  AOI220     u0274(.A0(men_men_n296_), .A1(i_8_), .B0(i_1_), .B1(men_men_n142_), .Y(men_men_n297_));
  NA2        u0275(.A(men_men_n283_), .B(men_men_n26_), .Y(men_men_n298_));
  NO2        u0276(.A(men_men_n298_), .B(men_men_n297_), .Y(men_men_n299_));
  NA2        u0277(.A(i_0_), .B(i_1_), .Y(men_men_n300_));
  NO2        u0278(.A(men_men_n300_), .B(i_2_), .Y(men_men_n301_));
  NO2        u0279(.A(men_men_n59_), .B(i_6_), .Y(men_men_n302_));
  NA3        u0280(.A(men_men_n302_), .B(men_men_n301_), .C(men_men_n164_), .Y(men_men_n303_));
  INV        u0281(.A(men_men_n303_), .Y(men_men_n304_));
  NO3        u0282(.A(men_men_n304_), .B(men_men_n299_), .C(men_men_n295_), .Y(men_men_n305_));
  NO2        u0283(.A(i_3_), .B(i_10_), .Y(men_men_n306_));
  NA3        u0284(.A(men_men_n306_), .B(men_men_n40_), .C(men_men_n44_), .Y(men_men_n307_));
  NO2        u0285(.A(i_2_), .B(men_men_n101_), .Y(men_men_n308_));
  NA2        u0286(.A(i_1_), .B(men_men_n36_), .Y(men_men_n309_));
  NOi21      u0287(.An(men_men_n220_), .B(men_men_n103_), .Y(men_men_n310_));
  NA3        u0288(.A(men_men_n310_), .B(men_men_n36_), .C(men_men_n308_), .Y(men_men_n311_));
  AN2        u0289(.A(i_3_), .B(i_10_), .Y(men_men_n312_));
  NA4        u0290(.A(men_men_n312_), .B(men_men_n200_), .C(men_men_n178_), .D(men_men_n176_), .Y(men_men_n313_));
  NO2        u0291(.A(i_5_), .B(men_men_n37_), .Y(men_men_n314_));
  NO2        u0292(.A(men_men_n46_), .B(men_men_n26_), .Y(men_men_n315_));
  OR2        u0293(.A(men_men_n311_), .B(men_men_n307_), .Y(men_men_n316_));
  OAI220     u0294(.A0(men_men_n316_), .A1(i_6_), .B0(men_men_n305_), .B1(men_men_n291_), .Y(men_men_n317_));
  NO4        u0295(.A(men_men_n317_), .B(men_men_n289_), .C(men_men_n216_), .D(men_men_n169_), .Y(men_men_n318_));
  NO3        u0296(.A(men_men_n44_), .B(i_13_), .C(i_9_), .Y(men_men_n319_));
  NO2        u0297(.A(men_men_n59_), .B(men_men_n85_), .Y(men_men_n320_));
  NA2        u0298(.A(men_men_n296_), .B(men_men_n320_), .Y(men_men_n321_));
  NO3        u0299(.A(i_6_), .B(men_men_n196_), .C(i_7_), .Y(men_men_n322_));
  NA2        u0300(.A(men_men_n322_), .B(men_men_n200_), .Y(men_men_n323_));
  AOI210     u0301(.A0(men_men_n323_), .A1(men_men_n321_), .B0(men_men_n171_), .Y(men_men_n324_));
  NO2        u0302(.A(i_2_), .B(i_3_), .Y(men_men_n325_));
  OR2        u0303(.A(i_0_), .B(i_5_), .Y(men_men_n326_));
  NA2        u0304(.A(men_men_n220_), .B(men_men_n326_), .Y(men_men_n327_));
  NA4        u0305(.A(men_men_n327_), .B(men_men_n236_), .C(men_men_n325_), .D(i_1_), .Y(men_men_n328_));
  NA3        u0306(.A(men_men_n296_), .B(men_men_n164_), .C(men_men_n112_), .Y(men_men_n329_));
  NAi21      u0307(.An(i_8_), .B(i_7_), .Y(men_men_n330_));
  NO2        u0308(.A(men_men_n330_), .B(i_6_), .Y(men_men_n331_));
  NO2        u0309(.A(men_men_n158_), .B(men_men_n46_), .Y(men_men_n332_));
  NA3        u0310(.A(men_men_n332_), .B(men_men_n331_), .C(men_men_n164_), .Y(men_men_n333_));
  NA3        u0311(.A(men_men_n333_), .B(men_men_n329_), .C(men_men_n328_), .Y(men_men_n334_));
  OAI210     u0312(.A0(men_men_n334_), .A1(men_men_n324_), .B0(i_4_), .Y(men_men_n335_));
  NO2        u0313(.A(i_12_), .B(i_10_), .Y(men_men_n336_));
  NOi21      u0314(.An(i_5_), .B(i_0_), .Y(men_men_n337_));
  NO2        u0315(.A(men_men_n309_), .B(men_men_n128_), .Y(men_men_n338_));
  NA2        u0316(.A(men_men_n338_), .B(men_men_n336_), .Y(men_men_n339_));
  NO2        u0317(.A(i_6_), .B(i_8_), .Y(men_men_n340_));
  NOi21      u0318(.An(i_0_), .B(i_2_), .Y(men_men_n341_));
  AN2        u0319(.A(men_men_n341_), .B(men_men_n340_), .Y(men_men_n342_));
  NO2        u0320(.A(i_1_), .B(i_7_), .Y(men_men_n343_));
  AO220      u0321(.A0(men_men_n343_), .A1(men_men_n342_), .B0(men_men_n331_), .B1(men_men_n237_), .Y(men_men_n344_));
  NA2        u0322(.A(men_men_n344_), .B(i_4_), .Y(men_men_n345_));
  NA3        u0323(.A(men_men_n345_), .B(men_men_n339_), .C(men_men_n335_), .Y(men_men_n346_));
  NO3        u0324(.A(men_men_n235_), .B(men_men_n46_), .C(i_1_), .Y(men_men_n347_));
  NO3        u0325(.A(men_men_n330_), .B(i_2_), .C(i_1_), .Y(men_men_n348_));
  OAI210     u0326(.A0(men_men_n348_), .A1(men_men_n347_), .B0(i_6_), .Y(men_men_n349_));
  NA2        u0327(.A(men_men_n255_), .B(men_men_n308_), .Y(men_men_n350_));
  AOI210     u0328(.A0(men_men_n350_), .A1(men_men_n349_), .B0(men_men_n327_), .Y(men_men_n351_));
  NOi21      u0329(.An(men_men_n154_), .B(men_men_n104_), .Y(men_men_n352_));
  NO2        u0330(.A(men_men_n352_), .B(men_men_n124_), .Y(men_men_n353_));
  OAI210     u0331(.A0(men_men_n353_), .A1(men_men_n351_), .B0(i_3_), .Y(men_men_n354_));
  INV        u0332(.A(men_men_n83_), .Y(men_men_n355_));
  NO2        u0333(.A(men_men_n300_), .B(men_men_n81_), .Y(men_men_n356_));
  NA2        u0334(.A(men_men_n356_), .B(men_men_n132_), .Y(men_men_n357_));
  NO2        u0335(.A(men_men_n92_), .B(men_men_n196_), .Y(men_men_n358_));
  NA3        u0336(.A(men_men_n310_), .B(men_men_n358_), .C(men_men_n63_), .Y(men_men_n359_));
  AOI210     u0337(.A0(men_men_n359_), .A1(men_men_n357_), .B0(men_men_n355_), .Y(men_men_n360_));
  NO2        u0338(.A(men_men_n196_), .B(i_9_), .Y(men_men_n361_));
  NO2        u0339(.A(men_men_n360_), .B(men_men_n299_), .Y(men_men_n362_));
  AOI210     u0340(.A0(men_men_n362_), .A1(men_men_n354_), .B0(men_men_n163_), .Y(men_men_n363_));
  AOI210     u0341(.A0(men_men_n346_), .A1(men_men_n319_), .B0(men_men_n363_), .Y(men_men_n364_));
  NOi32      u0342(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n365_));
  INV        u0343(.A(men_men_n365_), .Y(men_men_n366_));
  NAi21      u0344(.An(i_0_), .B(i_6_), .Y(men_men_n367_));
  NAi21      u0345(.An(i_1_), .B(i_5_), .Y(men_men_n368_));
  NA2        u0346(.A(men_men_n368_), .B(men_men_n367_), .Y(men_men_n369_));
  NA2        u0347(.A(men_men_n369_), .B(men_men_n25_), .Y(men_men_n370_));
  OAI210     u0348(.A0(men_men_n370_), .A1(men_men_n160_), .B0(men_men_n249_), .Y(men_men_n371_));
  NAi41      u0349(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n372_));
  AOI210     u0350(.A0(men_men_n372_), .A1(men_men_n160_), .B0(men_men_n158_), .Y(men_men_n373_));
  NOi32      u0351(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n374_));
  NO2        u0352(.A(i_1_), .B(men_men_n101_), .Y(men_men_n375_));
  NAi21      u0353(.An(i_3_), .B(i_4_), .Y(men_men_n376_));
  NO2        u0354(.A(men_men_n376_), .B(i_9_), .Y(men_men_n377_));
  AN2        u0355(.A(i_6_), .B(i_7_), .Y(men_men_n378_));
  OAI210     u0356(.A0(men_men_n378_), .A1(men_men_n375_), .B0(men_men_n377_), .Y(men_men_n379_));
  NA2        u0357(.A(i_2_), .B(i_7_), .Y(men_men_n380_));
  NO2        u0358(.A(men_men_n376_), .B(i_10_), .Y(men_men_n381_));
  NA3        u0359(.A(men_men_n381_), .B(men_men_n380_), .C(men_men_n247_), .Y(men_men_n382_));
  AOI210     u0360(.A0(men_men_n382_), .A1(men_men_n379_), .B0(men_men_n188_), .Y(men_men_n383_));
  AOI210     u0361(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n384_));
  AOI220     u0362(.A0(men_men_n381_), .A1(men_men_n343_), .B0(men_men_n241_), .B1(men_men_n191_), .Y(men_men_n385_));
  NO3        u0363(.A(men_men_n383_), .B(men_men_n373_), .C(men_men_n371_), .Y(men_men_n386_));
  NO2        u0364(.A(men_men_n386_), .B(men_men_n366_), .Y(men_men_n387_));
  NO2        u0365(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n388_));
  AN2        u0366(.A(i_12_), .B(i_5_), .Y(men_men_n389_));
  NO2        u0367(.A(i_4_), .B(men_men_n26_), .Y(men_men_n390_));
  NA2        u0368(.A(men_men_n390_), .B(men_men_n389_), .Y(men_men_n391_));
  NO2        u0369(.A(i_11_), .B(i_6_), .Y(men_men_n392_));
  NA3        u0370(.A(men_men_n392_), .B(men_men_n332_), .C(men_men_n227_), .Y(men_men_n393_));
  NO2        u0371(.A(men_men_n393_), .B(men_men_n391_), .Y(men_men_n394_));
  NO2        u0372(.A(men_men_n245_), .B(i_5_), .Y(men_men_n395_));
  NO2        u0373(.A(i_5_), .B(i_10_), .Y(men_men_n396_));
  NA2        u0374(.A(men_men_n395_), .B(men_men_n200_), .Y(men_men_n397_));
  NO2        u0375(.A(i_12_), .B(men_men_n397_), .Y(men_men_n398_));
  OAI210     u0376(.A0(men_men_n398_), .A1(men_men_n394_), .B0(men_men_n388_), .Y(men_men_n399_));
  NO2        u0377(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n400_));
  INV        u0378(.A(men_men_n150_), .Y(men_men_n401_));
  OAI210     u0379(.A0(men_men_n401_), .A1(men_men_n394_), .B0(men_men_n400_), .Y(men_men_n402_));
  NO3        u0380(.A(men_men_n85_), .B(men_men_n48_), .C(i_9_), .Y(men_men_n403_));
  NA2        u0381(.A(men_men_n306_), .B(men_men_n90_), .Y(men_men_n404_));
  NO2        u0382(.A(i_11_), .B(i_12_), .Y(men_men_n405_));
  NA2        u0383(.A(men_men_n405_), .B(men_men_n36_), .Y(men_men_n406_));
  NO2        u0384(.A(men_men_n404_), .B(men_men_n406_), .Y(men_men_n407_));
  NA2        u0385(.A(men_men_n396_), .B(men_men_n239_), .Y(men_men_n408_));
  NA3        u0386(.A(men_men_n112_), .B(i_4_), .C(i_11_), .Y(men_men_n409_));
  NO2        u0387(.A(men_men_n409_), .B(i_9_), .Y(men_men_n410_));
  NAi21      u0388(.An(i_13_), .B(i_0_), .Y(men_men_n411_));
  NO2        u0389(.A(men_men_n411_), .B(men_men_n242_), .Y(men_men_n412_));
  OAI210     u0390(.A0(men_men_n410_), .A1(men_men_n407_), .B0(men_men_n412_), .Y(men_men_n413_));
  NA3        u0391(.A(men_men_n413_), .B(men_men_n402_), .C(men_men_n399_), .Y(men_men_n414_));
  NO2        u0392(.A(i_0_), .B(i_11_), .Y(men_men_n415_));
  INV        u0393(.A(i_5_), .Y(men_men_n416_));
  AN2        u0394(.A(i_1_), .B(i_6_), .Y(men_men_n417_));
  NOi21      u0395(.An(i_2_), .B(i_12_), .Y(men_men_n418_));
  NA2        u0396(.A(men_men_n418_), .B(men_men_n417_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n419_), .B(men_men_n416_), .Y(men_men_n420_));
  NA2        u0398(.A(men_men_n142_), .B(i_9_), .Y(men_men_n421_));
  NO2        u0399(.A(men_men_n421_), .B(i_4_), .Y(men_men_n422_));
  NA2        u0400(.A(men_men_n420_), .B(men_men_n422_), .Y(men_men_n423_));
  NAi21      u0401(.An(i_9_), .B(i_4_), .Y(men_men_n424_));
  OR2        u0402(.A(i_13_), .B(i_10_), .Y(men_men_n425_));
  NO3        u0403(.A(men_men_n425_), .B(men_men_n117_), .C(men_men_n424_), .Y(men_men_n426_));
  NO2        u0404(.A(men_men_n174_), .B(men_men_n123_), .Y(men_men_n427_));
  NO2        u0405(.A(men_men_n101_), .B(men_men_n25_), .Y(men_men_n428_));
  NA2        u0406(.A(men_men_n290_), .B(men_men_n428_), .Y(men_men_n429_));
  NA2        u0407(.A(men_men_n283_), .B(men_men_n212_), .Y(men_men_n430_));
  OAI220     u0408(.A0(men_men_n430_), .A1(men_men_n218_), .B0(men_men_n429_), .B1(men_men_n352_), .Y(men_men_n431_));
  INV        u0409(.A(men_men_n431_), .Y(men_men_n432_));
  AOI210     u0410(.A0(men_men_n432_), .A1(men_men_n423_), .B0(men_men_n26_), .Y(men_men_n433_));
  NA2        u0411(.A(men_men_n329_), .B(men_men_n328_), .Y(men_men_n434_));
  AOI220     u0412(.A0(men_men_n302_), .A1(men_men_n293_), .B0(men_men_n296_), .B1(men_men_n320_), .Y(men_men_n435_));
  NO2        u0413(.A(men_men_n435_), .B(men_men_n171_), .Y(men_men_n436_));
  NO2        u0414(.A(men_men_n185_), .B(men_men_n85_), .Y(men_men_n437_));
  AOI220     u0415(.A0(men_men_n437_), .A1(men_men_n301_), .B0(men_men_n285_), .B1(men_men_n212_), .Y(men_men_n438_));
  NO2        u0416(.A(men_men_n438_), .B(men_men_n292_), .Y(men_men_n439_));
  NO3        u0417(.A(men_men_n439_), .B(men_men_n436_), .C(men_men_n434_), .Y(men_men_n440_));
  NA2        u0418(.A(men_men_n198_), .B(men_men_n96_), .Y(men_men_n441_));
  NA3        u0419(.A(men_men_n332_), .B(men_men_n164_), .C(men_men_n85_), .Y(men_men_n442_));
  AOI210     u0420(.A0(men_men_n442_), .A1(men_men_n441_), .B0(men_men_n330_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n302_), .B(men_men_n237_), .Y(men_men_n444_));
  NO2        u0422(.A(men_men_n444_), .B(men_men_n185_), .Y(men_men_n445_));
  NO2        u0423(.A(i_3_), .B(men_men_n48_), .Y(men_men_n446_));
  NO2        u0424(.A(men_men_n445_), .B(men_men_n443_), .Y(men_men_n447_));
  AOI210     u0425(.A0(men_men_n447_), .A1(men_men_n440_), .B0(men_men_n277_), .Y(men_men_n448_));
  NO4        u0426(.A(men_men_n448_), .B(men_men_n433_), .C(men_men_n414_), .D(men_men_n387_), .Y(men_men_n449_));
  NO2        u0427(.A(men_men_n63_), .B(i_4_), .Y(men_men_n450_));
  NO2        u0428(.A(men_men_n73_), .B(i_13_), .Y(men_men_n451_));
  NO2        u0429(.A(i_10_), .B(i_9_), .Y(men_men_n452_));
  NAi21      u0430(.An(i_12_), .B(i_8_), .Y(men_men_n453_));
  NO2        u0431(.A(men_men_n453_), .B(i_3_), .Y(men_men_n454_));
  NO2        u0432(.A(men_men_n46_), .B(i_4_), .Y(men_men_n455_));
  NA2        u0433(.A(men_men_n455_), .B(men_men_n104_), .Y(men_men_n456_));
  NO2        u0434(.A(men_men_n456_), .B(men_men_n207_), .Y(men_men_n457_));
  NA2        u0435(.A(men_men_n315_), .B(i_0_), .Y(men_men_n458_));
  NO3        u0436(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n459_));
  NA2        u0437(.A(men_men_n272_), .B(men_men_n97_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  NA2        u0439(.A(i_8_), .B(i_9_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n461_), .B(men_men_n458_), .Y(men_men_n463_));
  NO3        u0441(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n464_));
  NA3        u0442(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n465_));
  NA4        u0443(.A(men_men_n145_), .B(men_men_n115_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n466_));
  NO2        u0444(.A(men_men_n466_), .B(men_men_n465_), .Y(men_men_n467_));
  NO3        u0445(.A(men_men_n467_), .B(men_men_n463_), .C(men_men_n457_), .Y(men_men_n468_));
  OR2        u0446(.A(men_men_n300_), .B(men_men_n209_), .Y(men_men_n469_));
  BUFFER     u0447(.A(men_men_n303_), .Y(men_men_n470_));
  OA220      u0448(.A0(men_men_n470_), .A1(men_men_n163_), .B0(men_men_n469_), .B1(men_men_n234_), .Y(men_men_n471_));
  NA2        u0449(.A(men_men_n96_), .B(i_13_), .Y(men_men_n472_));
  NA2        u0450(.A(men_men_n437_), .B(men_men_n388_), .Y(men_men_n473_));
  NO2        u0451(.A(men_men_n473_), .B(men_men_n472_), .Y(men_men_n474_));
  NO3        u0452(.A(i_4_), .B(men_men_n48_), .C(i_8_), .Y(men_men_n475_));
  NO2        u0453(.A(i_6_), .B(i_7_), .Y(men_men_n476_));
  NA2        u0454(.A(men_men_n476_), .B(men_men_n475_), .Y(men_men_n477_));
  NO2        u0455(.A(i_11_), .B(i_1_), .Y(men_men_n478_));
  NO2        u0456(.A(men_men_n73_), .B(i_3_), .Y(men_men_n479_));
  NOi21      u0457(.An(i_2_), .B(i_7_), .Y(men_men_n480_));
  NAi31      u0458(.An(i_11_), .B(men_men_n480_), .C(men_men_n479_), .Y(men_men_n481_));
  NO2        u0459(.A(men_men_n425_), .B(i_6_), .Y(men_men_n482_));
  NA2        u0460(.A(men_men_n482_), .B(men_men_n450_), .Y(men_men_n483_));
  NO2        u0461(.A(men_men_n483_), .B(men_men_n481_), .Y(men_men_n484_));
  NO2        u0462(.A(i_6_), .B(i_10_), .Y(men_men_n485_));
  NA4        u0463(.A(men_men_n485_), .B(men_men_n319_), .C(i_8_), .D(men_men_n239_), .Y(men_men_n486_));
  NO2        u0464(.A(men_men_n486_), .B(men_men_n156_), .Y(men_men_n487_));
  NA2        u0465(.A(men_men_n46_), .B(men_men_n44_), .Y(men_men_n488_));
  NO2        u0466(.A(men_men_n158_), .B(i_3_), .Y(men_men_n489_));
  NAi31      u0467(.An(men_men_n488_), .B(men_men_n489_), .C(men_men_n228_), .Y(men_men_n490_));
  NA3        u0468(.A(men_men_n400_), .B(men_men_n181_), .C(men_men_n149_), .Y(men_men_n491_));
  NA2        u0469(.A(men_men_n491_), .B(men_men_n490_), .Y(men_men_n492_));
  NO4        u0470(.A(men_men_n492_), .B(men_men_n487_), .C(men_men_n484_), .D(men_men_n474_), .Y(men_men_n493_));
  NA2        u0471(.A(men_men_n464_), .B(men_men_n396_), .Y(men_men_n494_));
  NO2        u0472(.A(men_men_n494_), .B(men_men_n226_), .Y(men_men_n495_));
  NAi21      u0473(.An(men_men_n218_), .B(men_men_n405_), .Y(men_men_n496_));
  NA2        u0474(.A(men_men_n343_), .B(men_men_n220_), .Y(men_men_n497_));
  NO2        u0475(.A(men_men_n26_), .B(i_5_), .Y(men_men_n498_));
  NO2        u0476(.A(i_0_), .B(men_men_n85_), .Y(men_men_n499_));
  NA3        u0477(.A(men_men_n499_), .B(men_men_n498_), .C(men_men_n142_), .Y(men_men_n500_));
  OR3        u0478(.A(men_men_n309_), .B(men_men_n38_), .C(men_men_n46_), .Y(men_men_n501_));
  OAI220     u0479(.A0(men_men_n501_), .A1(men_men_n500_), .B0(men_men_n497_), .B1(men_men_n496_), .Y(men_men_n502_));
  NA2        u0480(.A(men_men_n27_), .B(i_10_), .Y(men_men_n503_));
  NO2        u0481(.A(men_men_n503_), .B(men_men_n472_), .Y(men_men_n504_));
  NA3        u0482(.A(men_men_n312_), .B(men_men_n225_), .C(men_men_n73_), .Y(men_men_n505_));
  NO2        u0483(.A(men_men_n505_), .B(men_men_n477_), .Y(men_men_n506_));
  NO4        u0484(.A(men_men_n506_), .B(men_men_n504_), .C(men_men_n502_), .D(men_men_n495_), .Y(men_men_n507_));
  NA4        u0485(.A(men_men_n507_), .B(men_men_n493_), .C(men_men_n471_), .D(men_men_n468_), .Y(men_men_n508_));
  NA3        u0486(.A(men_men_n312_), .B(men_men_n178_), .C(men_men_n176_), .Y(men_men_n509_));
  INV        u0487(.A(men_men_n509_), .Y(men_men_n510_));
  AN2        u0488(.A(men_men_n293_), .B(men_men_n236_), .Y(men_men_n511_));
  NA2        u0489(.A(men_men_n511_), .B(men_men_n510_), .Y(men_men_n512_));
  NA2        u0490(.A(men_men_n122_), .B(men_men_n111_), .Y(men_men_n513_));
  AN2        u0491(.A(men_men_n513_), .B(men_men_n459_), .Y(men_men_n514_));
  NA2        u0492(.A(men_men_n319_), .B(men_men_n165_), .Y(men_men_n515_));
  OAI210     u0493(.A0(men_men_n515_), .A1(men_men_n234_), .B0(men_men_n313_), .Y(men_men_n516_));
  AOI220     u0494(.A0(men_men_n516_), .A1(men_men_n331_), .B0(men_men_n514_), .B1(men_men_n315_), .Y(men_men_n517_));
  NA2        u0495(.A(men_men_n389_), .B(men_men_n227_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n365_), .B(men_men_n73_), .Y(men_men_n519_));
  NA2        u0497(.A(men_men_n378_), .B(men_men_n374_), .Y(men_men_n520_));
  AO210      u0498(.A0(men_men_n519_), .A1(men_men_n518_), .B0(men_men_n520_), .Y(men_men_n521_));
  NO2        u0499(.A(men_men_n36_), .B(i_8_), .Y(men_men_n522_));
  NAi41      u0500(.An(men_men_n519_), .B(men_men_n485_), .C(men_men_n522_), .D(men_men_n46_), .Y(men_men_n523_));
  AOI210     u0501(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n426_), .Y(men_men_n524_));
  NA3        u0502(.A(men_men_n524_), .B(men_men_n523_), .C(men_men_n521_), .Y(men_men_n525_));
  INV        u0503(.A(men_men_n525_), .Y(men_men_n526_));
  NA2        u0504(.A(men_men_n260_), .B(men_men_n64_), .Y(men_men_n527_));
  OAI210     u0505(.A0(i_8_), .A1(men_men_n527_), .B0(men_men_n134_), .Y(men_men_n528_));
  NO2        u0506(.A(i_7_), .B(men_men_n201_), .Y(men_men_n529_));
  OR2        u0507(.A(men_men_n185_), .B(i_4_), .Y(men_men_n530_));
  NO2        u0508(.A(men_men_n530_), .B(men_men_n85_), .Y(men_men_n531_));
  AOI220     u0509(.A0(men_men_n531_), .A1(men_men_n529_), .B0(men_men_n528_), .B1(men_men_n427_), .Y(men_men_n532_));
  NA4        u0510(.A(men_men_n532_), .B(men_men_n526_), .C(men_men_n517_), .D(men_men_n512_), .Y(men_men_n533_));
  NA2        u0511(.A(men_men_n395_), .B(men_men_n301_), .Y(men_men_n534_));
  OAI210     u0512(.A0(men_men_n391_), .A1(men_men_n170_), .B0(men_men_n534_), .Y(men_men_n535_));
  NA2        u0513(.A(men_men_n1041_), .B(men_men_n227_), .Y(men_men_n536_));
  NA2        u0514(.A(men_men_n485_), .B(men_men_n27_), .Y(men_men_n537_));
  NO2        u0515(.A(men_men_n537_), .B(men_men_n536_), .Y(men_men_n538_));
  NOi31      u0516(.An(men_men_n322_), .B(men_men_n425_), .C(men_men_n38_), .Y(men_men_n539_));
  OAI210     u0517(.A0(men_men_n539_), .A1(men_men_n538_), .B0(men_men_n535_), .Y(men_men_n540_));
  NO2        u0518(.A(i_8_), .B(i_7_), .Y(men_men_n541_));
  OAI210     u0519(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n542_));
  NA2        u0520(.A(men_men_n542_), .B(men_men_n225_), .Y(men_men_n543_));
  OAI220     u0521(.A0(men_men_n46_), .A1(men_men_n530_), .B0(men_men_n543_), .B1(men_men_n245_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n44_), .B(i_10_), .Y(men_men_n545_));
  NO2        u0523(.A(men_men_n545_), .B(i_6_), .Y(men_men_n546_));
  NA3        u0524(.A(men_men_n546_), .B(men_men_n544_), .C(men_men_n541_), .Y(men_men_n547_));
  AOI220     u0525(.A0(men_men_n437_), .A1(men_men_n332_), .B0(men_men_n250_), .B1(men_men_n247_), .Y(men_men_n548_));
  NO2        u0526(.A(men_men_n548_), .B(men_men_n268_), .Y(men_men_n549_));
  NA2        u0527(.A(men_men_n549_), .B(men_men_n271_), .Y(men_men_n550_));
  NO2        u0528(.A(men_men_n307_), .B(men_men_n183_), .Y(men_men_n551_));
  NA3        u0529(.A(men_men_n312_), .B(men_men_n176_), .C(men_men_n96_), .Y(men_men_n552_));
  NO2        u0530(.A(men_men_n223_), .B(men_men_n44_), .Y(men_men_n553_));
  NO2        u0531(.A(men_men_n158_), .B(i_5_), .Y(men_men_n554_));
  NA2        u0532(.A(men_men_n554_), .B(men_men_n325_), .Y(men_men_n555_));
  OAI210     u0533(.A0(men_men_n555_), .A1(men_men_n553_), .B0(men_men_n552_), .Y(men_men_n556_));
  OAI210     u0534(.A0(men_men_n556_), .A1(men_men_n551_), .B0(men_men_n464_), .Y(men_men_n557_));
  NA4        u0535(.A(men_men_n557_), .B(men_men_n550_), .C(men_men_n547_), .D(men_men_n540_), .Y(men_men_n558_));
  NA3        u0536(.A(men_men_n220_), .B(men_men_n71_), .C(men_men_n44_), .Y(men_men_n559_));
  NA2        u0537(.A(men_men_n290_), .B(men_men_n83_), .Y(men_men_n560_));
  AOI210     u0538(.A0(men_men_n559_), .A1(men_men_n357_), .B0(men_men_n560_), .Y(men_men_n561_));
  NA2        u0539(.A(men_men_n302_), .B(men_men_n293_), .Y(men_men_n562_));
  NO2        u0540(.A(men_men_n562_), .B(men_men_n175_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n564_));
  NA2        u0542(.A(men_men_n452_), .B(men_men_n223_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n564_), .B(men_men_n565_), .Y(men_men_n566_));
  NA2        u0544(.A(i_0_), .B(men_men_n48_), .Y(men_men_n567_));
  NO3        u0545(.A(men_men_n566_), .B(men_men_n563_), .C(men_men_n561_), .Y(men_men_n568_));
  NO4        u0546(.A(men_men_n255_), .B(men_men_n42_), .C(i_2_), .D(men_men_n48_), .Y(men_men_n569_));
  NO3        u0547(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n570_));
  NO2        u0548(.A(men_men_n235_), .B(men_men_n36_), .Y(men_men_n571_));
  AN2        u0549(.A(men_men_n571_), .B(men_men_n570_), .Y(men_men_n572_));
  OA210      u0550(.A0(men_men_n572_), .A1(men_men_n569_), .B0(men_men_n365_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n425_), .B(i_1_), .Y(men_men_n574_));
  NOi31      u0552(.An(men_men_n574_), .B(men_men_n460_), .C(men_men_n73_), .Y(men_men_n575_));
  AN4        u0553(.A(men_men_n575_), .B(men_men_n422_), .C(men_men_n498_), .D(i_2_), .Y(men_men_n576_));
  NO2        u0554(.A(men_men_n435_), .B(men_men_n179_), .Y(men_men_n577_));
  NO3        u0555(.A(men_men_n577_), .B(men_men_n576_), .C(men_men_n573_), .Y(men_men_n578_));
  NOi21      u0556(.An(i_10_), .B(i_6_), .Y(men_men_n579_));
  NO2        u0557(.A(men_men_n85_), .B(men_men_n25_), .Y(men_men_n580_));
  AOI220     u0558(.A0(men_men_n290_), .A1(men_men_n580_), .B0(men_men_n281_), .B1(men_men_n579_), .Y(men_men_n581_));
  NO2        u0559(.A(men_men_n581_), .B(men_men_n458_), .Y(men_men_n582_));
  NO2        u0560(.A(men_men_n114_), .B(men_men_n23_), .Y(men_men_n583_));
  NA2        u0561(.A(men_men_n322_), .B(men_men_n165_), .Y(men_men_n584_));
  AOI220     u0562(.A0(men_men_n584_), .A1(men_men_n444_), .B0(men_men_n186_), .B1(men_men_n184_), .Y(men_men_n585_));
  NO2        u0563(.A(men_men_n585_), .B(men_men_n582_), .Y(men_men_n586_));
  NO2        u0564(.A(men_men_n519_), .B(men_men_n385_), .Y(men_men_n587_));
  INV        u0565(.A(men_men_n325_), .Y(men_men_n588_));
  NO2        u0566(.A(i_12_), .B(men_men_n85_), .Y(men_men_n589_));
  NO3        u0567(.A(i_4_), .B(men_men_n349_), .C(men_men_n307_), .Y(men_men_n590_));
  OR2        u0568(.A(i_2_), .B(i_5_), .Y(men_men_n591_));
  OR2        u0569(.A(men_men_n591_), .B(men_men_n417_), .Y(men_men_n592_));
  NO2        u0570(.A(men_men_n592_), .B(men_men_n496_), .Y(men_men_n593_));
  NO3        u0571(.A(men_men_n593_), .B(men_men_n590_), .C(men_men_n587_), .Y(men_men_n594_));
  NA4        u0572(.A(men_men_n594_), .B(men_men_n586_), .C(men_men_n578_), .D(men_men_n568_), .Y(men_men_n595_));
  NO4        u0573(.A(men_men_n595_), .B(men_men_n558_), .C(men_men_n533_), .D(men_men_n508_), .Y(men_men_n596_));
  NA4        u0574(.A(men_men_n596_), .B(men_men_n449_), .C(men_men_n364_), .D(men_men_n318_), .Y(men7));
  NO2        u0575(.A(men_men_n92_), .B(men_men_n54_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n108_), .B(men_men_n89_), .Y(men_men_n599_));
  NA2        u0577(.A(i_11_), .B(men_men_n196_), .Y(men_men_n600_));
  NA3        u0578(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n601_));
  NO2        u0579(.A(men_men_n239_), .B(i_4_), .Y(men_men_n602_));
  NA2        u0580(.A(men_men_n602_), .B(i_8_), .Y(men_men_n603_));
  NO2        u0581(.A(men_men_n105_), .B(men_men_n601_), .Y(men_men_n604_));
  NA2        u0582(.A(i_2_), .B(men_men_n85_), .Y(men_men_n605_));
  OAI210     u0583(.A0(men_men_n86_), .A1(men_men_n205_), .B0(men_men_n206_), .Y(men_men_n606_));
  NO2        u0584(.A(i_7_), .B(men_men_n37_), .Y(men_men_n607_));
  NA2        u0585(.A(i_4_), .B(i_8_), .Y(men_men_n608_));
  AOI210     u0586(.A0(men_men_n608_), .A1(men_men_n312_), .B0(men_men_n607_), .Y(men_men_n609_));
  OAI220     u0587(.A0(men_men_n609_), .A1(men_men_n605_), .B0(men_men_n606_), .B1(i_13_), .Y(men_men_n610_));
  NO3        u0588(.A(men_men_n610_), .B(men_men_n604_), .C(men_men_n598_), .Y(men_men_n611_));
  OR2        u0589(.A(i_6_), .B(i_10_), .Y(men_men_n612_));
  NO2        u0590(.A(men_men_n612_), .B(men_men_n23_), .Y(men_men_n613_));
  OR3        u0591(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n614_));
  NO3        u0592(.A(men_men_n614_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n615_));
  INV        u0593(.A(men_men_n202_), .Y(men_men_n616_));
  NO2        u0594(.A(men_men_n615_), .B(men_men_n613_), .Y(men_men_n617_));
  OA220      u0595(.A0(men_men_n617_), .A1(men_men_n588_), .B0(men_men_n1043_), .B1(men_men_n273_), .Y(men_men_n618_));
  AOI210     u0596(.A0(men_men_n618_), .A1(men_men_n611_), .B0(men_men_n63_), .Y(men_men_n619_));
  NOi21      u0597(.An(i_11_), .B(i_7_), .Y(men_men_n620_));
  AO210      u0598(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n621_));
  NO2        u0599(.A(men_men_n621_), .B(men_men_n620_), .Y(men_men_n622_));
  NA2        u0600(.A(men_men_n622_), .B(men_men_n208_), .Y(men_men_n623_));
  NA3        u0601(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n624_));
  NAi31      u0602(.An(men_men_n624_), .B(men_men_n217_), .C(i_11_), .Y(men_men_n625_));
  AOI210     u0603(.A0(men_men_n625_), .A1(men_men_n623_), .B0(men_men_n63_), .Y(men_men_n626_));
  NO3        u0604(.A(men_men_n262_), .B(men_men_n210_), .C(men_men_n600_), .Y(men_men_n627_));
  OAI210     u0605(.A0(men_men_n627_), .A1(men_men_n228_), .B0(men_men_n63_), .Y(men_men_n628_));
  NA2        u0606(.A(men_men_n418_), .B(men_men_n31_), .Y(men_men_n629_));
  OR2        u0607(.A(men_men_n210_), .B(men_men_n108_), .Y(men_men_n630_));
  NA2        u0608(.A(men_men_n630_), .B(men_men_n629_), .Y(men_men_n631_));
  NO2        u0609(.A(men_men_n63_), .B(i_9_), .Y(men_men_n632_));
  NO2        u0610(.A(men_men_n632_), .B(i_4_), .Y(men_men_n633_));
  NA2        u0611(.A(men_men_n633_), .B(men_men_n631_), .Y(men_men_n634_));
  NO2        u0612(.A(i_1_), .B(i_12_), .Y(men_men_n635_));
  NA2        u0613(.A(men_men_n634_), .B(men_men_n628_), .Y(men_men_n636_));
  OAI210     u0614(.A0(men_men_n636_), .A1(men_men_n626_), .B0(i_6_), .Y(men_men_n637_));
  NO2        u0615(.A(men_men_n239_), .B(men_men_n85_), .Y(men_men_n638_));
  NO2        u0616(.A(men_men_n638_), .B(i_11_), .Y(men_men_n639_));
  INV        u0617(.A(men_men_n461_), .Y(men_men_n640_));
  NO4        u0618(.A(men_men_n217_), .B(men_men_n128_), .C(i_13_), .D(men_men_n85_), .Y(men_men_n641_));
  NA2        u0619(.A(men_men_n641_), .B(men_men_n632_), .Y(men_men_n642_));
  NA2        u0620(.A(men_men_n239_), .B(i_6_), .Y(men_men_n643_));
  NO3        u0621(.A(men_men_n612_), .B(men_men_n235_), .C(men_men_n23_), .Y(men_men_n644_));
  AOI210     u0622(.A0(i_1_), .A1(men_men_n263_), .B0(men_men_n644_), .Y(men_men_n645_));
  OAI210     u0623(.A0(men_men_n645_), .A1(men_men_n44_), .B0(men_men_n642_), .Y(men_men_n646_));
  NA3        u0624(.A(men_men_n541_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n647_));
  NA2        u0625(.A(men_men_n138_), .B(i_9_), .Y(men_men_n648_));
  NA3        u0626(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n649_));
  NO2        u0627(.A(men_men_n46_), .B(i_1_), .Y(men_men_n650_));
  NO2        u0628(.A(men_men_n648_), .B(men_men_n1040_), .Y(men_men_n651_));
  AOI210     u0629(.A0(men_men_n478_), .A1(men_men_n428_), .B0(men_men_n244_), .Y(men_men_n652_));
  NO2        u0630(.A(men_men_n652_), .B(men_men_n605_), .Y(men_men_n653_));
  NAi21      u0631(.An(men_men_n647_), .B(men_men_n91_), .Y(men_men_n654_));
  NA2        u0632(.A(men_men_n650_), .B(men_men_n272_), .Y(men_men_n655_));
  NO2        u0633(.A(i_11_), .B(men_men_n37_), .Y(men_men_n656_));
  NA2        u0634(.A(men_men_n656_), .B(men_men_n24_), .Y(men_men_n657_));
  OAI210     u0635(.A0(men_men_n657_), .A1(men_men_n655_), .B0(men_men_n654_), .Y(men_men_n658_));
  OR3        u0636(.A(men_men_n658_), .B(men_men_n653_), .C(men_men_n651_), .Y(men_men_n659_));
  NO3        u0637(.A(men_men_n659_), .B(men_men_n646_), .C(men_men_n640_), .Y(men_men_n660_));
  NO2        u0638(.A(men_men_n239_), .B(men_men_n101_), .Y(men_men_n661_));
  NO2        u0639(.A(men_men_n661_), .B(men_men_n620_), .Y(men_men_n662_));
  NA2        u0640(.A(men_men_n662_), .B(i_1_), .Y(men_men_n663_));
  NO2        u0641(.A(men_men_n663_), .B(men_men_n614_), .Y(men_men_n664_));
  NO2        u0642(.A(men_men_n424_), .B(men_men_n85_), .Y(men_men_n665_));
  NA2        u0643(.A(men_men_n664_), .B(men_men_n46_), .Y(men_men_n666_));
  NA2        u0644(.A(i_3_), .B(men_men_n196_), .Y(men_men_n667_));
  NO2        u0645(.A(men_men_n667_), .B(men_men_n114_), .Y(men_men_n668_));
  AN2        u0646(.A(men_men_n668_), .B(men_men_n546_), .Y(men_men_n669_));
  NO2        u0647(.A(men_men_n235_), .B(men_men_n44_), .Y(men_men_n670_));
  NO3        u0648(.A(men_men_n670_), .B(men_men_n315_), .C(men_men_n240_), .Y(men_men_n671_));
  NO2        u0649(.A(men_men_n117_), .B(men_men_n37_), .Y(men_men_n672_));
  NO2        u0650(.A(men_men_n672_), .B(i_6_), .Y(men_men_n673_));
  NO2        u0651(.A(men_men_n85_), .B(i_9_), .Y(men_men_n674_));
  NO2        u0652(.A(men_men_n674_), .B(men_men_n63_), .Y(men_men_n675_));
  NO2        u0653(.A(men_men_n675_), .B(men_men_n635_), .Y(men_men_n676_));
  NO4        u0654(.A(men_men_n676_), .B(men_men_n673_), .C(men_men_n671_), .D(i_4_), .Y(men_men_n677_));
  NA2        u0655(.A(i_1_), .B(i_3_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n462_), .B(men_men_n92_), .Y(men_men_n679_));
  AOI210     u0657(.A0(men_men_n670_), .A1(men_men_n579_), .B0(men_men_n679_), .Y(men_men_n680_));
  NO2        u0658(.A(men_men_n680_), .B(men_men_n678_), .Y(men_men_n681_));
  NO3        u0659(.A(men_men_n681_), .B(men_men_n677_), .C(men_men_n669_), .Y(men_men_n682_));
  NA4        u0660(.A(men_men_n682_), .B(men_men_n666_), .C(men_men_n660_), .D(men_men_n637_), .Y(men_men_n683_));
  NO3        u0661(.A(i_11_), .B(i_3_), .C(i_7_), .Y(men_men_n684_));
  NOi21      u0662(.An(men_men_n684_), .B(i_10_), .Y(men_men_n685_));
  OA210      u0663(.A0(men_men_n685_), .A1(men_men_n248_), .B0(men_men_n85_), .Y(men_men_n686_));
  NA2        u0664(.A(men_men_n378_), .B(men_men_n377_), .Y(men_men_n687_));
  NA3        u0665(.A(men_men_n485_), .B(men_men_n522_), .C(men_men_n46_), .Y(men_men_n688_));
  NO3        u0666(.A(men_men_n480_), .B(men_men_n608_), .C(men_men_n85_), .Y(men_men_n689_));
  NA2        u0667(.A(men_men_n689_), .B(men_men_n25_), .Y(men_men_n690_));
  NA3        u0668(.A(men_men_n690_), .B(men_men_n688_), .C(men_men_n687_), .Y(men_men_n691_));
  OAI210     u0669(.A0(men_men_n691_), .A1(men_men_n686_), .B0(i_1_), .Y(men_men_n692_));
  AOI210     u0670(.A0(men_men_n272_), .A1(men_men_n97_), .B0(i_1_), .Y(men_men_n693_));
  NO2        u0671(.A(men_men_n376_), .B(i_2_), .Y(men_men_n694_));
  NA2        u0672(.A(men_men_n694_), .B(men_men_n693_), .Y(men_men_n695_));
  AOI210     u0673(.A0(men_men_n695_), .A1(men_men_n692_), .B0(i_13_), .Y(men_men_n696_));
  OR2        u0674(.A(i_11_), .B(i_7_), .Y(men_men_n697_));
  NO2        u0675(.A(men_men_n54_), .B(i_12_), .Y(men_men_n698_));
  INV        u0676(.A(men_men_n698_), .Y(men_men_n699_));
  NO2        u0677(.A(men_men_n480_), .B(men_men_n24_), .Y(men_men_n700_));
  AOI220     u0678(.A0(men_men_n700_), .A1(men_men_n665_), .B0(men_men_n248_), .B1(men_men_n131_), .Y(men_men_n701_));
  OAI220     u0679(.A0(men_men_n701_), .A1(men_men_n41_), .B0(men_men_n699_), .B1(men_men_n92_), .Y(men_men_n702_));
  INV        u0680(.A(men_men_n702_), .Y(men_men_n703_));
  NA2        u0681(.A(men_men_n392_), .B(men_men_n650_), .Y(men_men_n704_));
  NO2        u0682(.A(men_men_n704_), .B(men_men_n245_), .Y(men_men_n705_));
  AOI210     u0683(.A0(men_men_n453_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n706_));
  NA2        u0684(.A(men_men_n127_), .B(i_13_), .Y(men_men_n707_));
  NO2        u0685(.A(men_men_n649_), .B(men_men_n114_), .Y(men_men_n708_));
  NO2        u0686(.A(men_men_n707_), .B(men_men_n693_), .Y(men_men_n709_));
  NA2        u0687(.A(men_men_n26_), .B(men_men_n196_), .Y(men_men_n710_));
  NA2        u0688(.A(men_men_n710_), .B(i_7_), .Y(men_men_n711_));
  NO3        u0689(.A(men_men_n480_), .B(men_men_n239_), .C(men_men_n85_), .Y(men_men_n712_));
  NA2        u0690(.A(men_men_n712_), .B(men_men_n711_), .Y(men_men_n713_));
  AOI220     u0691(.A0(men_men_n392_), .A1(men_men_n650_), .B0(men_men_n91_), .B1(men_men_n102_), .Y(men_men_n714_));
  OAI220     u0692(.A0(men_men_n714_), .A1(men_men_n603_), .B0(men_men_n713_), .B1(men_men_n616_), .Y(men_men_n715_));
  NO3        u0693(.A(men_men_n715_), .B(men_men_n709_), .C(men_men_n705_), .Y(men_men_n716_));
  OR2        u0694(.A(i_11_), .B(i_6_), .Y(men_men_n717_));
  NA3        u0695(.A(men_men_n418_), .B(men_men_n607_), .C(men_men_n97_), .Y(men_men_n718_));
  NA2        u0696(.A(men_men_n639_), .B(i_13_), .Y(men_men_n719_));
  NAi21      u0697(.An(i_11_), .B(i_12_), .Y(men_men_n720_));
  NA2        u0698(.A(men_men_n719_), .B(men_men_n718_), .Y(men_men_n721_));
  NA2        u0699(.A(men_men_n721_), .B(men_men_n63_), .Y(men_men_n722_));
  NO2        u0700(.A(i_2_), .B(i_12_), .Y(men_men_n723_));
  NA2        u0701(.A(men_men_n375_), .B(men_men_n723_), .Y(men_men_n724_));
  NA2        u0702(.A(i_8_), .B(men_men_n25_), .Y(men_men_n725_));
  NO3        u0703(.A(men_men_n725_), .B(men_men_n390_), .C(men_men_n602_), .Y(men_men_n726_));
  OAI210     u0704(.A0(men_men_n726_), .A1(men_men_n377_), .B0(men_men_n375_), .Y(men_men_n727_));
  NO2        u0705(.A(men_men_n128_), .B(i_2_), .Y(men_men_n728_));
  NA2        u0706(.A(men_men_n728_), .B(men_men_n635_), .Y(men_men_n729_));
  NA3        u0707(.A(men_men_n729_), .B(men_men_n727_), .C(men_men_n724_), .Y(men_men_n730_));
  NA3        u0708(.A(men_men_n730_), .B(men_men_n45_), .C(men_men_n227_), .Y(men_men_n731_));
  NA4        u0709(.A(men_men_n731_), .B(men_men_n722_), .C(men_men_n716_), .D(men_men_n703_), .Y(men_men_n732_));
  OR4        u0710(.A(men_men_n732_), .B(men_men_n696_), .C(men_men_n683_), .D(men_men_n619_), .Y(men5));
  AOI210     u0711(.A0(men_men_n662_), .A1(men_men_n275_), .B0(men_men_n427_), .Y(men_men_n734_));
  AN2        u0712(.A(men_men_n24_), .B(i_10_), .Y(men_men_n735_));
  NA3        u0713(.A(men_men_n735_), .B(men_men_n723_), .C(men_men_n108_), .Y(men_men_n736_));
  NO2        u0714(.A(men_men_n603_), .B(i_11_), .Y(men_men_n737_));
  NA2        u0715(.A(men_men_n86_), .B(men_men_n737_), .Y(men_men_n738_));
  NA3        u0716(.A(men_men_n738_), .B(men_men_n736_), .C(men_men_n734_), .Y(men_men_n739_));
  NO3        u0717(.A(i_11_), .B(men_men_n239_), .C(i_13_), .Y(men_men_n740_));
  NO2        u0718(.A(men_men_n124_), .B(men_men_n23_), .Y(men_men_n741_));
  NA2        u0719(.A(i_12_), .B(i_8_), .Y(men_men_n742_));
  OAI210     u0720(.A0(men_men_n46_), .A1(i_3_), .B0(men_men_n742_), .Y(men_men_n743_));
  INV        u0721(.A(men_men_n452_), .Y(men_men_n744_));
  AOI220     u0722(.A0(men_men_n325_), .A1(men_men_n583_), .B0(men_men_n743_), .B1(men_men_n741_), .Y(men_men_n745_));
  INV        u0723(.A(men_men_n745_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n746_), .B(men_men_n739_), .Y(men_men_n747_));
  INV        u0725(.A(men_men_n173_), .Y(men_men_n748_));
  INV        u0726(.A(men_men_n248_), .Y(men_men_n749_));
  OAI210     u0727(.A0(men_men_n694_), .A1(men_men_n454_), .B0(men_men_n110_), .Y(men_men_n750_));
  AOI210     u0728(.A0(men_men_n750_), .A1(men_men_n749_), .B0(men_men_n748_), .Y(men_men_n751_));
  NO2        u0729(.A(men_men_n462_), .B(men_men_n26_), .Y(men_men_n752_));
  NO2        u0730(.A(men_men_n752_), .B(men_men_n428_), .Y(men_men_n753_));
  NA2        u0731(.A(men_men_n753_), .B(i_2_), .Y(men_men_n754_));
  INV        u0732(.A(men_men_n754_), .Y(men_men_n755_));
  AOI210     u0733(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n425_), .Y(men_men_n756_));
  AOI210     u0734(.A0(men_men_n756_), .A1(men_men_n755_), .B0(men_men_n751_), .Y(men_men_n757_));
  NO2        u0735(.A(men_men_n193_), .B(men_men_n125_), .Y(men_men_n758_));
  OAI210     u0736(.A0(men_men_n758_), .A1(men_men_n741_), .B0(i_2_), .Y(men_men_n759_));
  NO2        u0737(.A(men_men_n759_), .B(men_men_n196_), .Y(men_men_n760_));
  OA210      u0738(.A0(men_men_n622_), .A1(men_men_n126_), .B0(i_13_), .Y(men_men_n761_));
  NA2        u0739(.A(men_men_n202_), .B(men_men_n205_), .Y(men_men_n762_));
  NA2        u0740(.A(men_men_n152_), .B(men_men_n600_), .Y(men_men_n763_));
  AOI210     u0741(.A0(men_men_n763_), .A1(men_men_n762_), .B0(men_men_n380_), .Y(men_men_n764_));
  AOI210     u0742(.A0(men_men_n210_), .A1(men_men_n148_), .B0(men_men_n522_), .Y(men_men_n765_));
  NA2        u0743(.A(men_men_n765_), .B(men_men_n428_), .Y(men_men_n766_));
  NO2        u0744(.A(men_men_n102_), .B(men_men_n44_), .Y(men_men_n767_));
  INV        u0745(.A(men_men_n308_), .Y(men_men_n768_));
  NA4        u0746(.A(men_men_n768_), .B(men_men_n312_), .C(men_men_n124_), .D(men_men_n42_), .Y(men_men_n769_));
  OAI210     u0747(.A0(men_men_n769_), .A1(men_men_n767_), .B0(men_men_n766_), .Y(men_men_n770_));
  NO4        u0748(.A(men_men_n770_), .B(men_men_n764_), .C(men_men_n761_), .D(men_men_n760_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n583_), .B(men_men_n28_), .Y(men_men_n772_));
  NA2        u0750(.A(men_men_n740_), .B(men_men_n282_), .Y(men_men_n773_));
  NA2        u0751(.A(men_men_n773_), .B(men_men_n772_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n62_), .B(i_12_), .Y(men_men_n775_));
  NO2        u0753(.A(men_men_n775_), .B(men_men_n126_), .Y(men_men_n776_));
  NO2        u0754(.A(men_men_n776_), .B(men_men_n600_), .Y(men_men_n777_));
  AOI220     u0755(.A0(men_men_n777_), .A1(men_men_n36_), .B0(men_men_n774_), .B1(men_men_n46_), .Y(men_men_n778_));
  NA4        u0756(.A(men_men_n778_), .B(men_men_n771_), .C(men_men_n757_), .D(men_men_n747_), .Y(men6));
  NO3        u0757(.A(i_9_), .B(men_men_n314_), .C(i_1_), .Y(men_men_n780_));
  NO2        u0758(.A(men_men_n188_), .B(men_men_n139_), .Y(men_men_n781_));
  OAI210     u0759(.A0(men_men_n781_), .A1(men_men_n780_), .B0(men_men_n728_), .Y(men_men_n782_));
  INV        u0760(.A(men_men_n337_), .Y(men_men_n783_));
  AO210      u0761(.A0(men_men_n783_), .A1(men_men_n782_), .B0(i_12_), .Y(men_men_n784_));
  NA2        u0762(.A(men_men_n589_), .B(men_men_n63_), .Y(men_men_n785_));
  NA2        u0763(.A(men_men_n685_), .B(men_men_n71_), .Y(men_men_n786_));
  NA2        u0764(.A(men_men_n786_), .B(men_men_n785_), .Y(men_men_n787_));
  NA2        u0765(.A(men_men_n787_), .B(men_men_n73_), .Y(men_men_n788_));
  INV        u0766(.A(men_men_n336_), .Y(men_men_n789_));
  NA2        u0767(.A(men_men_n75_), .B(men_men_n131_), .Y(men_men_n790_));
  NO2        u0768(.A(men_men_n790_), .B(men_men_n789_), .Y(men_men_n791_));
  NO2        u0769(.A(men_men_n255_), .B(i_9_), .Y(men_men_n792_));
  NA2        u0770(.A(men_men_n792_), .B(men_men_n775_), .Y(men_men_n793_));
  AOI210     u0771(.A0(men_men_n793_), .A1(men_men_n520_), .B0(men_men_n188_), .Y(men_men_n794_));
  NO2        u0772(.A(men_men_n32_), .B(i_11_), .Y(men_men_n795_));
  NA3        u0773(.A(men_men_n795_), .B(men_men_n476_), .C(men_men_n396_), .Y(men_men_n796_));
  NAi32      u0774(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n797_));
  NO2        u0775(.A(men_men_n717_), .B(men_men_n797_), .Y(men_men_n798_));
  OAI210     u0776(.A0(men_men_n684_), .A1(men_men_n571_), .B0(men_men_n570_), .Y(men_men_n799_));
  NAi31      u0777(.An(men_men_n798_), .B(men_men_n799_), .C(men_men_n796_), .Y(men_men_n800_));
  OR3        u0778(.A(men_men_n800_), .B(men_men_n794_), .C(men_men_n791_), .Y(men_men_n801_));
  NO2        u0779(.A(men_men_n697_), .B(i_2_), .Y(men_men_n802_));
  NA2        u0780(.A(men_men_n48_), .B(men_men_n37_), .Y(men_men_n803_));
  OAI210     u0781(.A0(men_men_n803_), .A1(men_men_n417_), .B0(men_men_n370_), .Y(men_men_n804_));
  NA2        u0782(.A(men_men_n804_), .B(men_men_n802_), .Y(men_men_n805_));
  AO210      u0783(.A0(men_men_n369_), .A1(men_men_n361_), .B0(men_men_n403_), .Y(men_men_n806_));
  NA3        u0784(.A(men_men_n806_), .B(men_men_n259_), .C(i_7_), .Y(men_men_n807_));
  NA3        u0785(.A(men_men_n454_), .B(men_men_n147_), .C(men_men_n69_), .Y(men_men_n808_));
  AO210      u0786(.A0(men_men_n494_), .A1(men_men_n744_), .B0(men_men_n36_), .Y(men_men_n809_));
  NA4        u0787(.A(men_men_n809_), .B(men_men_n808_), .C(men_men_n807_), .D(men_men_n805_), .Y(men_men_n810_));
  NO2        u0788(.A(men_men_n638_), .B(i_11_), .Y(men_men_n811_));
  NA2        u0789(.A(men_men_n811_), .B(men_men_n570_), .Y(men_men_n812_));
  NA3        u0790(.A(men_men_n380_), .B(men_men_n241_), .C(men_men_n147_), .Y(men_men_n813_));
  NA2        u0791(.A(men_men_n403_), .B(men_men_n70_), .Y(men_men_n814_));
  NA4        u0792(.A(men_men_n814_), .B(men_men_n813_), .C(men_men_n812_), .D(men_men_n606_), .Y(men_men_n815_));
  AN2        u0793(.A(men_men_n522_), .B(men_men_n46_), .Y(men_men_n816_));
  NA3        u0794(.A(men_men_n816_), .B(men_men_n485_), .C(men_men_n220_), .Y(men_men_n817_));
  AOI210     u0795(.A0(men_men_n454_), .A1(men_men_n452_), .B0(men_men_n569_), .Y(men_men_n818_));
  NA2        u0796(.A(men_men_n111_), .B(men_men_n415_), .Y(men_men_n819_));
  INV        u0797(.A(men_men_n592_), .Y(men_men_n820_));
  NA3        u0798(.A(men_men_n820_), .B(men_men_n336_), .C(i_7_), .Y(men_men_n821_));
  NA4        u0799(.A(men_men_n821_), .B(men_men_n819_), .C(men_men_n818_), .D(men_men_n817_), .Y(men_men_n822_));
  NO4        u0800(.A(men_men_n822_), .B(men_men_n815_), .C(men_men_n810_), .D(men_men_n801_), .Y(men_men_n823_));
  NA4        u0801(.A(men_men_n823_), .B(men_men_n788_), .C(men_men_n784_), .D(men_men_n386_), .Y(men3));
  NA2        u0802(.A(i_12_), .B(i_10_), .Y(men_men_n825_));
  NA2        u0803(.A(i_6_), .B(i_7_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n826_), .B(i_0_), .Y(men_men_n827_));
  NO2        u0805(.A(i_11_), .B(men_men_n239_), .Y(men_men_n828_));
  OAI210     u0806(.A0(men_men_n827_), .A1(men_men_n296_), .B0(men_men_n828_), .Y(men_men_n829_));
  NO2        u0807(.A(men_men_n829_), .B(men_men_n196_), .Y(men_men_n830_));
  NO3        u0808(.A(men_men_n458_), .B(men_men_n89_), .C(men_men_n44_), .Y(men_men_n831_));
  OA210      u0809(.A0(men_men_n831_), .A1(men_men_n830_), .B0(men_men_n176_), .Y(men_men_n832_));
  NA3        u0810(.A(men_men_n813_), .B(men_men_n606_), .C(men_men_n379_), .Y(men_men_n833_));
  NA2        u0811(.A(men_men_n833_), .B(men_men_n40_), .Y(men_men_n834_));
  NO3        u0812(.A(men_men_n630_), .B(men_men_n462_), .C(men_men_n131_), .Y(men_men_n835_));
  AN2        u0813(.A(men_men_n460_), .B(men_men_n55_), .Y(men_men_n836_));
  NO2        u0814(.A(men_men_n836_), .B(men_men_n835_), .Y(men_men_n837_));
  AOI210     u0815(.A0(men_men_n837_), .A1(men_men_n834_), .B0(men_men_n48_), .Y(men_men_n838_));
  NO4        u0816(.A(men_men_n384_), .B(men_men_n389_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n188_), .B(men_men_n579_), .Y(men_men_n840_));
  NOi21      u0818(.An(men_men_n840_), .B(men_men_n839_), .Y(men_men_n841_));
  NA2        u0819(.A(men_men_n706_), .B(men_men_n674_), .Y(men_men_n842_));
  NA2        u0820(.A(men_men_n341_), .B(men_men_n446_), .Y(men_men_n843_));
  OAI220     u0821(.A0(men_men_n843_), .A1(men_men_n842_), .B0(men_men_n841_), .B1(men_men_n63_), .Y(men_men_n844_));
  NOi21      u0822(.An(i_5_), .B(i_9_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n845_), .B(men_men_n451_), .Y(men_men_n846_));
  AOI210     u0824(.A0(men_men_n272_), .A1(men_men_n478_), .B0(men_men_n689_), .Y(men_men_n847_));
  NO3        u0825(.A(men_men_n421_), .B(men_men_n272_), .C(men_men_n73_), .Y(men_men_n848_));
  NO2        u0826(.A(men_men_n177_), .B(men_men_n148_), .Y(men_men_n849_));
  AOI210     u0827(.A0(men_men_n849_), .A1(men_men_n247_), .B0(men_men_n848_), .Y(men_men_n850_));
  OAI220     u0828(.A0(men_men_n850_), .A1(men_men_n183_), .B0(men_men_n847_), .B1(men_men_n846_), .Y(men_men_n851_));
  NO4        u0829(.A(men_men_n851_), .B(men_men_n844_), .C(men_men_n838_), .D(men_men_n832_), .Y(men_men_n852_));
  NA2        u0830(.A(men_men_n188_), .B(men_men_n24_), .Y(men_men_n853_));
  NA2        u0831(.A(men_men_n319_), .B(men_men_n129_), .Y(men_men_n854_));
  NAi21      u0832(.An(men_men_n163_), .B(men_men_n446_), .Y(men_men_n855_));
  NO2        u0833(.A(men_men_n854_), .B(men_men_n408_), .Y(men_men_n856_));
  INV        u0834(.A(men_men_n856_), .Y(men_men_n857_));
  NO2        u0835(.A(men_men_n396_), .B(men_men_n300_), .Y(men_men_n858_));
  NA2        u0836(.A(men_men_n858_), .B(men_men_n708_), .Y(men_men_n859_));
  NA2        u0837(.A(men_men_n580_), .B(i_0_), .Y(men_men_n860_));
  NO2        u0838(.A(men_men_n860_), .B(men_men_n391_), .Y(men_men_n861_));
  NO4        u0839(.A(men_men_n591_), .B(men_men_n217_), .C(men_men_n425_), .D(men_men_n417_), .Y(men_men_n862_));
  AOI210     u0840(.A0(men_men_n862_), .A1(i_11_), .B0(men_men_n861_), .Y(men_men_n863_));
  AN2        u0841(.A(men_men_n96_), .B(men_men_n246_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n740_), .B(men_men_n337_), .Y(men_men_n865_));
  INV        u0843(.A(men_men_n58_), .Y(men_men_n866_));
  OAI220     u0844(.A0(men_men_n866_), .A1(men_men_n865_), .B0(men_men_n657_), .B1(men_men_n543_), .Y(men_men_n867_));
  NO2        u0845(.A(men_men_n257_), .B(men_men_n154_), .Y(men_men_n868_));
  NA2        u0846(.A(i_0_), .B(i_10_), .Y(men_men_n869_));
  OAI210     u0847(.A0(men_men_n869_), .A1(men_men_n85_), .B0(men_men_n545_), .Y(men_men_n870_));
  NO4        u0848(.A(men_men_n114_), .B(men_men_n58_), .C(men_men_n667_), .D(i_5_), .Y(men_men_n871_));
  AO220      u0849(.A0(men_men_n871_), .A1(men_men_n870_), .B0(men_men_n868_), .B1(i_6_), .Y(men_men_n872_));
  AOI220     u0850(.A0(men_men_n341_), .A1(men_men_n98_), .B0(men_men_n188_), .B1(men_men_n83_), .Y(men_men_n873_));
  NA2        u0851(.A(men_men_n574_), .B(i_4_), .Y(men_men_n874_));
  NA2        u0852(.A(men_men_n191_), .B(men_men_n205_), .Y(men_men_n875_));
  OAI220     u0853(.A0(men_men_n875_), .A1(men_men_n865_), .B0(men_men_n874_), .B1(men_men_n873_), .Y(men_men_n876_));
  NO4        u0854(.A(men_men_n876_), .B(men_men_n872_), .C(men_men_n867_), .D(men_men_n864_), .Y(men_men_n877_));
  NA4        u0855(.A(men_men_n877_), .B(men_men_n863_), .C(men_men_n859_), .D(men_men_n857_), .Y(men_men_n878_));
  NO2        u0856(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n879_));
  NA2        u0857(.A(i_11_), .B(i_9_), .Y(men_men_n880_));
  NO3        u0858(.A(i_12_), .B(men_men_n880_), .C(men_men_n605_), .Y(men_men_n881_));
  AN2        u0859(.A(men_men_n881_), .B(men_men_n879_), .Y(men_men_n882_));
  NO2        u0860(.A(men_men_n48_), .B(i_7_), .Y(men_men_n883_));
  NA2        u0861(.A(men_men_n400_), .B(men_men_n181_), .Y(men_men_n884_));
  NA2        u0862(.A(men_men_n884_), .B(men_men_n161_), .Y(men_men_n885_));
  NO2        u0863(.A(men_men_n880_), .B(men_men_n73_), .Y(men_men_n886_));
  NO2        u0864(.A(men_men_n177_), .B(i_0_), .Y(men_men_n887_));
  INV        u0865(.A(men_men_n887_), .Y(men_men_n888_));
  NA2        u0866(.A(men_men_n476_), .B(men_men_n233_), .Y(men_men_n889_));
  NO2        u0867(.A(men_men_n889_), .B(men_men_n888_), .Y(men_men_n890_));
  NO3        u0868(.A(men_men_n890_), .B(men_men_n885_), .C(men_men_n882_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n656_), .B(men_men_n121_), .Y(men_men_n892_));
  NO2        u0870(.A(i_6_), .B(men_men_n892_), .Y(men_men_n893_));
  AOI210     u0871(.A0(men_men_n453_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n894_));
  NA2        u0872(.A(men_men_n173_), .B(men_men_n103_), .Y(men_men_n895_));
  NOi32      u0873(.An(men_men_n894_), .Bn(men_men_n191_), .C(men_men_n895_), .Y(men_men_n896_));
  NO2        u0874(.A(men_men_n896_), .B(men_men_n893_), .Y(men_men_n897_));
  NOi21      u0875(.An(i_7_), .B(i_5_), .Y(men_men_n898_));
  NOi31      u0876(.An(men_men_n898_), .B(i_0_), .C(men_men_n720_), .Y(men_men_n899_));
  NA3        u0877(.A(men_men_n899_), .B(men_men_n390_), .C(i_6_), .Y(men_men_n900_));
  OA210      u0878(.A0(men_men_n895_), .A1(men_men_n520_), .B0(men_men_n900_), .Y(men_men_n901_));
  NO3        u0879(.A(men_men_n411_), .B(men_men_n372_), .C(men_men_n368_), .Y(men_men_n902_));
  NO2        u0880(.A(men_men_n266_), .B(men_men_n326_), .Y(men_men_n903_));
  NO2        u0881(.A(men_men_n720_), .B(men_men_n261_), .Y(men_men_n904_));
  AOI210     u0882(.A0(men_men_n904_), .A1(men_men_n903_), .B0(men_men_n902_), .Y(men_men_n905_));
  NA4        u0883(.A(men_men_n905_), .B(men_men_n901_), .C(men_men_n897_), .D(men_men_n891_), .Y(men_men_n906_));
  NO2        u0884(.A(men_men_n853_), .B(men_men_n242_), .Y(men_men_n907_));
  AN2        u0885(.A(men_men_n340_), .B(men_men_n337_), .Y(men_men_n908_));
  AN2        u0886(.A(men_men_n908_), .B(men_men_n849_), .Y(men_men_n909_));
  OAI210     u0887(.A0(men_men_n909_), .A1(men_men_n907_), .B0(i_10_), .Y(men_men_n910_));
  NO2        u0888(.A(men_men_n825_), .B(men_men_n325_), .Y(men_men_n911_));
  NA2        u0889(.A(men_men_n911_), .B(men_men_n886_), .Y(men_men_n912_));
  NA3        u0890(.A(men_men_n475_), .B(men_men_n418_), .C(men_men_n45_), .Y(men_men_n913_));
  OAI210     u0891(.A0(men_men_n855_), .A1(i_6_), .B0(men_men_n913_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n259_), .B(men_men_n46_), .Y(men_men_n915_));
  NO2        u0893(.A(men_men_n915_), .B(men_men_n190_), .Y(men_men_n916_));
  AOI220     u0894(.A0(men_men_n916_), .A1(men_men_n476_), .B0(men_men_n914_), .B1(men_men_n73_), .Y(men_men_n917_));
  NA3        u0895(.A(men_men_n803_), .B(men_men_n388_), .C(men_men_n638_), .Y(men_men_n918_));
  NA2        u0896(.A(men_men_n92_), .B(men_men_n44_), .Y(men_men_n919_));
  NO2        u0897(.A(men_men_n75_), .B(men_men_n742_), .Y(men_men_n920_));
  AOI220     u0898(.A0(men_men_n920_), .A1(men_men_n919_), .B0(men_men_n176_), .B1(men_men_n599_), .Y(men_men_n921_));
  AOI210     u0899(.A0(men_men_n921_), .A1(men_men_n918_), .B0(men_men_n47_), .Y(men_men_n922_));
  NO3        u0900(.A(men_men_n591_), .B(men_men_n367_), .C(men_men_n24_), .Y(men_men_n923_));
  AOI210     u0901(.A0(men_men_n700_), .A1(men_men_n554_), .B0(men_men_n923_), .Y(men_men_n924_));
  NO2        u0902(.A(men_men_n601_), .B(men_men_n105_), .Y(men_men_n925_));
  NA2        u0903(.A(men_men_n925_), .B(i_0_), .Y(men_men_n926_));
  OAI220     u0904(.A0(men_men_n926_), .A1(men_men_n85_), .B0(men_men_n924_), .B1(men_men_n174_), .Y(men_men_n927_));
  NO3        u0905(.A(men_men_n927_), .B(men_men_n922_), .C(men_men_n525_), .Y(men_men_n928_));
  NA4        u0906(.A(men_men_n928_), .B(men_men_n917_), .C(men_men_n912_), .D(men_men_n910_), .Y(men_men_n929_));
  NO3        u0907(.A(men_men_n929_), .B(men_men_n906_), .C(men_men_n878_), .Y(men_men_n930_));
  NO2        u0908(.A(i_0_), .B(men_men_n720_), .Y(men_men_n931_));
  NA2        u0909(.A(men_men_n73_), .B(men_men_n44_), .Y(men_men_n932_));
  NA2        u0910(.A(men_men_n869_), .B(men_men_n932_), .Y(men_men_n933_));
  NO3        u0911(.A(men_men_n105_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n934_));
  AO220      u0912(.A0(men_men_n934_), .A1(men_men_n933_), .B0(men_men_n931_), .B1(men_men_n176_), .Y(men_men_n935_));
  AOI210     u0913(.A0(men_men_n785_), .A1(men_men_n687_), .B0(men_men_n895_), .Y(men_men_n936_));
  AOI210     u0914(.A0(men_men_n935_), .A1(men_men_n358_), .B0(men_men_n936_), .Y(men_men_n937_));
  NA2        u0915(.A(men_men_n728_), .B(men_men_n146_), .Y(men_men_n938_));
  INV        u0916(.A(men_men_n938_), .Y(men_men_n939_));
  NA3        u0917(.A(men_men_n939_), .B(men_men_n674_), .C(men_men_n73_), .Y(men_men_n940_));
  NO2        u0918(.A(men_men_n799_), .B(men_men_n411_), .Y(men_men_n941_));
  NA3        u0919(.A(men_men_n827_), .B(i_2_), .C(men_men_n48_), .Y(men_men_n942_));
  NA2        u0920(.A(men_men_n828_), .B(i_9_), .Y(men_men_n943_));
  AOI210     u0921(.A0(men_men_n942_), .A1(men_men_n500_), .B0(men_men_n943_), .Y(men_men_n944_));
  NA2        u0922(.A(men_men_n247_), .B(men_men_n232_), .Y(men_men_n945_));
  AOI210     u0923(.A0(men_men_n945_), .A1(men_men_n860_), .B0(men_men_n154_), .Y(men_men_n946_));
  NO3        u0924(.A(men_men_n946_), .B(men_men_n944_), .C(men_men_n941_), .Y(men_men_n947_));
  NA3        u0925(.A(men_men_n947_), .B(men_men_n940_), .C(men_men_n937_), .Y(men_men_n948_));
  NA2        u0926(.A(men_men_n908_), .B(men_men_n380_), .Y(men_men_n949_));
  AOI210     u0927(.A0(men_men_n307_), .A1(men_men_n163_), .B0(men_men_n949_), .Y(men_men_n950_));
  NA3        u0928(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n44_), .Y(men_men_n951_));
  NA2        u0929(.A(men_men_n883_), .B(men_men_n489_), .Y(men_men_n952_));
  AOI210     u0930(.A0(men_men_n951_), .A1(men_men_n163_), .B0(men_men_n952_), .Y(men_men_n953_));
  NO2        u0931(.A(men_men_n953_), .B(men_men_n950_), .Y(men_men_n954_));
  NO3        u0932(.A(men_men_n869_), .B(men_men_n845_), .C(men_men_n193_), .Y(men_men_n955_));
  AOI220     u0933(.A0(men_men_n955_), .A1(i_11_), .B0(men_men_n575_), .B1(men_men_n75_), .Y(men_men_n956_));
  NO3        u0934(.A(men_men_n211_), .B(men_men_n389_), .C(i_0_), .Y(men_men_n957_));
  OAI210     u0935(.A0(men_men_n957_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n958_));
  INV        u0936(.A(men_men_n220_), .Y(men_men_n959_));
  OAI220     u0937(.A0(men_men_n536_), .A1(men_men_n139_), .B0(men_men_n643_), .B1(men_men_n616_), .Y(men_men_n960_));
  NA3        u0938(.A(men_men_n960_), .B(i_7_), .C(men_men_n959_), .Y(men_men_n961_));
  NA4        u0939(.A(men_men_n961_), .B(men_men_n958_), .C(men_men_n956_), .D(men_men_n954_), .Y(men_men_n962_));
  NO2        u0940(.A(men_men_n245_), .B(men_men_n92_), .Y(men_men_n963_));
  NA2        u0941(.A(men_men_n963_), .B(men_men_n931_), .Y(men_men_n964_));
  AOI220     u0942(.A0(men_men_n898_), .A1(men_men_n489_), .B0(men_men_n827_), .B1(men_men_n164_), .Y(men_men_n965_));
  NA2        u0943(.A(men_men_n361_), .B(men_men_n178_), .Y(men_men_n966_));
  OA220      u0944(.A0(men_men_n966_), .A1(men_men_n965_), .B0(men_men_n964_), .B1(i_5_), .Y(men_men_n967_));
  AOI210     u0945(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n177_), .Y(men_men_n968_));
  NA3        u0946(.A(men_men_n613_), .B(men_men_n188_), .C(men_men_n83_), .Y(men_men_n969_));
  NA2        u0947(.A(men_men_n969_), .B(men_men_n552_), .Y(men_men_n970_));
  INV        u0948(.A(men_men_n970_), .Y(men_men_n971_));
  NA3        u0949(.A(men_men_n396_), .B(men_men_n342_), .C(men_men_n223_), .Y(men_men_n972_));
  INV        u0950(.A(men_men_n972_), .Y(men_men_n973_));
  NOi31      u0951(.An(men_men_n395_), .B(men_men_n932_), .C(men_men_n242_), .Y(men_men_n974_));
  NO2        u0952(.A(men_men_n974_), .B(men_men_n973_), .Y(men_men_n975_));
  NA3        u0953(.A(men_men_n975_), .B(men_men_n971_), .C(men_men_n967_), .Y(men_men_n976_));
  INV        u0954(.A(men_men_n615_), .Y(men_men_n977_));
  NO3        u0955(.A(men_men_n977_), .B(men_men_n567_), .C(men_men_n355_), .Y(men_men_n978_));
  NO2        u0956(.A(men_men_n85_), .B(i_5_), .Y(men_men_n979_));
  NA3        u0957(.A(men_men_n828_), .B(men_men_n109_), .C(men_men_n124_), .Y(men_men_n980_));
  INV        u0958(.A(men_men_n980_), .Y(men_men_n981_));
  AOI210     u0959(.A0(men_men_n981_), .A1(men_men_n979_), .B0(men_men_n978_), .Y(men_men_n982_));
  NA3        u0960(.A(men_men_n312_), .B(i_5_), .C(men_men_n196_), .Y(men_men_n983_));
  NAi31      u0961(.An(men_men_n244_), .B(men_men_n983_), .C(men_men_n245_), .Y(men_men_n984_));
  NO4        u0962(.A(men_men_n242_), .B(men_men_n211_), .C(i_0_), .D(i_12_), .Y(men_men_n985_));
  NA2        u0963(.A(men_men_n985_), .B(men_men_n984_), .Y(men_men_n986_));
  AN2        u0964(.A(men_men_n869_), .B(men_men_n154_), .Y(men_men_n987_));
  NO4        u0965(.A(men_men_n987_), .B(i_12_), .C(men_men_n647_), .D(men_men_n131_), .Y(men_men_n988_));
  NA2        u0966(.A(men_men_n988_), .B(men_men_n220_), .Y(men_men_n989_));
  NA3        u0967(.A(men_men_n98_), .B(men_men_n579_), .C(i_11_), .Y(men_men_n990_));
  NO2        u0968(.A(men_men_n990_), .B(men_men_n156_), .Y(men_men_n991_));
  NO2        u0969(.A(i_7_), .B(men_men_n983_), .Y(men_men_n992_));
  AOI210     u0970(.A0(men_men_n992_), .A1(men_men_n887_), .B0(men_men_n991_), .Y(men_men_n993_));
  NA4        u0971(.A(men_men_n993_), .B(men_men_n989_), .C(men_men_n986_), .D(men_men_n982_), .Y(men_men_n994_));
  NO4        u0972(.A(men_men_n994_), .B(men_men_n976_), .C(men_men_n962_), .D(men_men_n948_), .Y(men_men_n995_));
  OAI210     u0973(.A0(men_men_n802_), .A1(men_men_n795_), .B0(men_men_n37_), .Y(men_men_n996_));
  NA3        u0974(.A(men_men_n894_), .B(men_men_n375_), .C(i_5_), .Y(men_men_n997_));
  NA3        u0975(.A(men_men_n997_), .B(men_men_n996_), .C(men_men_n1043_), .Y(men_men_n998_));
  NA2        u0976(.A(men_men_n998_), .B(men_men_n208_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n189_), .B(men_men_n191_), .Y(men_men_n1000_));
  AO210      u0978(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  OAI210     u0979(.A0(men_men_n615_), .A1(men_men_n613_), .B0(men_men_n325_), .Y(men_men_n1002_));
  NAi31      u0980(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1003_));
  AOI210     u0981(.A0(men_men_n117_), .A1(men_men_n70_), .B0(men_men_n1003_), .Y(men_men_n1004_));
  NO2        u0982(.A(men_men_n1004_), .B(men_men_n644_), .Y(men_men_n1005_));
  NA3        u0983(.A(men_men_n1005_), .B(men_men_n1002_), .C(men_men_n1001_), .Y(men_men_n1006_));
  NO2        u0984(.A(men_men_n465_), .B(men_men_n272_), .Y(men_men_n1007_));
  NO4        u0985(.A(men_men_n235_), .B(men_men_n145_), .C(men_men_n678_), .D(men_men_n37_), .Y(men_men_n1008_));
  NO3        u0986(.A(men_men_n1008_), .B(men_men_n1007_), .C(men_men_n862_), .Y(men_men_n1009_));
  OAI210     u0987(.A0(men_men_n990_), .A1(men_men_n148_), .B0(men_men_n1009_), .Y(men_men_n1010_));
  AOI210     u0988(.A0(men_men_n1006_), .A1(men_men_n48_), .B0(men_men_n1010_), .Y(men_men_n1011_));
  AOI210     u0989(.A0(men_men_n1011_), .A1(men_men_n999_), .B0(men_men_n73_), .Y(men_men_n1012_));
  INV        u0990(.A(men_men_n572_), .Y(men_men_n1013_));
  NO2        u0991(.A(men_men_n1013_), .B(men_men_n748_), .Y(men_men_n1014_));
  OAI210     u0992(.A0(men_men_n80_), .A1(men_men_n54_), .B0(men_men_n108_), .Y(men_men_n1015_));
  NA2        u0993(.A(men_men_n1015_), .B(men_men_n76_), .Y(men_men_n1016_));
  AOI210     u0994(.A0(men_men_n968_), .A1(men_men_n883_), .B0(men_men_n899_), .Y(men_men_n1017_));
  AOI210     u0995(.A0(men_men_n1017_), .A1(men_men_n1016_), .B0(men_men_n678_), .Y(men_men_n1018_));
  NA2        u0996(.A(men_men_n266_), .B(men_men_n57_), .Y(men_men_n1019_));
  NA2        u0997(.A(men_men_n1019_), .B(men_men_n76_), .Y(men_men_n1020_));
  NO2        u0998(.A(men_men_n1020_), .B(men_men_n239_), .Y(men_men_n1021_));
  NA3        u0999(.A(men_men_n96_), .B(men_men_n314_), .C(men_men_n31_), .Y(men_men_n1022_));
  INV        u1000(.A(men_men_n1022_), .Y(men_men_n1023_));
  NO3        u1001(.A(men_men_n1023_), .B(men_men_n1021_), .C(men_men_n1018_), .Y(men_men_n1024_));
  OAI210     u1002(.A0(men_men_n274_), .A1(men_men_n159_), .B0(men_men_n86_), .Y(men_men_n1025_));
  NA3        u1003(.A(men_men_n752_), .B(men_men_n296_), .C(men_men_n80_), .Y(men_men_n1026_));
  AOI210     u1004(.A0(men_men_n1026_), .A1(men_men_n1025_), .B0(i_11_), .Y(men_men_n1027_));
  OAI210     u1005(.A0(men_men_n1042_), .A1(men_men_n894_), .B0(men_men_n208_), .Y(men_men_n1028_));
  NA2        u1006(.A(men_men_n165_), .B(i_5_), .Y(men_men_n1029_));
  NO2        u1007(.A(men_men_n1028_), .B(men_men_n1029_), .Y(men_men_n1030_));
  NO3        u1008(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1031_));
  OAI210     u1009(.A0(men_men_n903_), .A1(men_men_n314_), .B0(men_men_n1031_), .Y(men_men_n1032_));
  NO2        u1010(.A(men_men_n1032_), .B(men_men_n720_), .Y(men_men_n1033_));
  NO3        u1011(.A(men_men_n1033_), .B(men_men_n1030_), .C(men_men_n1027_), .Y(men_men_n1034_));
  OAI210     u1012(.A0(men_men_n1024_), .A1(i_4_), .B0(men_men_n1034_), .Y(men_men_n1035_));
  NO3        u1013(.A(men_men_n1035_), .B(men_men_n1014_), .C(men_men_n1012_), .Y(men_men_n1036_));
  NA4        u1014(.A(men_men_n1036_), .B(men_men_n995_), .C(men_men_n930_), .D(men_men_n852_), .Y(men4));
  INV        u1015(.A(i_2_), .Y(men_men_n1040_));
  INV        u1016(.A(i_12_), .Y(men_men_n1041_));
  INV        u1017(.A(i_12_), .Y(men_men_n1042_));
  INV        u1018(.A(men_men_n162_), .Y(men_men_n1043_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule