//Benchmark atmr_misex3_1774_0.125

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1045_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1092_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1118_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1161_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1226_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1291_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1340_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1059_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1101_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1124_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1178_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1244_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1314_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1370_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1573_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1582_, men_men_n1583_, men_men_n1585_, men_men_n1586_, men_men_n1587_, men_men_n1588_, men_men_n1589_, men_men_n1590_, men_men_n1591_, men_men_n1595_, men_men_n1596_, men_men_n1597_, men_men_n1598_, men_men_n1599_, men_men_n1600_, men_men_n1601_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o000(.A(j), .B(g), .Y(ori_ori_n29_));
  INV        o001(.A(i), .Y(ori_ori_n30_));
  NAi21      o002(.An(n), .B(m), .Y(ori_ori_n31_));
  NOi32      o003(.An(k), .Bn(h), .C(l), .Y(ori_ori_n32_));
  AN2        o004(.A(k), .B(h), .Y(ori_ori_n33_));
  INV        o005(.A(c), .Y(ori_ori_n34_));
  INV        o006(.A(d), .Y(ori_ori_n35_));
  NAi21      o007(.An(i), .B(h), .Y(ori_ori_n36_));
  INV        o008(.A(f), .Y(ori_ori_n37_));
  INV        o009(.A(m), .Y(ori_ori_n38_));
  INV        o010(.A(n), .Y(ori_ori_n39_));
  INV        o011(.A(j), .Y(ori_ori_n40_));
  NAi41      o012(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n41_));
  AN2        o013(.A(e), .B(b), .Y(ori_ori_n42_));
  NOi21      o014(.An(i), .B(h), .Y(ori_ori_n43_));
  INV        o015(.A(a), .Y(ori_ori_n44_));
  NA2        o016(.A(ori_ori_n42_), .B(ori_ori_n44_), .Y(ori_ori_n45_));
  NOi21      o017(.An(m), .B(n), .Y(ori_ori_n46_));
  AN2        o018(.A(k), .B(h), .Y(ori_ori_n47_));
  INV        o019(.A(b), .Y(ori_ori_n48_));
  AN2        o020(.A(k), .B(i), .Y(ori_ori_n49_));
  NOi32      o021(.An(f), .Bn(b), .C(e), .Y(ori_ori_n50_));
  NAi21      o022(.An(m), .B(n), .Y(ori_ori_n51_));
  NAi31      o023(.An(j), .B(k), .C(h), .Y(ori_ori_n52_));
  NAi21      o024(.An(e), .B(f), .Y(ori_ori_n53_));
  NAi21      o025(.An(c), .B(d), .Y(ori_ori_n54_));
  NOi21      o026(.An(h), .B(i), .Y(ori_ori_n55_));
  NOi21      o027(.An(k), .B(m), .Y(ori_ori_n56_));
  NA3        o028(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(n), .Y(ori_ori_n57_));
  NAi31      o029(.An(d), .B(f), .C(c), .Y(ori_ori_n58_));
  NAi31      o030(.An(e), .B(f), .C(c), .Y(ori_ori_n59_));
  NA2        o031(.A(ori_ori_n59_), .B(ori_ori_n58_), .Y(ori_ori_n60_));
  NA2        o032(.A(j), .B(h), .Y(ori_ori_n61_));
  OR3        o033(.A(n), .B(m), .C(k), .Y(ori_ori_n62_));
  NO2        o034(.A(ori_ori_n62_), .B(ori_ori_n61_), .Y(ori_ori_n63_));
  NAi32      o035(.An(m), .Bn(k), .C(n), .Y(ori_ori_n64_));
  NA2        o036(.A(ori_ori_n63_), .B(ori_ori_n60_), .Y(ori_ori_n65_));
  NO2        o037(.A(n), .B(m), .Y(ori_ori_n66_));
  NA2        o038(.A(ori_ori_n66_), .B(ori_ori_n32_), .Y(ori_ori_n67_));
  NAi21      o039(.An(f), .B(e), .Y(ori_ori_n68_));
  NA2        o040(.A(d), .B(c), .Y(ori_ori_n69_));
  NAi21      o041(.An(h), .B(f), .Y(ori_ori_n70_));
  NOi32      o042(.An(f), .Bn(c), .C(d), .Y(ori_ori_n71_));
  NOi32      o043(.An(f), .Bn(c), .C(e), .Y(ori_ori_n72_));
  NO2        o044(.A(ori_ori_n72_), .B(ori_ori_n71_), .Y(ori_ori_n73_));
  NO3        o045(.A(n), .B(m), .C(j), .Y(ori_ori_n74_));
  NA2        o046(.A(ori_ori_n74_), .B(ori_ori_n47_), .Y(ori_ori_n75_));
  AO210      o047(.A0(ori_ori_n75_), .A1(ori_ori_n67_), .B0(ori_ori_n73_), .Y(ori_ori_n76_));
  NA2        o048(.A(ori_ori_n76_), .B(ori_ori_n65_), .Y(ori_ori_n77_));
  INV        o049(.A(ori_ori_n77_), .Y(ori_ori_n78_));
  NAi31      o050(.An(n), .B(h), .C(g), .Y(ori_ori_n79_));
  BUFFER     o051(.A(k), .Y(ori_ori_n80_));
  NA3        o052(.A(ori_ori_n80_), .B(ori_ori_n46_), .C(g), .Y(ori_ori_n81_));
  INV        o053(.A(f), .Y(ori_ori_n82_));
  INV        o054(.A(g), .Y(ori_ori_n83_));
  NOi21      o055(.An(n), .B(m), .Y(ori_ori_n84_));
  NAi21      o056(.An(j), .B(h), .Y(ori_ori_n85_));
  XN2        o057(.A(i), .B(h), .Y(ori_ori_n86_));
  NA2        o058(.A(ori_ori_n86_), .B(ori_ori_n85_), .Y(ori_ori_n87_));
  NOi31      o059(.An(k), .B(n), .C(m), .Y(ori_ori_n88_));
  NOi31      o060(.An(ori_ori_n88_), .B(ori_ori_n69_), .C(ori_ori_n68_), .Y(ori_ori_n89_));
  NA2        o061(.A(ori_ori_n89_), .B(ori_ori_n87_), .Y(ori_ori_n90_));
  NAi31      o062(.An(f), .B(e), .C(c), .Y(ori_ori_n91_));
  NO4        o063(.A(ori_ori_n91_), .B(ori_ori_n62_), .C(ori_ori_n61_), .D(ori_ori_n35_), .Y(ori_ori_n92_));
  NAi32      o064(.An(m), .Bn(i), .C(k), .Y(ori_ori_n93_));
  INV        o065(.A(k), .Y(ori_ori_n94_));
  INV        o066(.A(ori_ori_n92_), .Y(ori_ori_n95_));
  NA3        o067(.A(m), .B(k), .C(h), .Y(ori_ori_n96_));
  AN2        o068(.A(ori_ori_n95_), .B(ori_ori_n90_), .Y(ori_ori_n97_));
  NO2        o069(.A(g), .B(ori_ori_n41_), .Y(ori_ori_n98_));
  NA2        o070(.A(ori_ori_n98_), .B(ori_ori_n50_), .Y(ori_ori_n99_));
  NA2        o071(.A(ori_ori_n56_), .B(ori_ori_n43_), .Y(ori_ori_n100_));
  INV        o072(.A(n), .Y(ori_ori_n101_));
  NAi31      o073(.An(ori_ori_n96_), .B(ori_ori_n101_), .C(ori_ori_n42_), .Y(ori_ori_n102_));
  NAi21      o074(.An(h), .B(i), .Y(ori_ori_n103_));
  NA2        o075(.A(ori_ori_n66_), .B(k), .Y(ori_ori_n104_));
  NO2        o076(.A(ori_ori_n104_), .B(ori_ori_n103_), .Y(ori_ori_n105_));
  NA2        o077(.A(ori_ori_n105_), .B(ori_ori_n71_), .Y(ori_ori_n106_));
  NA3        o078(.A(ori_ori_n106_), .B(ori_ori_n102_), .C(ori_ori_n99_), .Y(ori_ori_n107_));
  NOi21      o079(.An(ori_ori_n97_), .B(ori_ori_n107_), .Y(ori_ori_n108_));
  NA2        o080(.A(k), .B(h), .Y(ori_ori_n109_));
  NA3        o081(.A(ori_ori_n56_), .B(ori_ori_n55_), .C(ori_ori_n39_), .Y(ori_ori_n110_));
  NO2        o082(.A(ori_ori_n110_), .B(ori_ori_n73_), .Y(ori_ori_n111_));
  NA3        o083(.A(e), .B(c), .C(b), .Y(ori_ori_n112_));
  NAi21      o084(.An(m), .B(l), .Y(ori_ori_n113_));
  NAi32      o085(.An(n), .Bn(m), .C(l), .Y(ori_ori_n114_));
  INV        o086(.A(ori_ori_n111_), .Y(ori_ori_n115_));
  NA2        o087(.A(ori_ori_n105_), .B(ori_ori_n72_), .Y(ori_ori_n116_));
  NAi21      o088(.An(m), .B(k), .Y(ori_ori_n117_));
  NA2        o089(.A(e), .B(c), .Y(ori_ori_n118_));
  NO3        o090(.A(ori_ori_n118_), .B(n), .C(d), .Y(ori_ori_n119_));
  NOi31      o091(.An(l), .B(n), .C(m), .Y(ori_ori_n120_));
  NAi32      o092(.An(m), .Bn(j), .C(k), .Y(ori_ori_n121_));
  AN2        o093(.A(e), .B(b), .Y(ori_ori_n122_));
  NA2        o094(.A(ori_ori_n33_), .B(ori_ori_n46_), .Y(ori_ori_n123_));
  NA4        o095(.A(ori_ori_n116_), .B(ori_ori_n115_), .C(ori_ori_n108_), .D(ori_ori_n78_), .Y(ori10));
  NAi31      o096(.An(b), .B(f), .C(c), .Y(ori_ori_n125_));
  INV        o097(.A(ori_ori_n125_), .Y(ori_ori_n126_));
  NOi32      o098(.An(k), .Bn(h), .C(j), .Y(ori_ori_n127_));
  NA2        o099(.A(ori_ori_n127_), .B(ori_ori_n84_), .Y(ori_ori_n128_));
  NA2        o100(.A(ori_ori_n57_), .B(ori_ori_n128_), .Y(ori_ori_n129_));
  NA2        o101(.A(ori_ori_n129_), .B(ori_ori_n126_), .Y(ori_ori_n130_));
  AN2        o102(.A(j), .B(h), .Y(ori_ori_n131_));
  NO3        o103(.A(n), .B(m), .C(k), .Y(ori_ori_n132_));
  NA2        o104(.A(ori_ori_n132_), .B(ori_ori_n131_), .Y(ori_ori_n133_));
  NO3        o105(.A(ori_ori_n133_), .B(ori_ori_n54_), .C(ori_ori_n82_), .Y(ori_ori_n134_));
  OR2        o106(.A(m), .B(k), .Y(ori_ori_n135_));
  NO2        o107(.A(ori_ori_n61_), .B(ori_ori_n135_), .Y(ori_ori_n136_));
  NA4        o108(.A(n), .B(f), .C(c), .D(ori_ori_n48_), .Y(ori_ori_n137_));
  NOi21      o109(.An(ori_ori_n136_), .B(ori_ori_n137_), .Y(ori_ori_n138_));
  NO2        o110(.A(ori_ori_n138_), .B(ori_ori_n134_), .Y(ori_ori_n139_));
  NO2        o111(.A(ori_ori_n137_), .B(ori_ori_n113_), .Y(ori_ori_n140_));
  NOi32      o112(.An(f), .Bn(d), .C(c), .Y(ori_ori_n141_));
  NA2        o113(.A(ori_ori_n139_), .B(ori_ori_n130_), .Y(ori_ori_n142_));
  INV        o114(.A(e), .Y(ori_ori_n143_));
  INV        o115(.A(ori_ori_n142_), .Y(ori_ori_n144_));
  OR2        o116(.A(n), .B(m), .Y(ori_ori_n145_));
  NO2        o117(.A(ori_ori_n69_), .B(ori_ori_n53_), .Y(ori_ori_n146_));
  NA2        o118(.A(ori_ori_n63_), .B(ori_ori_n146_), .Y(ori_ori_n147_));
  INV        o119(.A(ori_ori_n123_), .Y(ori_ori_n148_));
  NA3        o120(.A(ori_ori_n148_), .B(ori_ori_n122_), .C(d), .Y(ori_ori_n149_));
  NAi21      o121(.An(k), .B(j), .Y(ori_ori_n150_));
  NAi21      o122(.An(e), .B(d), .Y(ori_ori_n151_));
  INV        o123(.A(ori_ori_n151_), .Y(ori_ori_n152_));
  NO2        o124(.A(ori_ori_n104_), .B(ori_ori_n82_), .Y(ori_ori_n153_));
  NA3        o125(.A(ori_ori_n153_), .B(ori_ori_n152_), .C(ori_ori_n87_), .Y(ori_ori_n154_));
  NA3        o126(.A(ori_ori_n154_), .B(ori_ori_n149_), .C(ori_ori_n147_), .Y(ori_ori_n155_));
  NOi31      o127(.An(n), .B(m), .C(k), .Y(ori_ori_n156_));
  AOI220     o128(.A0(ori_ori_n156_), .A1(ori_ori_n131_), .B0(ori_ori_n84_), .B1(ori_ori_n32_), .Y(ori_ori_n157_));
  NAi31      o129(.An(g), .B(f), .C(c), .Y(ori_ori_n158_));
  INV        o130(.A(ori_ori_n155_), .Y(ori_ori_n159_));
  AN2        o131(.A(e), .B(d), .Y(ori_ori_n160_));
  NO2        o132(.A(ori_ori_n37_), .B(e), .Y(ori_ori_n161_));
  NO4        o133(.A(ori_ori_n70_), .B(ori_ori_n41_), .C(ori_ori_n34_), .D(b), .Y(ori_ori_n162_));
  INV        o134(.A(ori_ori_n97_), .Y(ori_ori_n163_));
  XO2        o135(.A(i), .B(h), .Y(ori_ori_n164_));
  NA3        o136(.A(ori_ori_n164_), .B(ori_ori_n56_), .C(n), .Y(ori_ori_n165_));
  NA3        o137(.A(ori_ori_n165_), .B(ori_ori_n157_), .C(ori_ori_n128_), .Y(ori_ori_n166_));
  NOi32      o138(.An(ori_ori_n166_), .Bn(ori_ori_n161_), .C(ori_ori_n388_), .Y(ori_ori_n167_));
  NAi31      o139(.An(c), .B(f), .C(d), .Y(ori_ori_n168_));
  AOI210     o140(.A0(ori_ori_n110_), .A1(ori_ori_n75_), .B0(ori_ori_n168_), .Y(ori_ori_n169_));
  INV        o141(.A(ori_ori_n169_), .Y(ori_ori_n170_));
  NA2        o142(.A(ori_ori_n88_), .B(ori_ori_n43_), .Y(ori_ori_n171_));
  AOI210     o143(.A0(ori_ori_n171_), .A1(ori_ori_n67_), .B0(ori_ori_n168_), .Y(ori_ori_n172_));
  INV        o144(.A(ori_ori_n172_), .Y(ori_ori_n173_));
  NA2        o145(.A(ori_ori_n173_), .B(ori_ori_n170_), .Y(ori_ori_n174_));
  NO3        o146(.A(ori_ori_n174_), .B(ori_ori_n167_), .C(ori_ori_n163_), .Y(ori_ori_n175_));
  NA4        o147(.A(ori_ori_n175_), .B(ori_ori_n389_), .C(ori_ori_n159_), .D(ori_ori_n144_), .Y(ori11));
  NAi31      o148(.An(n), .B(m), .C(k), .Y(ori_ori_n177_));
  NO2        o149(.A(ori_ori_n109_), .B(ori_ori_n31_), .Y(ori_ori_n178_));
  INV        o150(.A(k), .Y(ori_ori_n179_));
  NO3        o151(.A(ori_ori_n117_), .B(ori_ori_n36_), .C(n), .Y(ori_ori_n180_));
  NA3        o152(.A(ori_ori_n168_), .B(ori_ori_n59_), .C(ori_ori_n58_), .Y(ori_ori_n181_));
  NA2        o153(.A(ori_ori_n158_), .B(ori_ori_n91_), .Y(ori_ori_n182_));
  OR2        o154(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n183_));
  NA2        o155(.A(ori_ori_n183_), .B(ori_ori_n180_), .Y(ori_ori_n184_));
  NO2        o156(.A(ori_ori_n184_), .B(ori_ori_n40_), .Y(ori_ori_n185_));
  NOi32      o157(.An(e), .Bn(c), .C(f), .Y(ori_ori_n186_));
  NA2        o158(.A(ori_ori_n186_), .B(ori_ori_n63_), .Y(ori_ori_n187_));
  NA2        o159(.A(ori_ori_n187_), .B(ori_ori_n65_), .Y(ori_ori_n188_));
  NOi31      o160(.An(m), .B(n), .C(k), .Y(ori_ori_n189_));
  NA2        o161(.A(ori_ori_n164_), .B(ori_ori_n56_), .Y(ori_ori_n190_));
  NO3        o162(.A(ori_ori_n137_), .B(ori_ori_n190_), .C(ori_ori_n40_), .Y(ori_ori_n191_));
  INV        o163(.A(ori_ori_n191_), .Y(ori_ori_n192_));
  AN3        o164(.A(f), .B(d), .C(b), .Y(ori_ori_n193_));
  OAI210     o165(.A0(ori_ori_n193_), .A1(ori_ori_n50_), .B0(n), .Y(ori_ori_n194_));
  NA3        o166(.A(ori_ori_n164_), .B(ori_ori_n56_), .C(ori_ori_n83_), .Y(ori_ori_n195_));
  NO2        o167(.A(ori_ori_n194_), .B(ori_ori_n195_), .Y(ori_ori_n196_));
  INV        o168(.A(ori_ori_n102_), .Y(ori_ori_n197_));
  OAI210     o169(.A0(ori_ori_n197_), .A1(ori_ori_n196_), .B0(j), .Y(ori_ori_n198_));
  NA2        o170(.A(ori_ori_n198_), .B(ori_ori_n192_), .Y(ori_ori_n199_));
  NO3        o171(.A(ori_ori_n199_), .B(ori_ori_n188_), .C(ori_ori_n185_), .Y(ori_ori_n200_));
  NA2        o172(.A(h), .B(f), .Y(ori_ori_n201_));
  NO3        o173(.A(g), .B(ori_ori_n82_), .C(ori_ori_n34_), .Y(ori_ori_n202_));
  NA2        o174(.A(ori_ori_n136_), .B(ori_ori_n202_), .Y(ori_ori_n203_));
  BUFFER     o175(.A(h), .Y(ori_ori_n204_));
  NA2        o176(.A(ori_ori_n204_), .B(ori_ori_n29_), .Y(ori_ori_n205_));
  INV        o177(.A(ori_ori_n203_), .Y(ori_ori_n206_));
  INV        o178(.A(ori_ori_n51_), .Y(ori_ori_n207_));
  NO3        o179(.A(ori_ori_n141_), .B(ori_ori_n72_), .C(ori_ori_n71_), .Y(ori_ori_n208_));
  NA2        o180(.A(ori_ori_n208_), .B(ori_ori_n91_), .Y(ori_ori_n209_));
  NA3        o181(.A(ori_ori_n209_), .B(ori_ori_n105_), .C(j), .Y(ori_ori_n210_));
  NO3        o182(.A(ori_ori_n158_), .B(ori_ori_n61_), .C(i), .Y(ori_ori_n211_));
  NA2        o183(.A(ori_ori_n210_), .B(ori_ori_n139_), .Y(ori_ori_n212_));
  NO2        o184(.A(ori_ori_n212_), .B(ori_ori_n206_), .Y(ori_ori_n213_));
  NA2        o185(.A(ori_ori_n213_), .B(ori_ori_n200_), .Y(ori08));
  NO2        o186(.A(k), .B(h), .Y(ori_ori_n215_));
  AO210      o187(.A0(ori_ori_n103_), .A1(ori_ori_n150_), .B0(ori_ori_n215_), .Y(ori_ori_n216_));
  NO2        o188(.A(ori_ori_n216_), .B(ori_ori_n113_), .Y(ori_ori_n217_));
  NA2        o189(.A(ori_ori_n186_), .B(ori_ori_n39_), .Y(ori_ori_n218_));
  NA2        o190(.A(ori_ori_n218_), .B(ori_ori_n158_), .Y(ori_ori_n219_));
  NA2        o191(.A(ori_ori_n219_), .B(ori_ori_n217_), .Y(ori_ori_n220_));
  INV        o192(.A(ori_ori_n220_), .Y(ori_ori_n221_));
  INV        o193(.A(ori_ori_n216_), .Y(ori_ori_n222_));
  NA2        o194(.A(ori_ori_n222_), .B(ori_ori_n140_), .Y(ori_ori_n223_));
  INV        o195(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NA3        o196(.A(ori_ori_n209_), .B(ori_ori_n120_), .C(ori_ori_n127_), .Y(ori_ori_n225_));
  INV        o197(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NO3        o198(.A(ori_ori_n226_), .B(ori_ori_n224_), .C(ori_ori_n221_), .Y(ori_ori_n227_));
  INV        o199(.A(ori_ori_n102_), .Y(ori_ori_n228_));
  NA2        o200(.A(l), .B(ori_ori_n38_), .Y(ori_ori_n229_));
  NO4        o201(.A(ori_ori_n208_), .B(ori_ori_n61_), .C(n), .D(i), .Y(ori_ori_n230_));
  BUFFER     o202(.A(h), .Y(ori_ori_n231_));
  NO2        o203(.A(ori_ori_n230_), .B(ori_ori_n211_), .Y(ori_ori_n232_));
  NO2        o204(.A(ori_ori_n232_), .B(ori_ori_n229_), .Y(ori_ori_n233_));
  AOI210     o205(.A0(ori_ori_n228_), .A1(l), .B0(ori_ori_n233_), .Y(ori_ori_n234_));
  NO2        o206(.A(ori_ori_n113_), .B(ori_ori_n52_), .Y(ori_ori_n235_));
  NO2        o207(.A(ori_ori_n208_), .B(n), .Y(ori_ori_n236_));
  BUFFER     o208(.A(ori_ori_n235_), .Y(ori_ori_n237_));
  AOI220     o209(.A0(ori_ori_n237_), .A1(ori_ori_n202_), .B0(ori_ori_n236_), .B1(ori_ori_n217_), .Y(ori_ori_n238_));
  NA3        o210(.A(ori_ori_n238_), .B(ori_ori_n234_), .C(ori_ori_n227_), .Y(ori09));
  INV        o211(.A(ori_ori_n187_), .Y(ori_ori_n240_));
  NA2        o212(.A(c), .B(ori_ori_n48_), .Y(ori_ori_n241_));
  NO2        o213(.A(ori_ori_n241_), .B(ori_ori_n143_), .Y(ori_ori_n242_));
  NA3        o214(.A(ori_ori_n242_), .B(ori_ori_n166_), .C(f), .Y(ori_ori_n243_));
  OR2        o215(.A(ori_ori_n201_), .B(ori_ori_n177_), .Y(ori_ori_n244_));
  INV        o216(.A(ori_ori_n244_), .Y(ori_ori_n245_));
  NA2        o217(.A(ori_ori_n42_), .B(ori_ori_n245_), .Y(ori_ori_n246_));
  NA2        o218(.A(ori_ori_n246_), .B(ori_ori_n243_), .Y(ori_ori_n247_));
  NO2        o219(.A(ori_ori_n247_), .B(ori_ori_n240_), .Y(ori_ori_n248_));
  NO2        o220(.A(ori_ori_n91_), .B(ori_ori_n85_), .Y(ori_ori_n249_));
  NA2        o221(.A(ori_ori_n249_), .B(ori_ori_n88_), .Y(ori_ori_n250_));
  NA2        o222(.A(e), .B(d), .Y(ori_ori_n251_));
  OAI220     o223(.A0(ori_ori_n251_), .A1(c), .B0(ori_ori_n118_), .B1(d), .Y(ori_ori_n252_));
  NA3        o224(.A(ori_ori_n252_), .B(ori_ori_n153_), .C(ori_ori_n164_), .Y(ori_ori_n253_));
  AOI210     o225(.A0(ori_ori_n171_), .A1(ori_ori_n67_), .B0(ori_ori_n91_), .Y(ori_ori_n254_));
  INV        o226(.A(ori_ori_n254_), .Y(ori_ori_n255_));
  NA2        o227(.A(ori_ori_n255_), .B(ori_ori_n253_), .Y(ori_ori_n256_));
  NO2        o228(.A(ori_ori_n256_), .B(ori_ori_n387_), .Y(ori_ori_n257_));
  NA2        o229(.A(ori_ori_n180_), .B(ori_ori_n186_), .Y(ori_ori_n258_));
  AO220      o230(.A0(ori_ori_n153_), .A1(ori_ori_n231_), .B0(ori_ori_n63_), .B1(f), .Y(ori_ori_n259_));
  NA2        o231(.A(ori_ori_n259_), .B(ori_ori_n252_), .Y(ori_ori_n260_));
  BUFFER     o232(.A(ori_ori_n260_), .Y(ori_ori_n261_));
  NA3        o233(.A(ori_ori_n261_), .B(ori_ori_n257_), .C(ori_ori_n248_), .Y(ori12));
  NO4        o234(.A(ori_ori_n145_), .B(ori_ori_n103_), .C(ori_ori_n179_), .D(ori_ori_n83_), .Y(ori_ori_n263_));
  AOI210     o235(.A0(ori_ori_n93_), .A1(ori_ori_n121_), .B0(ori_ori_n79_), .Y(ori_ori_n264_));
  OR2        o236(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n265_));
  NO2        o237(.A(ori_ori_n133_), .B(ori_ori_n83_), .Y(ori_ori_n266_));
  OAI210     o238(.A0(ori_ori_n266_), .A1(ori_ori_n265_), .B0(ori_ori_n141_), .Y(ori_ori_n267_));
  NO2        o239(.A(ori_ori_n102_), .B(ori_ori_n30_), .Y(ori_ori_n268_));
  INV        o240(.A(ori_ori_n268_), .Y(ori_ori_n269_));
  NA2        o241(.A(ori_ori_n49_), .B(g), .Y(ori_ori_n270_));
  AOI210     o242(.A0(ori_ori_n205_), .A1(ori_ori_n270_), .B0(m), .Y(ori_ori_n271_));
  NA2        o243(.A(ori_ori_n271_), .B(ori_ori_n119_), .Y(ori_ori_n272_));
  INV        o244(.A(ori_ori_n272_), .Y(ori_ori_n273_));
  NO2        o245(.A(ori_ori_n157_), .B(ori_ori_n83_), .Y(ori_ori_n274_));
  NA2        o246(.A(ori_ori_n274_), .B(ori_ori_n126_), .Y(ori_ori_n275_));
  INV        o247(.A(ori_ori_n275_), .Y(ori_ori_n276_));
  NO2        o248(.A(ori_ori_n276_), .B(ori_ori_n273_), .Y(ori_ori_n277_));
  NA2        o249(.A(ori_ori_n91_), .B(ori_ori_n59_), .Y(ori_ori_n278_));
  INV        o250(.A(ori_ori_n63_), .Y(ori_ori_n279_));
  NOi31      o251(.An(ori_ori_n278_), .B(ori_ori_n279_), .C(ori_ori_n83_), .Y(ori_ori_n280_));
  NA2        o252(.A(ori_ori_n162_), .B(g), .Y(ori_ori_n281_));
  INV        o253(.A(ori_ori_n281_), .Y(ori_ori_n282_));
  OAI210     o254(.A0(ori_ori_n264_), .A1(ori_ori_n263_), .B0(ori_ori_n278_), .Y(ori_ori_n283_));
  INV        o255(.A(ori_ori_n283_), .Y(ori_ori_n284_));
  NO3        o256(.A(ori_ori_n284_), .B(ori_ori_n282_), .C(ori_ori_n280_), .Y(ori_ori_n285_));
  NA4        o257(.A(ori_ori_n285_), .B(ori_ori_n277_), .C(ori_ori_n269_), .D(ori_ori_n267_), .Y(ori13));
  NAi21      o258(.An(c), .B(e), .Y(ori_ori_n287_));
  AN2        o259(.A(d), .B(c), .Y(ori_ori_n288_));
  NA2        o260(.A(ori_ori_n288_), .B(ori_ori_n48_), .Y(ori_ori_n289_));
  OR2        o261(.A(f), .B(e), .Y(ori_ori_n290_));
  NO3        o262(.A(m), .B(i), .C(h), .Y(ori_ori_n291_));
  NA3        o263(.A(k), .B(j), .C(i), .Y(ori_ori_n292_));
  NO2        o264(.A(f), .B(c), .Y(ori_ori_n293_));
  NOi21      o265(.An(ori_ori_n293_), .B(ori_ori_n145_), .Y(ori_ori_n294_));
  AN3        o266(.A(g), .B(f), .C(c), .Y(ori_ori_n295_));
  NA3        o267(.A(l), .B(k), .C(j), .Y(ori_ori_n296_));
  NA2        o268(.A(i), .B(h), .Y(ori_ori_n297_));
  NO3        o269(.A(ori_ori_n297_), .B(ori_ori_n296_), .C(ori_ori_n51_), .Y(ori_ori_n298_));
  NO2        o270(.A(ori_ori_n112_), .B(ori_ori_n83_), .Y(ori_ori_n299_));
  NOi21      o271(.An(m), .B(n), .Y(ori_ori_n300_));
  INV        o272(.A(ori_ori_n112_), .Y(ori_ori_n301_));
  NA2        o273(.A(ori_ori_n178_), .B(ori_ori_n301_), .Y(ori_ori_n302_));
  INV        o274(.A(ori_ori_n302_), .Y(ori00));
  NA2        o275(.A(ori_ori_n166_), .B(f), .Y(ori_ori_n304_));
  NO2        o276(.A(ori_ori_n304_), .B(ori_ori_n289_), .Y(ori_ori_n305_));
  INV        o277(.A(ori_ori_n305_), .Y(ori_ori_n306_));
  NO2        o278(.A(h), .B(g), .Y(ori_ori_n307_));
  NA2        o279(.A(ori_ori_n193_), .B(ori_ori_n98_), .Y(ori_ori_n308_));
  NA2        o280(.A(ori_ori_n308_), .B(ori_ori_n306_), .Y(ori01));
  INV        o281(.A(ori_ori_n111_), .Y(ori_ori_n310_));
  NA2        o282(.A(ori_ori_n138_), .B(i), .Y(ori_ori_n311_));
  NA2        o283(.A(ori_ori_n311_), .B(ori_ori_n310_), .Y(ori_ori_n312_));
  INV        o284(.A(ori_ori_n258_), .Y(ori_ori_n313_));
  INV        o285(.A(ori_ori_n250_), .Y(ori_ori_n314_));
  INV        o286(.A(ori_ori_n169_), .Y(ori_ori_n315_));
  OR2        o287(.A(ori_ori_n75_), .B(ori_ori_n73_), .Y(ori_ori_n316_));
  NA2        o288(.A(ori_ori_n316_), .B(ori_ori_n315_), .Y(ori_ori_n317_));
  NO4        o289(.A(ori_ori_n317_), .B(ori_ori_n314_), .C(ori_ori_n313_), .D(ori_ori_n312_), .Y(ori_ori_n318_));
  NA2        o290(.A(ori_ori_n110_), .B(ori_ori_n75_), .Y(ori_ori_n319_));
  NA2        o291(.A(ori_ori_n319_), .B(ori_ori_n202_), .Y(ori_ori_n320_));
  NO2        o292(.A(ori_ori_n81_), .B(ori_ori_n45_), .Y(ori_ori_n321_));
  INV        o293(.A(ori_ori_n130_), .Y(ori_ori_n322_));
  NO2        o294(.A(ori_ori_n322_), .B(ori_ori_n321_), .Y(ori_ori_n323_));
  NO3        o295(.A(ori_ori_n297_), .B(ori_ori_n64_), .C(ori_ori_n40_), .Y(ori_ori_n324_));
  NO2        o296(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n325_));
  NO4        o297(.A(ori_ori_n297_), .B(ori_ori_n325_), .C(ori_ori_n62_), .D(ori_ori_n40_), .Y(ori_ori_n326_));
  INV        o298(.A(ori_ori_n326_), .Y(ori_ori_n327_));
  NA4        o299(.A(ori_ori_n327_), .B(ori_ori_n323_), .C(ori_ori_n320_), .D(ori_ori_n318_), .Y(ori06));
  NO2        o300(.A(ori_ori_n85_), .B(ori_ori_n41_), .Y(ori_ori_n329_));
  OAI210     o301(.A0(ori_ori_n329_), .A1(ori_ori_n324_), .B0(ori_ori_n126_), .Y(ori_ori_n330_));
  INV        o302(.A(ori_ori_n330_), .Y(ori_ori_n331_));
  NO2        o303(.A(ori_ori_n331_), .B(ori_ori_n107_), .Y(ori_ori_n332_));
  NO2        o304(.A(ori_ori_n171_), .B(ori_ori_n59_), .Y(ori_ori_n333_));
  NO2        o305(.A(ori_ori_n158_), .B(ori_ori_n100_), .Y(ori_ori_n334_));
  NO2        o306(.A(ori_ori_n334_), .B(ori_ori_n333_), .Y(ori_ori_n335_));
  OAI220     o307(.A0(ori_ori_n218_), .A1(ori_ori_n100_), .B0(ori_ori_n168_), .B1(ori_ori_n171_), .Y(ori_ori_n336_));
  NAi21      o308(.An(j), .B(i), .Y(ori_ori_n337_));
  NO4        o309(.A(ori_ori_n325_), .B(ori_ori_n337_), .C(ori_ori_n145_), .D(ori_ori_n94_), .Y(ori_ori_n338_));
  NO3        o310(.A(ori_ori_n338_), .B(ori_ori_n162_), .C(ori_ori_n336_), .Y(ori_ori_n339_));
  NA4        o311(.A(ori_ori_n339_), .B(ori_ori_n335_), .C(ori_ori_n332_), .D(ori_ori_n327_), .Y(ori07));
  NOi31      o312(.An(n), .B(m), .C(b), .Y(ori_ori_n341_));
  NO2        o313(.A(ori_ori_n290_), .B(ori_ori_n145_), .Y(ori_ori_n342_));
  NO2        o314(.A(ori_ori_n292_), .B(ori_ori_n114_), .Y(ori_ori_n343_));
  INV        o315(.A(ori_ori_n342_), .Y(ori_ori_n344_));
  NO2        o316(.A(e), .B(c), .Y(ori_ori_n345_));
  NO2        o317(.A(ori_ori_n51_), .B(ori_ori_n83_), .Y(ori_ori_n346_));
  NA2        o318(.A(ori_ori_n346_), .B(ori_ori_n345_), .Y(ori_ori_n347_));
  INV        o319(.A(ori_ori_n347_), .Y(ori_ori_n348_));
  NA2        o320(.A(ori_ori_n215_), .B(ori_ori_n207_), .Y(ori_ori_n349_));
  INV        o321(.A(ori_ori_n349_), .Y(ori_ori_n350_));
  NO3        o322(.A(ori_ori_n145_), .B(d), .C(c), .Y(ori_ori_n351_));
  NO2        o323(.A(ori_ori_n350_), .B(ori_ori_n348_), .Y(ori_ori_n352_));
  NOi31      o324(.An(m), .B(n), .C(b), .Y(ori_ori_n353_));
  NA2        o325(.A(ori_ori_n295_), .B(ori_ori_n160_), .Y(ori_ori_n354_));
  NO2        o326(.A(ori_ori_n354_), .B(ori_ori_n145_), .Y(ori_ori_n355_));
  NO2        o327(.A(ori_ori_n291_), .B(ori_ori_n355_), .Y(ori_ori_n356_));
  NA2        o328(.A(ori_ori_n300_), .B(ori_ori_n143_), .Y(ori_ori_n357_));
  NO2        o329(.A(ori_ori_n390_), .B(ori_ori_n298_), .Y(ori_ori_n358_));
  NA4        o330(.A(ori_ori_n358_), .B(ori_ori_n356_), .C(ori_ori_n352_), .D(ori_ori_n344_), .Y(ori_ori_n359_));
  NO2        o331(.A(ori_ori_n135_), .B(j), .Y(ori_ori_n360_));
  NO2        o332(.A(ori_ori_n360_), .B(ori_ori_n294_), .Y(ori_ori_n361_));
  INV        o333(.A(ori_ori_n31_), .Y(ori_ori_n362_));
  NA2        o334(.A(ori_ori_n362_), .B(ori_ori_n307_), .Y(ori_ori_n363_));
  INV        o335(.A(a), .Y(ori_ori_n364_));
  NO2        o336(.A(ori_ori_n386_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  INV        o337(.A(ori_ori_n365_), .Y(ori_ori_n366_));
  NA3        o338(.A(ori_ori_n366_), .B(ori_ori_n363_), .C(ori_ori_n361_), .Y(ori_ori_n367_));
  NA2        o339(.A(h), .B(ori_ori_n343_), .Y(ori_ori_n368_));
  NA2        o340(.A(ori_ori_n341_), .B(ori_ori_n241_), .Y(ori_ori_n369_));
  NO2        o341(.A(ori_ori_n287_), .B(ori_ori_n51_), .Y(ori_ori_n370_));
  NA2        o342(.A(ori_ori_n370_), .B(f), .Y(ori_ori_n371_));
  NA3        o343(.A(ori_ori_n371_), .B(ori_ori_n369_), .C(ori_ori_n368_), .Y(ori_ori_n372_));
  NO2        o344(.A(ori_ori_n353_), .B(ori_ori_n372_), .Y(ori_ori_n373_));
  INV        o345(.A(ori_ori_n189_), .Y(ori_ori_n374_));
  BUFFER     o346(.A(ori_ori_n51_), .Y(ori_ori_n375_));
  OAI210     o347(.A0(ori_ori_n375_), .A1(f), .B0(ori_ori_n374_), .Y(ori_ori_n376_));
  INV        o348(.A(ori_ori_n376_), .Y(ori_ori_n377_));
  NO2        o349(.A(h), .B(ori_ori_n62_), .Y(ori_ori_n378_));
  NA2        o350(.A(ori_ori_n299_), .B(ori_ori_n84_), .Y(ori_ori_n379_));
  INV        o351(.A(ori_ori_n379_), .Y(ori_ori_n380_));
  NO3        o352(.A(ori_ori_n380_), .B(ori_ori_n378_), .C(ori_ori_n351_), .Y(ori_ori_n381_));
  NA3        o353(.A(ori_ori_n381_), .B(ori_ori_n377_), .C(ori_ori_n373_), .Y(ori_ori_n382_));
  OR3        o354(.A(ori_ori_n382_), .B(ori_ori_n367_), .C(ori_ori_n359_), .Y(ori04));
  INV        o355(.A(ori_ori_n46_), .Y(ori_ori_n386_));
  INV        o356(.A(ori_ori_n250_), .Y(ori_ori_n387_));
  INV        o357(.A(c), .Y(ori_ori_n388_));
  INV        o358(.A(ori_ori_n162_), .Y(ori_ori_n389_));
  INV        o359(.A(ori_ori_n357_), .Y(ori_ori_n390_));
  ZERO       o360(.Y(ori02));
  ZERO       o361(.Y(ori03));
  ZERO       o362(.Y(ori05));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  NO2        m0023(.A(mai_mai_n51_), .B(mai_mai_n50_), .Y(mai_mai_n52_));
  NO3        m0024(.A(mai_mai_n48_), .B(mai_mai_n43_), .C(mai_mai_n39_), .Y(mai_mai_n53_));
  NO2        m0025(.A(mai_mai_n53_), .B(mai_mai_n32_), .Y(mai_mai_n54_));
  INV        m0026(.A(c), .Y(mai_mai_n55_));
  NA2        m0027(.A(e), .B(b), .Y(mai_mai_n56_));
  NO2        m0028(.A(mai_mai_n56_), .B(mai_mai_n55_), .Y(mai_mai_n57_));
  INV        m0029(.A(d), .Y(mai_mai_n58_));
  NA2        m0030(.A(g), .B(mai_mai_n58_), .Y(mai_mai_n59_));
  NAi21      m0031(.An(i), .B(h), .Y(mai_mai_n60_));
  NAi31      m0032(.An(i), .B(l), .C(j), .Y(mai_mai_n61_));
  OAI220     m0033(.A0(mai_mai_n61_), .A1(mai_mai_n49_), .B0(mai_mai_n60_), .B1(mai_mai_n44_), .Y(mai_mai_n62_));
  NAi31      m0034(.An(mai_mai_n59_), .B(mai_mai_n62_), .C(mai_mai_n57_), .Y(mai_mai_n63_));
  NA2        m0035(.A(g), .B(f), .Y(mai_mai_n64_));
  NAi21      m0036(.An(i), .B(j), .Y(mai_mai_n65_));
  NAi32      m0037(.An(n), .Bn(k), .C(m), .Y(mai_mai_n66_));
  NAi31      m0038(.An(l), .B(m), .C(k), .Y(mai_mai_n67_));
  NAi21      m0039(.An(e), .B(h), .Y(mai_mai_n68_));
  NAi41      m0040(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n69_));
  INV        m0041(.A(m), .Y(mai_mai_n70_));
  NOi21      m0042(.An(k), .B(l), .Y(mai_mai_n71_));
  NA2        m0043(.A(mai_mai_n71_), .B(mai_mai_n70_), .Y(mai_mai_n72_));
  AN4        m0044(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n73_));
  NOi31      m0045(.An(h), .B(g), .C(f), .Y(mai_mai_n74_));
  NA2        m0046(.A(mai_mai_n74_), .B(mai_mai_n73_), .Y(mai_mai_n75_));
  NAi32      m0047(.An(m), .Bn(k), .C(j), .Y(mai_mai_n76_));
  NOi32      m0048(.An(h), .Bn(g), .C(f), .Y(mai_mai_n77_));
  NA2        m0049(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OA220      m0050(.A0(mai_mai_n78_), .A1(mai_mai_n76_), .B0(mai_mai_n75_), .B1(mai_mai_n72_), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n63_), .Y(mai_mai_n80_));
  INV        m0052(.A(n), .Y(mai_mai_n81_));
  NOi32      m0053(.An(e), .Bn(b), .C(d), .Y(mai_mai_n82_));
  NA2        m0054(.A(mai_mai_n82_), .B(mai_mai_n81_), .Y(mai_mai_n83_));
  INV        m0055(.A(j), .Y(mai_mai_n84_));
  AN3        m0056(.A(m), .B(k), .C(i), .Y(mai_mai_n85_));
  NA3        m0057(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .Y(mai_mai_n86_));
  NO2        m0058(.A(mai_mai_n86_), .B(f), .Y(mai_mai_n87_));
  NAi32      m0059(.An(g), .Bn(f), .C(h), .Y(mai_mai_n88_));
  NAi31      m0060(.An(j), .B(m), .C(l), .Y(mai_mai_n89_));
  NO2        m0061(.A(mai_mai_n89_), .B(mai_mai_n88_), .Y(mai_mai_n90_));
  NA2        m0062(.A(m), .B(l), .Y(mai_mai_n91_));
  NAi31      m0063(.An(k), .B(j), .C(g), .Y(mai_mai_n92_));
  NO3        m0064(.A(mai_mai_n92_), .B(mai_mai_n91_), .C(f), .Y(mai_mai_n93_));
  AN2        m0065(.A(j), .B(g), .Y(mai_mai_n94_));
  NOi32      m0066(.An(m), .Bn(l), .C(i), .Y(mai_mai_n95_));
  NOi21      m0067(.An(g), .B(i), .Y(mai_mai_n96_));
  NOi32      m0068(.An(m), .Bn(j), .C(k), .Y(mai_mai_n97_));
  AOI220     m0069(.A0(mai_mai_n97_), .A1(mai_mai_n96_), .B0(mai_mai_n95_), .B1(mai_mai_n94_), .Y(mai_mai_n98_));
  NO2        m0070(.A(mai_mai_n98_), .B(f), .Y(mai_mai_n99_));
  NO3        m0071(.A(mai_mai_n99_), .B(mai_mai_n93_), .C(mai_mai_n90_), .Y(mai_mai_n100_));
  NAi41      m0072(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n101_));
  AN2        m0073(.A(e), .B(b), .Y(mai_mai_n102_));
  NOi31      m0074(.An(c), .B(h), .C(f), .Y(mai_mai_n103_));
  NA2        m0075(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NO3        m0076(.A(mai_mai_n104_), .B(mai_mai_n101_), .C(g), .Y(mai_mai_n105_));
  NOi21      m0077(.An(i), .B(h), .Y(mai_mai_n106_));
  NA3        m0078(.A(mai_mai_n106_), .B(g), .C(mai_mai_n36_), .Y(mai_mai_n107_));
  INV        m0079(.A(a), .Y(mai_mai_n108_));
  NA2        m0080(.A(mai_mai_n102_), .B(mai_mai_n108_), .Y(mai_mai_n109_));
  INV        m0081(.A(l), .Y(mai_mai_n110_));
  NOi21      m0082(.An(m), .B(n), .Y(mai_mai_n111_));
  AN2        m0083(.A(k), .B(h), .Y(mai_mai_n112_));
  NO2        m0084(.A(mai_mai_n107_), .B(mai_mai_n83_), .Y(mai_mai_n113_));
  INV        m0085(.A(b), .Y(mai_mai_n114_));
  NA2        m0086(.A(l), .B(j), .Y(mai_mai_n115_));
  AN2        m0087(.A(k), .B(i), .Y(mai_mai_n116_));
  NA2        m0088(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NA2        m0089(.A(g), .B(e), .Y(mai_mai_n118_));
  NOi32      m0090(.An(c), .Bn(a), .C(d), .Y(mai_mai_n119_));
  NA2        m0091(.A(mai_mai_n119_), .B(mai_mai_n111_), .Y(mai_mai_n120_));
  NO4        m0092(.A(mai_mai_n120_), .B(mai_mai_n118_), .C(mai_mai_n117_), .D(mai_mai_n114_), .Y(mai_mai_n121_));
  NO3        m0093(.A(mai_mai_n121_), .B(mai_mai_n113_), .C(mai_mai_n105_), .Y(mai_mai_n122_));
  OAI210     m0094(.A0(mai_mai_n100_), .A1(mai_mai_n83_), .B0(mai_mai_n122_), .Y(mai_mai_n123_));
  NOi31      m0095(.An(k), .B(m), .C(j), .Y(mai_mai_n124_));
  NA3        m0096(.A(mai_mai_n124_), .B(mai_mai_n74_), .C(mai_mai_n73_), .Y(mai_mai_n125_));
  NOi31      m0097(.An(k), .B(m), .C(i), .Y(mai_mai_n126_));
  INV        m0098(.A(mai_mai_n125_), .Y(mai_mai_n127_));
  NOi32      m0099(.An(f), .Bn(b), .C(e), .Y(mai_mai_n128_));
  NAi21      m0100(.An(g), .B(h), .Y(mai_mai_n129_));
  NAi21      m0101(.An(m), .B(n), .Y(mai_mai_n130_));
  NAi21      m0102(.An(j), .B(k), .Y(mai_mai_n131_));
  NO3        m0103(.A(mai_mai_n131_), .B(mai_mai_n130_), .C(mai_mai_n129_), .Y(mai_mai_n132_));
  NAi41      m0104(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n133_));
  NAi31      m0105(.An(j), .B(k), .C(h), .Y(mai_mai_n134_));
  NO3        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n130_), .Y(mai_mai_n135_));
  AOI210     m0107(.A0(mai_mai_n132_), .A1(mai_mai_n128_), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  NO2        m0108(.A(k), .B(j), .Y(mai_mai_n137_));
  NO2        m0109(.A(mai_mai_n137_), .B(mai_mai_n130_), .Y(mai_mai_n138_));
  AN2        m0110(.A(k), .B(j), .Y(mai_mai_n139_));
  NAi21      m0111(.An(c), .B(b), .Y(mai_mai_n140_));
  NA2        m0112(.A(f), .B(d), .Y(mai_mai_n141_));
  NO4        m0113(.A(mai_mai_n141_), .B(mai_mai_n140_), .C(mai_mai_n139_), .D(mai_mai_n129_), .Y(mai_mai_n142_));
  NAi31      m0114(.An(f), .B(e), .C(b), .Y(mai_mai_n143_));
  NA2        m0115(.A(mai_mai_n142_), .B(mai_mai_n138_), .Y(mai_mai_n144_));
  NA2        m0116(.A(d), .B(b), .Y(mai_mai_n145_));
  NAi21      m0117(.An(e), .B(f), .Y(mai_mai_n146_));
  NO2        m0118(.A(mai_mai_n146_), .B(mai_mai_n145_), .Y(mai_mai_n147_));
  NA2        m0119(.A(b), .B(a), .Y(mai_mai_n148_));
  NAi21      m0120(.An(e), .B(g), .Y(mai_mai_n149_));
  NAi21      m0121(.An(c), .B(d), .Y(mai_mai_n150_));
  NAi31      m0122(.An(l), .B(k), .C(h), .Y(mai_mai_n151_));
  NO2        m0123(.A(mai_mai_n130_), .B(mai_mai_n151_), .Y(mai_mai_n152_));
  NA2        m0124(.A(mai_mai_n152_), .B(mai_mai_n147_), .Y(mai_mai_n153_));
  NAi41      m0125(.An(mai_mai_n127_), .B(mai_mai_n153_), .C(mai_mai_n144_), .D(mai_mai_n136_), .Y(mai_mai_n154_));
  NAi31      m0126(.An(e), .B(f), .C(b), .Y(mai_mai_n155_));
  NOi21      m0127(.An(g), .B(d), .Y(mai_mai_n156_));
  NO2        m0128(.A(mai_mai_n156_), .B(mai_mai_n155_), .Y(mai_mai_n157_));
  NOi21      m0129(.An(h), .B(i), .Y(mai_mai_n158_));
  NOi21      m0130(.An(k), .B(m), .Y(mai_mai_n159_));
  NA3        m0131(.A(mai_mai_n159_), .B(mai_mai_n158_), .C(n), .Y(mai_mai_n160_));
  NOi21      m0132(.An(mai_mai_n157_), .B(mai_mai_n160_), .Y(mai_mai_n161_));
  NOi21      m0133(.An(h), .B(g), .Y(mai_mai_n162_));
  NO2        m0134(.A(mai_mai_n141_), .B(mai_mai_n140_), .Y(mai_mai_n163_));
  NA2        m0135(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NOi32      m0136(.An(n), .Bn(k), .C(m), .Y(mai_mai_n165_));
  NA2        m0137(.A(l), .B(i), .Y(mai_mai_n166_));
  NA2        m0138(.A(mai_mai_n166_), .B(mai_mai_n165_), .Y(mai_mai_n167_));
  NO2        m0139(.A(mai_mai_n167_), .B(mai_mai_n164_), .Y(mai_mai_n168_));
  NAi31      m0140(.An(d), .B(f), .C(c), .Y(mai_mai_n169_));
  NAi31      m0141(.An(e), .B(f), .C(c), .Y(mai_mai_n170_));
  NA2        m0142(.A(mai_mai_n170_), .B(mai_mai_n169_), .Y(mai_mai_n171_));
  NA2        m0143(.A(j), .B(h), .Y(mai_mai_n172_));
  OR3        m0144(.A(n), .B(m), .C(k), .Y(mai_mai_n173_));
  NO2        m0145(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  NAi32      m0146(.An(m), .Bn(k), .C(n), .Y(mai_mai_n175_));
  NO2        m0147(.A(mai_mai_n175_), .B(mai_mai_n172_), .Y(mai_mai_n176_));
  AOI220     m0148(.A0(mai_mai_n176_), .A1(mai_mai_n157_), .B0(mai_mai_n174_), .B1(mai_mai_n171_), .Y(mai_mai_n177_));
  NO2        m0149(.A(n), .B(m), .Y(mai_mai_n178_));
  NA2        m0150(.A(mai_mai_n178_), .B(mai_mai_n50_), .Y(mai_mai_n179_));
  NAi21      m0151(.An(f), .B(e), .Y(mai_mai_n180_));
  NA2        m0152(.A(d), .B(c), .Y(mai_mai_n181_));
  NO2        m0153(.A(mai_mai_n181_), .B(mai_mai_n180_), .Y(mai_mai_n182_));
  NOi21      m0154(.An(mai_mai_n182_), .B(mai_mai_n179_), .Y(mai_mai_n183_));
  NAi31      m0155(.An(m), .B(n), .C(b), .Y(mai_mai_n184_));
  NA2        m0156(.A(k), .B(i), .Y(mai_mai_n185_));
  NAi21      m0157(.An(h), .B(f), .Y(mai_mai_n186_));
  NO2        m0158(.A(mai_mai_n186_), .B(mai_mai_n185_), .Y(mai_mai_n187_));
  NO2        m0159(.A(mai_mai_n184_), .B(mai_mai_n150_), .Y(mai_mai_n188_));
  NA2        m0160(.A(mai_mai_n188_), .B(mai_mai_n187_), .Y(mai_mai_n189_));
  NOi32      m0161(.An(f), .Bn(c), .C(d), .Y(mai_mai_n190_));
  NOi32      m0162(.An(f), .Bn(c), .C(e), .Y(mai_mai_n191_));
  NO2        m0163(.A(mai_mai_n191_), .B(mai_mai_n190_), .Y(mai_mai_n192_));
  NO3        m0164(.A(n), .B(m), .C(j), .Y(mai_mai_n193_));
  NA2        m0165(.A(mai_mai_n193_), .B(mai_mai_n112_), .Y(mai_mai_n194_));
  AO210      m0166(.A0(mai_mai_n194_), .A1(mai_mai_n179_), .B0(mai_mai_n192_), .Y(mai_mai_n195_));
  NAi41      m0167(.An(mai_mai_n183_), .B(mai_mai_n195_), .C(mai_mai_n189_), .D(mai_mai_n177_), .Y(mai_mai_n196_));
  OR4        m0168(.A(mai_mai_n196_), .B(mai_mai_n168_), .C(mai_mai_n161_), .D(mai_mai_n154_), .Y(mai_mai_n197_));
  NO4        m0169(.A(mai_mai_n197_), .B(mai_mai_n123_), .C(mai_mai_n80_), .D(mai_mai_n54_), .Y(mai_mai_n198_));
  NA3        m0170(.A(m), .B(mai_mai_n110_), .C(j), .Y(mai_mai_n199_));
  NAi31      m0171(.An(n), .B(h), .C(g), .Y(mai_mai_n200_));
  NO2        m0172(.A(mai_mai_n200_), .B(mai_mai_n199_), .Y(mai_mai_n201_));
  NOi32      m0173(.An(m), .Bn(k), .C(l), .Y(mai_mai_n202_));
  NA3        m0174(.A(mai_mai_n202_), .B(mai_mai_n84_), .C(g), .Y(mai_mai_n203_));
  NO2        m0175(.A(mai_mai_n203_), .B(n), .Y(mai_mai_n204_));
  NOi21      m0176(.An(k), .B(j), .Y(mai_mai_n205_));
  NA4        m0177(.A(mai_mai_n205_), .B(mai_mai_n111_), .C(i), .D(g), .Y(mai_mai_n206_));
  AN2        m0178(.A(i), .B(g), .Y(mai_mai_n207_));
  NA3        m0179(.A(mai_mai_n71_), .B(mai_mai_n207_), .C(mai_mai_n111_), .Y(mai_mai_n208_));
  NA2        m0180(.A(mai_mai_n208_), .B(mai_mai_n206_), .Y(mai_mai_n209_));
  NO3        m0181(.A(mai_mai_n209_), .B(mai_mai_n204_), .C(mai_mai_n201_), .Y(mai_mai_n210_));
  NAi41      m0182(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n211_));
  INV        m0183(.A(mai_mai_n211_), .Y(mai_mai_n212_));
  INV        m0184(.A(f), .Y(mai_mai_n213_));
  INV        m0185(.A(g), .Y(mai_mai_n214_));
  NOi31      m0186(.An(i), .B(j), .C(h), .Y(mai_mai_n215_));
  NOi21      m0187(.An(l), .B(m), .Y(mai_mai_n216_));
  NA2        m0188(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  NO3        m0189(.A(mai_mai_n217_), .B(mai_mai_n214_), .C(mai_mai_n213_), .Y(mai_mai_n218_));
  NA2        m0190(.A(mai_mai_n218_), .B(mai_mai_n212_), .Y(mai_mai_n219_));
  OAI210     m0191(.A0(mai_mai_n210_), .A1(mai_mai_n32_), .B0(mai_mai_n219_), .Y(mai_mai_n220_));
  NOi21      m0192(.An(n), .B(m), .Y(mai_mai_n221_));
  NOi32      m0193(.An(l), .Bn(i), .C(j), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n221_), .Y(mai_mai_n223_));
  OA220      m0195(.A0(mai_mai_n223_), .A1(mai_mai_n104_), .B0(mai_mai_n76_), .B1(mai_mai_n75_), .Y(mai_mai_n224_));
  NAi21      m0196(.An(j), .B(h), .Y(mai_mai_n225_));
  XN2        m0197(.A(i), .B(h), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n227_));
  NOi31      m0199(.An(k), .B(n), .C(m), .Y(mai_mai_n228_));
  NOi31      m0200(.An(mai_mai_n228_), .B(mai_mai_n181_), .C(mai_mai_n180_), .Y(mai_mai_n229_));
  NA2        m0201(.A(mai_mai_n229_), .B(mai_mai_n227_), .Y(mai_mai_n230_));
  NAi31      m0202(.An(f), .B(e), .C(c), .Y(mai_mai_n231_));
  NA4        m0203(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n232_));
  NAi32      m0204(.An(m), .Bn(i), .C(k), .Y(mai_mai_n233_));
  NO3        m0205(.A(mai_mai_n233_), .B(mai_mai_n88_), .C(mai_mai_n232_), .Y(mai_mai_n234_));
  INV        m0206(.A(k), .Y(mai_mai_n235_));
  INV        m0207(.A(mai_mai_n234_), .Y(mai_mai_n236_));
  NAi21      m0208(.An(n), .B(a), .Y(mai_mai_n237_));
  NO2        m0209(.A(mai_mai_n237_), .B(mai_mai_n145_), .Y(mai_mai_n238_));
  NAi41      m0210(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n239_));
  NO2        m0211(.A(mai_mai_n239_), .B(e), .Y(mai_mai_n240_));
  NA2        m0212(.A(mai_mai_n240_), .B(mai_mai_n238_), .Y(mai_mai_n241_));
  AN4        m0213(.A(mai_mai_n241_), .B(mai_mai_n236_), .C(mai_mai_n230_), .D(mai_mai_n224_), .Y(mai_mai_n242_));
  OR2        m0214(.A(h), .B(g), .Y(mai_mai_n243_));
  NO2        m0215(.A(mai_mai_n243_), .B(mai_mai_n101_), .Y(mai_mai_n244_));
  NAi41      m0216(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n245_));
  NO2        m0217(.A(mai_mai_n245_), .B(mai_mai_n213_), .Y(mai_mai_n246_));
  NA2        m0218(.A(mai_mai_n159_), .B(mai_mai_n106_), .Y(mai_mai_n247_));
  NAi21      m0219(.An(mai_mai_n247_), .B(mai_mai_n246_), .Y(mai_mai_n248_));
  NO2        m0220(.A(n), .B(a), .Y(mai_mai_n249_));
  NAi21      m0221(.An(h), .B(i), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n178_), .B(k), .Y(mai_mai_n251_));
  NO2        m0223(.A(mai_mai_n251_), .B(mai_mai_n250_), .Y(mai_mai_n252_));
  NA2        m0224(.A(mai_mai_n252_), .B(mai_mai_n190_), .Y(mai_mai_n253_));
  NA2        m0225(.A(mai_mai_n253_), .B(mai_mai_n248_), .Y(mai_mai_n254_));
  NO2        m0226(.A(mai_mai_n69_), .B(mai_mai_n70_), .Y(mai_mai_n255_));
  NOi32      m0227(.An(l), .Bn(j), .C(i), .Y(mai_mai_n256_));
  NAi21      m0228(.An(f), .B(g), .Y(mai_mai_n257_));
  NO2        m0229(.A(mai_mai_n66_), .B(mai_mai_n115_), .Y(mai_mai_n258_));
  NOi31      m0230(.An(mai_mai_n242_), .B(mai_mai_n254_), .C(mai_mai_n220_), .Y(mai_mai_n259_));
  NO4        m0231(.A(mai_mai_n201_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n260_), .B(mai_mai_n109_), .Y(mai_mai_n261_));
  NA3        m0233(.A(mai_mai_n58_), .B(c), .C(b), .Y(mai_mai_n262_));
  NAi21      m0234(.An(h), .B(g), .Y(mai_mai_n263_));
  OR3        m0235(.A(mai_mai_n263_), .B(mai_mai_n262_), .C(mai_mai_n223_), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n247_), .B(mai_mai_n257_), .Y(mai_mai_n265_));
  NA2        m0237(.A(mai_mai_n265_), .B(mai_mai_n73_), .Y(mai_mai_n266_));
  NAi31      m0238(.An(g), .B(k), .C(h), .Y(mai_mai_n267_));
  NAi31      m0239(.An(e), .B(d), .C(a), .Y(mai_mai_n268_));
  NA2        m0240(.A(mai_mai_n266_), .B(mai_mai_n264_), .Y(mai_mai_n269_));
  NA3        m0241(.A(mai_mai_n159_), .B(mai_mai_n77_), .C(mai_mai_n73_), .Y(mai_mai_n270_));
  BUFFER     m0242(.A(mai_mai_n270_), .Y(mai_mai_n271_));
  NA3        m0243(.A(e), .B(c), .C(b), .Y(mai_mai_n272_));
  NO2        m0244(.A(mai_mai_n59_), .B(mai_mai_n272_), .Y(mai_mai_n273_));
  NAi32      m0245(.An(k), .Bn(i), .C(j), .Y(mai_mai_n274_));
  NA3        m0246(.A(h), .B(mai_mai_n274_), .C(l), .Y(mai_mai_n275_));
  NOi21      m0247(.An(mai_mai_n275_), .B(mai_mai_n49_), .Y(mai_mai_n276_));
  NA2        m0248(.A(mai_mai_n273_), .B(mai_mai_n276_), .Y(mai_mai_n277_));
  NAi21      m0249(.An(l), .B(k), .Y(mai_mai_n278_));
  NO2        m0250(.A(mai_mai_n278_), .B(mai_mai_n49_), .Y(mai_mai_n279_));
  NOi21      m0251(.An(l), .B(j), .Y(mai_mai_n280_));
  NA2        m0252(.A(mai_mai_n162_), .B(mai_mai_n280_), .Y(mai_mai_n281_));
  OR3        m0253(.A(mai_mai_n69_), .B(mai_mai_n70_), .C(e), .Y(mai_mai_n282_));
  AOI210     m0254(.A0(mai_mai_n1430_), .A1(mai_mai_n281_), .B0(mai_mai_n282_), .Y(mai_mai_n283_));
  INV        m0255(.A(mai_mai_n283_), .Y(mai_mai_n284_));
  NAi32      m0256(.An(j), .Bn(h), .C(i), .Y(mai_mai_n285_));
  NAi21      m0257(.An(m), .B(l), .Y(mai_mai_n286_));
  NO3        m0258(.A(mai_mai_n286_), .B(mai_mai_n285_), .C(mai_mai_n81_), .Y(mai_mai_n287_));
  NA2        m0259(.A(h), .B(g), .Y(mai_mai_n288_));
  NA2        m0260(.A(mai_mai_n165_), .B(mai_mai_n45_), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n289_), .B(mai_mai_n288_), .Y(mai_mai_n290_));
  OAI210     m0262(.A0(mai_mai_n290_), .A1(mai_mai_n287_), .B0(mai_mai_n163_), .Y(mai_mai_n291_));
  NA4        m0263(.A(mai_mai_n291_), .B(mai_mai_n284_), .C(mai_mai_n277_), .D(mai_mai_n271_), .Y(mai_mai_n292_));
  NO2        m0264(.A(mai_mai_n143_), .B(d), .Y(mai_mai_n293_));
  NO2        m0265(.A(mai_mai_n104_), .B(mai_mai_n101_), .Y(mai_mai_n294_));
  NAi32      m0266(.An(n), .Bn(m), .C(l), .Y(mai_mai_n295_));
  NO2        m0267(.A(mai_mai_n295_), .B(mai_mai_n285_), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n296_), .B(mai_mai_n182_), .Y(mai_mai_n297_));
  NO2        m0269(.A(mai_mai_n120_), .B(mai_mai_n114_), .Y(mai_mai_n298_));
  NAi31      m0270(.An(k), .B(l), .C(j), .Y(mai_mai_n299_));
  OAI210     m0271(.A0(mai_mai_n278_), .A1(j), .B0(mai_mai_n299_), .Y(mai_mai_n300_));
  NOi21      m0272(.An(mai_mai_n300_), .B(mai_mai_n118_), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n301_), .B(mai_mai_n298_), .Y(mai_mai_n302_));
  NA2        m0274(.A(mai_mai_n302_), .B(mai_mai_n297_), .Y(mai_mai_n303_));
  NO4        m0275(.A(mai_mai_n303_), .B(mai_mai_n292_), .C(mai_mai_n269_), .D(mai_mai_n261_), .Y(mai_mai_n304_));
  NAi21      m0276(.An(m), .B(k), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n226_), .B(mai_mai_n305_), .Y(mai_mai_n306_));
  NAi41      m0278(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n307_), .B(mai_mai_n149_), .Y(mai_mai_n308_));
  NA2        m0280(.A(mai_mai_n308_), .B(mai_mai_n306_), .Y(mai_mai_n309_));
  NA2        m0281(.A(e), .B(c), .Y(mai_mai_n310_));
  NO3        m0282(.A(mai_mai_n310_), .B(n), .C(d), .Y(mai_mai_n311_));
  NOi21      m0283(.An(f), .B(h), .Y(mai_mai_n312_));
  NA2        m0284(.A(mai_mai_n312_), .B(mai_mai_n116_), .Y(mai_mai_n313_));
  NO2        m0285(.A(mai_mai_n313_), .B(mai_mai_n214_), .Y(mai_mai_n314_));
  NAi31      m0286(.An(d), .B(e), .C(b), .Y(mai_mai_n315_));
  NO2        m0287(.A(mai_mai_n130_), .B(mai_mai_n315_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n316_), .B(mai_mai_n314_), .Y(mai_mai_n317_));
  NA2        m0289(.A(mai_mai_n317_), .B(mai_mai_n309_), .Y(mai_mai_n318_));
  NO4        m0290(.A(mai_mai_n307_), .B(mai_mai_n76_), .C(mai_mai_n68_), .D(mai_mai_n214_), .Y(mai_mai_n319_));
  NA2        m0291(.A(mai_mai_n249_), .B(mai_mai_n102_), .Y(mai_mai_n320_));
  OR2        m0292(.A(mai_mai_n320_), .B(mai_mai_n203_), .Y(mai_mai_n321_));
  NOi31      m0293(.An(l), .B(n), .C(m), .Y(mai_mai_n322_));
  NA2        m0294(.A(mai_mai_n322_), .B(mai_mai_n215_), .Y(mai_mai_n323_));
  NO2        m0295(.A(mai_mai_n323_), .B(mai_mai_n192_), .Y(mai_mai_n324_));
  NAi32      m0296(.An(mai_mai_n324_), .Bn(mai_mai_n319_), .C(mai_mai_n321_), .Y(mai_mai_n325_));
  NAi32      m0297(.An(m), .Bn(j), .C(k), .Y(mai_mai_n326_));
  NAi41      m0298(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n327_));
  OAI210     m0299(.A0(mai_mai_n211_), .A1(mai_mai_n326_), .B0(mai_mai_n327_), .Y(mai_mai_n328_));
  NOi31      m0300(.An(j), .B(m), .C(k), .Y(mai_mai_n329_));
  NO2        m0301(.A(mai_mai_n124_), .B(mai_mai_n329_), .Y(mai_mai_n330_));
  AN3        m0302(.A(h), .B(g), .C(f), .Y(mai_mai_n331_));
  NAi31      m0303(.An(mai_mai_n330_), .B(mai_mai_n331_), .C(mai_mai_n328_), .Y(mai_mai_n332_));
  NOi32      m0304(.An(m), .Bn(j), .C(l), .Y(mai_mai_n333_));
  NO2        m0305(.A(mai_mai_n333_), .B(mai_mai_n95_), .Y(mai_mai_n334_));
  NAi32      m0306(.An(mai_mai_n334_), .Bn(mai_mai_n200_), .C(mai_mai_n293_), .Y(mai_mai_n335_));
  NO2        m0307(.A(mai_mai_n286_), .B(mai_mai_n285_), .Y(mai_mai_n336_));
  NO2        m0308(.A(mai_mai_n217_), .B(g), .Y(mai_mai_n337_));
  NO2        m0309(.A(mai_mai_n155_), .B(mai_mai_n81_), .Y(mai_mai_n338_));
  AOI220     m0310(.A0(mai_mai_n338_), .A1(mai_mai_n337_), .B0(mai_mai_n246_), .B1(mai_mai_n336_), .Y(mai_mai_n339_));
  NA2        m0311(.A(mai_mai_n233_), .B(mai_mai_n76_), .Y(mai_mai_n340_));
  NA3        m0312(.A(mai_mai_n340_), .B(mai_mai_n331_), .C(mai_mai_n212_), .Y(mai_mai_n341_));
  NA4        m0313(.A(mai_mai_n341_), .B(mai_mai_n339_), .C(mai_mai_n335_), .D(mai_mai_n332_), .Y(mai_mai_n342_));
  NA3        m0314(.A(h), .B(g), .C(f), .Y(mai_mai_n343_));
  NO2        m0315(.A(mai_mai_n343_), .B(mai_mai_n72_), .Y(mai_mai_n344_));
  NA2        m0316(.A(mai_mai_n327_), .B(mai_mai_n211_), .Y(mai_mai_n345_));
  NA2        m0317(.A(mai_mai_n162_), .B(e), .Y(mai_mai_n346_));
  NO2        m0318(.A(mai_mai_n346_), .B(mai_mai_n41_), .Y(mai_mai_n347_));
  AOI220     m0319(.A0(mai_mai_n347_), .A1(mai_mai_n298_), .B0(mai_mai_n345_), .B1(mai_mai_n344_), .Y(mai_mai_n348_));
  NOi32      m0320(.An(j), .Bn(g), .C(i), .Y(mai_mai_n349_));
  NA3        m0321(.A(mai_mai_n349_), .B(mai_mai_n278_), .C(mai_mai_n111_), .Y(mai_mai_n350_));
  AO210      m0322(.A0(mai_mai_n109_), .A1(mai_mai_n32_), .B0(mai_mai_n350_), .Y(mai_mai_n351_));
  NOi32      m0323(.An(e), .Bn(b), .C(a), .Y(mai_mai_n352_));
  INV        m0324(.A(mai_mai_n305_), .Y(mai_mai_n353_));
  NO3        m0325(.A(mai_mai_n307_), .B(mai_mai_n68_), .C(mai_mai_n214_), .Y(mai_mai_n354_));
  NA3        m0326(.A(mai_mai_n208_), .B(mai_mai_n206_), .C(mai_mai_n35_), .Y(mai_mai_n355_));
  AOI220     m0327(.A0(mai_mai_n355_), .A1(mai_mai_n352_), .B0(mai_mai_n354_), .B1(mai_mai_n353_), .Y(mai_mai_n356_));
  NO2        m0328(.A(mai_mai_n315_), .B(n), .Y(mai_mai_n357_));
  NA2        m0329(.A(mai_mai_n207_), .B(k), .Y(mai_mai_n358_));
  NA3        m0330(.A(m), .B(mai_mai_n110_), .C(mai_mai_n213_), .Y(mai_mai_n359_));
  NA4        m0331(.A(mai_mai_n202_), .B(mai_mai_n84_), .C(g), .D(mai_mai_n213_), .Y(mai_mai_n360_));
  OAI210     m0332(.A0(mai_mai_n359_), .A1(mai_mai_n358_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  NAi41      m0333(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n362_));
  NA2        m0334(.A(mai_mai_n51_), .B(mai_mai_n111_), .Y(mai_mai_n363_));
  NA2        m0335(.A(mai_mai_n361_), .B(mai_mai_n357_), .Y(mai_mai_n364_));
  NA4        m0336(.A(mai_mai_n364_), .B(mai_mai_n356_), .C(mai_mai_n351_), .D(mai_mai_n348_), .Y(mai_mai_n365_));
  NO4        m0337(.A(mai_mai_n365_), .B(mai_mai_n342_), .C(mai_mai_n325_), .D(mai_mai_n318_), .Y(mai_mai_n366_));
  NA4        m0338(.A(mai_mai_n366_), .B(mai_mai_n304_), .C(mai_mai_n259_), .D(mai_mai_n198_), .Y(mai10));
  NA3        m0339(.A(m), .B(k), .C(i), .Y(mai_mai_n368_));
  NO3        m0340(.A(mai_mai_n368_), .B(j), .C(mai_mai_n214_), .Y(mai_mai_n369_));
  NOi21      m0341(.An(e), .B(f), .Y(mai_mai_n370_));
  NO4        m0342(.A(mai_mai_n150_), .B(mai_mai_n370_), .C(n), .D(mai_mai_n108_), .Y(mai_mai_n371_));
  NAi31      m0343(.An(b), .B(f), .C(c), .Y(mai_mai_n372_));
  INV        m0344(.A(mai_mai_n372_), .Y(mai_mai_n373_));
  NOi32      m0345(.An(k), .Bn(h), .C(j), .Y(mai_mai_n374_));
  INV        m0346(.A(mai_mai_n160_), .Y(mai_mai_n375_));
  AOI220     m0347(.A0(mai_mai_n375_), .A1(mai_mai_n373_), .B0(mai_mai_n371_), .B1(mai_mai_n369_), .Y(mai_mai_n376_));
  AN2        m0348(.A(j), .B(h), .Y(mai_mai_n377_));
  OR2        m0349(.A(m), .B(k), .Y(mai_mai_n378_));
  NO2        m0350(.A(mai_mai_n172_), .B(mai_mai_n378_), .Y(mai_mai_n379_));
  NA4        m0351(.A(n), .B(f), .C(c), .D(mai_mai_n114_), .Y(mai_mai_n380_));
  NOi21      m0352(.An(mai_mai_n379_), .B(mai_mai_n380_), .Y(mai_mai_n381_));
  NOi32      m0353(.An(d), .Bn(a), .C(c), .Y(mai_mai_n382_));
  NA2        m0354(.A(mai_mai_n382_), .B(mai_mai_n180_), .Y(mai_mai_n383_));
  NAi21      m0355(.An(i), .B(g), .Y(mai_mai_n384_));
  NAi31      m0356(.An(k), .B(m), .C(j), .Y(mai_mai_n385_));
  NO3        m0357(.A(mai_mai_n385_), .B(mai_mai_n384_), .C(n), .Y(mai_mai_n386_));
  NOi21      m0358(.An(mai_mai_n386_), .B(mai_mai_n383_), .Y(mai_mai_n387_));
  NO2        m0359(.A(mai_mai_n387_), .B(mai_mai_n381_), .Y(mai_mai_n388_));
  NO2        m0360(.A(mai_mai_n380_), .B(mai_mai_n286_), .Y(mai_mai_n389_));
  NOi32      m0361(.An(f), .Bn(d), .C(c), .Y(mai_mai_n390_));
  AOI220     m0362(.A0(mai_mai_n390_), .A1(mai_mai_n296_), .B0(mai_mai_n389_), .B1(mai_mai_n215_), .Y(mai_mai_n391_));
  NA3        m0363(.A(mai_mai_n391_), .B(mai_mai_n388_), .C(mai_mai_n376_), .Y(mai_mai_n392_));
  NO2        m0364(.A(mai_mai_n58_), .B(mai_mai_n114_), .Y(mai_mai_n393_));
  NA2        m0365(.A(mai_mai_n249_), .B(mai_mai_n393_), .Y(mai_mai_n394_));
  INV        m0366(.A(e), .Y(mai_mai_n395_));
  NA2        m0367(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n396_));
  OAI220     m0368(.A0(mai_mai_n396_), .A1(mai_mai_n199_), .B0(mai_mai_n203_), .B1(mai_mai_n395_), .Y(mai_mai_n397_));
  AN2        m0369(.A(g), .B(e), .Y(mai_mai_n398_));
  NA3        m0370(.A(mai_mai_n398_), .B(mai_mai_n202_), .C(i), .Y(mai_mai_n399_));
  INV        m0371(.A(mai_mai_n399_), .Y(mai_mai_n400_));
  NO2        m0372(.A(mai_mai_n98_), .B(mai_mai_n395_), .Y(mai_mai_n401_));
  NO3        m0373(.A(mai_mai_n401_), .B(mai_mai_n400_), .C(mai_mai_n397_), .Y(mai_mai_n402_));
  NOi32      m0374(.An(h), .Bn(e), .C(g), .Y(mai_mai_n403_));
  NA3        m0375(.A(mai_mai_n403_), .B(mai_mai_n280_), .C(m), .Y(mai_mai_n404_));
  NOi21      m0376(.An(g), .B(h), .Y(mai_mai_n405_));
  AN3        m0377(.A(m), .B(l), .C(i), .Y(mai_mai_n406_));
  NA3        m0378(.A(mai_mai_n406_), .B(mai_mai_n405_), .C(e), .Y(mai_mai_n407_));
  AN3        m0379(.A(h), .B(g), .C(e), .Y(mai_mai_n408_));
  NA2        m0380(.A(mai_mai_n408_), .B(mai_mai_n95_), .Y(mai_mai_n409_));
  AN3        m0381(.A(mai_mai_n409_), .B(mai_mai_n407_), .C(mai_mai_n404_), .Y(mai_mai_n410_));
  AOI210     m0382(.A0(mai_mai_n410_), .A1(mai_mai_n402_), .B0(mai_mai_n394_), .Y(mai_mai_n411_));
  NA3        m0383(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(e), .Y(mai_mai_n412_));
  NO2        m0384(.A(mai_mai_n412_), .B(mai_mai_n394_), .Y(mai_mai_n413_));
  NA3        m0385(.A(mai_mai_n382_), .B(mai_mai_n180_), .C(mai_mai_n81_), .Y(mai_mai_n414_));
  NAi31      m0386(.An(b), .B(c), .C(a), .Y(mai_mai_n415_));
  NO2        m0387(.A(mai_mai_n415_), .B(n), .Y(mai_mai_n416_));
  OAI210     m0388(.A0(mai_mai_n51_), .A1(mai_mai_n50_), .B0(m), .Y(mai_mai_n417_));
  NO2        m0389(.A(mai_mai_n417_), .B(mai_mai_n146_), .Y(mai_mai_n418_));
  NA2        m0390(.A(mai_mai_n418_), .B(mai_mai_n416_), .Y(mai_mai_n419_));
  INV        m0391(.A(mai_mai_n419_), .Y(mai_mai_n420_));
  NO4        m0392(.A(mai_mai_n420_), .B(mai_mai_n413_), .C(mai_mai_n411_), .D(mai_mai_n392_), .Y(mai_mai_n421_));
  NA2        m0393(.A(i), .B(g), .Y(mai_mai_n422_));
  NO3        m0394(.A(mai_mai_n268_), .B(mai_mai_n422_), .C(c), .Y(mai_mai_n423_));
  NOi21      m0395(.An(a), .B(n), .Y(mai_mai_n424_));
  NOi21      m0396(.An(d), .B(c), .Y(mai_mai_n425_));
  NA2        m0397(.A(mai_mai_n425_), .B(mai_mai_n424_), .Y(mai_mai_n426_));
  NA3        m0398(.A(i), .B(g), .C(f), .Y(mai_mai_n427_));
  OR2        m0399(.A(mai_mai_n427_), .B(mai_mai_n67_), .Y(mai_mai_n428_));
  NA2        m0400(.A(mai_mai_n406_), .B(mai_mai_n405_), .Y(mai_mai_n429_));
  AOI210     m0401(.A0(mai_mai_n429_), .A1(mai_mai_n428_), .B0(mai_mai_n426_), .Y(mai_mai_n430_));
  AOI210     m0402(.A0(mai_mai_n423_), .A1(mai_mai_n279_), .B0(mai_mai_n430_), .Y(mai_mai_n431_));
  OR2        m0403(.A(n), .B(m), .Y(mai_mai_n432_));
  NO2        m0404(.A(mai_mai_n432_), .B(mai_mai_n151_), .Y(mai_mai_n433_));
  NO2        m0405(.A(mai_mai_n181_), .B(mai_mai_n146_), .Y(mai_mai_n434_));
  OAI210     m0406(.A0(mai_mai_n433_), .A1(mai_mai_n174_), .B0(mai_mai_n434_), .Y(mai_mai_n435_));
  NO2        m0407(.A(mai_mai_n415_), .B(mai_mai_n49_), .Y(mai_mai_n436_));
  NAi21      m0408(.An(k), .B(j), .Y(mai_mai_n437_));
  NAi21      m0409(.An(e), .B(d), .Y(mai_mai_n438_));
  NO2        m0410(.A(mai_mai_n251_), .B(mai_mai_n213_), .Y(mai_mai_n439_));
  NA3        m0411(.A(mai_mai_n439_), .B(d), .C(mai_mai_n227_), .Y(mai_mai_n440_));
  NA2        m0412(.A(mai_mai_n440_), .B(mai_mai_n435_), .Y(mai_mai_n441_));
  NO2        m0413(.A(mai_mai_n323_), .B(mai_mai_n213_), .Y(mai_mai_n442_));
  NA2        m0414(.A(mai_mai_n442_), .B(d), .Y(mai_mai_n443_));
  NOi31      m0415(.An(n), .B(m), .C(k), .Y(mai_mai_n444_));
  AOI220     m0416(.A0(mai_mai_n444_), .A1(mai_mai_n377_), .B0(mai_mai_n221_), .B1(mai_mai_n50_), .Y(mai_mai_n445_));
  NAi31      m0417(.An(g), .B(f), .C(c), .Y(mai_mai_n446_));
  NA2        m0418(.A(mai_mai_n443_), .B(mai_mai_n297_), .Y(mai_mai_n447_));
  NOi31      m0419(.An(mai_mai_n431_), .B(mai_mai_n447_), .C(mai_mai_n441_), .Y(mai_mai_n448_));
  NOi32      m0420(.An(c), .Bn(a), .C(b), .Y(mai_mai_n449_));
  NA2        m0421(.A(mai_mai_n449_), .B(mai_mai_n111_), .Y(mai_mai_n450_));
  INV        m0422(.A(mai_mai_n267_), .Y(mai_mai_n451_));
  AN2        m0423(.A(e), .B(d), .Y(mai_mai_n452_));
  NA2        m0424(.A(mai_mai_n452_), .B(mai_mai_n451_), .Y(mai_mai_n453_));
  INV        m0425(.A(mai_mai_n146_), .Y(mai_mai_n454_));
  NO2        m0426(.A(mai_mai_n129_), .B(mai_mai_n41_), .Y(mai_mai_n455_));
  NO2        m0427(.A(mai_mai_n64_), .B(e), .Y(mai_mai_n456_));
  AOI210     m0428(.A0(mai_mai_n455_), .A1(mai_mai_n454_), .B0(mai_mai_n456_), .Y(mai_mai_n457_));
  AOI210     m0429(.A0(mai_mai_n457_), .A1(mai_mai_n453_), .B0(mai_mai_n450_), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n209_), .B(mai_mai_n204_), .Y(mai_mai_n459_));
  NOi21      m0431(.An(a), .B(b), .Y(mai_mai_n460_));
  NA3        m0432(.A(e), .B(d), .C(c), .Y(mai_mai_n461_));
  NAi21      m0433(.An(mai_mai_n461_), .B(mai_mai_n460_), .Y(mai_mai_n462_));
  NO2        m0434(.A(mai_mai_n414_), .B(mai_mai_n203_), .Y(mai_mai_n463_));
  NOi21      m0435(.An(mai_mai_n462_), .B(mai_mai_n463_), .Y(mai_mai_n464_));
  AOI210     m0436(.A0(mai_mai_n260_), .A1(mai_mai_n459_), .B0(mai_mai_n464_), .Y(mai_mai_n465_));
  NO4        m0437(.A(mai_mai_n186_), .B(mai_mai_n101_), .C(mai_mai_n55_), .D(b), .Y(mai_mai_n466_));
  NA2        m0438(.A(mai_mai_n373_), .B(mai_mai_n152_), .Y(mai_mai_n467_));
  OR2        m0439(.A(k), .B(j), .Y(mai_mai_n468_));
  NA2        m0440(.A(l), .B(k), .Y(mai_mai_n469_));
  NA3        m0441(.A(mai_mai_n469_), .B(mai_mai_n468_), .C(mai_mai_n221_), .Y(mai_mai_n470_));
  AOI210     m0442(.A0(mai_mai_n233_), .A1(mai_mai_n326_), .B0(mai_mai_n81_), .Y(mai_mai_n471_));
  NOi21      m0443(.An(mai_mai_n470_), .B(mai_mai_n471_), .Y(mai_mai_n472_));
  NA2        m0444(.A(mai_mai_n270_), .B(mai_mai_n125_), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n382_), .B(mai_mai_n111_), .Y(mai_mai_n474_));
  NO3        m0446(.A(mai_mai_n474_), .B(mai_mai_n92_), .C(mai_mai_n110_), .Y(mai_mai_n475_));
  NO3        m0447(.A(mai_mai_n414_), .B(mai_mai_n89_), .C(mai_mai_n129_), .Y(mai_mai_n476_));
  NO3        m0448(.A(mai_mai_n476_), .B(mai_mai_n475_), .C(mai_mai_n473_), .Y(mai_mai_n477_));
  NA2        m0449(.A(mai_mai_n477_), .B(mai_mai_n467_), .Y(mai_mai_n478_));
  NO4        m0450(.A(mai_mai_n478_), .B(mai_mai_n466_), .C(mai_mai_n465_), .D(mai_mai_n458_), .Y(mai_mai_n479_));
  NOi21      m0451(.An(d), .B(e), .Y(mai_mai_n480_));
  NAi31      m0452(.An(j), .B(l), .C(i), .Y(mai_mai_n481_));
  OAI210     m0453(.A0(mai_mai_n481_), .A1(mai_mai_n130_), .B0(mai_mai_n101_), .Y(mai_mai_n482_));
  NO3        m0454(.A(mai_mai_n383_), .B(mai_mai_n334_), .C(mai_mai_n200_), .Y(mai_mai_n483_));
  NO2        m0455(.A(mai_mai_n383_), .B(mai_mai_n363_), .Y(mai_mai_n484_));
  NO4        m0456(.A(mai_mai_n484_), .B(mai_mai_n483_), .C(mai_mai_n183_), .D(mai_mai_n294_), .Y(mai_mai_n485_));
  NA2        m0457(.A(mai_mai_n485_), .B(mai_mai_n242_), .Y(mai_mai_n486_));
  OAI210     m0458(.A0(mai_mai_n126_), .A1(mai_mai_n124_), .B0(n), .Y(mai_mai_n487_));
  NO2        m0459(.A(mai_mai_n487_), .B(mai_mai_n129_), .Y(mai_mai_n488_));
  OA210      m0460(.A0(mai_mai_n287_), .A1(mai_mai_n488_), .B0(mai_mai_n191_), .Y(mai_mai_n489_));
  XO2        m0461(.A(i), .B(h), .Y(mai_mai_n490_));
  NA3        m0462(.A(mai_mai_n490_), .B(mai_mai_n159_), .C(n), .Y(mai_mai_n491_));
  NAi31      m0463(.An(mai_mai_n287_), .B(mai_mai_n491_), .C(mai_mai_n445_), .Y(mai_mai_n492_));
  NAi31      m0464(.An(c), .B(f), .C(d), .Y(mai_mai_n493_));
  NO2        m0465(.A(mai_mai_n194_), .B(mai_mai_n493_), .Y(mai_mai_n494_));
  BUFFER     m0466(.A(mai_mai_n79_), .Y(mai_mai_n495_));
  NA3        m0467(.A(mai_mai_n371_), .B(mai_mai_n95_), .C(mai_mai_n94_), .Y(mai_mai_n496_));
  NA2        m0468(.A(mai_mai_n228_), .B(mai_mai_n106_), .Y(mai_mai_n497_));
  AOI210     m0469(.A0(mai_mai_n350_), .A1(mai_mai_n35_), .B0(mai_mai_n462_), .Y(mai_mai_n498_));
  NOi21      m0470(.An(mai_mai_n496_), .B(mai_mai_n498_), .Y(mai_mai_n499_));
  NA3        m0471(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n500_));
  INV        m0472(.A(mai_mai_n283_), .Y(mai_mai_n501_));
  NA3        m0473(.A(mai_mai_n501_), .B(mai_mai_n499_), .C(mai_mai_n495_), .Y(mai_mai_n502_));
  NO3        m0474(.A(mai_mai_n502_), .B(mai_mai_n489_), .C(mai_mai_n486_), .Y(mai_mai_n503_));
  NA4        m0475(.A(mai_mai_n503_), .B(mai_mai_n479_), .C(mai_mai_n448_), .D(mai_mai_n421_), .Y(mai11));
  NO2        m0476(.A(mai_mai_n69_), .B(f), .Y(mai_mai_n505_));
  NA2        m0477(.A(j), .B(g), .Y(mai_mai_n506_));
  NAi31      m0478(.An(i), .B(m), .C(l), .Y(mai_mai_n507_));
  NA3        m0479(.A(m), .B(k), .C(j), .Y(mai_mai_n508_));
  OAI220     m0480(.A0(mai_mai_n508_), .A1(mai_mai_n129_), .B0(mai_mai_n507_), .B1(mai_mai_n506_), .Y(mai_mai_n509_));
  NA2        m0481(.A(mai_mai_n509_), .B(mai_mai_n505_), .Y(mai_mai_n510_));
  NOi32      m0482(.An(e), .Bn(b), .C(f), .Y(mai_mai_n511_));
  NA2        m0483(.A(mai_mai_n256_), .B(mai_mai_n111_), .Y(mai_mai_n512_));
  NA2        m0484(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n513_));
  NO2        m0485(.A(mai_mai_n513_), .B(mai_mai_n289_), .Y(mai_mai_n514_));
  NAi31      m0486(.An(d), .B(e), .C(a), .Y(mai_mai_n515_));
  NO2        m0487(.A(mai_mai_n515_), .B(n), .Y(mai_mai_n516_));
  AOI220     m0488(.A0(mai_mai_n516_), .A1(mai_mai_n99_), .B0(mai_mai_n514_), .B1(mai_mai_n511_), .Y(mai_mai_n517_));
  NAi41      m0489(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n518_));
  AN2        m0490(.A(mai_mai_n518_), .B(mai_mai_n362_), .Y(mai_mai_n519_));
  AOI210     m0491(.A0(mai_mai_n519_), .A1(mai_mai_n383_), .B0(mai_mai_n263_), .Y(mai_mai_n520_));
  NA2        m0492(.A(j), .B(i), .Y(mai_mai_n521_));
  NAi31      m0493(.An(n), .B(m), .C(k), .Y(mai_mai_n522_));
  NO3        m0494(.A(mai_mai_n522_), .B(mai_mai_n521_), .C(mai_mai_n110_), .Y(mai_mai_n523_));
  NO4        m0495(.A(n), .B(d), .C(mai_mai_n114_), .D(a), .Y(mai_mai_n524_));
  OR2        m0496(.A(n), .B(c), .Y(mai_mai_n525_));
  NO2        m0497(.A(mai_mai_n525_), .B(mai_mai_n148_), .Y(mai_mai_n526_));
  NO2        m0498(.A(mai_mai_n526_), .B(mai_mai_n524_), .Y(mai_mai_n527_));
  AOI220     m0499(.A0(g), .A1(mai_mai_n97_), .B0(mai_mai_n509_), .B1(f), .Y(mai_mai_n528_));
  NO2        m0500(.A(mai_mai_n528_), .B(mai_mai_n527_), .Y(mai_mai_n529_));
  AOI210     m0501(.A0(mai_mai_n523_), .A1(mai_mai_n520_), .B0(mai_mai_n529_), .Y(mai_mai_n530_));
  NA2        m0502(.A(mai_mai_n139_), .B(mai_mai_n34_), .Y(mai_mai_n531_));
  OAI220     m0503(.A0(mai_mai_n531_), .A1(m), .B0(mai_mai_n513_), .B1(mai_mai_n233_), .Y(mai_mai_n532_));
  NOi41      m0504(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n533_));
  NAi32      m0505(.An(e), .Bn(b), .C(c), .Y(mai_mai_n534_));
  OR2        m0506(.A(mai_mai_n534_), .B(mai_mai_n81_), .Y(mai_mai_n535_));
  AN2        m0507(.A(mai_mai_n327_), .B(mai_mai_n307_), .Y(mai_mai_n536_));
  NA2        m0508(.A(mai_mai_n536_), .B(mai_mai_n535_), .Y(mai_mai_n537_));
  OA210      m0509(.A0(mai_mai_n537_), .A1(mai_mai_n533_), .B0(mai_mai_n532_), .Y(mai_mai_n538_));
  OAI220     m0510(.A0(mai_mai_n385_), .A1(mai_mai_n384_), .B0(mai_mai_n507_), .B1(mai_mai_n506_), .Y(mai_mai_n539_));
  NAi31      m0511(.An(d), .B(c), .C(a), .Y(mai_mai_n540_));
  NO2        m0512(.A(mai_mai_n540_), .B(n), .Y(mai_mai_n541_));
  NA3        m0513(.A(mai_mai_n541_), .B(mai_mai_n539_), .C(e), .Y(mai_mai_n542_));
  NO3        m0514(.A(mai_mai_n61_), .B(mai_mai_n49_), .C(mai_mai_n214_), .Y(mai_mai_n543_));
  NO2        m0515(.A(mai_mai_n231_), .B(mai_mai_n108_), .Y(mai_mai_n544_));
  OAI210     m0516(.A0(mai_mai_n543_), .A1(mai_mai_n386_), .B0(mai_mai_n544_), .Y(mai_mai_n545_));
  NA2        m0517(.A(mai_mai_n545_), .B(mai_mai_n542_), .Y(mai_mai_n546_));
  NO2        m0518(.A(mai_mai_n268_), .B(n), .Y(mai_mai_n547_));
  NO2        m0519(.A(mai_mai_n416_), .B(mai_mai_n547_), .Y(mai_mai_n548_));
  NA2        m0520(.A(mai_mai_n539_), .B(f), .Y(mai_mai_n549_));
  NAi32      m0521(.An(d), .Bn(a), .C(b), .Y(mai_mai_n550_));
  NO2        m0522(.A(mai_mai_n550_), .B(mai_mai_n49_), .Y(mai_mai_n551_));
  NA2        m0523(.A(h), .B(f), .Y(mai_mai_n552_));
  NO2        m0524(.A(mai_mai_n552_), .B(mai_mai_n92_), .Y(mai_mai_n553_));
  NO3        m0525(.A(mai_mai_n175_), .B(mai_mai_n172_), .C(g), .Y(mai_mai_n554_));
  NA2        m0526(.A(mai_mai_n554_), .B(mai_mai_n57_), .Y(mai_mai_n555_));
  OAI210     m0527(.A0(mai_mai_n549_), .A1(mai_mai_n548_), .B0(mai_mai_n555_), .Y(mai_mai_n556_));
  AN3        m0528(.A(j), .B(h), .C(g), .Y(mai_mai_n557_));
  NO2        m0529(.A(mai_mai_n145_), .B(c), .Y(mai_mai_n558_));
  NA3        m0530(.A(mai_mai_n558_), .B(mai_mai_n557_), .C(mai_mai_n444_), .Y(mai_mai_n559_));
  NA3        m0531(.A(f), .B(d), .C(b), .Y(mai_mai_n560_));
  NO4        m0532(.A(mai_mai_n560_), .B(mai_mai_n175_), .C(mai_mai_n172_), .D(g), .Y(mai_mai_n561_));
  NAi21      m0533(.An(mai_mai_n561_), .B(mai_mai_n559_), .Y(mai_mai_n562_));
  NO4        m0534(.A(mai_mai_n562_), .B(mai_mai_n556_), .C(mai_mai_n546_), .D(mai_mai_n538_), .Y(mai_mai_n563_));
  AN4        m0535(.A(mai_mai_n563_), .B(mai_mai_n530_), .C(mai_mai_n517_), .D(mai_mai_n510_), .Y(mai_mai_n564_));
  INV        m0536(.A(k), .Y(mai_mai_n565_));
  NA3        m0537(.A(l), .B(mai_mai_n565_), .C(i), .Y(mai_mai_n566_));
  INV        m0538(.A(mai_mai_n566_), .Y(mai_mai_n567_));
  NA3        m0539(.A(mai_mai_n382_), .B(mai_mai_n405_), .C(mai_mai_n111_), .Y(mai_mai_n568_));
  NAi32      m0540(.An(h), .Bn(f), .C(g), .Y(mai_mai_n569_));
  NAi41      m0541(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n570_));
  OAI210     m0542(.A0(mai_mai_n515_), .A1(n), .B0(mai_mai_n570_), .Y(mai_mai_n571_));
  NA2        m0543(.A(mai_mai_n571_), .B(m), .Y(mai_mai_n572_));
  NAi31      m0544(.An(h), .B(g), .C(f), .Y(mai_mai_n573_));
  OR3        m0545(.A(mai_mai_n573_), .B(mai_mai_n268_), .C(mai_mai_n49_), .Y(mai_mai_n574_));
  NA4        m0546(.A(mai_mai_n405_), .B(mai_mai_n119_), .C(mai_mai_n111_), .D(e), .Y(mai_mai_n575_));
  AN2        m0547(.A(mai_mai_n575_), .B(mai_mai_n574_), .Y(mai_mai_n576_));
  OA210      m0548(.A0(mai_mai_n572_), .A1(mai_mai_n569_), .B0(mai_mai_n576_), .Y(mai_mai_n577_));
  NO3        m0549(.A(mai_mai_n569_), .B(mai_mai_n69_), .C(mai_mai_n70_), .Y(mai_mai_n578_));
  NO4        m0550(.A(mai_mai_n573_), .B(mai_mai_n525_), .C(mai_mai_n148_), .D(mai_mai_n70_), .Y(mai_mai_n579_));
  OR2        m0551(.A(mai_mai_n579_), .B(mai_mai_n578_), .Y(mai_mai_n580_));
  NAi31      m0552(.An(mai_mai_n580_), .B(mai_mai_n577_), .C(mai_mai_n568_), .Y(mai_mai_n581_));
  NAi31      m0553(.An(f), .B(h), .C(g), .Y(mai_mai_n582_));
  NO4        m0554(.A(mai_mai_n299_), .B(mai_mai_n582_), .C(mai_mai_n69_), .D(mai_mai_n70_), .Y(mai_mai_n583_));
  NOi21      m0555(.An(b), .B(c), .Y(mai_mai_n584_));
  NOi41      m0556(.An(mai_mai_n584_), .B(mai_mai_n343_), .C(mai_mai_n66_), .D(mai_mai_n115_), .Y(mai_mai_n585_));
  OR2        m0557(.A(mai_mai_n585_), .B(mai_mai_n583_), .Y(mai_mai_n586_));
  NOi32      m0558(.An(d), .Bn(a), .C(e), .Y(mai_mai_n587_));
  NA2        m0559(.A(mai_mai_n587_), .B(mai_mai_n111_), .Y(mai_mai_n588_));
  NO2        m0560(.A(n), .B(c), .Y(mai_mai_n589_));
  NA3        m0561(.A(mai_mai_n589_), .B(mai_mai_n29_), .C(m), .Y(mai_mai_n590_));
  NAi32      m0562(.An(n), .Bn(f), .C(m), .Y(mai_mai_n591_));
  NA3        m0563(.A(mai_mai_n591_), .B(mai_mai_n590_), .C(mai_mai_n588_), .Y(mai_mai_n592_));
  NOi32      m0564(.An(e), .Bn(a), .C(d), .Y(mai_mai_n593_));
  AOI210     m0565(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n593_), .Y(mai_mai_n594_));
  AOI210     m0566(.A0(mai_mai_n594_), .A1(mai_mai_n213_), .B0(mai_mai_n531_), .Y(mai_mai_n595_));
  AOI210     m0567(.A0(mai_mai_n595_), .A1(mai_mai_n592_), .B0(mai_mai_n586_), .Y(mai_mai_n596_));
  OAI210     m0568(.A0(mai_mai_n248_), .A1(mai_mai_n84_), .B0(mai_mai_n596_), .Y(mai_mai_n597_));
  AOI210     m0569(.A0(mai_mai_n581_), .A1(mai_mai_n567_), .B0(mai_mai_n597_), .Y(mai_mai_n598_));
  NO3        m0570(.A(mai_mai_n305_), .B(mai_mai_n60_), .C(n), .Y(mai_mai_n599_));
  NA3        m0571(.A(mai_mai_n493_), .B(mai_mai_n170_), .C(mai_mai_n169_), .Y(mai_mai_n600_));
  NA2        m0572(.A(mai_mai_n446_), .B(mai_mai_n231_), .Y(mai_mai_n601_));
  BUFFER     m0573(.A(mai_mai_n601_), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n71_), .B(mai_mai_n111_), .Y(mai_mai_n603_));
  NO2        m0575(.A(mai_mai_n603_), .B(mai_mai_n45_), .Y(mai_mai_n604_));
  AOI220     m0576(.A0(mai_mai_n604_), .A1(mai_mai_n520_), .B0(mai_mai_n602_), .B1(mai_mai_n599_), .Y(mai_mai_n605_));
  NO2        m0577(.A(mai_mai_n605_), .B(mai_mai_n84_), .Y(mai_mai_n606_));
  NA3        m0578(.A(mai_mai_n533_), .B(mai_mai_n329_), .C(mai_mai_n46_), .Y(mai_mai_n607_));
  NOi32      m0579(.An(e), .Bn(c), .C(f), .Y(mai_mai_n608_));
  INV        m0580(.A(mai_mai_n211_), .Y(mai_mai_n609_));
  AOI220     m0581(.A0(mai_mai_n609_), .A1(mai_mai_n379_), .B0(mai_mai_n608_), .B1(mai_mai_n174_), .Y(mai_mai_n610_));
  NA3        m0582(.A(mai_mai_n610_), .B(mai_mai_n607_), .C(mai_mai_n177_), .Y(mai_mai_n611_));
  AOI210     m0583(.A0(mai_mai_n519_), .A1(mai_mai_n383_), .B0(mai_mai_n288_), .Y(mai_mai_n612_));
  NA2        m0584(.A(mai_mai_n612_), .B(mai_mai_n258_), .Y(mai_mai_n613_));
  NOi21      m0585(.An(j), .B(l), .Y(mai_mai_n614_));
  NAi21      m0586(.An(k), .B(h), .Y(mai_mai_n615_));
  NO2        m0587(.A(mai_mai_n615_), .B(mai_mai_n257_), .Y(mai_mai_n616_));
  NA2        m0588(.A(mai_mai_n616_), .B(mai_mai_n614_), .Y(mai_mai_n617_));
  OR2        m0589(.A(mai_mai_n617_), .B(mai_mai_n572_), .Y(mai_mai_n618_));
  NOi31      m0590(.An(m), .B(n), .C(k), .Y(mai_mai_n619_));
  NA2        m0591(.A(mai_mai_n614_), .B(mai_mai_n619_), .Y(mai_mai_n620_));
  AOI210     m0592(.A0(mai_mai_n383_), .A1(mai_mai_n362_), .B0(mai_mai_n288_), .Y(mai_mai_n621_));
  NAi21      m0593(.An(mai_mai_n620_), .B(mai_mai_n621_), .Y(mai_mai_n622_));
  NO2        m0594(.A(mai_mai_n268_), .B(mai_mai_n49_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n299_), .B(mai_mai_n582_), .Y(mai_mai_n624_));
  NO2        m0596(.A(mai_mai_n515_), .B(mai_mai_n49_), .Y(mai_mai_n625_));
  AOI220     m0597(.A0(mai_mai_n625_), .A1(mai_mai_n624_), .B0(mai_mai_n623_), .B1(mai_mai_n553_), .Y(mai_mai_n626_));
  NA4        m0598(.A(mai_mai_n626_), .B(mai_mai_n622_), .C(mai_mai_n618_), .D(mai_mai_n613_), .Y(mai_mai_n627_));
  NA2        m0599(.A(mai_mai_n106_), .B(mai_mai_n36_), .Y(mai_mai_n628_));
  NO2        m0600(.A(mai_mai_n511_), .B(mai_mai_n352_), .Y(mai_mai_n629_));
  NO2        m0601(.A(mai_mai_n629_), .B(n), .Y(mai_mai_n630_));
  NAi31      m0602(.An(mai_mai_n628_), .B(mai_mai_n630_), .C(g), .Y(mai_mai_n631_));
  NO2        m0603(.A(mai_mai_n513_), .B(mai_mai_n175_), .Y(mai_mai_n632_));
  NA2        m0604(.A(mai_mai_n490_), .B(mai_mai_n159_), .Y(mai_mai_n633_));
  NO3        m0605(.A(mai_mai_n380_), .B(mai_mai_n633_), .C(mai_mai_n84_), .Y(mai_mai_n634_));
  AOI210     m0606(.A0(c), .A1(mai_mai_n632_), .B0(mai_mai_n634_), .Y(mai_mai_n635_));
  AN3        m0607(.A(f), .B(d), .C(b), .Y(mai_mai_n636_));
  NA3        m0608(.A(mai_mai_n490_), .B(mai_mai_n159_), .C(mai_mai_n214_), .Y(mai_mai_n637_));
  NO2        m0609(.A(mai_mai_n232_), .B(mai_mai_n637_), .Y(mai_mai_n638_));
  NAi31      m0610(.An(m), .B(n), .C(k), .Y(mai_mai_n639_));
  OR2        m0611(.A(mai_mai_n133_), .B(mai_mai_n60_), .Y(mai_mai_n640_));
  NO2        m0612(.A(mai_mai_n640_), .B(mai_mai_n639_), .Y(mai_mai_n641_));
  OAI210     m0613(.A0(mai_mai_n641_), .A1(mai_mai_n638_), .B0(j), .Y(mai_mai_n642_));
  NA3        m0614(.A(mai_mai_n642_), .B(mai_mai_n635_), .C(mai_mai_n631_), .Y(mai_mai_n643_));
  NO4        m0615(.A(mai_mai_n643_), .B(mai_mai_n627_), .C(mai_mai_n611_), .D(mai_mai_n606_), .Y(mai_mai_n644_));
  NA2        m0616(.A(mai_mai_n371_), .B(mai_mai_n162_), .Y(mai_mai_n645_));
  NAi31      m0617(.An(g), .B(h), .C(f), .Y(mai_mai_n646_));
  OR3        m0618(.A(mai_mai_n646_), .B(mai_mai_n268_), .C(n), .Y(mai_mai_n647_));
  OA210      m0619(.A0(mai_mai_n515_), .A1(n), .B0(mai_mai_n570_), .Y(mai_mai_n648_));
  NA3        m0620(.A(mai_mai_n403_), .B(mai_mai_n119_), .C(mai_mai_n81_), .Y(mai_mai_n649_));
  OAI210     m0621(.A0(mai_mai_n648_), .A1(mai_mai_n88_), .B0(mai_mai_n649_), .Y(mai_mai_n650_));
  NOi21      m0622(.An(mai_mai_n647_), .B(mai_mai_n650_), .Y(mai_mai_n651_));
  AOI210     m0623(.A0(mai_mai_n651_), .A1(mai_mai_n645_), .B0(mai_mai_n508_), .Y(mai_mai_n652_));
  NO3        m0624(.A(g), .B(mai_mai_n213_), .C(mai_mai_n55_), .Y(mai_mai_n653_));
  NO2        m0625(.A(mai_mai_n497_), .B(mai_mai_n84_), .Y(mai_mai_n654_));
  OAI210     m0626(.A0(mai_mai_n654_), .A1(mai_mai_n379_), .B0(mai_mai_n653_), .Y(mai_mai_n655_));
  NA2        m0627(.A(mai_mai_n584_), .B(mai_mai_n331_), .Y(mai_mai_n656_));
  OA220      m0628(.A0(mai_mai_n620_), .A1(mai_mai_n656_), .B0(mai_mai_n617_), .B1(mai_mai_n69_), .Y(mai_mai_n657_));
  NA3        m0629(.A(mai_mai_n505_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n658_));
  NA2        m0630(.A(h), .B(mai_mai_n37_), .Y(mai_mai_n659_));
  NA2        m0631(.A(mai_mai_n97_), .B(mai_mai_n46_), .Y(mai_mai_n660_));
  OAI220     m0632(.A0(mai_mai_n660_), .A1(mai_mai_n320_), .B0(mai_mai_n659_), .B1(mai_mai_n450_), .Y(mai_mai_n661_));
  AOI210     m0633(.A0(mai_mai_n550_), .A1(mai_mai_n415_), .B0(mai_mai_n49_), .Y(mai_mai_n662_));
  OAI220     m0634(.A0(mai_mai_n573_), .A1(mai_mai_n566_), .B0(mai_mai_n313_), .B1(mai_mai_n506_), .Y(mai_mai_n663_));
  AOI210     m0635(.A0(mai_mai_n663_), .A1(mai_mai_n662_), .B0(mai_mai_n661_), .Y(mai_mai_n664_));
  NA4        m0636(.A(mai_mai_n664_), .B(mai_mai_n658_), .C(mai_mai_n657_), .D(mai_mai_n655_), .Y(mai_mai_n665_));
  NO2        m0637(.A(mai_mai_n250_), .B(f), .Y(mai_mai_n666_));
  INV        m0638(.A(mai_mai_n60_), .Y(mai_mai_n667_));
  NO3        m0639(.A(mai_mai_n667_), .B(mai_mai_n666_), .C(mai_mai_n34_), .Y(mai_mai_n668_));
  NA2        m0640(.A(mai_mai_n316_), .B(mai_mai_n139_), .Y(mai_mai_n669_));
  NA2        m0641(.A(mai_mai_n130_), .B(mai_mai_n49_), .Y(mai_mai_n670_));
  AOI220     m0642(.A0(mai_mai_n670_), .A1(mai_mai_n511_), .B0(mai_mai_n352_), .B1(mai_mai_n111_), .Y(mai_mai_n671_));
  OA220      m0643(.A0(mai_mai_n671_), .A1(mai_mai_n531_), .B0(mai_mai_n350_), .B1(mai_mai_n109_), .Y(mai_mai_n672_));
  OAI210     m0644(.A0(mai_mai_n669_), .A1(mai_mai_n668_), .B0(mai_mai_n672_), .Y(mai_mai_n673_));
  NO3        m0645(.A(mai_mai_n390_), .B(mai_mai_n191_), .C(mai_mai_n190_), .Y(mai_mai_n674_));
  NA2        m0646(.A(mai_mai_n674_), .B(mai_mai_n231_), .Y(mai_mai_n675_));
  NA3        m0647(.A(mai_mai_n675_), .B(mai_mai_n252_), .C(j), .Y(mai_mai_n676_));
  NA2        m0648(.A(mai_mai_n449_), .B(mai_mai_n81_), .Y(mai_mai_n677_));
  NO3        m0649(.A(mai_mai_n508_), .B(mai_mai_n677_), .C(mai_mai_n129_), .Y(mai_mai_n678_));
  INV        m0650(.A(mai_mai_n678_), .Y(mai_mai_n679_));
  NA4        m0651(.A(mai_mai_n679_), .B(mai_mai_n676_), .C(mai_mai_n496_), .D(mai_mai_n388_), .Y(mai_mai_n680_));
  NO4        m0652(.A(mai_mai_n680_), .B(mai_mai_n673_), .C(mai_mai_n665_), .D(mai_mai_n652_), .Y(mai_mai_n681_));
  NA4        m0653(.A(mai_mai_n681_), .B(mai_mai_n644_), .C(mai_mai_n598_), .D(mai_mai_n564_), .Y(mai08));
  NO2        m0654(.A(k), .B(h), .Y(mai_mai_n683_));
  AO210      m0655(.A0(mai_mai_n250_), .A1(mai_mai_n437_), .B0(mai_mai_n683_), .Y(mai_mai_n684_));
  NO2        m0656(.A(mai_mai_n684_), .B(mai_mai_n286_), .Y(mai_mai_n685_));
  NA2        m0657(.A(mai_mai_n608_), .B(mai_mai_n81_), .Y(mai_mai_n686_));
  INV        m0658(.A(mai_mai_n686_), .Y(mai_mai_n687_));
  AOI210     m0659(.A0(mai_mai_n687_), .A1(mai_mai_n685_), .B0(mai_mai_n476_), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n81_), .B(mai_mai_n108_), .Y(mai_mai_n689_));
  NO2        m0661(.A(mai_mai_n689_), .B(mai_mai_n56_), .Y(mai_mai_n690_));
  NO4        m0662(.A(mai_mai_n368_), .B(mai_mai_n110_), .C(j), .D(mai_mai_n214_), .Y(mai_mai_n691_));
  NA2        m0663(.A(mai_mai_n560_), .B(mai_mai_n232_), .Y(mai_mai_n692_));
  AOI220     m0664(.A0(mai_mai_n692_), .A1(mai_mai_n337_), .B0(mai_mai_n691_), .B1(mai_mai_n690_), .Y(mai_mai_n693_));
  AOI210     m0665(.A0(mai_mai_n560_), .A1(mai_mai_n155_), .B0(mai_mai_n81_), .Y(mai_mai_n694_));
  NA4        m0666(.A(mai_mai_n216_), .B(mai_mai_n139_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n695_));
  AN2        m0667(.A(l), .B(k), .Y(mai_mai_n696_));
  NA4        m0668(.A(mai_mai_n696_), .B(mai_mai_n106_), .C(mai_mai_n70_), .D(mai_mai_n214_), .Y(mai_mai_n697_));
  OAI210     m0669(.A0(mai_mai_n695_), .A1(g), .B0(mai_mai_n697_), .Y(mai_mai_n698_));
  NA2        m0670(.A(mai_mai_n698_), .B(mai_mai_n694_), .Y(mai_mai_n699_));
  NA4        m0671(.A(mai_mai_n699_), .B(mai_mai_n693_), .C(mai_mai_n688_), .D(mai_mai_n339_), .Y(mai_mai_n700_));
  AN2        m0672(.A(mai_mai_n516_), .B(mai_mai_n93_), .Y(mai_mai_n701_));
  NO4        m0673(.A(mai_mai_n172_), .B(mai_mai_n378_), .C(mai_mai_n110_), .D(g), .Y(mai_mai_n702_));
  NA2        m0674(.A(mai_mai_n702_), .B(mai_mai_n692_), .Y(mai_mai_n703_));
  INV        m0675(.A(mai_mai_n38_), .Y(mai_mai_n704_));
  AOI220     m0676(.A0(mai_mai_n609_), .A1(mai_mai_n336_), .B0(mai_mai_n704_), .B1(mai_mai_n547_), .Y(mai_mai_n705_));
  NAi31      m0677(.An(mai_mai_n701_), .B(mai_mai_n705_), .C(mai_mai_n703_), .Y(mai_mai_n706_));
  NO2        m0678(.A(mai_mai_n519_), .B(mai_mai_n35_), .Y(mai_mai_n707_));
  OAI210     m0679(.A0(mai_mai_n534_), .A1(mai_mai_n47_), .B0(mai_mai_n640_), .Y(mai_mai_n708_));
  NO2        m0680(.A(mai_mai_n469_), .B(mai_mai_n130_), .Y(mai_mai_n709_));
  AOI210     m0681(.A0(mai_mai_n709_), .A1(mai_mai_n708_), .B0(mai_mai_n707_), .Y(mai_mai_n710_));
  NO3        m0682(.A(mai_mai_n305_), .B(mai_mai_n129_), .C(mai_mai_n41_), .Y(mai_mai_n711_));
  NAi21      m0683(.An(mai_mai_n711_), .B(mai_mai_n697_), .Y(mai_mai_n712_));
  NA2        m0684(.A(mai_mai_n684_), .B(mai_mai_n134_), .Y(mai_mai_n713_));
  AOI220     m0685(.A0(mai_mai_n713_), .A1(mai_mai_n389_), .B0(mai_mai_n712_), .B1(mai_mai_n73_), .Y(mai_mai_n714_));
  NA2        m0686(.A(mai_mai_n710_), .B(mai_mai_n714_), .Y(mai_mai_n715_));
  NA2        m0687(.A(mai_mai_n352_), .B(mai_mai_n43_), .Y(mai_mai_n716_));
  NA3        m0688(.A(mai_mai_n675_), .B(mai_mai_n322_), .C(mai_mai_n374_), .Y(mai_mai_n717_));
  NA2        m0689(.A(mai_mai_n696_), .B(mai_mai_n221_), .Y(mai_mai_n718_));
  NO2        m0690(.A(mai_mai_n718_), .B(mai_mai_n315_), .Y(mai_mai_n719_));
  AOI210     m0691(.A0(mai_mai_n719_), .A1(mai_mai_n666_), .B0(mai_mai_n475_), .Y(mai_mai_n720_));
  NA3        m0692(.A(m), .B(l), .C(k), .Y(mai_mai_n721_));
  AOI210     m0693(.A0(mai_mai_n649_), .A1(mai_mai_n647_), .B0(mai_mai_n721_), .Y(mai_mai_n722_));
  NO2        m0694(.A(mai_mai_n518_), .B(mai_mai_n263_), .Y(mai_mai_n723_));
  NOi21      m0695(.An(mai_mai_n723_), .B(mai_mai_n512_), .Y(mai_mai_n724_));
  NA4        m0696(.A(mai_mai_n111_), .B(l), .C(k), .D(mai_mai_n84_), .Y(mai_mai_n725_));
  NO2        m0697(.A(mai_mai_n724_), .B(mai_mai_n722_), .Y(mai_mai_n726_));
  NA4        m0698(.A(mai_mai_n726_), .B(mai_mai_n720_), .C(mai_mai_n717_), .D(mai_mai_n716_), .Y(mai_mai_n727_));
  NO4        m0699(.A(mai_mai_n727_), .B(mai_mai_n715_), .C(mai_mai_n706_), .D(mai_mai_n700_), .Y(mai_mai_n728_));
  NA2        m0700(.A(mai_mai_n609_), .B(mai_mai_n379_), .Y(mai_mai_n729_));
  NOi31      m0701(.An(g), .B(h), .C(f), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n625_), .B(mai_mai_n730_), .Y(mai_mai_n731_));
  AO210      m0703(.A0(mai_mai_n731_), .A1(mai_mai_n574_), .B0(mai_mai_n521_), .Y(mai_mai_n732_));
  NO3        m0704(.A(mai_mai_n383_), .B(mai_mai_n506_), .C(h), .Y(mai_mai_n733_));
  AOI210     m0705(.A0(mai_mai_n733_), .A1(mai_mai_n111_), .B0(mai_mai_n484_), .Y(mai_mai_n734_));
  NA4        m0706(.A(mai_mai_n734_), .B(mai_mai_n732_), .C(mai_mai_n729_), .D(mai_mai_n248_), .Y(mai_mai_n735_));
  NA2        m0707(.A(mai_mai_n696_), .B(mai_mai_n70_), .Y(mai_mai_n736_));
  NOi21      m0708(.An(h), .B(j), .Y(mai_mai_n737_));
  NA2        m0709(.A(mai_mai_n737_), .B(f), .Y(mai_mai_n738_));
  NO2        m0710(.A(mai_mai_n738_), .B(mai_mai_n245_), .Y(mai_mai_n739_));
  INV        m0711(.A(mai_mai_n739_), .Y(mai_mai_n740_));
  OAI220     m0712(.A0(mai_mai_n740_), .A1(mai_mai_n736_), .B0(mai_mai_n576_), .B1(mai_mai_n61_), .Y(mai_mai_n741_));
  AOI210     m0713(.A0(mai_mai_n735_), .A1(l), .B0(mai_mai_n741_), .Y(mai_mai_n742_));
  NO2        m0714(.A(j), .B(i), .Y(mai_mai_n743_));
  NA3        m0715(.A(mai_mai_n743_), .B(mai_mai_n77_), .C(l), .Y(mai_mai_n744_));
  NA2        m0716(.A(mai_mai_n743_), .B(mai_mai_n33_), .Y(mai_mai_n745_));
  NA2        m0717(.A(mai_mai_n408_), .B(mai_mai_n119_), .Y(mai_mai_n746_));
  OA220      m0718(.A0(mai_mai_n746_), .A1(mai_mai_n745_), .B0(mai_mai_n744_), .B1(mai_mai_n572_), .Y(mai_mai_n747_));
  NO3        m0719(.A(mai_mai_n150_), .B(mai_mai_n49_), .C(mai_mai_n108_), .Y(mai_mai_n748_));
  NO3        m0720(.A(mai_mai_n525_), .B(mai_mai_n148_), .C(mai_mai_n70_), .Y(mai_mai_n749_));
  NO3        m0721(.A(mai_mai_n469_), .B(mai_mai_n427_), .C(j), .Y(mai_mai_n750_));
  OAI210     m0722(.A0(mai_mai_n749_), .A1(mai_mai_n748_), .B0(mai_mai_n750_), .Y(mai_mai_n751_));
  OAI210     m0723(.A0(mai_mai_n731_), .A1(mai_mai_n61_), .B0(mai_mai_n751_), .Y(mai_mai_n752_));
  INV        m0724(.A(j), .Y(mai_mai_n753_));
  NO3        m0725(.A(mai_mai_n286_), .B(mai_mai_n753_), .C(mai_mai_n40_), .Y(mai_mai_n754_));
  AOI210     m0726(.A0(mai_mai_n511_), .A1(n), .B0(mai_mai_n533_), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n755_), .B(mai_mai_n536_), .Y(mai_mai_n756_));
  AN3        m0728(.A(mai_mai_n756_), .B(mai_mai_n754_), .C(mai_mai_n96_), .Y(mai_mai_n757_));
  NO3        m0729(.A(mai_mai_n172_), .B(mai_mai_n378_), .C(mai_mai_n110_), .Y(mai_mai_n758_));
  AOI220     m0730(.A0(mai_mai_n758_), .A1(mai_mai_n246_), .B0(mai_mai_n601_), .B1(mai_mai_n296_), .Y(mai_mai_n759_));
  NAi31      m0731(.An(mai_mai_n594_), .B(mai_mai_n90_), .C(mai_mai_n81_), .Y(mai_mai_n760_));
  NA2        m0732(.A(mai_mai_n760_), .B(mai_mai_n759_), .Y(mai_mai_n761_));
  NO2        m0733(.A(mai_mai_n286_), .B(mai_mai_n134_), .Y(mai_mai_n762_));
  AOI220     m0734(.A0(mai_mai_n762_), .A1(mai_mai_n609_), .B0(mai_mai_n711_), .B1(mai_mai_n694_), .Y(mai_mai_n763_));
  NO2        m0735(.A(mai_mai_n721_), .B(mai_mai_n88_), .Y(mai_mai_n764_));
  NA2        m0736(.A(mai_mai_n764_), .B(mai_mai_n571_), .Y(mai_mai_n765_));
  NO2        m0737(.A(mai_mai_n573_), .B(mai_mai_n115_), .Y(mai_mai_n766_));
  OAI210     m0738(.A0(mai_mai_n766_), .A1(mai_mai_n750_), .B0(mai_mai_n662_), .Y(mai_mai_n767_));
  NA3        m0739(.A(mai_mai_n767_), .B(mai_mai_n765_), .C(mai_mai_n763_), .Y(mai_mai_n768_));
  OR4        m0740(.A(mai_mai_n768_), .B(mai_mai_n761_), .C(mai_mai_n757_), .D(mai_mai_n752_), .Y(mai_mai_n769_));
  NA3        m0741(.A(mai_mai_n755_), .B(mai_mai_n536_), .C(mai_mai_n535_), .Y(mai_mai_n770_));
  NA4        m0742(.A(mai_mai_n770_), .B(mai_mai_n216_), .C(mai_mai_n437_), .D(mai_mai_n34_), .Y(mai_mai_n771_));
  NO4        m0743(.A(mai_mai_n469_), .B(mai_mai_n422_), .C(j), .D(f), .Y(mai_mai_n772_));
  OAI220     m0744(.A0(mai_mai_n695_), .A1(mai_mai_n686_), .B0(mai_mai_n320_), .B1(mai_mai_n38_), .Y(mai_mai_n773_));
  AOI210     m0745(.A0(mai_mai_n772_), .A1(mai_mai_n255_), .B0(mai_mai_n773_), .Y(mai_mai_n774_));
  NA3        m0746(.A(g), .B(mai_mai_n280_), .C(h), .Y(mai_mai_n775_));
  NOi21      m0747(.An(mai_mai_n662_), .B(mai_mai_n775_), .Y(mai_mai_n776_));
  NO2        m0748(.A(mai_mai_n89_), .B(mai_mai_n47_), .Y(mai_mai_n777_));
  OAI220     m0749(.A0(mai_mai_n775_), .A1(mai_mai_n590_), .B0(mai_mai_n744_), .B1(mai_mai_n69_), .Y(mai_mai_n778_));
  AOI210     m0750(.A0(mai_mai_n777_), .A1(mai_mai_n630_), .B0(mai_mai_n778_), .Y(mai_mai_n779_));
  NAi41      m0751(.An(mai_mai_n776_), .B(mai_mai_n779_), .C(mai_mai_n774_), .D(mai_mai_n771_), .Y(mai_mai_n780_));
  AOI220     m0752(.A0(mai_mai_n764_), .A1(mai_mai_n238_), .B0(mai_mai_n750_), .B1(mai_mai_n623_), .Y(mai_mai_n781_));
  NO2        m0753(.A(mai_mai_n648_), .B(mai_mai_n70_), .Y(mai_mai_n782_));
  AOI210     m0754(.A0(mai_mai_n772_), .A1(mai_mai_n782_), .B0(mai_mai_n324_), .Y(mai_mai_n783_));
  OAI210     m0755(.A0(mai_mai_n721_), .A1(mai_mai_n646_), .B0(mai_mai_n500_), .Y(mai_mai_n784_));
  NA3        m0756(.A(mai_mai_n249_), .B(mai_mai_n58_), .C(b), .Y(mai_mai_n785_));
  AOI220     m0757(.A0(mai_mai_n589_), .A1(mai_mai_n29_), .B0(mai_mai_n449_), .B1(mai_mai_n81_), .Y(mai_mai_n786_));
  NA2        m0758(.A(mai_mai_n786_), .B(mai_mai_n785_), .Y(mai_mai_n787_));
  NO2        m0759(.A(mai_mai_n775_), .B(mai_mai_n474_), .Y(mai_mai_n788_));
  AOI210     m0760(.A0(mai_mai_n787_), .A1(mai_mai_n784_), .B0(mai_mai_n788_), .Y(mai_mai_n789_));
  NA3        m0761(.A(mai_mai_n789_), .B(mai_mai_n783_), .C(mai_mai_n781_), .Y(mai_mai_n790_));
  NOi41      m0762(.An(mai_mai_n747_), .B(mai_mai_n790_), .C(mai_mai_n780_), .D(mai_mai_n769_), .Y(mai_mai_n791_));
  OR2        m0763(.A(mai_mai_n695_), .B(mai_mai_n232_), .Y(mai_mai_n792_));
  NO3        m0764(.A(mai_mai_n330_), .B(mai_mai_n288_), .C(mai_mai_n110_), .Y(mai_mai_n793_));
  NA2        m0765(.A(mai_mai_n793_), .B(mai_mai_n756_), .Y(mai_mai_n794_));
  INV        m0766(.A(mai_mai_n46_), .Y(mai_mai_n795_));
  NO3        m0767(.A(mai_mai_n795_), .B(mai_mai_n745_), .C(mai_mai_n268_), .Y(mai_mai_n796_));
  NO3        m0768(.A(mai_mai_n506_), .B(mai_mai_n91_), .C(h), .Y(mai_mai_n797_));
  AOI210     m0769(.A0(mai_mai_n797_), .A1(mai_mai_n690_), .B0(mai_mai_n796_), .Y(mai_mai_n798_));
  NA4        m0770(.A(mai_mai_n798_), .B(mai_mai_n794_), .C(mai_mai_n792_), .D(mai_mai_n391_), .Y(mai_mai_n799_));
  OR2        m0771(.A(mai_mai_n646_), .B(mai_mai_n89_), .Y(mai_mai_n800_));
  NOi31      m0772(.An(b), .B(d), .C(a), .Y(mai_mai_n801_));
  NO2        m0773(.A(mai_mai_n801_), .B(mai_mai_n587_), .Y(mai_mai_n802_));
  NO2        m0774(.A(mai_mai_n802_), .B(n), .Y(mai_mai_n803_));
  NOi21      m0775(.An(mai_mai_n786_), .B(mai_mai_n803_), .Y(mai_mai_n804_));
  NO2        m0776(.A(mai_mai_n804_), .B(mai_mai_n800_), .Y(mai_mai_n805_));
  NO2        m0777(.A(mai_mai_n534_), .B(mai_mai_n81_), .Y(mai_mai_n806_));
  NO2        m0778(.A(mai_mai_n315_), .B(mai_mai_n115_), .Y(mai_mai_n807_));
  NOi21      m0779(.An(mai_mai_n807_), .B(mai_mai_n160_), .Y(mai_mai_n808_));
  AOI210     m0780(.A0(mai_mai_n793_), .A1(mai_mai_n806_), .B0(mai_mai_n808_), .Y(mai_mai_n809_));
  OAI210     m0781(.A0(mai_mai_n695_), .A1(mai_mai_n380_), .B0(mai_mai_n809_), .Y(mai_mai_n810_));
  NO2        m0782(.A(mai_mai_n674_), .B(n), .Y(mai_mai_n811_));
  NA2        m0783(.A(mai_mai_n811_), .B(mai_mai_n685_), .Y(mai_mai_n812_));
  NO2        m0784(.A(mai_mai_n310_), .B(mai_mai_n237_), .Y(mai_mai_n813_));
  OAI210     m0785(.A0(mai_mai_n93_), .A1(mai_mai_n90_), .B0(mai_mai_n813_), .Y(mai_mai_n814_));
  NA2        m0786(.A(mai_mai_n119_), .B(mai_mai_n81_), .Y(mai_mai_n815_));
  AOI210     m0787(.A0(mai_mai_n412_), .A1(mai_mai_n404_), .B0(mai_mai_n815_), .Y(mai_mai_n816_));
  NAi21      m0788(.An(mai_mai_n816_), .B(mai_mai_n814_), .Y(mai_mai_n817_));
  NA2        m0789(.A(mai_mai_n719_), .B(mai_mai_n34_), .Y(mai_mai_n818_));
  NAi21      m0790(.An(mai_mai_n725_), .B(mai_mai_n423_), .Y(mai_mai_n819_));
  NO2        m0791(.A(mai_mai_n263_), .B(i), .Y(mai_mai_n820_));
  NA2        m0792(.A(mai_mai_n702_), .B(mai_mai_n338_), .Y(mai_mai_n821_));
  OAI210     m0793(.A0(mai_mai_n579_), .A1(mai_mai_n578_), .B0(l), .Y(mai_mai_n822_));
  AN3        m0794(.A(mai_mai_n822_), .B(mai_mai_n821_), .C(mai_mai_n819_), .Y(mai_mai_n823_));
  NAi41      m0795(.An(mai_mai_n817_), .B(mai_mai_n823_), .C(mai_mai_n818_), .D(mai_mai_n812_), .Y(mai_mai_n824_));
  NO4        m0796(.A(mai_mai_n824_), .B(mai_mai_n810_), .C(mai_mai_n805_), .D(mai_mai_n799_), .Y(mai_mai_n825_));
  NA4        m0797(.A(mai_mai_n825_), .B(mai_mai_n791_), .C(mai_mai_n742_), .D(mai_mai_n728_), .Y(mai09));
  INV        m0798(.A(mai_mai_n120_), .Y(mai_mai_n827_));
  NA2        m0799(.A(f), .B(e), .Y(mai_mai_n828_));
  NO2        m0800(.A(mai_mai_n226_), .B(mai_mai_n110_), .Y(mai_mai_n829_));
  NA2        m0801(.A(mai_mai_n829_), .B(g), .Y(mai_mai_n830_));
  NA4        m0802(.A(mai_mai_n299_), .B(l), .C(i), .D(mai_mai_n117_), .Y(mai_mai_n831_));
  AOI210     m0803(.A0(mai_mai_n831_), .A1(g), .B0(mai_mai_n455_), .Y(mai_mai_n832_));
  AOI210     m0804(.A0(mai_mai_n832_), .A1(mai_mai_n830_), .B0(mai_mai_n828_), .Y(mai_mai_n833_));
  NA2        m0805(.A(mai_mai_n833_), .B(mai_mai_n827_), .Y(mai_mai_n834_));
  NO2        m0806(.A(mai_mai_n203_), .B(mai_mai_n213_), .Y(mai_mai_n835_));
  NA3        m0807(.A(m), .B(l), .C(i), .Y(mai_mai_n836_));
  OAI220     m0808(.A0(mai_mai_n573_), .A1(mai_mai_n836_), .B0(mai_mai_n343_), .B1(mai_mai_n507_), .Y(mai_mai_n837_));
  NA4        m0809(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .D(f), .Y(mai_mai_n838_));
  NAi31      m0810(.An(mai_mai_n837_), .B(mai_mai_n838_), .C(mai_mai_n428_), .Y(mai_mai_n839_));
  OR2        m0811(.A(mai_mai_n839_), .B(mai_mai_n835_), .Y(mai_mai_n840_));
  NA3        m0812(.A(mai_mai_n800_), .B(mai_mai_n549_), .C(mai_mai_n500_), .Y(mai_mai_n841_));
  OA210      m0813(.A0(mai_mai_n841_), .A1(mai_mai_n840_), .B0(mai_mai_n803_), .Y(mai_mai_n842_));
  INV        m0814(.A(mai_mai_n327_), .Y(mai_mai_n843_));
  NO2        m0815(.A(mai_mai_n126_), .B(mai_mai_n124_), .Y(mai_mai_n844_));
  NOi31      m0816(.An(k), .B(m), .C(l), .Y(mai_mai_n845_));
  NO2        m0817(.A(m), .B(mai_mai_n582_), .Y(mai_mai_n846_));
  NA2        m0818(.A(mai_mai_n785_), .B(mai_mai_n320_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n331_), .B(mai_mai_n333_), .Y(mai_mai_n848_));
  OAI210     m0820(.A0(mai_mai_n203_), .A1(mai_mai_n213_), .B0(mai_mai_n848_), .Y(mai_mai_n849_));
  AOI220     m0821(.A0(mai_mai_n849_), .A1(mai_mai_n847_), .B0(mai_mai_n846_), .B1(mai_mai_n843_), .Y(mai_mai_n850_));
  NA2        m0822(.A(mai_mai_n166_), .B(mai_mai_n112_), .Y(mai_mai_n851_));
  NA3        m0823(.A(mai_mai_n851_), .B(mai_mai_n684_), .C(mai_mai_n134_), .Y(mai_mai_n852_));
  NA3        m0824(.A(mai_mai_n852_), .B(mai_mai_n188_), .C(mai_mai_n31_), .Y(mai_mai_n853_));
  NA4        m0825(.A(mai_mai_n853_), .B(mai_mai_n850_), .C(mai_mai_n610_), .D(mai_mai_n79_), .Y(mai_mai_n854_));
  NO2        m0826(.A(mai_mai_n569_), .B(mai_mai_n481_), .Y(mai_mai_n855_));
  NA2        m0827(.A(mai_mai_n855_), .B(mai_mai_n188_), .Y(mai_mai_n856_));
  NOi21      m0828(.An(f), .B(d), .Y(mai_mai_n857_));
  NA2        m0829(.A(mai_mai_n857_), .B(m), .Y(mai_mai_n858_));
  NO2        m0830(.A(mai_mai_n858_), .B(mai_mai_n52_), .Y(mai_mai_n859_));
  NOi32      m0831(.An(g), .Bn(f), .C(d), .Y(mai_mai_n860_));
  NA4        m0832(.A(mai_mai_n860_), .B(mai_mai_n589_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n861_));
  NOi21      m0833(.An(mai_mai_n300_), .B(mai_mai_n861_), .Y(mai_mai_n862_));
  AOI210     m0834(.A0(mai_mai_n859_), .A1(mai_mai_n526_), .B0(mai_mai_n862_), .Y(mai_mai_n863_));
  AN2        m0835(.A(f), .B(d), .Y(mai_mai_n864_));
  NA3        m0836(.A(mai_mai_n460_), .B(mai_mai_n864_), .C(mai_mai_n81_), .Y(mai_mai_n865_));
  NO3        m0837(.A(mai_mai_n865_), .B(mai_mai_n70_), .C(mai_mai_n214_), .Y(mai_mai_n866_));
  INV        m0838(.A(mai_mai_n274_), .Y(mai_mai_n867_));
  INV        m0839(.A(mai_mai_n866_), .Y(mai_mai_n868_));
  NAi41      m0840(.An(mai_mai_n473_), .B(mai_mai_n868_), .C(mai_mai_n863_), .D(mai_mai_n856_), .Y(mai_mai_n869_));
  NO3        m0841(.A(mai_mai_n130_), .B(mai_mai_n315_), .C(mai_mai_n151_), .Y(mai_mai_n870_));
  NO2        m0842(.A(mai_mai_n639_), .B(mai_mai_n315_), .Y(mai_mai_n871_));
  AN2        m0843(.A(mai_mai_n871_), .B(mai_mai_n666_), .Y(mai_mai_n872_));
  NO3        m0844(.A(mai_mai_n872_), .B(mai_mai_n870_), .C(mai_mai_n234_), .Y(mai_mai_n873_));
  NA2        m0845(.A(mai_mai_n587_), .B(mai_mai_n81_), .Y(mai_mai_n874_));
  NO2        m0846(.A(mai_mai_n848_), .B(mai_mai_n874_), .Y(mai_mai_n875_));
  NA3        m0847(.A(mai_mai_n159_), .B(mai_mai_n106_), .C(g), .Y(mai_mai_n876_));
  OAI220     m0848(.A0(mai_mai_n865_), .A1(mai_mai_n417_), .B0(mai_mai_n327_), .B1(mai_mai_n876_), .Y(mai_mai_n877_));
  NOi41      m0849(.An(mai_mai_n224_), .B(mai_mai_n877_), .C(mai_mai_n875_), .D(mai_mai_n294_), .Y(mai_mai_n878_));
  NA2        m0850(.A(c), .B(mai_mai_n114_), .Y(mai_mai_n879_));
  NO2        m0851(.A(mai_mai_n879_), .B(mai_mai_n395_), .Y(mai_mai_n880_));
  NA3        m0852(.A(mai_mai_n880_), .B(mai_mai_n492_), .C(f), .Y(mai_mai_n881_));
  OR2        m0853(.A(mai_mai_n646_), .B(mai_mai_n522_), .Y(mai_mai_n882_));
  INV        m0854(.A(mai_mai_n882_), .Y(mai_mai_n883_));
  NA2        m0855(.A(mai_mai_n802_), .B(mai_mai_n109_), .Y(mai_mai_n884_));
  NA2        m0856(.A(mai_mai_n884_), .B(mai_mai_n883_), .Y(mai_mai_n885_));
  NA4        m0857(.A(mai_mai_n885_), .B(mai_mai_n881_), .C(mai_mai_n878_), .D(mai_mai_n873_), .Y(mai_mai_n886_));
  NO4        m0858(.A(mai_mai_n886_), .B(mai_mai_n869_), .C(mai_mai_n854_), .D(mai_mai_n842_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n281_), .B(mai_mai_n865_), .Y(mai_mai_n888_));
  NO2        m0860(.A(mai_mai_n134_), .B(mai_mai_n130_), .Y(mai_mai_n889_));
  NO2        m0861(.A(mai_mai_n231_), .B(mai_mai_n225_), .Y(mai_mai_n890_));
  AOI220     m0862(.A0(mai_mai_n890_), .A1(mai_mai_n228_), .B0(mai_mai_n293_), .B1(mai_mai_n889_), .Y(mai_mai_n891_));
  NO2        m0863(.A(mai_mai_n417_), .B(mai_mai_n828_), .Y(mai_mai_n892_));
  NA2        m0864(.A(mai_mai_n892_), .B(mai_mai_n541_), .Y(mai_mai_n893_));
  NA2        m0865(.A(mai_mai_n893_), .B(mai_mai_n891_), .Y(mai_mai_n894_));
  NA2        m0866(.A(e), .B(d), .Y(mai_mai_n895_));
  OAI220     m0867(.A0(mai_mai_n895_), .A1(c), .B0(mai_mai_n310_), .B1(d), .Y(mai_mai_n896_));
  NA3        m0868(.A(mai_mai_n896_), .B(mai_mai_n439_), .C(mai_mai_n490_), .Y(mai_mai_n897_));
  AOI210     m0869(.A0(mai_mai_n497_), .A1(mai_mai_n179_), .B0(mai_mai_n231_), .Y(mai_mai_n898_));
  AOI210     m0870(.A0(mai_mai_n609_), .A1(mai_mai_n336_), .B0(mai_mai_n898_), .Y(mai_mai_n899_));
  NA3        m0871(.A(mai_mai_n165_), .B(mai_mai_n82_), .C(mai_mai_n34_), .Y(mai_mai_n900_));
  NA3        m0872(.A(mai_mai_n900_), .B(mai_mai_n899_), .C(mai_mai_n897_), .Y(mai_mai_n901_));
  NO3        m0873(.A(mai_mai_n901_), .B(mai_mai_n894_), .C(mai_mai_n888_), .Y(mai_mai_n902_));
  NA2        m0874(.A(mai_mai_n843_), .B(mai_mai_n31_), .Y(mai_mai_n903_));
  AO210      m0875(.A0(mai_mai_n903_), .A1(mai_mai_n686_), .B0(mai_mai_n217_), .Y(mai_mai_n904_));
  OAI210     m0876(.A0(mai_mai_n288_), .A1(j), .B0(mai_mai_n60_), .Y(mai_mai_n905_));
  AOI220     m0877(.A0(mai_mai_n905_), .A1(mai_mai_n871_), .B0(mai_mai_n599_), .B1(mai_mai_n608_), .Y(mai_mai_n906_));
  INV        m0878(.A(mai_mai_n906_), .Y(mai_mai_n907_));
  OAI210     m0879(.A0(mai_mai_n829_), .A1(mai_mai_n1434_), .B0(mai_mai_n860_), .Y(mai_mai_n908_));
  NO2        m0880(.A(mai_mai_n908_), .B(mai_mai_n590_), .Y(mai_mai_n909_));
  AOI210     m0881(.A0(mai_mai_n116_), .A1(mai_mai_n115_), .B0(mai_mai_n256_), .Y(mai_mai_n910_));
  NO2        m0882(.A(mai_mai_n910_), .B(mai_mai_n861_), .Y(mai_mai_n911_));
  AO210      m0883(.A0(mai_mai_n847_), .A1(mai_mai_n837_), .B0(mai_mai_n911_), .Y(mai_mai_n912_));
  NOi31      m0884(.An(mai_mai_n526_), .B(mai_mai_n858_), .C(mai_mai_n281_), .Y(mai_mai_n913_));
  NO4        m0885(.A(mai_mai_n913_), .B(mai_mai_n912_), .C(mai_mai_n909_), .D(mai_mai_n907_), .Y(mai_mai_n914_));
  AO220      m0886(.A0(mai_mai_n439_), .A1(mai_mai_n737_), .B0(mai_mai_n174_), .B1(f), .Y(mai_mai_n915_));
  OAI210     m0887(.A0(mai_mai_n915_), .A1(mai_mai_n442_), .B0(mai_mai_n896_), .Y(mai_mai_n916_));
  NO2        m0888(.A(mai_mai_n427_), .B(mai_mai_n67_), .Y(mai_mai_n917_));
  OAI210     m0889(.A0(mai_mai_n841_), .A1(mai_mai_n917_), .B0(mai_mai_n690_), .Y(mai_mai_n918_));
  AN4        m0890(.A(mai_mai_n918_), .B(mai_mai_n916_), .C(mai_mai_n914_), .D(mai_mai_n904_), .Y(mai_mai_n919_));
  NA4        m0891(.A(mai_mai_n919_), .B(mai_mai_n902_), .C(mai_mai_n887_), .D(mai_mai_n834_), .Y(mai12));
  NO2        m0892(.A(mai_mai_n438_), .B(c), .Y(mai_mai_n921_));
  NO4        m0893(.A(mai_mai_n432_), .B(mai_mai_n250_), .C(mai_mai_n565_), .D(mai_mai_n214_), .Y(mai_mai_n922_));
  NA2        m0894(.A(mai_mai_n922_), .B(mai_mai_n921_), .Y(mai_mai_n923_));
  NA2        m0895(.A(mai_mai_n526_), .B(mai_mai_n917_), .Y(mai_mai_n924_));
  NO2        m0896(.A(mai_mai_n438_), .B(mai_mai_n114_), .Y(mai_mai_n925_));
  NO2        m0897(.A(mai_mai_n844_), .B(mai_mai_n343_), .Y(mai_mai_n926_));
  NO2        m0898(.A(mai_mai_n646_), .B(mai_mai_n368_), .Y(mai_mai_n927_));
  AOI220     m0899(.A0(mai_mai_n927_), .A1(mai_mai_n524_), .B0(mai_mai_n926_), .B1(mai_mai_n925_), .Y(mai_mai_n928_));
  NA4        m0900(.A(mai_mai_n928_), .B(mai_mai_n924_), .C(mai_mai_n923_), .D(mai_mai_n431_), .Y(mai_mai_n929_));
  AOI210     m0901(.A0(mai_mai_n233_), .A1(mai_mai_n326_), .B0(mai_mai_n200_), .Y(mai_mai_n930_));
  BUFFER     m0902(.A(mai_mai_n922_), .Y(mai_mai_n931_));
  NO2        m0903(.A(mai_mai_n323_), .B(mai_mai_n214_), .Y(mai_mai_n932_));
  OAI210     m0904(.A0(mai_mai_n932_), .A1(mai_mai_n931_), .B0(mai_mai_n390_), .Y(mai_mai_n933_));
  NO2        m0905(.A(mai_mai_n628_), .B(mai_mai_n257_), .Y(mai_mai_n934_));
  NO2        m0906(.A(mai_mai_n573_), .B(mai_mai_n836_), .Y(mai_mai_n935_));
  AOI220     m0907(.A0(mai_mai_n935_), .A1(mai_mai_n547_), .B0(mai_mai_n813_), .B1(mai_mai_n934_), .Y(mai_mai_n936_));
  NO2        m0908(.A(mai_mai_n150_), .B(mai_mai_n237_), .Y(mai_mai_n937_));
  NA3        m0909(.A(mai_mai_n937_), .B(mai_mai_n240_), .C(i), .Y(mai_mai_n938_));
  NA3        m0910(.A(mai_mai_n938_), .B(mai_mai_n936_), .C(mai_mai_n933_), .Y(mai_mai_n939_));
  OR2        m0911(.A(mai_mai_n311_), .B(mai_mai_n925_), .Y(mai_mai_n940_));
  NA2        m0912(.A(mai_mai_n940_), .B(mai_mai_n344_), .Y(mai_mai_n941_));
  NO3        m0913(.A(mai_mai_n130_), .B(mai_mai_n151_), .C(mai_mai_n214_), .Y(mai_mai_n942_));
  NA2        m0914(.A(mai_mai_n942_), .B(mai_mai_n511_), .Y(mai_mai_n943_));
  NA4        m0915(.A(mai_mai_n433_), .B(mai_mai_n425_), .C(mai_mai_n180_), .D(g), .Y(mai_mai_n944_));
  NA3        m0916(.A(mai_mai_n944_), .B(mai_mai_n943_), .C(mai_mai_n941_), .Y(mai_mai_n945_));
  NO3        m0917(.A(mai_mai_n651_), .B(mai_mai_n89_), .C(mai_mai_n45_), .Y(mai_mai_n946_));
  NO4        m0918(.A(mai_mai_n946_), .B(mai_mai_n945_), .C(mai_mai_n939_), .D(mai_mai_n929_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n359_), .B(mai_mai_n358_), .Y(mai_mai_n948_));
  NA2        m0920(.A(mai_mai_n570_), .B(mai_mai_n69_), .Y(mai_mai_n949_));
  NOi21      m0921(.An(mai_mai_n34_), .B(mai_mai_n639_), .Y(mai_mai_n950_));
  AOI220     m0922(.A0(mai_mai_n950_), .A1(c), .B0(mai_mai_n949_), .B1(mai_mai_n948_), .Y(mai_mai_n951_));
  INV        m0923(.A(mai_mai_n951_), .Y(mai_mai_n952_));
  NA2        m0924(.A(mai_mai_n423_), .B(mai_mai_n258_), .Y(mai_mai_n953_));
  NO3        m0925(.A(mai_mai_n815_), .B(mai_mai_n86_), .C(mai_mai_n395_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n953_), .B(mai_mai_n309_), .Y(mai_mai_n955_));
  NO2        m0927(.A(mai_mai_n487_), .B(mai_mai_n288_), .Y(mai_mai_n956_));
  INV        m0928(.A(mai_mai_n619_), .Y(mai_mai_n957_));
  INV        m0929(.A(mai_mai_n356_), .Y(mai_mai_n958_));
  NO3        m0930(.A(mai_mai_n958_), .B(mai_mai_n955_), .C(mai_mai_n952_), .Y(mai_mai_n959_));
  NA2        m0931(.A(mai_mai_n336_), .B(g), .Y(mai_mai_n960_));
  NA2        m0932(.A(mai_mai_n162_), .B(i), .Y(mai_mai_n961_));
  NA2        m0933(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n962_));
  OAI220     m0934(.A0(mai_mai_n962_), .A1(mai_mai_n199_), .B0(mai_mai_n961_), .B1(mai_mai_n89_), .Y(mai_mai_n963_));
  AOI210     m0935(.A0(mai_mai_n406_), .A1(mai_mai_n37_), .B0(mai_mai_n963_), .Y(mai_mai_n964_));
  NO2        m0936(.A(mai_mai_n143_), .B(mai_mai_n81_), .Y(mai_mai_n965_));
  OR2        m0937(.A(mai_mai_n965_), .B(mai_mai_n533_), .Y(mai_mai_n966_));
  AOI210     m0938(.A0(c), .A1(n), .B0(mai_mai_n966_), .Y(mai_mai_n967_));
  OAI220     m0939(.A0(mai_mai_n967_), .A1(mai_mai_n960_), .B0(mai_mai_n964_), .B1(mai_mai_n320_), .Y(mai_mai_n968_));
  NO2        m0940(.A(mai_mai_n646_), .B(mai_mai_n481_), .Y(mai_mai_n969_));
  NA3        m0941(.A(mai_mai_n331_), .B(mai_mai_n614_), .C(i), .Y(mai_mai_n970_));
  OAI210     m0942(.A0(mai_mai_n427_), .A1(mai_mai_n299_), .B0(mai_mai_n970_), .Y(mai_mai_n971_));
  OAI220     m0943(.A0(mai_mai_n971_), .A1(mai_mai_n969_), .B0(mai_mai_n662_), .B1(mai_mai_n749_), .Y(mai_mai_n972_));
  NA2        m0944(.A(mai_mai_n593_), .B(mai_mai_n111_), .Y(mai_mai_n973_));
  OR3        m0945(.A(mai_mai_n299_), .B(mai_mai_n422_), .C(f), .Y(mai_mai_n974_));
  NA3        m0946(.A(mai_mai_n614_), .B(mai_mai_n77_), .C(i), .Y(mai_mai_n975_));
  OA220      m0947(.A0(mai_mai_n975_), .A1(mai_mai_n973_), .B0(mai_mai_n974_), .B1(mai_mai_n572_), .Y(mai_mai_n976_));
  NA3        m0948(.A(mai_mai_n312_), .B(mai_mai_n116_), .C(g), .Y(mai_mai_n977_));
  AOI210     m0949(.A0(mai_mai_n659_), .A1(mai_mai_n977_), .B0(m), .Y(mai_mai_n978_));
  OAI210     m0950(.A0(mai_mai_n978_), .A1(mai_mai_n926_), .B0(mai_mai_n311_), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n677_), .B(mai_mai_n874_), .Y(mai_mai_n980_));
  NA2        m0952(.A(mai_mai_n838_), .B(mai_mai_n428_), .Y(mai_mai_n981_));
  NA2        m0953(.A(mai_mai_n222_), .B(mai_mai_n74_), .Y(mai_mai_n982_));
  NA3        m0954(.A(mai_mai_n982_), .B(mai_mai_n975_), .C(mai_mai_n974_), .Y(mai_mai_n983_));
  AOI220     m0955(.A0(mai_mai_n983_), .A1(mai_mai_n255_), .B0(mai_mai_n981_), .B1(mai_mai_n980_), .Y(mai_mai_n984_));
  NA4        m0956(.A(mai_mai_n984_), .B(mai_mai_n979_), .C(mai_mai_n976_), .D(mai_mai_n972_), .Y(mai_mai_n985_));
  NO2        m0957(.A(mai_mai_n368_), .B(mai_mai_n88_), .Y(mai_mai_n986_));
  OAI210     m0958(.A0(mai_mai_n986_), .A1(mai_mai_n934_), .B0(mai_mai_n238_), .Y(mai_mai_n987_));
  NA2        m0959(.A(mai_mai_n650_), .B(mai_mai_n85_), .Y(mai_mai_n988_));
  NO2        m0960(.A(mai_mai_n445_), .B(mai_mai_n214_), .Y(mai_mai_n989_));
  AOI220     m0961(.A0(mai_mai_n989_), .A1(mai_mai_n373_), .B0(mai_mai_n940_), .B1(mai_mai_n218_), .Y(mai_mai_n990_));
  AOI220     m0962(.A0(mai_mai_n927_), .A1(mai_mai_n937_), .B0(mai_mai_n571_), .B1(mai_mai_n87_), .Y(mai_mai_n991_));
  NA4        m0963(.A(mai_mai_n991_), .B(mai_mai_n990_), .C(mai_mai_n988_), .D(mai_mai_n987_), .Y(mai_mai_n992_));
  OAI210     m0964(.A0(mai_mai_n981_), .A1(mai_mai_n935_), .B0(mai_mai_n524_), .Y(mai_mai_n993_));
  AOI210     m0965(.A0(mai_mai_n407_), .A1(mai_mai_n399_), .B0(mai_mai_n815_), .Y(mai_mai_n994_));
  OAI210     m0966(.A0(mai_mai_n359_), .A1(mai_mai_n358_), .B0(mai_mai_n107_), .Y(mai_mai_n995_));
  AOI210     m0967(.A0(mai_mai_n995_), .A1(mai_mai_n516_), .B0(mai_mai_n994_), .Y(mai_mai_n996_));
  NA2        m0968(.A(mai_mai_n978_), .B(mai_mai_n925_), .Y(mai_mai_n997_));
  NO3        m0969(.A(l), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n998_));
  AOI220     m0970(.A0(mai_mai_n998_), .A1(mai_mai_n612_), .B0(mai_mai_n632_), .B1(mai_mai_n511_), .Y(mai_mai_n999_));
  NA4        m0971(.A(mai_mai_n999_), .B(mai_mai_n997_), .C(mai_mai_n996_), .D(mai_mai_n993_), .Y(mai_mai_n1000_));
  NO4        m0972(.A(mai_mai_n1000_), .B(mai_mai_n992_), .C(mai_mai_n985_), .D(mai_mai_n968_), .Y(mai_mai_n1001_));
  NAi31      m0973(.An(mai_mai_n140_), .B(mai_mai_n408_), .C(n), .Y(mai_mai_n1002_));
  NO3        m0974(.A(mai_mai_n124_), .B(mai_mai_n329_), .C(mai_mai_n845_), .Y(mai_mai_n1003_));
  NO2        m0975(.A(mai_mai_n1003_), .B(mai_mai_n1002_), .Y(mai_mai_n1004_));
  NO3        m0976(.A(mai_mai_n263_), .B(mai_mai_n140_), .C(mai_mai_n395_), .Y(mai_mai_n1005_));
  AOI210     m0977(.A0(mai_mai_n1005_), .A1(mai_mai_n482_), .B0(mai_mai_n1004_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n476_), .B(i), .Y(mai_mai_n1007_));
  NA2        m0979(.A(mai_mai_n1007_), .B(mai_mai_n1006_), .Y(mai_mai_n1008_));
  NA2        m0980(.A(mai_mai_n231_), .B(mai_mai_n170_), .Y(mai_mai_n1009_));
  NO3        m0981(.A(mai_mai_n296_), .B(mai_mai_n433_), .C(mai_mai_n174_), .Y(mai_mai_n1010_));
  NOi31      m0982(.An(mai_mai_n1009_), .B(mai_mai_n1010_), .C(mai_mai_n214_), .Y(mai_mai_n1011_));
  NAi21      m0983(.An(mai_mai_n534_), .B(mai_mai_n989_), .Y(mai_mai_n1012_));
  NO3        m0984(.A(mai_mai_n427_), .B(mai_mai_n299_), .C(mai_mai_n70_), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n1013_), .B(mai_mai_n424_), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n1014_), .B(mai_mai_n1012_), .Y(mai_mai_n1015_));
  OAI220     m0987(.A0(mai_mai_n1002_), .A1(mai_mai_n233_), .B0(mai_mai_n970_), .B1(mai_mai_n588_), .Y(mai_mai_n1016_));
  NO2        m0988(.A(mai_mai_n647_), .B(mai_mai_n368_), .Y(mai_mai_n1017_));
  NA2        m0989(.A(mai_mai_n930_), .B(mai_mai_n921_), .Y(mai_mai_n1018_));
  NO2        m0990(.A(mai_mai_n525_), .B(mai_mai_n148_), .Y(mai_mai_n1019_));
  OAI210     m0991(.A0(mai_mai_n1019_), .A1(mai_mai_n505_), .B0(mai_mai_n369_), .Y(mai_mai_n1020_));
  OAI220     m0992(.A0(mai_mai_n927_), .A1(mai_mai_n935_), .B0(mai_mai_n526_), .B1(mai_mai_n416_), .Y(mai_mai_n1021_));
  NA4        m0993(.A(mai_mai_n1021_), .B(mai_mai_n1020_), .C(mai_mai_n1018_), .D(mai_mai_n607_), .Y(mai_mai_n1022_));
  OAI210     m0994(.A0(mai_mai_n930_), .A1(mai_mai_n922_), .B0(mai_mai_n1009_), .Y(mai_mai_n1023_));
  NA3        m0995(.A(c), .B(mai_mai_n471_), .C(mai_mai_n46_), .Y(mai_mai_n1024_));
  AOI210     m0996(.A0(mai_mai_n371_), .A1(mai_mai_n369_), .B0(mai_mai_n319_), .Y(mai_mai_n1025_));
  NA4        m0997(.A(mai_mai_n1025_), .B(mai_mai_n1024_), .C(mai_mai_n1023_), .D(mai_mai_n264_), .Y(mai_mai_n1026_));
  OR4        m0998(.A(mai_mai_n1026_), .B(mai_mai_n1022_), .C(mai_mai_n1017_), .D(mai_mai_n1016_), .Y(mai_mai_n1027_));
  NO4        m0999(.A(mai_mai_n1027_), .B(mai_mai_n1015_), .C(mai_mai_n1011_), .D(mai_mai_n1008_), .Y(mai_mai_n1028_));
  NA4        m1000(.A(mai_mai_n1028_), .B(mai_mai_n1001_), .C(mai_mai_n959_), .D(mai_mai_n947_), .Y(mai13));
  AN2        m1001(.A(c), .B(b), .Y(mai_mai_n1030_));
  NA3        m1002(.A(mai_mai_n249_), .B(mai_mai_n1030_), .C(m), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n480_), .B(f), .Y(mai_mai_n1032_));
  NO3        m1004(.A(mai_mai_n1032_), .B(mai_mai_n1031_), .C(mai_mai_n566_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n139_), .B(mai_mai_n45_), .Y(mai_mai_n1034_));
  NO4        m1006(.A(mai_mai_n1034_), .B(d), .C(mai_mai_n573_), .D(mai_mai_n295_), .Y(mai_mai_n1035_));
  NA2        m1007(.A(mai_mai_n398_), .B(mai_mai_n213_), .Y(mai_mai_n1036_));
  AN2        m1008(.A(d), .B(c), .Y(mai_mai_n1037_));
  NA2        m1009(.A(mai_mai_n1037_), .B(mai_mai_n114_), .Y(mai_mai_n1038_));
  NO4        m1010(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .C(mai_mai_n175_), .D(mai_mai_n166_), .Y(mai_mai_n1039_));
  NA2        m1011(.A(mai_mai_n480_), .B(c), .Y(mai_mai_n1040_));
  NO3        m1012(.A(mai_mai_n1034_), .B(mai_mai_n569_), .C(mai_mai_n295_), .Y(mai_mai_n1041_));
  OR2        m1013(.A(mai_mai_n1039_), .B(mai_mai_n1041_), .Y(mai_mai_n1042_));
  OR3        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1035_), .C(mai_mai_n1033_), .Y(mai_mai_n1043_));
  NO2        m1015(.A(f), .B(mai_mai_n145_), .Y(mai_mai_n1044_));
  NA2        m1016(.A(mai_mai_n1044_), .B(g), .Y(mai_mai_n1045_));
  OR2        m1017(.A(mai_mai_n225_), .B(mai_mai_n175_), .Y(mai_mai_n1046_));
  NO2        m1018(.A(mai_mai_n1046_), .B(mai_mai_n1045_), .Y(mai_mai_n1047_));
  NO2        m1019(.A(mai_mai_n1040_), .B(mai_mai_n295_), .Y(mai_mai_n1048_));
  NA2        m1020(.A(mai_mai_n616_), .B(mai_mai_n1429_), .Y(mai_mai_n1049_));
  NOi21      m1021(.An(mai_mai_n1048_), .B(mai_mai_n1049_), .Y(mai_mai_n1050_));
  NOi41      m1022(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1051_));
  NA2        m1023(.A(mai_mai_n1051_), .B(j), .Y(mai_mai_n1052_));
  NO2        m1024(.A(mai_mai_n1052_), .B(mai_mai_n1045_), .Y(mai_mai_n1053_));
  OR3        m1025(.A(e), .B(d), .C(c), .Y(mai_mai_n1054_));
  NA3        m1026(.A(k), .B(j), .C(i), .Y(mai_mai_n1055_));
  NO3        m1027(.A(mai_mai_n1055_), .B(mai_mai_n295_), .C(mai_mai_n88_), .Y(mai_mai_n1056_));
  NOi21      m1028(.An(mai_mai_n1056_), .B(mai_mai_n1054_), .Y(mai_mai_n1057_));
  OR4        m1029(.A(mai_mai_n1057_), .B(mai_mai_n1053_), .C(mai_mai_n1050_), .D(mai_mai_n1047_), .Y(mai_mai_n1058_));
  NA3        m1030(.A(mai_mai_n452_), .B(mai_mai_n322_), .C(mai_mai_n55_), .Y(mai_mai_n1059_));
  NO2        m1031(.A(mai_mai_n1059_), .B(mai_mai_n1049_), .Y(mai_mai_n1060_));
  NO3        m1032(.A(mai_mai_n1059_), .B(mai_mai_n569_), .C(mai_mai_n437_), .Y(mai_mai_n1061_));
  NO2        m1033(.A(f), .B(c), .Y(mai_mai_n1062_));
  NOi21      m1034(.An(mai_mai_n1062_), .B(mai_mai_n432_), .Y(mai_mai_n1063_));
  NA2        m1035(.A(mai_mai_n1063_), .B(mai_mai_n58_), .Y(mai_mai_n1064_));
  NO3        m1036(.A(i), .B(mai_mai_n243_), .C(l), .Y(mai_mai_n1065_));
  NOi31      m1037(.An(mai_mai_n1065_), .B(mai_mai_n1064_), .C(j), .Y(mai_mai_n1066_));
  OR3        m1038(.A(mai_mai_n1066_), .B(mai_mai_n1061_), .C(mai_mai_n1060_), .Y(mai_mai_n1067_));
  OR3        m1039(.A(mai_mai_n1067_), .B(mai_mai_n1058_), .C(mai_mai_n1043_), .Y(mai02));
  OR3        m1040(.A(h), .B(g), .C(f), .Y(mai_mai_n1069_));
  OR3        m1041(.A(n), .B(m), .C(i), .Y(mai_mai_n1070_));
  NO4        m1042(.A(mai_mai_n1070_), .B(mai_mai_n1069_), .C(l), .D(mai_mai_n1054_), .Y(mai_mai_n1071_));
  NOi31      m1043(.An(e), .B(d), .C(c), .Y(mai_mai_n1072_));
  AOI210     m1044(.A0(mai_mai_n1056_), .A1(mai_mai_n1072_), .B0(mai_mai_n1035_), .Y(mai_mai_n1073_));
  AN3        m1045(.A(g), .B(f), .C(c), .Y(mai_mai_n1074_));
  NA2        m1046(.A(mai_mai_n1074_), .B(mai_mai_n452_), .Y(mai_mai_n1075_));
  BUFFER     m1047(.A(mai_mai_n295_), .Y(mai_mai_n1076_));
  OR2        m1048(.A(mai_mai_n1076_), .B(mai_mai_n1075_), .Y(mai_mai_n1077_));
  NO3        m1049(.A(mai_mai_n1059_), .B(mai_mai_n1034_), .C(mai_mai_n569_), .Y(mai_mai_n1078_));
  NO2        m1050(.A(mai_mai_n1078_), .B(mai_mai_n1047_), .Y(mai_mai_n1079_));
  NA3        m1051(.A(l), .B(k), .C(j), .Y(mai_mai_n1080_));
  NA2        m1052(.A(i), .B(h), .Y(mai_mai_n1081_));
  NO3        m1053(.A(mai_mai_n1081_), .B(mai_mai_n1080_), .C(mai_mai_n130_), .Y(mai_mai_n1082_));
  NO3        m1054(.A(mai_mai_n141_), .B(mai_mai_n272_), .C(mai_mai_n214_), .Y(mai_mai_n1083_));
  AOI210     m1055(.A0(mai_mai_n1083_), .A1(mai_mai_n1082_), .B0(mai_mai_n1050_), .Y(mai_mai_n1084_));
  NA3        m1056(.A(c), .B(b), .C(a), .Y(mai_mai_n1085_));
  NO3        m1057(.A(mai_mai_n1085_), .B(mai_mai_n895_), .C(mai_mai_n213_), .Y(mai_mai_n1086_));
  NO3        m1058(.A(mai_mai_n288_), .B(mai_mai_n49_), .C(mai_mai_n110_), .Y(mai_mai_n1087_));
  AOI210     m1059(.A0(mai_mai_n1087_), .A1(mai_mai_n1086_), .B0(mai_mai_n1060_), .Y(mai_mai_n1088_));
  AN4        m1060(.A(mai_mai_n1088_), .B(mai_mai_n1084_), .C(mai_mai_n1079_), .D(mai_mai_n1077_), .Y(mai_mai_n1089_));
  NO2        m1061(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .Y(mai_mai_n1090_));
  NA2        m1062(.A(mai_mai_n1052_), .B(mai_mai_n1046_), .Y(mai_mai_n1091_));
  AOI210     m1063(.A0(mai_mai_n1091_), .A1(mai_mai_n1090_), .B0(mai_mai_n1033_), .Y(mai_mai_n1092_));
  NAi41      m1064(.An(mai_mai_n1071_), .B(mai_mai_n1092_), .C(mai_mai_n1089_), .D(mai_mai_n1073_), .Y(mai03));
  NO2        m1065(.A(mai_mai_n507_), .B(mai_mai_n582_), .Y(mai_mai_n1094_));
  NA4        m1066(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(g), .D(mai_mai_n213_), .Y(mai_mai_n1095_));
  NA4        m1067(.A(mai_mai_n557_), .B(m), .C(mai_mai_n110_), .D(mai_mai_n213_), .Y(mai_mai_n1096_));
  NA3        m1068(.A(mai_mai_n1096_), .B(mai_mai_n360_), .C(mai_mai_n1095_), .Y(mai_mai_n1097_));
  NO3        m1069(.A(mai_mai_n1097_), .B(mai_mai_n1094_), .C(mai_mai_n995_), .Y(mai_mai_n1098_));
  NOi41      m1070(.An(mai_mai_n800_), .B(mai_mai_n849_), .C(mai_mai_n839_), .D(mai_mai_n704_), .Y(mai_mai_n1099_));
  OAI220     m1071(.A0(mai_mai_n1099_), .A1(mai_mai_n677_), .B0(mai_mai_n1098_), .B1(mai_mai_n570_), .Y(mai_mai_n1100_));
  NA4        m1072(.A(i), .B(mai_mai_n1072_), .C(mai_mai_n331_), .D(mai_mai_n322_), .Y(mai_mai_n1101_));
  OAI210     m1073(.A0(mai_mai_n815_), .A1(mai_mai_n409_), .B0(mai_mai_n1101_), .Y(mai_mai_n1102_));
  NOi31      m1074(.An(m), .B(n), .C(f), .Y(mai_mai_n1103_));
  NA2        m1075(.A(mai_mai_n1103_), .B(mai_mai_n51_), .Y(mai_mai_n1104_));
  NA2        m1076(.A(c), .B(a), .Y(mai_mai_n1105_));
  OAI220     m1077(.A0(mai_mai_n1105_), .A1(mai_mai_n1104_), .B0(mai_mai_n882_), .B1(mai_mai_n415_), .Y(mai_mai_n1106_));
  NOi31      m1078(.An(mai_mai_n860_), .B(mai_mai_n1031_), .C(h), .Y(mai_mai_n1107_));
  NO4        m1079(.A(mai_mai_n1107_), .B(mai_mai_n1106_), .C(mai_mai_n1102_), .D(mai_mai_n994_), .Y(mai_mai_n1108_));
  NO2        m1080(.A(mai_mai_n272_), .B(a), .Y(mai_mai_n1109_));
  INV        m1081(.A(mai_mai_n1035_), .Y(mai_mai_n1110_));
  NO2        m1082(.A(mai_mai_n1081_), .B(mai_mai_n469_), .Y(mai_mai_n1111_));
  NO2        m1083(.A(mai_mai_n84_), .B(g), .Y(mai_mai_n1112_));
  AOI210     m1084(.A0(mai_mai_n1112_), .A1(mai_mai_n1111_), .B0(mai_mai_n1065_), .Y(mai_mai_n1113_));
  OR2        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1064_), .Y(mai_mai_n1114_));
  NA3        m1086(.A(mai_mai_n1114_), .B(mai_mai_n1110_), .C(mai_mai_n1108_), .Y(mai_mai_n1115_));
  NO4        m1087(.A(mai_mai_n1115_), .B(mai_mai_n1100_), .C(mai_mai_n817_), .D(mai_mai_n546_), .Y(mai_mai_n1116_));
  NA2        m1088(.A(c), .B(b), .Y(mai_mai_n1117_));
  NO2        m1089(.A(mai_mai_n689_), .B(mai_mai_n1117_), .Y(mai_mai_n1118_));
  OAI210     m1090(.A0(mai_mai_n858_), .A1(mai_mai_n832_), .B0(mai_mai_n402_), .Y(mai_mai_n1119_));
  OAI210     m1091(.A0(mai_mai_n1119_), .A1(mai_mai_n859_), .B0(mai_mai_n1118_), .Y(mai_mai_n1120_));
  NAi21      m1092(.An(mai_mai_n410_), .B(mai_mai_n1118_), .Y(mai_mai_n1121_));
  NA3        m1093(.A(mai_mai_n416_), .B(mai_mai_n539_), .C(f), .Y(mai_mai_n1122_));
  NA2        m1094(.A(mai_mai_n39_), .B(mai_mai_n1109_), .Y(mai_mai_n1123_));
  NA3        m1095(.A(mai_mai_n1123_), .B(mai_mai_n1122_), .C(mai_mai_n1121_), .Y(mai_mai_n1124_));
  NA2        m1096(.A(i), .B(mai_mai_n117_), .Y(mai_mai_n1125_));
  OAI210     m1097(.A0(mai_mai_n1125_), .A1(mai_mai_n275_), .B0(g), .Y(mai_mai_n1126_));
  NAi21      m1098(.An(f), .B(d), .Y(mai_mai_n1127_));
  NO2        m1099(.A(mai_mai_n1127_), .B(mai_mai_n1085_), .Y(mai_mai_n1128_));
  INV        m1100(.A(mai_mai_n1128_), .Y(mai_mai_n1129_));
  AOI210     m1101(.A0(mai_mai_n1126_), .A1(mai_mai_n281_), .B0(mai_mai_n1129_), .Y(mai_mai_n1130_));
  AOI210     m1102(.A0(mai_mai_n1130_), .A1(mai_mai_n111_), .B0(mai_mai_n1124_), .Y(mai_mai_n1131_));
  NA2        m1103(.A(mai_mai_n455_), .B(mai_mai_n454_), .Y(mai_mai_n1132_));
  NO2        m1104(.A(mai_mai_n181_), .B(mai_mai_n237_), .Y(mai_mai_n1133_));
  NA2        m1105(.A(mai_mai_n1133_), .B(m), .Y(mai_mai_n1134_));
  INV        m1106(.A(mai_mai_n456_), .Y(mai_mai_n1135_));
  AOI210     m1107(.A0(mai_mai_n1135_), .A1(mai_mai_n1132_), .B0(mai_mai_n1134_), .Y(mai_mai_n1136_));
  NA2        m1108(.A(mai_mai_n541_), .B(mai_mai_n397_), .Y(mai_mai_n1137_));
  NO2        m1109(.A(mai_mai_n957_), .B(mai_mai_n214_), .Y(mai_mai_n1138_));
  NA2        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1128_), .Y(mai_mai_n1139_));
  NO2        m1111(.A(mai_mai_n363_), .B(mai_mai_n362_), .Y(mai_mai_n1140_));
  NA2        m1112(.A(mai_mai_n1133_), .B(mai_mai_n418_), .Y(mai_mai_n1141_));
  NA3        m1113(.A(mai_mai_n1141_), .B(mai_mai_n1139_), .C(mai_mai_n1137_), .Y(mai_mai_n1142_));
  NO2        m1114(.A(mai_mai_n1142_), .B(mai_mai_n1136_), .Y(mai_mai_n1143_));
  NA4        m1115(.A(mai_mai_n1143_), .B(mai_mai_n1131_), .C(mai_mai_n1120_), .D(mai_mai_n1116_), .Y(mai00));
  INV        m1116(.A(mai_mai_n287_), .Y(mai_mai_n1145_));
  NO2        m1117(.A(mai_mai_n1145_), .B(mai_mai_n560_), .Y(mai_mai_n1146_));
  AOI210     m1118(.A0(mai_mai_n892_), .A1(mai_mai_n937_), .B0(mai_mai_n1102_), .Y(mai_mai_n1147_));
  NO2        m1119(.A(mai_mai_n954_), .B(mai_mai_n701_), .Y(mai_mai_n1148_));
  NA3        m1120(.A(mai_mai_n1148_), .B(mai_mai_n1147_), .C(mai_mai_n996_), .Y(mai_mai_n1149_));
  NA2        m1121(.A(mai_mai_n492_), .B(f), .Y(mai_mai_n1150_));
  OAI210     m1122(.A0(mai_mai_n1003_), .A1(mai_mai_n40_), .B0(mai_mai_n633_), .Y(mai_mai_n1151_));
  NA3        m1123(.A(mai_mai_n1151_), .B(g), .C(n), .Y(mai_mai_n1152_));
  AOI210     m1124(.A0(mai_mai_n1152_), .A1(mai_mai_n1150_), .B0(mai_mai_n1038_), .Y(mai_mai_n1153_));
  NO4        m1125(.A(mai_mai_n1153_), .B(mai_mai_n1149_), .C(mai_mai_n1146_), .D(mai_mai_n1058_), .Y(mai_mai_n1154_));
  NA3        m1126(.A(mai_mai_n165_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1155_));
  NA2        m1127(.A(d), .B(b), .Y(mai_mai_n1156_));
  NOi31      m1128(.An(n), .B(m), .C(i), .Y(mai_mai_n1157_));
  NA3        m1129(.A(mai_mai_n1157_), .B(mai_mai_n636_), .C(mai_mai_n51_), .Y(mai_mai_n1158_));
  OAI210     m1130(.A0(mai_mai_n1156_), .A1(mai_mai_n1155_), .B0(mai_mai_n1158_), .Y(mai_mai_n1159_));
  INV        m1131(.A(mai_mai_n559_), .Y(mai_mai_n1160_));
  NO4        m1132(.A(mai_mai_n1160_), .B(mai_mai_n1159_), .C(mai_mai_n1140_), .D(mai_mai_n913_), .Y(mai_mai_n1161_));
  NO4        m1133(.A(mai_mai_n472_), .B(mai_mai_n346_), .C(mai_mai_n1117_), .D(mai_mai_n58_), .Y(mai_mai_n1162_));
  NA3        m1134(.A(mai_mai_n374_), .B(mai_mai_n221_), .C(g), .Y(mai_mai_n1163_));
  OR2        m1135(.A(mai_mai_n1163_), .B(mai_mai_n1156_), .Y(mai_mai_n1164_));
  NO2        m1136(.A(h), .B(g), .Y(mai_mai_n1165_));
  NA4        m1137(.A(mai_mai_n482_), .B(mai_mai_n452_), .C(mai_mai_n1165_), .D(mai_mai_n1030_), .Y(mai_mai_n1166_));
  OAI220     m1138(.A0(mai_mai_n507_), .A1(mai_mai_n582_), .B0(mai_mai_n89_), .B1(mai_mai_n88_), .Y(mai_mai_n1167_));
  AOI220     m1139(.A0(mai_mai_n1167_), .A1(mai_mai_n516_), .B0(mai_mai_n942_), .B1(mai_mai_n558_), .Y(mai_mai_n1168_));
  AOI220     m1140(.A0(mai_mai_n306_), .A1(mai_mai_n246_), .B0(mai_mai_n176_), .B1(mai_mai_n147_), .Y(mai_mai_n1169_));
  NA4        m1141(.A(mai_mai_n1169_), .B(mai_mai_n1168_), .C(mai_mai_n1166_), .D(mai_mai_n1164_), .Y(mai_mai_n1170_));
  NO2        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1162_), .Y(mai_mai_n1171_));
  AOI210     m1143(.A0(mai_mai_n246_), .A1(mai_mai_n336_), .B0(mai_mai_n561_), .Y(mai_mai_n1172_));
  NA2        m1144(.A(mai_mai_n1172_), .B(mai_mai_n153_), .Y(mai_mai_n1173_));
  NO2        m1145(.A(mai_mai_n239_), .B(mai_mai_n180_), .Y(mai_mai_n1174_));
  NA2        m1146(.A(mai_mai_n1174_), .B(mai_mai_n416_), .Y(mai_mai_n1175_));
  NA3        m1147(.A(mai_mai_n178_), .B(mai_mai_n110_), .C(g), .Y(mai_mai_n1176_));
  NA3        m1148(.A(mai_mai_n452_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1177_));
  NOi31      m1149(.An(mai_mai_n867_), .B(mai_mai_n1177_), .C(mai_mai_n1176_), .Y(mai_mai_n1178_));
  NAi31      m1150(.An(mai_mai_n184_), .B(mai_mai_n855_), .C(mai_mai_n452_), .Y(mai_mai_n1179_));
  NAi31      m1151(.An(mai_mai_n1178_), .B(mai_mai_n1179_), .C(mai_mai_n1175_), .Y(mai_mai_n1180_));
  NO2        m1152(.A(mai_mai_n267_), .B(mai_mai_n70_), .Y(mai_mai_n1181_));
  NO3        m1153(.A(mai_mai_n415_), .B(mai_mai_n828_), .C(n), .Y(mai_mai_n1182_));
  AOI210     m1154(.A0(mai_mai_n1182_), .A1(mai_mai_n1181_), .B0(mai_mai_n1071_), .Y(mai_mai_n1183_));
  NAi21      m1155(.An(mai_mai_n1041_), .B(mai_mai_n1183_), .Y(mai_mai_n1184_));
  NO3        m1156(.A(mai_mai_n1184_), .B(mai_mai_n1180_), .C(mai_mai_n1173_), .Y(mai_mai_n1185_));
  AN3        m1157(.A(mai_mai_n1185_), .B(mai_mai_n1171_), .C(mai_mai_n1161_), .Y(mai_mai_n1186_));
  NA2        m1158(.A(mai_mai_n516_), .B(mai_mai_n99_), .Y(mai_mai_n1187_));
  NA3        m1159(.A(mai_mai_n1103_), .B(mai_mai_n593_), .C(mai_mai_n451_), .Y(mai_mai_n1188_));
  NA4        m1160(.A(mai_mai_n1188_), .B(mai_mai_n542_), .C(mai_mai_n1187_), .D(mai_mai_n241_), .Y(mai_mai_n1189_));
  NA2        m1161(.A(mai_mai_n1097_), .B(mai_mai_n516_), .Y(mai_mai_n1190_));
  NA4        m1162(.A(mai_mai_n636_), .B(mai_mai_n205_), .C(mai_mai_n221_), .D(mai_mai_n162_), .Y(mai_mai_n1191_));
  NA2        m1163(.A(mai_mai_n1190_), .B(mai_mai_n284_), .Y(mai_mai_n1192_));
  OAI210     m1164(.A0(mai_mai_n450_), .A1(mai_mai_n118_), .B0(mai_mai_n861_), .Y(mai_mai_n1193_));
  AOI210     m1165(.A0(mai_mai_n541_), .A1(mai_mai_n397_), .B0(mai_mai_n1193_), .Y(mai_mai_n1194_));
  OR3        m1166(.A(mai_mai_n1038_), .B(mai_mai_n263_), .C(mai_mai_n223_), .Y(mai_mai_n1195_));
  NO2        m1167(.A(mai_mai_n217_), .B(mai_mai_n214_), .Y(mai_mai_n1196_));
  NA2        m1168(.A(n), .B(e), .Y(mai_mai_n1197_));
  NO2        m1169(.A(mai_mai_n1197_), .B(mai_mai_n145_), .Y(mai_mai_n1198_));
  AOI220     m1170(.A0(mai_mai_n1198_), .A1(mai_mai_n265_), .B0(mai_mai_n843_), .B1(mai_mai_n1196_), .Y(mai_mai_n1199_));
  NA2        m1171(.A(mai_mai_n347_), .B(mai_mai_n436_), .Y(mai_mai_n1200_));
  NA4        m1172(.A(mai_mai_n1200_), .B(mai_mai_n1199_), .C(mai_mai_n1195_), .D(mai_mai_n1194_), .Y(mai_mai_n1201_));
  AOI210     m1173(.A0(mai_mai_n1198_), .A1(mai_mai_n846_), .B0(mai_mai_n816_), .Y(mai_mai_n1202_));
  AOI220     m1174(.A0(mai_mai_n950_), .A1(mai_mai_n558_), .B0(mai_mai_n636_), .B1(mai_mai_n244_), .Y(mai_mai_n1203_));
  NO2        m1175(.A(mai_mai_n65_), .B(h), .Y(mai_mai_n1204_));
  NO3        m1176(.A(mai_mai_n1038_), .B(mai_mai_n1036_), .C(mai_mai_n718_), .Y(mai_mai_n1205_));
  OAI210     m1177(.A0(mai_mai_n1083_), .A1(mai_mai_n1205_), .B0(mai_mai_n1204_), .Y(mai_mai_n1206_));
  NA4        m1178(.A(mai_mai_n1206_), .B(mai_mai_n1203_), .C(mai_mai_n1202_), .D(mai_mai_n863_), .Y(mai_mai_n1207_));
  NO4        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1201_), .C(mai_mai_n1192_), .D(mai_mai_n1189_), .Y(mai_mai_n1208_));
  NA2        m1180(.A(mai_mai_n833_), .B(mai_mai_n748_), .Y(mai_mai_n1209_));
  NA4        m1181(.A(mai_mai_n1209_), .B(mai_mai_n1208_), .C(mai_mai_n1186_), .D(mai_mai_n1154_), .Y(mai01));
  NO3        m1182(.A(mai_mai_n796_), .B(mai_mai_n788_), .C(mai_mai_n463_), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n575_), .B(mai_mai_n278_), .Y(mai_mai_n1212_));
  OAI210     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n381_), .B0(i), .Y(mai_mai_n1213_));
  NA3        m1185(.A(mai_mai_n1213_), .B(mai_mai_n1211_), .C(mai_mai_n1018_), .Y(mai_mai_n1214_));
  NA2        m1186(.A(mai_mai_n571_), .B(mai_mai_n87_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n956_), .B(c), .Y(mai_mai_n1216_));
  NA4        m1188(.A(mai_mai_n1216_), .B(mai_mai_n1215_), .C(mai_mai_n906_), .D(mai_mai_n321_), .Y(mai_mai_n1217_));
  NA2        m1189(.A(mai_mai_n696_), .B(mai_mai_n94_), .Y(mai_mai_n1218_));
  NO2        m1190(.A(mai_mai_n1218_), .B(i), .Y(mai_mai_n1219_));
  OAI210     m1191(.A0(mai_mai_n775_), .A1(mai_mai_n588_), .B0(mai_mai_n1191_), .Y(mai_mai_n1220_));
  AOI210     m1192(.A0(mai_mai_n1219_), .A1(mai_mai_n623_), .B0(mai_mai_n1220_), .Y(mai_mai_n1221_));
  NA2        m1193(.A(mai_mai_n116_), .B(l), .Y(mai_mai_n1222_));
  OA220      m1194(.A0(mai_mai_n1222_), .A1(mai_mai_n568_), .B0(mai_mai_n648_), .B1(mai_mai_n360_), .Y(mai_mai_n1223_));
  NAi41      m1195(.An(mai_mai_n161_), .B(mai_mai_n1223_), .C(mai_mai_n1221_), .D(mai_mai_n891_), .Y(mai_mai_n1224_));
  NO3        m1196(.A(mai_mai_n776_), .B(mai_mai_n661_), .C(mai_mai_n494_), .Y(mai_mai_n1225_));
  NA4        m1197(.A(mai_mai_n696_), .B(mai_mai_n94_), .C(mai_mai_n45_), .D(mai_mai_n213_), .Y(mai_mai_n1226_));
  OR2        m1198(.A(mai_mai_n194_), .B(mai_mai_n192_), .Y(mai_mai_n1227_));
  NA3        m1199(.A(mai_mai_n1227_), .B(mai_mai_n1225_), .C(mai_mai_n136_), .Y(mai_mai_n1228_));
  NO4        m1200(.A(mai_mai_n1228_), .B(mai_mai_n1224_), .C(mai_mai_n1217_), .D(mai_mai_n1214_), .Y(mai_mai_n1229_));
  NA2        m1201(.A(mai_mai_n519_), .B(mai_mai_n383_), .Y(mai_mai_n1230_));
  AOI210     m1202(.A0(mai_mai_n574_), .A1(mai_mai_n568_), .B0(mai_mai_n1433_), .Y(mai_mai_n1231_));
  AOI210     m1203(.A0(mai_mai_n543_), .A1(mai_mai_n1230_), .B0(mai_mai_n1231_), .Y(mai_mai_n1232_));
  AOI210     m1204(.A0(mai_mai_n203_), .A1(mai_mai_n86_), .B0(mai_mai_n213_), .Y(mai_mai_n1233_));
  OAI210     m1205(.A0(mai_mai_n803_), .A1(mai_mai_n416_), .B0(mai_mai_n1233_), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n1234_), .B(mai_mai_n1232_), .Y(mai_mai_n1235_));
  AOI210     m1207(.A0(mai_mai_n580_), .A1(mai_mai_n116_), .B0(mai_mai_n586_), .Y(mai_mai_n1236_));
  OAI210     m1208(.A0(mai_mai_n1222_), .A1(mai_mai_n577_), .B0(mai_mai_n1236_), .Y(mai_mai_n1237_));
  NO2        m1209(.A(mai_mai_n815_), .B(mai_mai_n203_), .Y(mai_mai_n1238_));
  NO2        m1210(.A(mai_mai_n1238_), .B(mai_mai_n954_), .Y(mai_mai_n1239_));
  OAI210     m1211(.A0(mai_mai_n1219_), .A1(mai_mai_n314_), .B0(mai_mai_n662_), .Y(mai_mai_n1240_));
  NA3        m1212(.A(mai_mai_n1240_), .B(mai_mai_n1239_), .C(mai_mai_n779_), .Y(mai_mai_n1241_));
  NO3        m1213(.A(mai_mai_n1241_), .B(mai_mai_n1237_), .C(mai_mai_n1235_), .Y(mai_mai_n1242_));
  NA3        m1214(.A(mai_mai_n589_), .B(mai_mai_n29_), .C(f), .Y(mai_mai_n1243_));
  NO2        m1215(.A(mai_mai_n1243_), .B(mai_mai_n203_), .Y(mai_mai_n1244_));
  AOI210     m1216(.A0(mai_mai_n488_), .A1(mai_mai_n57_), .B0(mai_mai_n1244_), .Y(mai_mai_n1245_));
  OR2        m1217(.A(mai_mai_n1218_), .B(mai_mai_n590_), .Y(mai_mai_n1246_));
  NA3        m1218(.A(mai_mai_n730_), .B(mai_mai_n71_), .C(i), .Y(mai_mai_n1247_));
  AOI210     m1219(.A0(mai_mai_n1247_), .A1(mai_mai_n1226_), .B0(mai_mai_n973_), .Y(mai_mai_n1248_));
  NO2        m1220(.A(mai_mai_n1248_), .B(mai_mai_n1159_), .Y(mai_mai_n1249_));
  NA4        m1221(.A(mai_mai_n1249_), .B(mai_mai_n1246_), .C(mai_mai_n1245_), .D(mai_mai_n747_), .Y(mai_mai_n1250_));
  NO2        m1222(.A(mai_mai_n961_), .B(mai_mai_n232_), .Y(mai_mai_n1251_));
  NO2        m1223(.A(mai_mai_n962_), .B(mai_mai_n536_), .Y(mai_mai_n1252_));
  OAI210     m1224(.A0(mai_mai_n1252_), .A1(mai_mai_n1251_), .B0(mai_mai_n329_), .Y(mai_mai_n1253_));
  NA2        m1225(.A(mai_mai_n553_), .B(mai_mai_n551_), .Y(mai_mai_n1254_));
  NO3        m1226(.A(mai_mai_n76_), .B(mai_mai_n288_), .C(mai_mai_n45_), .Y(mai_mai_n1255_));
  NA2        m1227(.A(mai_mai_n1255_), .B(mai_mai_n533_), .Y(mai_mai_n1256_));
  NA3        m1228(.A(mai_mai_n1256_), .B(mai_mai_n1254_), .C(mai_mai_n657_), .Y(mai_mai_n1257_));
  OR2        m1229(.A(mai_mai_n1163_), .B(mai_mai_n1156_), .Y(mai_mai_n1258_));
  NO2        m1230(.A(mai_mai_n360_), .B(mai_mai_n69_), .Y(mai_mai_n1259_));
  AOI210     m1231(.A0(mai_mai_n723_), .A1(mai_mai_n604_), .B0(mai_mai_n1259_), .Y(mai_mai_n1260_));
  NA2        m1232(.A(mai_mai_n1255_), .B(mai_mai_n806_), .Y(mai_mai_n1261_));
  NA4        m1233(.A(mai_mai_n1261_), .B(mai_mai_n1260_), .C(mai_mai_n1258_), .D(mai_mai_n376_), .Y(mai_mai_n1262_));
  NOi41      m1234(.An(mai_mai_n1253_), .B(mai_mai_n1262_), .C(mai_mai_n1257_), .D(mai_mai_n1250_), .Y(mai_mai_n1263_));
  NO2        m1235(.A(mai_mai_n129_), .B(mai_mai_n45_), .Y(mai_mai_n1264_));
  NO2        m1236(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1265_));
  AO220      m1237(.A0(mai_mai_n1265_), .A1(mai_mai_n609_), .B0(mai_mai_n1264_), .B1(mai_mai_n694_), .Y(mai_mai_n1266_));
  NA2        m1238(.A(mai_mai_n1266_), .B(mai_mai_n329_), .Y(mai_mai_n1267_));
  INV        m1239(.A(mai_mai_n133_), .Y(mai_mai_n1268_));
  NO3        m1240(.A(mai_mai_n1081_), .B(mai_mai_n175_), .C(mai_mai_n84_), .Y(mai_mai_n1269_));
  AOI220     m1241(.A0(mai_mai_n1269_), .A1(mai_mai_n1268_), .B0(mai_mai_n1255_), .B1(mai_mai_n965_), .Y(mai_mai_n1270_));
  NA2        m1242(.A(mai_mai_n1270_), .B(mai_mai_n1267_), .Y(mai_mai_n1271_));
  NO2        m1243(.A(mai_mai_n601_), .B(mai_mai_n600_), .Y(mai_mai_n1272_));
  NO4        m1244(.A(mai_mai_n1081_), .B(mai_mai_n1272_), .C(mai_mai_n173_), .D(mai_mai_n84_), .Y(mai_mai_n1273_));
  NO3        m1245(.A(mai_mai_n1273_), .B(mai_mai_n1271_), .C(mai_mai_n627_), .Y(mai_mai_n1274_));
  NA4        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1263_), .C(mai_mai_n1242_), .D(mai_mai_n1229_), .Y(mai06));
  NA2        m1247(.A(mai_mai_n1269_), .B(mai_mai_n373_), .Y(mai_mai_n1276_));
  NO3        m1248(.A(mai_mai_n584_), .B(mai_mai_n801_), .C(mai_mai_n587_), .Y(mai_mai_n1277_));
  OR2        m1249(.A(mai_mai_n1277_), .B(mai_mai_n882_), .Y(mai_mai_n1278_));
  NA3        m1250(.A(mai_mai_n1278_), .B(mai_mai_n1276_), .C(mai_mai_n1253_), .Y(mai_mai_n1279_));
  NO3        m1251(.A(mai_mai_n1279_), .B(mai_mai_n1257_), .C(mai_mai_n254_), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n288_), .B(mai_mai_n45_), .Y(mai_mai_n1281_));
  AOI210     m1253(.A0(mai_mai_n1281_), .A1(mai_mai_n966_), .B0(mai_mai_n1251_), .Y(mai_mai_n1282_));
  AOI210     m1254(.A0(mai_mai_n1281_), .A1(mai_mai_n537_), .B0(mai_mai_n1266_), .Y(mai_mai_n1283_));
  AOI210     m1255(.A0(mai_mai_n1283_), .A1(mai_mai_n1282_), .B0(mai_mai_n326_), .Y(mai_mai_n1284_));
  OAI210     m1256(.A0(mai_mai_n86_), .A1(mai_mai_n40_), .B0(mai_mai_n660_), .Y(mai_mai_n1285_));
  NA2        m1257(.A(mai_mai_n1285_), .B(mai_mai_n630_), .Y(mai_mai_n1286_));
  NO2        m1258(.A(mai_mai_n594_), .B(mai_mai_n1104_), .Y(mai_mai_n1287_));
  INV        m1259(.A(mai_mai_n900_), .Y(mai_mai_n1288_));
  NO3        m1260(.A(mai_mai_n1288_), .B(mai_mai_n1287_), .C(mai_mai_n135_), .Y(mai_mai_n1289_));
  OR2        m1261(.A(mai_mai_n585_), .B(mai_mai_n583_), .Y(mai_mai_n1290_));
  INV        m1262(.A(mai_mai_n1290_), .Y(mai_mai_n1291_));
  NA3        m1263(.A(mai_mai_n1291_), .B(mai_mai_n1289_), .C(mai_mai_n1286_), .Y(mai_mai_n1292_));
  AN2        m1264(.A(mai_mai_n950_), .B(c), .Y(mai_mai_n1293_));
  NO3        m1265(.A(mai_mai_n1293_), .B(mai_mai_n1292_), .C(mai_mai_n1284_), .Y(mai_mai_n1294_));
  NO2        m1266(.A(mai_mai_n225_), .B(mai_mai_n603_), .Y(mai_mai_n1295_));
  NA2        m1267(.A(mai_mai_n1432_), .B(mai_mai_n1295_), .Y(mai_mai_n1296_));
  NO3        m1268(.A(mai_mai_n243_), .B(mai_mai_n101_), .C(mai_mai_n272_), .Y(mai_mai_n1297_));
  OAI220     m1269(.A0(mai_mai_n686_), .A1(mai_mai_n247_), .B0(mai_mai_n493_), .B1(mai_mai_n497_), .Y(mai_mai_n1298_));
  NO2        m1270(.A(mai_mai_n582_), .B(j), .Y(mai_mai_n1299_));
  NO3        m1271(.A(mai_mai_n1298_), .B(mai_mai_n1297_), .C(mai_mai_n1106_), .Y(mai_mai_n1300_));
  NA4        m1272(.A(mai_mai_n786_), .B(mai_mai_n785_), .C(mai_mai_n426_), .D(mai_mai_n874_), .Y(mai_mai_n1301_));
  NAi31      m1273(.An(mai_mai_n738_), .B(mai_mai_n1301_), .C(mai_mai_n202_), .Y(mai_mai_n1302_));
  NA4        m1274(.A(mai_mai_n1302_), .B(mai_mai_n1300_), .C(mai_mai_n1296_), .D(mai_mai_n1203_), .Y(mai_mai_n1303_));
  NOi31      m1275(.An(mai_mai_n1277_), .B(mai_mai_n449_), .C(mai_mai_n382_), .Y(mai_mai_n1304_));
  OR3        m1276(.A(mai_mai_n1304_), .B(mai_mai_n775_), .C(mai_mai_n522_), .Y(mai_mai_n1305_));
  NA2        m1277(.A(mai_mai_n553_), .B(mai_mai_n436_), .Y(mai_mai_n1306_));
  NA2        m1278(.A(mai_mai_n1299_), .B(mai_mai_n782_), .Y(mai_mai_n1307_));
  NA3        m1279(.A(mai_mai_n1307_), .B(mai_mai_n1306_), .C(mai_mai_n1305_), .Y(mai_mai_n1308_));
  AN2        m1280(.A(mai_mai_n922_), .B(mai_mai_n921_), .Y(mai_mai_n1309_));
  NO4        m1281(.A(mai_mai_n1309_), .B(mai_mai_n872_), .C(mai_mai_n484_), .D(mai_mai_n466_), .Y(mai_mai_n1310_));
  NA2        m1282(.A(mai_mai_n1310_), .B(mai_mai_n1261_), .Y(mai_mai_n1311_));
  NAi21      m1283(.An(j), .B(i), .Y(mai_mai_n1312_));
  NO4        m1284(.A(mai_mai_n1272_), .B(mai_mai_n1312_), .C(mai_mai_n432_), .D(mai_mai_n235_), .Y(mai_mai_n1313_));
  NO4        m1285(.A(mai_mai_n1313_), .B(mai_mai_n1311_), .C(mai_mai_n1308_), .D(mai_mai_n1303_), .Y(mai_mai_n1314_));
  NA4        m1286(.A(mai_mai_n1314_), .B(mai_mai_n1294_), .C(mai_mai_n1280_), .D(mai_mai_n1274_), .Y(mai07));
  NAi32      m1287(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1316_));
  NO3        m1288(.A(mai_mai_n1316_), .B(g), .C(f), .Y(mai_mai_n1317_));
  OAI210     m1289(.A0(i), .A1(mai_mai_n468_), .B0(mai_mai_n1317_), .Y(mai_mai_n1318_));
  NAi21      m1290(.An(f), .B(c), .Y(mai_mai_n1319_));
  OR2        m1291(.A(e), .B(d), .Y(mai_mai_n1320_));
  OAI220     m1292(.A0(mai_mai_n1320_), .A1(mai_mai_n1319_), .B0(mai_mai_n615_), .B1(mai_mai_n310_), .Y(mai_mai_n1321_));
  NA3        m1293(.A(mai_mai_n1321_), .B(mai_mai_n1429_), .C(mai_mai_n178_), .Y(mai_mai_n1322_));
  NOi31      m1294(.An(n), .B(m), .C(b), .Y(mai_mai_n1323_));
  NO3        m1295(.A(mai_mai_n130_), .B(mai_mai_n437_), .C(h), .Y(mai_mai_n1324_));
  NA2        m1296(.A(mai_mai_n1322_), .B(mai_mai_n1318_), .Y(mai_mai_n1325_));
  NOi41      m1297(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1326_));
  NO2        m1298(.A(mai_mai_n1055_), .B(mai_mai_n295_), .Y(mai_mai_n1327_));
  NA2        m1299(.A(mai_mai_n523_), .B(mai_mai_n77_), .Y(mai_mai_n1328_));
  NA2        m1300(.A(mai_mai_n1204_), .B(mai_mai_n279_), .Y(mai_mai_n1329_));
  NA2        m1301(.A(mai_mai_n1329_), .B(mai_mai_n1328_), .Y(mai_mai_n1330_));
  NO2        m1302(.A(mai_mai_n1330_), .B(mai_mai_n1325_), .Y(mai_mai_n1331_));
  NO3        m1303(.A(e), .B(d), .C(c), .Y(mai_mai_n1332_));
  OAI210     m1304(.A0(mai_mai_n130_), .A1(mai_mai_n214_), .B0(mai_mai_n591_), .Y(mai_mai_n1333_));
  NA2        m1305(.A(mai_mai_n1333_), .B(mai_mai_n1332_), .Y(mai_mai_n1334_));
  INV        m1306(.A(mai_mai_n1334_), .Y(mai_mai_n1335_));
  NA3        m1307(.A(mai_mai_n683_), .B(mai_mai_n670_), .C(mai_mai_n110_), .Y(mai_mai_n1336_));
  NO2        m1308(.A(mai_mai_n1336_), .B(mai_mai_n45_), .Y(mai_mai_n1337_));
  NO2        m1309(.A(l), .B(k), .Y(mai_mai_n1338_));
  NO3        m1310(.A(mai_mai_n432_), .B(d), .C(c), .Y(mai_mai_n1339_));
  NO2        m1311(.A(mai_mai_n1337_), .B(mai_mai_n1335_), .Y(mai_mai_n1340_));
  NO2        m1312(.A(mai_mai_n146_), .B(h), .Y(mai_mai_n1341_));
  NO2        m1313(.A(g), .B(c), .Y(mai_mai_n1342_));
  NA3        m1314(.A(mai_mai_n1342_), .B(mai_mai_n141_), .C(mai_mai_n185_), .Y(mai_mai_n1343_));
  NO2        m1315(.A(mai_mai_n1343_), .B(mai_mai_n1428_), .Y(mai_mai_n1344_));
  NA2        m1316(.A(mai_mai_n1344_), .B(mai_mai_n178_), .Y(mai_mai_n1345_));
  NO2        m1317(.A(i), .B(h), .Y(mai_mai_n1346_));
  AOI210     m1318(.A0(mai_mai_n1127_), .A1(h), .B0(mai_mai_n403_), .Y(mai_mai_n1347_));
  NA2        m1319(.A(mai_mai_n137_), .B(mai_mai_n221_), .Y(mai_mai_n1348_));
  NO2        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1347_), .Y(mai_mai_n1349_));
  NO2        m1321(.A(mai_mai_n745_), .B(mai_mai_n186_), .Y(mai_mai_n1350_));
  NOi31      m1322(.An(m), .B(n), .C(b), .Y(mai_mai_n1351_));
  NOi31      m1323(.An(f), .B(d), .C(c), .Y(mai_mai_n1352_));
  NA2        m1324(.A(mai_mai_n1352_), .B(mai_mai_n1351_), .Y(mai_mai_n1353_));
  INV        m1325(.A(mai_mai_n1353_), .Y(mai_mai_n1354_));
  NO3        m1326(.A(mai_mai_n1354_), .B(mai_mai_n1350_), .C(mai_mai_n1349_), .Y(mai_mai_n1355_));
  NA2        m1327(.A(mai_mai_n1074_), .B(mai_mai_n452_), .Y(mai_mai_n1356_));
  OAI210     m1328(.A0(mai_mai_n181_), .A1(mai_mai_n506_), .B0(mai_mai_n1051_), .Y(mai_mai_n1357_));
  NO3        m1329(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1358_));
  AN3        m1330(.A(mai_mai_n1357_), .B(mai_mai_n1355_), .C(mai_mai_n1345_), .Y(mai_mai_n1359_));
  NA2        m1331(.A(mai_mai_n1339_), .B(mai_mai_n215_), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n1082_), .B(mai_mai_n1356_), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n1361_), .B(mai_mai_n1360_), .Y(mai_mai_n1362_));
  NO4        m1334(.A(mai_mai_n130_), .B(g), .C(f), .D(e), .Y(mai_mai_n1363_));
  NA2        m1335(.A(mai_mai_n280_), .B(h), .Y(mai_mai_n1364_));
  OR2        m1336(.A(e), .B(a), .Y(mai_mai_n1365_));
  NA2        m1337(.A(mai_mai_n30_), .B(h), .Y(mai_mai_n1366_));
  NO2        m1338(.A(mai_mai_n1366_), .B(mai_mai_n1070_), .Y(mai_mai_n1367_));
  NA2        m1339(.A(mai_mai_n1326_), .B(mai_mai_n1338_), .Y(mai_mai_n1368_));
  OR3        m1340(.A(mai_mai_n522_), .B(mai_mai_n521_), .C(mai_mai_n110_), .Y(mai_mai_n1369_));
  NO3        m1341(.A(mai_mai_n1431_), .B(mai_mai_n1367_), .C(mai_mai_n1362_), .Y(mai_mai_n1370_));
  NA4        m1342(.A(mai_mai_n1370_), .B(mai_mai_n1359_), .C(mai_mai_n1340_), .D(mai_mai_n1331_), .Y(mai_mai_n1371_));
  NA3        m1343(.A(mai_mai_n1358_), .B(mai_mai_n1320_), .C(mai_mai_n1103_), .Y(mai_mai_n1372_));
  NAi41      m1344(.An(mai_mai_n1346_), .B(mai_mai_n1063_), .C(mai_mai_n166_), .D(mai_mai_n149_), .Y(mai_mai_n1373_));
  NA2        m1345(.A(mai_mai_n1373_), .B(mai_mai_n1372_), .Y(mai_mai_n1374_));
  NO3        m1346(.A(mai_mai_n738_), .B(mai_mai_n173_), .C(mai_mai_n398_), .Y(mai_mai_n1375_));
  NO2        m1347(.A(mai_mai_n1375_), .B(mai_mai_n1374_), .Y(mai_mai_n1376_));
  OR2        m1348(.A(n), .B(i), .Y(mai_mai_n1377_));
  OAI210     m1349(.A0(mai_mai_n1377_), .A1(mai_mai_n1062_), .B0(mai_mai_n49_), .Y(mai_mai_n1378_));
  AOI220     m1350(.A0(mai_mai_n1378_), .A1(mai_mai_n1165_), .B0(mai_mai_n820_), .B1(mai_mai_n193_), .Y(mai_mai_n1379_));
  NO3        m1351(.A(mai_mai_n1085_), .B(mai_mai_n1320_), .C(mai_mai_n49_), .Y(mai_mai_n1380_));
  NA2        m1352(.A(mai_mai_n178_), .B(mai_mai_n110_), .Y(mai_mai_n1381_));
  NOi21      m1353(.An(d), .B(f), .Y(mai_mai_n1382_));
  NO2        m1354(.A(mai_mai_n1320_), .B(f), .Y(mai_mai_n1383_));
  NA2        m1355(.A(mai_mai_n1379_), .B(mai_mai_n1376_), .Y(mai_mai_n1384_));
  NO3        m1356(.A(mai_mai_n1074_), .B(mai_mai_n1062_), .C(mai_mai_n40_), .Y(mai_mai_n1385_));
  NA2        m1357(.A(mai_mai_n1385_), .B(mai_mai_n1327_), .Y(mai_mai_n1386_));
  OAI210     m1358(.A0(mai_mai_n1363_), .A1(mai_mai_n1323_), .B0(mai_mai_n879_), .Y(mai_mai_n1387_));
  NA2        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1386_), .Y(mai_mai_n1388_));
  NA2        m1360(.A(mai_mai_n1342_), .B(mai_mai_n1382_), .Y(mai_mai_n1389_));
  NO2        m1361(.A(mai_mai_n1389_), .B(m), .Y(mai_mai_n1390_));
  NA2        m1362(.A(mai_mai_n108_), .B(mai_mai_n1351_), .Y(mai_mai_n1391_));
  INV        m1363(.A(mai_mai_n1391_), .Y(mai_mai_n1392_));
  NO3        m1364(.A(mai_mai_n1392_), .B(mai_mai_n1390_), .C(mai_mai_n1388_), .Y(mai_mai_n1393_));
  NO2        m1365(.A(mai_mai_n1319_), .B(e), .Y(mai_mai_n1394_));
  NA2        m1366(.A(mai_mai_n1112_), .B(mai_mai_n619_), .Y(mai_mai_n1395_));
  NO2        m1367(.A(mai_mai_n1395_), .B(mai_mai_n434_), .Y(mai_mai_n1396_));
  NO3        m1368(.A(mai_mai_n1369_), .B(mai_mai_n343_), .C(a), .Y(mai_mai_n1397_));
  NO2        m1369(.A(mai_mai_n1397_), .B(mai_mai_n1396_), .Y(mai_mai_n1398_));
  NO2        m1370(.A(mai_mai_n180_), .B(c), .Y(mai_mai_n1399_));
  OAI210     m1371(.A0(mai_mai_n1399_), .A1(mai_mai_n1394_), .B0(mai_mai_n178_), .Y(mai_mai_n1400_));
  AOI220     m1372(.A0(mai_mai_n1400_), .A1(mai_mai_n1064_), .B0(mai_mai_n513_), .B1(mai_mai_n358_), .Y(mai_mai_n1401_));
  AOI210     m1373(.A0(mai_mai_n895_), .A1(mai_mai_n405_), .B0(mai_mai_n103_), .Y(mai_mai_n1402_));
  OR2        m1374(.A(mai_mai_n1402_), .B(mai_mai_n521_), .Y(mai_mai_n1403_));
  NO2        m1375(.A(mai_mai_n1403_), .B(mai_mai_n173_), .Y(mai_mai_n1404_));
  NA2        m1376(.A(mai_mai_n1324_), .B(mai_mai_n181_), .Y(mai_mai_n1405_));
  NO2        m1377(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1406_));
  OAI210     m1378(.A0(mai_mai_n1365_), .A1(mai_mai_n857_), .B0(mai_mai_n468_), .Y(mai_mai_n1407_));
  OAI210     m1379(.A0(mai_mai_n1407_), .A1(mai_mai_n1086_), .B0(mai_mai_n1406_), .Y(mai_mai_n1408_));
  NO2        m1380(.A(m), .B(i), .Y(mai_mai_n1409_));
  NA2        m1381(.A(mai_mai_n1409_), .B(mai_mai_n1341_), .Y(mai_mai_n1410_));
  NA3        m1382(.A(mai_mai_n1410_), .B(mai_mai_n1408_), .C(mai_mai_n1405_), .Y(mai_mai_n1411_));
  NO4        m1383(.A(mai_mai_n1411_), .B(mai_mai_n1404_), .C(mai_mai_n1380_), .D(mai_mai_n1401_), .Y(mai_mai_n1412_));
  NA3        m1384(.A(mai_mai_n1412_), .B(mai_mai_n1398_), .C(mai_mai_n1393_), .Y(mai_mai_n1413_));
  AOI210     m1385(.A0(mai_mai_n156_), .A1(mai_mai_n55_), .B0(mai_mai_n1394_), .Y(mai_mai_n1414_));
  NO2        m1386(.A(mai_mai_n1414_), .B(mai_mai_n1381_), .Y(mai_mai_n1415_));
  OR4        m1387(.A(mai_mai_n1415_), .B(mai_mai_n1413_), .C(mai_mai_n1384_), .D(mai_mai_n1371_), .Y(mai04));
  NOi31      m1388(.An(mai_mai_n1363_), .B(mai_mai_n1364_), .C(mai_mai_n1038_), .Y(mai_mai_n1417_));
  NA2        m1389(.A(mai_mai_n1383_), .B(mai_mai_n820_), .Y(mai_mai_n1418_));
  NO2        m1390(.A(mai_mai_n1418_), .B(mai_mai_n1031_), .Y(mai_mai_n1419_));
  OR3        m1391(.A(mai_mai_n1419_), .B(mai_mai_n1417_), .C(mai_mai_n1053_), .Y(mai_mai_n1420_));
  NO2        m1392(.A(mai_mai_n88_), .B(k), .Y(mai_mai_n1421_));
  AOI210     m1393(.A0(mai_mai_n1421_), .A1(mai_mai_n1048_), .B0(mai_mai_n1178_), .Y(mai_mai_n1422_));
  NA2        m1394(.A(mai_mai_n1422_), .B(mai_mai_n1206_), .Y(mai_mai_n1423_));
  NO4        m1395(.A(mai_mai_n1423_), .B(mai_mai_n1420_), .C(mai_mai_n1061_), .D(mai_mai_n1043_), .Y(mai_mai_n1424_));
  NA4        m1396(.A(mai_mai_n1424_), .B(mai_mai_n1114_), .C(mai_mai_n1101_), .D(mai_mai_n1089_), .Y(mai05));
  INV        m1397(.A(l), .Y(mai_mai_n1428_));
  INV        m1398(.A(j), .Y(mai_mai_n1429_));
  INV        m1399(.A(g), .Y(mai_mai_n1430_));
  INV        m1400(.A(mai_mai_n1368_), .Y(mai_mai_n1431_));
  INV        m1401(.A(mai_mai_n268_), .Y(mai_mai_n1432_));
  INV        m1402(.A(k), .Y(mai_mai_n1433_));
  INV        m1403(.A(k), .Y(mai_mai_n1434_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  NO2        u0023(.A(men_men_n51_), .B(men_men_n50_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NAi31      u0033(.An(i), .B(l), .C(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(g), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(g), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(g), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n103_), .B(f), .Y(men_men_n104_));
  NO4        u0076(.A(men_men_n104_), .B(men_men_n98_), .C(men_men_n95_), .D(men_men_n92_), .Y(men_men_n105_));
  NAi41      u0077(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n106_));
  AN2        u0078(.A(e), .B(b), .Y(men_men_n107_));
  NOi31      u0079(.An(c), .B(h), .C(f), .Y(men_men_n108_));
  NA2        u0080(.A(men_men_n108_), .B(men_men_n107_), .Y(men_men_n109_));
  NO3        u0081(.A(men_men_n109_), .B(men_men_n106_), .C(g), .Y(men_men_n110_));
  NOi21      u0082(.An(g), .B(f), .Y(men_men_n111_));
  NOi21      u0083(.An(i), .B(h), .Y(men_men_n112_));
  NA3        u0084(.A(men_men_n112_), .B(men_men_n111_), .C(men_men_n36_), .Y(men_men_n113_));
  INV        u0085(.A(a), .Y(men_men_n114_));
  NA2        u0086(.A(men_men_n107_), .B(men_men_n114_), .Y(men_men_n115_));
  INV        u0087(.A(l), .Y(men_men_n116_));
  NOi21      u0088(.An(m), .B(n), .Y(men_men_n117_));
  AN2        u0089(.A(k), .B(h), .Y(men_men_n118_));
  NO2        u0090(.A(men_men_n113_), .B(men_men_n88_), .Y(men_men_n119_));
  INV        u0091(.A(b), .Y(men_men_n120_));
  NA2        u0092(.A(l), .B(j), .Y(men_men_n121_));
  AN2        u0093(.A(k), .B(i), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n121_), .Y(men_men_n123_));
  NA2        u0095(.A(g), .B(e), .Y(men_men_n124_));
  NOi32      u0096(.An(c), .Bn(a), .C(d), .Y(men_men_n125_));
  NA2        u0097(.A(men_men_n125_), .B(men_men_n117_), .Y(men_men_n126_));
  NO4        u0098(.A(men_men_n126_), .B(men_men_n124_), .C(men_men_n123_), .D(men_men_n120_), .Y(men_men_n127_));
  NO3        u0099(.A(men_men_n127_), .B(men_men_n119_), .C(men_men_n110_), .Y(men_men_n128_));
  OAI210     u0100(.A0(men_men_n105_), .A1(men_men_n88_), .B0(men_men_n128_), .Y(men_men_n129_));
  NOi31      u0101(.An(k), .B(m), .C(j), .Y(men_men_n130_));
  NA3        u0102(.A(men_men_n130_), .B(men_men_n79_), .C(men_men_n78_), .Y(men_men_n131_));
  NOi31      u0103(.An(k), .B(m), .C(i), .Y(men_men_n132_));
  NA3        u0104(.A(men_men_n132_), .B(men_men_n82_), .C(men_men_n78_), .Y(men_men_n133_));
  NA2        u0105(.A(men_men_n133_), .B(men_men_n131_), .Y(men_men_n134_));
  NOi32      u0106(.An(f), .Bn(b), .C(e), .Y(men_men_n135_));
  NAi21      u0107(.An(g), .B(h), .Y(men_men_n136_));
  NAi21      u0108(.An(m), .B(n), .Y(men_men_n137_));
  NAi21      u0109(.An(j), .B(k), .Y(men_men_n138_));
  NO3        u0110(.A(men_men_n138_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n139_));
  NAi41      u0111(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n140_));
  NAi31      u0112(.An(j), .B(k), .C(h), .Y(men_men_n141_));
  NO3        u0113(.A(men_men_n141_), .B(men_men_n140_), .C(men_men_n137_), .Y(men_men_n142_));
  AOI210     u0114(.A0(men_men_n139_), .A1(men_men_n135_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u0115(.A(k), .B(j), .Y(men_men_n144_));
  INV        u0116(.A(men_men_n137_), .Y(men_men_n145_));
  AN2        u0117(.A(k), .B(j), .Y(men_men_n146_));
  NAi21      u0118(.An(c), .B(b), .Y(men_men_n147_));
  NA2        u0119(.A(f), .B(d), .Y(men_men_n148_));
  NO4        u0120(.A(men_men_n148_), .B(men_men_n147_), .C(men_men_n146_), .D(men_men_n136_), .Y(men_men_n149_));
  NA2        u0121(.A(h), .B(c), .Y(men_men_n150_));
  NAi31      u0122(.An(f), .B(e), .C(b), .Y(men_men_n151_));
  NA2        u0123(.A(men_men_n149_), .B(men_men_n145_), .Y(men_men_n152_));
  NA2        u0124(.A(d), .B(b), .Y(men_men_n153_));
  NAi21      u0125(.An(e), .B(f), .Y(men_men_n154_));
  NO2        u0126(.A(men_men_n154_), .B(men_men_n153_), .Y(men_men_n155_));
  NA2        u0127(.A(b), .B(a), .Y(men_men_n156_));
  NAi21      u0128(.An(c), .B(d), .Y(men_men_n157_));
  NAi31      u0129(.An(l), .B(k), .C(h), .Y(men_men_n158_));
  NO2        u0130(.A(men_men_n137_), .B(men_men_n158_), .Y(men_men_n159_));
  NA2        u0131(.A(men_men_n159_), .B(men_men_n155_), .Y(men_men_n160_));
  NAi41      u0132(.An(men_men_n134_), .B(men_men_n160_), .C(men_men_n152_), .D(men_men_n143_), .Y(men_men_n161_));
  NAi31      u0133(.An(e), .B(f), .C(b), .Y(men_men_n162_));
  NOi21      u0134(.An(g), .B(d), .Y(men_men_n163_));
  NO2        u0135(.A(men_men_n163_), .B(men_men_n162_), .Y(men_men_n164_));
  NOi21      u0136(.An(h), .B(i), .Y(men_men_n165_));
  NOi21      u0137(.An(k), .B(m), .Y(men_men_n166_));
  NA2        u0138(.A(men_men_n166_), .B(men_men_n165_), .Y(men_men_n167_));
  NOi21      u0139(.An(men_men_n164_), .B(men_men_n167_), .Y(men_men_n168_));
  NOi21      u0140(.An(h), .B(g), .Y(men_men_n169_));
  NO2        u0141(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n170_));
  NA2        u0142(.A(men_men_n170_), .B(men_men_n169_), .Y(men_men_n171_));
  NAi31      u0143(.An(l), .B(j), .C(h), .Y(men_men_n172_));
  NO2        u0144(.A(men_men_n172_), .B(men_men_n49_), .Y(men_men_n173_));
  NA2        u0145(.A(men_men_n173_), .B(men_men_n67_), .Y(men_men_n174_));
  NOi32      u0146(.An(n), .Bn(k), .C(m), .Y(men_men_n175_));
  NA2        u0147(.A(l), .B(i), .Y(men_men_n176_));
  NA2        u0148(.A(men_men_n176_), .B(men_men_n175_), .Y(men_men_n177_));
  OAI210     u0149(.A0(men_men_n177_), .A1(men_men_n171_), .B0(men_men_n174_), .Y(men_men_n178_));
  NAi31      u0150(.An(e), .B(f), .C(c), .Y(men_men_n179_));
  NA2        u0151(.A(j), .B(h), .Y(men_men_n180_));
  OR3        u0152(.A(n), .B(m), .C(k), .Y(men_men_n181_));
  NAi32      u0153(.An(m), .Bn(k), .C(n), .Y(men_men_n182_));
  NO2        u0154(.A(men_men_n182_), .B(men_men_n180_), .Y(men_men_n183_));
  NA2        u0155(.A(men_men_n183_), .B(men_men_n164_), .Y(men_men_n184_));
  NO2        u0156(.A(n), .B(m), .Y(men_men_n185_));
  NA2        u0157(.A(men_men_n185_), .B(men_men_n50_), .Y(men_men_n186_));
  NAi21      u0158(.An(f), .B(e), .Y(men_men_n187_));
  NA2        u0159(.A(d), .B(c), .Y(men_men_n188_));
  NO2        u0160(.A(men_men_n188_), .B(men_men_n187_), .Y(men_men_n189_));
  NOi21      u0161(.An(men_men_n189_), .B(men_men_n186_), .Y(men_men_n190_));
  NAi21      u0162(.An(d), .B(c), .Y(men_men_n191_));
  NAi31      u0163(.An(m), .B(n), .C(b), .Y(men_men_n192_));
  NA2        u0164(.A(k), .B(i), .Y(men_men_n193_));
  NAi21      u0165(.An(h), .B(f), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(men_men_n193_), .Y(men_men_n195_));
  NO2        u0167(.A(men_men_n192_), .B(men_men_n157_), .Y(men_men_n196_));
  NA2        u0168(.A(men_men_n196_), .B(men_men_n195_), .Y(men_men_n197_));
  NOi32      u0169(.An(f), .Bn(c), .C(d), .Y(men_men_n198_));
  NOi32      u0170(.An(f), .Bn(c), .C(e), .Y(men_men_n199_));
  NO2        u0171(.A(men_men_n199_), .B(men_men_n198_), .Y(men_men_n200_));
  NO3        u0172(.A(n), .B(m), .C(j), .Y(men_men_n201_));
  NA2        u0173(.A(men_men_n201_), .B(men_men_n118_), .Y(men_men_n202_));
  NAi31      u0174(.An(men_men_n190_), .B(men_men_n197_), .C(men_men_n184_), .Y(men_men_n203_));
  OR4        u0175(.A(men_men_n203_), .B(men_men_n178_), .C(men_men_n168_), .D(men_men_n161_), .Y(men_men_n204_));
  NO4        u0176(.A(men_men_n204_), .B(men_men_n129_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n205_));
  NA3        u0177(.A(m), .B(men_men_n116_), .C(j), .Y(men_men_n206_));
  NAi31      u0178(.An(n), .B(h), .C(g), .Y(men_men_n207_));
  NO2        u0179(.A(men_men_n207_), .B(men_men_n206_), .Y(men_men_n208_));
  NOi32      u0180(.An(m), .Bn(k), .C(l), .Y(men_men_n209_));
  NA3        u0181(.A(men_men_n209_), .B(men_men_n89_), .C(g), .Y(men_men_n210_));
  NO2        u0182(.A(men_men_n210_), .B(n), .Y(men_men_n211_));
  NOi21      u0183(.An(k), .B(j), .Y(men_men_n212_));
  NA4        u0184(.A(men_men_n212_), .B(men_men_n117_), .C(i), .D(g), .Y(men_men_n213_));
  AN2        u0185(.A(i), .B(g), .Y(men_men_n214_));
  NA3        u0186(.A(men_men_n76_), .B(men_men_n214_), .C(men_men_n117_), .Y(men_men_n215_));
  NA2        u0187(.A(men_men_n215_), .B(men_men_n213_), .Y(men_men_n216_));
  NO3        u0188(.A(men_men_n216_), .B(men_men_n211_), .C(men_men_n208_), .Y(men_men_n217_));
  NAi41      u0189(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n218_));
  INV        u0190(.A(men_men_n218_), .Y(men_men_n219_));
  INV        u0191(.A(f), .Y(men_men_n220_));
  INV        u0192(.A(g), .Y(men_men_n221_));
  NOi31      u0193(.An(i), .B(j), .C(h), .Y(men_men_n222_));
  NOi21      u0194(.An(l), .B(m), .Y(men_men_n223_));
  NA2        u0195(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n224_));
  NO3        u0196(.A(men_men_n224_), .B(men_men_n221_), .C(men_men_n220_), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n219_), .Y(men_men_n226_));
  OAI210     u0198(.A0(men_men_n217_), .A1(men_men_n32_), .B0(men_men_n226_), .Y(men_men_n227_));
  NOi21      u0199(.An(n), .B(m), .Y(men_men_n228_));
  NOi32      u0200(.An(l), .Bn(i), .C(j), .Y(men_men_n229_));
  NA2        u0201(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  OA220      u0202(.A0(men_men_n230_), .A1(men_men_n109_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n231_));
  NAi21      u0203(.An(j), .B(h), .Y(men_men_n232_));
  XN2        u0204(.A(i), .B(h), .Y(men_men_n233_));
  NOi31      u0205(.An(k), .B(n), .C(m), .Y(men_men_n234_));
  NAi31      u0206(.An(f), .B(e), .C(c), .Y(men_men_n235_));
  NO4        u0207(.A(men_men_n235_), .B(men_men_n181_), .C(men_men_n180_), .D(men_men_n59_), .Y(men_men_n236_));
  NA4        u0208(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n237_));
  NAi32      u0209(.An(m), .Bn(i), .C(k), .Y(men_men_n238_));
  NO3        u0210(.A(men_men_n238_), .B(men_men_n93_), .C(men_men_n237_), .Y(men_men_n239_));
  NO2        u0211(.A(men_men_n239_), .B(men_men_n236_), .Y(men_men_n240_));
  NAi21      u0212(.An(n), .B(a), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n153_), .Y(men_men_n242_));
  NAi41      u0214(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n243_), .B(e), .Y(men_men_n244_));
  NO3        u0216(.A(men_men_n154_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n245_));
  OAI210     u0217(.A0(men_men_n245_), .A1(men_men_n244_), .B0(men_men_n242_), .Y(men_men_n246_));
  AN3        u0218(.A(men_men_n246_), .B(men_men_n240_), .C(men_men_n231_), .Y(men_men_n247_));
  OR2        u0219(.A(h), .B(g), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n248_), .B(men_men_n106_), .Y(men_men_n249_));
  NA2        u0221(.A(men_men_n249_), .B(men_men_n135_), .Y(men_men_n250_));
  NAi41      u0222(.An(e), .B(n), .C(d), .D(b), .Y(men_men_n251_));
  NO2        u0223(.A(men_men_n251_), .B(men_men_n220_), .Y(men_men_n252_));
  NA2        u0224(.A(men_men_n166_), .B(men_men_n112_), .Y(men_men_n253_));
  NAi21      u0225(.An(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NO2        u0226(.A(n), .B(a), .Y(men_men_n255_));
  NAi31      u0227(.An(men_men_n243_), .B(men_men_n255_), .C(men_men_n107_), .Y(men_men_n256_));
  AN2        u0228(.A(men_men_n256_), .B(men_men_n254_), .Y(men_men_n257_));
  NAi21      u0229(.An(h), .B(i), .Y(men_men_n258_));
  NA2        u0230(.A(men_men_n185_), .B(k), .Y(men_men_n259_));
  NO2        u0231(.A(men_men_n259_), .B(men_men_n258_), .Y(men_men_n260_));
  NA2        u0232(.A(men_men_n257_), .B(men_men_n250_), .Y(men_men_n261_));
  NOi21      u0233(.An(g), .B(e), .Y(men_men_n262_));
  NO2        u0234(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n263_));
  NA2        u0235(.A(men_men_n263_), .B(men_men_n262_), .Y(men_men_n264_));
  NOi32      u0236(.An(l), .Bn(j), .C(i), .Y(men_men_n265_));
  AOI210     u0237(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n265_), .Y(men_men_n266_));
  NO2        u0238(.A(men_men_n258_), .B(men_men_n44_), .Y(men_men_n267_));
  NAi21      u0239(.An(f), .B(g), .Y(men_men_n268_));
  NO2        u0240(.A(men_men_n268_), .B(men_men_n65_), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n69_), .B(men_men_n121_), .Y(men_men_n270_));
  AOI220     u0242(.A0(men_men_n270_), .A1(men_men_n269_), .B0(men_men_n267_), .B1(men_men_n67_), .Y(men_men_n271_));
  OAI210     u0243(.A0(men_men_n266_), .A1(men_men_n264_), .B0(men_men_n271_), .Y(men_men_n272_));
  NO3        u0244(.A(men_men_n138_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n273_));
  NOi41      u0245(.An(men_men_n247_), .B(men_men_n272_), .C(men_men_n261_), .D(men_men_n227_), .Y(men_men_n274_));
  NO4        u0246(.A(men_men_n208_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n275_));
  NO2        u0247(.A(men_men_n275_), .B(men_men_n115_), .Y(men_men_n276_));
  NA3        u0248(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n277_));
  NAi21      u0249(.An(h), .B(g), .Y(men_men_n278_));
  OR4        u0250(.A(men_men_n278_), .B(men_men_n277_), .C(men_men_n230_), .D(e), .Y(men_men_n279_));
  NO2        u0251(.A(men_men_n253_), .B(men_men_n268_), .Y(men_men_n280_));
  NA2        u0252(.A(men_men_n280_), .B(men_men_n78_), .Y(men_men_n281_));
  NAi31      u0253(.An(g), .B(k), .C(h), .Y(men_men_n282_));
  NO3        u0254(.A(men_men_n137_), .B(men_men_n282_), .C(l), .Y(men_men_n283_));
  NAi31      u0255(.An(e), .B(d), .C(a), .Y(men_men_n284_));
  NA2        u0256(.A(men_men_n283_), .B(men_men_n135_), .Y(men_men_n285_));
  NA3        u0257(.A(men_men_n285_), .B(men_men_n281_), .C(men_men_n279_), .Y(men_men_n286_));
  NA4        u0258(.A(men_men_n166_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n121_), .Y(men_men_n287_));
  NA3        u0259(.A(men_men_n166_), .B(men_men_n165_), .C(men_men_n86_), .Y(men_men_n288_));
  NO2        u0260(.A(men_men_n288_), .B(men_men_n200_), .Y(men_men_n289_));
  NOi21      u0261(.An(men_men_n287_), .B(men_men_n289_), .Y(men_men_n290_));
  NA3        u0262(.A(e), .B(c), .C(b), .Y(men_men_n291_));
  NO2        u0263(.A(men_men_n60_), .B(men_men_n291_), .Y(men_men_n292_));
  NAi32      u0264(.An(k), .Bn(i), .C(j), .Y(men_men_n293_));
  NAi31      u0265(.An(h), .B(l), .C(i), .Y(men_men_n294_));
  NA3        u0266(.A(men_men_n294_), .B(men_men_n293_), .C(men_men_n172_), .Y(men_men_n295_));
  NOi21      u0267(.An(men_men_n295_), .B(men_men_n49_), .Y(men_men_n296_));
  OAI210     u0268(.A0(men_men_n269_), .A1(men_men_n292_), .B0(men_men_n296_), .Y(men_men_n297_));
  NAi21      u0269(.An(l), .B(k), .Y(men_men_n298_));
  NO2        u0270(.A(men_men_n298_), .B(men_men_n49_), .Y(men_men_n299_));
  NOi21      u0271(.An(l), .B(j), .Y(men_men_n300_));
  NA2        u0272(.A(men_men_n169_), .B(men_men_n300_), .Y(men_men_n301_));
  NA3        u0273(.A(men_men_n122_), .B(men_men_n121_), .C(g), .Y(men_men_n302_));
  OR3        u0274(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n303_));
  AOI210     u0275(.A0(men_men_n302_), .A1(men_men_n301_), .B0(men_men_n303_), .Y(men_men_n304_));
  INV        u0276(.A(men_men_n304_), .Y(men_men_n305_));
  NAi32      u0277(.An(j), .Bn(h), .C(i), .Y(men_men_n306_));
  NAi21      u0278(.An(m), .B(l), .Y(men_men_n307_));
  NO3        u0279(.A(men_men_n307_), .B(men_men_n306_), .C(men_men_n86_), .Y(men_men_n308_));
  NA2        u0280(.A(h), .B(g), .Y(men_men_n309_));
  NA2        u0281(.A(men_men_n175_), .B(men_men_n45_), .Y(men_men_n310_));
  NO2        u0282(.A(men_men_n310_), .B(men_men_n309_), .Y(men_men_n311_));
  OAI210     u0283(.A0(men_men_n311_), .A1(men_men_n308_), .B0(men_men_n170_), .Y(men_men_n312_));
  NA4        u0284(.A(men_men_n312_), .B(men_men_n305_), .C(men_men_n297_), .D(men_men_n290_), .Y(men_men_n313_));
  NO2        u0285(.A(men_men_n151_), .B(d), .Y(men_men_n314_));
  NA2        u0286(.A(men_men_n314_), .B(men_men_n53_), .Y(men_men_n315_));
  NO2        u0287(.A(men_men_n109_), .B(men_men_n106_), .Y(men_men_n316_));
  NAi32      u0288(.An(n), .Bn(m), .C(l), .Y(men_men_n317_));
  NO2        u0289(.A(men_men_n317_), .B(men_men_n306_), .Y(men_men_n318_));
  NA2        u0290(.A(men_men_n318_), .B(men_men_n189_), .Y(men_men_n319_));
  NO2        u0291(.A(men_men_n126_), .B(men_men_n120_), .Y(men_men_n320_));
  NAi31      u0292(.An(k), .B(l), .C(j), .Y(men_men_n321_));
  OAI210     u0293(.A0(men_men_n298_), .A1(j), .B0(men_men_n321_), .Y(men_men_n322_));
  NOi21      u0294(.An(men_men_n322_), .B(men_men_n124_), .Y(men_men_n323_));
  NA2        u0295(.A(men_men_n323_), .B(men_men_n320_), .Y(men_men_n324_));
  NA3        u0296(.A(men_men_n324_), .B(men_men_n319_), .C(men_men_n315_), .Y(men_men_n325_));
  NO4        u0297(.A(men_men_n325_), .B(men_men_n313_), .C(men_men_n286_), .D(men_men_n276_), .Y(men_men_n326_));
  NA2        u0298(.A(men_men_n260_), .B(men_men_n199_), .Y(men_men_n327_));
  NAi21      u0299(.An(m), .B(k), .Y(men_men_n328_));
  NO2        u0300(.A(men_men_n233_), .B(men_men_n328_), .Y(men_men_n329_));
  NAi41      u0301(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n330_));
  NO2        u0302(.A(men_men_n330_), .B(e), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n331_), .B(men_men_n329_), .Y(men_men_n332_));
  NAi31      u0304(.An(i), .B(l), .C(h), .Y(men_men_n333_));
  NO4        u0305(.A(men_men_n333_), .B(e), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n334_));
  NA2        u0306(.A(e), .B(c), .Y(men_men_n335_));
  NO3        u0307(.A(men_men_n335_), .B(n), .C(d), .Y(men_men_n336_));
  NOi21      u0308(.An(f), .B(h), .Y(men_men_n337_));
  NA2        u0309(.A(men_men_n337_), .B(men_men_n122_), .Y(men_men_n338_));
  NO2        u0310(.A(men_men_n338_), .B(men_men_n221_), .Y(men_men_n339_));
  NAi31      u0311(.An(d), .B(e), .C(b), .Y(men_men_n340_));
  NO2        u0312(.A(men_men_n137_), .B(men_men_n340_), .Y(men_men_n341_));
  NA2        u0313(.A(men_men_n341_), .B(men_men_n339_), .Y(men_men_n342_));
  NAi41      u0314(.An(men_men_n334_), .B(men_men_n342_), .C(men_men_n332_), .D(men_men_n327_), .Y(men_men_n343_));
  NO4        u0315(.A(men_men_n330_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n221_), .Y(men_men_n344_));
  NA2        u0316(.A(men_men_n255_), .B(men_men_n107_), .Y(men_men_n345_));
  OR2        u0317(.A(men_men_n345_), .B(men_men_n210_), .Y(men_men_n346_));
  NOi31      u0318(.An(l), .B(n), .C(m), .Y(men_men_n347_));
  NA2        u0319(.A(men_men_n347_), .B(men_men_n222_), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n200_), .Y(men_men_n349_));
  NAi32      u0321(.An(men_men_n349_), .Bn(men_men_n344_), .C(men_men_n346_), .Y(men_men_n350_));
  NAi32      u0322(.An(m), .Bn(j), .C(k), .Y(men_men_n351_));
  NAi41      u0323(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n352_));
  OAI210     u0324(.A0(men_men_n218_), .A1(men_men_n351_), .B0(men_men_n352_), .Y(men_men_n353_));
  NOi31      u0325(.An(j), .B(m), .C(k), .Y(men_men_n354_));
  NO2        u0326(.A(men_men_n130_), .B(men_men_n354_), .Y(men_men_n355_));
  AN3        u0327(.A(h), .B(g), .C(f), .Y(men_men_n356_));
  NAi31      u0328(.An(men_men_n355_), .B(men_men_n356_), .C(men_men_n353_), .Y(men_men_n357_));
  NOi32      u0329(.An(m), .Bn(j), .C(l), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n358_), .B(men_men_n100_), .Y(men_men_n359_));
  NAi32      u0331(.An(men_men_n359_), .Bn(men_men_n207_), .C(men_men_n314_), .Y(men_men_n360_));
  NO2        u0332(.A(men_men_n307_), .B(men_men_n306_), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n224_), .B(g), .Y(men_men_n362_));
  INV        u0334(.A(men_men_n162_), .Y(men_men_n363_));
  AOI220     u0335(.A0(men_men_n363_), .A1(men_men_n362_), .B0(men_men_n252_), .B1(men_men_n361_), .Y(men_men_n364_));
  NA2        u0336(.A(men_men_n238_), .B(men_men_n81_), .Y(men_men_n365_));
  NA3        u0337(.A(men_men_n365_), .B(men_men_n356_), .C(men_men_n219_), .Y(men_men_n366_));
  NA4        u0338(.A(men_men_n366_), .B(men_men_n364_), .C(men_men_n360_), .D(men_men_n357_), .Y(men_men_n367_));
  NA3        u0339(.A(h), .B(g), .C(f), .Y(men_men_n368_));
  NO2        u0340(.A(men_men_n368_), .B(men_men_n77_), .Y(men_men_n369_));
  NA2        u0341(.A(men_men_n169_), .B(e), .Y(men_men_n370_));
  NO2        u0342(.A(men_men_n370_), .B(men_men_n41_), .Y(men_men_n371_));
  AOI220     u0343(.A0(men_men_n371_), .A1(men_men_n320_), .B0(b), .B1(men_men_n369_), .Y(men_men_n372_));
  NOi32      u0344(.An(j), .Bn(g), .C(i), .Y(men_men_n373_));
  NA3        u0345(.A(men_men_n373_), .B(men_men_n298_), .C(men_men_n117_), .Y(men_men_n374_));
  AO210      u0346(.A0(men_men_n115_), .A1(men_men_n32_), .B0(men_men_n374_), .Y(men_men_n375_));
  NOi32      u0347(.An(e), .Bn(b), .C(a), .Y(men_men_n376_));
  AN2        u0348(.A(l), .B(j), .Y(men_men_n377_));
  NO2        u0349(.A(men_men_n328_), .B(men_men_n377_), .Y(men_men_n378_));
  NO3        u0350(.A(men_men_n330_), .B(men_men_n72_), .C(men_men_n221_), .Y(men_men_n379_));
  NA3        u0351(.A(men_men_n215_), .B(men_men_n213_), .C(men_men_n35_), .Y(men_men_n380_));
  AOI220     u0352(.A0(men_men_n380_), .A1(men_men_n376_), .B0(men_men_n379_), .B1(men_men_n378_), .Y(men_men_n381_));
  NO2        u0353(.A(men_men_n340_), .B(n), .Y(men_men_n382_));
  NA2        u0354(.A(men_men_n214_), .B(k), .Y(men_men_n383_));
  NA3        u0355(.A(m), .B(men_men_n116_), .C(men_men_n220_), .Y(men_men_n384_));
  NA4        u0356(.A(men_men_n209_), .B(men_men_n89_), .C(g), .D(men_men_n220_), .Y(men_men_n385_));
  OAI210     u0357(.A0(men_men_n384_), .A1(men_men_n383_), .B0(men_men_n385_), .Y(men_men_n386_));
  NAi41      u0358(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n387_));
  NA2        u0359(.A(men_men_n51_), .B(men_men_n117_), .Y(men_men_n388_));
  NO2        u0360(.A(men_men_n388_), .B(men_men_n387_), .Y(men_men_n389_));
  AOI220     u0361(.A0(men_men_n389_), .A1(b), .B0(men_men_n386_), .B1(men_men_n382_), .Y(men_men_n390_));
  NA4        u0362(.A(men_men_n390_), .B(men_men_n381_), .C(men_men_n375_), .D(men_men_n372_), .Y(men_men_n391_));
  NO4        u0363(.A(men_men_n391_), .B(men_men_n367_), .C(men_men_n350_), .D(men_men_n343_), .Y(men_men_n392_));
  NA4        u0364(.A(men_men_n392_), .B(men_men_n326_), .C(men_men_n274_), .D(men_men_n205_), .Y(men10));
  NA3        u0365(.A(m), .B(k), .C(i), .Y(men_men_n394_));
  NO3        u0366(.A(men_men_n394_), .B(j), .C(men_men_n221_), .Y(men_men_n395_));
  NOi21      u0367(.An(e), .B(f), .Y(men_men_n396_));
  NO4        u0368(.A(men_men_n157_), .B(men_men_n396_), .C(n), .D(men_men_n114_), .Y(men_men_n397_));
  NAi31      u0369(.An(b), .B(f), .C(c), .Y(men_men_n398_));
  INV        u0370(.A(men_men_n398_), .Y(men_men_n399_));
  NOi32      u0371(.An(k), .Bn(h), .C(j), .Y(men_men_n400_));
  NA2        u0372(.A(men_men_n400_), .B(men_men_n228_), .Y(men_men_n401_));
  INV        u0373(.A(men_men_n401_), .Y(men_men_n402_));
  AOI220     u0374(.A0(men_men_n402_), .A1(men_men_n399_), .B0(men_men_n397_), .B1(men_men_n395_), .Y(men_men_n403_));
  AN2        u0375(.A(j), .B(h), .Y(men_men_n404_));
  NO3        u0376(.A(n), .B(m), .C(k), .Y(men_men_n405_));
  NA2        u0377(.A(men_men_n405_), .B(men_men_n404_), .Y(men_men_n406_));
  NO3        u0378(.A(men_men_n406_), .B(men_men_n157_), .C(men_men_n220_), .Y(men_men_n407_));
  OR2        u0379(.A(m), .B(k), .Y(men_men_n408_));
  NO2        u0380(.A(men_men_n180_), .B(men_men_n408_), .Y(men_men_n409_));
  NA4        u0381(.A(n), .B(f), .C(c), .D(men_men_n120_), .Y(men_men_n410_));
  NOi32      u0382(.An(d), .Bn(a), .C(c), .Y(men_men_n411_));
  NA2        u0383(.A(men_men_n411_), .B(men_men_n187_), .Y(men_men_n412_));
  NAi21      u0384(.An(i), .B(g), .Y(men_men_n413_));
  NAi31      u0385(.An(k), .B(m), .C(j), .Y(men_men_n414_));
  NO3        u0386(.A(men_men_n414_), .B(men_men_n413_), .C(n), .Y(men_men_n415_));
  NOi21      u0387(.An(men_men_n415_), .B(men_men_n412_), .Y(men_men_n416_));
  NO2        u0388(.A(men_men_n416_), .B(men_men_n407_), .Y(men_men_n417_));
  NO2        u0389(.A(men_men_n410_), .B(men_men_n307_), .Y(men_men_n418_));
  NOi32      u0390(.An(f), .Bn(d), .C(c), .Y(men_men_n419_));
  AOI220     u0391(.A0(men_men_n419_), .A1(men_men_n318_), .B0(men_men_n418_), .B1(men_men_n222_), .Y(men_men_n420_));
  NA3        u0392(.A(men_men_n420_), .B(men_men_n417_), .C(men_men_n403_), .Y(men_men_n421_));
  NO2        u0393(.A(men_men_n59_), .B(men_men_n120_), .Y(men_men_n422_));
  NA2        u0394(.A(men_men_n255_), .B(men_men_n422_), .Y(men_men_n423_));
  INV        u0395(.A(e), .Y(men_men_n424_));
  NA2        u0396(.A(men_men_n46_), .B(e), .Y(men_men_n425_));
  OAI220     u0397(.A0(men_men_n425_), .A1(men_men_n206_), .B0(men_men_n210_), .B1(men_men_n424_), .Y(men_men_n426_));
  AN2        u0398(.A(g), .B(e), .Y(men_men_n427_));
  NA3        u0399(.A(men_men_n427_), .B(men_men_n209_), .C(i), .Y(men_men_n428_));
  OAI210     u0400(.A0(men_men_n91_), .A1(men_men_n424_), .B0(men_men_n428_), .Y(men_men_n429_));
  NO2        u0401(.A(men_men_n103_), .B(men_men_n424_), .Y(men_men_n430_));
  NO3        u0402(.A(men_men_n430_), .B(men_men_n429_), .C(men_men_n426_), .Y(men_men_n431_));
  NOi32      u0403(.An(h), .Bn(e), .C(g), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n432_), .B(men_men_n300_), .C(m), .Y(men_men_n433_));
  NOi21      u0405(.An(g), .B(h), .Y(men_men_n434_));
  AN3        u0406(.A(m), .B(l), .C(i), .Y(men_men_n435_));
  NA3        u0407(.A(men_men_n435_), .B(men_men_n434_), .C(e), .Y(men_men_n436_));
  AN3        u0408(.A(h), .B(g), .C(e), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n437_), .B(men_men_n100_), .Y(men_men_n438_));
  AN3        u0410(.A(men_men_n438_), .B(men_men_n436_), .C(men_men_n433_), .Y(men_men_n439_));
  AOI210     u0411(.A0(men_men_n439_), .A1(men_men_n431_), .B0(men_men_n423_), .Y(men_men_n440_));
  NA3        u0412(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n441_));
  NO2        u0413(.A(men_men_n441_), .B(men_men_n423_), .Y(men_men_n442_));
  NA3        u0414(.A(men_men_n411_), .B(men_men_n187_), .C(men_men_n86_), .Y(men_men_n443_));
  NAi31      u0415(.An(b), .B(c), .C(a), .Y(men_men_n444_));
  NO2        u0416(.A(men_men_n444_), .B(n), .Y(men_men_n445_));
  OAI210     u0417(.A0(men_men_n51_), .A1(men_men_n50_), .B0(m), .Y(men_men_n446_));
  NO2        u0418(.A(men_men_n446_), .B(men_men_n154_), .Y(men_men_n447_));
  NA2        u0419(.A(men_men_n447_), .B(men_men_n445_), .Y(men_men_n448_));
  INV        u0420(.A(men_men_n448_), .Y(men_men_n449_));
  NO4        u0421(.A(men_men_n449_), .B(men_men_n442_), .C(men_men_n440_), .D(men_men_n421_), .Y(men_men_n450_));
  NA2        u0422(.A(i), .B(g), .Y(men_men_n451_));
  NO3        u0423(.A(men_men_n284_), .B(men_men_n451_), .C(c), .Y(men_men_n452_));
  NOi21      u0424(.An(a), .B(n), .Y(men_men_n453_));
  NOi21      u0425(.An(d), .B(c), .Y(men_men_n454_));
  NA2        u0426(.A(men_men_n454_), .B(men_men_n453_), .Y(men_men_n455_));
  NA3        u0427(.A(i), .B(g), .C(f), .Y(men_men_n456_));
  OR2        u0428(.A(men_men_n456_), .B(men_men_n71_), .Y(men_men_n457_));
  NA3        u0429(.A(men_men_n435_), .B(men_men_n434_), .C(men_men_n187_), .Y(men_men_n458_));
  AOI210     u0430(.A0(men_men_n458_), .A1(men_men_n457_), .B0(men_men_n455_), .Y(men_men_n459_));
  AOI210     u0431(.A0(men_men_n452_), .A1(men_men_n299_), .B0(men_men_n459_), .Y(men_men_n460_));
  OR2        u0432(.A(n), .B(m), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n461_), .B(men_men_n158_), .Y(men_men_n462_));
  NO2        u0434(.A(men_men_n188_), .B(men_men_n154_), .Y(men_men_n463_));
  NA2        u0435(.A(men_men_n462_), .B(men_men_n463_), .Y(men_men_n464_));
  INV        u0436(.A(men_men_n388_), .Y(men_men_n465_));
  NA3        u0437(.A(men_men_n465_), .B(men_men_n376_), .C(d), .Y(men_men_n466_));
  NO2        u0438(.A(men_men_n444_), .B(men_men_n49_), .Y(men_men_n467_));
  NO3        u0439(.A(men_men_n66_), .B(men_men_n116_), .C(e), .Y(men_men_n468_));
  NAi21      u0440(.An(k), .B(j), .Y(men_men_n469_));
  NA2        u0441(.A(men_men_n258_), .B(men_men_n469_), .Y(men_men_n470_));
  NA3        u0442(.A(men_men_n470_), .B(men_men_n468_), .C(men_men_n467_), .Y(men_men_n471_));
  NAi21      u0443(.An(e), .B(d), .Y(men_men_n472_));
  NO2        u0444(.A(men_men_n472_), .B(men_men_n56_), .Y(men_men_n473_));
  NA3        u0445(.A(men_men_n471_), .B(men_men_n466_), .C(men_men_n464_), .Y(men_men_n474_));
  NO2        u0446(.A(men_men_n348_), .B(men_men_n220_), .Y(men_men_n475_));
  NA2        u0447(.A(men_men_n475_), .B(men_men_n473_), .Y(men_men_n476_));
  NOi31      u0448(.An(n), .B(m), .C(k), .Y(men_men_n477_));
  AOI220     u0449(.A0(men_men_n477_), .A1(men_men_n404_), .B0(men_men_n228_), .B1(men_men_n50_), .Y(men_men_n478_));
  NAi31      u0450(.An(g), .B(f), .C(c), .Y(men_men_n479_));
  OR3        u0451(.A(men_men_n479_), .B(men_men_n478_), .C(e), .Y(men_men_n480_));
  NA3        u0452(.A(men_men_n480_), .B(men_men_n476_), .C(men_men_n319_), .Y(men_men_n481_));
  NOi41      u0453(.An(men_men_n460_), .B(men_men_n481_), .C(men_men_n474_), .D(men_men_n272_), .Y(men_men_n482_));
  NOi32      u0454(.An(c), .Bn(a), .C(b), .Y(men_men_n483_));
  NA2        u0455(.A(men_men_n483_), .B(men_men_n117_), .Y(men_men_n484_));
  INV        u0456(.A(men_men_n282_), .Y(men_men_n485_));
  AN2        u0457(.A(e), .B(d), .Y(men_men_n486_));
  NA2        u0458(.A(men_men_n486_), .B(men_men_n485_), .Y(men_men_n487_));
  INV        u0459(.A(men_men_n154_), .Y(men_men_n488_));
  NO2        u0460(.A(men_men_n136_), .B(men_men_n41_), .Y(men_men_n489_));
  NO2        u0461(.A(men_men_n66_), .B(e), .Y(men_men_n490_));
  NOi31      u0462(.An(j), .B(k), .C(i), .Y(men_men_n491_));
  NOi21      u0463(.An(men_men_n172_), .B(men_men_n491_), .Y(men_men_n492_));
  NA4        u0464(.A(men_men_n333_), .B(men_men_n492_), .C(men_men_n266_), .D(men_men_n123_), .Y(men_men_n493_));
  AOI220     u0465(.A0(men_men_n493_), .A1(men_men_n490_), .B0(men_men_n489_), .B1(men_men_n488_), .Y(men_men_n494_));
  AOI210     u0466(.A0(men_men_n494_), .A1(men_men_n487_), .B0(men_men_n484_), .Y(men_men_n495_));
  NO2        u0467(.A(men_men_n216_), .B(men_men_n211_), .Y(men_men_n496_));
  NOi21      u0468(.An(a), .B(b), .Y(men_men_n497_));
  NA3        u0469(.A(e), .B(d), .C(c), .Y(men_men_n498_));
  NAi21      u0470(.An(men_men_n498_), .B(men_men_n497_), .Y(men_men_n499_));
  NO2        u0471(.A(men_men_n443_), .B(men_men_n210_), .Y(men_men_n500_));
  NOi21      u0472(.An(men_men_n499_), .B(men_men_n500_), .Y(men_men_n501_));
  AOI210     u0473(.A0(men_men_n275_), .A1(men_men_n496_), .B0(men_men_n501_), .Y(men_men_n502_));
  NA2        u0474(.A(men_men_n399_), .B(men_men_n159_), .Y(men_men_n503_));
  OR2        u0475(.A(k), .B(j), .Y(men_men_n504_));
  NA2        u0476(.A(l), .B(k), .Y(men_men_n505_));
  NA3        u0477(.A(men_men_n505_), .B(men_men_n504_), .C(men_men_n228_), .Y(men_men_n506_));
  NA2        u0478(.A(men_men_n238_), .B(men_men_n351_), .Y(men_men_n507_));
  NOi21      u0479(.An(men_men_n506_), .B(men_men_n507_), .Y(men_men_n508_));
  OR3        u0480(.A(men_men_n508_), .B(men_men_n150_), .C(men_men_n140_), .Y(men_men_n509_));
  NA3        u0481(.A(men_men_n287_), .B(men_men_n133_), .C(men_men_n131_), .Y(men_men_n510_));
  NA2        u0482(.A(men_men_n411_), .B(men_men_n117_), .Y(men_men_n511_));
  NO4        u0483(.A(men_men_n511_), .B(men_men_n97_), .C(men_men_n116_), .D(e), .Y(men_men_n512_));
  NO3        u0484(.A(men_men_n443_), .B(men_men_n94_), .C(men_men_n136_), .Y(men_men_n513_));
  NO4        u0485(.A(men_men_n513_), .B(men_men_n512_), .C(men_men_n510_), .D(men_men_n334_), .Y(men_men_n514_));
  NA3        u0486(.A(men_men_n514_), .B(men_men_n509_), .C(men_men_n503_), .Y(men_men_n515_));
  NO3        u0487(.A(men_men_n515_), .B(men_men_n502_), .C(men_men_n495_), .Y(men_men_n516_));
  NA2        u0488(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n517_));
  NOi21      u0489(.An(d), .B(e), .Y(men_men_n518_));
  NO2        u0490(.A(men_men_n194_), .B(men_men_n56_), .Y(men_men_n519_));
  NAi31      u0491(.An(j), .B(l), .C(i), .Y(men_men_n520_));
  OAI210     u0492(.A0(men_men_n520_), .A1(men_men_n137_), .B0(men_men_n106_), .Y(men_men_n521_));
  NA4        u0493(.A(men_men_n521_), .B(men_men_n519_), .C(men_men_n518_), .D(b), .Y(men_men_n522_));
  NO3        u0494(.A(men_men_n412_), .B(men_men_n359_), .C(men_men_n207_), .Y(men_men_n523_));
  NO2        u0495(.A(men_men_n412_), .B(men_men_n388_), .Y(men_men_n524_));
  NO4        u0496(.A(men_men_n524_), .B(men_men_n523_), .C(men_men_n190_), .D(men_men_n316_), .Y(men_men_n525_));
  NA4        u0497(.A(men_men_n525_), .B(men_men_n522_), .C(men_men_n517_), .D(men_men_n247_), .Y(men_men_n526_));
  OAI210     u0498(.A0(men_men_n132_), .A1(men_men_n130_), .B0(n), .Y(men_men_n527_));
  NO2        u0499(.A(men_men_n527_), .B(men_men_n136_), .Y(men_men_n528_));
  OR2        u0500(.A(men_men_n308_), .B(men_men_n249_), .Y(men_men_n529_));
  AN2        u0501(.A(men_men_n529_), .B(men_men_n199_), .Y(men_men_n530_));
  XO2        u0502(.A(i), .B(h), .Y(men_men_n531_));
  NA3        u0503(.A(men_men_n531_), .B(men_men_n166_), .C(n), .Y(men_men_n532_));
  NAi41      u0504(.An(men_men_n308_), .B(men_men_n532_), .C(men_men_n478_), .D(men_men_n401_), .Y(men_men_n533_));
  NOi32      u0505(.An(men_men_n533_), .Bn(men_men_n490_), .C(men_men_n277_), .Y(men_men_n534_));
  NAi31      u0506(.An(c), .B(f), .C(d), .Y(men_men_n535_));
  NO2        u0507(.A(men_men_n288_), .B(men_men_n535_), .Y(men_men_n536_));
  BUFFER     u0508(.A(men_men_n84_), .Y(men_men_n537_));
  NA3        u0509(.A(men_men_n397_), .B(men_men_n100_), .C(men_men_n99_), .Y(men_men_n538_));
  NA2        u0510(.A(men_men_n234_), .B(men_men_n112_), .Y(men_men_n539_));
  AOI210     u0511(.A0(men_men_n539_), .A1(men_men_n186_), .B0(men_men_n535_), .Y(men_men_n540_));
  AOI210     u0512(.A0(men_men_n374_), .A1(men_men_n35_), .B0(men_men_n499_), .Y(men_men_n541_));
  NOi31      u0513(.An(men_men_n538_), .B(men_men_n541_), .C(men_men_n540_), .Y(men_men_n542_));
  AO220      u0514(.A0(men_men_n296_), .A1(men_men_n269_), .B0(men_men_n173_), .B1(men_men_n67_), .Y(men_men_n543_));
  NA3        u0515(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n544_));
  NO2        u0516(.A(men_men_n544_), .B(men_men_n455_), .Y(men_men_n545_));
  NO2        u0517(.A(men_men_n545_), .B(men_men_n304_), .Y(men_men_n546_));
  NAi41      u0518(.An(men_men_n543_), .B(men_men_n546_), .C(men_men_n542_), .D(men_men_n537_), .Y(men_men_n547_));
  NO4        u0519(.A(men_men_n547_), .B(men_men_n534_), .C(men_men_n530_), .D(men_men_n526_), .Y(men_men_n548_));
  NA4        u0520(.A(men_men_n548_), .B(men_men_n516_), .C(men_men_n482_), .D(men_men_n450_), .Y(men11));
  NO2        u0521(.A(men_men_n73_), .B(f), .Y(men_men_n550_));
  NA2        u0522(.A(j), .B(g), .Y(men_men_n551_));
  NAi31      u0523(.An(i), .B(m), .C(l), .Y(men_men_n552_));
  NA3        u0524(.A(m), .B(k), .C(j), .Y(men_men_n553_));
  OAI220     u0525(.A0(men_men_n553_), .A1(men_men_n136_), .B0(men_men_n552_), .B1(men_men_n551_), .Y(men_men_n554_));
  NA2        u0526(.A(men_men_n554_), .B(men_men_n550_), .Y(men_men_n555_));
  NOi32      u0527(.An(e), .Bn(b), .C(f), .Y(men_men_n556_));
  NA2        u0528(.A(men_men_n265_), .B(men_men_n117_), .Y(men_men_n557_));
  NA2        u0529(.A(men_men_n46_), .B(j), .Y(men_men_n558_));
  NO2        u0530(.A(men_men_n558_), .B(men_men_n310_), .Y(men_men_n559_));
  NAi31      u0531(.An(d), .B(e), .C(a), .Y(men_men_n560_));
  NO2        u0532(.A(men_men_n560_), .B(n), .Y(men_men_n561_));
  AOI220     u0533(.A0(men_men_n561_), .A1(men_men_n104_), .B0(men_men_n559_), .B1(men_men_n556_), .Y(men_men_n562_));
  NAi41      u0534(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n563_));
  AN2        u0535(.A(men_men_n563_), .B(men_men_n387_), .Y(men_men_n564_));
  AOI210     u0536(.A0(men_men_n564_), .A1(men_men_n412_), .B0(men_men_n278_), .Y(men_men_n565_));
  NA2        u0537(.A(j), .B(i), .Y(men_men_n566_));
  NAi31      u0538(.An(n), .B(m), .C(k), .Y(men_men_n567_));
  NO3        u0539(.A(men_men_n567_), .B(men_men_n566_), .C(men_men_n116_), .Y(men_men_n568_));
  NO4        u0540(.A(n), .B(d), .C(men_men_n120_), .D(a), .Y(men_men_n569_));
  OR2        u0541(.A(n), .B(c), .Y(men_men_n570_));
  NO2        u0542(.A(men_men_n570_), .B(men_men_n156_), .Y(men_men_n571_));
  NO2        u0543(.A(men_men_n571_), .B(men_men_n569_), .Y(men_men_n572_));
  NOi32      u0544(.An(g), .Bn(f), .C(i), .Y(men_men_n573_));
  AOI220     u0545(.A0(men_men_n573_), .A1(men_men_n102_), .B0(men_men_n554_), .B1(f), .Y(men_men_n574_));
  NO2        u0546(.A(men_men_n282_), .B(men_men_n49_), .Y(men_men_n575_));
  NO2        u0547(.A(men_men_n574_), .B(men_men_n572_), .Y(men_men_n576_));
  AOI210     u0548(.A0(men_men_n568_), .A1(men_men_n565_), .B0(men_men_n576_), .Y(men_men_n577_));
  NA2        u0549(.A(men_men_n146_), .B(men_men_n34_), .Y(men_men_n578_));
  OAI220     u0550(.A0(men_men_n578_), .A1(m), .B0(men_men_n558_), .B1(men_men_n238_), .Y(men_men_n579_));
  NOi41      u0551(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n580_));
  NAi32      u0552(.An(e), .Bn(b), .C(c), .Y(men_men_n581_));
  AN2        u0553(.A(men_men_n352_), .B(men_men_n330_), .Y(men_men_n582_));
  NA2        u0554(.A(men_men_n582_), .B(men_men_n581_), .Y(men_men_n583_));
  OA210      u0555(.A0(men_men_n583_), .A1(men_men_n580_), .B0(men_men_n579_), .Y(men_men_n584_));
  OAI220     u0556(.A0(men_men_n414_), .A1(men_men_n413_), .B0(men_men_n552_), .B1(men_men_n551_), .Y(men_men_n585_));
  NAi31      u0557(.An(d), .B(c), .C(a), .Y(men_men_n586_));
  NO2        u0558(.A(men_men_n586_), .B(n), .Y(men_men_n587_));
  NA3        u0559(.A(men_men_n587_), .B(men_men_n585_), .C(e), .Y(men_men_n588_));
  NO3        u0560(.A(men_men_n62_), .B(men_men_n49_), .C(men_men_n221_), .Y(men_men_n589_));
  NO2        u0561(.A(men_men_n235_), .B(men_men_n114_), .Y(men_men_n590_));
  OAI210     u0562(.A0(men_men_n589_), .A1(men_men_n415_), .B0(men_men_n590_), .Y(men_men_n591_));
  NA2        u0563(.A(men_men_n591_), .B(men_men_n588_), .Y(men_men_n592_));
  NO2        u0564(.A(men_men_n284_), .B(n), .Y(men_men_n593_));
  NO2        u0565(.A(men_men_n445_), .B(men_men_n593_), .Y(men_men_n594_));
  NA2        u0566(.A(men_men_n585_), .B(f), .Y(men_men_n595_));
  NAi32      u0567(.An(d), .Bn(a), .C(b), .Y(men_men_n596_));
  NO2        u0568(.A(men_men_n596_), .B(men_men_n49_), .Y(men_men_n597_));
  NA2        u0569(.A(h), .B(f), .Y(men_men_n598_));
  NO2        u0570(.A(men_men_n598_), .B(men_men_n97_), .Y(men_men_n599_));
  NO3        u0571(.A(men_men_n182_), .B(men_men_n180_), .C(g), .Y(men_men_n600_));
  AOI220     u0572(.A0(men_men_n600_), .A1(men_men_n58_), .B0(men_men_n599_), .B1(men_men_n597_), .Y(men_men_n601_));
  OAI210     u0573(.A0(men_men_n595_), .A1(men_men_n594_), .B0(men_men_n601_), .Y(men_men_n602_));
  AN3        u0574(.A(j), .B(h), .C(g), .Y(men_men_n603_));
  NO2        u0575(.A(men_men_n153_), .B(c), .Y(men_men_n604_));
  NA3        u0576(.A(men_men_n604_), .B(men_men_n603_), .C(men_men_n477_), .Y(men_men_n605_));
  NA3        u0577(.A(f), .B(d), .C(b), .Y(men_men_n606_));
  NO4        u0578(.A(men_men_n606_), .B(men_men_n182_), .C(men_men_n180_), .D(g), .Y(men_men_n607_));
  NAi21      u0579(.An(men_men_n607_), .B(men_men_n605_), .Y(men_men_n608_));
  NO4        u0580(.A(men_men_n608_), .B(men_men_n602_), .C(men_men_n592_), .D(men_men_n584_), .Y(men_men_n609_));
  AN4        u0581(.A(men_men_n609_), .B(men_men_n577_), .C(men_men_n562_), .D(men_men_n555_), .Y(men_men_n610_));
  INV        u0582(.A(k), .Y(men_men_n611_));
  NA3        u0583(.A(l), .B(men_men_n611_), .C(i), .Y(men_men_n612_));
  INV        u0584(.A(men_men_n612_), .Y(men_men_n613_));
  NA4        u0585(.A(men_men_n411_), .B(men_men_n434_), .C(men_men_n187_), .D(men_men_n117_), .Y(men_men_n614_));
  NAi32      u0586(.An(h), .Bn(f), .C(g), .Y(men_men_n615_));
  NAi41      u0587(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n616_));
  OAI210     u0588(.A0(men_men_n560_), .A1(n), .B0(men_men_n616_), .Y(men_men_n617_));
  NA2        u0589(.A(men_men_n617_), .B(m), .Y(men_men_n618_));
  NAi31      u0590(.An(h), .B(g), .C(f), .Y(men_men_n619_));
  OR3        u0591(.A(men_men_n619_), .B(men_men_n284_), .C(men_men_n49_), .Y(men_men_n620_));
  NA4        u0592(.A(men_men_n434_), .B(men_men_n125_), .C(men_men_n117_), .D(e), .Y(men_men_n621_));
  AN2        u0593(.A(men_men_n621_), .B(men_men_n620_), .Y(men_men_n622_));
  OA210      u0594(.A0(men_men_n618_), .A1(men_men_n615_), .B0(men_men_n622_), .Y(men_men_n623_));
  NO3        u0595(.A(men_men_n615_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n624_));
  NO4        u0596(.A(men_men_n619_), .B(men_men_n570_), .C(men_men_n156_), .D(men_men_n75_), .Y(men_men_n625_));
  OR2        u0597(.A(men_men_n625_), .B(men_men_n624_), .Y(men_men_n626_));
  NAi31      u0598(.An(men_men_n626_), .B(men_men_n623_), .C(men_men_n614_), .Y(men_men_n627_));
  NAi31      u0599(.An(f), .B(h), .C(g), .Y(men_men_n628_));
  NO4        u0600(.A(men_men_n321_), .B(men_men_n628_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n629_));
  NOi32      u0601(.An(b), .Bn(a), .C(c), .Y(men_men_n630_));
  NOi41      u0602(.An(men_men_n630_), .B(men_men_n368_), .C(men_men_n69_), .D(men_men_n121_), .Y(men_men_n631_));
  OR2        u0603(.A(men_men_n631_), .B(men_men_n629_), .Y(men_men_n632_));
  NOi32      u0604(.An(d), .Bn(a), .C(e), .Y(men_men_n633_));
  NA2        u0605(.A(men_men_n633_), .B(men_men_n117_), .Y(men_men_n634_));
  NO2        u0606(.A(n), .B(c), .Y(men_men_n635_));
  NA3        u0607(.A(men_men_n635_), .B(men_men_n29_), .C(m), .Y(men_men_n636_));
  NOi32      u0608(.An(e), .Bn(a), .C(d), .Y(men_men_n637_));
  AOI210     u0609(.A0(men_men_n29_), .A1(d), .B0(men_men_n637_), .Y(men_men_n638_));
  AOI210     u0610(.A0(men_men_n638_), .A1(men_men_n220_), .B0(men_men_n578_), .Y(men_men_n639_));
  AOI210     u0611(.A0(men_men_n639_), .A1(men_men_n117_), .B0(men_men_n632_), .Y(men_men_n640_));
  INV        u0612(.A(men_men_n640_), .Y(men_men_n641_));
  AOI210     u0613(.A0(men_men_n627_), .A1(men_men_n613_), .B0(men_men_n641_), .Y(men_men_n642_));
  NO3        u0614(.A(men_men_n328_), .B(men_men_n61_), .C(n), .Y(men_men_n643_));
  NA2        u0615(.A(men_men_n76_), .B(men_men_n117_), .Y(men_men_n644_));
  NO2        u0616(.A(men_men_n644_), .B(men_men_n45_), .Y(men_men_n645_));
  AOI220     u0617(.A0(men_men_n645_), .A1(men_men_n565_), .B0(f), .B1(men_men_n643_), .Y(men_men_n646_));
  NO2        u0618(.A(men_men_n646_), .B(men_men_n89_), .Y(men_men_n647_));
  NA3        u0619(.A(men_men_n580_), .B(men_men_n354_), .C(men_men_n46_), .Y(men_men_n648_));
  NOi32      u0620(.An(e), .Bn(c), .C(f), .Y(men_men_n649_));
  NOi21      u0621(.An(f), .B(g), .Y(men_men_n650_));
  NO2        u0622(.A(men_men_n650_), .B(men_men_n218_), .Y(men_men_n651_));
  NA2        u0623(.A(men_men_n651_), .B(men_men_n409_), .Y(men_men_n652_));
  NA3        u0624(.A(men_men_n652_), .B(men_men_n648_), .C(men_men_n184_), .Y(men_men_n653_));
  AOI210     u0625(.A0(men_men_n564_), .A1(men_men_n412_), .B0(men_men_n309_), .Y(men_men_n654_));
  NA2        u0626(.A(men_men_n654_), .B(men_men_n270_), .Y(men_men_n655_));
  NOi21      u0627(.An(j), .B(l), .Y(men_men_n656_));
  NAi21      u0628(.An(k), .B(h), .Y(men_men_n657_));
  NO2        u0629(.A(men_men_n657_), .B(men_men_n268_), .Y(men_men_n658_));
  NA2        u0630(.A(men_men_n658_), .B(men_men_n656_), .Y(men_men_n659_));
  OR2        u0631(.A(men_men_n659_), .B(men_men_n618_), .Y(men_men_n660_));
  NOi31      u0632(.An(m), .B(n), .C(k), .Y(men_men_n661_));
  NA2        u0633(.A(men_men_n656_), .B(men_men_n661_), .Y(men_men_n662_));
  AOI210     u0634(.A0(men_men_n412_), .A1(men_men_n387_), .B0(men_men_n309_), .Y(men_men_n663_));
  NAi21      u0635(.An(men_men_n662_), .B(men_men_n663_), .Y(men_men_n664_));
  NO2        u0636(.A(men_men_n284_), .B(men_men_n49_), .Y(men_men_n665_));
  NO2        u0637(.A(men_men_n321_), .B(men_men_n628_), .Y(men_men_n666_));
  NO2        u0638(.A(men_men_n560_), .B(men_men_n49_), .Y(men_men_n667_));
  AOI220     u0639(.A0(men_men_n667_), .A1(men_men_n666_), .B0(men_men_n665_), .B1(men_men_n599_), .Y(men_men_n668_));
  NA4        u0640(.A(men_men_n668_), .B(men_men_n664_), .C(men_men_n660_), .D(men_men_n655_), .Y(men_men_n669_));
  NA2        u0641(.A(men_men_n112_), .B(men_men_n36_), .Y(men_men_n670_));
  NO2        u0642(.A(k), .B(men_men_n221_), .Y(men_men_n671_));
  NO2        u0643(.A(men_men_n556_), .B(men_men_n376_), .Y(men_men_n672_));
  NO2        u0644(.A(men_men_n672_), .B(n), .Y(men_men_n673_));
  NAi31      u0645(.An(men_men_n670_), .B(men_men_n673_), .C(men_men_n671_), .Y(men_men_n674_));
  NO2        u0646(.A(men_men_n558_), .B(men_men_n182_), .Y(men_men_n675_));
  NA3        u0647(.A(men_men_n581_), .B(men_men_n277_), .C(men_men_n151_), .Y(men_men_n676_));
  NA2        u0648(.A(men_men_n531_), .B(men_men_n166_), .Y(men_men_n677_));
  NA2        u0649(.A(men_men_n676_), .B(men_men_n675_), .Y(men_men_n678_));
  AN3        u0650(.A(f), .B(d), .C(b), .Y(men_men_n679_));
  NO2        u0651(.A(men_men_n679_), .B(men_men_n135_), .Y(men_men_n680_));
  NA3        u0652(.A(men_men_n531_), .B(men_men_n166_), .C(men_men_n221_), .Y(men_men_n681_));
  AOI210     u0653(.A0(men_men_n680_), .A1(men_men_n237_), .B0(men_men_n681_), .Y(men_men_n682_));
  NAi31      u0654(.An(m), .B(n), .C(k), .Y(men_men_n683_));
  OAI210     u0655(.A0(men_men_n140_), .A1(men_men_n683_), .B0(men_men_n256_), .Y(men_men_n684_));
  OAI210     u0656(.A0(men_men_n684_), .A1(men_men_n682_), .B0(j), .Y(men_men_n685_));
  NA3        u0657(.A(men_men_n685_), .B(men_men_n678_), .C(men_men_n674_), .Y(men_men_n686_));
  NO4        u0658(.A(men_men_n686_), .B(men_men_n669_), .C(men_men_n653_), .D(men_men_n647_), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n397_), .B(men_men_n169_), .Y(men_men_n688_));
  NAi31      u0660(.An(g), .B(h), .C(f), .Y(men_men_n689_));
  OR3        u0661(.A(men_men_n689_), .B(men_men_n284_), .C(n), .Y(men_men_n690_));
  OA210      u0662(.A0(men_men_n560_), .A1(n), .B0(men_men_n616_), .Y(men_men_n691_));
  NA3        u0663(.A(men_men_n432_), .B(men_men_n125_), .C(men_men_n86_), .Y(men_men_n692_));
  OAI210     u0664(.A0(men_men_n691_), .A1(men_men_n93_), .B0(men_men_n692_), .Y(men_men_n693_));
  NOi21      u0665(.An(men_men_n690_), .B(men_men_n693_), .Y(men_men_n694_));
  AOI210     u0666(.A0(men_men_n694_), .A1(men_men_n688_), .B0(men_men_n553_), .Y(men_men_n695_));
  NO3        u0667(.A(g), .B(men_men_n220_), .C(men_men_n56_), .Y(men_men_n696_));
  NAi21      u0668(.An(h), .B(j), .Y(men_men_n697_));
  NO2        u0669(.A(men_men_n539_), .B(men_men_n89_), .Y(men_men_n698_));
  OAI210     u0670(.A0(men_men_n698_), .A1(men_men_n409_), .B0(men_men_n696_), .Y(men_men_n699_));
  OR2        u0671(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n700_));
  NA2        u0672(.A(men_men_n630_), .B(men_men_n356_), .Y(men_men_n701_));
  OA220      u0673(.A0(men_men_n662_), .A1(men_men_n701_), .B0(men_men_n659_), .B1(men_men_n700_), .Y(men_men_n702_));
  NA3        u0674(.A(men_men_n550_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n703_));
  AN2        u0675(.A(h), .B(f), .Y(men_men_n704_));
  NA2        u0676(.A(men_men_n704_), .B(men_men_n37_), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n706_));
  OAI220     u0678(.A0(men_men_n706_), .A1(men_men_n345_), .B0(men_men_n705_), .B1(men_men_n484_), .Y(men_men_n707_));
  AOI210     u0679(.A0(men_men_n596_), .A1(men_men_n444_), .B0(men_men_n49_), .Y(men_men_n708_));
  NO2        u0680(.A(men_men_n619_), .B(men_men_n612_), .Y(men_men_n709_));
  AOI210     u0681(.A0(men_men_n709_), .A1(men_men_n708_), .B0(men_men_n707_), .Y(men_men_n710_));
  NA4        u0682(.A(men_men_n710_), .B(men_men_n703_), .C(men_men_n702_), .D(men_men_n699_), .Y(men_men_n711_));
  NO2        u0683(.A(men_men_n258_), .B(f), .Y(men_men_n712_));
  NA2        u0684(.A(men_men_n341_), .B(men_men_n146_), .Y(men_men_n713_));
  NA2        u0685(.A(men_men_n137_), .B(men_men_n49_), .Y(men_men_n714_));
  OA220      u0686(.A0(men_men_n1595_), .A1(men_men_n578_), .B0(men_men_n374_), .B1(men_men_n115_), .Y(men_men_n715_));
  OAI210     u0687(.A0(men_men_n713_), .A1(men_men_n650_), .B0(men_men_n715_), .Y(men_men_n716_));
  NA2        u0688(.A(men_men_n483_), .B(men_men_n86_), .Y(men_men_n717_));
  NO4        u0689(.A(men_men_n553_), .B(men_men_n717_), .C(men_men_n136_), .D(men_men_n220_), .Y(men_men_n718_));
  INV        u0690(.A(men_men_n718_), .Y(men_men_n719_));
  NA3        u0691(.A(men_men_n719_), .B(men_men_n538_), .C(men_men_n417_), .Y(men_men_n720_));
  NO4        u0692(.A(men_men_n720_), .B(men_men_n716_), .C(men_men_n711_), .D(men_men_n695_), .Y(men_men_n721_));
  NA4        u0693(.A(men_men_n721_), .B(men_men_n687_), .C(men_men_n642_), .D(men_men_n610_), .Y(men08));
  NO2        u0694(.A(k), .B(h), .Y(men_men_n723_));
  AO210      u0695(.A0(men_men_n258_), .A1(men_men_n469_), .B0(men_men_n723_), .Y(men_men_n724_));
  NO2        u0696(.A(men_men_n724_), .B(men_men_n307_), .Y(men_men_n725_));
  NA2        u0697(.A(men_men_n649_), .B(men_men_n86_), .Y(men_men_n726_));
  AOI210     u0698(.A0(men_men_n1600_), .A1(men_men_n725_), .B0(men_men_n513_), .Y(men_men_n727_));
  NA2        u0699(.A(men_men_n86_), .B(men_men_n114_), .Y(men_men_n728_));
  NO2        u0700(.A(men_men_n728_), .B(men_men_n57_), .Y(men_men_n729_));
  NO4        u0701(.A(men_men_n394_), .B(men_men_n116_), .C(j), .D(men_men_n221_), .Y(men_men_n730_));
  NA2        u0702(.A(men_men_n606_), .B(men_men_n237_), .Y(men_men_n731_));
  AOI220     u0703(.A0(men_men_n731_), .A1(men_men_n362_), .B0(men_men_n730_), .B1(men_men_n729_), .Y(men_men_n732_));
  AOI210     u0704(.A0(men_men_n606_), .A1(men_men_n162_), .B0(men_men_n86_), .Y(men_men_n733_));
  NA4        u0705(.A(men_men_n223_), .B(men_men_n146_), .C(men_men_n45_), .D(h), .Y(men_men_n734_));
  AN2        u0706(.A(l), .B(k), .Y(men_men_n735_));
  NA4        u0707(.A(men_men_n735_), .B(men_men_n112_), .C(men_men_n75_), .D(men_men_n221_), .Y(men_men_n736_));
  OAI210     u0708(.A0(men_men_n734_), .A1(g), .B0(men_men_n736_), .Y(men_men_n737_));
  NA2        u0709(.A(men_men_n737_), .B(men_men_n733_), .Y(men_men_n738_));
  NA4        u0710(.A(men_men_n738_), .B(men_men_n732_), .C(men_men_n727_), .D(men_men_n364_), .Y(men_men_n739_));
  AN2        u0711(.A(men_men_n561_), .B(men_men_n98_), .Y(men_men_n740_));
  NO4        u0712(.A(men_men_n180_), .B(men_men_n408_), .C(men_men_n116_), .D(g), .Y(men_men_n741_));
  AOI210     u0713(.A0(men_men_n741_), .A1(men_men_n731_), .B0(men_men_n545_), .Y(men_men_n742_));
  NO2        u0714(.A(men_men_n38_), .B(men_men_n220_), .Y(men_men_n743_));
  AOI220     u0715(.A0(men_men_n651_), .A1(men_men_n361_), .B0(men_men_n743_), .B1(men_men_n593_), .Y(men_men_n744_));
  NAi31      u0716(.An(men_men_n740_), .B(men_men_n744_), .C(men_men_n742_), .Y(men_men_n745_));
  NO2        u0717(.A(men_men_n564_), .B(men_men_n35_), .Y(men_men_n746_));
  OAI210     u0718(.A0(men_men_n581_), .A1(men_men_n47_), .B0(men_men_n140_), .Y(men_men_n747_));
  NO2        u0719(.A(men_men_n505_), .B(men_men_n137_), .Y(men_men_n748_));
  AOI210     u0720(.A0(men_men_n748_), .A1(men_men_n747_), .B0(men_men_n746_), .Y(men_men_n749_));
  NO3        u0721(.A(men_men_n328_), .B(men_men_n136_), .C(men_men_n41_), .Y(men_men_n750_));
  NAi21      u0722(.An(men_men_n750_), .B(men_men_n736_), .Y(men_men_n751_));
  AOI220     u0723(.A0(men_men_n1596_), .A1(men_men_n418_), .B0(men_men_n751_), .B1(men_men_n78_), .Y(men_men_n752_));
  OAI210     u0724(.A0(men_men_n749_), .A1(men_men_n89_), .B0(men_men_n752_), .Y(men_men_n753_));
  NA2        u0725(.A(men_men_n376_), .B(men_men_n43_), .Y(men_men_n754_));
  NA2        u0726(.A(men_men_n735_), .B(men_men_n228_), .Y(men_men_n755_));
  NO2        u0727(.A(men_men_n755_), .B(men_men_n340_), .Y(men_men_n756_));
  AOI210     u0728(.A0(men_men_n756_), .A1(men_men_n712_), .B0(men_men_n512_), .Y(men_men_n757_));
  NA3        u0729(.A(m), .B(l), .C(k), .Y(men_men_n758_));
  AOI210     u0730(.A0(men_men_n692_), .A1(men_men_n690_), .B0(men_men_n758_), .Y(men_men_n759_));
  NO2        u0731(.A(men_men_n563_), .B(men_men_n278_), .Y(men_men_n760_));
  NOi21      u0732(.An(men_men_n760_), .B(men_men_n557_), .Y(men_men_n761_));
  NA4        u0733(.A(men_men_n117_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n762_));
  NA3        u0734(.A(men_men_n125_), .B(men_men_n427_), .C(i), .Y(men_men_n763_));
  NO2        u0735(.A(men_men_n763_), .B(men_men_n762_), .Y(men_men_n764_));
  NO3        u0736(.A(men_men_n764_), .B(men_men_n761_), .C(men_men_n759_), .Y(men_men_n765_));
  NA3        u0737(.A(men_men_n765_), .B(men_men_n757_), .C(men_men_n754_), .Y(men_men_n766_));
  NO4        u0738(.A(men_men_n766_), .B(men_men_n753_), .C(men_men_n745_), .D(men_men_n739_), .Y(men_men_n767_));
  NA2        u0739(.A(men_men_n651_), .B(men_men_n409_), .Y(men_men_n768_));
  NOi31      u0740(.An(g), .B(h), .C(f), .Y(men_men_n769_));
  NA2        u0741(.A(men_men_n667_), .B(men_men_n769_), .Y(men_men_n770_));
  AO210      u0742(.A0(men_men_n770_), .A1(men_men_n620_), .B0(men_men_n566_), .Y(men_men_n771_));
  NO3        u0743(.A(men_men_n412_), .B(men_men_n551_), .C(h), .Y(men_men_n772_));
  AOI210     u0744(.A0(men_men_n772_), .A1(men_men_n117_), .B0(men_men_n524_), .Y(men_men_n773_));
  NA4        u0745(.A(men_men_n773_), .B(men_men_n771_), .C(men_men_n768_), .D(men_men_n257_), .Y(men_men_n774_));
  NA2        u0746(.A(men_men_n735_), .B(men_men_n75_), .Y(men_men_n775_));
  NO4        u0747(.A(men_men_n1599_), .B(men_men_n180_), .C(n), .D(i), .Y(men_men_n776_));
  NOi21      u0748(.An(h), .B(j), .Y(men_men_n777_));
  NA2        u0749(.A(men_men_n777_), .B(f), .Y(men_men_n778_));
  NO2        u0750(.A(men_men_n778_), .B(men_men_n251_), .Y(men_men_n779_));
  NO2        u0751(.A(men_men_n779_), .B(men_men_n776_), .Y(men_men_n780_));
  OAI220     u0752(.A0(men_men_n780_), .A1(men_men_n775_), .B0(men_men_n622_), .B1(men_men_n62_), .Y(men_men_n781_));
  AOI210     u0753(.A0(men_men_n774_), .A1(l), .B0(men_men_n781_), .Y(men_men_n782_));
  NO2        u0754(.A(j), .B(i), .Y(men_men_n783_));
  NA3        u0755(.A(men_men_n783_), .B(men_men_n82_), .C(l), .Y(men_men_n784_));
  NA2        u0756(.A(men_men_n783_), .B(men_men_n33_), .Y(men_men_n785_));
  NA2        u0757(.A(men_men_n437_), .B(men_men_n125_), .Y(men_men_n786_));
  OA220      u0758(.A0(men_men_n786_), .A1(men_men_n785_), .B0(men_men_n784_), .B1(men_men_n618_), .Y(men_men_n787_));
  NO3        u0759(.A(men_men_n157_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n788_));
  NO3        u0760(.A(men_men_n570_), .B(men_men_n156_), .C(men_men_n75_), .Y(men_men_n789_));
  NO3        u0761(.A(men_men_n505_), .B(men_men_n456_), .C(j), .Y(men_men_n790_));
  OAI210     u0762(.A0(men_men_n789_), .A1(men_men_n788_), .B0(men_men_n790_), .Y(men_men_n791_));
  OAI210     u0763(.A0(men_men_n770_), .A1(men_men_n62_), .B0(men_men_n791_), .Y(men_men_n792_));
  NA2        u0764(.A(k), .B(j), .Y(men_men_n793_));
  NO3        u0765(.A(men_men_n307_), .B(men_men_n793_), .C(men_men_n40_), .Y(men_men_n794_));
  AOI210     u0766(.A0(men_men_n556_), .A1(n), .B0(men_men_n580_), .Y(men_men_n795_));
  NA2        u0767(.A(men_men_n795_), .B(men_men_n582_), .Y(men_men_n796_));
  AN3        u0768(.A(men_men_n796_), .B(men_men_n794_), .C(men_men_n101_), .Y(men_men_n797_));
  NO3        u0769(.A(men_men_n180_), .B(men_men_n408_), .C(men_men_n116_), .Y(men_men_n798_));
  AOI220     u0770(.A0(men_men_n798_), .A1(men_men_n252_), .B0(c), .B1(men_men_n318_), .Y(men_men_n799_));
  NAi31      u0771(.An(men_men_n638_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n800_));
  NA2        u0772(.A(men_men_n800_), .B(men_men_n799_), .Y(men_men_n801_));
  NO2        u0773(.A(men_men_n307_), .B(men_men_n141_), .Y(men_men_n802_));
  AOI220     u0774(.A0(men_men_n802_), .A1(men_men_n651_), .B0(men_men_n750_), .B1(men_men_n733_), .Y(men_men_n803_));
  NO2        u0775(.A(men_men_n758_), .B(men_men_n93_), .Y(men_men_n804_));
  NA2        u0776(.A(men_men_n804_), .B(men_men_n617_), .Y(men_men_n805_));
  NO2        u0777(.A(men_men_n619_), .B(men_men_n121_), .Y(men_men_n806_));
  OAI210     u0778(.A0(men_men_n806_), .A1(men_men_n790_), .B0(men_men_n708_), .Y(men_men_n807_));
  NA3        u0779(.A(men_men_n807_), .B(men_men_n805_), .C(men_men_n803_), .Y(men_men_n808_));
  OR4        u0780(.A(men_men_n808_), .B(men_men_n801_), .C(men_men_n797_), .D(men_men_n792_), .Y(men_men_n809_));
  NA3        u0781(.A(men_men_n795_), .B(men_men_n582_), .C(men_men_n581_), .Y(men_men_n810_));
  NA4        u0782(.A(men_men_n810_), .B(men_men_n223_), .C(men_men_n469_), .D(men_men_n34_), .Y(men_men_n811_));
  NO4        u0783(.A(men_men_n505_), .B(men_men_n451_), .C(j), .D(f), .Y(men_men_n812_));
  OAI220     u0784(.A0(men_men_n734_), .A1(men_men_n726_), .B0(men_men_n345_), .B1(men_men_n38_), .Y(men_men_n813_));
  AOI210     u0785(.A0(men_men_n812_), .A1(men_men_n263_), .B0(men_men_n813_), .Y(men_men_n814_));
  NA3        u0786(.A(men_men_n573_), .B(men_men_n300_), .C(h), .Y(men_men_n815_));
  NOi21      u0787(.An(men_men_n708_), .B(men_men_n815_), .Y(men_men_n816_));
  NO2        u0788(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n817_));
  OAI220     u0789(.A0(men_men_n815_), .A1(men_men_n636_), .B0(men_men_n784_), .B1(men_men_n700_), .Y(men_men_n818_));
  AOI210     u0790(.A0(men_men_n817_), .A1(men_men_n673_), .B0(men_men_n818_), .Y(men_men_n819_));
  NAi41      u0791(.An(men_men_n816_), .B(men_men_n819_), .C(men_men_n814_), .D(men_men_n811_), .Y(men_men_n820_));
  OR2        u0792(.A(men_men_n804_), .B(men_men_n98_), .Y(men_men_n821_));
  AOI220     u0793(.A0(men_men_n821_), .A1(men_men_n242_), .B0(men_men_n790_), .B1(men_men_n665_), .Y(men_men_n822_));
  NO2        u0794(.A(men_men_n691_), .B(men_men_n75_), .Y(men_men_n823_));
  AOI210     u0795(.A0(men_men_n812_), .A1(men_men_n823_), .B0(men_men_n349_), .Y(men_men_n824_));
  OAI210     u0796(.A0(men_men_n758_), .A1(men_men_n689_), .B0(men_men_n544_), .Y(men_men_n825_));
  NA3        u0797(.A(men_men_n255_), .B(men_men_n59_), .C(b), .Y(men_men_n826_));
  AOI220     u0798(.A0(men_men_n635_), .A1(men_men_n29_), .B0(men_men_n483_), .B1(men_men_n86_), .Y(men_men_n827_));
  NA2        u0799(.A(men_men_n827_), .B(men_men_n826_), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n815_), .B(men_men_n511_), .Y(men_men_n829_));
  AOI210     u0801(.A0(men_men_n828_), .A1(men_men_n825_), .B0(men_men_n829_), .Y(men_men_n830_));
  NA3        u0802(.A(men_men_n830_), .B(men_men_n824_), .C(men_men_n822_), .Y(men_men_n831_));
  NOi41      u0803(.An(men_men_n787_), .B(men_men_n831_), .C(men_men_n820_), .D(men_men_n809_), .Y(men_men_n832_));
  OR3        u0804(.A(men_men_n734_), .B(men_men_n237_), .C(g), .Y(men_men_n833_));
  NO3        u0805(.A(men_men_n355_), .B(men_men_n309_), .C(men_men_n116_), .Y(men_men_n834_));
  NA2        u0806(.A(men_men_n834_), .B(men_men_n796_), .Y(men_men_n835_));
  NA2        u0807(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n836_));
  NO3        u0808(.A(men_men_n836_), .B(men_men_n785_), .C(men_men_n284_), .Y(men_men_n837_));
  NO3        u0809(.A(men_men_n551_), .B(men_men_n96_), .C(h), .Y(men_men_n838_));
  AOI210     u0810(.A0(men_men_n838_), .A1(men_men_n729_), .B0(men_men_n837_), .Y(men_men_n839_));
  NA4        u0811(.A(men_men_n839_), .B(men_men_n835_), .C(men_men_n833_), .D(men_men_n420_), .Y(men_men_n840_));
  OR2        u0812(.A(men_men_n689_), .B(men_men_n94_), .Y(men_men_n841_));
  NOi31      u0813(.An(b), .B(d), .C(a), .Y(men_men_n842_));
  NO2        u0814(.A(men_men_n842_), .B(men_men_n633_), .Y(men_men_n843_));
  NO2        u0815(.A(men_men_n843_), .B(n), .Y(men_men_n844_));
  NOi21      u0816(.An(men_men_n827_), .B(men_men_n844_), .Y(men_men_n845_));
  OAI220     u0817(.A0(men_men_n845_), .A1(men_men_n841_), .B0(men_men_n815_), .B1(men_men_n634_), .Y(men_men_n846_));
  INV        u0818(.A(men_men_n581_), .Y(men_men_n847_));
  NO3        u0819(.A(men_men_n650_), .B(men_men_n340_), .C(men_men_n121_), .Y(men_men_n848_));
  NOi21      u0820(.An(men_men_n848_), .B(men_men_n167_), .Y(men_men_n849_));
  AOI210     u0821(.A0(men_men_n834_), .A1(men_men_n847_), .B0(men_men_n849_), .Y(men_men_n850_));
  OAI210     u0822(.A0(men_men_n734_), .A1(men_men_n410_), .B0(men_men_n850_), .Y(men_men_n851_));
  NA2        u0823(.A(men_men_n802_), .B(men_men_n696_), .Y(men_men_n852_));
  NO2        u0824(.A(men_men_n335_), .B(men_men_n241_), .Y(men_men_n853_));
  OAI210     u0825(.A0(men_men_n98_), .A1(men_men_n95_), .B0(men_men_n853_), .Y(men_men_n854_));
  NA2        u0826(.A(men_men_n125_), .B(men_men_n86_), .Y(men_men_n855_));
  AOI210     u0827(.A0(men_men_n441_), .A1(men_men_n433_), .B0(men_men_n855_), .Y(men_men_n856_));
  NAi21      u0828(.An(men_men_n856_), .B(men_men_n854_), .Y(men_men_n857_));
  NA2        u0829(.A(men_men_n756_), .B(men_men_n34_), .Y(men_men_n858_));
  NAi21      u0830(.An(men_men_n762_), .B(men_men_n452_), .Y(men_men_n859_));
  NA2        u0831(.A(men_men_n741_), .B(men_men_n363_), .Y(men_men_n860_));
  OAI210     u0832(.A0(men_men_n625_), .A1(men_men_n624_), .B0(men_men_n377_), .Y(men_men_n861_));
  AN3        u0833(.A(men_men_n861_), .B(men_men_n860_), .C(men_men_n859_), .Y(men_men_n862_));
  NAi41      u0834(.An(men_men_n857_), .B(men_men_n862_), .C(men_men_n858_), .D(men_men_n852_), .Y(men_men_n863_));
  NO4        u0835(.A(men_men_n863_), .B(men_men_n851_), .C(men_men_n846_), .D(men_men_n840_), .Y(men_men_n864_));
  NA4        u0836(.A(men_men_n864_), .B(men_men_n832_), .C(men_men_n782_), .D(men_men_n767_), .Y(men09));
  INV        u0837(.A(men_men_n126_), .Y(men_men_n866_));
  NA2        u0838(.A(f), .B(e), .Y(men_men_n867_));
  NO2        u0839(.A(men_men_n233_), .B(men_men_n116_), .Y(men_men_n868_));
  NA2        u0840(.A(men_men_n868_), .B(g), .Y(men_men_n869_));
  NA4        u0841(.A(men_men_n321_), .B(men_men_n492_), .C(men_men_n266_), .D(men_men_n123_), .Y(men_men_n870_));
  AOI210     u0842(.A0(men_men_n870_), .A1(g), .B0(men_men_n489_), .Y(men_men_n871_));
  AOI210     u0843(.A0(men_men_n871_), .A1(men_men_n869_), .B0(men_men_n867_), .Y(men_men_n872_));
  NA2        u0844(.A(men_men_n462_), .B(e), .Y(men_men_n873_));
  NO2        u0845(.A(men_men_n873_), .B(men_men_n535_), .Y(men_men_n874_));
  AOI210     u0846(.A0(men_men_n872_), .A1(men_men_n866_), .B0(men_men_n874_), .Y(men_men_n875_));
  NO2        u0847(.A(men_men_n210_), .B(men_men_n220_), .Y(men_men_n876_));
  NA3        u0848(.A(m), .B(l), .C(i), .Y(men_men_n877_));
  OAI220     u0849(.A0(men_men_n619_), .A1(men_men_n877_), .B0(men_men_n368_), .B1(men_men_n552_), .Y(men_men_n878_));
  NA4        u0850(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n879_));
  NAi31      u0851(.An(men_men_n878_), .B(men_men_n879_), .C(men_men_n457_), .Y(men_men_n880_));
  OR2        u0852(.A(men_men_n880_), .B(men_men_n876_), .Y(men_men_n881_));
  NA3        u0853(.A(men_men_n841_), .B(men_men_n595_), .C(men_men_n544_), .Y(men_men_n882_));
  OA210      u0854(.A0(men_men_n882_), .A1(men_men_n881_), .B0(men_men_n844_), .Y(men_men_n883_));
  INV        u0855(.A(men_men_n352_), .Y(men_men_n884_));
  NO2        u0856(.A(men_men_n132_), .B(men_men_n130_), .Y(men_men_n885_));
  NOi31      u0857(.An(k), .B(m), .C(l), .Y(men_men_n886_));
  NO2        u0858(.A(men_men_n354_), .B(men_men_n886_), .Y(men_men_n887_));
  AOI210     u0859(.A0(men_men_n887_), .A1(men_men_n885_), .B0(men_men_n628_), .Y(men_men_n888_));
  NA2        u0860(.A(men_men_n826_), .B(men_men_n345_), .Y(men_men_n889_));
  NA2        u0861(.A(men_men_n356_), .B(men_men_n358_), .Y(men_men_n890_));
  OAI210     u0862(.A0(men_men_n210_), .A1(men_men_n220_), .B0(men_men_n890_), .Y(men_men_n891_));
  AOI220     u0863(.A0(men_men_n891_), .A1(men_men_n889_), .B0(men_men_n888_), .B1(men_men_n884_), .Y(men_men_n892_));
  NA3        u0864(.A(men_men_n1597_), .B(men_men_n196_), .C(men_men_n31_), .Y(men_men_n893_));
  NA4        u0865(.A(men_men_n893_), .B(men_men_n892_), .C(men_men_n652_), .D(men_men_n84_), .Y(men_men_n894_));
  NO2        u0866(.A(men_men_n615_), .B(men_men_n520_), .Y(men_men_n895_));
  NA2        u0867(.A(men_men_n895_), .B(men_men_n196_), .Y(men_men_n896_));
  NOi21      u0868(.An(f), .B(d), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n897_), .B(m), .Y(men_men_n898_));
  NO2        u0870(.A(men_men_n898_), .B(men_men_n52_), .Y(men_men_n899_));
  NOi32      u0871(.An(g), .Bn(f), .C(d), .Y(men_men_n900_));
  NA4        u0872(.A(men_men_n900_), .B(men_men_n635_), .C(men_men_n29_), .D(m), .Y(men_men_n901_));
  NOi21      u0873(.An(men_men_n322_), .B(men_men_n901_), .Y(men_men_n902_));
  AOI210     u0874(.A0(men_men_n899_), .A1(men_men_n571_), .B0(men_men_n902_), .Y(men_men_n903_));
  NA3        u0875(.A(men_men_n321_), .B(men_men_n266_), .C(men_men_n123_), .Y(men_men_n904_));
  AN2        u0876(.A(f), .B(d), .Y(men_men_n905_));
  NA3        u0877(.A(men_men_n497_), .B(men_men_n905_), .C(men_men_n86_), .Y(men_men_n906_));
  NO3        u0878(.A(men_men_n906_), .B(men_men_n75_), .C(men_men_n221_), .Y(men_men_n907_));
  NO2        u0879(.A(men_men_n293_), .B(men_men_n56_), .Y(men_men_n908_));
  NA2        u0880(.A(men_men_n904_), .B(men_men_n907_), .Y(men_men_n909_));
  NAi41      u0881(.An(men_men_n510_), .B(men_men_n909_), .C(men_men_n903_), .D(men_men_n896_), .Y(men_men_n910_));
  NO4        u0882(.A(men_men_n650_), .B(men_men_n137_), .C(men_men_n340_), .D(men_men_n158_), .Y(men_men_n911_));
  NO2        u0883(.A(men_men_n683_), .B(men_men_n340_), .Y(men_men_n912_));
  AN2        u0884(.A(men_men_n912_), .B(men_men_n712_), .Y(men_men_n913_));
  NO3        u0885(.A(men_men_n913_), .B(men_men_n911_), .C(men_men_n239_), .Y(men_men_n914_));
  NA2        u0886(.A(men_men_n633_), .B(men_men_n86_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n890_), .B(men_men_n915_), .Y(men_men_n916_));
  NA3        u0888(.A(men_men_n166_), .B(men_men_n112_), .C(men_men_n111_), .Y(men_men_n917_));
  OAI220     u0889(.A0(men_men_n906_), .A1(men_men_n446_), .B0(men_men_n352_), .B1(men_men_n917_), .Y(men_men_n918_));
  NOi41      u0890(.An(men_men_n231_), .B(men_men_n918_), .C(men_men_n916_), .D(men_men_n316_), .Y(men_men_n919_));
  NA2        u0891(.A(c), .B(men_men_n120_), .Y(men_men_n920_));
  NO2        u0892(.A(men_men_n920_), .B(men_men_n424_), .Y(men_men_n921_));
  NA3        u0893(.A(men_men_n921_), .B(men_men_n533_), .C(f), .Y(men_men_n922_));
  OR2        u0894(.A(men_men_n689_), .B(men_men_n567_), .Y(men_men_n923_));
  INV        u0895(.A(men_men_n923_), .Y(men_men_n924_));
  NA2        u0896(.A(men_men_n843_), .B(men_men_n115_), .Y(men_men_n925_));
  NA2        u0897(.A(men_men_n925_), .B(men_men_n924_), .Y(men_men_n926_));
  NA4        u0898(.A(men_men_n926_), .B(men_men_n922_), .C(men_men_n919_), .D(men_men_n914_), .Y(men_men_n927_));
  NO4        u0899(.A(men_men_n927_), .B(men_men_n910_), .C(men_men_n894_), .D(men_men_n883_), .Y(men_men_n928_));
  OR2        u0900(.A(men_men_n906_), .B(men_men_n75_), .Y(men_men_n929_));
  NA2        u0901(.A(men_men_n116_), .B(j), .Y(men_men_n930_));
  NA2        u0902(.A(men_men_n868_), .B(g), .Y(men_men_n931_));
  AOI210     u0903(.A0(men_men_n931_), .A1(men_men_n301_), .B0(men_men_n929_), .Y(men_men_n932_));
  NO2        u0904(.A(men_men_n345_), .B(men_men_n879_), .Y(men_men_n933_));
  NO2        u0905(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n934_));
  NA2        u0906(.A(men_men_n314_), .B(men_men_n934_), .Y(men_men_n935_));
  NO2        u0907(.A(men_men_n446_), .B(men_men_n867_), .Y(men_men_n936_));
  NA2        u0908(.A(men_men_n936_), .B(men_men_n587_), .Y(men_men_n937_));
  NA2        u0909(.A(men_men_n937_), .B(men_men_n935_), .Y(men_men_n938_));
  NA2        u0910(.A(e), .B(d), .Y(men_men_n939_));
  NA2        u0911(.A(men_men_n651_), .B(men_men_n361_), .Y(men_men_n940_));
  NA2        u0912(.A(men_men_n293_), .B(men_men_n172_), .Y(men_men_n941_));
  NA2        u0913(.A(men_men_n907_), .B(men_men_n941_), .Y(men_men_n942_));
  NA3        u0914(.A(men_men_n175_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n943_));
  NA3        u0915(.A(men_men_n943_), .B(men_men_n942_), .C(men_men_n940_), .Y(men_men_n944_));
  NO4        u0916(.A(men_men_n944_), .B(men_men_n938_), .C(men_men_n933_), .D(men_men_n932_), .Y(men_men_n945_));
  NA2        u0917(.A(men_men_n884_), .B(men_men_n31_), .Y(men_men_n946_));
  AO210      u0918(.A0(men_men_n946_), .A1(men_men_n726_), .B0(men_men_n224_), .Y(men_men_n947_));
  OAI220     u0919(.A0(men_men_n650_), .A1(men_men_n61_), .B0(men_men_n309_), .B1(j), .Y(men_men_n948_));
  AOI220     u0920(.A0(men_men_n948_), .A1(men_men_n912_), .B0(men_men_n643_), .B1(men_men_n649_), .Y(men_men_n949_));
  OAI210     u0921(.A0(men_men_n873_), .A1(d), .B0(men_men_n949_), .Y(men_men_n950_));
  OAI210     u0922(.A0(men_men_n868_), .A1(men_men_n941_), .B0(men_men_n900_), .Y(men_men_n951_));
  NO2        u0923(.A(men_men_n951_), .B(men_men_n636_), .Y(men_men_n952_));
  AOI210     u0924(.A0(men_men_n122_), .A1(men_men_n121_), .B0(men_men_n265_), .Y(men_men_n953_));
  NO2        u0925(.A(men_men_n953_), .B(men_men_n901_), .Y(men_men_n954_));
  AO210      u0926(.A0(men_men_n889_), .A1(men_men_n878_), .B0(men_men_n954_), .Y(men_men_n955_));
  NOi31      u0927(.An(men_men_n571_), .B(men_men_n898_), .C(men_men_n301_), .Y(men_men_n956_));
  NO4        u0928(.A(men_men_n956_), .B(men_men_n955_), .C(men_men_n952_), .D(men_men_n950_), .Y(men_men_n957_));
  NA2        u0929(.A(men_men_n475_), .B(e), .Y(men_men_n958_));
  NO2        u0930(.A(men_men_n456_), .B(men_men_n71_), .Y(men_men_n959_));
  OAI210     u0931(.A0(men_men_n882_), .A1(men_men_n959_), .B0(men_men_n729_), .Y(men_men_n960_));
  AN4        u0932(.A(men_men_n960_), .B(men_men_n958_), .C(men_men_n957_), .D(men_men_n947_), .Y(men_men_n961_));
  NA4        u0933(.A(men_men_n961_), .B(men_men_n945_), .C(men_men_n928_), .D(men_men_n875_), .Y(men12));
  NO2        u0934(.A(men_men_n472_), .B(c), .Y(men_men_n963_));
  NO4        u0935(.A(men_men_n461_), .B(men_men_n258_), .C(men_men_n611_), .D(men_men_n221_), .Y(men_men_n964_));
  NA2        u0936(.A(men_men_n964_), .B(men_men_n963_), .Y(men_men_n965_));
  NA2        u0937(.A(men_men_n571_), .B(men_men_n959_), .Y(men_men_n966_));
  NO2        u0938(.A(men_men_n472_), .B(men_men_n120_), .Y(men_men_n967_));
  NO2        u0939(.A(men_men_n885_), .B(men_men_n368_), .Y(men_men_n968_));
  NO2        u0940(.A(men_men_n689_), .B(men_men_n394_), .Y(men_men_n969_));
  AOI220     u0941(.A0(men_men_n969_), .A1(men_men_n569_), .B0(men_men_n968_), .B1(men_men_n967_), .Y(men_men_n970_));
  NA4        u0942(.A(men_men_n970_), .B(men_men_n966_), .C(men_men_n965_), .D(men_men_n460_), .Y(men_men_n971_));
  AOI210     u0943(.A0(men_men_n238_), .A1(men_men_n351_), .B0(men_men_n207_), .Y(men_men_n972_));
  AOI210     u0944(.A0(men_men_n348_), .A1(men_men_n406_), .B0(men_men_n221_), .Y(men_men_n973_));
  OAI210     u0945(.A0(men_men_n973_), .A1(men_men_n972_), .B0(men_men_n419_), .Y(men_men_n974_));
  NO2        u0946(.A(men_men_n670_), .B(men_men_n268_), .Y(men_men_n975_));
  NO2        u0947(.A(men_men_n619_), .B(men_men_n877_), .Y(men_men_n976_));
  AOI220     u0948(.A0(men_men_n976_), .A1(men_men_n593_), .B0(men_men_n853_), .B1(men_men_n975_), .Y(men_men_n977_));
  NO2        u0949(.A(men_men_n157_), .B(men_men_n241_), .Y(men_men_n978_));
  NA3        u0950(.A(men_men_n978_), .B(men_men_n244_), .C(i), .Y(men_men_n979_));
  NA3        u0951(.A(men_men_n979_), .B(men_men_n977_), .C(men_men_n974_), .Y(men_men_n980_));
  BUFFER     u0952(.A(men_men_n967_), .Y(men_men_n981_));
  NA2        u0953(.A(men_men_n981_), .B(men_men_n369_), .Y(men_men_n982_));
  NO3        u0954(.A(men_men_n137_), .B(men_men_n158_), .C(men_men_n221_), .Y(men_men_n983_));
  NA2        u0955(.A(men_men_n983_), .B(men_men_n556_), .Y(men_men_n984_));
  NA4        u0956(.A(men_men_n462_), .B(men_men_n454_), .C(men_men_n187_), .D(g), .Y(men_men_n985_));
  NA3        u0957(.A(men_men_n985_), .B(men_men_n984_), .C(men_men_n982_), .Y(men_men_n986_));
  NO3        u0958(.A(men_men_n694_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n987_));
  NO4        u0959(.A(men_men_n987_), .B(men_men_n986_), .C(men_men_n980_), .D(men_men_n971_), .Y(men_men_n988_));
  NO2        u0960(.A(men_men_n384_), .B(men_men_n383_), .Y(men_men_n989_));
  NA2        u0961(.A(men_men_n616_), .B(men_men_n73_), .Y(men_men_n990_));
  NA2        u0962(.A(men_men_n581_), .B(men_men_n151_), .Y(men_men_n991_));
  NOi21      u0963(.An(men_men_n34_), .B(men_men_n683_), .Y(men_men_n992_));
  AOI220     u0964(.A0(men_men_n992_), .A1(men_men_n991_), .B0(men_men_n990_), .B1(men_men_n989_), .Y(men_men_n993_));
  OAI210     u0965(.A0(men_men_n256_), .A1(men_men_n45_), .B0(men_men_n993_), .Y(men_men_n994_));
  NA2        u0966(.A(men_men_n452_), .B(men_men_n270_), .Y(men_men_n995_));
  NO3        u0967(.A(men_men_n855_), .B(men_men_n91_), .C(men_men_n424_), .Y(men_men_n996_));
  NAi31      u0968(.An(men_men_n996_), .B(men_men_n995_), .C(men_men_n332_), .Y(men_men_n997_));
  NO2        u0969(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n998_));
  NO2        u0970(.A(men_men_n527_), .B(men_men_n309_), .Y(men_men_n999_));
  NO2        u0971(.A(men_men_n999_), .B(men_men_n380_), .Y(men_men_n1000_));
  NO2        u0972(.A(men_men_n1000_), .B(men_men_n151_), .Y(men_men_n1001_));
  NA2        u0973(.A(men_men_n661_), .B(men_men_n377_), .Y(men_men_n1002_));
  OAI210     u0974(.A0(men_men_n763_), .A1(men_men_n1002_), .B0(men_men_n381_), .Y(men_men_n1003_));
  NO4        u0975(.A(men_men_n1003_), .B(men_men_n1001_), .C(men_men_n997_), .D(men_men_n994_), .Y(men_men_n1004_));
  NA2        u0976(.A(men_men_n361_), .B(g), .Y(men_men_n1005_));
  NA2        u0977(.A(men_men_n169_), .B(i), .Y(men_men_n1006_));
  NA2        u0978(.A(men_men_n46_), .B(i), .Y(men_men_n1007_));
  OAI220     u0979(.A0(men_men_n1007_), .A1(men_men_n206_), .B0(men_men_n1006_), .B1(men_men_n94_), .Y(men_men_n1008_));
  AOI210     u0980(.A0(men_men_n435_), .A1(men_men_n37_), .B0(men_men_n1008_), .Y(men_men_n1009_));
  NO2        u0981(.A(men_men_n151_), .B(men_men_n86_), .Y(men_men_n1010_));
  OR2        u0982(.A(men_men_n1010_), .B(men_men_n580_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n581_), .B(men_men_n398_), .Y(men_men_n1012_));
  NO2        u0984(.A(men_men_n1012_), .B(men_men_n1011_), .Y(men_men_n1013_));
  OAI220     u0985(.A0(men_men_n1013_), .A1(men_men_n1005_), .B0(men_men_n1009_), .B1(men_men_n345_), .Y(men_men_n1014_));
  NO2        u0986(.A(men_men_n689_), .B(men_men_n520_), .Y(men_men_n1015_));
  NA3        u0987(.A(men_men_n356_), .B(men_men_n656_), .C(i), .Y(men_men_n1016_));
  OAI210     u0988(.A0(men_men_n456_), .A1(men_men_n321_), .B0(men_men_n1016_), .Y(men_men_n1017_));
  OAI220     u0989(.A0(men_men_n1017_), .A1(men_men_n1015_), .B0(men_men_n708_), .B1(men_men_n789_), .Y(men_men_n1018_));
  NA2        u0990(.A(men_men_n637_), .B(men_men_n117_), .Y(men_men_n1019_));
  OR3        u0991(.A(men_men_n321_), .B(men_men_n451_), .C(f), .Y(men_men_n1020_));
  NA3        u0992(.A(men_men_n656_), .B(men_men_n82_), .C(i), .Y(men_men_n1021_));
  OA220      u0993(.A0(men_men_n1021_), .A1(men_men_n1019_), .B0(men_men_n1020_), .B1(men_men_n618_), .Y(men_men_n1022_));
  NA3        u0994(.A(men_men_n337_), .B(men_men_n122_), .C(g), .Y(men_men_n1023_));
  AOI210     u0995(.A0(men_men_n705_), .A1(men_men_n1023_), .B0(m), .Y(men_men_n1024_));
  NA2        u0996(.A(men_men_n968_), .B(men_men_n336_), .Y(men_men_n1025_));
  NA2        u0997(.A(men_men_n717_), .B(men_men_n915_), .Y(men_men_n1026_));
  NA2        u0998(.A(men_men_n879_), .B(men_men_n457_), .Y(men_men_n1027_));
  NA2        u0999(.A(men_men_n229_), .B(men_men_n79_), .Y(men_men_n1028_));
  NA3        u1000(.A(men_men_n1028_), .B(men_men_n1021_), .C(men_men_n1020_), .Y(men_men_n1029_));
  AOI220     u1001(.A0(men_men_n1029_), .A1(men_men_n263_), .B0(men_men_n1027_), .B1(men_men_n1026_), .Y(men_men_n1030_));
  NA4        u1002(.A(men_men_n1030_), .B(men_men_n1025_), .C(men_men_n1022_), .D(men_men_n1018_), .Y(men_men_n1031_));
  NO2        u1003(.A(men_men_n394_), .B(men_men_n93_), .Y(men_men_n1032_));
  OAI210     u1004(.A0(men_men_n1032_), .A1(men_men_n975_), .B0(men_men_n242_), .Y(men_men_n1033_));
  NA2        u1005(.A(men_men_n693_), .B(men_men_n90_), .Y(men_men_n1034_));
  NO2        u1006(.A(men_men_n478_), .B(men_men_n221_), .Y(men_men_n1035_));
  NA2        u1007(.A(men_men_n981_), .B(men_men_n225_), .Y(men_men_n1036_));
  AOI220     u1008(.A0(men_men_n969_), .A1(men_men_n978_), .B0(men_men_n617_), .B1(men_men_n92_), .Y(men_men_n1037_));
  NA4        u1009(.A(men_men_n1037_), .B(men_men_n1036_), .C(men_men_n1034_), .D(men_men_n1033_), .Y(men_men_n1038_));
  OAI210     u1010(.A0(men_men_n1027_), .A1(men_men_n976_), .B0(men_men_n569_), .Y(men_men_n1039_));
  AOI210     u1011(.A0(men_men_n436_), .A1(men_men_n428_), .B0(men_men_n855_), .Y(men_men_n1040_));
  OAI210     u1012(.A0(men_men_n384_), .A1(men_men_n383_), .B0(men_men_n113_), .Y(men_men_n1041_));
  AOI210     u1013(.A0(men_men_n1041_), .A1(men_men_n561_), .B0(men_men_n1040_), .Y(men_men_n1042_));
  NA2        u1014(.A(men_men_n1024_), .B(men_men_n967_), .Y(men_men_n1043_));
  NO3        u1015(.A(men_men_n930_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1044_));
  AOI220     u1016(.A0(men_men_n1044_), .A1(men_men_n654_), .B0(men_men_n675_), .B1(men_men_n556_), .Y(men_men_n1045_));
  NA4        u1017(.A(men_men_n1045_), .B(men_men_n1043_), .C(men_men_n1042_), .D(men_men_n1039_), .Y(men_men_n1046_));
  NO4        u1018(.A(men_men_n1046_), .B(men_men_n1038_), .C(men_men_n1031_), .D(men_men_n1014_), .Y(men_men_n1047_));
  NAi31      u1019(.An(men_men_n147_), .B(men_men_n437_), .C(n), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n130_), .B(men_men_n354_), .C(men_men_n886_), .Y(men_men_n1049_));
  NO2        u1021(.A(men_men_n1049_), .B(men_men_n1048_), .Y(men_men_n1050_));
  NO2        u1022(.A(men_men_n278_), .B(men_men_n147_), .Y(men_men_n1051_));
  AOI210     u1023(.A0(men_men_n1051_), .A1(men_men_n521_), .B0(men_men_n1050_), .Y(men_men_n1052_));
  NA2        u1024(.A(men_men_n513_), .B(i), .Y(men_men_n1053_));
  NA2        u1025(.A(men_men_n1053_), .B(men_men_n1052_), .Y(men_men_n1054_));
  NO2        u1026(.A(men_men_n318_), .B(men_men_n462_), .Y(men_men_n1055_));
  NOi31      u1027(.An(c), .B(men_men_n1055_), .C(men_men_n221_), .Y(men_men_n1056_));
  NAi21      u1028(.An(men_men_n581_), .B(men_men_n1035_), .Y(men_men_n1057_));
  NA2        u1029(.A(men_men_n455_), .B(men_men_n915_), .Y(men_men_n1058_));
  NO3        u1030(.A(men_men_n456_), .B(men_men_n321_), .C(men_men_n75_), .Y(men_men_n1059_));
  NA2        u1031(.A(men_men_n1059_), .B(men_men_n1058_), .Y(men_men_n1060_));
  NA2        u1032(.A(men_men_n1060_), .B(men_men_n1057_), .Y(men_men_n1061_));
  OAI220     u1033(.A0(men_men_n1048_), .A1(men_men_n238_), .B0(men_men_n1016_), .B1(men_men_n634_), .Y(men_men_n1062_));
  NO2        u1034(.A(men_men_n690_), .B(men_men_n394_), .Y(men_men_n1063_));
  NA2        u1035(.A(men_men_n972_), .B(men_men_n963_), .Y(men_men_n1064_));
  NO3        u1036(.A(men_men_n570_), .B(men_men_n156_), .C(men_men_n220_), .Y(men_men_n1065_));
  OAI210     u1037(.A0(men_men_n1065_), .A1(men_men_n550_), .B0(men_men_n395_), .Y(men_men_n1066_));
  OAI220     u1038(.A0(men_men_n969_), .A1(men_men_n976_), .B0(men_men_n571_), .B1(men_men_n445_), .Y(men_men_n1067_));
  NA4        u1039(.A(men_men_n1067_), .B(men_men_n1066_), .C(men_men_n1064_), .D(men_men_n648_), .Y(men_men_n1068_));
  NA3        u1040(.A(men_men_n1012_), .B(men_men_n507_), .C(men_men_n46_), .Y(men_men_n1069_));
  AOI210     u1041(.A0(men_men_n397_), .A1(men_men_n395_), .B0(men_men_n344_), .Y(men_men_n1070_));
  NA3        u1042(.A(men_men_n1070_), .B(men_men_n1069_), .C(men_men_n279_), .Y(men_men_n1071_));
  OR4        u1043(.A(men_men_n1071_), .B(men_men_n1068_), .C(men_men_n1063_), .D(men_men_n1062_), .Y(men_men_n1072_));
  NO4        u1044(.A(men_men_n1072_), .B(men_men_n1061_), .C(men_men_n1056_), .D(men_men_n1054_), .Y(men_men_n1073_));
  NA4        u1045(.A(men_men_n1073_), .B(men_men_n1047_), .C(men_men_n1004_), .D(men_men_n988_), .Y(men13));
  NA2        u1046(.A(men_men_n46_), .B(men_men_n89_), .Y(men_men_n1075_));
  AN2        u1047(.A(c), .B(b), .Y(men_men_n1076_));
  NA3        u1048(.A(men_men_n255_), .B(men_men_n1076_), .C(m), .Y(men_men_n1077_));
  NO4        u1049(.A(e), .B(men_men_n1077_), .C(men_men_n1075_), .D(men_men_n612_), .Y(men_men_n1078_));
  INV        u1050(.A(men_men_n270_), .Y(men_men_n1079_));
  NO4        u1051(.A(men_men_n1079_), .B(e), .C(men_men_n1006_), .D(a), .Y(men_men_n1080_));
  NAi32      u1052(.An(d), .Bn(c), .C(e), .Y(men_men_n1081_));
  NO4        u1053(.A(men_men_n1601_), .B(men_men_n1081_), .C(men_men_n619_), .D(men_men_n317_), .Y(men_men_n1082_));
  NA2        u1054(.A(men_men_n697_), .B(men_men_n232_), .Y(men_men_n1083_));
  NA2        u1055(.A(men_men_n427_), .B(men_men_n220_), .Y(men_men_n1084_));
  AN2        u1056(.A(d), .B(c), .Y(men_men_n1085_));
  NA2        u1057(.A(men_men_n1085_), .B(men_men_n120_), .Y(men_men_n1086_));
  NO4        u1058(.A(men_men_n1086_), .B(men_men_n1084_), .C(men_men_n182_), .D(men_men_n176_), .Y(men_men_n1087_));
  NA2        u1059(.A(men_men_n518_), .B(c), .Y(men_men_n1088_));
  NO4        u1060(.A(men_men_n1601_), .B(men_men_n615_), .C(men_men_n1088_), .D(men_men_n317_), .Y(men_men_n1089_));
  AO210      u1061(.A0(men_men_n1087_), .A1(men_men_n1083_), .B0(men_men_n1089_), .Y(men_men_n1090_));
  OR4        u1062(.A(men_men_n1090_), .B(men_men_n1082_), .C(men_men_n1080_), .D(men_men_n1078_), .Y(men_men_n1091_));
  NAi32      u1063(.An(f), .Bn(e), .C(c), .Y(men_men_n1092_));
  NO2        u1064(.A(men_men_n1092_), .B(men_men_n153_), .Y(men_men_n1093_));
  NA2        u1065(.A(men_men_n1093_), .B(g), .Y(men_men_n1094_));
  OR3        u1066(.A(men_men_n232_), .B(men_men_n182_), .C(men_men_n176_), .Y(men_men_n1095_));
  NO2        u1067(.A(men_men_n1095_), .B(men_men_n1094_), .Y(men_men_n1096_));
  NO2        u1068(.A(men_men_n1088_), .B(men_men_n317_), .Y(men_men_n1097_));
  NO2        u1069(.A(j), .B(men_men_n45_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n658_), .B(men_men_n1098_), .Y(men_men_n1099_));
  NOi21      u1071(.An(men_men_n1097_), .B(men_men_n1099_), .Y(men_men_n1100_));
  NO2        u1072(.A(men_men_n793_), .B(men_men_n116_), .Y(men_men_n1101_));
  NOi41      u1073(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1102_));
  NA2        u1074(.A(men_men_n1102_), .B(men_men_n1101_), .Y(men_men_n1103_));
  NO2        u1075(.A(men_men_n1103_), .B(men_men_n1094_), .Y(men_men_n1104_));
  OR3        u1076(.A(e), .B(d), .C(c), .Y(men_men_n1105_));
  NA3        u1077(.A(k), .B(j), .C(i), .Y(men_men_n1106_));
  NO3        u1078(.A(men_men_n1106_), .B(men_men_n317_), .C(men_men_n93_), .Y(men_men_n1107_));
  BUFFER     u1079(.A(men_men_n1107_), .Y(men_men_n1108_));
  OR4        u1080(.A(men_men_n1108_), .B(men_men_n1104_), .C(men_men_n1100_), .D(men_men_n1096_), .Y(men_men_n1109_));
  NA3        u1081(.A(men_men_n486_), .B(men_men_n347_), .C(men_men_n56_), .Y(men_men_n1110_));
  NO2        u1082(.A(men_men_n1110_), .B(men_men_n1099_), .Y(men_men_n1111_));
  NO3        u1083(.A(men_men_n1110_), .B(men_men_n615_), .C(men_men_n45_), .Y(men_men_n1112_));
  NO2        u1084(.A(f), .B(c), .Y(men_men_n1113_));
  NOi21      u1085(.An(men_men_n1113_), .B(men_men_n461_), .Y(men_men_n1114_));
  NA2        u1086(.A(men_men_n1114_), .B(men_men_n59_), .Y(men_men_n1115_));
  OR2        u1087(.A(k), .B(i), .Y(men_men_n1116_));
  NO3        u1088(.A(men_men_n1116_), .B(men_men_n248_), .C(l), .Y(men_men_n1117_));
  NOi21      u1089(.An(men_men_n1117_), .B(men_men_n1115_), .Y(men_men_n1118_));
  OR3        u1090(.A(men_men_n1118_), .B(men_men_n1112_), .C(men_men_n1111_), .Y(men_men_n1119_));
  OR3        u1091(.A(men_men_n1119_), .B(men_men_n1109_), .C(men_men_n1091_), .Y(men02));
  OR2        u1092(.A(l), .B(k), .Y(men_men_n1121_));
  OR3        u1093(.A(n), .B(m), .C(i), .Y(men_men_n1122_));
  NO4        u1094(.A(men_men_n1122_), .B(h), .C(men_men_n1121_), .D(men_men_n1105_), .Y(men_men_n1123_));
  NOi31      u1095(.An(e), .B(d), .C(c), .Y(men_men_n1124_));
  NO2        u1096(.A(men_men_n1107_), .B(men_men_n1082_), .Y(men_men_n1125_));
  AN3        u1097(.A(g), .B(f), .C(c), .Y(men_men_n1126_));
  NA3        u1098(.A(men_men_n1126_), .B(men_men_n486_), .C(h), .Y(men_men_n1127_));
  OR2        u1099(.A(men_men_n1106_), .B(men_men_n1127_), .Y(men_men_n1128_));
  NO3        u1100(.A(men_men_n1110_), .B(men_men_n1601_), .C(men_men_n615_), .Y(men_men_n1129_));
  NO2        u1101(.A(men_men_n1129_), .B(men_men_n1096_), .Y(men_men_n1130_));
  NA3        u1102(.A(l), .B(k), .C(j), .Y(men_men_n1131_));
  NA2        u1103(.A(i), .B(h), .Y(men_men_n1132_));
  NO3        u1104(.A(men_men_n148_), .B(men_men_n291_), .C(men_men_n221_), .Y(men_men_n1133_));
  INV        u1105(.A(men_men_n1100_), .Y(men_men_n1134_));
  NA3        u1106(.A(c), .B(b), .C(a), .Y(men_men_n1135_));
  NO3        u1107(.A(men_men_n1135_), .B(men_men_n939_), .C(men_men_n220_), .Y(men_men_n1136_));
  INV        u1108(.A(men_men_n1111_), .Y(men_men_n1137_));
  AN4        u1109(.A(men_men_n1137_), .B(men_men_n1134_), .C(men_men_n1130_), .D(men_men_n1128_), .Y(men_men_n1138_));
  NO2        u1110(.A(men_men_n1086_), .B(men_men_n1084_), .Y(men_men_n1139_));
  NA2        u1111(.A(men_men_n1103_), .B(men_men_n1095_), .Y(men_men_n1140_));
  AOI210     u1112(.A0(men_men_n1140_), .A1(men_men_n1139_), .B0(men_men_n1078_), .Y(men_men_n1141_));
  NAi41      u1113(.An(men_men_n1123_), .B(men_men_n1141_), .C(men_men_n1138_), .D(men_men_n1125_), .Y(men03));
  NO2        u1114(.A(men_men_n552_), .B(men_men_n628_), .Y(men_men_n1143_));
  NA4        u1115(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n220_), .Y(men_men_n1144_));
  NA4        u1116(.A(men_men_n603_), .B(m), .C(men_men_n116_), .D(men_men_n220_), .Y(men_men_n1145_));
  NA3        u1117(.A(men_men_n1145_), .B(men_men_n385_), .C(men_men_n1144_), .Y(men_men_n1146_));
  NO3        u1118(.A(men_men_n1146_), .B(men_men_n1143_), .C(men_men_n1041_), .Y(men_men_n1147_));
  NOi41      u1119(.An(men_men_n841_), .B(men_men_n891_), .C(men_men_n880_), .D(men_men_n743_), .Y(men_men_n1148_));
  OAI220     u1120(.A0(men_men_n1148_), .A1(men_men_n717_), .B0(men_men_n1147_), .B1(men_men_n616_), .Y(men_men_n1149_));
  NOi31      u1121(.An(i), .B(k), .C(j), .Y(men_men_n1150_));
  NA4        u1122(.A(men_men_n1150_), .B(men_men_n1124_), .C(men_men_n356_), .D(men_men_n347_), .Y(men_men_n1151_));
  OAI210     u1123(.A0(men_men_n855_), .A1(men_men_n438_), .B0(men_men_n1151_), .Y(men_men_n1152_));
  NOi31      u1124(.An(m), .B(n), .C(f), .Y(men_men_n1153_));
  NA2        u1125(.A(men_men_n1153_), .B(men_men_n51_), .Y(men_men_n1154_));
  AN2        u1126(.A(e), .B(c), .Y(men_men_n1155_));
  NA2        u1127(.A(men_men_n1155_), .B(a), .Y(men_men_n1156_));
  OAI220     u1128(.A0(men_men_n1156_), .A1(men_men_n1154_), .B0(men_men_n923_), .B1(men_men_n444_), .Y(men_men_n1157_));
  NA2        u1129(.A(men_men_n531_), .B(l), .Y(men_men_n1158_));
  NOi31      u1130(.An(men_men_n900_), .B(men_men_n1077_), .C(men_men_n1158_), .Y(men_men_n1159_));
  NO4        u1131(.A(men_men_n1159_), .B(men_men_n1157_), .C(men_men_n1152_), .D(men_men_n1040_), .Y(men_men_n1160_));
  NO2        u1132(.A(men_men_n291_), .B(a), .Y(men_men_n1161_));
  INV        u1133(.A(men_men_n1082_), .Y(men_men_n1162_));
  NO2        u1134(.A(men_men_n1132_), .B(men_men_n505_), .Y(men_men_n1163_));
  NO2        u1135(.A(men_men_n89_), .B(g), .Y(men_men_n1164_));
  AOI210     u1136(.A0(men_men_n1164_), .A1(men_men_n1163_), .B0(men_men_n1117_), .Y(men_men_n1165_));
  OR2        u1137(.A(men_men_n1165_), .B(men_men_n1115_), .Y(men_men_n1166_));
  NA3        u1138(.A(men_men_n1166_), .B(men_men_n1162_), .C(men_men_n1160_), .Y(men_men_n1167_));
  NO4        u1139(.A(men_men_n1167_), .B(men_men_n1149_), .C(men_men_n857_), .D(men_men_n592_), .Y(men_men_n1168_));
  NA2        u1140(.A(c), .B(b), .Y(men_men_n1169_));
  NO2        u1141(.A(men_men_n728_), .B(men_men_n1169_), .Y(men_men_n1170_));
  OAI210     u1142(.A0(men_men_n898_), .A1(men_men_n871_), .B0(men_men_n431_), .Y(men_men_n1171_));
  OAI210     u1143(.A0(men_men_n1171_), .A1(men_men_n899_), .B0(men_men_n1170_), .Y(men_men_n1172_));
  NAi21      u1144(.An(men_men_n439_), .B(men_men_n1170_), .Y(men_men_n1173_));
  NA3        u1145(.A(men_men_n445_), .B(men_men_n585_), .C(f), .Y(men_men_n1174_));
  OAI210     u1146(.A0(men_men_n575_), .A1(men_men_n39_), .B0(men_men_n1161_), .Y(men_men_n1175_));
  NA3        u1147(.A(men_men_n1175_), .B(men_men_n1174_), .C(men_men_n1173_), .Y(men_men_n1176_));
  NA2        u1148(.A(men_men_n266_), .B(men_men_n123_), .Y(men_men_n1177_));
  OAI210     u1149(.A0(men_men_n1177_), .A1(men_men_n295_), .B0(g), .Y(men_men_n1178_));
  NAi21      u1150(.An(f), .B(d), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n1179_), .B(men_men_n1135_), .Y(men_men_n1180_));
  INV        u1152(.A(men_men_n1180_), .Y(men_men_n1181_));
  AOI210     u1153(.A0(men_men_n1178_), .A1(men_men_n301_), .B0(men_men_n1181_), .Y(men_men_n1182_));
  AOI210     u1154(.A0(men_men_n1182_), .A1(men_men_n117_), .B0(men_men_n1176_), .Y(men_men_n1183_));
  NA2        u1155(.A(men_men_n489_), .B(men_men_n488_), .Y(men_men_n1184_));
  NO2        u1156(.A(men_men_n188_), .B(men_men_n241_), .Y(men_men_n1185_));
  NA2        u1157(.A(men_men_n1185_), .B(m), .Y(men_men_n1186_));
  NA3        u1158(.A(men_men_n953_), .B(men_men_n1158_), .C(men_men_n492_), .Y(men_men_n1187_));
  OAI210     u1159(.A0(men_men_n1187_), .A1(men_men_n322_), .B0(men_men_n490_), .Y(men_men_n1188_));
  AOI210     u1160(.A0(men_men_n1188_), .A1(men_men_n1184_), .B0(men_men_n1186_), .Y(men_men_n1189_));
  NA2        u1161(.A(men_men_n587_), .B(men_men_n426_), .Y(men_men_n1190_));
  NA2        u1162(.A(men_men_n165_), .B(men_men_n33_), .Y(men_men_n1191_));
  AOI210     u1163(.A0(men_men_n1002_), .A1(men_men_n1191_), .B0(men_men_n221_), .Y(men_men_n1192_));
  OAI210     u1164(.A0(men_men_n1192_), .A1(men_men_n465_), .B0(men_men_n1180_), .Y(men_men_n1193_));
  NO2        u1165(.A(men_men_n388_), .B(men_men_n387_), .Y(men_men_n1194_));
  AOI210     u1166(.A0(men_men_n1185_), .A1(men_men_n447_), .B0(men_men_n996_), .Y(men_men_n1195_));
  NAi41      u1167(.An(men_men_n1194_), .B(men_men_n1195_), .C(men_men_n1193_), .D(men_men_n1190_), .Y(men_men_n1196_));
  NO2        u1168(.A(men_men_n1196_), .B(men_men_n1189_), .Y(men_men_n1197_));
  NA4        u1169(.A(men_men_n1197_), .B(men_men_n1183_), .C(men_men_n1172_), .D(men_men_n1168_), .Y(men00));
  AOI210     u1170(.A0(men_men_n308_), .A1(men_men_n221_), .B0(men_men_n283_), .Y(men_men_n1199_));
  NO2        u1171(.A(men_men_n1199_), .B(men_men_n606_), .Y(men_men_n1200_));
  AOI210     u1172(.A0(men_men_n936_), .A1(men_men_n978_), .B0(men_men_n1152_), .Y(men_men_n1201_));
  NO3        u1173(.A(men_men_n1129_), .B(men_men_n996_), .C(men_men_n740_), .Y(men_men_n1202_));
  NA3        u1174(.A(men_men_n1202_), .B(men_men_n1201_), .C(men_men_n1042_), .Y(men_men_n1203_));
  NA2        u1175(.A(men_men_n533_), .B(f), .Y(men_men_n1204_));
  OAI210     u1176(.A0(men_men_n1049_), .A1(men_men_n40_), .B0(men_men_n677_), .Y(men_men_n1205_));
  NA2        u1177(.A(men_men_n1205_), .B(men_men_n262_), .Y(men_men_n1206_));
  AOI210     u1178(.A0(men_men_n1206_), .A1(men_men_n1204_), .B0(men_men_n1086_), .Y(men_men_n1207_));
  NO4        u1179(.A(men_men_n1207_), .B(men_men_n1203_), .C(men_men_n1200_), .D(men_men_n1109_), .Y(men_men_n1208_));
  NA3        u1180(.A(men_men_n175_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1209_));
  NA3        u1181(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1210_));
  NOi31      u1182(.An(n), .B(m), .C(i), .Y(men_men_n1211_));
  NA3        u1183(.A(men_men_n1211_), .B(men_men_n679_), .C(men_men_n51_), .Y(men_men_n1212_));
  OAI210     u1184(.A0(men_men_n1210_), .A1(men_men_n1209_), .B0(men_men_n1212_), .Y(men_men_n1213_));
  INV        u1185(.A(men_men_n605_), .Y(men_men_n1214_));
  NO4        u1186(.A(men_men_n1214_), .B(men_men_n1213_), .C(men_men_n1194_), .D(men_men_n956_), .Y(men_men_n1215_));
  NO4        u1187(.A(men_men_n508_), .B(men_men_n370_), .C(men_men_n1169_), .D(men_men_n59_), .Y(men_men_n1216_));
  NA3        u1188(.A(men_men_n400_), .B(men_men_n228_), .C(g), .Y(men_men_n1217_));
  OA220      u1189(.A0(men_men_n1217_), .A1(men_men_n1210_), .B0(men_men_n401_), .B1(men_men_n140_), .Y(men_men_n1218_));
  NO2        u1190(.A(h), .B(g), .Y(men_men_n1219_));
  NA4        u1191(.A(men_men_n521_), .B(men_men_n486_), .C(men_men_n1219_), .D(men_men_n1076_), .Y(men_men_n1220_));
  OAI220     u1192(.A0(men_men_n552_), .A1(men_men_n628_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1221_));
  AOI220     u1193(.A0(men_men_n1221_), .A1(men_men_n561_), .B0(men_men_n983_), .B1(men_men_n604_), .Y(men_men_n1222_));
  AOI220     u1194(.A0(men_men_n329_), .A1(men_men_n252_), .B0(men_men_n183_), .B1(men_men_n155_), .Y(men_men_n1223_));
  NA4        u1195(.A(men_men_n1223_), .B(men_men_n1222_), .C(men_men_n1220_), .D(men_men_n1218_), .Y(men_men_n1224_));
  NO3        u1196(.A(men_men_n1224_), .B(men_men_n1216_), .C(men_men_n272_), .Y(men_men_n1225_));
  INV        u1197(.A(men_men_n334_), .Y(men_men_n1226_));
  AOI210     u1198(.A0(men_men_n252_), .A1(men_men_n361_), .B0(men_men_n607_), .Y(men_men_n1227_));
  NA3        u1199(.A(men_men_n1227_), .B(men_men_n1226_), .C(men_men_n160_), .Y(men_men_n1228_));
  NO2        u1200(.A(men_men_n243_), .B(men_men_n187_), .Y(men_men_n1229_));
  NA2        u1201(.A(men_men_n1229_), .B(men_men_n445_), .Y(men_men_n1230_));
  NA3        u1202(.A(men_men_n185_), .B(men_men_n116_), .C(g), .Y(men_men_n1231_));
  NOi31      u1203(.An(men_men_n908_), .B(h), .C(men_men_n1231_), .Y(men_men_n1232_));
  NAi31      u1204(.An(men_men_n192_), .B(men_men_n895_), .C(men_men_n486_), .Y(men_men_n1233_));
  NAi31      u1205(.An(men_men_n1232_), .B(men_men_n1233_), .C(men_men_n1230_), .Y(men_men_n1234_));
  NO2        u1206(.A(men_men_n282_), .B(men_men_n75_), .Y(men_men_n1235_));
  NO3        u1207(.A(men_men_n444_), .B(men_men_n867_), .C(n), .Y(men_men_n1236_));
  AOI210     u1208(.A0(men_men_n1236_), .A1(men_men_n1235_), .B0(men_men_n1123_), .Y(men_men_n1237_));
  NAi31      u1209(.An(men_men_n1089_), .B(men_men_n1237_), .C(men_men_n74_), .Y(men_men_n1238_));
  NO4        u1210(.A(men_men_n1238_), .B(men_men_n1234_), .C(men_men_n1228_), .D(men_men_n543_), .Y(men_men_n1239_));
  AN3        u1211(.A(men_men_n1239_), .B(men_men_n1225_), .C(men_men_n1215_), .Y(men_men_n1240_));
  NA2        u1212(.A(men_men_n561_), .B(men_men_n104_), .Y(men_men_n1241_));
  NA3        u1213(.A(men_men_n1153_), .B(men_men_n637_), .C(men_men_n485_), .Y(men_men_n1242_));
  NA4        u1214(.A(men_men_n1242_), .B(men_men_n588_), .C(men_men_n1241_), .D(men_men_n246_), .Y(men_men_n1243_));
  NA2        u1215(.A(men_men_n1146_), .B(men_men_n561_), .Y(men_men_n1244_));
  NA4        u1216(.A(men_men_n679_), .B(men_men_n212_), .C(men_men_n228_), .D(men_men_n169_), .Y(men_men_n1245_));
  NA3        u1217(.A(men_men_n1245_), .B(men_men_n1244_), .C(men_men_n305_), .Y(men_men_n1246_));
  OAI210     u1218(.A0(men_men_n484_), .A1(men_men_n124_), .B0(men_men_n901_), .Y(men_men_n1247_));
  AOI220     u1219(.A0(men_men_n1247_), .A1(men_men_n1187_), .B0(men_men_n587_), .B1(men_men_n426_), .Y(men_men_n1248_));
  OR3        u1220(.A(men_men_n1086_), .B(men_men_n230_), .C(e), .Y(men_men_n1249_));
  NO2        u1221(.A(men_men_n224_), .B(men_men_n221_), .Y(men_men_n1250_));
  NA2        u1222(.A(n), .B(e), .Y(men_men_n1251_));
  NO2        u1223(.A(men_men_n1251_), .B(men_men_n153_), .Y(men_men_n1252_));
  AOI220     u1224(.A0(men_men_n1252_), .A1(men_men_n280_), .B0(men_men_n884_), .B1(men_men_n1250_), .Y(men_men_n1253_));
  OAI210     u1225(.A0(men_men_n371_), .A1(men_men_n323_), .B0(men_men_n467_), .Y(men_men_n1254_));
  NA4        u1226(.A(men_men_n1254_), .B(men_men_n1253_), .C(men_men_n1249_), .D(men_men_n1248_), .Y(men_men_n1255_));
  AOI210     u1227(.A0(men_men_n1252_), .A1(men_men_n888_), .B0(men_men_n856_), .Y(men_men_n1256_));
  AOI220     u1228(.A0(men_men_n992_), .A1(men_men_n604_), .B0(men_men_n679_), .B1(men_men_n249_), .Y(men_men_n1257_));
  NO2        u1229(.A(men_men_n68_), .B(h), .Y(men_men_n1258_));
  NO3        u1230(.A(men_men_n1086_), .B(men_men_n1084_), .C(men_men_n755_), .Y(men_men_n1259_));
  NO2        u1231(.A(men_men_n1121_), .B(men_men_n137_), .Y(men_men_n1260_));
  AN2        u1232(.A(men_men_n1260_), .B(men_men_n1133_), .Y(men_men_n1261_));
  OAI210     u1233(.A0(men_men_n1261_), .A1(men_men_n1259_), .B0(men_men_n1258_), .Y(men_men_n1262_));
  NA4        u1234(.A(men_men_n1262_), .B(men_men_n1257_), .C(men_men_n1256_), .D(men_men_n903_), .Y(men_men_n1263_));
  NO4        u1235(.A(men_men_n1263_), .B(men_men_n1255_), .C(men_men_n1246_), .D(men_men_n1243_), .Y(men_men_n1264_));
  NA2        u1236(.A(men_men_n872_), .B(men_men_n788_), .Y(men_men_n1265_));
  NA4        u1237(.A(men_men_n1265_), .B(men_men_n1264_), .C(men_men_n1240_), .D(men_men_n1208_), .Y(men01));
  AN2        u1238(.A(men_men_n1066_), .B(men_men_n1064_), .Y(men_men_n1267_));
  NO4        u1239(.A(men_men_n837_), .B(men_men_n829_), .C(men_men_n500_), .D(men_men_n289_), .Y(men_men_n1268_));
  NO2        u1240(.A(men_men_n621_), .B(men_men_n298_), .Y(men_men_n1269_));
  INV        u1241(.A(men_men_n1269_), .Y(men_men_n1270_));
  NA3        u1242(.A(men_men_n1270_), .B(men_men_n1268_), .C(men_men_n1267_), .Y(men_men_n1271_));
  NA2        u1243(.A(men_men_n617_), .B(men_men_n92_), .Y(men_men_n1272_));
  NA2        u1244(.A(men_men_n581_), .B(men_men_n277_), .Y(men_men_n1273_));
  NA2        u1245(.A(men_men_n999_), .B(men_men_n1273_), .Y(men_men_n1274_));
  NA4        u1246(.A(men_men_n1274_), .B(men_men_n1272_), .C(men_men_n949_), .D(men_men_n346_), .Y(men_men_n1275_));
  NA2        u1247(.A(men_men_n45_), .B(f), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n735_), .B(men_men_n99_), .Y(men_men_n1277_));
  NO2        u1249(.A(men_men_n1277_), .B(men_men_n1276_), .Y(men_men_n1278_));
  OAI210     u1250(.A0(men_men_n815_), .A1(men_men_n634_), .B0(men_men_n1245_), .Y(men_men_n1279_));
  AOI210     u1251(.A0(men_men_n1278_), .A1(men_men_n665_), .B0(men_men_n1279_), .Y(men_men_n1280_));
  NA2        u1252(.A(men_men_n122_), .B(l), .Y(men_men_n1281_));
  OA220      u1253(.A0(men_men_n1281_), .A1(men_men_n614_), .B0(men_men_n691_), .B1(men_men_n385_), .Y(men_men_n1282_));
  NAi41      u1254(.An(men_men_n168_), .B(men_men_n1282_), .C(men_men_n1280_), .D(men_men_n935_), .Y(men_men_n1283_));
  NO3        u1255(.A(men_men_n816_), .B(men_men_n707_), .C(men_men_n536_), .Y(men_men_n1284_));
  NA4        u1256(.A(men_men_n735_), .B(men_men_n99_), .C(men_men_n45_), .D(men_men_n220_), .Y(men_men_n1285_));
  OR2        u1257(.A(men_men_n1285_), .B(men_men_n700_), .Y(men_men_n1286_));
  NA3        u1258(.A(men_men_n1286_), .B(men_men_n1284_), .C(men_men_n143_), .Y(men_men_n1287_));
  NO4        u1259(.A(men_men_n1287_), .B(men_men_n1283_), .C(men_men_n1275_), .D(men_men_n1271_), .Y(men_men_n1288_));
  NA2        u1260(.A(men_men_n1217_), .B(men_men_n213_), .Y(men_men_n1289_));
  OAI210     u1261(.A0(men_men_n1289_), .A1(men_men_n311_), .B0(men_men_n556_), .Y(men_men_n1290_));
  NA2        u1262(.A(men_men_n564_), .B(men_men_n412_), .Y(men_men_n1291_));
  NA2        u1263(.A(men_men_n76_), .B(i), .Y(men_men_n1292_));
  AOI210     u1264(.A0(men_men_n620_), .A1(men_men_n614_), .B0(men_men_n1292_), .Y(men_men_n1293_));
  NOi21      u1265(.An(men_men_n589_), .B(men_men_n611_), .Y(men_men_n1294_));
  AOI210     u1266(.A0(men_men_n1294_), .A1(men_men_n1291_), .B0(men_men_n1293_), .Y(men_men_n1295_));
  AOI210     u1267(.A0(men_men_n210_), .A1(men_men_n91_), .B0(men_men_n220_), .Y(men_men_n1296_));
  OAI210     u1268(.A0(men_men_n844_), .A1(men_men_n445_), .B0(men_men_n1296_), .Y(men_men_n1297_));
  AN3        u1269(.A(m), .B(l), .C(k), .Y(men_men_n1298_));
  OAI210     u1270(.A0(men_men_n373_), .A1(men_men_n34_), .B0(men_men_n1298_), .Y(men_men_n1299_));
  NA2        u1271(.A(men_men_n209_), .B(men_men_n34_), .Y(men_men_n1300_));
  AO210      u1272(.A0(men_men_n1300_), .A1(men_men_n1299_), .B0(men_men_n345_), .Y(men_men_n1301_));
  NA4        u1273(.A(men_men_n1301_), .B(men_men_n1297_), .C(men_men_n1295_), .D(men_men_n1290_), .Y(men_men_n1302_));
  AOI210     u1274(.A0(men_men_n626_), .A1(men_men_n122_), .B0(men_men_n632_), .Y(men_men_n1303_));
  OAI210     u1275(.A0(men_men_n1281_), .A1(men_men_n623_), .B0(men_men_n1303_), .Y(men_men_n1304_));
  NA2        u1276(.A(men_men_n288_), .B(men_men_n202_), .Y(men_men_n1305_));
  OAI210     u1277(.A0(men_men_n1305_), .A1(men_men_n402_), .B0(men_men_n696_), .Y(men_men_n1306_));
  NO3        u1278(.A(men_men_n855_), .B(men_men_n210_), .C(men_men_n424_), .Y(men_men_n1307_));
  NO2        u1279(.A(men_men_n1307_), .B(men_men_n996_), .Y(men_men_n1308_));
  OAI210     u1280(.A0(men_men_n1278_), .A1(men_men_n339_), .B0(men_men_n708_), .Y(men_men_n1309_));
  NA4        u1281(.A(men_men_n1309_), .B(men_men_n1308_), .C(men_men_n1306_), .D(men_men_n819_), .Y(men_men_n1310_));
  NO3        u1282(.A(men_men_n1310_), .B(men_men_n1304_), .C(men_men_n1302_), .Y(men_men_n1311_));
  NA3        u1283(.A(men_men_n635_), .B(men_men_n29_), .C(f), .Y(men_men_n1312_));
  NO2        u1284(.A(men_men_n1312_), .B(men_men_n210_), .Y(men_men_n1313_));
  AOI210     u1285(.A0(men_men_n528_), .A1(men_men_n58_), .B0(men_men_n1313_), .Y(men_men_n1314_));
  OR3        u1286(.A(men_men_n1277_), .B(men_men_n636_), .C(men_men_n1276_), .Y(men_men_n1315_));
  NA3        u1287(.A(men_men_n769_), .B(men_men_n76_), .C(i), .Y(men_men_n1316_));
  AOI210     u1288(.A0(men_men_n1316_), .A1(men_men_n1285_), .B0(men_men_n1019_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n213_), .B(men_men_n115_), .Y(men_men_n1318_));
  NO3        u1290(.A(men_men_n1318_), .B(men_men_n1317_), .C(men_men_n1213_), .Y(men_men_n1319_));
  NA4        u1291(.A(men_men_n1319_), .B(men_men_n1315_), .C(men_men_n1314_), .D(men_men_n787_), .Y(men_men_n1320_));
  NO2        u1292(.A(men_men_n1006_), .B(men_men_n237_), .Y(men_men_n1321_));
  NO2        u1293(.A(men_men_n1007_), .B(men_men_n582_), .Y(men_men_n1322_));
  OAI210     u1294(.A0(men_men_n1322_), .A1(men_men_n1321_), .B0(men_men_n354_), .Y(men_men_n1323_));
  NA2        u1295(.A(men_men_n599_), .B(men_men_n597_), .Y(men_men_n1324_));
  NO3        u1296(.A(men_men_n81_), .B(men_men_n309_), .C(men_men_n45_), .Y(men_men_n1325_));
  NA2        u1297(.A(men_men_n1325_), .B(men_men_n580_), .Y(men_men_n1326_));
  NA3        u1298(.A(men_men_n1326_), .B(men_men_n1324_), .C(men_men_n702_), .Y(men_men_n1327_));
  OR2        u1299(.A(men_men_n1217_), .B(men_men_n1210_), .Y(men_men_n1328_));
  NO2        u1300(.A(men_men_n385_), .B(men_men_n73_), .Y(men_men_n1329_));
  AOI210     u1301(.A0(men_men_n760_), .A1(men_men_n645_), .B0(men_men_n1329_), .Y(men_men_n1330_));
  NA2        u1302(.A(men_men_n1325_), .B(men_men_n847_), .Y(men_men_n1331_));
  NA4        u1303(.A(men_men_n1331_), .B(men_men_n1330_), .C(men_men_n1328_), .D(men_men_n403_), .Y(men_men_n1332_));
  NOi41      u1304(.An(men_men_n1323_), .B(men_men_n1332_), .C(men_men_n1327_), .D(men_men_n1320_), .Y(men_men_n1333_));
  NO2        u1305(.A(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1334_));
  AO220      u1306(.A0(i), .A1(men_men_n651_), .B0(men_men_n1334_), .B1(men_men_n733_), .Y(men_men_n1335_));
  NA2        u1307(.A(men_men_n1335_), .B(men_men_n354_), .Y(men_men_n1336_));
  NA2        u1308(.A(men_men_n479_), .B(men_men_n140_), .Y(men_men_n1337_));
  NO3        u1309(.A(men_men_n1132_), .B(men_men_n182_), .C(men_men_n89_), .Y(men_men_n1338_));
  AOI220     u1310(.A0(men_men_n1338_), .A1(men_men_n1337_), .B0(men_men_n1325_), .B1(men_men_n1010_), .Y(men_men_n1339_));
  NA2        u1311(.A(men_men_n1339_), .B(men_men_n1336_), .Y(men_men_n1340_));
  NO2        u1312(.A(men_men_n1340_), .B(men_men_n669_), .Y(men_men_n1341_));
  NA4        u1313(.A(men_men_n1341_), .B(men_men_n1333_), .C(men_men_n1311_), .D(men_men_n1288_), .Y(men06));
  NO2        u1314(.A(men_men_n425_), .B(men_men_n586_), .Y(men_men_n1343_));
  NO2        u1315(.A(men_men_n762_), .B(i), .Y(men_men_n1344_));
  OAI210     u1316(.A0(men_men_n1344_), .A1(men_men_n273_), .B0(men_men_n1343_), .Y(men_men_n1345_));
  NO2        u1317(.A(men_men_n232_), .B(men_men_n106_), .Y(men_men_n1346_));
  NA2        u1318(.A(men_men_n1346_), .B(men_men_n399_), .Y(men_men_n1347_));
  NO3        u1319(.A(men_men_n630_), .B(men_men_n842_), .C(men_men_n633_), .Y(men_men_n1348_));
  OR2        u1320(.A(men_men_n1348_), .B(men_men_n923_), .Y(men_men_n1349_));
  NA4        u1321(.A(men_men_n1349_), .B(men_men_n1347_), .C(men_men_n1345_), .D(men_men_n1323_), .Y(men_men_n1350_));
  NO3        u1322(.A(men_men_n1350_), .B(men_men_n1327_), .C(men_men_n261_), .Y(men_men_n1351_));
  NO2        u1323(.A(men_men_n309_), .B(men_men_n45_), .Y(men_men_n1352_));
  AOI210     u1324(.A0(men_men_n1352_), .A1(men_men_n1011_), .B0(men_men_n1321_), .Y(men_men_n1353_));
  AOI210     u1325(.A0(men_men_n1352_), .A1(men_men_n583_), .B0(men_men_n1335_), .Y(men_men_n1354_));
  AOI210     u1326(.A0(men_men_n1354_), .A1(men_men_n1353_), .B0(men_men_n351_), .Y(men_men_n1355_));
  OAI210     u1327(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n706_), .Y(men_men_n1356_));
  NA2        u1328(.A(men_men_n1356_), .B(men_men_n673_), .Y(men_men_n1357_));
  NO2        u1329(.A(men_men_n539_), .B(men_men_n179_), .Y(men_men_n1358_));
  NOi21      u1330(.An(men_men_n142_), .B(men_men_n45_), .Y(men_men_n1359_));
  NO2        u1331(.A(men_men_n638_), .B(men_men_n1154_), .Y(men_men_n1360_));
  OAI210     u1332(.A0(men_men_n479_), .A1(men_men_n253_), .B0(men_men_n943_), .Y(men_men_n1361_));
  NO4        u1333(.A(men_men_n1361_), .B(men_men_n1360_), .C(men_men_n1359_), .D(men_men_n1358_), .Y(men_men_n1362_));
  OR2        u1334(.A(men_men_n631_), .B(men_men_n629_), .Y(men_men_n1363_));
  NO2        u1335(.A(men_men_n384_), .B(men_men_n141_), .Y(men_men_n1364_));
  AOI210     u1336(.A0(men_men_n1364_), .A1(men_men_n617_), .B0(men_men_n1363_), .Y(men_men_n1365_));
  NA3        u1337(.A(men_men_n1365_), .B(men_men_n1362_), .C(men_men_n1357_), .Y(men_men_n1366_));
  NO2        u1338(.A(men_men_n778_), .B(men_men_n383_), .Y(men_men_n1367_));
  NO3        u1339(.A(men_men_n708_), .B(men_men_n789_), .C(men_men_n665_), .Y(men_men_n1368_));
  NOi21      u1340(.An(men_men_n1367_), .B(men_men_n1368_), .Y(men_men_n1369_));
  AN2        u1341(.A(men_men_n992_), .B(men_men_n676_), .Y(men_men_n1370_));
  NO4        u1342(.A(men_men_n1370_), .B(men_men_n1369_), .C(men_men_n1366_), .D(men_men_n1355_), .Y(men_men_n1371_));
  NO2        u1343(.A(men_men_n836_), .B(men_men_n284_), .Y(men_men_n1372_));
  OAI220     u1344(.A0(men_men_n762_), .A1(men_men_n47_), .B0(men_men_n232_), .B1(men_men_n644_), .Y(men_men_n1373_));
  OAI210     u1345(.A0(men_men_n284_), .A1(c), .B0(men_men_n672_), .Y(men_men_n1374_));
  AOI220     u1346(.A0(men_men_n1374_), .A1(men_men_n1373_), .B0(men_men_n1372_), .B1(men_men_n273_), .Y(men_men_n1375_));
  NO3        u1347(.A(men_men_n248_), .B(men_men_n106_), .C(men_men_n291_), .Y(men_men_n1376_));
  OAI210     u1348(.A0(l), .A1(i), .B0(k), .Y(men_men_n1377_));
  NO3        u1349(.A(men_men_n1377_), .B(men_men_n628_), .C(j), .Y(men_men_n1378_));
  NOi21      u1350(.An(men_men_n1378_), .B(men_men_n700_), .Y(men_men_n1379_));
  NO3        u1351(.A(men_men_n1379_), .B(men_men_n1376_), .C(men_men_n1157_), .Y(men_men_n1380_));
  NA4        u1352(.A(men_men_n827_), .B(men_men_n826_), .C(men_men_n455_), .D(men_men_n915_), .Y(men_men_n1381_));
  NAi31      u1353(.An(men_men_n778_), .B(men_men_n1381_), .C(men_men_n209_), .Y(men_men_n1382_));
  NA4        u1354(.A(men_men_n1382_), .B(men_men_n1380_), .C(men_men_n1375_), .D(men_men_n1257_), .Y(men_men_n1383_));
  NOi31      u1355(.An(men_men_n1348_), .B(men_men_n483_), .C(men_men_n411_), .Y(men_men_n1384_));
  OR3        u1356(.A(men_men_n1384_), .B(men_men_n815_), .C(men_men_n567_), .Y(men_men_n1385_));
  OR3        u1357(.A(men_men_n387_), .B(men_men_n232_), .C(men_men_n644_), .Y(men_men_n1386_));
  AOI210     u1358(.A0(men_men_n599_), .A1(men_men_n467_), .B0(men_men_n389_), .Y(men_men_n1387_));
  NA2        u1359(.A(men_men_n1378_), .B(men_men_n823_), .Y(men_men_n1388_));
  NA4        u1360(.A(men_men_n1388_), .B(men_men_n1387_), .C(men_men_n1386_), .D(men_men_n1385_), .Y(men_men_n1389_));
  AOI220     u1361(.A0(men_men_n1367_), .A1(men_men_n788_), .B0(men_men_n1364_), .B1(men_men_n242_), .Y(men_men_n1390_));
  AN2        u1362(.A(men_men_n964_), .B(men_men_n963_), .Y(men_men_n1391_));
  NO3        u1363(.A(men_men_n1391_), .B(men_men_n913_), .C(men_men_n524_), .Y(men_men_n1392_));
  NA3        u1364(.A(men_men_n1392_), .B(men_men_n1390_), .C(men_men_n1331_), .Y(men_men_n1393_));
  NO3        u1365(.A(men_men_n1393_), .B(men_men_n1389_), .C(men_men_n1383_), .Y(men_men_n1394_));
  NA4        u1366(.A(men_men_n1394_), .B(men_men_n1371_), .C(men_men_n1351_), .D(men_men_n1341_), .Y(men07));
  NOi21      u1367(.An(j), .B(k), .Y(men_men_n1396_));
  NA4        u1368(.A(men_men_n185_), .B(men_men_n112_), .C(men_men_n1396_), .D(f), .Y(men_men_n1397_));
  NAi32      u1369(.An(m), .Bn(b), .C(n), .Y(men_men_n1398_));
  NAi21      u1370(.An(f), .B(c), .Y(men_men_n1399_));
  NOi31      u1371(.An(n), .B(m), .C(b), .Y(men_men_n1400_));
  NO3        u1372(.A(men_men_n137_), .B(men_men_n469_), .C(h), .Y(men_men_n1401_));
  NOi41      u1373(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1402_));
  NA3        u1374(.A(men_men_n1402_), .B(men_men_n905_), .C(men_men_n427_), .Y(men_men_n1403_));
  NOi21      u1375(.An(h), .B(k), .Y(men_men_n1404_));
  NO2        u1376(.A(men_men_n1403_), .B(men_men_n56_), .Y(men_men_n1405_));
  NA2        u1377(.A(men_men_n1133_), .B(men_men_n228_), .Y(men_men_n1406_));
  NO2        u1378(.A(men_men_n1406_), .B(men_men_n61_), .Y(men_men_n1407_));
  NO2        u1379(.A(k), .B(i), .Y(men_men_n1408_));
  NA2        u1380(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1409_));
  NO2        u1381(.A(men_men_n1092_), .B(men_men_n461_), .Y(men_men_n1410_));
  NA3        u1382(.A(men_men_n1410_), .B(men_men_n1409_), .C(men_men_n221_), .Y(men_men_n1411_));
  NO2        u1383(.A(men_men_n1106_), .B(men_men_n317_), .Y(men_men_n1412_));
  NA2        u1384(.A(men_men_n568_), .B(men_men_n82_), .Y(men_men_n1413_));
  NA2        u1385(.A(men_men_n1258_), .B(men_men_n299_), .Y(men_men_n1414_));
  NA3        u1386(.A(men_men_n1414_), .B(men_men_n1413_), .C(men_men_n1411_), .Y(men_men_n1415_));
  NO4        u1387(.A(men_men_n1415_), .B(men_men_n1407_), .C(men_men_n1405_), .D(men_men_n1598_), .Y(men_men_n1416_));
  OR2        u1388(.A(h), .B(f), .Y(men_men_n1417_));
  NO3        u1389(.A(n), .B(m), .C(i), .Y(men_men_n1418_));
  OAI210     u1390(.A0(men_men_n1155_), .A1(men_men_n163_), .B0(men_men_n1418_), .Y(men_men_n1419_));
  NO2        u1391(.A(i), .B(g), .Y(men_men_n1420_));
  OR3        u1392(.A(men_men_n1420_), .B(men_men_n1398_), .C(men_men_n72_), .Y(men_men_n1421_));
  OAI220     u1393(.A0(men_men_n1421_), .A1(men_men_n504_), .B0(men_men_n1419_), .B1(men_men_n1417_), .Y(men_men_n1422_));
  NA3        u1394(.A(men_men_n723_), .B(men_men_n714_), .C(men_men_n116_), .Y(men_men_n1423_));
  NA3        u1395(.A(men_men_n1400_), .B(men_men_n1101_), .C(men_men_n704_), .Y(men_men_n1424_));
  AOI210     u1396(.A0(men_men_n1424_), .A1(men_men_n1423_), .B0(men_men_n45_), .Y(men_men_n1425_));
  NA2        u1397(.A(men_men_n1418_), .B(men_men_n671_), .Y(men_men_n1426_));
  NO2        u1398(.A(l), .B(k), .Y(men_men_n1427_));
  NOi41      u1399(.An(men_men_n573_), .B(men_men_n1427_), .C(men_men_n498_), .D(men_men_n461_), .Y(men_men_n1428_));
  NO3        u1400(.A(men_men_n461_), .B(d), .C(c), .Y(men_men_n1429_));
  NO3        u1401(.A(men_men_n1428_), .B(men_men_n1425_), .C(men_men_n1422_), .Y(men_men_n1430_));
  NO2        u1402(.A(men_men_n154_), .B(h), .Y(men_men_n1431_));
  NO2        u1403(.A(g), .B(c), .Y(men_men_n1432_));
  OAI210     u1404(.A0(men_men_n1404_), .A1(men_men_n220_), .B0(men_men_n1116_), .Y(men_men_n1433_));
  NO2        u1405(.A(men_men_n472_), .B(a), .Y(men_men_n1434_));
  NA3        u1406(.A(men_men_n1434_), .B(men_men_n1433_), .C(men_men_n117_), .Y(men_men_n1435_));
  NO2        u1407(.A(i), .B(h), .Y(men_men_n1436_));
  NA2        u1408(.A(men_men_n1436_), .B(men_men_n228_), .Y(men_men_n1437_));
  AOI210     u1409(.A0(men_men_n262_), .A1(men_men_n120_), .B0(men_men_n556_), .Y(men_men_n1438_));
  NO2        u1410(.A(men_men_n1438_), .B(men_men_n1437_), .Y(men_men_n1439_));
  NO2        u1411(.A(men_men_n785_), .B(men_men_n194_), .Y(men_men_n1440_));
  NOi31      u1412(.An(m), .B(n), .C(b), .Y(men_men_n1441_));
  NOi31      u1413(.An(f), .B(d), .C(c), .Y(men_men_n1442_));
  NA2        u1414(.A(men_men_n1442_), .B(men_men_n1441_), .Y(men_men_n1443_));
  INV        u1415(.A(men_men_n1443_), .Y(men_men_n1444_));
  NO3        u1416(.A(men_men_n1444_), .B(men_men_n1440_), .C(men_men_n1439_), .Y(men_men_n1445_));
  NA2        u1417(.A(men_men_n1126_), .B(men_men_n486_), .Y(men_men_n1446_));
  NO4        u1418(.A(men_men_n1446_), .B(men_men_n1101_), .C(men_men_n461_), .D(men_men_n45_), .Y(men_men_n1447_));
  OAI210     u1419(.A0(men_men_n188_), .A1(men_men_n551_), .B0(men_men_n1102_), .Y(men_men_n1448_));
  NO3        u1420(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1449_));
  INV        u1421(.A(men_men_n1448_), .Y(men_men_n1450_));
  NO2        u1422(.A(men_men_n1450_), .B(men_men_n1447_), .Y(men_men_n1451_));
  AN3        u1423(.A(men_men_n1451_), .B(men_men_n1445_), .C(men_men_n1435_), .Y(men_men_n1452_));
  NA2        u1424(.A(men_men_n1400_), .B(men_men_n396_), .Y(men_men_n1453_));
  NO2        u1425(.A(men_men_n1453_), .B(men_men_n1083_), .Y(men_men_n1454_));
  NO2        u1426(.A(men_men_n194_), .B(b), .Y(men_men_n1455_));
  NA2        u1427(.A(men_men_n1211_), .B(men_men_n1455_), .Y(men_men_n1456_));
  NO2        u1428(.A(i), .B(men_men_n220_), .Y(men_men_n1457_));
  NA4        u1429(.A(men_men_n1185_), .B(men_men_n1457_), .C(men_men_n107_), .D(m), .Y(men_men_n1458_));
  NAi31      u1430(.An(men_men_n1454_), .B(men_men_n1458_), .C(men_men_n1456_), .Y(men_men_n1459_));
  NO4        u1431(.A(men_men_n137_), .B(g), .C(f), .D(e), .Y(men_men_n1460_));
  NA2        u1432(.A(men_men_n1408_), .B(h), .Y(men_men_n1461_));
  NA2        u1433(.A(men_men_n201_), .B(men_men_n101_), .Y(men_men_n1462_));
  OR2        u1434(.A(e), .B(a), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n30_), .B(h), .Y(men_men_n1464_));
  NO2        u1436(.A(men_men_n1464_), .B(men_men_n1122_), .Y(men_men_n1465_));
  NOi41      u1437(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1466_));
  NA2        u1438(.A(men_men_n1466_), .B(men_men_n117_), .Y(men_men_n1467_));
  NA2        u1439(.A(men_men_n1402_), .B(men_men_n1427_), .Y(men_men_n1468_));
  NA2        u1440(.A(men_men_n1468_), .B(men_men_n1467_), .Y(men_men_n1469_));
  OR3        u1441(.A(men_men_n567_), .B(men_men_n566_), .C(men_men_n116_), .Y(men_men_n1470_));
  NA2        u1442(.A(men_men_n1153_), .B(men_men_n424_), .Y(men_men_n1471_));
  OAI220     u1443(.A0(men_men_n1471_), .A1(men_men_n454_), .B0(men_men_n1470_), .B1(men_men_n309_), .Y(men_men_n1472_));
  AO210      u1444(.A0(men_men_n1472_), .A1(men_men_n120_), .B0(men_men_n1469_), .Y(men_men_n1473_));
  NO3        u1445(.A(men_men_n1473_), .B(men_men_n1465_), .C(men_men_n1459_), .Y(men_men_n1474_));
  NA4        u1446(.A(men_men_n1474_), .B(men_men_n1452_), .C(men_men_n1430_), .D(men_men_n1416_), .Y(men_men_n1475_));
  NO2        u1447(.A(men_men_n1169_), .B(men_men_n114_), .Y(men_men_n1476_));
  NA2        u1448(.A(men_men_n396_), .B(men_men_n56_), .Y(men_men_n1477_));
  AOI210     u1449(.A0(men_men_n1477_), .A1(men_men_n1092_), .B0(men_men_n1426_), .Y(men_men_n1478_));
  NA2        u1450(.A(men_men_n222_), .B(men_men_n185_), .Y(men_men_n1479_));
  AOI210     u1451(.A0(men_men_n1479_), .A1(men_men_n1231_), .B0(men_men_n1477_), .Y(men_men_n1480_));
  NO2        u1452(.A(men_men_n1127_), .B(men_men_n1122_), .Y(men_men_n1481_));
  NO3        u1453(.A(men_men_n1481_), .B(men_men_n1480_), .C(men_men_n1478_), .Y(men_men_n1482_));
  NO2        u1454(.A(men_men_n408_), .B(j), .Y(men_men_n1483_));
  NA3        u1455(.A(men_men_n1449_), .B(e), .C(men_men_n1153_), .Y(men_men_n1484_));
  INV        u1456(.A(men_men_n1484_), .Y(men_men_n1485_));
  NA3        u1457(.A(g), .B(men_men_n1483_), .C(men_men_n165_), .Y(men_men_n1486_));
  INV        u1458(.A(men_men_n1486_), .Y(men_men_n1487_));
  NO2        u1459(.A(men_men_n1487_), .B(men_men_n1485_), .Y(men_men_n1488_));
  NO3        u1460(.A(men_men_n1122_), .B(men_men_n611_), .C(g), .Y(men_men_n1489_));
  NOi21      u1461(.An(men_men_n1479_), .B(men_men_n1489_), .Y(men_men_n1490_));
  AOI210     u1462(.A0(men_men_n1490_), .A1(men_men_n1462_), .B0(men_men_n1092_), .Y(men_men_n1491_));
  INV        u1463(.A(men_men_n49_), .Y(men_men_n1492_));
  NA2        u1464(.A(men_men_n1492_), .B(men_men_n1219_), .Y(men_men_n1493_));
  INV        u1465(.A(men_men_n1493_), .Y(men_men_n1494_));
  OAI220     u1466(.A0(men_men_n697_), .A1(g), .B0(men_men_n232_), .B1(c), .Y(men_men_n1495_));
  AOI210     u1467(.A0(men_men_n1455_), .A1(men_men_n41_), .B0(men_men_n1495_), .Y(men_men_n1496_));
  NO2        u1468(.A(men_men_n137_), .B(l), .Y(men_men_n1497_));
  NO2        u1469(.A(men_men_n232_), .B(k), .Y(men_men_n1498_));
  OAI210     u1470(.A0(men_men_n1498_), .A1(men_men_n1436_), .B0(men_men_n1497_), .Y(men_men_n1499_));
  OAI220     u1471(.A0(men_men_n1499_), .A1(men_men_n31_), .B0(men_men_n1496_), .B1(men_men_n182_), .Y(men_men_n1500_));
  NO3        u1472(.A(men_men_n1470_), .B(men_men_n486_), .C(men_men_n368_), .Y(men_men_n1501_));
  NO4        u1473(.A(men_men_n1501_), .B(men_men_n1500_), .C(men_men_n1494_), .D(men_men_n1491_), .Y(men_men_n1502_));
  NO2        u1474(.A(men_men_n49_), .B(men_men_n611_), .Y(men_men_n1503_));
  NA2        u1475(.A(men_men_n1136_), .B(men_men_n1503_), .Y(men_men_n1504_));
  NO2        u1476(.A(men_men_n1122_), .B(h), .Y(men_men_n1505_));
  NA3        u1477(.A(men_men_n1505_), .B(d), .C(men_men_n1084_), .Y(men_men_n1506_));
  OAI220     u1478(.A0(men_men_n1506_), .A1(c), .B0(men_men_n1504_), .B1(j), .Y(men_men_n1507_));
  NA3        u1479(.A(men_men_n1476_), .B(men_men_n486_), .C(f), .Y(men_men_n1508_));
  NO2        u1480(.A(men_men_n1396_), .B(men_men_n42_), .Y(men_men_n1509_));
  AOI210     u1481(.A0(men_men_n117_), .A1(men_men_n40_), .B0(men_men_n1509_), .Y(men_men_n1510_));
  NO2        u1482(.A(men_men_n1510_), .B(men_men_n1508_), .Y(men_men_n1511_));
  AOI210     u1483(.A0(men_men_n551_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1512_));
  NA2        u1484(.A(men_men_n1512_), .B(men_men_n1434_), .Y(men_men_n1513_));
  NO2        u1485(.A(j), .B(men_men_n181_), .Y(men_men_n1514_));
  NOi21      u1486(.An(d), .B(f), .Y(men_men_n1515_));
  NO3        u1487(.A(men_men_n1442_), .B(men_men_n1515_), .C(men_men_n40_), .Y(men_men_n1516_));
  NA2        u1488(.A(men_men_n1516_), .B(men_men_n1514_), .Y(men_men_n1517_));
  NA2        u1489(.A(men_men_n1434_), .B(men_men_n1509_), .Y(men_men_n1518_));
  NO2        u1490(.A(men_men_n309_), .B(c), .Y(men_men_n1519_));
  NA2        u1491(.A(men_men_n1519_), .B(men_men_n568_), .Y(men_men_n1520_));
  NA4        u1492(.A(men_men_n1520_), .B(men_men_n1518_), .C(men_men_n1517_), .D(men_men_n1513_), .Y(men_men_n1521_));
  NO3        u1493(.A(men_men_n1521_), .B(men_men_n1511_), .C(men_men_n1507_), .Y(men_men_n1522_));
  NA4        u1494(.A(men_men_n1522_), .B(men_men_n1502_), .C(men_men_n1488_), .D(men_men_n1482_), .Y(men_men_n1523_));
  OAI220     u1495(.A0(men_men_n486_), .A1(men_men_n309_), .B0(men_men_n136_), .B1(men_men_n59_), .Y(men_men_n1524_));
  NA2        u1496(.A(men_men_n1524_), .B(men_men_n1412_), .Y(men_men_n1525_));
  OAI210     u1497(.A0(men_men_n1460_), .A1(men_men_n1400_), .B0(men_men_n920_), .Y(men_men_n1526_));
  NO2        u1498(.A(men_men_n1081_), .B(men_men_n137_), .Y(men_men_n1527_));
  NA2        u1499(.A(men_men_n1527_), .B(men_men_n650_), .Y(men_men_n1528_));
  NA3        u1500(.A(men_men_n1528_), .B(men_men_n1526_), .C(men_men_n1525_), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n1432_), .B(men_men_n1515_), .Y(men_men_n1530_));
  NO2        u1502(.A(men_men_n1530_), .B(m), .Y(men_men_n1531_));
  NA3        u1503(.A(men_men_n1133_), .B(men_men_n112_), .C(men_men_n228_), .Y(men_men_n1532_));
  OAI220     u1504(.A0(men_men_n157_), .A1(men_men_n187_), .B0(men_men_n469_), .B1(g), .Y(men_men_n1533_));
  OAI210     u1505(.A0(men_men_n1533_), .A1(men_men_n114_), .B0(men_men_n1441_), .Y(men_men_n1534_));
  NA2        u1506(.A(men_men_n1534_), .B(men_men_n1532_), .Y(men_men_n1535_));
  NO3        u1507(.A(men_men_n1535_), .B(men_men_n1531_), .C(men_men_n1529_), .Y(men_men_n1536_));
  NO2        u1508(.A(men_men_n1399_), .B(e), .Y(men_men_n1537_));
  NA2        u1509(.A(men_men_n1537_), .B(men_men_n422_), .Y(men_men_n1538_));
  OR3        u1510(.A(men_men_n1498_), .B(men_men_n1258_), .C(men_men_n137_), .Y(men_men_n1539_));
  NO2        u1511(.A(men_men_n1539_), .B(men_men_n1538_), .Y(men_men_n1540_));
  NO3        u1512(.A(men_men_n1470_), .B(men_men_n368_), .C(a), .Y(men_men_n1541_));
  NO2        u1513(.A(men_men_n1541_), .B(men_men_n1540_), .Y(men_men_n1542_));
  NA2        u1514(.A(men_men_n566_), .B(g), .Y(men_men_n1543_));
  NA2        u1515(.A(men_men_n1543_), .B(men_men_n1429_), .Y(men_men_n1544_));
  NO2        u1516(.A(men_men_n1463_), .B(f), .Y(men_men_n1545_));
  AOI210     u1517(.A0(men_men_n1164_), .A1(a), .B0(men_men_n1545_), .Y(men_men_n1546_));
  OAI220     u1518(.A0(men_men_n1546_), .A1(men_men_n69_), .B0(men_men_n1544_), .B1(men_men_n220_), .Y(men_men_n1547_));
  NA2        u1519(.A(men_men_n1545_), .B(men_men_n1409_), .Y(men_men_n1548_));
  NO2        u1520(.A(men_men_n1548_), .B(men_men_n49_), .Y(men_men_n1549_));
  NA4        u1521(.A(men_men_n1133_), .B(men_men_n1131_), .C(men_men_n228_), .D(men_men_n68_), .Y(men_men_n1550_));
  NO2        u1522(.A(men_men_n49_), .B(l), .Y(men_men_n1551_));
  INV        u1523(.A(men_men_n504_), .Y(men_men_n1552_));
  NA2        u1524(.A(men_men_n1552_), .B(men_men_n1551_), .Y(men_men_n1553_));
  NO2        u1525(.A(men_men_n258_), .B(g), .Y(men_men_n1554_));
  NO2        u1526(.A(m), .B(i), .Y(men_men_n1555_));
  AOI220     u1527(.A0(men_men_n1555_), .A1(men_men_n1431_), .B0(men_men_n1114_), .B1(men_men_n1554_), .Y(men_men_n1556_));
  NA3        u1528(.A(men_men_n1556_), .B(men_men_n1553_), .C(men_men_n1550_), .Y(men_men_n1557_));
  NO3        u1529(.A(men_men_n1557_), .B(men_men_n1549_), .C(men_men_n1547_), .Y(men_men_n1558_));
  NA3        u1530(.A(men_men_n1558_), .B(men_men_n1542_), .C(men_men_n1536_), .Y(men_men_n1559_));
  NA3        u1531(.A(men_men_n998_), .B(men_men_n144_), .C(men_men_n46_), .Y(men_men_n1560_));
  AOI210     u1532(.A0(men_men_n155_), .A1(c), .B0(men_men_n1560_), .Y(men_men_n1561_));
  OAI210     u1533(.A0(men_men_n611_), .A1(g), .B0(men_men_n191_), .Y(men_men_n1562_));
  NA2        u1534(.A(men_men_n1562_), .B(men_men_n1505_), .Y(men_men_n1563_));
  AO210      u1535(.A0(men_men_n138_), .A1(l), .B0(men_men_n1453_), .Y(men_men_n1564_));
  NO2        u1536(.A(men_men_n72_), .B(c), .Y(men_men_n1565_));
  NO4        u1537(.A(men_men_n1417_), .B(men_men_n192_), .C(men_men_n469_), .D(men_men_n45_), .Y(men_men_n1566_));
  AOI210     u1538(.A0(men_men_n1514_), .A1(men_men_n1565_), .B0(men_men_n1566_), .Y(men_men_n1567_));
  NA3        u1539(.A(men_men_n1567_), .B(men_men_n1564_), .C(men_men_n1563_), .Y(men_men_n1568_));
  NO2        u1540(.A(men_men_n1568_), .B(men_men_n1561_), .Y(men_men_n1569_));
  NO4        u1541(.A(men_men_n232_), .B(men_men_n192_), .C(men_men_n262_), .D(k), .Y(men_men_n1570_));
  NO2        u1542(.A(men_men_n1560_), .B(men_men_n114_), .Y(men_men_n1571_));
  NOi21      u1543(.An(men_men_n1401_), .B(e), .Y(men_men_n1572_));
  NO3        u1544(.A(men_men_n1572_), .B(men_men_n1571_), .C(men_men_n1570_), .Y(men_men_n1573_));
  AN2        u1545(.A(men_men_n1133_), .B(men_men_n1121_), .Y(men_men_n1574_));
  AOI220     u1546(.A0(men_men_n1555_), .A1(men_men_n671_), .B0(men_men_n1098_), .B1(men_men_n166_), .Y(men_men_n1575_));
  NOi31      u1547(.An(men_men_n30_), .B(men_men_n1575_), .C(n), .Y(men_men_n1576_));
  AOI210     u1548(.A0(men_men_n1574_), .A1(men_men_n1211_), .B0(men_men_n1576_), .Y(men_men_n1577_));
  NO2        u1549(.A(men_men_n1508_), .B(men_men_n69_), .Y(men_men_n1578_));
  NA2        u1550(.A(men_men_n59_), .B(a), .Y(men_men_n1579_));
  NO2        u1551(.A(men_men_n1408_), .B(men_men_n122_), .Y(men_men_n1580_));
  OAI220     u1552(.A0(men_men_n1580_), .A1(men_men_n1453_), .B0(men_men_n1471_), .B1(men_men_n1579_), .Y(men_men_n1581_));
  NO2        u1553(.A(men_men_n1581_), .B(men_men_n1578_), .Y(men_men_n1582_));
  NA4        u1554(.A(men_men_n1582_), .B(men_men_n1577_), .C(men_men_n1573_), .D(men_men_n1569_), .Y(men_men_n1583_));
  OR4        u1555(.A(men_men_n1583_), .B(men_men_n1559_), .C(men_men_n1523_), .D(men_men_n1475_), .Y(men04));
  NOi31      u1556(.An(men_men_n1460_), .B(men_men_n1461_), .C(men_men_n1086_), .Y(men_men_n1585_));
  NO4        u1557(.A(men_men_n278_), .B(men_men_n1077_), .C(men_men_n505_), .D(j), .Y(men_men_n1586_));
  OR3        u1558(.A(men_men_n1586_), .B(men_men_n1585_), .C(men_men_n1104_), .Y(men_men_n1587_));
  NO3        u1559(.A(men_men_n1409_), .B(men_men_n93_), .C(k), .Y(men_men_n1588_));
  AOI210     u1560(.A0(men_men_n1588_), .A1(men_men_n1097_), .B0(men_men_n1232_), .Y(men_men_n1589_));
  NA2        u1561(.A(men_men_n1589_), .B(men_men_n1262_), .Y(men_men_n1590_));
  NO4        u1562(.A(men_men_n1590_), .B(men_men_n1587_), .C(men_men_n1112_), .D(men_men_n1091_), .Y(men_men_n1591_));
  NA4        u1563(.A(men_men_n1591_), .B(men_men_n1166_), .C(men_men_n1151_), .D(men_men_n1138_), .Y(men05));
  INV        u1564(.A(men_men_n556_), .Y(men_men_n1595_));
  INV        u1565(.A(men_men_n141_), .Y(men_men_n1596_));
  INV        u1566(.A(men_men_n723_), .Y(men_men_n1597_));
  INV        u1567(.A(men_men_n1397_), .Y(men_men_n1598_));
  INV        u1568(.A(f), .Y(men_men_n1599_));
  INV        u1569(.A(men_men_n479_), .Y(men_men_n1600_));
  INV        u1570(.A(k), .Y(men_men_n1601_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule