library verilog;
use verilog.vl_types.all;
entity sum_difabs_vlg_vec_tst is
end sum_difabs_vlg_vec_tst;
