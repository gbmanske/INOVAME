// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n141_, new_new_n143_,
    new_new_n144_, new_new_n145_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n737_, new_new_n738_,
    new_new_n739_, new_new_n740_, new_new_n741_, new_new_n742_,
    new_new_n743_, new_new_n744_, new_new_n745_, new_new_n746_,
    new_new_n747_, new_new_n748_, new_new_n749_, new_new_n750_,
    new_new_n751_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n786_, new_new_n787_,
    new_new_n788_, new_new_n789_, new_new_n790_, new_new_n791_,
    new_new_n792_, new_new_n793_, new_new_n794_, new_new_n795_,
    new_new_n796_, new_new_n797_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1048_, new_new_n1049_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(mai1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NO2        g0033(.A(new_new_n55_), .B(new_new_n54_), .Y(new_new_n56_));
  NA2        g0034(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n57_));
  NA3        g0035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n58_));
  NO2        g0036(.A(i_1_), .B(i_6_), .Y(new_new_n59_));
  NA2        g0037(.A(i_8_), .B(i_7_), .Y(new_new_n60_));
  OAI210     g0038(.A0(new_new_n60_), .A1(new_new_n59_), .B0(new_new_n58_), .Y(new_new_n61_));
  NA2        g0039(.A(new_new_n61_), .B(i_12_), .Y(new_new_n62_));
  NAi21      g0040(.An(i_2_), .B(i_7_), .Y(new_new_n63_));
  INV        g0041(.A(i_1_), .Y(new_new_n64_));
  NA2        g0042(.A(new_new_n64_), .B(i_6_), .Y(new_new_n65_));
  NA3        g0043(.A(new_new_n65_), .B(new_new_n63_), .C(new_new_n31_), .Y(new_new_n66_));
  NA2        g0044(.A(i_1_), .B(i_10_), .Y(new_new_n67_));
  NO2        g0045(.A(new_new_n67_), .B(i_6_), .Y(new_new_n68_));
  NAi31      g0046(.An(new_new_n68_), .B(new_new_n66_), .C(new_new_n62_), .Y(new_new_n69_));
  NA2        g0047(.A(new_new_n51_), .B(i_2_), .Y(new_new_n70_));
  AOI210     g0048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n71_));
  NA2        g0049(.A(i_1_), .B(i_6_), .Y(new_new_n72_));
  NO2        g0050(.A(new_new_n72_), .B(new_new_n25_), .Y(new_new_n73_));
  INV        g0051(.A(i_0_), .Y(new_new_n74_));
  NAi21      g0052(.An(i_5_), .B(i_10_), .Y(new_new_n75_));
  NA2        g0053(.A(i_5_), .B(i_9_), .Y(new_new_n76_));
  AOI210     g0054(.A0(new_new_n76_), .A1(new_new_n75_), .B0(new_new_n74_), .Y(new_new_n77_));
  NO2        g0055(.A(new_new_n77_), .B(new_new_n73_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n71_), .A1(new_new_n70_), .B0(new_new_n78_), .Y(new_new_n79_));
  OAI210     g0057(.A0(new_new_n79_), .A1(new_new_n69_), .B0(i_0_), .Y(new_new_n80_));
  NA2        g0058(.A(i_12_), .B(i_5_), .Y(new_new_n81_));
  NA2        g0059(.A(i_2_), .B(i_8_), .Y(new_new_n82_));
  NO2        g0060(.A(new_new_n82_), .B(new_new_n59_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_9_), .Y(new_new_n84_));
  NO2        g0062(.A(i_3_), .B(i_7_), .Y(new_new_n85_));
  NO3        g0063(.A(new_new_n85_), .B(new_new_n84_), .C(new_new_n64_), .Y(new_new_n86_));
  INV        g0064(.A(i_6_), .Y(new_new_n87_));
  OR4        g0065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n88_));
  INV        g0066(.A(new_new_n88_), .Y(new_new_n89_));
  NO2        g0067(.A(i_2_), .B(i_7_), .Y(new_new_n90_));
  NO2        g0068(.A(new_new_n89_), .B(new_new_n90_), .Y(new_new_n91_));
  OAI210     g0069(.A0(new_new_n86_), .A1(new_new_n83_), .B0(new_new_n91_), .Y(new_new_n92_));
  NAi21      g0070(.An(i_6_), .B(i_10_), .Y(new_new_n93_));
  NA2        g0071(.A(i_6_), .B(i_9_), .Y(new_new_n94_));
  AOI210     g0072(.A0(new_new_n94_), .A1(new_new_n93_), .B0(new_new_n64_), .Y(new_new_n95_));
  NA2        g0073(.A(i_2_), .B(i_6_), .Y(new_new_n96_));
  NO3        g0074(.A(new_new_n96_), .B(new_new_n50_), .C(new_new_n25_), .Y(new_new_n97_));
  NO2        g0075(.A(new_new_n97_), .B(new_new_n95_), .Y(new_new_n98_));
  AOI210     g0076(.A0(new_new_n98_), .A1(new_new_n92_), .B0(new_new_n81_), .Y(new_new_n99_));
  AN3        g0077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n100_));
  NAi21      g0078(.An(i_6_), .B(i_11_), .Y(new_new_n101_));
  NO2        g0079(.A(i_5_), .B(i_8_), .Y(new_new_n102_));
  NOi21      g0080(.An(new_new_n102_), .B(new_new_n101_), .Y(new_new_n103_));
  AOI220     g0081(.A0(new_new_n103_), .A1(new_new_n63_), .B0(new_new_n100_), .B1(new_new_n32_), .Y(new_new_n104_));
  INV        g0082(.A(i_7_), .Y(new_new_n105_));
  NA2        g0083(.A(new_new_n47_), .B(new_new_n105_), .Y(new_new_n106_));
  NO2        g0084(.A(i_0_), .B(i_5_), .Y(new_new_n107_));
  NO2        g0085(.A(new_new_n107_), .B(new_new_n87_), .Y(new_new_n108_));
  NA2        g0086(.A(i_12_), .B(i_3_), .Y(new_new_n109_));
  INV        g0087(.A(new_new_n109_), .Y(new_new_n110_));
  NA3        g0088(.A(new_new_n110_), .B(new_new_n108_), .C(new_new_n106_), .Y(new_new_n111_));
  NAi21      g0089(.An(i_7_), .B(i_11_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n93_), .C(new_new_n54_), .Y(new_new_n113_));
  AN2        g0091(.A(i_2_), .B(i_10_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n114_), .B(i_7_), .Y(new_new_n115_));
  OR2        g0093(.A(new_new_n81_), .B(new_new_n59_), .Y(new_new_n116_));
  NO2        g0094(.A(i_8_), .B(new_new_n105_), .Y(new_new_n117_));
  NO3        g0095(.A(new_new_n117_), .B(new_new_n116_), .C(new_new_n115_), .Y(new_new_n118_));
  NA2        g0096(.A(i_12_), .B(i_7_), .Y(new_new_n119_));
  NO2        g0097(.A(new_new_n64_), .B(new_new_n26_), .Y(new_new_n120_));
  NA2        g0098(.A(new_new_n120_), .B(i_0_), .Y(new_new_n121_));
  NA2        g0099(.A(i_11_), .B(i_12_), .Y(new_new_n122_));
  OAI210     g0100(.A0(new_new_n121_), .A1(new_new_n119_), .B0(new_new_n122_), .Y(new_new_n123_));
  NO2        g0101(.A(new_new_n123_), .B(new_new_n118_), .Y(new_new_n124_));
  NAi41      g0102(.An(new_new_n113_), .B(new_new_n124_), .C(new_new_n111_), .D(new_new_n104_), .Y(new_new_n125_));
  NOi21      g0103(.An(i_1_), .B(i_5_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n126_), .B(i_11_), .Y(new_new_n127_));
  NA2        g0105(.A(new_new_n105_), .B(new_new_n37_), .Y(new_new_n128_));
  NA2        g0106(.A(i_7_), .B(new_new_n25_), .Y(new_new_n129_));
  NA2        g0107(.A(new_new_n129_), .B(new_new_n128_), .Y(new_new_n130_));
  NO2        g0108(.A(new_new_n130_), .B(new_new_n47_), .Y(new_new_n131_));
  NA2        g0109(.A(new_new_n94_), .B(new_new_n93_), .Y(new_new_n132_));
  NAi21      g0110(.An(i_3_), .B(i_8_), .Y(new_new_n133_));
  NA2        g0111(.A(new_new_n133_), .B(new_new_n63_), .Y(new_new_n134_));
  NOi31      g0112(.An(new_new_n134_), .B(new_new_n132_), .C(new_new_n131_), .Y(new_new_n135_));
  NO2        g0113(.A(i_1_), .B(new_new_n87_), .Y(new_new_n136_));
  NO2        g0114(.A(i_6_), .B(i_5_), .Y(new_new_n137_));
  NA2        g0115(.A(new_new_n137_), .B(i_3_), .Y(new_new_n138_));
  AO210      g0116(.A0(new_new_n138_), .A1(new_new_n48_), .B0(new_new_n136_), .Y(new_new_n139_));
  OAI220     g0117(.A0(new_new_n139_), .A1(new_new_n112_), .B0(new_new_n135_), .B1(new_new_n127_), .Y(new_new_n140_));
  NO3        g0118(.A(new_new_n140_), .B(new_new_n125_), .C(new_new_n99_), .Y(new_new_n141_));
  NA3        g0119(.A(new_new_n141_), .B(new_new_n80_), .C(new_new_n57_), .Y(mai2));
  NO2        g0120(.A(new_new_n64_), .B(new_new_n37_), .Y(new_new_n143_));
  NA2        g0121(.A(i_6_), .B(new_new_n25_), .Y(new_new_n144_));
  NA2        g0122(.A(new_new_n144_), .B(new_new_n143_), .Y(new_new_n145_));
  NA4        g0123(.A(new_new_n145_), .B(new_new_n78_), .C(new_new_n70_), .D(new_new_n30_), .Y(mai0));
  AN2        g0124(.A(i_8_), .B(i_7_), .Y(new_new_n147_));
  NA2        g0125(.A(new_new_n147_), .B(i_6_), .Y(new_new_n148_));
  NO2        g0126(.A(i_12_), .B(i_13_), .Y(new_new_n149_));
  NAi21      g0127(.An(i_5_), .B(i_11_), .Y(new_new_n150_));
  NOi21      g0128(.An(new_new_n149_), .B(new_new_n150_), .Y(new_new_n151_));
  NO2        g0129(.A(i_0_), .B(i_1_), .Y(new_new_n152_));
  NA2        g0130(.A(i_2_), .B(i_3_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n153_), .B(i_4_), .Y(new_new_n154_));
  NA3        g0132(.A(new_new_n154_), .B(new_new_n152_), .C(new_new_n151_), .Y(new_new_n155_));
  OR2        g0133(.A(new_new_n155_), .B(new_new_n25_), .Y(new_new_n156_));
  AN2        g0134(.A(new_new_n149_), .B(new_new_n84_), .Y(new_new_n157_));
  NO2        g0135(.A(new_new_n157_), .B(new_new_n27_), .Y(new_new_n158_));
  NA2        g0136(.A(i_1_), .B(i_5_), .Y(new_new_n159_));
  NO2        g0137(.A(new_new_n74_), .B(new_new_n47_), .Y(new_new_n160_));
  NA2        g0138(.A(new_new_n160_), .B(new_new_n36_), .Y(new_new_n161_));
  NO3        g0139(.A(new_new_n161_), .B(new_new_n159_), .C(new_new_n158_), .Y(new_new_n162_));
  OR2        g0140(.A(i_0_), .B(i_1_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n163_), .B(new_new_n81_), .C(i_13_), .Y(new_new_n164_));
  NAi32      g0142(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n165_));
  NAi21      g0143(.An(new_new_n165_), .B(new_new_n164_), .Y(new_new_n166_));
  NOi21      g0144(.An(i_4_), .B(i_10_), .Y(new_new_n167_));
  NA2        g0145(.A(new_new_n167_), .B(new_new_n40_), .Y(new_new_n168_));
  NO2        g0146(.A(i_3_), .B(i_5_), .Y(new_new_n169_));
  INV        g0147(.A(new_new_n162_), .Y(new_new_n170_));
  AOI210     g0148(.A0(new_new_n170_), .A1(new_new_n156_), .B0(new_new_n148_), .Y(new_new_n171_));
  NA3        g0149(.A(new_new_n74_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n172_));
  NA2        g0150(.A(i_3_), .B(new_new_n49_), .Y(new_new_n173_));
  NOi21      g0151(.An(i_4_), .B(i_9_), .Y(new_new_n174_));
  NOi21      g0152(.An(i_11_), .B(i_13_), .Y(new_new_n175_));
  NA2        g0153(.A(new_new_n175_), .B(new_new_n174_), .Y(new_new_n176_));
  OR2        g0154(.A(new_new_n176_), .B(new_new_n173_), .Y(new_new_n177_));
  NO2        g0155(.A(i_4_), .B(i_5_), .Y(new_new_n178_));
  NAi21      g0156(.An(i_12_), .B(i_11_), .Y(new_new_n179_));
  NO2        g0157(.A(new_new_n179_), .B(i_13_), .Y(new_new_n180_));
  NA3        g0158(.A(new_new_n180_), .B(new_new_n178_), .C(new_new_n84_), .Y(new_new_n181_));
  AOI210     g0159(.A0(new_new_n181_), .A1(new_new_n177_), .B0(new_new_n172_), .Y(new_new_n182_));
  NO2        g0160(.A(new_new_n74_), .B(new_new_n64_), .Y(new_new_n183_));
  NA2        g0161(.A(new_new_n183_), .B(new_new_n47_), .Y(new_new_n184_));
  NA2        g0162(.A(new_new_n36_), .B(i_5_), .Y(new_new_n185_));
  NA2        g0163(.A(i_3_), .B(i_5_), .Y(new_new_n186_));
  NO2        g0164(.A(new_new_n74_), .B(i_5_), .Y(new_new_n187_));
  NO2        g0165(.A(i_13_), .B(i_10_), .Y(new_new_n188_));
  NA3        g0166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n45_), .Y(new_new_n189_));
  NO2        g0167(.A(i_2_), .B(i_1_), .Y(new_new_n190_));
  NA2        g0168(.A(new_new_n190_), .B(i_3_), .Y(new_new_n191_));
  NAi21      g0169(.An(i_4_), .B(i_12_), .Y(new_new_n192_));
  NO4        g0170(.A(new_new_n192_), .B(new_new_n191_), .C(new_new_n189_), .D(new_new_n25_), .Y(new_new_n193_));
  NO2        g0171(.A(new_new_n193_), .B(new_new_n182_), .Y(new_new_n194_));
  INV        g0172(.A(i_8_), .Y(new_new_n195_));
  NO2        g0173(.A(new_new_n195_), .B(i_7_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(i_6_), .Y(new_new_n197_));
  NO3        g0175(.A(i_3_), .B(new_new_n87_), .C(new_new_n49_), .Y(new_new_n198_));
  NA2        g0176(.A(new_new_n198_), .B(new_new_n117_), .Y(new_new_n199_));
  NO3        g0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n200_));
  NA3        g0178(.A(new_new_n200_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n201_));
  NO3        g0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n202_));
  OAI210     g0180(.A0(new_new_n100_), .A1(i_12_), .B0(new_new_n202_), .Y(new_new_n203_));
  AOI210     g0181(.A0(new_new_n203_), .A1(new_new_n201_), .B0(new_new_n199_), .Y(new_new_n204_));
  NO2        g0182(.A(i_3_), .B(i_8_), .Y(new_new_n205_));
  NO3        g0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n206_));
  NA3        g0184(.A(new_new_n206_), .B(new_new_n205_), .C(new_new_n40_), .Y(new_new_n207_));
  NO2        g0185(.A(new_new_n107_), .B(new_new_n59_), .Y(new_new_n208_));
  INV        g0186(.A(new_new_n208_), .Y(new_new_n209_));
  NO2        g0187(.A(i_13_), .B(i_9_), .Y(new_new_n210_));
  NA3        g0188(.A(new_new_n210_), .B(i_6_), .C(new_new_n195_), .Y(new_new_n211_));
  NAi21      g0189(.An(i_12_), .B(i_3_), .Y(new_new_n212_));
  OR2        g0190(.A(new_new_n212_), .B(new_new_n211_), .Y(new_new_n213_));
  NO2        g0191(.A(new_new_n45_), .B(i_5_), .Y(new_new_n214_));
  NO3        g0192(.A(i_0_), .B(i_2_), .C(new_new_n64_), .Y(new_new_n215_));
  NA3        g0193(.A(new_new_n215_), .B(new_new_n214_), .C(i_10_), .Y(new_new_n216_));
  OAI220     g0194(.A0(new_new_n216_), .A1(new_new_n213_), .B0(new_new_n209_), .B1(new_new_n207_), .Y(new_new_n217_));
  AOI210     g0195(.A0(new_new_n217_), .A1(i_7_), .B0(new_new_n204_), .Y(new_new_n218_));
  OAI220     g0196(.A0(new_new_n218_), .A1(i_4_), .B0(new_new_n197_), .B1(new_new_n194_), .Y(new_new_n219_));
  NAi21      g0197(.An(i_12_), .B(i_7_), .Y(new_new_n220_));
  NA3        g0198(.A(i_13_), .B(new_new_n195_), .C(i_10_), .Y(new_new_n221_));
  NO2        g0199(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n222_));
  NA2        g0200(.A(i_0_), .B(i_5_), .Y(new_new_n223_));
  NA2        g0201(.A(new_new_n223_), .B(new_new_n108_), .Y(new_new_n224_));
  OAI220     g0202(.A0(new_new_n224_), .A1(new_new_n191_), .B0(new_new_n184_), .B1(new_new_n138_), .Y(new_new_n225_));
  NAi31      g0203(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n226_));
  NO2        g0204(.A(new_new_n36_), .B(i_13_), .Y(new_new_n227_));
  NO2        g0205(.A(new_new_n74_), .B(new_new_n26_), .Y(new_new_n228_));
  NO2        g0206(.A(new_new_n47_), .B(new_new_n64_), .Y(new_new_n229_));
  INV        g0207(.A(i_13_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n230_), .Y(new_new_n231_));
  NA2        g0209(.A(new_new_n225_), .B(new_new_n222_), .Y(new_new_n232_));
  NO2        g0210(.A(i_12_), .B(new_new_n37_), .Y(new_new_n233_));
  NO2        g0211(.A(new_new_n186_), .B(i_4_), .Y(new_new_n234_));
  NA2        g0212(.A(new_new_n234_), .B(new_new_n233_), .Y(new_new_n235_));
  OR2        g0213(.A(i_8_), .B(i_7_), .Y(new_new_n236_));
  NO2        g0214(.A(new_new_n236_), .B(new_new_n87_), .Y(new_new_n237_));
  NO2        g0215(.A(new_new_n54_), .B(i_1_), .Y(new_new_n238_));
  NA2        g0216(.A(new_new_n238_), .B(new_new_n237_), .Y(new_new_n239_));
  INV        g0217(.A(i_12_), .Y(new_new_n240_));
  NO2        g0218(.A(new_new_n45_), .B(new_new_n240_), .Y(new_new_n241_));
  NO3        g0219(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n242_));
  NA2        g0220(.A(i_2_), .B(i_1_), .Y(new_new_n243_));
  NO2        g0221(.A(new_new_n239_), .B(new_new_n235_), .Y(new_new_n244_));
  NO3        g0222(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n245_));
  NAi21      g0223(.An(i_4_), .B(i_3_), .Y(new_new_n246_));
  NO2        g0224(.A(i_0_), .B(i_6_), .Y(new_new_n247_));
  NOi41      g0225(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n248_));
  NA2        g0226(.A(new_new_n248_), .B(new_new_n247_), .Y(new_new_n249_));
  NO2        g0227(.A(new_new_n243_), .B(new_new_n186_), .Y(new_new_n250_));
  NAi21      g0228(.An(new_new_n249_), .B(new_new_n250_), .Y(new_new_n251_));
  INV        g0229(.A(new_new_n251_), .Y(new_new_n252_));
  AOI220     g0230(.A0(new_new_n252_), .A1(new_new_n40_), .B0(new_new_n244_), .B1(new_new_n210_), .Y(new_new_n253_));
  NO2        g0231(.A(i_11_), .B(new_new_n230_), .Y(new_new_n254_));
  NOi21      g0232(.An(i_1_), .B(i_6_), .Y(new_new_n255_));
  NAi21      g0233(.An(i_3_), .B(i_7_), .Y(new_new_n256_));
  NA2        g0234(.A(new_new_n240_), .B(i_9_), .Y(new_new_n257_));
  OR4        g0235(.A(new_new_n257_), .B(new_new_n256_), .C(new_new_n255_), .D(new_new_n187_), .Y(new_new_n258_));
  NO2        g0236(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n259_));
  NO2        g0237(.A(i_12_), .B(i_3_), .Y(new_new_n260_));
  NA2        g0238(.A(new_new_n74_), .B(i_5_), .Y(new_new_n261_));
  NA2        g0239(.A(i_3_), .B(i_9_), .Y(new_new_n262_));
  NAi21      g0240(.An(i_7_), .B(i_10_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n263_), .B(new_new_n262_), .Y(new_new_n264_));
  NA3        g0242(.A(new_new_n264_), .B(new_new_n261_), .C(new_new_n65_), .Y(new_new_n265_));
  NA2        g0243(.A(new_new_n265_), .B(new_new_n258_), .Y(new_new_n266_));
  NA3        g0244(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n267_));
  INV        g0245(.A(new_new_n148_), .Y(new_new_n268_));
  NA2        g0246(.A(new_new_n240_), .B(i_13_), .Y(new_new_n269_));
  NO2        g0247(.A(new_new_n269_), .B(new_new_n76_), .Y(new_new_n270_));
  AOI220     g0248(.A0(new_new_n270_), .A1(new_new_n268_), .B0(new_new_n266_), .B1(new_new_n254_), .Y(new_new_n271_));
  NO2        g0249(.A(new_new_n236_), .B(new_new_n37_), .Y(new_new_n272_));
  NA2        g0250(.A(i_12_), .B(i_6_), .Y(new_new_n273_));
  OR2        g0251(.A(i_13_), .B(i_9_), .Y(new_new_n274_));
  NO3        g0252(.A(new_new_n274_), .B(new_new_n273_), .C(new_new_n49_), .Y(new_new_n275_));
  NO2        g0253(.A(new_new_n246_), .B(i_2_), .Y(new_new_n276_));
  NA3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n45_), .Y(new_new_n277_));
  NA2        g0255(.A(new_new_n254_), .B(i_9_), .Y(new_new_n278_));
  NA2        g0256(.A(new_new_n261_), .B(new_new_n65_), .Y(new_new_n279_));
  OAI210     g0257(.A0(new_new_n279_), .A1(new_new_n278_), .B0(new_new_n277_), .Y(new_new_n280_));
  NO3        g0258(.A(i_11_), .B(new_new_n230_), .C(new_new_n25_), .Y(new_new_n281_));
  NO2        g0259(.A(new_new_n256_), .B(i_8_), .Y(new_new_n282_));
  NO2        g0260(.A(i_6_), .B(new_new_n49_), .Y(new_new_n283_));
  NA2        g0261(.A(new_new_n280_), .B(new_new_n272_), .Y(new_new_n284_));
  NA4        g0262(.A(new_new_n284_), .B(new_new_n271_), .C(new_new_n253_), .D(new_new_n232_), .Y(new_new_n285_));
  NO3        g0263(.A(i_12_), .B(new_new_n230_), .C(new_new_n37_), .Y(new_new_n286_));
  INV        g0264(.A(new_new_n286_), .Y(new_new_n287_));
  NO3        g0265(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n288_));
  NO2        g0266(.A(new_new_n243_), .B(i_0_), .Y(new_new_n289_));
  NA2        g0267(.A(i_0_), .B(i_1_), .Y(new_new_n290_));
  NO2        g0268(.A(new_new_n290_), .B(i_2_), .Y(new_new_n291_));
  NO2        g0269(.A(new_new_n60_), .B(i_6_), .Y(new_new_n292_));
  NA3        g0270(.A(new_new_n292_), .B(new_new_n291_), .C(new_new_n169_), .Y(new_new_n293_));
  NO2        g0271(.A(i_3_), .B(i_10_), .Y(new_new_n294_));
  NA3        g0272(.A(new_new_n294_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n295_));
  NO2        g0273(.A(i_2_), .B(new_new_n105_), .Y(new_new_n296_));
  NA2        g0274(.A(i_1_), .B(new_new_n36_), .Y(new_new_n297_));
  NO2        g0275(.A(new_new_n297_), .B(i_8_), .Y(new_new_n298_));
  NOi21      g0276(.An(new_new_n223_), .B(new_new_n107_), .Y(new_new_n299_));
  NA3        g0277(.A(new_new_n299_), .B(new_new_n298_), .C(new_new_n296_), .Y(new_new_n300_));
  AN2        g0278(.A(i_3_), .B(i_10_), .Y(new_new_n301_));
  NA4        g0279(.A(new_new_n301_), .B(new_new_n200_), .C(new_new_n180_), .D(new_new_n178_), .Y(new_new_n302_));
  NO2        g0280(.A(i_5_), .B(new_new_n37_), .Y(new_new_n303_));
  NO2        g0281(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n304_));
  OR2        g0282(.A(new_new_n300_), .B(new_new_n295_), .Y(new_new_n305_));
  OAI220     g0283(.A0(new_new_n305_), .A1(i_6_), .B0(new_new_n293_), .B1(new_new_n287_), .Y(new_new_n306_));
  NO4        g0284(.A(new_new_n306_), .B(new_new_n285_), .C(new_new_n219_), .D(new_new_n171_), .Y(new_new_n307_));
  NO3        g0285(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n308_));
  NO2        g0286(.A(new_new_n60_), .B(new_new_n87_), .Y(new_new_n309_));
  NO3        g0287(.A(i_6_), .B(new_new_n195_), .C(i_7_), .Y(new_new_n310_));
  NO2        g0288(.A(i_2_), .B(i_3_), .Y(new_new_n311_));
  OR2        g0289(.A(i_0_), .B(i_5_), .Y(new_new_n312_));
  NA2        g0290(.A(new_new_n223_), .B(new_new_n312_), .Y(new_new_n313_));
  NA4        g0291(.A(new_new_n313_), .B(new_new_n237_), .C(new_new_n311_), .D(i_1_), .Y(new_new_n314_));
  NAi21      g0292(.An(i_8_), .B(i_7_), .Y(new_new_n315_));
  NO2        g0293(.A(new_new_n315_), .B(i_6_), .Y(new_new_n316_));
  NO2        g0294(.A(new_new_n163_), .B(new_new_n47_), .Y(new_new_n317_));
  NA3        g0295(.A(new_new_n317_), .B(new_new_n316_), .C(new_new_n169_), .Y(new_new_n318_));
  NA2        g0296(.A(new_new_n318_), .B(new_new_n314_), .Y(new_new_n319_));
  NA2        g0297(.A(new_new_n319_), .B(i_4_), .Y(new_new_n320_));
  NO2        g0298(.A(i_12_), .B(i_10_), .Y(new_new_n321_));
  NOi21      g0299(.An(i_5_), .B(i_0_), .Y(new_new_n322_));
  NA4        g0300(.A(new_new_n85_), .B(new_new_n36_), .C(new_new_n87_), .D(i_8_), .Y(new_new_n323_));
  NO2        g0301(.A(i_6_), .B(i_8_), .Y(new_new_n324_));
  NOi21      g0302(.An(i_0_), .B(i_2_), .Y(new_new_n325_));
  AN2        g0303(.A(new_new_n325_), .B(new_new_n324_), .Y(new_new_n326_));
  NO2        g0304(.A(i_1_), .B(i_7_), .Y(new_new_n327_));
  AO220      g0305(.A0(new_new_n327_), .A1(new_new_n326_), .B0(new_new_n316_), .B1(new_new_n238_), .Y(new_new_n328_));
  NA3        g0306(.A(new_new_n328_), .B(new_new_n42_), .C(i_5_), .Y(new_new_n329_));
  NA2        g0307(.A(new_new_n329_), .B(new_new_n320_), .Y(new_new_n330_));
  NO3        g0308(.A(new_new_n236_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n331_));
  NO3        g0309(.A(new_new_n315_), .B(i_2_), .C(i_1_), .Y(new_new_n332_));
  OAI210     g0310(.A0(new_new_n332_), .A1(new_new_n331_), .B0(i_6_), .Y(new_new_n333_));
  NA3        g0311(.A(new_new_n255_), .B(new_new_n296_), .C(new_new_n195_), .Y(new_new_n334_));
  AOI210     g0312(.A0(new_new_n334_), .A1(new_new_n333_), .B0(new_new_n313_), .Y(new_new_n335_));
  NOi21      g0313(.An(new_new_n159_), .B(new_new_n108_), .Y(new_new_n336_));
  NO2        g0314(.A(new_new_n336_), .B(new_new_n129_), .Y(new_new_n337_));
  OAI210     g0315(.A0(new_new_n337_), .A1(new_new_n335_), .B0(i_3_), .Y(new_new_n338_));
  INV        g0316(.A(new_new_n85_), .Y(new_new_n339_));
  NO2        g0317(.A(new_new_n290_), .B(new_new_n82_), .Y(new_new_n340_));
  NA2        g0318(.A(new_new_n340_), .B(new_new_n137_), .Y(new_new_n341_));
  NO2        g0319(.A(new_new_n96_), .B(new_new_n195_), .Y(new_new_n342_));
  NA3        g0320(.A(new_new_n299_), .B(new_new_n342_), .C(new_new_n64_), .Y(new_new_n343_));
  AOI210     g0321(.A0(new_new_n343_), .A1(new_new_n341_), .B0(new_new_n339_), .Y(new_new_n344_));
  NO2        g0322(.A(new_new_n195_), .B(i_9_), .Y(new_new_n345_));
  NA2        g0323(.A(new_new_n345_), .B(new_new_n208_), .Y(new_new_n346_));
  NO2        g0324(.A(new_new_n346_), .B(new_new_n47_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n347_), .B(new_new_n344_), .Y(new_new_n348_));
  AOI210     g0326(.A0(new_new_n348_), .A1(new_new_n338_), .B0(new_new_n168_), .Y(new_new_n349_));
  AOI210     g0327(.A0(new_new_n330_), .A1(new_new_n308_), .B0(new_new_n349_), .Y(new_new_n350_));
  NOi32      g0328(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n351_));
  INV        g0329(.A(new_new_n351_), .Y(new_new_n352_));
  NAi21      g0330(.An(i_0_), .B(i_6_), .Y(new_new_n353_));
  NAi21      g0331(.An(i_1_), .B(i_5_), .Y(new_new_n354_));
  NA2        g0332(.A(new_new_n354_), .B(new_new_n353_), .Y(new_new_n355_));
  NA2        g0333(.A(new_new_n355_), .B(new_new_n25_), .Y(new_new_n356_));
  OAI210     g0334(.A0(new_new_n356_), .A1(new_new_n165_), .B0(new_new_n249_), .Y(new_new_n357_));
  NAi41      g0335(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n358_));
  OAI220     g0336(.A0(new_new_n358_), .A1(new_new_n354_), .B0(new_new_n226_), .B1(new_new_n165_), .Y(new_new_n359_));
  AOI210     g0337(.A0(new_new_n358_), .A1(new_new_n165_), .B0(new_new_n163_), .Y(new_new_n360_));
  NOi32      g0338(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n361_));
  OR2        g0339(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n362_));
  NO2        g0340(.A(i_1_), .B(new_new_n105_), .Y(new_new_n363_));
  NAi21      g0341(.An(i_3_), .B(i_4_), .Y(new_new_n364_));
  NO2        g0342(.A(new_new_n364_), .B(i_9_), .Y(new_new_n365_));
  AN2        g0343(.A(i_6_), .B(i_7_), .Y(new_new_n366_));
  OAI210     g0344(.A0(new_new_n366_), .A1(new_new_n363_), .B0(new_new_n365_), .Y(new_new_n367_));
  NA2        g0345(.A(i_2_), .B(i_7_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n364_), .B(i_10_), .Y(new_new_n369_));
  NA3        g0347(.A(new_new_n369_), .B(new_new_n368_), .C(new_new_n247_), .Y(new_new_n370_));
  AOI210     g0348(.A0(new_new_n370_), .A1(new_new_n367_), .B0(new_new_n187_), .Y(new_new_n371_));
  AOI210     g0349(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n372_));
  OAI210     g0350(.A0(new_new_n372_), .A1(new_new_n190_), .B0(new_new_n369_), .Y(new_new_n373_));
  AOI220     g0351(.A0(new_new_n369_), .A1(new_new_n327_), .B0(new_new_n242_), .B1(new_new_n190_), .Y(new_new_n374_));
  AOI210     g0352(.A0(new_new_n374_), .A1(new_new_n373_), .B0(i_5_), .Y(new_new_n375_));
  NO4        g0353(.A(new_new_n375_), .B(new_new_n371_), .C(new_new_n362_), .D(new_new_n357_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n376_), .B(new_new_n352_), .Y(new_new_n377_));
  AN2        g0355(.A(i_12_), .B(i_5_), .Y(new_new_n378_));
  NO2        g0356(.A(i_4_), .B(new_new_n26_), .Y(new_new_n379_));
  NA2        g0357(.A(new_new_n379_), .B(new_new_n378_), .Y(new_new_n380_));
  NO2        g0358(.A(i_11_), .B(i_6_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n246_), .B(i_5_), .Y(new_new_n382_));
  NO2        g0360(.A(i_5_), .B(i_10_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n384_));
  NO3        g0362(.A(new_new_n87_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n385_));
  NO2        g0363(.A(i_3_), .B(new_new_n105_), .Y(new_new_n386_));
  NA4        g0364(.A(new_new_n294_), .B(new_new_n94_), .C(new_new_n76_), .D(new_new_n55_), .Y(new_new_n387_));
  NO2        g0365(.A(i_11_), .B(i_12_), .Y(new_new_n388_));
  NA2        g0366(.A(new_new_n388_), .B(new_new_n36_), .Y(new_new_n389_));
  NO2        g0367(.A(new_new_n387_), .B(new_new_n389_), .Y(new_new_n390_));
  NA3        g0368(.A(new_new_n117_), .B(new_new_n42_), .C(i_11_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n391_), .B(new_new_n226_), .Y(new_new_n392_));
  NAi21      g0370(.An(i_13_), .B(i_0_), .Y(new_new_n393_));
  NO2        g0371(.A(new_new_n393_), .B(new_new_n243_), .Y(new_new_n394_));
  OAI210     g0372(.A0(new_new_n392_), .A1(new_new_n390_), .B0(new_new_n394_), .Y(new_new_n395_));
  INV        g0373(.A(new_new_n395_), .Y(new_new_n396_));
  NA2        g0374(.A(new_new_n45_), .B(new_new_n230_), .Y(new_new_n397_));
  NO3        g0375(.A(i_1_), .B(i_12_), .C(new_new_n87_), .Y(new_new_n398_));
  NO2        g0376(.A(i_0_), .B(i_11_), .Y(new_new_n399_));
  INV        g0377(.A(i_5_), .Y(new_new_n400_));
  AN2        g0378(.A(i_1_), .B(i_6_), .Y(new_new_n401_));
  NOi21      g0379(.An(i_2_), .B(i_12_), .Y(new_new_n402_));
  NA2        g0380(.A(new_new_n402_), .B(new_new_n401_), .Y(new_new_n403_));
  NO2        g0381(.A(new_new_n403_), .B(new_new_n400_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n147_), .B(i_9_), .Y(new_new_n405_));
  NO2        g0383(.A(new_new_n405_), .B(i_4_), .Y(new_new_n406_));
  NA2        g0384(.A(new_new_n404_), .B(new_new_n406_), .Y(new_new_n407_));
  NAi21      g0385(.An(i_9_), .B(i_4_), .Y(new_new_n408_));
  OR2        g0386(.A(i_13_), .B(i_10_), .Y(new_new_n409_));
  NO3        g0387(.A(new_new_n409_), .B(new_new_n122_), .C(new_new_n408_), .Y(new_new_n410_));
  NO2        g0388(.A(new_new_n176_), .B(new_new_n128_), .Y(new_new_n411_));
  OR2        g0389(.A(new_new_n221_), .B(new_new_n220_), .Y(new_new_n412_));
  NO2        g0390(.A(new_new_n105_), .B(new_new_n25_), .Y(new_new_n413_));
  NA2        g0391(.A(new_new_n286_), .B(new_new_n413_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n283_), .B(new_new_n215_), .Y(new_new_n415_));
  OAI220     g0393(.A0(new_new_n415_), .A1(new_new_n412_), .B0(new_new_n414_), .B1(new_new_n336_), .Y(new_new_n416_));
  INV        g0394(.A(new_new_n416_), .Y(new_new_n417_));
  AOI210     g0395(.A0(new_new_n417_), .A1(new_new_n407_), .B0(new_new_n26_), .Y(new_new_n418_));
  INV        g0396(.A(new_new_n314_), .Y(new_new_n419_));
  AOI220     g0397(.A0(new_new_n292_), .A1(new_new_n288_), .B0(new_new_n289_), .B1(new_new_n309_), .Y(new_new_n420_));
  NO2        g0398(.A(new_new_n420_), .B(new_new_n173_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n186_), .B(new_new_n87_), .Y(new_new_n422_));
  NO2        g0400(.A(new_new_n421_), .B(new_new_n419_), .Y(new_new_n423_));
  NA2        g0401(.A(new_new_n195_), .B(i_10_), .Y(new_new_n424_));
  NA3        g0402(.A(new_new_n261_), .B(new_new_n65_), .C(i_2_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(new_new_n424_), .Y(new_new_n426_));
  NA2        g0404(.A(new_new_n310_), .B(new_new_n313_), .Y(new_new_n427_));
  NO2        g0405(.A(new_new_n427_), .B(new_new_n191_), .Y(new_new_n428_));
  NO2        g0406(.A(new_new_n428_), .B(new_new_n426_), .Y(new_new_n429_));
  AOI210     g0407(.A0(new_new_n429_), .A1(new_new_n423_), .B0(new_new_n278_), .Y(new_new_n430_));
  NO4        g0408(.A(new_new_n430_), .B(new_new_n418_), .C(new_new_n396_), .D(new_new_n377_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n64_), .B(i_4_), .Y(new_new_n432_));
  NO2        g0410(.A(new_new_n74_), .B(i_13_), .Y(new_new_n433_));
  NO2        g0411(.A(i_10_), .B(i_9_), .Y(new_new_n434_));
  NAi21      g0412(.An(i_12_), .B(i_8_), .Y(new_new_n435_));
  NO2        g0413(.A(new_new_n435_), .B(i_3_), .Y(new_new_n436_));
  NO2        g0414(.A(new_new_n47_), .B(i_4_), .Y(new_new_n437_));
  NA2        g0415(.A(new_new_n437_), .B(new_new_n108_), .Y(new_new_n438_));
  NO2        g0416(.A(new_new_n438_), .B(new_new_n207_), .Y(new_new_n439_));
  NA2        g0417(.A(new_new_n304_), .B(i_0_), .Y(new_new_n440_));
  NO3        g0418(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n441_));
  NA2        g0419(.A(new_new_n273_), .B(new_new_n101_), .Y(new_new_n442_));
  NA2        g0420(.A(new_new_n442_), .B(new_new_n441_), .Y(new_new_n443_));
  NA2        g0421(.A(i_8_), .B(i_9_), .Y(new_new_n444_));
  AOI210     g0422(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n445_));
  OR2        g0423(.A(new_new_n445_), .B(new_new_n444_), .Y(new_new_n446_));
  NA2        g0424(.A(new_new_n286_), .B(new_new_n208_), .Y(new_new_n447_));
  OAI220     g0425(.A0(new_new_n447_), .A1(new_new_n446_), .B0(new_new_n443_), .B1(new_new_n440_), .Y(new_new_n448_));
  NA2        g0426(.A(new_new_n254_), .B(new_new_n303_), .Y(new_new_n449_));
  NO3        g0427(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n450_));
  INV        g0428(.A(new_new_n450_), .Y(new_new_n451_));
  NA3        g0429(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n452_));
  NA4        g0430(.A(new_new_n150_), .B(new_new_n120_), .C(new_new_n81_), .D(new_new_n23_), .Y(new_new_n453_));
  OAI220     g0431(.A0(new_new_n453_), .A1(new_new_n452_), .B0(new_new_n451_), .B1(new_new_n449_), .Y(new_new_n454_));
  NO3        g0432(.A(new_new_n454_), .B(new_new_n448_), .C(new_new_n439_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n291_), .B(new_new_n112_), .Y(new_new_n456_));
  OR2        g0434(.A(new_new_n456_), .B(new_new_n211_), .Y(new_new_n457_));
  OA210      g0435(.A0(new_new_n346_), .A1(new_new_n105_), .B0(new_new_n293_), .Y(new_new_n458_));
  OA220      g0436(.A0(new_new_n458_), .A1(new_new_n168_), .B0(new_new_n457_), .B1(new_new_n235_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n100_), .B(i_13_), .Y(new_new_n460_));
  NO2        g0438(.A(i_2_), .B(i_13_), .Y(new_new_n461_));
  NA3        g0439(.A(new_new_n461_), .B(new_new_n167_), .C(new_new_n103_), .Y(new_new_n462_));
  NO2        g0440(.A(new_new_n462_), .B(new_new_n240_), .Y(new_new_n463_));
  NO3        g0441(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n464_));
  NO2        g0442(.A(i_6_), .B(i_7_), .Y(new_new_n465_));
  NA2        g0443(.A(new_new_n465_), .B(new_new_n464_), .Y(new_new_n466_));
  NO2        g0444(.A(i_11_), .B(i_1_), .Y(new_new_n467_));
  NO2        g0445(.A(new_new_n74_), .B(i_3_), .Y(new_new_n468_));
  OR2        g0446(.A(i_11_), .B(i_8_), .Y(new_new_n469_));
  NOi21      g0447(.An(i_2_), .B(i_7_), .Y(new_new_n470_));
  NAi31      g0448(.An(new_new_n469_), .B(new_new_n470_), .C(new_new_n468_), .Y(new_new_n471_));
  NO2        g0449(.A(new_new_n409_), .B(i_6_), .Y(new_new_n472_));
  NA3        g0450(.A(new_new_n472_), .B(new_new_n432_), .C(new_new_n76_), .Y(new_new_n473_));
  NO2        g0451(.A(new_new_n473_), .B(new_new_n471_), .Y(new_new_n474_));
  NO2        g0452(.A(i_3_), .B(new_new_n195_), .Y(new_new_n475_));
  NO2        g0453(.A(i_6_), .B(i_10_), .Y(new_new_n476_));
  NA4        g0454(.A(new_new_n476_), .B(new_new_n308_), .C(new_new_n475_), .D(new_new_n240_), .Y(new_new_n477_));
  NO2        g0455(.A(new_new_n477_), .B(new_new_n161_), .Y(new_new_n478_));
  NA3        g0456(.A(new_new_n248_), .B(new_new_n175_), .C(new_new_n137_), .Y(new_new_n479_));
  NA2        g0457(.A(new_new_n47_), .B(new_new_n45_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n163_), .B(i_3_), .Y(new_new_n481_));
  NAi31      g0459(.An(new_new_n480_), .B(new_new_n481_), .C(new_new_n231_), .Y(new_new_n482_));
  NA3        g0460(.A(new_new_n384_), .B(new_new_n183_), .C(new_new_n154_), .Y(new_new_n483_));
  NA3        g0461(.A(new_new_n483_), .B(new_new_n482_), .C(new_new_n479_), .Y(new_new_n484_));
  NO4        g0462(.A(new_new_n484_), .B(new_new_n478_), .C(new_new_n474_), .D(new_new_n463_), .Y(new_new_n485_));
  NA2        g0463(.A(new_new_n441_), .B(new_new_n378_), .Y(new_new_n486_));
  NA2        g0464(.A(new_new_n450_), .B(new_new_n383_), .Y(new_new_n487_));
  NAi21      g0465(.An(new_new_n221_), .B(new_new_n388_), .Y(new_new_n488_));
  NA2        g0466(.A(new_new_n327_), .B(new_new_n223_), .Y(new_new_n489_));
  NO2        g0467(.A(new_new_n26_), .B(i_5_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n489_), .B(new_new_n488_), .Y(new_new_n491_));
  NA2        g0469(.A(new_new_n27_), .B(i_10_), .Y(new_new_n492_));
  NA2        g0470(.A(new_new_n308_), .B(new_new_n242_), .Y(new_new_n493_));
  OAI220     g0471(.A0(new_new_n493_), .A1(new_new_n425_), .B0(new_new_n492_), .B1(new_new_n460_), .Y(new_new_n494_));
  NA4        g0472(.A(new_new_n301_), .B(new_new_n229_), .C(new_new_n74_), .D(new_new_n240_), .Y(new_new_n495_));
  NO2        g0473(.A(new_new_n495_), .B(new_new_n466_), .Y(new_new_n496_));
  NO3        g0474(.A(new_new_n496_), .B(new_new_n494_), .C(new_new_n491_), .Y(new_new_n497_));
  NA4        g0475(.A(new_new_n497_), .B(new_new_n485_), .C(new_new_n459_), .D(new_new_n455_), .Y(new_new_n498_));
  NA3        g0476(.A(new_new_n301_), .B(new_new_n180_), .C(new_new_n178_), .Y(new_new_n499_));
  OAI210     g0477(.A0(new_new_n295_), .A1(new_new_n185_), .B0(new_new_n499_), .Y(new_new_n500_));
  AN2        g0478(.A(new_new_n288_), .B(new_new_n237_), .Y(new_new_n501_));
  NA2        g0479(.A(new_new_n501_), .B(new_new_n500_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n127_), .B(new_new_n116_), .Y(new_new_n503_));
  AN2        g0481(.A(new_new_n503_), .B(new_new_n441_), .Y(new_new_n504_));
  NA2        g0482(.A(new_new_n308_), .B(i_0_), .Y(new_new_n505_));
  OAI210     g0483(.A0(new_new_n505_), .A1(new_new_n235_), .B0(new_new_n302_), .Y(new_new_n506_));
  AOI220     g0484(.A0(new_new_n506_), .A1(new_new_n316_), .B0(new_new_n504_), .B1(new_new_n304_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n378_), .B(new_new_n230_), .Y(new_new_n508_));
  NA2        g0486(.A(new_new_n351_), .B(new_new_n74_), .Y(new_new_n509_));
  NA2        g0487(.A(new_new_n366_), .B(new_new_n361_), .Y(new_new_n510_));
  OR2        g0488(.A(new_new_n508_), .B(new_new_n510_), .Y(new_new_n511_));
  NO2        g0489(.A(new_new_n36_), .B(i_8_), .Y(new_new_n512_));
  AOI210     g0490(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n410_), .Y(new_new_n513_));
  NA2        g0491(.A(new_new_n513_), .B(new_new_n511_), .Y(new_new_n514_));
  INV        g0492(.A(new_new_n514_), .Y(new_new_n515_));
  INV        g0493(.A(new_new_n139_), .Y(new_new_n516_));
  NO2        g0494(.A(i_7_), .B(new_new_n201_), .Y(new_new_n517_));
  OR2        g0495(.A(new_new_n186_), .B(i_4_), .Y(new_new_n518_));
  NO2        g0496(.A(new_new_n518_), .B(new_new_n87_), .Y(new_new_n519_));
  AOI220     g0497(.A0(new_new_n519_), .A1(new_new_n517_), .B0(new_new_n516_), .B1(new_new_n411_), .Y(new_new_n520_));
  NA4        g0498(.A(new_new_n520_), .B(new_new_n515_), .C(new_new_n507_), .D(new_new_n502_), .Y(new_new_n521_));
  NA2        g0499(.A(new_new_n382_), .B(new_new_n291_), .Y(new_new_n522_));
  OAI210     g0500(.A0(new_new_n380_), .A1(new_new_n172_), .B0(new_new_n522_), .Y(new_new_n523_));
  NO2        g0501(.A(i_12_), .B(new_new_n195_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n524_), .B(new_new_n230_), .Y(new_new_n525_));
  NO3        g0503(.A(new_new_n1049_), .B(new_new_n525_), .C(new_new_n456_), .Y(new_new_n526_));
  NOi31      g0504(.An(new_new_n310_), .B(new_new_n409_), .C(new_new_n38_), .Y(new_new_n527_));
  OAI210     g0505(.A0(new_new_n527_), .A1(new_new_n526_), .B0(new_new_n523_), .Y(new_new_n528_));
  NO2        g0506(.A(i_8_), .B(i_7_), .Y(new_new_n529_));
  AOI220     g0507(.A0(new_new_n317_), .A1(new_new_n40_), .B0(new_new_n238_), .B1(new_new_n210_), .Y(new_new_n530_));
  NO2        g0508(.A(new_new_n530_), .B(new_new_n518_), .Y(new_new_n531_));
  NA2        g0509(.A(new_new_n45_), .B(i_10_), .Y(new_new_n532_));
  NO2        g0510(.A(new_new_n532_), .B(i_6_), .Y(new_new_n533_));
  NA3        g0511(.A(new_new_n533_), .B(new_new_n531_), .C(new_new_n529_), .Y(new_new_n534_));
  AOI220     g0512(.A0(new_new_n422_), .A1(new_new_n317_), .B0(new_new_n250_), .B1(new_new_n247_), .Y(new_new_n535_));
  OAI220     g0513(.A0(new_new_n535_), .A1(new_new_n269_), .B0(new_new_n460_), .B1(new_new_n138_), .Y(new_new_n536_));
  NA2        g0514(.A(new_new_n536_), .B(new_new_n272_), .Y(new_new_n537_));
  NOi31      g0515(.An(new_new_n289_), .B(new_new_n295_), .C(new_new_n185_), .Y(new_new_n538_));
  NA3        g0516(.A(new_new_n301_), .B(new_new_n178_), .C(new_new_n100_), .Y(new_new_n539_));
  NO2        g0517(.A(new_new_n227_), .B(new_new_n45_), .Y(new_new_n540_));
  NO2        g0518(.A(new_new_n163_), .B(i_5_), .Y(new_new_n541_));
  NA3        g0519(.A(new_new_n541_), .B(new_new_n397_), .C(new_new_n311_), .Y(new_new_n542_));
  OAI210     g0520(.A0(new_new_n542_), .A1(new_new_n540_), .B0(new_new_n539_), .Y(new_new_n543_));
  OAI210     g0521(.A0(new_new_n543_), .A1(new_new_n538_), .B0(new_new_n450_), .Y(new_new_n544_));
  NA4        g0522(.A(new_new_n544_), .B(new_new_n537_), .C(new_new_n534_), .D(new_new_n528_), .Y(new_new_n545_));
  NA3        g0523(.A(new_new_n223_), .B(new_new_n72_), .C(new_new_n45_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n286_), .B(new_new_n85_), .Y(new_new_n547_));
  AOI210     g0525(.A0(new_new_n546_), .A1(new_new_n341_), .B0(new_new_n547_), .Y(new_new_n548_));
  NA2        g0526(.A(new_new_n292_), .B(new_new_n288_), .Y(new_new_n549_));
  NO2        g0527(.A(new_new_n549_), .B(new_new_n177_), .Y(new_new_n550_));
  NA2        g0528(.A(new_new_n229_), .B(new_new_n228_), .Y(new_new_n551_));
  NA2        g0529(.A(new_new_n434_), .B(new_new_n227_), .Y(new_new_n552_));
  NO2        g0530(.A(new_new_n551_), .B(new_new_n552_), .Y(new_new_n553_));
  AOI210     g0531(.A0(i_6_), .A1(new_new_n47_), .B0(new_new_n363_), .Y(new_new_n554_));
  NA2        g0532(.A(i_0_), .B(new_new_n49_), .Y(new_new_n555_));
  NA3        g0533(.A(new_new_n524_), .B(new_new_n281_), .C(new_new_n555_), .Y(new_new_n556_));
  NO2        g0534(.A(new_new_n554_), .B(new_new_n556_), .Y(new_new_n557_));
  NO4        g0535(.A(new_new_n557_), .B(new_new_n553_), .C(new_new_n550_), .D(new_new_n548_), .Y(new_new_n558_));
  NO4        g0536(.A(new_new_n255_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n559_));
  NO3        g0537(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n560_));
  NO2        g0538(.A(new_new_n236_), .B(new_new_n36_), .Y(new_new_n561_));
  AN2        g0539(.A(new_new_n561_), .B(new_new_n560_), .Y(new_new_n562_));
  OA210      g0540(.A0(new_new_n562_), .A1(new_new_n559_), .B0(new_new_n351_), .Y(new_new_n563_));
  NO2        g0541(.A(new_new_n409_), .B(i_1_), .Y(new_new_n564_));
  NOi31      g0542(.An(new_new_n564_), .B(new_new_n442_), .C(new_new_n74_), .Y(new_new_n565_));
  AN4        g0543(.A(new_new_n565_), .B(new_new_n406_), .C(new_new_n490_), .D(i_2_), .Y(new_new_n566_));
  NO2        g0544(.A(new_new_n420_), .B(new_new_n181_), .Y(new_new_n567_));
  NO3        g0545(.A(new_new_n567_), .B(new_new_n566_), .C(new_new_n563_), .Y(new_new_n568_));
  NOi21      g0546(.An(i_10_), .B(i_6_), .Y(new_new_n569_));
  NO2        g0547(.A(new_new_n87_), .B(new_new_n25_), .Y(new_new_n570_));
  AOI220     g0548(.A0(new_new_n286_), .A1(new_new_n570_), .B0(new_new_n281_), .B1(new_new_n569_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n571_), .B(new_new_n440_), .Y(new_new_n572_));
  NO2        g0550(.A(new_new_n119_), .B(new_new_n23_), .Y(new_new_n573_));
  NO2        g0551(.A(new_new_n200_), .B(new_new_n37_), .Y(new_new_n574_));
  NOi31      g0552(.An(new_new_n151_), .B(new_new_n574_), .C(new_new_n323_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n575_), .B(new_new_n572_), .Y(new_new_n576_));
  NO2        g0554(.A(new_new_n509_), .B(new_new_n374_), .Y(new_new_n577_));
  INV        g0555(.A(new_new_n311_), .Y(new_new_n578_));
  NO2        g0556(.A(i_12_), .B(new_new_n87_), .Y(new_new_n579_));
  NA2        g0557(.A(new_new_n178_), .B(i_0_), .Y(new_new_n580_));
  NO3        g0558(.A(new_new_n580_), .B(new_new_n333_), .C(new_new_n295_), .Y(new_new_n581_));
  OR2        g0559(.A(i_2_), .B(i_5_), .Y(new_new_n582_));
  OR2        g0560(.A(new_new_n582_), .B(new_new_n401_), .Y(new_new_n583_));
  NO2        g0561(.A(new_new_n583_), .B(new_new_n488_), .Y(new_new_n584_));
  NO3        g0562(.A(new_new_n584_), .B(new_new_n581_), .C(new_new_n577_), .Y(new_new_n585_));
  NA4        g0563(.A(new_new_n585_), .B(new_new_n576_), .C(new_new_n568_), .D(new_new_n558_), .Y(new_new_n586_));
  NO4        g0564(.A(new_new_n586_), .B(new_new_n545_), .C(new_new_n521_), .D(new_new_n498_), .Y(new_new_n587_));
  NA4        g0565(.A(new_new_n587_), .B(new_new_n431_), .C(new_new_n350_), .D(new_new_n307_), .Y(mai7));
  NO2        g0566(.A(new_new_n96_), .B(new_new_n55_), .Y(new_new_n589_));
  NO2        g0567(.A(new_new_n112_), .B(new_new_n93_), .Y(new_new_n590_));
  NA2        g0568(.A(new_new_n476_), .B(new_new_n85_), .Y(new_new_n591_));
  NA2        g0569(.A(i_11_), .B(new_new_n195_), .Y(new_new_n592_));
  NA3        g0570(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n240_), .B(i_4_), .Y(new_new_n594_));
  NA2        g0572(.A(new_new_n594_), .B(i_8_), .Y(new_new_n595_));
  NO2        g0573(.A(new_new_n109_), .B(new_new_n593_), .Y(new_new_n596_));
  NA2        g0574(.A(i_2_), .B(new_new_n87_), .Y(new_new_n597_));
  OAI210     g0575(.A0(new_new_n90_), .A1(new_new_n205_), .B0(new_new_n206_), .Y(new_new_n598_));
  NO2        g0576(.A(i_7_), .B(new_new_n37_), .Y(new_new_n599_));
  NA2        g0577(.A(i_4_), .B(i_8_), .Y(new_new_n600_));
  AOI210     g0578(.A0(new_new_n600_), .A1(new_new_n301_), .B0(new_new_n599_), .Y(new_new_n601_));
  OAI220     g0579(.A0(new_new_n601_), .A1(new_new_n597_), .B0(new_new_n598_), .B1(i_13_), .Y(new_new_n602_));
  NO3        g0580(.A(new_new_n602_), .B(new_new_n596_), .C(new_new_n589_), .Y(new_new_n603_));
  AOI210     g0581(.A0(new_new_n133_), .A1(new_new_n63_), .B0(i_10_), .Y(new_new_n604_));
  AOI210     g0582(.A0(new_new_n604_), .A1(new_new_n240_), .B0(new_new_n167_), .Y(new_new_n605_));
  OR2        g0583(.A(i_6_), .B(i_10_), .Y(new_new_n606_));
  NO2        g0584(.A(new_new_n606_), .B(new_new_n23_), .Y(new_new_n607_));
  OR3        g0585(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n608_));
  NO3        g0586(.A(new_new_n608_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n609_));
  INV        g0587(.A(new_new_n202_), .Y(new_new_n610_));
  NO2        g0588(.A(new_new_n609_), .B(new_new_n607_), .Y(new_new_n611_));
  OA220      g0589(.A0(new_new_n611_), .A1(new_new_n578_), .B0(new_new_n605_), .B1(new_new_n274_), .Y(new_new_n612_));
  AOI210     g0590(.A0(new_new_n612_), .A1(new_new_n603_), .B0(new_new_n64_), .Y(new_new_n613_));
  NOi21      g0591(.An(i_11_), .B(i_7_), .Y(new_new_n614_));
  AO210      g0592(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n615_));
  NO2        g0593(.A(new_new_n615_), .B(new_new_n614_), .Y(new_new_n616_));
  NA2        g0594(.A(new_new_n616_), .B(new_new_n210_), .Y(new_new_n617_));
  NO2        g0595(.A(new_new_n617_), .B(new_new_n64_), .Y(new_new_n618_));
  NA2        g0596(.A(new_new_n89_), .B(new_new_n64_), .Y(new_new_n619_));
  AO210      g0597(.A0(new_new_n619_), .A1(new_new_n374_), .B0(new_new_n41_), .Y(new_new_n620_));
  NO3        g0598(.A(new_new_n263_), .B(new_new_n212_), .C(new_new_n592_), .Y(new_new_n621_));
  OAI210     g0599(.A0(new_new_n621_), .A1(new_new_n231_), .B0(new_new_n64_), .Y(new_new_n622_));
  NA2        g0600(.A(new_new_n402_), .B(new_new_n31_), .Y(new_new_n623_));
  OR2        g0601(.A(new_new_n212_), .B(new_new_n112_), .Y(new_new_n624_));
  NA2        g0602(.A(new_new_n624_), .B(new_new_n623_), .Y(new_new_n625_));
  NO2        g0603(.A(new_new_n64_), .B(i_9_), .Y(new_new_n626_));
  NO2        g0604(.A(new_new_n626_), .B(i_4_), .Y(new_new_n627_));
  NA2        g0605(.A(new_new_n627_), .B(new_new_n625_), .Y(new_new_n628_));
  NO2        g0606(.A(i_1_), .B(i_12_), .Y(new_new_n629_));
  NA3        g0607(.A(new_new_n629_), .B(new_new_n114_), .C(new_new_n24_), .Y(new_new_n630_));
  BUFFER     g0608(.A(new_new_n630_), .Y(new_new_n631_));
  NA4        g0609(.A(new_new_n631_), .B(new_new_n628_), .C(new_new_n622_), .D(new_new_n620_), .Y(new_new_n632_));
  OAI210     g0610(.A0(new_new_n632_), .A1(new_new_n618_), .B0(i_6_), .Y(new_new_n633_));
  NO2        g0611(.A(i_6_), .B(i_11_), .Y(new_new_n634_));
  INV        g0612(.A(new_new_n443_), .Y(new_new_n635_));
  NO4        g0613(.A(new_new_n220_), .B(new_new_n133_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n636_));
  NA2        g0614(.A(new_new_n636_), .B(new_new_n626_), .Y(new_new_n637_));
  NA2        g0615(.A(new_new_n240_), .B(i_6_), .Y(new_new_n638_));
  NO3        g0616(.A(new_new_n606_), .B(new_new_n236_), .C(new_new_n23_), .Y(new_new_n639_));
  AOI210     g0617(.A0(i_1_), .A1(new_new_n264_), .B0(new_new_n639_), .Y(new_new_n640_));
  OAI210     g0618(.A0(new_new_n640_), .A1(new_new_n45_), .B0(new_new_n637_), .Y(new_new_n641_));
  INV        g0619(.A(i_2_), .Y(new_new_n642_));
  NA2        g0620(.A(new_new_n143_), .B(i_9_), .Y(new_new_n643_));
  NA3        g0621(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n644_));
  NO2        g0622(.A(new_new_n47_), .B(i_1_), .Y(new_new_n645_));
  NA3        g0623(.A(new_new_n645_), .B(new_new_n273_), .C(new_new_n45_), .Y(new_new_n646_));
  OAI220     g0624(.A0(new_new_n646_), .A1(new_new_n644_), .B0(new_new_n643_), .B1(new_new_n642_), .Y(new_new_n647_));
  NA3        g0625(.A(new_new_n626_), .B(new_new_n311_), .C(i_6_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n648_), .B(new_new_n23_), .Y(new_new_n649_));
  AOI210     g0627(.A0(new_new_n467_), .A1(new_new_n413_), .B0(new_new_n245_), .Y(new_new_n650_));
  NO2        g0628(.A(new_new_n650_), .B(new_new_n597_), .Y(new_new_n651_));
  NO2        g0629(.A(i_11_), .B(new_new_n37_), .Y(new_new_n652_));
  OR3        g0630(.A(new_new_n651_), .B(new_new_n649_), .C(new_new_n647_), .Y(new_new_n653_));
  NO3        g0631(.A(new_new_n653_), .B(new_new_n641_), .C(new_new_n635_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n240_), .B(new_new_n105_), .Y(new_new_n655_));
  NO2        g0633(.A(new_new_n655_), .B(new_new_n614_), .Y(new_new_n656_));
  NA2        g0634(.A(new_new_n656_), .B(i_1_), .Y(new_new_n657_));
  NO2        g0635(.A(new_new_n657_), .B(new_new_n608_), .Y(new_new_n658_));
  NO2        g0636(.A(new_new_n408_), .B(new_new_n87_), .Y(new_new_n659_));
  NA2        g0637(.A(new_new_n658_), .B(new_new_n47_), .Y(new_new_n660_));
  NA2        g0638(.A(i_3_), .B(new_new_n195_), .Y(new_new_n661_));
  NO2        g0639(.A(new_new_n661_), .B(new_new_n119_), .Y(new_new_n662_));
  AN2        g0640(.A(new_new_n662_), .B(new_new_n533_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n236_), .B(new_new_n45_), .Y(new_new_n664_));
  NO3        g0642(.A(new_new_n664_), .B(new_new_n304_), .C(new_new_n241_), .Y(new_new_n665_));
  NO2        g0643(.A(new_new_n122_), .B(new_new_n37_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n666_), .B(i_6_), .Y(new_new_n667_));
  NO2        g0645(.A(new_new_n87_), .B(i_9_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n64_), .Y(new_new_n669_));
  NO2        g0647(.A(new_new_n669_), .B(new_new_n629_), .Y(new_new_n670_));
  NO4        g0648(.A(new_new_n670_), .B(new_new_n667_), .C(new_new_n665_), .D(i_4_), .Y(new_new_n671_));
  NA2        g0649(.A(i_1_), .B(i_3_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n444_), .B(new_new_n96_), .Y(new_new_n673_));
  AOI210     g0651(.A0(new_new_n664_), .A1(new_new_n569_), .B0(new_new_n673_), .Y(new_new_n674_));
  NO2        g0652(.A(new_new_n674_), .B(new_new_n672_), .Y(new_new_n675_));
  NO3        g0653(.A(new_new_n675_), .B(new_new_n671_), .C(new_new_n663_), .Y(new_new_n676_));
  NA4        g0654(.A(new_new_n676_), .B(new_new_n660_), .C(new_new_n654_), .D(new_new_n633_), .Y(new_new_n677_));
  NO3        g0655(.A(new_new_n469_), .B(i_3_), .C(i_7_), .Y(new_new_n678_));
  NOi21      g0656(.An(new_new_n678_), .B(i_10_), .Y(new_new_n679_));
  OA210      g0657(.A0(new_new_n679_), .A1(new_new_n248_), .B0(new_new_n87_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n366_), .B(new_new_n365_), .Y(new_new_n681_));
  NA3        g0659(.A(new_new_n476_), .B(new_new_n512_), .C(new_new_n47_), .Y(new_new_n682_));
  NA3        g0660(.A(new_new_n167_), .B(new_new_n85_), .C(new_new_n87_), .Y(new_new_n683_));
  NA3        g0661(.A(new_new_n683_), .B(new_new_n682_), .C(new_new_n681_), .Y(new_new_n684_));
  OAI210     g0662(.A0(new_new_n684_), .A1(new_new_n680_), .B0(i_1_), .Y(new_new_n685_));
  AOI210     g0663(.A0(new_new_n273_), .A1(new_new_n101_), .B0(i_1_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n364_), .B(i_2_), .Y(new_new_n687_));
  NA2        g0665(.A(new_new_n687_), .B(new_new_n686_), .Y(new_new_n688_));
  OAI210     g0666(.A0(new_new_n648_), .A1(new_new_n435_), .B0(new_new_n688_), .Y(new_new_n689_));
  INV        g0667(.A(new_new_n689_), .Y(new_new_n690_));
  AOI210     g0668(.A0(new_new_n690_), .A1(new_new_n685_), .B0(i_13_), .Y(new_new_n691_));
  OR2        g0669(.A(i_11_), .B(i_7_), .Y(new_new_n692_));
  AOI210     g0670(.A0(new_new_n644_), .A1(new_new_n55_), .B0(i_12_), .Y(new_new_n693_));
  NO2        g0671(.A(new_new_n470_), .B(new_new_n24_), .Y(new_new_n694_));
  AOI220     g0672(.A0(new_new_n694_), .A1(new_new_n659_), .B0(new_new_n248_), .B1(new_new_n136_), .Y(new_new_n695_));
  OAI220     g0673(.A0(new_new_n695_), .A1(new_new_n41_), .B0(new_new_n1048_), .B1(new_new_n96_), .Y(new_new_n696_));
  INV        g0674(.A(new_new_n696_), .Y(new_new_n697_));
  INV        g0675(.A(new_new_n119_), .Y(new_new_n698_));
  AOI220     g0676(.A0(new_new_n698_), .A1(new_new_n73_), .B0(new_new_n381_), .B1(new_new_n645_), .Y(new_new_n699_));
  NO2        g0677(.A(new_new_n699_), .B(new_new_n246_), .Y(new_new_n700_));
  AOI210     g0678(.A0(new_new_n435_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n701_));
  NOi31      g0679(.An(new_new_n701_), .B(new_new_n591_), .C(new_new_n45_), .Y(new_new_n702_));
  NA2        g0680(.A(new_new_n132_), .B(i_13_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n644_), .B(new_new_n119_), .Y(new_new_n704_));
  INV        g0682(.A(new_new_n704_), .Y(new_new_n705_));
  OAI220     g0683(.A0(new_new_n705_), .A1(new_new_n72_), .B0(new_new_n703_), .B1(new_new_n686_), .Y(new_new_n706_));
  NO3        g0684(.A(new_new_n72_), .B(new_new_n32_), .C(new_new_n105_), .Y(new_new_n707_));
  NA2        g0685(.A(new_new_n26_), .B(new_new_n195_), .Y(new_new_n708_));
  NA2        g0686(.A(new_new_n708_), .B(i_7_), .Y(new_new_n709_));
  NO3        g0687(.A(new_new_n470_), .B(new_new_n240_), .C(new_new_n87_), .Y(new_new_n710_));
  AOI210     g0688(.A0(new_new_n710_), .A1(new_new_n709_), .B0(new_new_n707_), .Y(new_new_n711_));
  AOI220     g0689(.A0(new_new_n381_), .A1(new_new_n645_), .B0(new_new_n95_), .B1(new_new_n106_), .Y(new_new_n712_));
  OAI220     g0690(.A0(new_new_n712_), .A1(new_new_n595_), .B0(new_new_n711_), .B1(new_new_n610_), .Y(new_new_n713_));
  NO4        g0691(.A(new_new_n713_), .B(new_new_n706_), .C(new_new_n702_), .D(new_new_n700_), .Y(new_new_n714_));
  OR2        g0692(.A(i_11_), .B(i_6_), .Y(new_new_n715_));
  NA3        g0693(.A(new_new_n594_), .B(new_new_n708_), .C(i_7_), .Y(new_new_n716_));
  AOI210     g0694(.A0(new_new_n716_), .A1(new_new_n705_), .B0(new_new_n715_), .Y(new_new_n717_));
  NA3        g0695(.A(new_new_n402_), .B(new_new_n599_), .C(new_new_n101_), .Y(new_new_n718_));
  NA2        g0696(.A(new_new_n634_), .B(i_13_), .Y(new_new_n719_));
  NA2        g0697(.A(new_new_n106_), .B(new_new_n708_), .Y(new_new_n720_));
  NAi21      g0698(.An(i_11_), .B(i_12_), .Y(new_new_n721_));
  NOi41      g0699(.An(new_new_n115_), .B(new_new_n721_), .C(i_13_), .D(new_new_n87_), .Y(new_new_n722_));
  NA2        g0700(.A(new_new_n722_), .B(new_new_n720_), .Y(new_new_n723_));
  NA3        g0701(.A(new_new_n723_), .B(new_new_n719_), .C(new_new_n718_), .Y(new_new_n724_));
  OAI210     g0702(.A0(new_new_n724_), .A1(new_new_n717_), .B0(new_new_n64_), .Y(new_new_n725_));
  NO2        g0703(.A(i_2_), .B(i_12_), .Y(new_new_n726_));
  NA2        g0704(.A(new_new_n363_), .B(new_new_n726_), .Y(new_new_n727_));
  NA2        g0705(.A(i_8_), .B(new_new_n25_), .Y(new_new_n728_));
  NO3        g0706(.A(new_new_n728_), .B(new_new_n379_), .C(new_new_n594_), .Y(new_new_n729_));
  OAI210     g0707(.A0(new_new_n729_), .A1(new_new_n365_), .B0(new_new_n363_), .Y(new_new_n730_));
  NO2        g0708(.A(new_new_n133_), .B(i_2_), .Y(new_new_n731_));
  NA2        g0709(.A(new_new_n731_), .B(new_new_n629_), .Y(new_new_n732_));
  NA3        g0710(.A(new_new_n732_), .B(new_new_n730_), .C(new_new_n727_), .Y(new_new_n733_));
  NA3        g0711(.A(new_new_n733_), .B(new_new_n46_), .C(new_new_n230_), .Y(new_new_n734_));
  NA4        g0712(.A(new_new_n734_), .B(new_new_n725_), .C(new_new_n714_), .D(new_new_n697_), .Y(new_new_n735_));
  OR4        g0713(.A(new_new_n735_), .B(new_new_n691_), .C(new_new_n677_), .D(new_new_n613_), .Y(mai5));
  NA2        g0714(.A(new_new_n656_), .B(new_new_n276_), .Y(new_new_n737_));
  AN2        g0715(.A(new_new_n24_), .B(i_10_), .Y(new_new_n738_));
  NA3        g0716(.A(new_new_n738_), .B(new_new_n726_), .C(new_new_n112_), .Y(new_new_n739_));
  NO2        g0717(.A(new_new_n595_), .B(i_11_), .Y(new_new_n740_));
  NA2        g0718(.A(new_new_n90_), .B(new_new_n740_), .Y(new_new_n741_));
  NA3        g0719(.A(new_new_n741_), .B(new_new_n739_), .C(new_new_n737_), .Y(new_new_n742_));
  NO3        g0720(.A(i_11_), .B(new_new_n240_), .C(i_13_), .Y(new_new_n743_));
  NO2        g0721(.A(new_new_n129_), .B(new_new_n23_), .Y(new_new_n744_));
  NA2        g0722(.A(i_12_), .B(i_8_), .Y(new_new_n745_));
  OAI210     g0723(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n745_), .Y(new_new_n746_));
  INV        g0724(.A(new_new_n434_), .Y(new_new_n747_));
  AOI220     g0725(.A0(new_new_n311_), .A1(new_new_n573_), .B0(new_new_n746_), .B1(new_new_n744_), .Y(new_new_n748_));
  INV        g0726(.A(new_new_n748_), .Y(new_new_n749_));
  NO2        g0727(.A(new_new_n749_), .B(new_new_n742_), .Y(new_new_n750_));
  INV        g0728(.A(new_new_n175_), .Y(new_new_n751_));
  INV        g0729(.A(new_new_n248_), .Y(new_new_n752_));
  OAI210     g0730(.A0(new_new_n687_), .A1(new_new_n436_), .B0(new_new_n115_), .Y(new_new_n753_));
  AOI210     g0731(.A0(new_new_n753_), .A1(new_new_n752_), .B0(new_new_n751_), .Y(new_new_n754_));
  NO2        g0732(.A(new_new_n444_), .B(new_new_n26_), .Y(new_new_n755_));
  NO2        g0733(.A(new_new_n755_), .B(new_new_n413_), .Y(new_new_n756_));
  NA2        g0734(.A(new_new_n756_), .B(i_2_), .Y(new_new_n757_));
  INV        g0735(.A(new_new_n757_), .Y(new_new_n758_));
  AOI210     g0736(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n409_), .Y(new_new_n759_));
  AOI210     g0737(.A0(new_new_n759_), .A1(new_new_n758_), .B0(new_new_n754_), .Y(new_new_n760_));
  NO2        g0738(.A(new_new_n192_), .B(new_new_n130_), .Y(new_new_n761_));
  OAI210     g0739(.A0(new_new_n761_), .A1(new_new_n744_), .B0(i_2_), .Y(new_new_n762_));
  INV        g0740(.A(new_new_n176_), .Y(new_new_n763_));
  NO3        g0741(.A(new_new_n615_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n764_));
  AOI210     g0742(.A0(new_new_n763_), .A1(new_new_n90_), .B0(new_new_n764_), .Y(new_new_n765_));
  AOI210     g0743(.A0(new_new_n765_), .A1(new_new_n762_), .B0(new_new_n195_), .Y(new_new_n766_));
  OA210      g0744(.A0(new_new_n616_), .A1(new_new_n131_), .B0(i_13_), .Y(new_new_n767_));
  NA2        g0745(.A(new_new_n202_), .B(new_new_n205_), .Y(new_new_n768_));
  NA2        g0746(.A(new_new_n157_), .B(new_new_n592_), .Y(new_new_n769_));
  AOI210     g0747(.A0(new_new_n769_), .A1(new_new_n768_), .B0(new_new_n368_), .Y(new_new_n770_));
  AOI210     g0748(.A0(new_new_n212_), .A1(new_new_n153_), .B0(new_new_n512_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(new_new_n413_), .Y(new_new_n772_));
  NO2        g0750(.A(new_new_n106_), .B(new_new_n45_), .Y(new_new_n773_));
  INV        g0751(.A(new_new_n296_), .Y(new_new_n774_));
  NA4        g0752(.A(new_new_n774_), .B(new_new_n301_), .C(new_new_n129_), .D(new_new_n43_), .Y(new_new_n775_));
  OAI210     g0753(.A0(new_new_n775_), .A1(new_new_n773_), .B0(new_new_n772_), .Y(new_new_n776_));
  NO4        g0754(.A(new_new_n776_), .B(new_new_n770_), .C(new_new_n767_), .D(new_new_n766_), .Y(new_new_n777_));
  NA2        g0755(.A(new_new_n573_), .B(new_new_n28_), .Y(new_new_n778_));
  NA2        g0756(.A(new_new_n743_), .B(new_new_n282_), .Y(new_new_n779_));
  NA2        g0757(.A(new_new_n779_), .B(new_new_n778_), .Y(new_new_n780_));
  NO2        g0758(.A(new_new_n63_), .B(i_12_), .Y(new_new_n781_));
  NO2        g0759(.A(new_new_n781_), .B(new_new_n131_), .Y(new_new_n782_));
  NO2        g0760(.A(new_new_n782_), .B(new_new_n592_), .Y(new_new_n783_));
  AOI220     g0761(.A0(new_new_n783_), .A1(new_new_n36_), .B0(new_new_n780_), .B1(new_new_n47_), .Y(new_new_n784_));
  NA4        g0762(.A(new_new_n784_), .B(new_new_n777_), .C(new_new_n760_), .D(new_new_n750_), .Y(mai6));
  NO2        g0763(.A(new_new_n187_), .B(new_new_n144_), .Y(new_new_n786_));
  NA2        g0764(.A(new_new_n786_), .B(new_new_n731_), .Y(new_new_n787_));
  NA4        g0765(.A(new_new_n383_), .B(new_new_n475_), .C(new_new_n72_), .D(new_new_n105_), .Y(new_new_n788_));
  INV        g0766(.A(new_new_n788_), .Y(new_new_n789_));
  NO2        g0767(.A(new_new_n226_), .B(new_new_n480_), .Y(new_new_n790_));
  NO2        g0768(.A(i_11_), .B(i_9_), .Y(new_new_n791_));
  NO2        g0769(.A(new_new_n789_), .B(new_new_n322_), .Y(new_new_n792_));
  AO210      g0770(.A0(new_new_n792_), .A1(new_new_n787_), .B0(i_12_), .Y(new_new_n793_));
  NA2        g0771(.A(new_new_n369_), .B(new_new_n327_), .Y(new_new_n794_));
  NA2        g0772(.A(new_new_n579_), .B(new_new_n64_), .Y(new_new_n795_));
  NA2        g0773(.A(new_new_n679_), .B(new_new_n72_), .Y(new_new_n796_));
  BUFFER     g0774(.A(new_new_n619_), .Y(new_new_n797_));
  NA4        g0775(.A(new_new_n797_), .B(new_new_n796_), .C(new_new_n795_), .D(new_new_n794_), .Y(new_new_n798_));
  INV        g0776(.A(new_new_n199_), .Y(new_new_n799_));
  AOI220     g0777(.A0(new_new_n799_), .A1(new_new_n791_), .B0(new_new_n798_), .B1(new_new_n74_), .Y(new_new_n800_));
  INV        g0778(.A(new_new_n321_), .Y(new_new_n801_));
  NA2        g0779(.A(new_new_n76_), .B(new_new_n136_), .Y(new_new_n802_));
  INV        g0780(.A(new_new_n129_), .Y(new_new_n803_));
  NA2        g0781(.A(new_new_n803_), .B(new_new_n47_), .Y(new_new_n804_));
  AOI210     g0782(.A0(new_new_n804_), .A1(new_new_n802_), .B0(new_new_n801_), .Y(new_new_n805_));
  NO3        g0783(.A(new_new_n255_), .B(new_new_n137_), .C(i_9_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n806_), .B(new_new_n781_), .Y(new_new_n807_));
  AOI210     g0785(.A0(new_new_n807_), .A1(new_new_n510_), .B0(new_new_n187_), .Y(new_new_n808_));
  NO2        g0786(.A(new_new_n32_), .B(i_11_), .Y(new_new_n809_));
  NA3        g0787(.A(new_new_n809_), .B(new_new_n465_), .C(new_new_n383_), .Y(new_new_n810_));
  NAi32      g0788(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n811_));
  NO2        g0789(.A(new_new_n715_), .B(new_new_n811_), .Y(new_new_n812_));
  OAI210     g0790(.A0(new_new_n678_), .A1(new_new_n561_), .B0(new_new_n560_), .Y(new_new_n813_));
  NAi31      g0791(.An(new_new_n812_), .B(new_new_n813_), .C(new_new_n810_), .Y(new_new_n814_));
  OR3        g0792(.A(new_new_n814_), .B(new_new_n808_), .C(new_new_n805_), .Y(new_new_n815_));
  NO2        g0793(.A(new_new_n692_), .B(i_2_), .Y(new_new_n816_));
  NA2        g0794(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n817_), .B(new_new_n401_), .Y(new_new_n818_));
  NA2        g0796(.A(new_new_n818_), .B(new_new_n816_), .Y(new_new_n819_));
  AO220      g0797(.A0(new_new_n355_), .A1(new_new_n345_), .B0(new_new_n385_), .B1(new_new_n592_), .Y(new_new_n820_));
  NA3        g0798(.A(new_new_n820_), .B(new_new_n260_), .C(i_7_), .Y(new_new_n821_));
  NA3        g0799(.A(new_new_n616_), .B(new_new_n152_), .C(new_new_n70_), .Y(new_new_n822_));
  AO210      g0800(.A0(new_new_n487_), .A1(new_new_n747_), .B0(new_new_n36_), .Y(new_new_n823_));
  NA4        g0801(.A(new_new_n823_), .B(new_new_n822_), .C(new_new_n821_), .D(new_new_n819_), .Y(new_new_n824_));
  OAI210     g0802(.A0(i_6_), .A1(i_11_), .B0(new_new_n88_), .Y(new_new_n825_));
  AOI220     g0803(.A0(new_new_n825_), .A1(new_new_n560_), .B0(new_new_n790_), .B1(new_new_n709_), .Y(new_new_n826_));
  NA3        g0804(.A(new_new_n368_), .B(new_new_n242_), .C(new_new_n152_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n385_), .B(new_new_n71_), .Y(new_new_n828_));
  NA4        g0806(.A(new_new_n828_), .B(new_new_n827_), .C(new_new_n826_), .D(new_new_n598_), .Y(new_new_n829_));
  AO210      g0807(.A0(new_new_n512_), .A1(new_new_n47_), .B0(new_new_n89_), .Y(new_new_n830_));
  NA3        g0808(.A(new_new_n830_), .B(new_new_n476_), .C(new_new_n223_), .Y(new_new_n831_));
  AOI210     g0809(.A0(new_new_n436_), .A1(new_new_n434_), .B0(new_new_n559_), .Y(new_new_n832_));
  NO2        g0810(.A(new_new_n606_), .B(new_new_n106_), .Y(new_new_n833_));
  OAI210     g0811(.A0(new_new_n833_), .A1(new_new_n116_), .B0(new_new_n399_), .Y(new_new_n834_));
  INV        g0812(.A(new_new_n583_), .Y(new_new_n835_));
  NA3        g0813(.A(new_new_n835_), .B(new_new_n321_), .C(i_7_), .Y(new_new_n836_));
  NA4        g0814(.A(new_new_n836_), .B(new_new_n834_), .C(new_new_n832_), .D(new_new_n831_), .Y(new_new_n837_));
  NO4        g0815(.A(new_new_n837_), .B(new_new_n829_), .C(new_new_n824_), .D(new_new_n815_), .Y(new_new_n838_));
  NA4        g0816(.A(new_new_n838_), .B(new_new_n800_), .C(new_new_n793_), .D(new_new_n376_), .Y(mai3));
  NA2        g0817(.A(i_6_), .B(i_7_), .Y(new_new_n840_));
  NO2        g0818(.A(new_new_n840_), .B(i_0_), .Y(new_new_n841_));
  NO2        g0819(.A(i_11_), .B(new_new_n240_), .Y(new_new_n842_));
  OAI210     g0820(.A0(new_new_n841_), .A1(new_new_n289_), .B0(new_new_n842_), .Y(new_new_n843_));
  NO2        g0821(.A(new_new_n843_), .B(new_new_n195_), .Y(new_new_n844_));
  NO3        g0822(.A(new_new_n440_), .B(new_new_n93_), .C(new_new_n45_), .Y(new_new_n845_));
  OA210      g0823(.A0(new_new_n845_), .A1(new_new_n844_), .B0(new_new_n178_), .Y(new_new_n846_));
  NA3        g0824(.A(new_new_n827_), .B(new_new_n598_), .C(new_new_n367_), .Y(new_new_n847_));
  NA2        g0825(.A(new_new_n847_), .B(new_new_n40_), .Y(new_new_n848_));
  NOi21      g0826(.An(new_new_n100_), .B(new_new_n756_), .Y(new_new_n849_));
  NO3        g0827(.A(new_new_n624_), .B(new_new_n444_), .C(new_new_n136_), .Y(new_new_n850_));
  NA2        g0828(.A(new_new_n402_), .B(new_new_n46_), .Y(new_new_n851_));
  AN2        g0829(.A(new_new_n442_), .B(new_new_n56_), .Y(new_new_n852_));
  NO3        g0830(.A(new_new_n852_), .B(new_new_n850_), .C(new_new_n849_), .Y(new_new_n853_));
  AOI210     g0831(.A0(new_new_n853_), .A1(new_new_n848_), .B0(new_new_n49_), .Y(new_new_n854_));
  NO4        g0832(.A(new_new_n372_), .B(new_new_n378_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n855_));
  NA2        g0833(.A(new_new_n187_), .B(new_new_n569_), .Y(new_new_n856_));
  NOi21      g0834(.An(new_new_n856_), .B(new_new_n855_), .Y(new_new_n857_));
  NO2        g0835(.A(new_new_n857_), .B(new_new_n64_), .Y(new_new_n858_));
  NOi21      g0836(.An(i_5_), .B(i_9_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n859_), .B(new_new_n433_), .Y(new_new_n860_));
  BUFFER     g0838(.A(new_new_n273_), .Y(new_new_n861_));
  NA2        g0839(.A(new_new_n861_), .B(new_new_n467_), .Y(new_new_n862_));
  NO3        g0840(.A(new_new_n405_), .B(new_new_n273_), .C(new_new_n74_), .Y(new_new_n863_));
  NO2        g0841(.A(new_new_n179_), .B(new_new_n153_), .Y(new_new_n864_));
  AOI210     g0842(.A0(new_new_n864_), .A1(new_new_n247_), .B0(new_new_n863_), .Y(new_new_n865_));
  OAI220     g0843(.A0(new_new_n865_), .A1(new_new_n185_), .B0(new_new_n862_), .B1(new_new_n860_), .Y(new_new_n866_));
  NO4        g0844(.A(new_new_n866_), .B(new_new_n858_), .C(new_new_n854_), .D(new_new_n846_), .Y(new_new_n867_));
  NA2        g0845(.A(new_new_n187_), .B(new_new_n24_), .Y(new_new_n868_));
  NO2        g0846(.A(new_new_n666_), .B(new_new_n590_), .Y(new_new_n869_));
  NO2        g0847(.A(new_new_n869_), .B(new_new_n868_), .Y(new_new_n870_));
  INV        g0848(.A(new_new_n870_), .Y(new_new_n871_));
  NO2        g0849(.A(new_new_n383_), .B(new_new_n290_), .Y(new_new_n872_));
  NA2        g0850(.A(new_new_n872_), .B(new_new_n704_), .Y(new_new_n873_));
  NA2        g0851(.A(new_new_n570_), .B(i_0_), .Y(new_new_n874_));
  NO3        g0852(.A(new_new_n874_), .B(new_new_n380_), .C(new_new_n90_), .Y(new_new_n875_));
  NO4        g0853(.A(new_new_n582_), .B(new_new_n220_), .C(new_new_n409_), .D(new_new_n401_), .Y(new_new_n876_));
  AOI210     g0854(.A0(new_new_n876_), .A1(i_11_), .B0(new_new_n875_), .Y(new_new_n877_));
  NA2        g0855(.A(new_new_n743_), .B(new_new_n322_), .Y(new_new_n878_));
  AOI210     g0856(.A0(new_new_n476_), .A1(new_new_n90_), .B0(new_new_n59_), .Y(new_new_n879_));
  NO2        g0857(.A(new_new_n879_), .B(new_new_n878_), .Y(new_new_n880_));
  NO2        g0858(.A(new_new_n257_), .B(new_new_n159_), .Y(new_new_n881_));
  NA2        g0859(.A(i_0_), .B(i_10_), .Y(new_new_n882_));
  INV        g0860(.A(new_new_n532_), .Y(new_new_n883_));
  NO4        g0861(.A(new_new_n119_), .B(new_new_n59_), .C(new_new_n661_), .D(i_5_), .Y(new_new_n884_));
  AO220      g0862(.A0(new_new_n884_), .A1(new_new_n883_), .B0(new_new_n881_), .B1(i_6_), .Y(new_new_n885_));
  AOI220     g0863(.A0(new_new_n325_), .A1(new_new_n102_), .B0(new_new_n187_), .B1(new_new_n85_), .Y(new_new_n886_));
  NA2        g0864(.A(new_new_n564_), .B(i_4_), .Y(new_new_n887_));
  NA2        g0865(.A(new_new_n190_), .B(new_new_n205_), .Y(new_new_n888_));
  OAI220     g0866(.A0(new_new_n888_), .A1(new_new_n878_), .B0(new_new_n887_), .B1(new_new_n886_), .Y(new_new_n889_));
  NO3        g0867(.A(new_new_n889_), .B(new_new_n885_), .C(new_new_n880_), .Y(new_new_n890_));
  NA4        g0868(.A(new_new_n890_), .B(new_new_n877_), .C(new_new_n873_), .D(new_new_n871_), .Y(new_new_n891_));
  NO2        g0869(.A(new_new_n107_), .B(new_new_n37_), .Y(new_new_n892_));
  NA2        g0870(.A(i_11_), .B(i_9_), .Y(new_new_n893_));
  NO3        g0871(.A(i_12_), .B(new_new_n893_), .C(new_new_n597_), .Y(new_new_n894_));
  AN2        g0872(.A(new_new_n894_), .B(new_new_n892_), .Y(new_new_n895_));
  NO2        g0873(.A(new_new_n49_), .B(i_7_), .Y(new_new_n896_));
  NA2        g0874(.A(new_new_n384_), .B(new_new_n183_), .Y(new_new_n897_));
  NA2        g0875(.A(new_new_n897_), .B(new_new_n166_), .Y(new_new_n898_));
  NO2        g0876(.A(new_new_n893_), .B(new_new_n74_), .Y(new_new_n899_));
  NO2        g0877(.A(new_new_n179_), .B(i_0_), .Y(new_new_n900_));
  INV        g0878(.A(new_new_n900_), .Y(new_new_n901_));
  NA2        g0879(.A(new_new_n465_), .B(new_new_n234_), .Y(new_new_n902_));
  AOI210     g0880(.A0(new_new_n366_), .A1(new_new_n42_), .B0(new_new_n398_), .Y(new_new_n903_));
  OAI220     g0881(.A0(new_new_n903_), .A1(new_new_n860_), .B0(new_new_n902_), .B1(new_new_n901_), .Y(new_new_n904_));
  NO3        g0882(.A(new_new_n904_), .B(new_new_n898_), .C(new_new_n895_), .Y(new_new_n905_));
  NA2        g0883(.A(new_new_n652_), .B(new_new_n126_), .Y(new_new_n906_));
  NO2        g0884(.A(i_6_), .B(new_new_n906_), .Y(new_new_n907_));
  NA2        g0885(.A(new_new_n175_), .B(new_new_n107_), .Y(new_new_n908_));
  INV        g0886(.A(new_new_n907_), .Y(new_new_n909_));
  NOi21      g0887(.An(i_7_), .B(i_5_), .Y(new_new_n910_));
  NOi31      g0888(.An(new_new_n910_), .B(i_0_), .C(new_new_n721_), .Y(new_new_n911_));
  NA3        g0889(.A(new_new_n911_), .B(new_new_n379_), .C(i_6_), .Y(new_new_n912_));
  BUFFER     g0890(.A(new_new_n912_), .Y(new_new_n913_));
  NO3        g0891(.A(new_new_n393_), .B(new_new_n358_), .C(new_new_n354_), .Y(new_new_n914_));
  NO2        g0892(.A(new_new_n267_), .B(new_new_n312_), .Y(new_new_n915_));
  NO2        g0893(.A(new_new_n721_), .B(new_new_n262_), .Y(new_new_n916_));
  AOI210     g0894(.A0(new_new_n916_), .A1(new_new_n915_), .B0(new_new_n914_), .Y(new_new_n917_));
  NA4        g0895(.A(new_new_n917_), .B(new_new_n913_), .C(new_new_n909_), .D(new_new_n905_), .Y(new_new_n918_));
  NO2        g0896(.A(new_new_n868_), .B(new_new_n243_), .Y(new_new_n919_));
  AN2        g0897(.A(new_new_n324_), .B(new_new_n322_), .Y(new_new_n920_));
  AN2        g0898(.A(new_new_n920_), .B(new_new_n864_), .Y(new_new_n921_));
  OAI210     g0899(.A0(new_new_n921_), .A1(new_new_n919_), .B0(i_10_), .Y(new_new_n922_));
  OA210      g0900(.A0(new_new_n465_), .A1(new_new_n229_), .B0(new_new_n464_), .Y(new_new_n923_));
  NO2        g0901(.A(new_new_n260_), .B(new_new_n47_), .Y(new_new_n924_));
  NA2        g0902(.A(new_new_n899_), .B(new_new_n301_), .Y(new_new_n925_));
  OAI210     g0903(.A0(new_new_n924_), .A1(new_new_n189_), .B0(new_new_n925_), .Y(new_new_n926_));
  NA2        g0904(.A(new_new_n926_), .B(new_new_n465_), .Y(new_new_n927_));
  NA2        g0905(.A(new_new_n96_), .B(new_new_n45_), .Y(new_new_n928_));
  NO2        g0906(.A(new_new_n76_), .B(new_new_n745_), .Y(new_new_n929_));
  AOI220     g0907(.A0(new_new_n929_), .A1(new_new_n928_), .B0(new_new_n178_), .B1(new_new_n590_), .Y(new_new_n930_));
  NO2        g0908(.A(new_new_n930_), .B(new_new_n48_), .Y(new_new_n931_));
  NO3        g0909(.A(new_new_n582_), .B(new_new_n353_), .C(new_new_n24_), .Y(new_new_n932_));
  AOI210     g0910(.A0(new_new_n694_), .A1(new_new_n541_), .B0(new_new_n932_), .Y(new_new_n933_));
  NAi21      g0911(.An(i_9_), .B(i_5_), .Y(new_new_n934_));
  NO2        g0912(.A(new_new_n934_), .B(new_new_n393_), .Y(new_new_n935_));
  NO2        g0913(.A(new_new_n593_), .B(new_new_n109_), .Y(new_new_n936_));
  AOI220     g0914(.A0(new_new_n936_), .A1(i_0_), .B0(new_new_n935_), .B1(new_new_n616_), .Y(new_new_n937_));
  OAI220     g0915(.A0(new_new_n937_), .A1(new_new_n87_), .B0(new_new_n933_), .B1(new_new_n176_), .Y(new_new_n938_));
  NO3        g0916(.A(new_new_n938_), .B(new_new_n931_), .C(new_new_n514_), .Y(new_new_n939_));
  NA3        g0917(.A(new_new_n939_), .B(new_new_n927_), .C(new_new_n922_), .Y(new_new_n940_));
  NO3        g0918(.A(new_new_n940_), .B(new_new_n918_), .C(new_new_n891_), .Y(new_new_n941_));
  NO2        g0919(.A(i_0_), .B(new_new_n721_), .Y(new_new_n942_));
  NA2        g0920(.A(new_new_n74_), .B(new_new_n45_), .Y(new_new_n943_));
  INV        g0921(.A(new_new_n943_), .Y(new_new_n944_));
  NO3        g0922(.A(new_new_n109_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n945_));
  AO220      g0923(.A0(new_new_n945_), .A1(new_new_n944_), .B0(new_new_n942_), .B1(new_new_n178_), .Y(new_new_n946_));
  AOI210     g0924(.A0(new_new_n795_), .A1(new_new_n681_), .B0(new_new_n908_), .Y(new_new_n947_));
  AOI210     g0925(.A0(new_new_n946_), .A1(new_new_n342_), .B0(new_new_n947_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n731_), .B(new_new_n151_), .Y(new_new_n949_));
  INV        g0927(.A(new_new_n949_), .Y(new_new_n950_));
  NA3        g0928(.A(new_new_n950_), .B(new_new_n668_), .C(new_new_n74_), .Y(new_new_n951_));
  NO2        g0929(.A(new_new_n813_), .B(new_new_n393_), .Y(new_new_n952_));
  NA3        g0930(.A(new_new_n841_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n953_));
  NA2        g0931(.A(new_new_n842_), .B(i_9_), .Y(new_new_n954_));
  NO2        g0932(.A(new_new_n953_), .B(new_new_n954_), .Y(new_new_n955_));
  OAI210     g0933(.A0(new_new_n247_), .A1(i_9_), .B0(new_new_n233_), .Y(new_new_n956_));
  AOI210     g0934(.A0(new_new_n956_), .A1(new_new_n874_), .B0(new_new_n159_), .Y(new_new_n957_));
  NO3        g0935(.A(new_new_n957_), .B(new_new_n955_), .C(new_new_n952_), .Y(new_new_n958_));
  NA3        g0936(.A(new_new_n958_), .B(new_new_n951_), .C(new_new_n948_), .Y(new_new_n959_));
  NA2        g0937(.A(new_new_n920_), .B(new_new_n368_), .Y(new_new_n960_));
  AOI210     g0938(.A0(new_new_n295_), .A1(new_new_n168_), .B0(new_new_n960_), .Y(new_new_n961_));
  NA3        g0939(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n962_));
  NA2        g0940(.A(new_new_n896_), .B(new_new_n481_), .Y(new_new_n963_));
  AOI210     g0941(.A0(new_new_n962_), .A1(new_new_n168_), .B0(new_new_n963_), .Y(new_new_n964_));
  NO2        g0942(.A(new_new_n964_), .B(new_new_n961_), .Y(new_new_n965_));
  NO3        g0943(.A(new_new_n882_), .B(new_new_n859_), .C(new_new_n192_), .Y(new_new_n966_));
  AOI220     g0944(.A0(new_new_n966_), .A1(i_11_), .B0(new_new_n565_), .B1(new_new_n76_), .Y(new_new_n967_));
  NO3        g0945(.A(new_new_n214_), .B(new_new_n378_), .C(i_0_), .Y(new_new_n968_));
  OAI210     g0946(.A0(new_new_n968_), .A1(new_new_n77_), .B0(i_13_), .Y(new_new_n969_));
  INV        g0947(.A(new_new_n223_), .Y(new_new_n970_));
  OAI220     g0948(.A0(new_new_n525_), .A1(new_new_n144_), .B0(new_new_n638_), .B1(new_new_n610_), .Y(new_new_n971_));
  NA3        g0949(.A(new_new_n971_), .B(new_new_n386_), .C(new_new_n970_), .Y(new_new_n972_));
  NA4        g0950(.A(new_new_n972_), .B(new_new_n969_), .C(new_new_n967_), .D(new_new_n965_), .Y(new_new_n973_));
  NO2        g0951(.A(new_new_n246_), .B(new_new_n96_), .Y(new_new_n974_));
  AOI210     g0952(.A0(new_new_n974_), .A1(new_new_n942_), .B0(new_new_n113_), .Y(new_new_n975_));
  AOI220     g0953(.A0(new_new_n910_), .A1(new_new_n481_), .B0(new_new_n841_), .B1(new_new_n169_), .Y(new_new_n976_));
  NA2        g0954(.A(new_new_n345_), .B(new_new_n180_), .Y(new_new_n977_));
  OA220      g0955(.A0(new_new_n977_), .A1(new_new_n976_), .B0(new_new_n975_), .B1(i_5_), .Y(new_new_n978_));
  AOI210     g0956(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n179_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n979_), .B(new_new_n923_), .Y(new_new_n980_));
  NA3        g0958(.A(new_new_n607_), .B(new_new_n187_), .C(new_new_n85_), .Y(new_new_n981_));
  NA2        g0959(.A(new_new_n981_), .B(new_new_n539_), .Y(new_new_n982_));
  NO3        g0960(.A(new_new_n851_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n983_));
  NA3        g0961(.A(new_new_n486_), .B(new_new_n479_), .C(new_new_n462_), .Y(new_new_n984_));
  NO3        g0962(.A(new_new_n984_), .B(new_new_n983_), .C(new_new_n982_), .Y(new_new_n985_));
  NA3        g0963(.A(new_new_n383_), .B(new_new_n175_), .C(new_new_n174_), .Y(new_new_n986_));
  NA3        g0964(.A(new_new_n896_), .B(new_new_n289_), .C(new_new_n233_), .Y(new_new_n987_));
  NA2        g0965(.A(new_new_n987_), .B(new_new_n986_), .Y(new_new_n988_));
  NO3        g0966(.A(new_new_n893_), .B(new_new_n223_), .C(new_new_n192_), .Y(new_new_n989_));
  NO2        g0967(.A(new_new_n989_), .B(new_new_n988_), .Y(new_new_n990_));
  NA4        g0968(.A(new_new_n990_), .B(new_new_n985_), .C(new_new_n980_), .D(new_new_n978_), .Y(new_new_n991_));
  INV        g0969(.A(new_new_n609_), .Y(new_new_n992_));
  NO3        g0970(.A(new_new_n992_), .B(new_new_n555_), .C(new_new_n339_), .Y(new_new_n993_));
  NO2        g0971(.A(new_new_n87_), .B(i_5_), .Y(new_new_n994_));
  NA3        g0972(.A(new_new_n842_), .B(new_new_n114_), .C(new_new_n129_), .Y(new_new_n995_));
  INV        g0973(.A(new_new_n995_), .Y(new_new_n996_));
  AOI210     g0974(.A0(new_new_n996_), .A1(new_new_n994_), .B0(new_new_n993_), .Y(new_new_n997_));
  NA3        g0975(.A(new_new_n301_), .B(i_5_), .C(new_new_n195_), .Y(new_new_n998_));
  NAi31      g0976(.An(new_new_n245_), .B(new_new_n998_), .C(new_new_n246_), .Y(new_new_n999_));
  NO4        g0977(.A(new_new_n243_), .B(new_new_n214_), .C(i_0_), .D(i_12_), .Y(new_new_n1000_));
  AOI220     g0978(.A0(new_new_n1000_), .A1(new_new_n999_), .B0(new_new_n789_), .B1(new_new_n180_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n910_), .B(new_new_n461_), .Y(new_new_n1002_));
  NA2        g0980(.A(new_new_n65_), .B(new_new_n105_), .Y(new_new_n1003_));
  OAI220     g0981(.A0(new_new_n1003_), .A1(new_new_n998_), .B0(new_new_n1002_), .B1(new_new_n669_), .Y(new_new_n1004_));
  NA2        g0982(.A(new_new_n1004_), .B(new_new_n900_), .Y(new_new_n1005_));
  NA3        g0983(.A(new_new_n1005_), .B(new_new_n1001_), .C(new_new_n997_), .Y(new_new_n1006_));
  NO4        g0984(.A(new_new_n1006_), .B(new_new_n991_), .C(new_new_n973_), .D(new_new_n959_), .Y(new_new_n1007_));
  OAI210     g0985(.A0(new_new_n816_), .A1(new_new_n809_), .B0(new_new_n37_), .Y(new_new_n1008_));
  NA2        g0986(.A(new_new_n1008_), .B(new_new_n605_), .Y(new_new_n1009_));
  NA2        g0987(.A(new_new_n1009_), .B(new_new_n210_), .Y(new_new_n1010_));
  OAI210     g0988(.A0(new_new_n609_), .A1(new_new_n607_), .B0(new_new_n311_), .Y(new_new_n1011_));
  NAi31      g0989(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n1012_));
  AOI210     g0990(.A0(new_new_n122_), .A1(new_new_n71_), .B0(new_new_n1012_), .Y(new_new_n1013_));
  INV        g0991(.A(new_new_n1013_), .Y(new_new_n1014_));
  NA2        g0992(.A(new_new_n1014_), .B(new_new_n1011_), .Y(new_new_n1015_));
  NO2        g0993(.A(new_new_n452_), .B(new_new_n273_), .Y(new_new_n1016_));
  NO4        g0994(.A(new_new_n236_), .B(new_new_n150_), .C(new_new_n672_), .D(new_new_n37_), .Y(new_new_n1017_));
  NO3        g0995(.A(new_new_n1017_), .B(new_new_n1016_), .C(new_new_n876_), .Y(new_new_n1018_));
  INV        g0996(.A(new_new_n1018_), .Y(new_new_n1019_));
  AOI210     g0997(.A0(new_new_n1015_), .A1(new_new_n49_), .B0(new_new_n1019_), .Y(new_new_n1020_));
  AOI210     g0998(.A0(new_new_n1020_), .A1(new_new_n1010_), .B0(new_new_n74_), .Y(new_new_n1021_));
  NO2        g0999(.A(new_new_n562_), .B(new_new_n375_), .Y(new_new_n1022_));
  NO2        g1000(.A(new_new_n1022_), .B(new_new_n751_), .Y(new_new_n1023_));
  AOI210     g1001(.A0(new_new_n979_), .A1(new_new_n896_), .B0(new_new_n911_), .Y(new_new_n1024_));
  NO2        g1002(.A(new_new_n1024_), .B(new_new_n672_), .Y(new_new_n1025_));
  NA2        g1003(.A(new_new_n267_), .B(new_new_n58_), .Y(new_new_n1026_));
  AOI220     g1004(.A0(new_new_n1026_), .A1(new_new_n77_), .B0(new_new_n340_), .B1(new_new_n259_), .Y(new_new_n1027_));
  NO2        g1005(.A(new_new_n1027_), .B(new_new_n240_), .Y(new_new_n1028_));
  NA3        g1006(.A(new_new_n100_), .B(new_new_n303_), .C(new_new_n31_), .Y(new_new_n1029_));
  INV        g1007(.A(new_new_n1029_), .Y(new_new_n1030_));
  NO3        g1008(.A(new_new_n1030_), .B(new_new_n1028_), .C(new_new_n1025_), .Y(new_new_n1031_));
  OAI210     g1009(.A0(new_new_n275_), .A1(new_new_n164_), .B0(new_new_n90_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n755_), .B(new_new_n289_), .C(new_new_n81_), .Y(new_new_n1033_));
  AOI210     g1011(.A0(new_new_n1033_), .A1(new_new_n1032_), .B0(i_11_), .Y(new_new_n1034_));
  NO3        g1012(.A(new_new_n60_), .B(new_new_n59_), .C(i_4_), .Y(new_new_n1035_));
  OAI210     g1013(.A0(new_new_n915_), .A1(new_new_n303_), .B0(new_new_n1035_), .Y(new_new_n1036_));
  NO2        g1014(.A(new_new_n1036_), .B(new_new_n721_), .Y(new_new_n1037_));
  NO4        g1015(.A(new_new_n934_), .B(new_new_n469_), .C(new_new_n256_), .D(new_new_n255_), .Y(new_new_n1038_));
  NO2        g1016(.A(new_new_n1038_), .B(new_new_n559_), .Y(new_new_n1039_));
  INV        g1017(.A(new_new_n359_), .Y(new_new_n1040_));
  AOI210     g1018(.A0(new_new_n1040_), .A1(new_new_n1039_), .B0(new_new_n41_), .Y(new_new_n1041_));
  NO3        g1019(.A(new_new_n1041_), .B(new_new_n1037_), .C(new_new_n1034_), .Y(new_new_n1042_));
  OAI210     g1020(.A0(new_new_n1031_), .A1(i_4_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  NO3        g1021(.A(new_new_n1043_), .B(new_new_n1023_), .C(new_new_n1021_), .Y(new_new_n1044_));
  NA4        g1022(.A(new_new_n1044_), .B(new_new_n1007_), .C(new_new_n941_), .D(new_new_n867_), .Y(mai4));
  INV        g1023(.A(new_new_n693_), .Y(new_new_n1048_));
  INV        g1024(.A(new_new_n476_), .Y(new_new_n1049_));
endmodule


