//Benchmark atmr_intb_466_0.5

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n200_, ori_ori_n204_, ori_ori_n205_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n261_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n347_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  INV        o007(.A(x03), .Y(ori_ori_n30_));
  NA2        o008(.A(x10), .B(ori_ori_n30_), .Y(ori_ori_n31_));
  INV        o009(.A(x04), .Y(ori_ori_n32_));
  INV        o010(.A(x08), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(x02), .Y(ori_ori_n34_));
  NA2        o012(.A(x08), .B(x03), .Y(ori_ori_n35_));
  AOI210     o013(.A0(ori_ori_n35_), .A1(ori_ori_n34_), .B0(ori_ori_n32_), .Y(ori_ori_n36_));
  INV        o014(.A(x05), .Y(ori_ori_n37_));
  NO2        o015(.A(ori_ori_n36_), .B(ori_ori_n26_), .Y(ori00));
  INV        o016(.A(x01), .Y(ori_ori_n39_));
  INV        o017(.A(x06), .Y(ori_ori_n40_));
  INV        o018(.A(x09), .Y(ori_ori_n41_));
  NO2        o019(.A(x10), .B(x02), .Y(ori_ori_n42_));
  NOi21      o020(.An(x01), .B(x09), .Y(ori_ori_n43_));
  INV        o021(.A(x00), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n41_), .B(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o023(.A(ori_ori_n45_), .B(ori_ori_n43_), .Y(ori_ori_n46_));
  NA2        o024(.A(x09), .B(ori_ori_n44_), .Y(ori_ori_n47_));
  INV        o025(.A(x07), .Y(ori_ori_n48_));
  INV        o026(.A(ori_ori_n46_), .Y(ori_ori_n49_));
  NA2        o027(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n50_));
  NA2        o028(.A(ori_ori_n50_), .B(ori_ori_n24_), .Y(ori_ori_n51_));
  NO2        o029(.A(ori_ori_n51_), .B(ori_ori_n49_), .Y(ori_ori_n52_));
  INV        o030(.A(ori_ori_n52_), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n53_), .B(x05), .Y(ori_ori_n54_));
  NA2        o032(.A(x09), .B(x05), .Y(ori_ori_n55_));
  NOi31      o033(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n56_));
  NO2        o034(.A(ori_ori_n33_), .B(x00), .Y(ori_ori_n57_));
  NO2        o035(.A(x08), .B(x01), .Y(ori_ori_n58_));
  OAI210     o036(.A0(ori_ori_n58_), .A1(ori_ori_n57_), .B0(ori_ori_n32_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n41_), .B(ori_ori_n33_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n59_), .B(x02), .Y(ori_ori_n61_));
  INV        o039(.A(ori_ori_n59_), .Y(ori_ori_n62_));
  NA2        o040(.A(x11), .B(x00), .Y(ori_ori_n63_));
  NO2        o041(.A(x11), .B(ori_ori_n39_), .Y(ori_ori_n64_));
  NOi21      o042(.An(ori_ori_n63_), .B(ori_ori_n64_), .Y(ori_ori_n65_));
  INV        o043(.A(ori_ori_n65_), .Y(ori_ori_n66_));
  NOi21      o044(.An(x01), .B(x10), .Y(ori_ori_n67_));
  NO2        o045(.A(ori_ori_n29_), .B(ori_ori_n44_), .Y(ori_ori_n68_));
  NO3        o046(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(x06), .Y(ori_ori_n69_));
  NA2        o047(.A(ori_ori_n69_), .B(ori_ori_n27_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n66_), .A1(x07), .B0(ori_ori_n70_), .Y(ori_ori_n71_));
  NO3        o049(.A(ori_ori_n71_), .B(ori_ori_n61_), .C(ori_ori_n54_), .Y(ori01));
  INV        o050(.A(x12), .Y(ori_ori_n73_));
  INV        o051(.A(x13), .Y(ori_ori_n74_));
  NO2        o052(.A(x10), .B(x01), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n43_), .B(x05), .Y(ori_ori_n76_));
  NOi21      o054(.An(ori_ori_n76_), .B(ori_ori_n45_), .Y(ori_ori_n77_));
  NO2        o055(.A(x04), .B(x05), .Y(ori_ori_n78_));
  NA2        o056(.A(ori_ori_n29_), .B(ori_ori_n39_), .Y(ori_ori_n79_));
  NA2        o057(.A(x10), .B(ori_ori_n44_), .Y(ori_ori_n80_));
  NA2        o058(.A(ori_ori_n80_), .B(ori_ori_n79_), .Y(ori_ori_n81_));
  NO2        o059(.A(ori_ori_n47_), .B(x05), .Y(ori_ori_n82_));
  NO3        o060(.A(ori_ori_n79_), .B(x06), .C(x03), .Y(ori_ori_n83_));
  INV        o061(.A(ori_ori_n83_), .Y(ori_ori_n84_));
  OAI210     o062(.A0(ori_ori_n58_), .A1(x13), .B0(ori_ori_n32_), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n86_));
  NO2        o064(.A(x09), .B(x05), .Y(ori_ori_n87_));
  NA2        o065(.A(ori_ori_n87_), .B(ori_ori_n39_), .Y(ori_ori_n88_));
  NA2        o066(.A(x09), .B(x00), .Y(ori_ori_n89_));
  NA2        o067(.A(ori_ori_n76_), .B(ori_ori_n89_), .Y(ori_ori_n90_));
  NO2        o068(.A(x03), .B(x02), .Y(ori_ori_n91_));
  NA2        o069(.A(ori_ori_n59_), .B(ori_ori_n74_), .Y(ori_ori_n92_));
  OAI210     o070(.A0(ori_ori_n92_), .A1(ori_ori_n77_), .B0(ori_ori_n91_), .Y(ori_ori_n93_));
  OAI210     o071(.A0(ori_ori_n84_), .A1(ori_ori_n23_), .B0(ori_ori_n93_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n95_));
  NO2        o073(.A(x13), .B(x08), .Y(ori_ori_n96_));
  INV        o074(.A(ori_ori_n68_), .Y(ori_ori_n97_));
  NOi21      o075(.An(x09), .B(x00), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n98_), .B(ori_ori_n39_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n99_), .B(ori_ori_n80_), .Y(ori_ori_n100_));
  NA2        o078(.A(x06), .B(x05), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n101_), .B(ori_ori_n73_), .Y(ori_ori_n102_));
  AOI210     o080(.A0(x10), .A1(ori_ori_n45_), .B0(ori_ori_n102_), .Y(ori_ori_n103_));
  NA2        o081(.A(ori_ori_n103_), .B(ori_ori_n100_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n74_), .B(x12), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n32_), .B(ori_ori_n30_), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n107_), .B(x02), .Y(ori_ori_n108_));
  NA2        o086(.A(ori_ori_n106_), .B(ori_ori_n104_), .Y(ori_ori_n109_));
  INV        o087(.A(ori_ori_n109_), .Y(ori_ori_n110_));
  AOI210     o088(.A0(ori_ori_n94_), .A1(ori_ori_n73_), .B0(ori_ori_n110_), .Y(ori_ori_n111_));
  NA2        o089(.A(ori_ori_n41_), .B(ori_ori_n39_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(ori_ori_n85_), .Y(ori_ori_n113_));
  NO2        o091(.A(x06), .B(x05), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n114_), .B(ori_ori_n113_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n115_), .B(x12), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n67_), .B(x06), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n117_), .B(ori_ori_n37_), .Y(ori_ori_n118_));
  INV        o096(.A(ori_ori_n86_), .Y(ori_ori_n119_));
  OAI210     o097(.A0(ori_ori_n119_), .A1(ori_ori_n118_), .B0(x02), .Y(ori_ori_n120_));
  AOI210     o098(.A0(ori_ori_n120_), .A1(ori_ori_n44_), .B0(ori_ori_n23_), .Y(ori_ori_n121_));
  OAI210     o099(.A0(ori_ori_n116_), .A1(ori_ori_n44_), .B0(ori_ori_n121_), .Y(ori_ori_n122_));
  INV        o100(.A(ori_ori_n86_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n31_), .B(x06), .Y(ori_ori_n124_));
  NOi21      o102(.An(x13), .B(x04), .Y(ori_ori_n125_));
  NO3        o103(.A(ori_ori_n125_), .B(ori_ori_n56_), .C(ori_ori_n98_), .Y(ori_ori_n126_));
  NO2        o104(.A(ori_ori_n126_), .B(x05), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n127_), .B(ori_ori_n124_), .Y(ori_ori_n128_));
  INV        o106(.A(ori_ori_n128_), .Y(ori_ori_n129_));
  INV        o107(.A(ori_ori_n64_), .Y(ori_ori_n130_));
  NA2        o108(.A(ori_ori_n23_), .B(ori_ori_n39_), .Y(ori_ori_n131_));
  NO2        o109(.A(ori_ori_n41_), .B(ori_ori_n33_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n29_), .B(ori_ori_n40_), .Y(ori_ori_n133_));
  NA2        o111(.A(x13), .B(ori_ori_n73_), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n102_), .B(ori_ori_n65_), .Y(ori_ori_n135_));
  INV        o113(.A(ori_ori_n135_), .Y(ori_ori_n136_));
  AOI210     o114(.A0(ori_ori_n64_), .A1(ori_ori_n129_), .B0(ori_ori_n136_), .Y(ori_ori_n137_));
  AOI210     o115(.A0(ori_ori_n137_), .A1(ori_ori_n122_), .B0(x07), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n55_), .B(ori_ori_n29_), .Y(ori_ori_n139_));
  NO2        o117(.A(ori_ori_n125_), .B(ori_ori_n98_), .Y(ori_ori_n140_));
  NO2        o118(.A(ori_ori_n140_), .B(ori_ori_n139_), .Y(ori_ori_n141_));
  NO2        o119(.A(x02), .B(ori_ori_n130_), .Y(ori_ori_n142_));
  AN2        o120(.A(ori_ori_n141_), .B(ori_ori_n142_), .Y(ori_ori_n143_));
  NOi21      o121(.An(ori_ori_n139_), .B(ori_ori_n117_), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n145_));
  NA2        o123(.A(ori_ori_n144_), .B(ori_ori_n145_), .Y(ori_ori_n146_));
  NO2        o124(.A(ori_ori_n45_), .B(x05), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n147_), .B(ori_ori_n97_), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n131_), .B(ori_ori_n28_), .Y(ori_ori_n149_));
  OAI210     o127(.A0(ori_ori_n148_), .A1(ori_ori_n123_), .B0(ori_ori_n149_), .Y(ori_ori_n150_));
  NA2        o128(.A(ori_ori_n150_), .B(ori_ori_n146_), .Y(ori_ori_n151_));
  NO3        o129(.A(ori_ori_n151_), .B(ori_ori_n143_), .C(ori_ori_n138_), .Y(ori_ori_n152_));
  OAI210     o130(.A0(ori_ori_n111_), .A1(ori_ori_n48_), .B0(ori_ori_n152_), .Y(ori02));
  NA2        o131(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n154_), .B(ori_ori_n40_), .Y(ori_ori_n155_));
  NO2        o133(.A(x05), .B(x02), .Y(ori_ori_n156_));
  OAI210     o134(.A0(ori_ori_n113_), .A1(ori_ori_n98_), .B0(ori_ori_n156_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n157_), .B(ori_ori_n86_), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n133_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n159_), .B(ori_ori_n127_), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n204_), .B(ori_ori_n68_), .Y(ori_ori_n161_));
  INV        o139(.A(ori_ori_n91_), .Y(ori_ori_n162_));
  NO2        o140(.A(ori_ori_n162_), .B(ori_ori_n81_), .Y(ori_ori_n163_));
  NA2        o141(.A(ori_ori_n163_), .B(x13), .Y(ori_ori_n164_));
  NA3        o142(.A(ori_ori_n164_), .B(ori_ori_n161_), .C(ori_ori_n160_), .Y(ori_ori_n165_));
  NO3        o143(.A(ori_ori_n165_), .B(ori_ori_n158_), .C(ori_ori_n155_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n205_), .B(ori_ori_n75_), .Y(ori_ori_n167_));
  NA2        o145(.A(x12), .B(ori_ori_n81_), .Y(ori_ori_n168_));
  NA3        o146(.A(ori_ori_n168_), .B(ori_ori_n167_), .C(ori_ori_n40_), .Y(ori_ori_n169_));
  INV        o147(.A(ori_ori_n107_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n31_), .B(x05), .Y(ori_ori_n171_));
  OAI210     o149(.A0(ori_ori_n170_), .A1(ori_ori_n46_), .B0(ori_ori_n171_), .Y(ori_ori_n172_));
  NA2        o150(.A(ori_ori_n172_), .B(x02), .Y(ori_ori_n173_));
  INV        o151(.A(ori_ori_n132_), .Y(ori_ori_n174_));
  NA2        o152(.A(ori_ori_n105_), .B(x04), .Y(ori_ori_n175_));
  NO3        o153(.A(ori_ori_n105_), .B(ori_ori_n95_), .C(ori_ori_n42_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n89_), .B(ori_ori_n73_), .Y(ori_ori_n177_));
  OAI210     o155(.A0(ori_ori_n177_), .A1(ori_ori_n99_), .B0(ori_ori_n176_), .Y(ori_ori_n178_));
  NA3        o156(.A(ori_ori_n178_), .B(ori_ori_n173_), .C(x06), .Y(ori_ori_n179_));
  NA2        o157(.A(x09), .B(x03), .Y(ori_ori_n180_));
  OAI220     o158(.A0(ori_ori_n180_), .A1(ori_ori_n80_), .B0(ori_ori_n112_), .B1(ori_ori_n50_), .Y(ori_ori_n181_));
  NO3        o159(.A(ori_ori_n76_), .B(ori_ori_n80_), .C(ori_ori_n35_), .Y(ori_ori_n182_));
  AO220      o160(.A0(ori_ori_n182_), .A1(x04), .B0(ori_ori_n181_), .B1(x05), .Y(ori_ori_n183_));
  AOI210     o161(.A0(ori_ori_n179_), .A1(ori_ori_n169_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  OAI210     o162(.A0(ori_ori_n166_), .A1(x12), .B0(ori_ori_n184_), .Y(ori03));
  AO210      o163(.A0(ori_ori_n174_), .A1(ori_ori_n60_), .B0(ori_ori_n175_), .Y(ori_ori_n186_));
  NA2        o164(.A(ori_ori_n105_), .B(ori_ori_n91_), .Y(ori_ori_n187_));
  NA3        o165(.A(ori_ori_n187_), .B(ori_ori_n186_), .C(ori_ori_n108_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n188_), .B(x05), .Y(ori_ori_n189_));
  INV        o167(.A(ori_ori_n78_), .Y(ori_ori_n190_));
  NO2        o168(.A(ori_ori_n190_), .B(ori_ori_n46_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n191_), .B(ori_ori_n73_), .Y(ori_ori_n192_));
  AOI210     o170(.A0(ori_ori_n88_), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n90_), .B(x13), .Y(ori_ori_n194_));
  OAI210     o172(.A0(ori_ori_n194_), .A1(ori_ori_n193_), .B0(x04), .Y(ori_ori_n195_));
  NO2        o173(.A(ori_ori_n73_), .B(ori_ori_n88_), .Y(ori_ori_n196_));
  OA210      o174(.A0(ori_ori_n96_), .A1(x12), .B0(ori_ori_n82_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n197_), .B(ori_ori_n196_), .Y(ori_ori_n198_));
  NA4        o176(.A(ori_ori_n198_), .B(ori_ori_n195_), .C(ori_ori_n192_), .D(ori_ori_n189_), .Y(ori04));
  NO2        o177(.A(ori_ori_n62_), .B(ori_ori_n36_), .Y(ori_ori_n200_));
  XO2        o178(.A(ori_ori_n200_), .B(ori_ori_n134_), .Y(ori05));
  INV        o179(.A(ori_ori_n88_), .Y(ori_ori_n204_));
  INV        o180(.A(x13), .Y(ori_ori_n205_));
  ZERO       o181(.Y(ori06));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  NO2        m032(.A(mai_mai_n54_), .B(mai_mai_n50_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  NA2        m040(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n63_), .B(mai_mai_n24_), .Y(mai_mai_n64_));
  OAI220     m042(.A0(mai_mai_n64_), .A1(mai_mai_n58_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n65_));
  NA2        m043(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n66_));
  OAI210     m044(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n66_), .Y(mai_mai_n67_));
  AOI220     m045(.A0(mai_mai_n67_), .A1(mai_mai_n59_), .B0(mai_mai_n65_), .B1(mai_mai_n31_), .Y(mai_mai_n68_));
  AOI210     m046(.A0(mai_mai_n68_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n69_));
  NA2        m047(.A(x09), .B(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x10), .B(x06), .Y(mai_mai_n71_));
  NA3        m049(.A(mai_mai_n71_), .B(mai_mai_n70_), .C(mai_mai_n28_), .Y(mai_mai_n72_));
  OAI210     m050(.A0(mai_mai_n72_), .A1(x11), .B0(x03), .Y(mai_mai_n73_));
  NOi31      m051(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n74_));
  NO2        m052(.A(mai_mai_n301_), .B(mai_mai_n24_), .Y(mai_mai_n75_));
  NA2        m053(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n48_), .B(mai_mai_n76_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n78_));
  NO2        m056(.A(x08), .B(x01), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n79_), .A1(mai_mai_n78_), .B0(mai_mai_n35_), .Y(mai_mai_n80_));
  NO3        m058(.A(mai_mai_n80_), .B(mai_mai_n77_), .C(mai_mai_n75_), .Y(mai_mai_n81_));
  AN2        m059(.A(mai_mai_n81_), .B(mai_mai_n73_), .Y(mai_mai_n82_));
  INV        m060(.A(mai_mai_n80_), .Y(mai_mai_n83_));
  NO2        m061(.A(x06), .B(x05), .Y(mai_mai_n84_));
  NA2        m062(.A(x11), .B(x00), .Y(mai_mai_n85_));
  NO2        m063(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n86_));
  NOi21      m064(.An(mai_mai_n85_), .B(mai_mai_n86_), .Y(mai_mai_n87_));
  AOI210     m065(.A0(mai_mai_n84_), .A1(mai_mai_n83_), .B0(mai_mai_n87_), .Y(mai_mai_n88_));
  NOi21      m066(.An(x01), .B(x10), .Y(mai_mai_n89_));
  NO2        m067(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n90_));
  NO3        m068(.A(mai_mai_n90_), .B(mai_mai_n89_), .C(x06), .Y(mai_mai_n91_));
  NA2        m069(.A(mai_mai_n91_), .B(mai_mai_n27_), .Y(mai_mai_n92_));
  OAI210     m070(.A0(mai_mai_n88_), .A1(x07), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  NO3        m071(.A(mai_mai_n93_), .B(mai_mai_n82_), .C(mai_mai_n69_), .Y(mai01));
  INV        m072(.A(x12), .Y(mai_mai_n95_));
  INV        m073(.A(x13), .Y(mai_mai_n96_));
  NA2        m074(.A(x08), .B(x04), .Y(mai_mai_n97_));
  NA2        m075(.A(mai_mai_n89_), .B(mai_mai_n28_), .Y(mai_mai_n98_));
  NO2        m076(.A(x10), .B(x01), .Y(mai_mai_n99_));
  NO2        m077(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n100_));
  NO2        m078(.A(mai_mai_n100_), .B(mai_mai_n99_), .Y(mai_mai_n101_));
  NA2        m079(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(mai_mai_n36_), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n104_));
  NO2        m082(.A(mai_mai_n96_), .B(mai_mai_n36_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n106_));
  NA2        m084(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n107_), .B(x01), .Y(mai_mai_n108_));
  NA2        m086(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n110_));
  NO2        m088(.A(x06), .B(x03), .Y(mai_mai_n111_));
  NO3        m089(.A(mai_mai_n111_), .B(mai_mai_n303_), .C(mai_mai_n103_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n114_));
  AOI210     m092(.A0(mai_mai_n114_), .A1(mai_mai_n49_), .B0(mai_mai_n113_), .Y(mai_mai_n115_));
  NO2        m093(.A(x09), .B(x05), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(mai_mai_n47_), .Y(mai_mai_n117_));
  NO2        m095(.A(mai_mai_n101_), .B(mai_mai_n49_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n118_), .B(mai_mai_n115_), .Y(mai_mai_n119_));
  OR2        m097(.A(mai_mai_n119_), .B(x11), .Y(mai_mai_n120_));
  OAI210     m098(.A0(mai_mai_n112_), .A1(mai_mai_n23_), .B0(mai_mai_n120_), .Y(mai_mai_n121_));
  NA2        m099(.A(mai_mai_n101_), .B(mai_mai_n40_), .Y(mai_mai_n122_));
  NAi21      m100(.An(x06), .B(x10), .Y(mai_mai_n123_));
  NOi21      m101(.An(x01), .B(x13), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n125_));
  NO2        m103(.A(mai_mai_n122_), .B(mai_mai_n41_), .Y(mai_mai_n126_));
  NO2        m104(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n127_));
  NA2        m105(.A(mai_mai_n96_), .B(x01), .Y(mai_mai_n128_));
  NO2        m106(.A(mai_mai_n128_), .B(x08), .Y(mai_mai_n129_));
  OAI210     m107(.A0(x05), .A1(mai_mai_n129_), .B0(mai_mai_n51_), .Y(mai_mai_n130_));
  AOI210     m108(.A0(mai_mai_n130_), .A1(mai_mai_n127_), .B0(mai_mai_n48_), .Y(mai_mai_n131_));
  OAI210     m109(.A0(mai_mai_n131_), .A1(mai_mai_n126_), .B0(x02), .Y(mai_mai_n132_));
  NA2        m110(.A(x04), .B(x02), .Y(mai_mai_n133_));
  NA2        m111(.A(x10), .B(x05), .Y(mai_mai_n134_));
  NO2        m112(.A(mai_mai_n104_), .B(x08), .Y(mai_mai_n135_));
  NA3        m113(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n51_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n89_), .B(x05), .Y(mai_mai_n137_));
  OAI210     m115(.A0(mai_mai_n137_), .A1(mai_mai_n105_), .B0(mai_mai_n136_), .Y(mai_mai_n138_));
  AOI210     m116(.A0(mai_mai_n135_), .A1(x06), .B0(mai_mai_n138_), .Y(mai_mai_n139_));
  NO2        m117(.A(mai_mai_n139_), .B(x11), .Y(mai_mai_n140_));
  NAi21      m118(.An(mai_mai_n133_), .B(mai_mai_n140_), .Y(mai_mai_n141_));
  NAi21      m119(.An(x13), .B(x00), .Y(mai_mai_n142_));
  AOI210     m120(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n142_), .Y(mai_mai_n143_));
  AOI220     m121(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n144_));
  AN2        m122(.A(x04), .B(mai_mai_n143_), .Y(mai_mai_n145_));
  INV        m123(.A(x06), .Y(mai_mai_n146_));
  NO2        m124(.A(mai_mai_n142_), .B(mai_mai_n36_), .Y(mai_mai_n147_));
  OAI210     m125(.A0(mai_mai_n147_), .A1(mai_mai_n145_), .B0(x11), .Y(mai_mai_n148_));
  NO2        m126(.A(mai_mai_n78_), .B(mai_mai_n47_), .Y(mai_mai_n149_));
  NA2        m127(.A(mai_mai_n149_), .B(mai_mai_n107_), .Y(mai_mai_n150_));
  NA2        m128(.A(mai_mai_n95_), .B(mai_mai_n150_), .Y(mai_mai_n151_));
  NO2        m129(.A(mai_mai_n96_), .B(x12), .Y(mai_mai_n152_));
  AOI210     m130(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n152_), .Y(mai_mai_n153_));
  NO2        m131(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n154_));
  NA2        m132(.A(mai_mai_n153_), .B(mai_mai_n151_), .Y(mai_mai_n155_));
  NA4        m133(.A(mai_mai_n155_), .B(mai_mai_n148_), .C(mai_mai_n141_), .D(mai_mai_n132_), .Y(mai_mai_n156_));
  AOI210     m134(.A0(mai_mai_n121_), .A1(mai_mai_n95_), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  INV        m135(.A(mai_mai_n74_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n125_), .B(mai_mai_n57_), .Y(mai_mai_n159_));
  NA2        m137(.A(mai_mai_n159_), .B(mai_mai_n158_), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n161_));
  NA2        m139(.A(mai_mai_n56_), .B(x02), .Y(mai_mai_n162_));
  AOI210     m140(.A0(mai_mai_n162_), .A1(mai_mai_n160_), .B0(mai_mai_n23_), .Y(mai_mai_n163_));
  INV        m141(.A(mai_mai_n163_), .Y(mai_mai_n164_));
  INV        m142(.A(mai_mai_n114_), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n96_), .B(x03), .Y(mai_mai_n167_));
  OAI210     m145(.A0(x03), .A1(mai_mai_n165_), .B0(mai_mai_n123_), .Y(mai_mai_n168_));
  INV        m146(.A(mai_mai_n86_), .Y(mai_mai_n169_));
  NO2        m147(.A(mai_mai_n169_), .B(x12), .Y(mai_mai_n170_));
  OAI210     m148(.A0(x08), .A1(x04), .B0(mai_mai_n143_), .Y(mai_mai_n171_));
  AOI210     m149(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n172_));
  NO2        m150(.A(mai_mai_n172_), .B(mai_mai_n41_), .Y(mai_mai_n173_));
  NA2        m151(.A(mai_mai_n97_), .B(mai_mai_n71_), .Y(mai_mai_n174_));
  NO2        m152(.A(mai_mai_n174_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NA2        m153(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n176_));
  NA2        m154(.A(mai_mai_n176_), .B(x03), .Y(mai_mai_n177_));
  OA210      m155(.A0(mai_mai_n177_), .A1(mai_mai_n175_), .B0(mai_mai_n171_), .Y(mai_mai_n178_));
  NA2        m156(.A(x13), .B(mai_mai_n95_), .Y(mai_mai_n179_));
  NA2        m157(.A(x12), .B(mai_mai_n87_), .Y(mai_mai_n180_));
  OAI210     m158(.A0(mai_mai_n178_), .A1(x01), .B0(mai_mai_n180_), .Y(mai_mai_n181_));
  AOI210     m159(.A0(mai_mai_n170_), .A1(mai_mai_n168_), .B0(mai_mai_n181_), .Y(mai_mai_n182_));
  AOI210     m160(.A0(mai_mai_n182_), .A1(mai_mai_n164_), .B0(x07), .Y(mai_mai_n183_));
  NA2        m161(.A(mai_mai_n70_), .B(mai_mai_n29_), .Y(mai_mai_n184_));
  INV        m162(.A(mai_mai_n184_), .Y(mai_mai_n185_));
  NO2        m163(.A(x12), .B(x02), .Y(mai_mai_n186_));
  INV        m164(.A(mai_mai_n186_), .Y(mai_mai_n187_));
  NO2        m165(.A(mai_mai_n187_), .B(mai_mai_n169_), .Y(mai_mai_n188_));
  OA210      m166(.A0(mai_mai_n31_), .A1(mai_mai_n185_), .B0(mai_mai_n188_), .Y(mai_mai_n189_));
  NA2        m167(.A(mai_mai_n96_), .B(x04), .Y(mai_mai_n190_));
  INV        m168(.A(mai_mai_n97_), .Y(mai_mai_n191_));
  INV        m169(.A(mai_mai_n25_), .Y(mai_mai_n192_));
  NA2        m170(.A(mai_mai_n191_), .B(mai_mai_n192_), .Y(mai_mai_n193_));
  NO2        m171(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n194_));
  NO3        m172(.A(mai_mai_n194_), .B(mai_mai_n161_), .C(mai_mai_n146_), .Y(mai_mai_n195_));
  NO2        m173(.A(x01), .B(mai_mai_n28_), .Y(mai_mai_n196_));
  OAI210     m174(.A0(mai_mai_n195_), .A1(mai_mai_n165_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  NA2        m175(.A(mai_mai_n197_), .B(mai_mai_n193_), .Y(mai_mai_n198_));
  NO3        m176(.A(mai_mai_n198_), .B(mai_mai_n189_), .C(mai_mai_n183_), .Y(mai_mai_n199_));
  OAI210     m177(.A0(mai_mai_n157_), .A1(mai_mai_n61_), .B0(mai_mai_n199_), .Y(mai02));
  INV        m178(.A(mai_mai_n109_), .Y(mai_mai_n201_));
  NA3        m179(.A(x04), .B(x10), .C(mai_mai_n56_), .Y(mai_mai_n202_));
  OAI210     m180(.A0(x00), .A1(mai_mai_n32_), .B0(mai_mai_n202_), .Y(mai_mai_n203_));
  OAI210     m181(.A0(mai_mai_n203_), .A1(mai_mai_n201_), .B0(mai_mai_n134_), .Y(mai_mai_n204_));
  INV        m182(.A(mai_mai_n134_), .Y(mai_mai_n205_));
  AOI210     m183(.A0(x04), .A1(x08), .B0(mai_mai_n161_), .Y(mai_mai_n206_));
  OAI220     m184(.A0(mai_mai_n206_), .A1(mai_mai_n96_), .B0(mai_mai_n80_), .B1(mai_mai_n51_), .Y(mai_mai_n207_));
  NA2        m185(.A(mai_mai_n207_), .B(mai_mai_n205_), .Y(mai_mai_n208_));
  AOI210     m186(.A0(mai_mai_n208_), .A1(mai_mai_n204_), .B0(mai_mai_n48_), .Y(mai_mai_n209_));
  NOi21      m187(.An(x04), .B(x08), .Y(mai_mai_n210_));
  INV        m188(.A(mai_mai_n210_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n211_), .B(mai_mai_n114_), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n176_), .B(mai_mai_n47_), .Y(mai_mai_n213_));
  INV        m191(.A(mai_mai_n213_), .Y(mai_mai_n214_));
  OAI210     m192(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n215_));
  AN2        m193(.A(x08), .B(mai_mai_n117_), .Y(mai_mai_n216_));
  AOI210     m194(.A0(mai_mai_n216_), .A1(x04), .B0(mai_mai_n215_), .Y(mai_mai_n217_));
  OAI210     m195(.A0(mai_mai_n217_), .A1(mai_mai_n167_), .B0(mai_mai_n90_), .Y(mai_mai_n218_));
  NA3        m196(.A(mai_mai_n90_), .B(mai_mai_n79_), .C(mai_mai_n166_), .Y(mai_mai_n219_));
  NO2        m197(.A(mai_mai_n219_), .B(x04), .Y(mai_mai_n220_));
  INV        m198(.A(mai_mai_n98_), .Y(mai_mai_n221_));
  NO2        m199(.A(mai_mai_n221_), .B(mai_mai_n220_), .Y(mai_mai_n222_));
  NA3        m200(.A(mai_mai_n222_), .B(mai_mai_n218_), .C(mai_mai_n214_), .Y(mai_mai_n223_));
  NO3        m201(.A(mai_mai_n223_), .B(mai_mai_n212_), .C(mai_mai_n209_), .Y(mai_mai_n224_));
  NA2        m202(.A(mai_mai_n113_), .B(x03), .Y(mai_mai_n225_));
  OAI210     m203(.A0(mai_mai_n35_), .A1(mai_mai_n194_), .B0(mai_mai_n225_), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n226_), .B(mai_mai_n99_), .Y(mai_mai_n227_));
  NA2        m205(.A(mai_mai_n133_), .B(mai_mai_n128_), .Y(mai_mai_n228_));
  AN2        m206(.A(mai_mai_n228_), .B(mai_mai_n135_), .Y(mai_mai_n229_));
  OAI220     m207(.A0(mai_mai_n190_), .A1(x09), .B0(mai_mai_n109_), .B1(mai_mai_n28_), .Y(mai_mai_n230_));
  OAI210     m208(.A0(mai_mai_n230_), .A1(mai_mai_n229_), .B0(mai_mai_n100_), .Y(mai_mai_n231_));
  NA2        m209(.A(mai_mai_n190_), .B(mai_mai_n95_), .Y(mai_mai_n232_));
  NA2        m210(.A(mai_mai_n95_), .B(mai_mai_n41_), .Y(mai_mai_n233_));
  NA3        m211(.A(mai_mai_n233_), .B(mai_mai_n232_), .C(mai_mai_n108_), .Y(mai_mai_n234_));
  NA4        m212(.A(mai_mai_n234_), .B(mai_mai_n231_), .C(mai_mai_n227_), .D(mai_mai_n48_), .Y(mai_mai_n235_));
  INV        m213(.A(mai_mai_n154_), .Y(mai_mai_n236_));
  OAI220     m214(.A0(mai_mai_n302_), .A1(mai_mai_n31_), .B0(mai_mai_n236_), .B1(mai_mai_n59_), .Y(mai_mai_n237_));
  NA2        m215(.A(mai_mai_n237_), .B(x02), .Y(mai_mai_n238_));
  NA2        m216(.A(mai_mai_n152_), .B(x04), .Y(mai_mai_n239_));
  NO2        m217(.A(mai_mai_n144_), .B(mai_mai_n31_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n240_), .B(mai_mai_n90_), .Y(mai_mai_n241_));
  NO3        m219(.A(mai_mai_n152_), .B(mai_mai_n127_), .C(mai_mai_n52_), .Y(mai_mai_n242_));
  OAI210     m220(.A0(x12), .A1(mai_mai_n149_), .B0(mai_mai_n242_), .Y(mai_mai_n243_));
  NA4        m221(.A(mai_mai_n243_), .B(mai_mai_n241_), .C(mai_mai_n238_), .D(x06), .Y(mai_mai_n244_));
  NO2        m222(.A(x09), .B(mai_mai_n63_), .Y(mai_mai_n245_));
  NA2        m223(.A(mai_mai_n242_), .B(x05), .Y(mai_mai_n246_));
  INV        m224(.A(mai_mai_n246_), .Y(mai_mai_n247_));
  AO220      m225(.A0(mai_mai_n247_), .A1(x04), .B0(mai_mai_n245_), .B1(x05), .Y(mai_mai_n248_));
  AOI210     m226(.A0(mai_mai_n244_), .A1(mai_mai_n235_), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  OAI210     m227(.A0(mai_mai_n224_), .A1(x12), .B0(mai_mai_n249_), .Y(mai03));
  OR2        m228(.A(mai_mai_n42_), .B(mai_mai_n166_), .Y(mai_mai_n251_));
  INV        m229(.A(mai_mai_n251_), .Y(mai_mai_n252_));
  NA2        m230(.A(mai_mai_n252_), .B(x05), .Y(mai_mai_n253_));
  OAI210     m231(.A0(x13), .A1(x05), .B0(mai_mai_n95_), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n104_), .B(x04), .Y(mai_mai_n255_));
  NO3        m233(.A(mai_mai_n233_), .B(mai_mai_n80_), .C(mai_mai_n59_), .Y(mai_mai_n256_));
  AOI210     m234(.A0(mai_mai_n36_), .A1(mai_mai_n95_), .B0(mai_mai_n117_), .Y(mai_mai_n257_));
  OA210      m235(.A0(mai_mai_n129_), .A1(x12), .B0(mai_mai_n110_), .Y(mai_mai_n258_));
  NO3        m236(.A(mai_mai_n258_), .B(mai_mai_n257_), .C(mai_mai_n256_), .Y(mai_mai_n259_));
  NA4        m237(.A(mai_mai_n259_), .B(mai_mai_n255_), .C(mai_mai_n254_), .D(mai_mai_n253_), .Y(mai04));
  NO2        m238(.A(mai_mai_n83_), .B(mai_mai_n39_), .Y(mai_mai_n261_));
  XO2        m239(.A(mai_mai_n261_), .B(mai_mai_n179_), .Y(mai05));
  NA2        m240(.A(mai_mai_n70_), .B(mai_mai_n52_), .Y(mai_mai_n263_));
  AOI210     m241(.A0(mai_mai_n263_), .A1(mai_mai_n215_), .B0(mai_mai_n25_), .Y(mai_mai_n264_));
  NA3        m242(.A(mai_mai_n114_), .B(mai_mai_n109_), .C(mai_mai_n31_), .Y(mai_mai_n265_));
  INV        m243(.A(mai_mai_n84_), .Y(mai_mai_n266_));
  AOI210     m244(.A0(mai_mai_n266_), .A1(mai_mai_n265_), .B0(mai_mai_n24_), .Y(mai_mai_n267_));
  OAI210     m245(.A0(mai_mai_n267_), .A1(mai_mai_n264_), .B0(mai_mai_n95_), .Y(mai_mai_n268_));
  NA2        m246(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n269_));
  NA2        m247(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n270_));
  NA2        m248(.A(mai_mai_n184_), .B(x03), .Y(mai_mai_n271_));
  OAI220     m249(.A0(mai_mai_n271_), .A1(mai_mai_n270_), .B0(mai_mai_n269_), .B1(mai_mai_n76_), .Y(mai_mai_n272_));
  OAI210     m250(.A0(mai_mai_n26_), .A1(mai_mai_n95_), .B0(x07), .Y(mai_mai_n273_));
  AOI210     m251(.A0(mai_mai_n272_), .A1(x06), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  NA2        m252(.A(mai_mai_n33_), .B(mai_mai_n95_), .Y(mai_mai_n275_));
  AOI210     m253(.A0(mai_mai_n275_), .A1(mai_mai_n86_), .B0(x07), .Y(mai_mai_n276_));
  AOI210     m254(.A0(mai_mai_n274_), .A1(mai_mai_n268_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  INV        m255(.A(mai_mai_n113_), .Y(mai_mai_n278_));
  OR2        m256(.A(mai_mai_n278_), .B(x03), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n116_), .B(mai_mai_n28_), .Y(mai_mai_n280_));
  AOI210     m258(.A0(mai_mai_n280_), .A1(mai_mai_n279_), .B0(mai_mai_n47_), .Y(mai_mai_n281_));
  NA2        m259(.A(mai_mai_n281_), .B(mai_mai_n96_), .Y(mai_mai_n282_));
  AOI210     m260(.A0(mai_mai_n239_), .A1(mai_mai_n102_), .B0(mai_mai_n186_), .Y(mai_mai_n283_));
  NOi21      m261(.An(mai_mai_n225_), .B(mai_mai_n110_), .Y(mai_mai_n284_));
  NO2        m262(.A(mai_mai_n284_), .B(mai_mai_n187_), .Y(mai_mai_n285_));
  OAI210     m263(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n286_));
  AOI210     m264(.A0(mai_mai_n179_), .A1(mai_mai_n47_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  NO4        m265(.A(mai_mai_n287_), .B(mai_mai_n285_), .C(mai_mai_n283_), .D(x08), .Y(mai_mai_n288_));
  NA3        m266(.A(mai_mai_n236_), .B(mai_mai_n106_), .C(x12), .Y(mai_mai_n289_));
  AO210      m267(.A0(mai_mai_n236_), .A1(mai_mai_n106_), .B0(mai_mai_n179_), .Y(mai_mai_n290_));
  NA3        m268(.A(mai_mai_n290_), .B(mai_mai_n289_), .C(x08), .Y(mai_mai_n291_));
  INV        m269(.A(mai_mai_n291_), .Y(mai_mai_n292_));
  AOI210     m270(.A0(mai_mai_n288_), .A1(mai_mai_n282_), .B0(mai_mai_n292_), .Y(mai_mai_n293_));
  NA2        m271(.A(mai_mai_n275_), .B(mai_mai_n61_), .Y(mai_mai_n294_));
  NO2        m272(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n295_));
  NA2        m273(.A(mai_mai_n295_), .B(mai_mai_n95_), .Y(mai_mai_n296_));
  OAI210     m274(.A0(mai_mai_n294_), .A1(mai_mai_n85_), .B0(mai_mai_n296_), .Y(mai_mai_n297_));
  NO4        m275(.A(mai_mai_n297_), .B(mai_mai_n304_), .C(mai_mai_n293_), .D(mai_mai_n277_), .Y(mai06));
  INV        m276(.A(x07), .Y(mai_mai_n301_));
  INV        m277(.A(x05), .Y(mai_mai_n302_));
  INV        m278(.A(mai_mai_n71_), .Y(mai_mai_n303_));
  INV        m279(.A(x14), .Y(mai_mai_n304_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  INV        u003(.A(x02), .Y(men_men_n26_));
  INV        u004(.A(x10), .Y(men_men_n27_));
  NA2        u005(.A(men_men_n27_), .B(men_men_n26_), .Y(men_men_n28_));
  INV        u006(.A(x03), .Y(men_men_n29_));
  NA2        u007(.A(x10), .B(men_men_n29_), .Y(men_men_n30_));
  NA3        u008(.A(men_men_n30_), .B(men_men_n28_), .C(x06), .Y(men_men_n31_));
  INV        u009(.A(men_men_n31_), .Y(men_men_n32_));
  INV        u010(.A(x04), .Y(men_men_n33_));
  INV        u011(.A(x08), .Y(men_men_n34_));
  NA2        u012(.A(men_men_n34_), .B(x02), .Y(men_men_n35_));
  NA2        u013(.A(x08), .B(x03), .Y(men_men_n36_));
  AOI210     u014(.A0(men_men_n36_), .A1(men_men_n35_), .B0(men_men_n33_), .Y(men_men_n37_));
  NA2        u015(.A(x09), .B(men_men_n29_), .Y(men_men_n38_));
  INV        u016(.A(x05), .Y(men_men_n39_));
  NO2        u017(.A(x09), .B(x02), .Y(men_men_n40_));
  NO2        u018(.A(men_men_n40_), .B(men_men_n39_), .Y(men_men_n41_));
  NA2        u019(.A(men_men_n41_), .B(men_men_n38_), .Y(men_men_n42_));
  INV        u020(.A(men_men_n42_), .Y(men_men_n43_));
  NO3        u021(.A(men_men_n43_), .B(men_men_n37_), .C(men_men_n32_), .Y(men00));
  INV        u022(.A(x01), .Y(men_men_n45_));
  INV        u023(.A(x06), .Y(men_men_n46_));
  NO2        u024(.A(x06), .B(x11), .Y(men_men_n47_));
  INV        u025(.A(x09), .Y(men_men_n48_));
  NO2        u026(.A(x10), .B(x02), .Y(men_men_n49_));
  NO2        u027(.A(x10), .B(x07), .Y(men_men_n50_));
  OAI210     u028(.A0(men_men_n50_), .A1(men_men_n47_), .B0(men_men_n45_), .Y(men_men_n51_));
  NOi21      u029(.An(x01), .B(x09), .Y(men_men_n52_));
  INV        u030(.A(x00), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n48_), .B(men_men_n53_), .Y(men_men_n54_));
  NO2        u032(.A(men_men_n54_), .B(men_men_n52_), .Y(men_men_n55_));
  NA2        u033(.A(x09), .B(men_men_n53_), .Y(men_men_n56_));
  INV        u034(.A(x07), .Y(men_men_n57_));
  NA2        u035(.A(men_men_n57_), .B(men_men_n46_), .Y(men_men_n58_));
  OAI210     u036(.A0(men_men_n28_), .A1(x11), .B0(men_men_n58_), .Y(men_men_n59_));
  AOI220     u037(.A0(men_men_n59_), .A1(men_men_n55_), .B0(men_men_n55_), .B1(men_men_n29_), .Y(men_men_n60_));
  AOI210     u038(.A0(men_men_n60_), .A1(men_men_n51_), .B0(x05), .Y(men_men_n61_));
  NA2        u039(.A(x10), .B(x09), .Y(men_men_n62_));
  NA2        u040(.A(x09), .B(x05), .Y(men_men_n63_));
  NA2        u041(.A(x10), .B(x06), .Y(men_men_n64_));
  NA3        u042(.A(men_men_n64_), .B(men_men_n63_), .C(men_men_n26_), .Y(men_men_n65_));
  NO2        u043(.A(men_men_n57_), .B(men_men_n39_), .Y(men_men_n66_));
  OAI210     u044(.A0(men_men_n65_), .A1(x07), .B0(x03), .Y(men_men_n67_));
  NOi31      u045(.An(x08), .B(x04), .C(x00), .Y(men_men_n68_));
  NO2        u046(.A(x09), .B(men_men_n39_), .Y(men_men_n69_));
  NO2        u047(.A(men_men_n69_), .B(men_men_n34_), .Y(men_men_n70_));
  OAI210     u048(.A0(men_men_n69_), .A1(men_men_n27_), .B0(x02), .Y(men_men_n71_));
  AOI210     u049(.A0(men_men_n70_), .A1(men_men_n46_), .B0(men_men_n71_), .Y(men_men_n72_));
  NO2        u050(.A(men_men_n34_), .B(x00), .Y(men_men_n73_));
  NO2        u051(.A(x08), .B(x01), .Y(men_men_n74_));
  OAI210     u052(.A0(men_men_n74_), .A1(men_men_n73_), .B0(men_men_n33_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n75_), .B(men_men_n72_), .Y(men_men_n76_));
  AN2        u054(.A(men_men_n76_), .B(men_men_n67_), .Y(men_men_n77_));
  INV        u055(.A(men_men_n75_), .Y(men_men_n78_));
  NO2        u056(.A(x06), .B(x05), .Y(men_men_n79_));
  NA2        u057(.A(x11), .B(x00), .Y(men_men_n80_));
  NO2        u058(.A(x11), .B(men_men_n45_), .Y(men_men_n81_));
  NOi21      u059(.An(men_men_n80_), .B(men_men_n81_), .Y(men_men_n82_));
  AOI210     u060(.A0(men_men_n79_), .A1(men_men_n78_), .B0(men_men_n82_), .Y(men_men_n83_));
  NOi21      u061(.An(x01), .B(x10), .Y(men_men_n84_));
  NO2        u062(.A(men_men_n27_), .B(men_men_n53_), .Y(men_men_n85_));
  NO2        u063(.A(men_men_n83_), .B(x07), .Y(men_men_n86_));
  NO3        u064(.A(men_men_n86_), .B(men_men_n77_), .C(men_men_n61_), .Y(men01));
  INV        u065(.A(x12), .Y(men_men_n88_));
  INV        u066(.A(x13), .Y(men_men_n89_));
  NA2        u067(.A(x08), .B(x04), .Y(men_men_n90_));
  NA2        u068(.A(men_men_n84_), .B(men_men_n26_), .Y(men_men_n91_));
  NO2        u069(.A(men_men_n91_), .B(men_men_n63_), .Y(men_men_n92_));
  NO2        u070(.A(x10), .B(x01), .Y(men_men_n93_));
  NO2        u071(.A(men_men_n27_), .B(x00), .Y(men_men_n94_));
  NO2        u072(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u073(.A(x04), .B(men_men_n26_), .Y(men_men_n96_));
  NO3        u074(.A(men_men_n96_), .B(men_men_n34_), .C(men_men_n39_), .Y(men_men_n97_));
  AOI210     u075(.A0(men_men_n97_), .A1(men_men_n95_), .B0(men_men_n92_), .Y(men_men_n98_));
  NO2        u076(.A(men_men_n98_), .B(men_men_n89_), .Y(men_men_n99_));
  NO2        u077(.A(men_men_n52_), .B(x05), .Y(men_men_n100_));
  NOi21      u078(.An(men_men_n100_), .B(men_men_n54_), .Y(men_men_n101_));
  NO2        u079(.A(men_men_n33_), .B(x02), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n89_), .B(men_men_n34_), .Y(men_men_n103_));
  NA3        u081(.A(men_men_n103_), .B(men_men_n102_), .C(x06), .Y(men_men_n104_));
  NO2        u082(.A(men_men_n104_), .B(men_men_n101_), .Y(men_men_n105_));
  NO2        u083(.A(men_men_n74_), .B(x13), .Y(men_men_n106_));
  NA2        u084(.A(x09), .B(men_men_n33_), .Y(men_men_n107_));
  NO2        u085(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NA2        u086(.A(x13), .B(men_men_n33_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(x05), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n110_), .B(men_men_n108_), .Y(men_men_n111_));
  NA2        u089(.A(men_men_n33_), .B(men_men_n53_), .Y(men_men_n112_));
  NA2        u090(.A(men_men_n112_), .B(men_men_n89_), .Y(men_men_n113_));
  AOI210     u091(.A0(men_men_n113_), .A1(men_men_n70_), .B0(men_men_n101_), .Y(men_men_n114_));
  AOI210     u092(.A0(men_men_n114_), .A1(men_men_n111_), .B0(men_men_n64_), .Y(men_men_n115_));
  NA2        u093(.A(men_men_n27_), .B(men_men_n45_), .Y(men_men_n116_));
  NA2        u094(.A(x10), .B(men_men_n53_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NA2        u096(.A(men_men_n48_), .B(x05), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n34_), .B(x04), .Y(men_men_n120_));
  NA3        u098(.A(men_men_n120_), .B(men_men_n119_), .C(x13), .Y(men_men_n121_));
  NO3        u099(.A(men_men_n112_), .B(men_men_n69_), .C(men_men_n34_), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n56_), .B(x05), .Y(men_men_n123_));
  NOi41      u101(.An(men_men_n121_), .B(men_men_n123_), .C(men_men_n122_), .D(men_men_n118_), .Y(men_men_n124_));
  NO3        u102(.A(men_men_n124_), .B(x06), .C(x03), .Y(men_men_n125_));
  NO4        u103(.A(men_men_n125_), .B(men_men_n115_), .C(men_men_n105_), .D(men_men_n99_), .Y(men_men_n126_));
  NA2        u104(.A(x13), .B(men_men_n34_), .Y(men_men_n127_));
  OAI210     u105(.A0(men_men_n74_), .A1(x13), .B0(men_men_n33_), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n129_));
  NO2        u107(.A(men_men_n48_), .B(men_men_n39_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n27_), .B(x06), .Y(men_men_n131_));
  OA210      u109(.A0(men_men_n26_), .A1(x04), .B0(men_men_n129_), .Y(men_men_n132_));
  NO2        u110(.A(x09), .B(x05), .Y(men_men_n133_));
  NA2        u111(.A(men_men_n133_), .B(men_men_n45_), .Y(men_men_n134_));
  AOI210     u112(.A0(men_men_n134_), .A1(men_men_n95_), .B0(x06), .Y(men_men_n135_));
  NA2        u113(.A(x09), .B(x00), .Y(men_men_n136_));
  NA2        u114(.A(men_men_n100_), .B(men_men_n136_), .Y(men_men_n137_));
  NA2        u115(.A(men_men_n68_), .B(men_men_n48_), .Y(men_men_n138_));
  AOI210     u116(.A0(men_men_n138_), .A1(men_men_n137_), .B0(men_men_n131_), .Y(men_men_n139_));
  NO3        u117(.A(men_men_n139_), .B(men_men_n135_), .C(men_men_n132_), .Y(men_men_n140_));
  NO2        u118(.A(x03), .B(x02), .Y(men_men_n141_));
  NA2        u119(.A(men_men_n75_), .B(men_men_n89_), .Y(men_men_n142_));
  OAI210     u120(.A0(men_men_n142_), .A1(men_men_n101_), .B0(men_men_n141_), .Y(men_men_n143_));
  OA210      u121(.A0(men_men_n140_), .A1(x11), .B0(men_men_n143_), .Y(men_men_n144_));
  OAI210     u122(.A0(men_men_n126_), .A1(men_men_n23_), .B0(men_men_n144_), .Y(men_men_n145_));
  NA2        u123(.A(men_men_n95_), .B(men_men_n38_), .Y(men_men_n146_));
  NAi21      u124(.An(x06), .B(x10), .Y(men_men_n147_));
  NOi21      u125(.An(x01), .B(x13), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n148_), .B(men_men_n147_), .Y(men_men_n149_));
  OR2        u127(.A(men_men_n149_), .B(x08), .Y(men_men_n150_));
  AOI210     u128(.A0(men_men_n150_), .A1(men_men_n146_), .B0(men_men_n39_), .Y(men_men_n151_));
  NO2        u129(.A(men_men_n27_), .B(x03), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n89_), .B(x01), .Y(men_men_n153_));
  NO2        u131(.A(men_men_n152_), .B(men_men_n46_), .Y(men_men_n154_));
  AOI210     u132(.A0(x11), .A1(men_men_n29_), .B0(men_men_n26_), .Y(men_men_n155_));
  OAI210     u133(.A0(men_men_n154_), .A1(men_men_n151_), .B0(men_men_n155_), .Y(men_men_n156_));
  NA2        u134(.A(x04), .B(x02), .Y(men_men_n157_));
  NA2        u135(.A(x10), .B(x05), .Y(men_men_n158_));
  NA2        u136(.A(x09), .B(x06), .Y(men_men_n159_));
  NO2        u137(.A(x09), .B(x01), .Y(men_men_n160_));
  NO3        u138(.A(men_men_n160_), .B(men_men_n93_), .C(men_men_n29_), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n161_), .B(x00), .Y(men_men_n162_));
  NA3        u140(.A(men_men_n148_), .B(men_men_n147_), .C(men_men_n48_), .Y(men_men_n163_));
  OAI210     u141(.A0(men_men_n418_), .A1(men_men_n103_), .B0(men_men_n163_), .Y(men_men_n164_));
  INV        u142(.A(men_men_n164_), .Y(men_men_n165_));
  OAI210     u143(.A0(men_men_n165_), .A1(x11), .B0(men_men_n162_), .Y(men_men_n166_));
  NAi21      u144(.An(men_men_n157_), .B(men_men_n166_), .Y(men_men_n167_));
  INV        u145(.A(men_men_n25_), .Y(men_men_n168_));
  NAi21      u146(.An(x13), .B(x00), .Y(men_men_n169_));
  AOI210     u147(.A0(men_men_n27_), .A1(men_men_n46_), .B0(men_men_n169_), .Y(men_men_n170_));
  AOI220     u148(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n171_));
  OAI210     u149(.A0(men_men_n158_), .A1(men_men_n33_), .B0(men_men_n171_), .Y(men_men_n172_));
  AN2        u150(.A(men_men_n172_), .B(men_men_n170_), .Y(men_men_n173_));
  NO2        u151(.A(men_men_n85_), .B(x06), .Y(men_men_n174_));
  NO2        u152(.A(men_men_n169_), .B(men_men_n34_), .Y(men_men_n175_));
  OAI220     u153(.A0(men_men_n169_), .A1(men_men_n159_), .B0(men_men_n174_), .B1(men_men_n63_), .Y(men_men_n176_));
  OAI210     u154(.A0(men_men_n176_), .A1(men_men_n173_), .B0(men_men_n168_), .Y(men_men_n177_));
  NOi21      u155(.An(x09), .B(x00), .Y(men_men_n178_));
  NO3        u156(.A(men_men_n73_), .B(men_men_n178_), .C(men_men_n45_), .Y(men_men_n179_));
  INV        u157(.A(men_men_n179_), .Y(men_men_n180_));
  NA2        u158(.A(x10), .B(x08), .Y(men_men_n181_));
  INV        u159(.A(men_men_n181_), .Y(men_men_n182_));
  NA2        u160(.A(x06), .B(x05), .Y(men_men_n183_));
  OAI210     u161(.A0(men_men_n183_), .A1(men_men_n33_), .B0(men_men_n88_), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n182_), .A1(men_men_n54_), .B0(men_men_n184_), .Y(men_men_n185_));
  NA2        u163(.A(men_men_n185_), .B(men_men_n180_), .Y(men_men_n186_));
  AOI210     u164(.A0(men_men_n25_), .A1(men_men_n24_), .B0(x13), .Y(men_men_n187_));
  NA2        u165(.A(men_men_n84_), .B(men_men_n48_), .Y(men_men_n188_));
  NO2        u166(.A(men_men_n33_), .B(men_men_n29_), .Y(men_men_n189_));
  NA2        u167(.A(men_men_n189_), .B(x02), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n190_), .B(men_men_n188_), .Y(men_men_n191_));
  AOI210     u169(.A0(men_men_n187_), .A1(men_men_n186_), .B0(men_men_n191_), .Y(men_men_n192_));
  NA4        u170(.A(men_men_n192_), .B(men_men_n177_), .C(men_men_n167_), .D(men_men_n156_), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n145_), .A1(men_men_n88_), .B0(men_men_n193_), .Y(men_men_n194_));
  AOI210     u172(.A0(men_men_n127_), .A1(x09), .B0(men_men_n65_), .Y(men_men_n195_));
  NA2        u173(.A(men_men_n195_), .B(men_men_n129_), .Y(men_men_n196_));
  NA2        u174(.A(men_men_n48_), .B(men_men_n45_), .Y(men_men_n197_));
  NA2        u175(.A(men_men_n197_), .B(men_men_n128_), .Y(men_men_n198_));
  AOI210     u176(.A0(men_men_n28_), .A1(x06), .B0(x05), .Y(men_men_n199_));
  NO2        u177(.A(men_men_n116_), .B(x06), .Y(men_men_n200_));
  AOI210     u178(.A0(men_men_n199_), .A1(men_men_n198_), .B0(men_men_n200_), .Y(men_men_n201_));
  AOI210     u179(.A0(men_men_n201_), .A1(men_men_n196_), .B0(x12), .Y(men_men_n202_));
  INV        u180(.A(men_men_n68_), .Y(men_men_n203_));
  AOI210     u181(.A0(men_men_n181_), .A1(x05), .B0(men_men_n48_), .Y(men_men_n204_));
  OAI210     u182(.A0(men_men_n204_), .A1(men_men_n149_), .B0(men_men_n53_), .Y(men_men_n205_));
  NA2        u183(.A(men_men_n205_), .B(men_men_n203_), .Y(men_men_n206_));
  NO2        u184(.A(men_men_n84_), .B(x06), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n34_), .A1(x04), .B0(men_men_n48_), .Y(men_men_n208_));
  NO3        u186(.A(men_men_n208_), .B(men_men_n207_), .C(men_men_n39_), .Y(men_men_n209_));
  NA4        u187(.A(men_men_n147_), .B(men_men_n52_), .C(men_men_n34_), .D(x04), .Y(men_men_n210_));
  NA2        u188(.A(men_men_n210_), .B(men_men_n131_), .Y(men_men_n211_));
  OAI210     u189(.A0(men_men_n211_), .A1(men_men_n209_), .B0(x02), .Y(men_men_n212_));
  AOI210     u190(.A0(men_men_n212_), .A1(men_men_n206_), .B0(men_men_n23_), .Y(men_men_n213_));
  OAI210     u191(.A0(men_men_n202_), .A1(men_men_n53_), .B0(men_men_n213_), .Y(men_men_n214_));
  INV        u192(.A(men_men_n131_), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n48_), .B(x03), .Y(men_men_n216_));
  OAI210     u194(.A0(men_men_n69_), .A1(men_men_n34_), .B0(men_men_n107_), .Y(men_men_n217_));
  NO2        u195(.A(men_men_n89_), .B(x03), .Y(men_men_n218_));
  AOI220     u196(.A0(men_men_n218_), .A1(men_men_n217_), .B0(men_men_n68_), .B1(men_men_n216_), .Y(men_men_n219_));
  INV        u197(.A(men_men_n147_), .Y(men_men_n220_));
  NOi21      u198(.An(x13), .B(x04), .Y(men_men_n221_));
  NO3        u199(.A(men_men_n221_), .B(men_men_n68_), .C(men_men_n178_), .Y(men_men_n222_));
  NO2        u200(.A(men_men_n222_), .B(x05), .Y(men_men_n223_));
  AOI210     u201(.A0(men_men_n220_), .A1(men_men_n53_), .B0(men_men_n223_), .Y(men_men_n224_));
  NA2        u202(.A(men_men_n219_), .B(men_men_n224_), .Y(men_men_n225_));
  INV        u203(.A(men_men_n81_), .Y(men_men_n226_));
  NO2        u204(.A(men_men_n226_), .B(x12), .Y(men_men_n227_));
  NA2        u205(.A(men_men_n23_), .B(men_men_n45_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n48_), .B(men_men_n34_), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n229_), .A1(men_men_n172_), .B0(men_men_n170_), .Y(men_men_n230_));
  AOI210     u208(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n231_));
  NO2        u209(.A(x06), .B(x00), .Y(men_men_n232_));
  NO3        u210(.A(men_men_n232_), .B(men_men_n231_), .C(men_men_n39_), .Y(men_men_n233_));
  OAI210     u211(.A0(men_men_n90_), .A1(men_men_n136_), .B0(men_men_n64_), .Y(men_men_n234_));
  NO2        u212(.A(men_men_n234_), .B(men_men_n233_), .Y(men_men_n235_));
  INV        u213(.A(x03), .Y(men_men_n236_));
  OA210      u214(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n230_), .Y(men_men_n237_));
  NA2        u215(.A(x13), .B(men_men_n88_), .Y(men_men_n238_));
  NA3        u216(.A(men_men_n238_), .B(men_men_n184_), .C(men_men_n82_), .Y(men_men_n239_));
  OAI210     u217(.A0(men_men_n237_), .A1(men_men_n228_), .B0(men_men_n239_), .Y(men_men_n240_));
  AOI210     u218(.A0(men_men_n227_), .A1(men_men_n225_), .B0(men_men_n240_), .Y(men_men_n241_));
  AOI210     u219(.A0(men_men_n241_), .A1(men_men_n214_), .B0(x07), .Y(men_men_n242_));
  NA2        u220(.A(men_men_n63_), .B(men_men_n27_), .Y(men_men_n243_));
  AOI210     u221(.A0(men_men_n417_), .A1(men_men_n138_), .B0(men_men_n243_), .Y(men_men_n244_));
  NO2        u222(.A(men_men_n89_), .B(x06), .Y(men_men_n245_));
  NO2        u223(.A(x08), .B(x05), .Y(men_men_n246_));
  NO2        u224(.A(men_men_n246_), .B(men_men_n231_), .Y(men_men_n247_));
  OAI210     u225(.A0(men_men_n68_), .A1(x13), .B0(men_men_n29_), .Y(men_men_n248_));
  OAI210     u226(.A0(men_men_n247_), .A1(men_men_n89_), .B0(men_men_n248_), .Y(men_men_n249_));
  NO2        u227(.A(x12), .B(x02), .Y(men_men_n250_));
  INV        u228(.A(men_men_n250_), .Y(men_men_n251_));
  NO2        u229(.A(men_men_n251_), .B(men_men_n226_), .Y(men_men_n252_));
  OA210      u230(.A0(men_men_n249_), .A1(men_men_n244_), .B0(men_men_n252_), .Y(men_men_n253_));
  NA2        u231(.A(men_men_n48_), .B(men_men_n39_), .Y(men_men_n254_));
  NO2        u232(.A(men_men_n254_), .B(x01), .Y(men_men_n255_));
  NOi21      u233(.An(men_men_n74_), .B(men_men_n107_), .Y(men_men_n256_));
  NO2        u234(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  AOI210     u235(.A0(men_men_n257_), .A1(men_men_n121_), .B0(men_men_n27_), .Y(men_men_n258_));
  NA2        u236(.A(men_men_n245_), .B(men_men_n217_), .Y(men_men_n259_));
  NA2        u237(.A(men_men_n89_), .B(x04), .Y(men_men_n260_));
  NA2        u238(.A(men_men_n260_), .B(men_men_n26_), .Y(men_men_n261_));
  OAI210     u239(.A0(men_men_n261_), .A1(men_men_n106_), .B0(men_men_n259_), .Y(men_men_n262_));
  NO3        u240(.A(men_men_n80_), .B(x12), .C(x03), .Y(men_men_n263_));
  OAI210     u241(.A0(men_men_n262_), .A1(men_men_n258_), .B0(men_men_n263_), .Y(men_men_n264_));
  AOI210     u242(.A0(men_men_n188_), .A1(men_men_n183_), .B0(men_men_n90_), .Y(men_men_n265_));
  NOi21      u243(.An(men_men_n243_), .B(men_men_n207_), .Y(men_men_n266_));
  NO2        u244(.A(men_men_n25_), .B(x00), .Y(men_men_n267_));
  OAI210     u245(.A0(men_men_n266_), .A1(men_men_n265_), .B0(men_men_n267_), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n54_), .B(x05), .Y(men_men_n269_));
  NO3        u247(.A(men_men_n269_), .B(men_men_n208_), .C(men_men_n174_), .Y(men_men_n270_));
  NO2        u248(.A(men_men_n228_), .B(men_men_n26_), .Y(men_men_n271_));
  NA2        u249(.A(men_men_n270_), .B(men_men_n271_), .Y(men_men_n272_));
  NA3        u250(.A(men_men_n272_), .B(men_men_n268_), .C(men_men_n264_), .Y(men_men_n273_));
  NO3        u251(.A(men_men_n273_), .B(men_men_n253_), .C(men_men_n242_), .Y(men_men_n274_));
  OAI210     u252(.A0(men_men_n194_), .A1(men_men_n57_), .B0(men_men_n274_), .Y(men02));
  AOI210     u253(.A0(men_men_n127_), .A1(men_men_n75_), .B0(men_men_n119_), .Y(men_men_n276_));
  NOi21      u254(.An(men_men_n222_), .B(men_men_n160_), .Y(men_men_n277_));
  NA3        u255(.A(x13), .B(men_men_n182_), .C(men_men_n52_), .Y(men_men_n278_));
  OAI210     u256(.A0(men_men_n277_), .A1(men_men_n30_), .B0(men_men_n278_), .Y(men_men_n279_));
  OAI210     u257(.A0(men_men_n279_), .A1(men_men_n276_), .B0(men_men_n158_), .Y(men_men_n280_));
  INV        u258(.A(men_men_n158_), .Y(men_men_n281_));
  NO2        u259(.A(men_men_n102_), .B(men_men_n208_), .Y(men_men_n282_));
  OAI220     u260(.A0(men_men_n282_), .A1(men_men_n89_), .B0(men_men_n75_), .B1(men_men_n48_), .Y(men_men_n283_));
  AOI220     u261(.A0(men_men_n283_), .A1(men_men_n281_), .B0(men_men_n142_), .B1(men_men_n141_), .Y(men_men_n284_));
  AOI210     u262(.A0(men_men_n284_), .A1(men_men_n280_), .B0(men_men_n46_), .Y(men_men_n285_));
  NO2        u263(.A(x05), .B(x02), .Y(men_men_n286_));
  OAI210     u264(.A0(men_men_n198_), .A1(men_men_n178_), .B0(men_men_n286_), .Y(men_men_n287_));
  AOI220     u265(.A0(men_men_n246_), .A1(men_men_n54_), .B0(men_men_n52_), .B1(men_men_n34_), .Y(men_men_n288_));
  NOi21      u266(.An(x13), .B(men_men_n288_), .Y(men_men_n289_));
  AOI210     u267(.A0(men_men_n221_), .A1(men_men_n69_), .B0(men_men_n289_), .Y(men_men_n290_));
  AOI210     u268(.A0(men_men_n290_), .A1(men_men_n287_), .B0(men_men_n131_), .Y(men_men_n291_));
  NAi21      u269(.An(men_men_n223_), .B(men_men_n219_), .Y(men_men_n292_));
  NO2        u270(.A(x06), .B(men_men_n45_), .Y(men_men_n293_));
  NA2        u271(.A(men_men_n293_), .B(men_men_n292_), .Y(men_men_n294_));
  AN2        u272(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n295_));
  OAI210     u273(.A0(men_men_n40_), .A1(men_men_n39_), .B0(men_men_n46_), .Y(men_men_n296_));
  NA2        u274(.A(x13), .B(men_men_n26_), .Y(men_men_n297_));
  AOI210     u275(.A0(men_men_n297_), .A1(men_men_n128_), .B0(men_men_n296_), .Y(men_men_n298_));
  OAI210     u276(.A0(men_men_n298_), .A1(men_men_n295_), .B0(men_men_n85_), .Y(men_men_n299_));
  NA3        u277(.A(men_men_n85_), .B(men_men_n74_), .C(men_men_n216_), .Y(men_men_n300_));
  NA3        u278(.A(men_men_n84_), .B(men_men_n73_), .C(men_men_n40_), .Y(men_men_n301_));
  AOI210     u279(.A0(men_men_n301_), .A1(men_men_n300_), .B0(x04), .Y(men_men_n302_));
  NO2        u280(.A(men_men_n247_), .B(men_men_n91_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n303_), .A1(x13), .B0(men_men_n302_), .Y(men_men_n304_));
  NA3        u282(.A(men_men_n304_), .B(men_men_n299_), .C(men_men_n294_), .Y(men_men_n305_));
  NO3        u283(.A(men_men_n305_), .B(men_men_n291_), .C(men_men_n285_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n130_), .B(x03), .Y(men_men_n307_));
  INV        u285(.A(men_men_n169_), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n48_), .A1(men_men_n33_), .B0(men_men_n34_), .Y(men_men_n309_));
  AOI220     u287(.A0(men_men_n309_), .A1(men_men_n308_), .B0(men_men_n189_), .B1(x08), .Y(men_men_n310_));
  OAI210     u288(.A0(men_men_n310_), .A1(men_men_n269_), .B0(men_men_n307_), .Y(men_men_n311_));
  NA2        u289(.A(men_men_n311_), .B(men_men_n93_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n52_), .A1(x05), .B0(men_men_n94_), .Y(men_men_n313_));
  NA2        u291(.A(men_men_n260_), .B(men_men_n88_), .Y(men_men_n314_));
  NA2        u292(.A(men_men_n88_), .B(men_men_n39_), .Y(men_men_n315_));
  NA3        u293(.A(men_men_n313_), .B(men_men_n312_), .C(men_men_n46_), .Y(men_men_n316_));
  NO3        u294(.A(men_men_n171_), .B(x13), .C(men_men_n29_), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n317_), .A1(men_men_n229_), .B0(men_men_n85_), .Y(men_men_n318_));
  NO3        u296(.A(x13), .B(men_men_n152_), .C(men_men_n49_), .Y(men_men_n319_));
  OAI210     u297(.A0(men_men_n136_), .A1(men_men_n34_), .B0(men_men_n88_), .Y(men_men_n320_));
  NA2        u298(.A(men_men_n320_), .B(men_men_n319_), .Y(men_men_n321_));
  NA3        u299(.A(men_men_n321_), .B(men_men_n318_), .C(x06), .Y(men_men_n322_));
  OAI220     u300(.A0(men_men_n153_), .A1(x09), .B0(x08), .B1(men_men_n39_), .Y(men_men_n323_));
  NO3        u301(.A(men_men_n269_), .B(men_men_n116_), .C(x08), .Y(men_men_n324_));
  AOI210     u302(.A0(men_men_n323_), .A1(men_men_n215_), .B0(men_men_n324_), .Y(men_men_n325_));
  NO2        u303(.A(men_men_n46_), .B(men_men_n39_), .Y(men_men_n326_));
  NO3        u304(.A(men_men_n100_), .B(men_men_n117_), .C(men_men_n36_), .Y(men_men_n327_));
  AOI210     u305(.A0(men_men_n319_), .A1(men_men_n326_), .B0(men_men_n327_), .Y(men_men_n328_));
  OAI210     u306(.A0(men_men_n325_), .A1(men_men_n26_), .B0(men_men_n328_), .Y(men_men_n329_));
  AN2        u307(.A(men_men_n329_), .B(x04), .Y(men_men_n330_));
  AOI210     u308(.A0(men_men_n322_), .A1(men_men_n316_), .B0(men_men_n330_), .Y(men_men_n331_));
  OAI210     u309(.A0(men_men_n306_), .A1(x12), .B0(men_men_n331_), .Y(men03));
  OR2        u310(.A(men_men_n40_), .B(men_men_n216_), .Y(men_men_n333_));
  AOI210     u311(.A0(men_men_n142_), .A1(men_men_n88_), .B0(men_men_n333_), .Y(men_men_n334_));
  NA2        u312(.A(men_men_n334_), .B(x05), .Y(men_men_n335_));
  NA2        u313(.A(men_men_n333_), .B(x05), .Y(men_men_n336_));
  AOI210     u314(.A0(men_men_n128_), .A1(men_men_n203_), .B0(men_men_n336_), .Y(men_men_n337_));
  AOI210     u315(.A0(men_men_n218_), .A1(men_men_n70_), .B0(men_men_n110_), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n55_), .B0(men_men_n297_), .B1(men_men_n288_), .Y(men_men_n339_));
  OAI210     u317(.A0(men_men_n339_), .A1(men_men_n337_), .B0(men_men_n88_), .Y(men_men_n340_));
  AOI210     u318(.A0(men_men_n134_), .A1(men_men_n56_), .B0(men_men_n36_), .Y(men_men_n341_));
  NO2        u319(.A(men_men_n160_), .B(men_men_n123_), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n35_), .Y(men_men_n343_));
  OAI210     u321(.A0(men_men_n343_), .A1(men_men_n341_), .B0(x04), .Y(men_men_n344_));
  AOI210     u322(.A0(men_men_n169_), .A1(men_men_n88_), .B0(men_men_n134_), .Y(men_men_n345_));
  NA4        u323(.A(men_men_n420_), .B(men_men_n344_), .C(men_men_n340_), .D(men_men_n335_), .Y(men04));
  NO2        u324(.A(men_men_n78_), .B(men_men_n37_), .Y(men_men_n347_));
  XO2        u325(.A(men_men_n347_), .B(men_men_n238_), .Y(men05));
  AOI210     u326(.A0(men_men_n63_), .A1(men_men_n49_), .B0(men_men_n200_), .Y(men_men_n349_));
  AOI210     u327(.A0(men_men_n349_), .A1(men_men_n296_), .B0(men_men_n25_), .Y(men_men_n350_));
  NA3        u328(.A(men_men_n131_), .B(men_men_n119_), .C(men_men_n29_), .Y(men_men_n351_));
  AOI210     u329(.A0(men_men_n220_), .A1(men_men_n53_), .B0(men_men_n79_), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n352_), .A1(men_men_n351_), .B0(men_men_n24_), .Y(men_men_n353_));
  OAI210     u331(.A0(men_men_n353_), .A1(men_men_n350_), .B0(men_men_n88_), .Y(men_men_n354_));
  NA2        u332(.A(x11), .B(men_men_n29_), .Y(men_men_n355_));
  NA2        u333(.A(men_men_n23_), .B(men_men_n26_), .Y(men_men_n356_));
  NA2        u334(.A(men_men_n243_), .B(x03), .Y(men_men_n357_));
  OAI220     u335(.A0(men_men_n357_), .A1(men_men_n356_), .B0(men_men_n355_), .B1(men_men_n71_), .Y(men_men_n358_));
  INV        u336(.A(x07), .Y(men_men_n359_));
  AOI210     u337(.A0(men_men_n358_), .A1(x06), .B0(men_men_n359_), .Y(men_men_n360_));
  AOI220     u338(.A0(men_men_n71_), .A1(men_men_n29_), .B0(men_men_n49_), .B1(men_men_n48_), .Y(men_men_n361_));
  NO3        u339(.A(men_men_n361_), .B(men_men_n23_), .C(x00), .Y(men_men_n362_));
  NA2        u340(.A(men_men_n62_), .B(x02), .Y(men_men_n363_));
  AOI210     u341(.A0(men_men_n363_), .A1(men_men_n357_), .B0(men_men_n245_), .Y(men_men_n364_));
  OR2        u342(.A(men_men_n364_), .B(men_men_n228_), .Y(men_men_n365_));
  NA2        u343(.A(men_men_n148_), .B(x05), .Y(men_men_n366_));
  NA3        u344(.A(men_men_n366_), .B(men_men_n232_), .C(men_men_n226_), .Y(men_men_n367_));
  NO2        u345(.A(men_men_n23_), .B(x10), .Y(men_men_n368_));
  OAI210     u346(.A0(x11), .A1(men_men_n27_), .B0(men_men_n46_), .Y(men_men_n369_));
  OR3        u347(.A(men_men_n369_), .B(men_men_n368_), .C(men_men_n42_), .Y(men_men_n370_));
  NA3        u348(.A(men_men_n370_), .B(men_men_n367_), .C(men_men_n365_), .Y(men_men_n371_));
  OAI210     u349(.A0(men_men_n371_), .A1(men_men_n362_), .B0(men_men_n88_), .Y(men_men_n372_));
  INV        u350(.A(x07), .Y(men_men_n373_));
  AOI220     u351(.A0(men_men_n373_), .A1(men_men_n372_), .B0(men_men_n360_), .B1(men_men_n354_), .Y(men_men_n374_));
  NA3        u352(.A(men_men_n23_), .B(men_men_n57_), .C(men_men_n46_), .Y(men_men_n375_));
  AO210      u353(.A0(men_men_n375_), .A1(men_men_n254_), .B0(men_men_n251_), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n368_), .A1(men_men_n66_), .B0(men_men_n130_), .Y(men_men_n377_));
  OR2        u355(.A(men_men_n377_), .B(x03), .Y(men_men_n378_));
  NA2        u356(.A(men_men_n326_), .B(men_men_n57_), .Y(men_men_n379_));
  NO2        u357(.A(men_men_n379_), .B(x11), .Y(men_men_n380_));
  NO3        u358(.A(men_men_n380_), .B(men_men_n133_), .C(men_men_n26_), .Y(men_men_n381_));
  AOI220     u359(.A0(men_men_n381_), .A1(men_men_n378_), .B0(men_men_n376_), .B1(men_men_n45_), .Y(men_men_n382_));
  NO4        u360(.A(men_men_n315_), .B(men_men_n30_), .C(x11), .D(x09), .Y(men_men_n383_));
  OAI210     u361(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n89_), .Y(men_men_n384_));
  NOi21      u362(.An(men_men_n307_), .B(men_men_n123_), .Y(men_men_n385_));
  AOI210     u363(.A0(men_men_n368_), .A1(men_men_n26_), .B0(men_men_n29_), .Y(men_men_n386_));
  NA2        u364(.A(x09), .B(men_men_n39_), .Y(men_men_n387_));
  OAI220     u365(.A0(men_men_n387_), .A1(men_men_n386_), .B0(men_men_n355_), .B1(men_men_n58_), .Y(men_men_n388_));
  NO2        u366(.A(x13), .B(x12), .Y(men_men_n389_));
  NO2        u367(.A(men_men_n119_), .B(men_men_n26_), .Y(men_men_n390_));
  NO2        u368(.A(men_men_n390_), .B(men_men_n255_), .Y(men_men_n391_));
  OR3        u369(.A(men_men_n391_), .B(x12), .C(x03), .Y(men_men_n392_));
  NA2        u370(.A(men_men_n392_), .B(x08), .Y(men_men_n393_));
  AOI210     u371(.A0(men_men_n389_), .A1(men_men_n388_), .B0(men_men_n393_), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n419_), .A1(men_men_n384_), .B0(men_men_n394_), .Y(men_men_n395_));
  OAI210     u373(.A0(men_men_n379_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n396_));
  NA2        u374(.A(men_men_n281_), .B(x07), .Y(men_men_n397_));
  OAI220     u375(.A0(men_men_n397_), .A1(men_men_n356_), .B0(men_men_n133_), .B1(men_men_n41_), .Y(men_men_n398_));
  OAI210     u376(.A0(men_men_n398_), .A1(men_men_n396_), .B0(men_men_n175_), .Y(men_men_n399_));
  NA3        u377(.A(men_men_n391_), .B(men_men_n385_), .C(men_men_n314_), .Y(men_men_n400_));
  INV        u378(.A(x14), .Y(men_men_n401_));
  NO3        u379(.A(men_men_n307_), .B(men_men_n91_), .C(x11), .Y(men_men_n402_));
  NO3        u380(.A(men_men_n153_), .B(men_men_n66_), .C(men_men_n53_), .Y(men_men_n403_));
  NO3        u381(.A(men_men_n375_), .B(men_men_n315_), .C(men_men_n169_), .Y(men_men_n404_));
  NO4        u382(.A(men_men_n404_), .B(men_men_n403_), .C(men_men_n402_), .D(men_men_n401_), .Y(men_men_n405_));
  NA3        u383(.A(men_men_n405_), .B(men_men_n400_), .C(men_men_n399_), .Y(men_men_n406_));
  NA2        u384(.A(men_men_n390_), .B(men_men_n152_), .Y(men_men_n407_));
  NOi21      u385(.An(men_men_n260_), .B(men_men_n137_), .Y(men_men_n408_));
  NO3        u386(.A(men_men_n116_), .B(men_men_n24_), .C(x06), .Y(men_men_n409_));
  AOI210     u387(.A0(men_men_n267_), .A1(men_men_n220_), .B0(men_men_n409_), .Y(men_men_n410_));
  INV        u388(.A(men_men_n410_), .Y(men_men_n411_));
  OAI210     u389(.A0(men_men_n411_), .A1(men_men_n408_), .B0(men_men_n88_), .Y(men_men_n412_));
  OAI210     u390(.A0(men_men_n407_), .A1(men_men_n80_), .B0(men_men_n412_), .Y(men_men_n413_));
  NO4        u391(.A(men_men_n413_), .B(men_men_n406_), .C(men_men_n395_), .D(men_men_n374_), .Y(men06));
  INV        u392(.A(men_men_n178_), .Y(men_men_n417_));
  INV        u393(.A(x05), .Y(men_men_n418_));
  INV        u394(.A(x08), .Y(men_men_n419_));
  INV        u395(.A(men_men_n345_), .Y(men_men_n420_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule