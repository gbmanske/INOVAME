library verilog;
use verilog.vl_types.all;
entity fulladder_vlg_vec_tst is
end fulladder_vlg_vec_tst;
