//Benchmark atmr_intb_466_0.0313

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n331_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n374_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n381_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  INV        o035(.A(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(ori_ori_n24_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n60_), .B(ori_ori_n58_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n62_));
  OAI210     o040(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o041(.A0(ori_ori_n63_), .A1(ori_ori_n55_), .B0(ori_ori_n61_), .B1(ori_ori_n31_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(x05), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n57_), .B(ori_ori_n23_), .Y(ori_ori_n66_));
  NA2        o044(.A(x09), .B(x05), .Y(ori_ori_n67_));
  NA2        o045(.A(x10), .B(x06), .Y(ori_ori_n68_));
  NA3        o046(.A(ori_ori_n68_), .B(ori_ori_n67_), .C(ori_ori_n28_), .Y(ori_ori_n69_));
  NO2        o047(.A(ori_ori_n57_), .B(ori_ori_n41_), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n69_), .A1(ori_ori_n66_), .B0(x03), .Y(ori_ori_n71_));
  NOi31      o049(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n72_));
  INV        o050(.A(x07), .Y(ori_ori_n73_));
  NO2        o051(.A(ori_ori_n73_), .B(ori_ori_n24_), .Y(ori_ori_n74_));
  NO2        o052(.A(x09), .B(ori_ori_n41_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n36_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n75_), .A1(ori_ori_n29_), .B0(x02), .Y(ori_ori_n77_));
  AOI210     o055(.A0(ori_ori_n76_), .A1(ori_ori_n48_), .B0(ori_ori_n77_), .Y(ori_ori_n78_));
  NO2        o056(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n79_));
  NO2        o057(.A(x08), .B(x01), .Y(ori_ori_n80_));
  OAI210     o058(.A0(ori_ori_n80_), .A1(ori_ori_n79_), .B0(ori_ori_n35_), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n82_));
  NO3        o060(.A(ori_ori_n81_), .B(ori_ori_n78_), .C(ori_ori_n74_), .Y(ori_ori_n83_));
  AN2        o061(.A(ori_ori_n83_), .B(ori_ori_n71_), .Y(ori_ori_n84_));
  INV        o062(.A(ori_ori_n81_), .Y(ori_ori_n85_));
  NA2        o063(.A(x11), .B(x00), .Y(ori_ori_n86_));
  NO2        o064(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n87_));
  NOi21      o065(.An(ori_ori_n86_), .B(ori_ori_n87_), .Y(ori_ori_n88_));
  NOi21      o066(.An(x01), .B(x10), .Y(ori_ori_n89_));
  NO2        o067(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n90_));
  NO3        o068(.A(ori_ori_n90_), .B(ori_ori_n89_), .C(x06), .Y(ori_ori_n91_));
  NA2        o069(.A(ori_ori_n91_), .B(ori_ori_n27_), .Y(ori_ori_n92_));
  OAI210     o070(.A0(ori_ori_n381_), .A1(x07), .B0(ori_ori_n92_), .Y(ori_ori_n93_));
  NO3        o071(.A(ori_ori_n93_), .B(ori_ori_n84_), .C(ori_ori_n65_), .Y(ori01));
  INV        o072(.A(x12), .Y(ori_ori_n95_));
  INV        o073(.A(x13), .Y(ori_ori_n96_));
  NA2        o074(.A(ori_ori_n89_), .B(ori_ori_n28_), .Y(ori_ori_n97_));
  NO2        o075(.A(x10), .B(x01), .Y(ori_ori_n98_));
  NO2        o076(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  NA2        o078(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n101_));
  NO2        o079(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n102_));
  NOi21      o080(.An(ori_ori_n102_), .B(ori_ori_n54_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n35_), .B(x02), .Y(ori_ori_n104_));
  NA2        o082(.A(x09), .B(ori_ori_n35_), .Y(ori_ori_n105_));
  NA2        o083(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n106_));
  NO2        o084(.A(ori_ori_n106_), .B(x05), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n108_));
  INV        o086(.A(ori_ori_n103_), .Y(ori_ori_n109_));
  NO2        o087(.A(ori_ori_n109_), .B(ori_ori_n68_), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n111_));
  NA2        o089(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(ori_ori_n111_), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n114_));
  NA2        o092(.A(ori_ori_n36_), .B(x04), .Y(ori_ori_n115_));
  NA3        o093(.A(ori_ori_n115_), .B(ori_ori_n114_), .C(x13), .Y(ori_ori_n116_));
  NO2        o094(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n117_));
  NOi31      o095(.An(ori_ori_n116_), .B(ori_ori_n117_), .C(ori_ori_n113_), .Y(ori_ori_n118_));
  NO3        o096(.A(ori_ori_n118_), .B(x06), .C(x03), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n119_), .B(ori_ori_n110_), .Y(ori_ori_n120_));
  NA2        o098(.A(x13), .B(ori_ori_n36_), .Y(ori_ori_n121_));
  OAI210     o099(.A0(ori_ori_n80_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n122_), .B(ori_ori_n121_), .Y(ori_ori_n123_));
  NO2        o101(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n124_));
  NA2        o102(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n125_));
  AOI210     o103(.A0(ori_ori_n125_), .A1(ori_ori_n49_), .B0(ori_ori_n124_), .Y(ori_ori_n126_));
  AN2        o104(.A(ori_ori_n126_), .B(ori_ori_n123_), .Y(ori_ori_n127_));
  NO2        o105(.A(x09), .B(x05), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n47_), .Y(ori_ori_n129_));
  NO2        o107(.A(ori_ori_n100_), .B(ori_ori_n49_), .Y(ori_ori_n130_));
  NA2        o108(.A(x09), .B(x00), .Y(ori_ori_n131_));
  NA2        o109(.A(ori_ori_n102_), .B(ori_ori_n131_), .Y(ori_ori_n132_));
  NO2        o110(.A(ori_ori_n132_), .B(ori_ori_n125_), .Y(ori_ori_n133_));
  NO3        o111(.A(ori_ori_n133_), .B(ori_ori_n130_), .C(ori_ori_n127_), .Y(ori_ori_n134_));
  NO2        o112(.A(x03), .B(x02), .Y(ori_ori_n135_));
  NA2        o113(.A(ori_ori_n81_), .B(ori_ori_n96_), .Y(ori_ori_n136_));
  OAI210     o114(.A0(ori_ori_n136_), .A1(ori_ori_n103_), .B0(ori_ori_n135_), .Y(ori_ori_n137_));
  OA210      o115(.A0(ori_ori_n134_), .A1(x11), .B0(ori_ori_n137_), .Y(ori_ori_n138_));
  OAI210     o116(.A0(ori_ori_n120_), .A1(ori_ori_n23_), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  NA2        o117(.A(ori_ori_n100_), .B(ori_ori_n40_), .Y(ori_ori_n140_));
  NAi21      o118(.An(x06), .B(x10), .Y(ori_ori_n141_));
  NO2        o119(.A(ori_ori_n140_), .B(ori_ori_n41_), .Y(ori_ori_n142_));
  NO2        o120(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n96_), .B(x01), .Y(ori_ori_n144_));
  NO2        o122(.A(ori_ori_n144_), .B(x08), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n143_), .B(ori_ori_n48_), .Y(ori_ori_n146_));
  AOI210     o124(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n147_));
  OAI210     o125(.A0(ori_ori_n146_), .A1(ori_ori_n142_), .B0(ori_ori_n147_), .Y(ori_ori_n148_));
  NA2        o126(.A(x04), .B(x02), .Y(ori_ori_n149_));
  NA2        o127(.A(x10), .B(x05), .Y(ori_ori_n150_));
  NO2        o128(.A(x09), .B(x01), .Y(ori_ori_n151_));
  NO2        o129(.A(ori_ori_n102_), .B(x08), .Y(ori_ori_n152_));
  INV        o130(.A(ori_ori_n25_), .Y(ori_ori_n153_));
  NAi21      o131(.An(x13), .B(x00), .Y(ori_ori_n154_));
  AN2        o132(.A(ori_ori_n68_), .B(ori_ori_n67_), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n90_), .B(x06), .Y(ori_ori_n156_));
  NO2        o134(.A(ori_ori_n154_), .B(ori_ori_n36_), .Y(ori_ori_n157_));
  INV        o135(.A(ori_ori_n157_), .Y(ori_ori_n158_));
  NO2        o136(.A(ori_ori_n156_), .B(ori_ori_n155_), .Y(ori_ori_n159_));
  NA2        o137(.A(ori_ori_n159_), .B(ori_ori_n153_), .Y(ori_ori_n160_));
  NOi21      o138(.An(x09), .B(x00), .Y(ori_ori_n161_));
  NO3        o139(.A(ori_ori_n79_), .B(ori_ori_n161_), .C(ori_ori_n47_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n162_), .B(ori_ori_n112_), .Y(ori_ori_n163_));
  NA2        o141(.A(x06), .B(x05), .Y(ori_ori_n164_));
  OAI210     o142(.A0(ori_ori_n164_), .A1(ori_ori_n35_), .B0(ori_ori_n95_), .Y(ori_ori_n165_));
  AOI210     o143(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n165_), .Y(ori_ori_n166_));
  NA2        o144(.A(ori_ori_n166_), .B(ori_ori_n163_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n96_), .B(x12), .Y(ori_ori_n168_));
  AOI210     o146(.A0(ori_ori_n25_), .A1(ori_ori_n24_), .B0(ori_ori_n168_), .Y(ori_ori_n169_));
  NO2        o147(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n170_));
  NA2        o148(.A(ori_ori_n170_), .B(x02), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n169_), .B(ori_ori_n167_), .Y(ori_ori_n172_));
  NA3        o150(.A(ori_ori_n172_), .B(ori_ori_n160_), .C(ori_ori_n148_), .Y(ori_ori_n173_));
  AOI210     o151(.A0(ori_ori_n139_), .A1(ori_ori_n95_), .B0(ori_ori_n173_), .Y(ori_ori_n174_));
  INV        o152(.A(ori_ori_n69_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n123_), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n177_));
  NA2        o155(.A(ori_ori_n177_), .B(ori_ori_n122_), .Y(ori_ori_n178_));
  AOI210     o156(.A0(ori_ori_n30_), .A1(x06), .B0(x05), .Y(ori_ori_n179_));
  NO2        o157(.A(ori_ori_n111_), .B(x06), .Y(ori_ori_n180_));
  AOI210     o158(.A0(ori_ori_n179_), .A1(ori_ori_n178_), .B0(ori_ori_n180_), .Y(ori_ori_n181_));
  AOI210     o159(.A0(ori_ori_n181_), .A1(ori_ori_n176_), .B0(x12), .Y(ori_ori_n182_));
  INV        o160(.A(ori_ori_n72_), .Y(ori_ori_n183_));
  NO2        o161(.A(ori_ori_n89_), .B(x06), .Y(ori_ori_n184_));
  AOI210     o162(.A0(ori_ori_n36_), .A1(x04), .B0(ori_ori_n50_), .Y(ori_ori_n185_));
  NO3        o163(.A(ori_ori_n185_), .B(ori_ori_n184_), .C(ori_ori_n41_), .Y(ori_ori_n186_));
  INV        o164(.A(ori_ori_n125_), .Y(ori_ori_n187_));
  OAI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n186_), .B0(x02), .Y(ori_ori_n188_));
  AOI210     o166(.A0(ori_ori_n188_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n189_));
  OAI210     o167(.A0(ori_ori_n182_), .A1(ori_ori_n53_), .B0(ori_ori_n189_), .Y(ori_ori_n190_));
  INV        o168(.A(ori_ori_n125_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n192_));
  OAI210     o170(.A0(ori_ori_n75_), .A1(ori_ori_n36_), .B0(ori_ori_n105_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n96_), .B(x03), .Y(ori_ori_n194_));
  AOI220     o172(.A0(ori_ori_n194_), .A1(ori_ori_n193_), .B0(ori_ori_n72_), .B1(ori_ori_n192_), .Y(ori_ori_n195_));
  NA2        o173(.A(ori_ori_n32_), .B(x06), .Y(ori_ori_n196_));
  INV        o174(.A(ori_ori_n141_), .Y(ori_ori_n197_));
  NOi21      o175(.An(x13), .B(x04), .Y(ori_ori_n198_));
  NO3        o176(.A(ori_ori_n198_), .B(ori_ori_n72_), .C(ori_ori_n161_), .Y(ori_ori_n199_));
  NO2        o177(.A(ori_ori_n199_), .B(x05), .Y(ori_ori_n200_));
  AOI220     o178(.A0(ori_ori_n200_), .A1(ori_ori_n196_), .B0(ori_ori_n197_), .B1(ori_ori_n53_), .Y(ori_ori_n201_));
  OAI210     o179(.A0(ori_ori_n195_), .A1(ori_ori_n191_), .B0(ori_ori_n201_), .Y(ori_ori_n202_));
  INV        o180(.A(ori_ori_n87_), .Y(ori_ori_n203_));
  NO2        o181(.A(ori_ori_n203_), .B(x12), .Y(ori_ori_n204_));
  NA2        o182(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n205_));
  NO2        o183(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n206_));
  AOI210     o184(.A0(x08), .A1(x04), .B0(x09), .Y(ori_ori_n207_));
  NO2        o185(.A(x06), .B(x00), .Y(ori_ori_n208_));
  NO3        o186(.A(ori_ori_n208_), .B(ori_ori_n207_), .C(ori_ori_n41_), .Y(ori_ori_n209_));
  INV        o187(.A(ori_ori_n68_), .Y(ori_ori_n210_));
  NO2        o188(.A(ori_ori_n210_), .B(ori_ori_n209_), .Y(ori_ori_n211_));
  NA2        o189(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n212_));
  NA2        o190(.A(ori_ori_n212_), .B(x03), .Y(ori_ori_n213_));
  OR2        o191(.A(ori_ori_n213_), .B(ori_ori_n211_), .Y(ori_ori_n214_));
  NA2        o192(.A(x13), .B(ori_ori_n95_), .Y(ori_ori_n215_));
  NA3        o193(.A(ori_ori_n215_), .B(ori_ori_n165_), .C(ori_ori_n88_), .Y(ori_ori_n216_));
  OAI210     o194(.A0(ori_ori_n214_), .A1(ori_ori_n205_), .B0(ori_ori_n216_), .Y(ori_ori_n217_));
  AOI210     o195(.A0(ori_ori_n204_), .A1(ori_ori_n202_), .B0(ori_ori_n217_), .Y(ori_ori_n218_));
  AOI210     o196(.A0(ori_ori_n218_), .A1(ori_ori_n190_), .B0(x07), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n67_), .B(ori_ori_n29_), .Y(ori_ori_n220_));
  NOi31      o198(.An(ori_ori_n121_), .B(ori_ori_n198_), .C(ori_ori_n161_), .Y(ori_ori_n221_));
  NO2        o199(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NO2        o200(.A(x08), .B(x05), .Y(ori_ori_n223_));
  NO2        o201(.A(ori_ori_n223_), .B(ori_ori_n207_), .Y(ori_ori_n224_));
  OAI210     o202(.A0(ori_ori_n72_), .A1(x13), .B0(ori_ori_n31_), .Y(ori_ori_n225_));
  INV        o203(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  NO2        o204(.A(x12), .B(x02), .Y(ori_ori_n227_));
  INV        o205(.A(ori_ori_n227_), .Y(ori_ori_n228_));
  NO2        o206(.A(ori_ori_n228_), .B(ori_ori_n203_), .Y(ori_ori_n229_));
  OA210      o207(.A0(ori_ori_n226_), .A1(ori_ori_n222_), .B0(ori_ori_n229_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n231_));
  NO2        o209(.A(ori_ori_n231_), .B(x01), .Y(ori_ori_n232_));
  INV        o210(.A(ori_ori_n232_), .Y(ori_ori_n233_));
  AOI210     o211(.A0(ori_ori_n233_), .A1(ori_ori_n116_), .B0(ori_ori_n29_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n96_), .B(x04), .Y(ori_ori_n235_));
  NA2        o213(.A(ori_ori_n235_), .B(ori_ori_n28_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n383_), .Y(ori_ori_n237_));
  NO3        o215(.A(ori_ori_n86_), .B(x12), .C(x03), .Y(ori_ori_n238_));
  OAI210     o216(.A0(ori_ori_n237_), .A1(ori_ori_n234_), .B0(ori_ori_n238_), .Y(ori_ori_n239_));
  NOi21      o217(.An(ori_ori_n220_), .B(ori_ori_n184_), .Y(ori_ori_n240_));
  NO2        o218(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n241_));
  NA2        o219(.A(ori_ori_n240_), .B(ori_ori_n241_), .Y(ori_ori_n242_));
  NO2        o220(.A(ori_ori_n54_), .B(x05), .Y(ori_ori_n243_));
  NO3        o221(.A(ori_ori_n243_), .B(ori_ori_n185_), .C(ori_ori_n156_), .Y(ori_ori_n244_));
  NO2        o222(.A(ori_ori_n205_), .B(ori_ori_n28_), .Y(ori_ori_n245_));
  OAI210     o223(.A0(ori_ori_n244_), .A1(ori_ori_n191_), .B0(ori_ori_n245_), .Y(ori_ori_n246_));
  NA3        o224(.A(ori_ori_n246_), .B(ori_ori_n242_), .C(ori_ori_n239_), .Y(ori_ori_n247_));
  NO3        o225(.A(ori_ori_n247_), .B(ori_ori_n230_), .C(ori_ori_n219_), .Y(ori_ori_n248_));
  OAI210     o226(.A0(ori_ori_n174_), .A1(ori_ori_n57_), .B0(ori_ori_n248_), .Y(ori02));
  AOI210     o227(.A0(ori_ori_n121_), .A1(ori_ori_n81_), .B0(ori_ori_n114_), .Y(ori_ori_n250_));
  NOi21      o228(.An(ori_ori_n199_), .B(ori_ori_n151_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n251_), .B(ori_ori_n32_), .Y(ori_ori_n252_));
  OAI210     o230(.A0(ori_ori_n252_), .A1(ori_ori_n250_), .B0(ori_ori_n150_), .Y(ori_ori_n253_));
  INV        o231(.A(ori_ori_n150_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n104_), .A1(ori_ori_n82_), .B0(ori_ori_n185_), .Y(ori_ori_n255_));
  OAI220     o233(.A0(ori_ori_n255_), .A1(ori_ori_n96_), .B0(ori_ori_n81_), .B1(ori_ori_n50_), .Y(ori_ori_n256_));
  AOI220     o234(.A0(ori_ori_n256_), .A1(ori_ori_n254_), .B0(ori_ori_n136_), .B1(ori_ori_n135_), .Y(ori_ori_n257_));
  AOI210     o235(.A0(ori_ori_n257_), .A1(ori_ori_n253_), .B0(ori_ori_n48_), .Y(ori_ori_n258_));
  NO2        o236(.A(x05), .B(x02), .Y(ori_ori_n259_));
  OAI210     o237(.A0(ori_ori_n178_), .A1(ori_ori_n161_), .B0(ori_ori_n259_), .Y(ori_ori_n260_));
  AOI220     o238(.A0(ori_ori_n223_), .A1(ori_ori_n54_), .B0(ori_ori_n52_), .B1(ori_ori_n36_), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n260_), .B(ori_ori_n125_), .Y(ori_ori_n262_));
  NAi21      o240(.An(ori_ori_n200_), .B(ori_ori_n195_), .Y(ori_ori_n263_));
  NO2        o241(.A(ori_ori_n212_), .B(ori_ori_n47_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n265_));
  AN2        o243(.A(ori_ori_n194_), .B(ori_ori_n193_), .Y(ori_ori_n266_));
  OAI210     o244(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n267_));
  NA2        o245(.A(x13), .B(ori_ori_n28_), .Y(ori_ori_n268_));
  OA210      o246(.A0(ori_ori_n268_), .A1(x08), .B0(ori_ori_n129_), .Y(ori_ori_n269_));
  AOI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n122_), .B0(ori_ori_n267_), .Y(ori_ori_n270_));
  OAI210     o248(.A0(ori_ori_n270_), .A1(ori_ori_n266_), .B0(ori_ori_n90_), .Y(ori_ori_n271_));
  INV        o249(.A(ori_ori_n135_), .Y(ori_ori_n272_));
  OAI220     o250(.A0(ori_ori_n224_), .A1(ori_ori_n97_), .B0(ori_ori_n272_), .B1(ori_ori_n113_), .Y(ori_ori_n273_));
  NA2        o251(.A(ori_ori_n273_), .B(x13), .Y(ori_ori_n274_));
  NA3        o252(.A(ori_ori_n274_), .B(ori_ori_n271_), .C(ori_ori_n265_), .Y(ori_ori_n275_));
  NO3        o253(.A(ori_ori_n275_), .B(ori_ori_n262_), .C(ori_ori_n258_), .Y(ori_ori_n276_));
  NA2        o254(.A(ori_ori_n124_), .B(x03), .Y(ori_ori_n277_));
  INV        o255(.A(ori_ori_n154_), .Y(ori_ori_n278_));
  AOI220     o256(.A0(x08), .A1(ori_ori_n278_), .B0(ori_ori_n170_), .B1(x08), .Y(ori_ori_n279_));
  OAI210     o257(.A0(ori_ori_n279_), .A1(ori_ori_n243_), .B0(ori_ori_n277_), .Y(ori_ori_n280_));
  NA2        o258(.A(ori_ori_n280_), .B(ori_ori_n98_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n149_), .B(ori_ori_n144_), .Y(ori_ori_n282_));
  AN2        o260(.A(ori_ori_n282_), .B(ori_ori_n152_), .Y(ori_ori_n283_));
  NO2        o261(.A(ori_ori_n114_), .B(ori_ori_n28_), .Y(ori_ori_n284_));
  OAI210     o262(.A0(ori_ori_n284_), .A1(ori_ori_n283_), .B0(ori_ori_n99_), .Y(ori_ori_n285_));
  NA2        o263(.A(ori_ori_n235_), .B(ori_ori_n95_), .Y(ori_ori_n286_));
  NA2        o264(.A(ori_ori_n95_), .B(ori_ori_n41_), .Y(ori_ori_n287_));
  NA3        o265(.A(ori_ori_n287_), .B(ori_ori_n286_), .C(ori_ori_n113_), .Y(ori_ori_n288_));
  NA4        o266(.A(ori_ori_n288_), .B(ori_ori_n285_), .C(ori_ori_n281_), .D(ori_ori_n48_), .Y(ori_ori_n289_));
  INV        o267(.A(ori_ori_n170_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n291_));
  OAI220     o269(.A0(ori_ori_n291_), .A1(ori_ori_n382_), .B0(ori_ori_n290_), .B1(ori_ori_n55_), .Y(ori_ori_n292_));
  NA2        o270(.A(ori_ori_n292_), .B(x02), .Y(ori_ori_n293_));
  INV        o271(.A(ori_ori_n206_), .Y(ori_ori_n294_));
  NA2        o272(.A(ori_ori_n168_), .B(x04), .Y(ori_ori_n295_));
  NO3        o273(.A(ori_ori_n168_), .B(ori_ori_n143_), .C(ori_ori_n51_), .Y(ori_ori_n296_));
  OAI210     o274(.A0(ori_ori_n131_), .A1(ori_ori_n36_), .B0(ori_ori_n95_), .Y(ori_ori_n297_));
  OAI210     o275(.A0(ori_ori_n297_), .A1(ori_ori_n162_), .B0(ori_ori_n296_), .Y(ori_ori_n298_));
  NA3        o276(.A(ori_ori_n298_), .B(ori_ori_n293_), .C(x06), .Y(ori_ori_n299_));
  NA2        o277(.A(x09), .B(x03), .Y(ori_ori_n300_));
  OAI220     o278(.A0(ori_ori_n300_), .A1(ori_ori_n112_), .B0(ori_ori_n177_), .B1(ori_ori_n59_), .Y(ori_ori_n301_));
  NO3        o279(.A(ori_ori_n243_), .B(ori_ori_n111_), .C(x08), .Y(ori_ori_n302_));
  INV        o280(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  NO2        o281(.A(ori_ori_n48_), .B(ori_ori_n41_), .Y(ori_ori_n304_));
  NO3        o282(.A(ori_ori_n102_), .B(ori_ori_n112_), .C(ori_ori_n38_), .Y(ori_ori_n305_));
  AOI210     o283(.A0(ori_ori_n296_), .A1(ori_ori_n304_), .B0(ori_ori_n305_), .Y(ori_ori_n306_));
  OAI210     o284(.A0(ori_ori_n303_), .A1(ori_ori_n28_), .B0(ori_ori_n306_), .Y(ori_ori_n307_));
  AO220      o285(.A0(ori_ori_n307_), .A1(x04), .B0(ori_ori_n301_), .B1(x05), .Y(ori_ori_n308_));
  AOI210     o286(.A0(ori_ori_n299_), .A1(ori_ori_n289_), .B0(ori_ori_n308_), .Y(ori_ori_n309_));
  OAI210     o287(.A0(ori_ori_n276_), .A1(x12), .B0(ori_ori_n309_), .Y(ori03));
  OR2        o288(.A(ori_ori_n42_), .B(ori_ori_n192_), .Y(ori_ori_n311_));
  AOI210     o289(.A0(ori_ori_n136_), .A1(ori_ori_n95_), .B0(ori_ori_n311_), .Y(ori_ori_n312_));
  AO210      o290(.A0(ori_ori_n294_), .A1(ori_ori_n82_), .B0(ori_ori_n295_), .Y(ori_ori_n313_));
  NA2        o291(.A(ori_ori_n168_), .B(ori_ori_n135_), .Y(ori_ori_n314_));
  NA3        o292(.A(ori_ori_n314_), .B(ori_ori_n313_), .C(ori_ori_n171_), .Y(ori_ori_n315_));
  OAI210     o293(.A0(ori_ori_n315_), .A1(ori_ori_n312_), .B0(x05), .Y(ori_ori_n316_));
  NA2        o294(.A(ori_ori_n311_), .B(x05), .Y(ori_ori_n317_));
  AOI210     o295(.A0(ori_ori_n122_), .A1(ori_ori_n183_), .B0(ori_ori_n317_), .Y(ori_ori_n318_));
  AOI210     o296(.A0(ori_ori_n194_), .A1(ori_ori_n76_), .B0(ori_ori_n107_), .Y(ori_ori_n319_));
  OAI220     o297(.A0(ori_ori_n319_), .A1(ori_ori_n55_), .B0(ori_ori_n268_), .B1(ori_ori_n261_), .Y(ori_ori_n320_));
  OAI210     o298(.A0(ori_ori_n320_), .A1(ori_ori_n318_), .B0(ori_ori_n95_), .Y(ori_ori_n321_));
  AOI210     o299(.A0(ori_ori_n129_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n322_));
  NO2        o300(.A(ori_ori_n151_), .B(ori_ori_n117_), .Y(ori_ori_n323_));
  OAI220     o301(.A0(ori_ori_n323_), .A1(ori_ori_n37_), .B0(ori_ori_n132_), .B1(x13), .Y(ori_ori_n324_));
  OAI210     o302(.A0(ori_ori_n324_), .A1(ori_ori_n322_), .B0(x04), .Y(ori_ori_n325_));
  NO3        o303(.A(ori_ori_n287_), .B(ori_ori_n81_), .C(ori_ori_n55_), .Y(ori_ori_n326_));
  AOI210     o304(.A0(ori_ori_n158_), .A1(ori_ori_n95_), .B0(ori_ori_n129_), .Y(ori_ori_n327_));
  OA210      o305(.A0(ori_ori_n145_), .A1(x12), .B0(ori_ori_n117_), .Y(ori_ori_n328_));
  NO3        o306(.A(ori_ori_n328_), .B(ori_ori_n327_), .C(ori_ori_n326_), .Y(ori_ori_n329_));
  NA4        o307(.A(ori_ori_n329_), .B(ori_ori_n325_), .C(ori_ori_n321_), .D(ori_ori_n316_), .Y(ori04));
  NO2        o308(.A(ori_ori_n85_), .B(ori_ori_n39_), .Y(ori_ori_n331_));
  XO2        o309(.A(ori_ori_n331_), .B(ori_ori_n215_), .Y(ori05));
  NO2        o310(.A(ori_ori_n51_), .B(ori_ori_n180_), .Y(ori_ori_n333_));
  AOI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n267_), .B0(ori_ori_n25_), .Y(ori_ori_n334_));
  NO2        o312(.A(x06), .B(ori_ori_n24_), .Y(ori_ori_n335_));
  OAI210     o313(.A0(ori_ori_n335_), .A1(ori_ori_n334_), .B0(ori_ori_n95_), .Y(ori_ori_n336_));
  OAI210     o314(.A0(ori_ori_n26_), .A1(ori_ori_n95_), .B0(x07), .Y(ori_ori_n337_));
  INV        o315(.A(ori_ori_n337_), .Y(ori_ori_n338_));
  AOI210     o316(.A0(ori_ori_n77_), .A1(ori_ori_n31_), .B0(ori_ori_n51_), .Y(ori_ori_n339_));
  NO3        o317(.A(ori_ori_n339_), .B(ori_ori_n23_), .C(x00), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n208_), .B(ori_ori_n203_), .Y(ori_ori_n341_));
  NA2        o319(.A(ori_ori_n341_), .B(ori_ori_n205_), .Y(ori_ori_n342_));
  OAI210     o320(.A0(ori_ori_n342_), .A1(ori_ori_n340_), .B0(ori_ori_n95_), .Y(ori_ori_n343_));
  NA2        o321(.A(ori_ori_n33_), .B(ori_ori_n95_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n344_), .A1(ori_ori_n87_), .B0(x07), .Y(ori_ori_n345_));
  AOI220     o323(.A0(ori_ori_n345_), .A1(ori_ori_n343_), .B0(ori_ori_n338_), .B1(ori_ori_n336_), .Y(ori_ori_n346_));
  OR2        o324(.A(ori_ori_n231_), .B(ori_ori_n228_), .Y(ori_ori_n347_));
  NO2        o325(.A(ori_ori_n128_), .B(ori_ori_n28_), .Y(ori_ori_n348_));
  AOI210     o326(.A0(ori_ori_n347_), .A1(ori_ori_n47_), .B0(ori_ori_n348_), .Y(ori_ori_n349_));
  NA2        o327(.A(ori_ori_n349_), .B(ori_ori_n96_), .Y(ori_ori_n350_));
  AOI210     o328(.A0(ori_ori_n295_), .A1(ori_ori_n101_), .B0(ori_ori_n227_), .Y(ori_ori_n351_));
  NOi21      o329(.An(ori_ori_n277_), .B(ori_ori_n117_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n228_), .Y(ori_ori_n353_));
  OAI210     o331(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n354_));
  AOI210     o332(.A0(ori_ori_n215_), .A1(ori_ori_n47_), .B0(ori_ori_n354_), .Y(ori_ori_n355_));
  NO4        o333(.A(ori_ori_n355_), .B(ori_ori_n353_), .C(ori_ori_n351_), .D(x08), .Y(ori_ori_n356_));
  NO2        o334(.A(ori_ori_n114_), .B(ori_ori_n28_), .Y(ori_ori_n357_));
  NO2        o335(.A(ori_ori_n357_), .B(ori_ori_n232_), .Y(ori_ori_n358_));
  OR3        o336(.A(ori_ori_n358_), .B(x12), .C(x03), .Y(ori_ori_n359_));
  NA3        o337(.A(ori_ori_n290_), .B(ori_ori_n108_), .C(x12), .Y(ori_ori_n360_));
  AO210      o338(.A0(ori_ori_n290_), .A1(ori_ori_n108_), .B0(ori_ori_n215_), .Y(ori_ori_n361_));
  NA4        o339(.A(ori_ori_n361_), .B(ori_ori_n360_), .C(ori_ori_n359_), .D(x08), .Y(ori_ori_n362_));
  INV        o340(.A(ori_ori_n362_), .Y(ori_ori_n363_));
  AOI210     o341(.A0(ori_ori_n356_), .A1(ori_ori_n350_), .B0(ori_ori_n363_), .Y(ori_ori_n364_));
  INV        o342(.A(x03), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n128_), .B(ori_ori_n43_), .Y(ori_ori_n366_));
  OAI210     o344(.A0(ori_ori_n366_), .A1(ori_ori_n365_), .B0(ori_ori_n157_), .Y(ori_ori_n367_));
  NA3        o345(.A(ori_ori_n358_), .B(ori_ori_n352_), .C(ori_ori_n286_), .Y(ori_ori_n368_));
  INV        o346(.A(x14), .Y(ori_ori_n369_));
  NO3        o347(.A(ori_ori_n144_), .B(ori_ori_n70_), .C(ori_ori_n53_), .Y(ori_ori_n370_));
  NO2        o348(.A(ori_ori_n370_), .B(ori_ori_n369_), .Y(ori_ori_n371_));
  NA3        o349(.A(ori_ori_n371_), .B(ori_ori_n368_), .C(ori_ori_n367_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n344_), .B(ori_ori_n57_), .Y(ori_ori_n373_));
  NOi21      o351(.An(ori_ori_n235_), .B(ori_ori_n132_), .Y(ori_ori_n374_));
  NO2        o352(.A(ori_ori_n44_), .B(x04), .Y(ori_ori_n375_));
  OAI210     o353(.A0(ori_ori_n375_), .A1(ori_ori_n374_), .B0(ori_ori_n95_), .Y(ori_ori_n376_));
  OAI210     o354(.A0(ori_ori_n373_), .A1(ori_ori_n86_), .B0(ori_ori_n376_), .Y(ori_ori_n377_));
  NO4        o355(.A(ori_ori_n377_), .B(ori_ori_n372_), .C(ori_ori_n364_), .D(ori_ori_n346_), .Y(ori06));
  INV        o356(.A(ori_ori_n88_), .Y(ori_ori_n381_));
  INV        o357(.A(ori_ori_n40_), .Y(ori_ori_n382_));
  INV        o358(.A(x13), .Y(ori_ori_n383_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NA2        m044(.A(mai_mai_n61_), .B(mai_mai_n48_), .Y(mai_mai_n67_));
  OAI210     m045(.A0(mai_mai_n30_), .A1(x11), .B0(mai_mai_n67_), .Y(mai_mai_n68_));
  AOI220     m046(.A0(mai_mai_n68_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n69_));
  AOI210     m047(.A0(mai_mai_n69_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA3        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n28_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(x11), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  NO2        m053(.A(x10), .B(x09), .Y(mai_mai_n76_));
  NO2        m054(.A(mai_mai_n437_), .B(mai_mai_n24_), .Y(mai_mai_n77_));
  NO2        m055(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n78_));
  NO2        m056(.A(mai_mai_n78_), .B(mai_mai_n36_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n78_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n80_));
  AOI210     m058(.A0(mai_mai_n79_), .A1(mai_mai_n48_), .B0(mai_mai_n80_), .Y(mai_mai_n81_));
  NO2        m059(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n82_));
  NO2        m060(.A(x08), .B(x01), .Y(mai_mai_n83_));
  OAI210     m061(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n35_), .Y(mai_mai_n84_));
  NA2        m062(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n84_), .B(mai_mai_n81_), .C(mai_mai_n77_), .Y(mai_mai_n86_));
  AN2        m064(.A(mai_mai_n86_), .B(mai_mai_n74_), .Y(mai_mai_n87_));
  INV        m065(.A(mai_mai_n84_), .Y(mai_mai_n88_));
  NO2        m066(.A(x06), .B(x05), .Y(mai_mai_n89_));
  NA2        m067(.A(x11), .B(x00), .Y(mai_mai_n90_));
  NO2        m068(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n91_));
  NOi21      m069(.An(mai_mai_n90_), .B(mai_mai_n91_), .Y(mai_mai_n92_));
  AOI210     m070(.A0(mai_mai_n89_), .A1(mai_mai_n88_), .B0(mai_mai_n92_), .Y(mai_mai_n93_));
  NOi21      m071(.An(x01), .B(x10), .Y(mai_mai_n94_));
  NO2        m072(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n95_));
  NO3        m073(.A(mai_mai_n95_), .B(mai_mai_n94_), .C(x06), .Y(mai_mai_n96_));
  NA2        m074(.A(mai_mai_n96_), .B(mai_mai_n27_), .Y(mai_mai_n97_));
  OAI210     m075(.A0(mai_mai_n93_), .A1(x07), .B0(mai_mai_n97_), .Y(mai_mai_n98_));
  NO3        m076(.A(mai_mai_n98_), .B(mai_mai_n87_), .C(mai_mai_n70_), .Y(mai01));
  INV        m077(.A(x12), .Y(mai_mai_n100_));
  INV        m078(.A(x13), .Y(mai_mai_n101_));
  NA2        m079(.A(x08), .B(x04), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n102_), .B(mai_mai_n57_), .Y(mai_mai_n103_));
  NA2        m081(.A(mai_mai_n103_), .B(mai_mai_n89_), .Y(mai_mai_n104_));
  NA2        m082(.A(mai_mai_n94_), .B(mai_mai_n28_), .Y(mai_mai_n105_));
  NO2        m083(.A(mai_mai_n105_), .B(mai_mai_n71_), .Y(mai_mai_n106_));
  NO2        m084(.A(x10), .B(x01), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n108_));
  NO2        m086(.A(mai_mai_n108_), .B(mai_mai_n107_), .Y(mai_mai_n109_));
  NA2        m087(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n110_));
  NO3        m088(.A(mai_mai_n110_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n111_));
  AOI210     m089(.A0(mai_mai_n111_), .A1(mai_mai_n109_), .B0(mai_mai_n106_), .Y(mai_mai_n112_));
  AOI210     m090(.A0(mai_mai_n112_), .A1(mai_mai_n104_), .B0(mai_mai_n101_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n114_));
  NOi21      m092(.An(mai_mai_n114_), .B(mai_mai_n58_), .Y(mai_mai_n115_));
  NO2        m093(.A(mai_mai_n35_), .B(x02), .Y(mai_mai_n116_));
  NO2        m094(.A(mai_mai_n101_), .B(mai_mai_n36_), .Y(mai_mai_n117_));
  NA3        m095(.A(mai_mai_n117_), .B(mai_mai_n116_), .C(x06), .Y(mai_mai_n118_));
  INV        m096(.A(mai_mai_n118_), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n83_), .B(x13), .Y(mai_mai_n120_));
  NA2        m098(.A(x09), .B(mai_mai_n35_), .Y(mai_mai_n121_));
  NO2        m099(.A(mai_mai_n121_), .B(mai_mai_n120_), .Y(mai_mai_n122_));
  NA2        m100(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n123_));
  NO2        m101(.A(mai_mai_n123_), .B(x05), .Y(mai_mai_n124_));
  NO2        m102(.A(mai_mai_n124_), .B(mai_mai_n122_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n126_));
  AOI210     m104(.A0(mai_mai_n57_), .A1(mai_mai_n79_), .B0(mai_mai_n115_), .Y(mai_mai_n127_));
  AOI210     m105(.A0(mai_mai_n127_), .A1(mai_mai_n125_), .B0(mai_mai_n72_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n129_));
  NA2        m107(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(mai_mai_n129_), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n132_));
  NO3        m110(.A(mai_mai_n126_), .B(mai_mai_n78_), .C(mai_mai_n36_), .Y(mai_mai_n133_));
  NO2        m111(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n134_));
  NO3        m112(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n131_), .Y(mai_mai_n135_));
  NO3        m113(.A(mai_mai_n135_), .B(x06), .C(x03), .Y(mai_mai_n136_));
  NO4        m114(.A(mai_mai_n136_), .B(mai_mai_n128_), .C(mai_mai_n119_), .D(mai_mai_n113_), .Y(mai_mai_n137_));
  NA2        m115(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n138_));
  OAI210     m116(.A0(mai_mai_n83_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n139_));
  NO2        m117(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n140_));
  NA2        m118(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n141_));
  AN2        m119(.A(x01), .B(mai_mai_n83_), .Y(mai_mai_n142_));
  NO2        m120(.A(x09), .B(x05), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(mai_mai_n47_), .Y(mai_mai_n144_));
  AOI210     m122(.A0(mai_mai_n144_), .A1(mai_mai_n109_), .B0(mai_mai_n49_), .Y(mai_mai_n145_));
  NA2        m123(.A(x09), .B(x00), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n114_), .B(mai_mai_n146_), .Y(mai_mai_n147_));
  NA2        m125(.A(mai_mai_n75_), .B(mai_mai_n51_), .Y(mai_mai_n148_));
  AOI210     m126(.A0(mai_mai_n148_), .A1(mai_mai_n147_), .B0(mai_mai_n141_), .Y(mai_mai_n149_));
  NO3        m127(.A(mai_mai_n149_), .B(mai_mai_n145_), .C(mai_mai_n142_), .Y(mai_mai_n150_));
  NO2        m128(.A(x03), .B(x02), .Y(mai_mai_n151_));
  NA2        m129(.A(mai_mai_n84_), .B(mai_mai_n101_), .Y(mai_mai_n152_));
  OAI210     m130(.A0(mai_mai_n152_), .A1(mai_mai_n115_), .B0(mai_mai_n151_), .Y(mai_mai_n153_));
  OA210      m131(.A0(mai_mai_n150_), .A1(x11), .B0(mai_mai_n153_), .Y(mai_mai_n154_));
  OAI210     m132(.A0(mai_mai_n137_), .A1(mai_mai_n23_), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  NA2        m133(.A(mai_mai_n109_), .B(mai_mai_n40_), .Y(mai_mai_n156_));
  NAi21      m134(.An(x06), .B(x10), .Y(mai_mai_n157_));
  NOi21      m135(.An(x01), .B(x13), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  BUFFER     m137(.A(mai_mai_n159_), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n160_), .A1(mai_mai_n156_), .B0(mai_mai_n41_), .Y(mai_mai_n161_));
  NO2        m139(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n162_));
  NA2        m140(.A(mai_mai_n101_), .B(x01), .Y(mai_mai_n163_));
  NO2        m141(.A(mai_mai_n163_), .B(x08), .Y(mai_mai_n164_));
  OAI210     m142(.A0(x05), .A1(mai_mai_n164_), .B0(mai_mai_n51_), .Y(mai_mai_n165_));
  AOI210     m143(.A0(mai_mai_n165_), .A1(mai_mai_n162_), .B0(mai_mai_n48_), .Y(mai_mai_n166_));
  AOI210     m144(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n167_));
  OAI210     m145(.A0(mai_mai_n166_), .A1(mai_mai_n161_), .B0(mai_mai_n167_), .Y(mai_mai_n168_));
  NA2        m146(.A(x04), .B(x02), .Y(mai_mai_n169_));
  NA2        m147(.A(x10), .B(x05), .Y(mai_mai_n170_));
  NA2        m148(.A(x09), .B(x06), .Y(mai_mai_n171_));
  AOI210     m149(.A0(mai_mai_n171_), .A1(mai_mai_n170_), .B0(x11), .Y(mai_mai_n172_));
  NO2        m150(.A(x09), .B(x01), .Y(mai_mai_n173_));
  NO3        m151(.A(mai_mai_n173_), .B(mai_mai_n107_), .C(mai_mai_n31_), .Y(mai_mai_n174_));
  OAI210     m152(.A0(mai_mai_n174_), .A1(mai_mai_n172_), .B0(x00), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n114_), .B(x08), .Y(mai_mai_n176_));
  OAI210     m154(.A0(mai_mai_n441_), .A1(x11), .B0(mai_mai_n175_), .Y(mai_mai_n177_));
  NAi21      m155(.An(mai_mai_n169_), .B(mai_mai_n177_), .Y(mai_mai_n178_));
  INV        m156(.A(mai_mai_n25_), .Y(mai_mai_n179_));
  NAi21      m157(.An(x13), .B(x00), .Y(mai_mai_n180_));
  AOI210     m158(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n180_), .Y(mai_mai_n181_));
  AOI220     m159(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n182_));
  OAI210     m160(.A0(mai_mai_n170_), .A1(mai_mai_n35_), .B0(mai_mai_n182_), .Y(mai_mai_n183_));
  AN2        m161(.A(mai_mai_n183_), .B(mai_mai_n181_), .Y(mai_mai_n184_));
  NO2        m162(.A(mai_mai_n180_), .B(mai_mai_n36_), .Y(mai_mai_n185_));
  INV        m163(.A(mai_mai_n185_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n186_), .B(mai_mai_n171_), .Y(mai_mai_n187_));
  OAI210     m165(.A0(mai_mai_n187_), .A1(mai_mai_n184_), .B0(mai_mai_n179_), .Y(mai_mai_n188_));
  NOi21      m166(.An(x09), .B(x00), .Y(mai_mai_n189_));
  NO3        m167(.A(mai_mai_n82_), .B(mai_mai_n189_), .C(mai_mai_n47_), .Y(mai_mai_n190_));
  NA2        m168(.A(mai_mai_n190_), .B(mai_mai_n130_), .Y(mai_mai_n191_));
  NA2        m169(.A(x10), .B(x08), .Y(mai_mai_n192_));
  INV        m170(.A(mai_mai_n192_), .Y(mai_mai_n193_));
  NA2        m171(.A(x06), .B(x05), .Y(mai_mai_n194_));
  OAI210     m172(.A0(mai_mai_n194_), .A1(mai_mai_n35_), .B0(mai_mai_n100_), .Y(mai_mai_n195_));
  NA2        m173(.A(mai_mai_n100_), .B(mai_mai_n191_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n101_), .B(x12), .Y(mai_mai_n197_));
  AOI210     m175(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n197_), .Y(mai_mai_n198_));
  NA2        m176(.A(mai_mai_n94_), .B(mai_mai_n51_), .Y(mai_mai_n199_));
  NO2        m177(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n200_));
  NA2        m178(.A(mai_mai_n200_), .B(x02), .Y(mai_mai_n201_));
  NO2        m179(.A(mai_mai_n201_), .B(mai_mai_n199_), .Y(mai_mai_n202_));
  AOI210     m180(.A0(mai_mai_n198_), .A1(mai_mai_n196_), .B0(mai_mai_n202_), .Y(mai_mai_n203_));
  NA4        m181(.A(mai_mai_n203_), .B(mai_mai_n188_), .C(mai_mai_n178_), .D(mai_mai_n168_), .Y(mai_mai_n204_));
  AOI210     m182(.A0(mai_mai_n155_), .A1(mai_mai_n100_), .B0(mai_mai_n204_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n206_));
  NA2        m184(.A(mai_mai_n206_), .B(mai_mai_n139_), .Y(mai_mai_n207_));
  AOI210     m185(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n208_));
  NO2        m186(.A(mai_mai_n129_), .B(x06), .Y(mai_mai_n209_));
  AOI210     m187(.A0(mai_mai_n208_), .A1(mai_mai_n207_), .B0(mai_mai_n209_), .Y(mai_mai_n210_));
  NO2        m188(.A(mai_mai_n210_), .B(x12), .Y(mai_mai_n211_));
  INV        m189(.A(mai_mai_n75_), .Y(mai_mai_n212_));
  AOI210     m190(.A0(mai_mai_n192_), .A1(x05), .B0(mai_mai_n51_), .Y(mai_mai_n213_));
  OAI210     m191(.A0(mai_mai_n213_), .A1(mai_mai_n159_), .B0(mai_mai_n57_), .Y(mai_mai_n214_));
  NA2        m192(.A(mai_mai_n214_), .B(mai_mai_n212_), .Y(mai_mai_n215_));
  NO2        m193(.A(mai_mai_n94_), .B(x06), .Y(mai_mai_n216_));
  NA4        m194(.A(mai_mai_n157_), .B(mai_mai_n56_), .C(mai_mai_n36_), .D(x04), .Y(mai_mai_n217_));
  NA2        m195(.A(mai_mai_n217_), .B(mai_mai_n141_), .Y(mai_mai_n218_));
  NA2        m196(.A(mai_mai_n218_), .B(x02), .Y(mai_mai_n219_));
  AOI210     m197(.A0(mai_mai_n219_), .A1(mai_mai_n215_), .B0(mai_mai_n23_), .Y(mai_mai_n220_));
  OAI210     m198(.A0(mai_mai_n211_), .A1(mai_mai_n57_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  INV        m199(.A(mai_mai_n141_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n223_));
  OAI210     m201(.A0(mai_mai_n78_), .A1(mai_mai_n36_), .B0(mai_mai_n121_), .Y(mai_mai_n224_));
  NO2        m202(.A(mai_mai_n101_), .B(x03), .Y(mai_mai_n225_));
  AOI220     m203(.A0(mai_mai_n225_), .A1(mai_mai_n224_), .B0(mai_mai_n75_), .B1(mai_mai_n223_), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n32_), .B(x06), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n157_), .Y(mai_mai_n228_));
  NOi21      m206(.An(x13), .B(x04), .Y(mai_mai_n229_));
  NO3        m207(.A(mai_mai_n229_), .B(mai_mai_n75_), .C(mai_mai_n189_), .Y(mai_mai_n230_));
  NO2        m208(.A(mai_mai_n230_), .B(x05), .Y(mai_mai_n231_));
  AOI220     m209(.A0(mai_mai_n231_), .A1(mai_mai_n227_), .B0(mai_mai_n228_), .B1(mai_mai_n57_), .Y(mai_mai_n232_));
  OAI210     m210(.A0(mai_mai_n226_), .A1(mai_mai_n222_), .B0(mai_mai_n232_), .Y(mai_mai_n233_));
  INV        m211(.A(mai_mai_n91_), .Y(mai_mai_n234_));
  NO2        m212(.A(mai_mai_n234_), .B(x12), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n51_), .B(mai_mai_n36_), .Y(mai_mai_n237_));
  OAI210     m215(.A0(mai_mai_n237_), .A1(mai_mai_n183_), .B0(mai_mai_n181_), .Y(mai_mai_n238_));
  AOI210     m216(.A0(x08), .A1(x04), .B0(x09), .Y(mai_mai_n239_));
  NO2        m217(.A(x06), .B(x00), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n146_), .B(mai_mai_n72_), .Y(mai_mai_n241_));
  INV        m219(.A(mai_mai_n241_), .Y(mai_mai_n242_));
  NA2        m220(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n243_));
  NA2        m221(.A(mai_mai_n243_), .B(x03), .Y(mai_mai_n244_));
  OA210      m222(.A0(mai_mai_n244_), .A1(mai_mai_n242_), .B0(mai_mai_n238_), .Y(mai_mai_n245_));
  NA2        m223(.A(x13), .B(mai_mai_n100_), .Y(mai_mai_n246_));
  NA3        m224(.A(mai_mai_n246_), .B(mai_mai_n195_), .C(mai_mai_n92_), .Y(mai_mai_n247_));
  OAI210     m225(.A0(mai_mai_n245_), .A1(mai_mai_n236_), .B0(mai_mai_n247_), .Y(mai_mai_n248_));
  AOI210     m226(.A0(mai_mai_n235_), .A1(mai_mai_n233_), .B0(mai_mai_n248_), .Y(mai_mai_n249_));
  AOI210     m227(.A0(mai_mai_n249_), .A1(mai_mai_n221_), .B0(x07), .Y(mai_mai_n250_));
  NA2        m228(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n251_));
  AOI210     m229(.A0(mai_mai_n138_), .A1(mai_mai_n148_), .B0(mai_mai_n251_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n101_), .B(x06), .Y(mai_mai_n253_));
  INV        m231(.A(mai_mai_n253_), .Y(mai_mai_n254_));
  NO2        m232(.A(x08), .B(x05), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n255_), .B(mai_mai_n239_), .Y(mai_mai_n256_));
  OAI210     m234(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n257_));
  OAI210     m235(.A0(mai_mai_n256_), .A1(mai_mai_n254_), .B0(mai_mai_n257_), .Y(mai_mai_n258_));
  NO2        m236(.A(x12), .B(x02), .Y(mai_mai_n259_));
  INV        m237(.A(mai_mai_n259_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n260_), .B(mai_mai_n234_), .Y(mai_mai_n261_));
  OA210      m239(.A0(mai_mai_n258_), .A1(mai_mai_n252_), .B0(mai_mai_n261_), .Y(mai_mai_n262_));
  NA2        m240(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n263_));
  NO2        m241(.A(mai_mai_n263_), .B(x01), .Y(mai_mai_n264_));
  NOi21      m242(.An(mai_mai_n83_), .B(mai_mai_n121_), .Y(mai_mai_n265_));
  NO2        m243(.A(mai_mai_n265_), .B(mai_mai_n264_), .Y(mai_mai_n266_));
  NO2        m244(.A(mai_mai_n266_), .B(mai_mai_n29_), .Y(mai_mai_n267_));
  NA2        m245(.A(mai_mai_n253_), .B(mai_mai_n224_), .Y(mai_mai_n268_));
  NA2        m246(.A(mai_mai_n101_), .B(x04), .Y(mai_mai_n269_));
  NA2        m247(.A(mai_mai_n269_), .B(mai_mai_n28_), .Y(mai_mai_n270_));
  OAI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n120_), .B0(mai_mai_n268_), .Y(mai_mai_n271_));
  NO3        m249(.A(mai_mai_n90_), .B(x12), .C(x03), .Y(mai_mai_n272_));
  OAI210     m250(.A0(mai_mai_n271_), .A1(mai_mai_n267_), .B0(mai_mai_n272_), .Y(mai_mai_n273_));
  AOI210     m251(.A0(mai_mai_n199_), .A1(mai_mai_n194_), .B0(mai_mai_n102_), .Y(mai_mai_n274_));
  NOi21      m252(.An(mai_mai_n251_), .B(mai_mai_n216_), .Y(mai_mai_n275_));
  NO2        m253(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n276_));
  OAI210     m254(.A0(mai_mai_n275_), .A1(mai_mai_n274_), .B0(mai_mai_n276_), .Y(mai_mai_n277_));
  NO2        m255(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n236_), .B(mai_mai_n28_), .Y(mai_mai_n279_));
  NA2        m257(.A(mai_mai_n222_), .B(mai_mai_n279_), .Y(mai_mai_n280_));
  NA3        m258(.A(mai_mai_n280_), .B(mai_mai_n277_), .C(mai_mai_n273_), .Y(mai_mai_n281_));
  NO3        m259(.A(mai_mai_n281_), .B(mai_mai_n262_), .C(mai_mai_n250_), .Y(mai_mai_n282_));
  OAI210     m260(.A0(mai_mai_n205_), .A1(mai_mai_n61_), .B0(mai_mai_n282_), .Y(mai02));
  NOi21      m261(.An(mai_mai_n230_), .B(mai_mai_n173_), .Y(mai_mai_n284_));
  NO2        m262(.A(mai_mai_n101_), .B(mai_mai_n35_), .Y(mai_mai_n285_));
  NA3        m263(.A(mai_mai_n285_), .B(mai_mai_n193_), .C(mai_mai_n56_), .Y(mai_mai_n286_));
  OAI210     m264(.A0(mai_mai_n284_), .A1(mai_mai_n32_), .B0(mai_mai_n286_), .Y(mai_mai_n287_));
  NA2        m265(.A(mai_mai_n287_), .B(mai_mai_n170_), .Y(mai_mai_n288_));
  INV        m266(.A(mai_mai_n170_), .Y(mai_mai_n289_));
  AOI210     m267(.A0(mai_mai_n116_), .A1(mai_mai_n85_), .B0(x09), .Y(mai_mai_n290_));
  OAI220     m268(.A0(mai_mai_n290_), .A1(mai_mai_n101_), .B0(mai_mai_n84_), .B1(mai_mai_n51_), .Y(mai_mai_n291_));
  AOI220     m269(.A0(mai_mai_n291_), .A1(mai_mai_n289_), .B0(mai_mai_n152_), .B1(mai_mai_n151_), .Y(mai_mai_n292_));
  AOI210     m270(.A0(mai_mai_n292_), .A1(mai_mai_n288_), .B0(mai_mai_n48_), .Y(mai_mai_n293_));
  NO2        m271(.A(x05), .B(x02), .Y(mai_mai_n294_));
  OAI210     m272(.A0(mai_mai_n207_), .A1(mai_mai_n189_), .B0(mai_mai_n294_), .Y(mai_mai_n295_));
  AOI220     m273(.A0(mai_mai_n255_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n296_));
  NOi21      m274(.An(mai_mai_n285_), .B(mai_mai_n296_), .Y(mai_mai_n297_));
  AOI210     m275(.A0(mai_mai_n229_), .A1(mai_mai_n78_), .B0(mai_mai_n297_), .Y(mai_mai_n298_));
  AOI210     m276(.A0(mai_mai_n298_), .A1(mai_mai_n295_), .B0(mai_mai_n141_), .Y(mai_mai_n299_));
  NAi21      m277(.An(mai_mai_n231_), .B(mai_mai_n226_), .Y(mai_mai_n300_));
  NO2        m278(.A(mai_mai_n243_), .B(mai_mai_n47_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n301_), .B(mai_mai_n300_), .Y(mai_mai_n302_));
  AN2        m280(.A(mai_mai_n225_), .B(mai_mai_n224_), .Y(mai_mai_n303_));
  OAI210     m281(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n304_));
  NA2        m282(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n305_));
  BUFFER     m283(.A(mai_mai_n144_), .Y(mai_mai_n306_));
  AOI210     m284(.A0(mai_mai_n306_), .A1(mai_mai_n139_), .B0(mai_mai_n304_), .Y(mai_mai_n307_));
  OAI210     m285(.A0(mai_mai_n307_), .A1(mai_mai_n303_), .B0(mai_mai_n95_), .Y(mai_mai_n308_));
  NA3        m286(.A(mai_mai_n95_), .B(mai_mai_n83_), .C(mai_mai_n223_), .Y(mai_mai_n309_));
  NA3        m287(.A(mai_mai_n94_), .B(mai_mai_n82_), .C(mai_mai_n42_), .Y(mai_mai_n310_));
  AOI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n309_), .B0(x04), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n151_), .Y(mai_mai_n312_));
  OAI220     m290(.A0(mai_mai_n256_), .A1(mai_mai_n105_), .B0(mai_mai_n312_), .B1(mai_mai_n131_), .Y(mai_mai_n313_));
  AOI210     m291(.A0(mai_mai_n313_), .A1(x13), .B0(mai_mai_n311_), .Y(mai_mai_n314_));
  NA3        m292(.A(mai_mai_n314_), .B(mai_mai_n308_), .C(mai_mai_n302_), .Y(mai_mai_n315_));
  NO3        m293(.A(mai_mai_n315_), .B(mai_mai_n299_), .C(mai_mai_n293_), .Y(mai_mai_n316_));
  NA2        m294(.A(mai_mai_n140_), .B(x03), .Y(mai_mai_n317_));
  INV        m295(.A(mai_mai_n180_), .Y(mai_mai_n318_));
  OAI210     m296(.A0(mai_mai_n51_), .A1(mai_mai_n35_), .B0(mai_mai_n36_), .Y(mai_mai_n319_));
  AOI220     m297(.A0(mai_mai_n319_), .A1(mai_mai_n318_), .B0(mai_mai_n200_), .B1(x08), .Y(mai_mai_n320_));
  OAI210     m298(.A0(mai_mai_n320_), .A1(mai_mai_n278_), .B0(mai_mai_n317_), .Y(mai_mai_n321_));
  NA2        m299(.A(mai_mai_n321_), .B(mai_mai_n107_), .Y(mai_mai_n322_));
  NA2        m300(.A(mai_mai_n169_), .B(mai_mai_n163_), .Y(mai_mai_n323_));
  AN2        m301(.A(mai_mai_n323_), .B(mai_mai_n176_), .Y(mai_mai_n324_));
  INV        m302(.A(mai_mai_n56_), .Y(mai_mai_n325_));
  OAI220     m303(.A0(mai_mai_n269_), .A1(mai_mai_n325_), .B0(mai_mai_n132_), .B1(mai_mai_n28_), .Y(mai_mai_n326_));
  OAI210     m304(.A0(mai_mai_n326_), .A1(mai_mai_n324_), .B0(mai_mai_n108_), .Y(mai_mai_n327_));
  NA2        m305(.A(mai_mai_n269_), .B(mai_mai_n100_), .Y(mai_mai_n328_));
  NA2        m306(.A(mai_mai_n100_), .B(mai_mai_n41_), .Y(mai_mai_n329_));
  NA3        m307(.A(mai_mai_n329_), .B(mai_mai_n328_), .C(mai_mai_n131_), .Y(mai_mai_n330_));
  NA4        m308(.A(mai_mai_n330_), .B(mai_mai_n327_), .C(mai_mai_n322_), .D(mai_mai_n48_), .Y(mai_mai_n331_));
  INV        m309(.A(mai_mai_n200_), .Y(mai_mai_n332_));
  NO2        m310(.A(mai_mai_n164_), .B(mai_mai_n40_), .Y(mai_mai_n333_));
  NA2        m311(.A(mai_mai_n32_), .B(x05), .Y(mai_mai_n334_));
  OAI220     m312(.A0(mai_mai_n334_), .A1(mai_mai_n333_), .B0(mai_mai_n332_), .B1(mai_mai_n59_), .Y(mai_mai_n335_));
  NA2        m313(.A(mai_mai_n335_), .B(x02), .Y(mai_mai_n336_));
  INV        m314(.A(mai_mai_n237_), .Y(mai_mai_n337_));
  NA2        m315(.A(mai_mai_n197_), .B(x04), .Y(mai_mai_n338_));
  NO2        m316(.A(mai_mai_n338_), .B(mai_mai_n337_), .Y(mai_mai_n339_));
  NO3        m317(.A(mai_mai_n182_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n340_));
  OAI210     m318(.A0(mai_mai_n340_), .A1(mai_mai_n339_), .B0(mai_mai_n95_), .Y(mai_mai_n341_));
  NO3        m319(.A(mai_mai_n197_), .B(mai_mai_n162_), .C(mai_mai_n52_), .Y(mai_mai_n342_));
  OAI210     m320(.A0(mai_mai_n146_), .A1(mai_mai_n36_), .B0(mai_mai_n100_), .Y(mai_mai_n343_));
  OAI210     m321(.A0(mai_mai_n343_), .A1(mai_mai_n190_), .B0(mai_mai_n342_), .Y(mai_mai_n344_));
  NA4        m322(.A(mai_mai_n344_), .B(mai_mai_n341_), .C(mai_mai_n336_), .D(x06), .Y(mai_mai_n345_));
  NA2        m323(.A(x09), .B(x03), .Y(mai_mai_n346_));
  OAI220     m324(.A0(mai_mai_n346_), .A1(mai_mai_n130_), .B0(mai_mai_n206_), .B1(mai_mai_n64_), .Y(mai_mai_n347_));
  OAI220     m325(.A0(mai_mai_n163_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n348_));
  NA2        m326(.A(mai_mai_n348_), .B(mai_mai_n222_), .Y(mai_mai_n349_));
  NO2        m327(.A(mai_mai_n349_), .B(mai_mai_n28_), .Y(mai_mai_n350_));
  AO220      m328(.A0(mai_mai_n350_), .A1(x04), .B0(mai_mai_n347_), .B1(x05), .Y(mai_mai_n351_));
  AOI210     m329(.A0(mai_mai_n345_), .A1(mai_mai_n331_), .B0(mai_mai_n351_), .Y(mai_mai_n352_));
  OAI210     m330(.A0(mai_mai_n316_), .A1(x12), .B0(mai_mai_n352_), .Y(mai03));
  OR2        m331(.A(mai_mai_n42_), .B(mai_mai_n223_), .Y(mai_mai_n354_));
  AOI210     m332(.A0(mai_mai_n152_), .A1(mai_mai_n100_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  AO210      m333(.A0(mai_mai_n337_), .A1(mai_mai_n85_), .B0(mai_mai_n338_), .Y(mai_mai_n356_));
  NA2        m334(.A(mai_mai_n197_), .B(mai_mai_n151_), .Y(mai_mai_n357_));
  NA3        m335(.A(mai_mai_n357_), .B(mai_mai_n356_), .C(mai_mai_n201_), .Y(mai_mai_n358_));
  OAI210     m336(.A0(mai_mai_n358_), .A1(mai_mai_n355_), .B0(x05), .Y(mai_mai_n359_));
  NA2        m337(.A(mai_mai_n354_), .B(x05), .Y(mai_mai_n360_));
  AOI210     m338(.A0(mai_mai_n139_), .A1(mai_mai_n212_), .B0(mai_mai_n360_), .Y(mai_mai_n361_));
  AOI210     m339(.A0(mai_mai_n225_), .A1(mai_mai_n79_), .B0(mai_mai_n124_), .Y(mai_mai_n362_));
  OAI220     m340(.A0(mai_mai_n362_), .A1(mai_mai_n59_), .B0(mai_mai_n305_), .B1(mai_mai_n296_), .Y(mai_mai_n363_));
  OAI210     m341(.A0(mai_mai_n363_), .A1(mai_mai_n361_), .B0(mai_mai_n100_), .Y(mai_mai_n364_));
  AOI210     m342(.A0(mai_mai_n144_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n365_));
  NO2        m343(.A(mai_mai_n173_), .B(mai_mai_n134_), .Y(mai_mai_n366_));
  OAI220     m344(.A0(mai_mai_n366_), .A1(mai_mai_n37_), .B0(mai_mai_n147_), .B1(x13), .Y(mai_mai_n367_));
  OAI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n365_), .B0(x04), .Y(mai_mai_n368_));
  NO3        m346(.A(mai_mai_n329_), .B(mai_mai_n84_), .C(mai_mai_n59_), .Y(mai_mai_n369_));
  AOI210     m347(.A0(mai_mai_n186_), .A1(mai_mai_n100_), .B0(mai_mai_n144_), .Y(mai_mai_n370_));
  OA210      m348(.A0(mai_mai_n164_), .A1(x12), .B0(mai_mai_n134_), .Y(mai_mai_n371_));
  NO3        m349(.A(mai_mai_n371_), .B(mai_mai_n370_), .C(mai_mai_n369_), .Y(mai_mai_n372_));
  NA4        m350(.A(mai_mai_n372_), .B(mai_mai_n368_), .C(mai_mai_n364_), .D(mai_mai_n359_), .Y(mai04));
  NO2        m351(.A(mai_mai_n88_), .B(mai_mai_n39_), .Y(mai_mai_n374_));
  XO2        m352(.A(mai_mai_n374_), .B(mai_mai_n246_), .Y(mai05));
  NO2        m353(.A(mai_mai_n304_), .B(mai_mai_n25_), .Y(mai_mai_n376_));
  NAi41      m354(.An(mai_mai_n76_), .B(mai_mai_n141_), .C(mai_mai_n132_), .D(mai_mai_n31_), .Y(mai_mai_n377_));
  AOI210     m355(.A0(mai_mai_n439_), .A1(mai_mai_n377_), .B0(mai_mai_n24_), .Y(mai_mai_n378_));
  OAI210     m356(.A0(mai_mai_n378_), .A1(mai_mai_n376_), .B0(mai_mai_n100_), .Y(mai_mai_n379_));
  NA2        m357(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n380_));
  NA2        m358(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n381_));
  NA2        m359(.A(mai_mai_n251_), .B(x03), .Y(mai_mai_n382_));
  OAI220     m360(.A0(mai_mai_n382_), .A1(mai_mai_n381_), .B0(mai_mai_n380_), .B1(mai_mai_n80_), .Y(mai_mai_n383_));
  OAI210     m361(.A0(mai_mai_n26_), .A1(mai_mai_n100_), .B0(x07), .Y(mai_mai_n384_));
  AOI210     m362(.A0(mai_mai_n383_), .A1(x06), .B0(mai_mai_n384_), .Y(mai_mai_n385_));
  NA2        m363(.A(mai_mai_n440_), .B(mai_mai_n382_), .Y(mai_mai_n386_));
  OR2        m364(.A(mai_mai_n386_), .B(mai_mai_n236_), .Y(mai_mai_n387_));
  NA2        m365(.A(mai_mai_n158_), .B(x05), .Y(mai_mai_n388_));
  NA3        m366(.A(mai_mai_n388_), .B(mai_mai_n240_), .C(mai_mai_n234_), .Y(mai_mai_n389_));
  NO2        m367(.A(mai_mai_n23_), .B(x10), .Y(mai_mai_n390_));
  OAI210     m368(.A0(x11), .A1(mai_mai_n29_), .B0(mai_mai_n48_), .Y(mai_mai_n391_));
  OR3        m369(.A(mai_mai_n391_), .B(mai_mai_n390_), .C(mai_mai_n44_), .Y(mai_mai_n392_));
  NA3        m370(.A(mai_mai_n392_), .B(mai_mai_n389_), .C(mai_mai_n387_), .Y(mai_mai_n393_));
  NA2        m371(.A(mai_mai_n393_), .B(mai_mai_n100_), .Y(mai_mai_n394_));
  NA2        m372(.A(mai_mai_n33_), .B(mai_mai_n100_), .Y(mai_mai_n395_));
  AOI210     m373(.A0(mai_mai_n395_), .A1(mai_mai_n91_), .B0(x07), .Y(mai_mai_n396_));
  AOI220     m374(.A0(mai_mai_n396_), .A1(mai_mai_n394_), .B0(mai_mai_n385_), .B1(mai_mai_n379_), .Y(mai_mai_n397_));
  AOI210     m375(.A0(mai_mai_n390_), .A1(x07), .B0(mai_mai_n140_), .Y(mai_mai_n398_));
  OR2        m376(.A(mai_mai_n398_), .B(x03), .Y(mai_mai_n399_));
  NO2        m377(.A(x07), .B(x11), .Y(mai_mai_n400_));
  NO3        m378(.A(mai_mai_n400_), .B(mai_mai_n143_), .C(mai_mai_n28_), .Y(mai_mai_n401_));
  AOI210     m379(.A0(mai_mai_n401_), .A1(mai_mai_n399_), .B0(mai_mai_n47_), .Y(mai_mai_n402_));
  NA2        m380(.A(mai_mai_n402_), .B(mai_mai_n101_), .Y(mai_mai_n403_));
  AOI210     m381(.A0(mai_mai_n338_), .A1(mai_mai_n110_), .B0(mai_mai_n259_), .Y(mai_mai_n404_));
  NOi21      m382(.An(mai_mai_n317_), .B(mai_mai_n134_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n405_), .B(mai_mai_n260_), .Y(mai_mai_n406_));
  OAI210     m384(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n407_));
  AOI210     m385(.A0(mai_mai_n246_), .A1(mai_mai_n47_), .B0(mai_mai_n407_), .Y(mai_mai_n408_));
  NO4        m386(.A(mai_mai_n408_), .B(mai_mai_n406_), .C(mai_mai_n404_), .D(x08), .Y(mai_mai_n409_));
  NO2        m387(.A(x05), .B(x03), .Y(mai_mai_n410_));
  NO2        m388(.A(x13), .B(x12), .Y(mai_mai_n411_));
  NO2        m389(.A(mai_mai_n132_), .B(mai_mai_n28_), .Y(mai_mai_n412_));
  NO2        m390(.A(mai_mai_n412_), .B(mai_mai_n264_), .Y(mai_mai_n413_));
  OR3        m391(.A(mai_mai_n413_), .B(x12), .C(x03), .Y(mai_mai_n414_));
  NA3        m392(.A(mai_mai_n332_), .B(mai_mai_n126_), .C(x12), .Y(mai_mai_n415_));
  AO210      m393(.A0(mai_mai_n332_), .A1(mai_mai_n126_), .B0(mai_mai_n246_), .Y(mai_mai_n416_));
  NA4        m394(.A(mai_mai_n416_), .B(mai_mai_n415_), .C(mai_mai_n414_), .D(x08), .Y(mai_mai_n417_));
  AOI210     m395(.A0(mai_mai_n411_), .A1(mai_mai_n410_), .B0(mai_mai_n417_), .Y(mai_mai_n418_));
  AOI210     m396(.A0(mai_mai_n409_), .A1(mai_mai_n403_), .B0(mai_mai_n418_), .Y(mai_mai_n419_));
  OAI210     m397(.A0(x07), .A1(mai_mai_n23_), .B0(x03), .Y(mai_mai_n420_));
  OAI220     m398(.A0(mai_mai_n438_), .A1(mai_mai_n381_), .B0(mai_mai_n143_), .B1(mai_mai_n43_), .Y(mai_mai_n421_));
  OAI210     m399(.A0(mai_mai_n421_), .A1(mai_mai_n420_), .B0(mai_mai_n185_), .Y(mai_mai_n422_));
  NA3        m400(.A(mai_mai_n413_), .B(mai_mai_n405_), .C(mai_mai_n328_), .Y(mai_mai_n423_));
  INV        m401(.A(x14), .Y(mai_mai_n424_));
  NO3        m402(.A(mai_mai_n317_), .B(mai_mai_n105_), .C(x11), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n425_), .B(mai_mai_n424_), .Y(mai_mai_n426_));
  NA3        m404(.A(mai_mai_n426_), .B(mai_mai_n423_), .C(mai_mai_n422_), .Y(mai_mai_n427_));
  AOI220     m405(.A0(mai_mai_n395_), .A1(mai_mai_n61_), .B0(mai_mai_n412_), .B1(mai_mai_n162_), .Y(mai_mai_n428_));
  NOi21      m406(.An(mai_mai_n269_), .B(mai_mai_n147_), .Y(mai_mai_n429_));
  NA2        m407(.A(mai_mai_n276_), .B(mai_mai_n228_), .Y(mai_mai_n430_));
  OAI210     m408(.A0(mai_mai_n44_), .A1(x04), .B0(mai_mai_n430_), .Y(mai_mai_n431_));
  OAI210     m409(.A0(mai_mai_n431_), .A1(mai_mai_n429_), .B0(mai_mai_n100_), .Y(mai_mai_n432_));
  OAI210     m410(.A0(mai_mai_n428_), .A1(mai_mai_n90_), .B0(mai_mai_n432_), .Y(mai_mai_n433_));
  NO4        m411(.A(mai_mai_n433_), .B(mai_mai_n427_), .C(mai_mai_n419_), .D(mai_mai_n397_), .Y(mai06));
  INV        m412(.A(x07), .Y(mai_mai_n437_));
  INV        m413(.A(x07), .Y(mai_mai_n438_));
  INV        m414(.A(mai_mai_n89_), .Y(mai_mai_n439_));
  INV        m415(.A(x02), .Y(mai_mai_n440_));
  INV        m416(.A(x01), .Y(mai_mai_n441_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  AOI220     u039(.A0(x11), .A1(men_men_n48_), .B0(x10), .B1(men_men_n61_), .Y(men_men_n62_));
  INV        u040(.A(men_men_n59_), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n29_), .B(x02), .Y(men_men_n64_));
  NA2        u042(.A(men_men_n64_), .B(men_men_n24_), .Y(men_men_n65_));
  OAI220     u043(.A0(men_men_n65_), .A1(men_men_n63_), .B0(men_men_n62_), .B1(men_men_n60_), .Y(men_men_n66_));
  NA2        u044(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n67_));
  OAI210     u045(.A0(men_men_n30_), .A1(x11), .B0(men_men_n67_), .Y(men_men_n68_));
  AOI220     u046(.A0(men_men_n68_), .A1(men_men_n59_), .B0(men_men_n66_), .B1(men_men_n31_), .Y(men_men_n69_));
  AOI210     u047(.A0(men_men_n69_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n70_));
  NA2        u048(.A(x10), .B(x09), .Y(men_men_n71_));
  AOI210     u049(.A0(men_men_n71_), .A1(men_men_n61_), .B0(men_men_n23_), .Y(men_men_n72_));
  NA2        u050(.A(x09), .B(x05), .Y(men_men_n73_));
  NA2        u051(.A(x10), .B(x06), .Y(men_men_n74_));
  NA3        u052(.A(men_men_n74_), .B(men_men_n73_), .C(men_men_n28_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n76_));
  OAI210     u054(.A0(men_men_n75_), .A1(men_men_n72_), .B0(x03), .Y(men_men_n77_));
  NOi31      u055(.An(x08), .B(x04), .C(x00), .Y(men_men_n78_));
  NO2        u056(.A(x10), .B(x09), .Y(men_men_n79_));
  INV        u057(.A(men_men_n24_), .Y(men_men_n80_));
  NO2        u058(.A(x09), .B(men_men_n41_), .Y(men_men_n81_));
  NO2        u059(.A(men_men_n81_), .B(men_men_n36_), .Y(men_men_n82_));
  OAI210     u060(.A0(men_men_n81_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n83_));
  AOI210     u061(.A0(men_men_n82_), .A1(men_men_n48_), .B0(men_men_n83_), .Y(men_men_n84_));
  NO2        u062(.A(men_men_n36_), .B(x00), .Y(men_men_n85_));
  NO2        u063(.A(x08), .B(x01), .Y(men_men_n86_));
  OAI210     u064(.A0(men_men_n86_), .A1(men_men_n85_), .B0(men_men_n35_), .Y(men_men_n87_));
  NA2        u065(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n88_));
  NO3        u066(.A(men_men_n87_), .B(men_men_n84_), .C(men_men_n80_), .Y(men_men_n89_));
  AN2        u067(.A(men_men_n89_), .B(men_men_n77_), .Y(men_men_n90_));
  INV        u068(.A(men_men_n87_), .Y(men_men_n91_));
  NO2        u069(.A(x06), .B(x05), .Y(men_men_n92_));
  NA2        u070(.A(x11), .B(x00), .Y(men_men_n93_));
  NO2        u071(.A(x11), .B(men_men_n47_), .Y(men_men_n94_));
  NOi21      u072(.An(men_men_n93_), .B(men_men_n94_), .Y(men_men_n95_));
  AOI210     u073(.A0(men_men_n92_), .A1(men_men_n91_), .B0(men_men_n95_), .Y(men_men_n96_));
  NOi21      u074(.An(x01), .B(x10), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n98_));
  NO3        u076(.A(men_men_n98_), .B(men_men_n97_), .C(x06), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n99_), .B(men_men_n27_), .Y(men_men_n100_));
  OAI210     u078(.A0(men_men_n96_), .A1(x07), .B0(men_men_n100_), .Y(men_men_n101_));
  NO3        u079(.A(men_men_n101_), .B(men_men_n90_), .C(men_men_n70_), .Y(men01));
  INV        u080(.A(x12), .Y(men_men_n103_));
  INV        u081(.A(x13), .Y(men_men_n104_));
  NA2        u082(.A(men_men_n456_), .B(men_men_n71_), .Y(men_men_n105_));
  NA2        u083(.A(x08), .B(x04), .Y(men_men_n106_));
  NO2        u084(.A(men_men_n106_), .B(men_men_n57_), .Y(men_men_n107_));
  NA2        u085(.A(men_men_n107_), .B(men_men_n105_), .Y(men_men_n108_));
  NA2        u086(.A(men_men_n97_), .B(men_men_n28_), .Y(men_men_n109_));
  NO2        u087(.A(men_men_n109_), .B(men_men_n73_), .Y(men_men_n110_));
  NO2        u088(.A(x10), .B(x01), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n29_), .B(x00), .Y(men_men_n112_));
  NO2        u090(.A(men_men_n112_), .B(men_men_n111_), .Y(men_men_n113_));
  NA2        u091(.A(x04), .B(men_men_n28_), .Y(men_men_n114_));
  NO3        u092(.A(men_men_n114_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n115_));
  AOI210     u093(.A0(men_men_n115_), .A1(men_men_n113_), .B0(men_men_n110_), .Y(men_men_n116_));
  AOI210     u094(.A0(men_men_n116_), .A1(men_men_n108_), .B0(men_men_n104_), .Y(men_men_n117_));
  NO2        u095(.A(men_men_n56_), .B(x05), .Y(men_men_n118_));
  NOi21      u096(.An(men_men_n118_), .B(men_men_n58_), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n35_), .B(x02), .Y(men_men_n120_));
  NO2        u098(.A(men_men_n104_), .B(men_men_n36_), .Y(men_men_n121_));
  NA3        u099(.A(men_men_n121_), .B(men_men_n120_), .C(x06), .Y(men_men_n122_));
  NO2        u100(.A(men_men_n122_), .B(men_men_n119_), .Y(men_men_n123_));
  NO2        u101(.A(men_men_n86_), .B(x13), .Y(men_men_n124_));
  NA2        u102(.A(x13), .B(men_men_n35_), .Y(men_men_n125_));
  NO2        u103(.A(men_men_n125_), .B(x05), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n127_), .B(men_men_n104_), .Y(men_men_n128_));
  AOI210     u106(.A0(men_men_n128_), .A1(men_men_n82_), .B0(men_men_n119_), .Y(men_men_n129_));
  AOI210     u107(.A0(men_men_n129_), .A1(men_men_n124_), .B0(men_men_n74_), .Y(men_men_n130_));
  NA2        u108(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n131_));
  NA2        u109(.A(x10), .B(men_men_n57_), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n132_), .B(men_men_n131_), .Y(men_men_n133_));
  NA2        u111(.A(men_men_n51_), .B(x05), .Y(men_men_n134_));
  NO2        u112(.A(men_men_n60_), .B(x05), .Y(men_men_n135_));
  NOi41      u113(.An(men_men_n458_), .B(men_men_n135_), .C(men_men_n57_), .D(men_men_n133_), .Y(men_men_n136_));
  NO3        u114(.A(men_men_n136_), .B(x06), .C(x03), .Y(men_men_n137_));
  NO4        u115(.A(men_men_n137_), .B(men_men_n130_), .C(men_men_n123_), .D(men_men_n117_), .Y(men_men_n138_));
  NA2        u116(.A(x13), .B(men_men_n36_), .Y(men_men_n139_));
  OAI210     u117(.A0(men_men_n86_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n140_));
  NA2        u118(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n141_));
  NO2        u119(.A(men_men_n35_), .B(men_men_n47_), .Y(men_men_n142_));
  OA210      u120(.A0(x00), .A1(men_men_n79_), .B0(men_men_n142_), .Y(men_men_n143_));
  NO2        u121(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n144_));
  NA2        u122(.A(men_men_n29_), .B(x06), .Y(men_men_n145_));
  AOI210     u123(.A0(men_men_n145_), .A1(men_men_n49_), .B0(men_men_n144_), .Y(men_men_n146_));
  OA210      u124(.A0(men_men_n146_), .A1(men_men_n143_), .B0(men_men_n141_), .Y(men_men_n147_));
  NO2        u125(.A(x09), .B(x05), .Y(men_men_n148_));
  NA2        u126(.A(men_men_n148_), .B(men_men_n47_), .Y(men_men_n149_));
  AOI210     u127(.A0(men_men_n149_), .A1(men_men_n113_), .B0(men_men_n49_), .Y(men_men_n150_));
  NA2        u128(.A(x09), .B(x00), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n118_), .B(men_men_n151_), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n78_), .B(men_men_n51_), .Y(men_men_n153_));
  AOI210     u131(.A0(men_men_n153_), .A1(men_men_n152_), .B0(men_men_n145_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n154_), .B(men_men_n150_), .C(men_men_n147_), .Y(men_men_n155_));
  NO2        u133(.A(x03), .B(x02), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n87_), .B(men_men_n104_), .Y(men_men_n157_));
  OAI210     u135(.A0(men_men_n157_), .A1(men_men_n119_), .B0(men_men_n156_), .Y(men_men_n158_));
  OA210      u136(.A0(men_men_n155_), .A1(x11), .B0(men_men_n158_), .Y(men_men_n159_));
  OAI210     u137(.A0(men_men_n138_), .A1(men_men_n23_), .B0(men_men_n159_), .Y(men_men_n160_));
  NA2        u138(.A(men_men_n113_), .B(men_men_n40_), .Y(men_men_n161_));
  NA2        u139(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n162_));
  NAi21      u140(.An(x06), .B(x10), .Y(men_men_n163_));
  NOi21      u141(.An(x01), .B(x13), .Y(men_men_n164_));
  NA2        u142(.A(men_men_n164_), .B(men_men_n163_), .Y(men_men_n165_));
  OR2        u143(.A(men_men_n165_), .B(men_men_n162_), .Y(men_men_n166_));
  AOI210     u144(.A0(men_men_n166_), .A1(men_men_n161_), .B0(men_men_n41_), .Y(men_men_n167_));
  NO2        u145(.A(men_men_n29_), .B(x03), .Y(men_men_n168_));
  NA2        u146(.A(men_men_n104_), .B(x01), .Y(men_men_n169_));
  NO2        u147(.A(men_men_n169_), .B(x08), .Y(men_men_n170_));
  OAI210     u148(.A0(x05), .A1(men_men_n170_), .B0(men_men_n51_), .Y(men_men_n171_));
  AOI210     u149(.A0(men_men_n171_), .A1(men_men_n168_), .B0(men_men_n48_), .Y(men_men_n172_));
  AOI210     u150(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n173_));
  OAI210     u151(.A0(men_men_n172_), .A1(men_men_n167_), .B0(men_men_n173_), .Y(men_men_n174_));
  NA2        u152(.A(x04), .B(x02), .Y(men_men_n175_));
  NA2        u153(.A(x10), .B(x05), .Y(men_men_n176_));
  NA2        u154(.A(x09), .B(x06), .Y(men_men_n177_));
  AOI210     u155(.A0(men_men_n177_), .A1(men_men_n176_), .B0(men_men_n162_), .Y(men_men_n178_));
  NO2        u156(.A(x09), .B(x01), .Y(men_men_n179_));
  NO3        u157(.A(men_men_n179_), .B(men_men_n111_), .C(men_men_n31_), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(men_men_n178_), .B0(x00), .Y(men_men_n181_));
  NO2        u159(.A(men_men_n118_), .B(x08), .Y(men_men_n182_));
  NA3        u160(.A(men_men_n164_), .B(men_men_n163_), .C(men_men_n51_), .Y(men_men_n183_));
  NA2        u161(.A(men_men_n97_), .B(x05), .Y(men_men_n184_));
  OAI210     u162(.A0(men_men_n184_), .A1(men_men_n121_), .B0(men_men_n183_), .Y(men_men_n185_));
  AOI210     u163(.A0(men_men_n182_), .A1(x06), .B0(men_men_n185_), .Y(men_men_n186_));
  OAI210     u164(.A0(men_men_n186_), .A1(x11), .B0(men_men_n181_), .Y(men_men_n187_));
  NAi21      u165(.An(men_men_n175_), .B(men_men_n187_), .Y(men_men_n188_));
  INV        u166(.A(men_men_n25_), .Y(men_men_n189_));
  NAi21      u167(.An(x13), .B(x00), .Y(men_men_n190_));
  AOI210     u168(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n190_), .Y(men_men_n191_));
  AOI220     u169(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n192_));
  OAI210     u170(.A0(men_men_n176_), .A1(men_men_n35_), .B0(men_men_n192_), .Y(men_men_n193_));
  AN2        u171(.A(men_men_n193_), .B(men_men_n191_), .Y(men_men_n194_));
  AN2        u172(.A(men_men_n74_), .B(men_men_n73_), .Y(men_men_n195_));
  NO2        u173(.A(men_men_n98_), .B(x06), .Y(men_men_n196_));
  NO2        u174(.A(men_men_n190_), .B(men_men_n36_), .Y(men_men_n197_));
  INV        u175(.A(men_men_n197_), .Y(men_men_n198_));
  OAI220     u176(.A0(men_men_n198_), .A1(men_men_n177_), .B0(men_men_n196_), .B1(men_men_n195_), .Y(men_men_n199_));
  OAI210     u177(.A0(men_men_n199_), .A1(men_men_n194_), .B0(men_men_n189_), .Y(men_men_n200_));
  NOi21      u178(.An(x09), .B(x00), .Y(men_men_n201_));
  NO3        u179(.A(men_men_n85_), .B(men_men_n201_), .C(men_men_n47_), .Y(men_men_n202_));
  NA2        u180(.A(men_men_n202_), .B(men_men_n132_), .Y(men_men_n203_));
  NA2        u181(.A(x10), .B(x08), .Y(men_men_n204_));
  INV        u182(.A(men_men_n204_), .Y(men_men_n205_));
  NA2        u183(.A(x06), .B(x05), .Y(men_men_n206_));
  OAI210     u184(.A0(men_men_n206_), .A1(men_men_n35_), .B0(men_men_n103_), .Y(men_men_n207_));
  AOI210     u185(.A0(men_men_n205_), .A1(men_men_n58_), .B0(men_men_n207_), .Y(men_men_n208_));
  NA2        u186(.A(men_men_n208_), .B(men_men_n203_), .Y(men_men_n209_));
  NO2        u187(.A(men_men_n104_), .B(x12), .Y(men_men_n210_));
  AOI210     u188(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n210_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n97_), .B(men_men_n51_), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n213_));
  NA2        u191(.A(men_men_n213_), .B(x02), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n214_), .B(men_men_n212_), .Y(men_men_n215_));
  AOI210     u193(.A0(men_men_n211_), .A1(men_men_n209_), .B0(men_men_n215_), .Y(men_men_n216_));
  NA4        u194(.A(men_men_n216_), .B(men_men_n200_), .C(men_men_n188_), .D(men_men_n174_), .Y(men_men_n217_));
  AOI210     u195(.A0(men_men_n160_), .A1(men_men_n103_), .B0(men_men_n217_), .Y(men_men_n218_));
  INV        u196(.A(men_men_n75_), .Y(men_men_n219_));
  NA2        u197(.A(men_men_n219_), .B(men_men_n141_), .Y(men_men_n220_));
  NA2        u198(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n221_));
  NA2        u199(.A(men_men_n221_), .B(men_men_n140_), .Y(men_men_n222_));
  NO2        u200(.A(men_men_n131_), .B(x06), .Y(men_men_n223_));
  INV        u201(.A(men_men_n223_), .Y(men_men_n224_));
  AOI210     u202(.A0(men_men_n224_), .A1(men_men_n220_), .B0(x12), .Y(men_men_n225_));
  INV        u203(.A(men_men_n78_), .Y(men_men_n226_));
  NA2        u204(.A(men_men_n165_), .B(men_men_n57_), .Y(men_men_n227_));
  NA2        u205(.A(men_men_n227_), .B(men_men_n226_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n97_), .B(x06), .Y(men_men_n229_));
  AOI210     u207(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n230_));
  NO3        u208(.A(men_men_n230_), .B(men_men_n229_), .C(men_men_n41_), .Y(men_men_n231_));
  NA4        u209(.A(men_men_n163_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n232_), .B(men_men_n145_), .Y(men_men_n233_));
  OAI210     u211(.A0(men_men_n233_), .A1(men_men_n231_), .B0(x02), .Y(men_men_n234_));
  AOI210     u212(.A0(men_men_n234_), .A1(men_men_n228_), .B0(men_men_n23_), .Y(men_men_n235_));
  OAI210     u213(.A0(men_men_n225_), .A1(men_men_n57_), .B0(men_men_n235_), .Y(men_men_n236_));
  INV        u214(.A(men_men_n145_), .Y(men_men_n237_));
  NO2        u215(.A(men_men_n51_), .B(x03), .Y(men_men_n238_));
  NO2        u216(.A(men_men_n104_), .B(x03), .Y(men_men_n239_));
  INV        u217(.A(men_men_n163_), .Y(men_men_n240_));
  NOi21      u218(.An(x13), .B(x04), .Y(men_men_n241_));
  NO3        u219(.A(men_men_n241_), .B(men_men_n78_), .C(men_men_n201_), .Y(men_men_n242_));
  NO2        u220(.A(men_men_n242_), .B(x05), .Y(men_men_n243_));
  AOI220     u221(.A0(men_men_n243_), .A1(men_men_n460_), .B0(men_men_n240_), .B1(men_men_n57_), .Y(men_men_n244_));
  INV        u222(.A(men_men_n244_), .Y(men_men_n245_));
  INV        u223(.A(men_men_n94_), .Y(men_men_n246_));
  NO2        u224(.A(men_men_n246_), .B(x12), .Y(men_men_n247_));
  NA2        u225(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n248_));
  NO2        u226(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n249_));
  OAI210     u227(.A0(men_men_n249_), .A1(men_men_n193_), .B0(men_men_n191_), .Y(men_men_n250_));
  AOI210     u228(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n251_));
  NO2        u229(.A(men_men_n251_), .B(men_men_n41_), .Y(men_men_n252_));
  OAI210     u230(.A0(men_men_n106_), .A1(men_men_n151_), .B0(men_men_n74_), .Y(men_men_n253_));
  NO2        u231(.A(men_men_n253_), .B(men_men_n252_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n255_));
  NA2        u233(.A(men_men_n255_), .B(x03), .Y(men_men_n256_));
  OA210      u234(.A0(men_men_n256_), .A1(men_men_n254_), .B0(men_men_n250_), .Y(men_men_n257_));
  NA2        u235(.A(x13), .B(men_men_n103_), .Y(men_men_n258_));
  NA3        u236(.A(men_men_n258_), .B(men_men_n207_), .C(men_men_n95_), .Y(men_men_n259_));
  OAI210     u237(.A0(men_men_n257_), .A1(men_men_n248_), .B0(men_men_n259_), .Y(men_men_n260_));
  AOI210     u238(.A0(men_men_n247_), .A1(men_men_n245_), .B0(men_men_n260_), .Y(men_men_n261_));
  AOI210     u239(.A0(men_men_n261_), .A1(men_men_n236_), .B0(x07), .Y(men_men_n262_));
  NA2        u240(.A(men_men_n73_), .B(men_men_n29_), .Y(men_men_n263_));
  NOi31      u241(.An(men_men_n139_), .B(men_men_n241_), .C(men_men_n201_), .Y(men_men_n264_));
  AOI210     u242(.A0(men_men_n264_), .A1(men_men_n153_), .B0(men_men_n263_), .Y(men_men_n265_));
  NO2        u243(.A(men_men_n104_), .B(x06), .Y(men_men_n266_));
  INV        u244(.A(men_men_n266_), .Y(men_men_n267_));
  NO2        u245(.A(x08), .B(x05), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n268_), .B(men_men_n251_), .Y(men_men_n269_));
  OAI210     u247(.A0(men_men_n78_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n270_));
  OAI210     u248(.A0(men_men_n269_), .A1(men_men_n267_), .B0(men_men_n270_), .Y(men_men_n271_));
  NO2        u249(.A(x12), .B(x02), .Y(men_men_n272_));
  INV        u250(.A(men_men_n272_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n273_), .B(men_men_n246_), .Y(men_men_n274_));
  OA210      u252(.A0(men_men_n271_), .A1(men_men_n265_), .B0(men_men_n274_), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n276_));
  NO2        u254(.A(men_men_n276_), .B(x01), .Y(men_men_n277_));
  AOI210     u255(.A0(men_men_n459_), .A1(men_men_n458_), .B0(men_men_n29_), .Y(men_men_n278_));
  NA2        u256(.A(men_men_n104_), .B(x04), .Y(men_men_n279_));
  OAI210     u257(.A0(x02), .A1(men_men_n124_), .B0(men_men_n457_), .Y(men_men_n280_));
  NO3        u258(.A(men_men_n93_), .B(x12), .C(x03), .Y(men_men_n281_));
  OAI210     u259(.A0(men_men_n280_), .A1(men_men_n278_), .B0(men_men_n281_), .Y(men_men_n282_));
  AOI210     u260(.A0(men_men_n212_), .A1(men_men_n206_), .B0(men_men_n106_), .Y(men_men_n283_));
  NOi21      u261(.An(men_men_n263_), .B(men_men_n229_), .Y(men_men_n284_));
  NO2        u262(.A(men_men_n25_), .B(x00), .Y(men_men_n285_));
  OAI210     u263(.A0(men_men_n284_), .A1(men_men_n283_), .B0(men_men_n285_), .Y(men_men_n286_));
  NO2        u264(.A(men_men_n58_), .B(x05), .Y(men_men_n287_));
  NO3        u265(.A(men_men_n287_), .B(men_men_n230_), .C(men_men_n196_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n248_), .B(men_men_n28_), .Y(men_men_n289_));
  OAI210     u267(.A0(men_men_n288_), .A1(men_men_n237_), .B0(men_men_n289_), .Y(men_men_n290_));
  NA3        u268(.A(men_men_n290_), .B(men_men_n286_), .C(men_men_n282_), .Y(men_men_n291_));
  NO3        u269(.A(men_men_n291_), .B(men_men_n275_), .C(men_men_n262_), .Y(men_men_n292_));
  OAI210     u270(.A0(men_men_n218_), .A1(men_men_n61_), .B0(men_men_n292_), .Y(men02));
  AOI210     u271(.A0(men_men_n139_), .A1(men_men_n87_), .B0(men_men_n134_), .Y(men_men_n294_));
  NOi21      u272(.An(men_men_n242_), .B(men_men_n179_), .Y(men_men_n295_));
  NO2        u273(.A(men_men_n104_), .B(men_men_n35_), .Y(men_men_n296_));
  NA3        u274(.A(men_men_n296_), .B(men_men_n205_), .C(men_men_n56_), .Y(men_men_n297_));
  OAI210     u275(.A0(men_men_n295_), .A1(men_men_n32_), .B0(men_men_n297_), .Y(men_men_n298_));
  OAI210     u276(.A0(men_men_n298_), .A1(men_men_n294_), .B0(men_men_n176_), .Y(men_men_n299_));
  INV        u277(.A(men_men_n176_), .Y(men_men_n300_));
  AOI210     u278(.A0(men_men_n120_), .A1(men_men_n88_), .B0(men_men_n230_), .Y(men_men_n301_));
  OAI220     u279(.A0(men_men_n301_), .A1(men_men_n104_), .B0(men_men_n87_), .B1(men_men_n51_), .Y(men_men_n302_));
  AOI220     u280(.A0(men_men_n302_), .A1(men_men_n300_), .B0(men_men_n157_), .B1(men_men_n156_), .Y(men_men_n303_));
  AOI210     u281(.A0(men_men_n303_), .A1(men_men_n299_), .B0(men_men_n48_), .Y(men_men_n304_));
  NO2        u282(.A(x05), .B(x02), .Y(men_men_n305_));
  OAI210     u283(.A0(men_men_n222_), .A1(men_men_n201_), .B0(men_men_n305_), .Y(men_men_n306_));
  AOI220     u284(.A0(men_men_n268_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n307_));
  NOi21      u285(.An(men_men_n296_), .B(men_men_n307_), .Y(men_men_n308_));
  AOI210     u286(.A0(men_men_n241_), .A1(men_men_n81_), .B0(men_men_n308_), .Y(men_men_n309_));
  AOI210     u287(.A0(men_men_n309_), .A1(men_men_n306_), .B0(men_men_n145_), .Y(men_men_n310_));
  NO2        u288(.A(men_men_n255_), .B(men_men_n47_), .Y(men_men_n311_));
  NA2        u289(.A(men_men_n311_), .B(men_men_n243_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n313_));
  NA2        u291(.A(x13), .B(men_men_n28_), .Y(men_men_n314_));
  OA210      u292(.A0(men_men_n314_), .A1(x08), .B0(men_men_n149_), .Y(men_men_n315_));
  AOI210     u293(.A0(men_men_n315_), .A1(men_men_n140_), .B0(men_men_n313_), .Y(men_men_n316_));
  NA2        u294(.A(men_men_n316_), .B(men_men_n98_), .Y(men_men_n317_));
  NA3        u295(.A(men_men_n98_), .B(men_men_n86_), .C(men_men_n238_), .Y(men_men_n318_));
  NA3        u296(.A(men_men_n97_), .B(men_men_n85_), .C(men_men_n42_), .Y(men_men_n319_));
  AOI210     u297(.A0(men_men_n319_), .A1(men_men_n318_), .B0(x04), .Y(men_men_n320_));
  INV        u298(.A(men_men_n156_), .Y(men_men_n321_));
  OAI220     u299(.A0(men_men_n269_), .A1(men_men_n109_), .B0(men_men_n321_), .B1(men_men_n133_), .Y(men_men_n322_));
  AOI210     u300(.A0(men_men_n322_), .A1(x13), .B0(men_men_n320_), .Y(men_men_n323_));
  NA3        u301(.A(men_men_n323_), .B(men_men_n317_), .C(men_men_n312_), .Y(men_men_n324_));
  NO3        u302(.A(men_men_n324_), .B(men_men_n310_), .C(men_men_n304_), .Y(men_men_n325_));
  NA2        u303(.A(men_men_n144_), .B(x03), .Y(men_men_n326_));
  OAI210     u304(.A0(men_men_n190_), .A1(men_men_n287_), .B0(men_men_n326_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n327_), .B(men_men_n111_), .Y(men_men_n328_));
  INV        u306(.A(men_men_n56_), .Y(men_men_n329_));
  OAI220     u307(.A0(men_men_n279_), .A1(men_men_n329_), .B0(men_men_n134_), .B1(men_men_n28_), .Y(men_men_n330_));
  NA2        u308(.A(men_men_n330_), .B(men_men_n112_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n279_), .B(men_men_n103_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n103_), .B(men_men_n41_), .Y(men_men_n333_));
  NA3        u311(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n133_), .Y(men_men_n334_));
  NA4        u312(.A(men_men_n334_), .B(men_men_n331_), .C(men_men_n328_), .D(men_men_n48_), .Y(men_men_n335_));
  INV        u313(.A(men_men_n213_), .Y(men_men_n336_));
  NO2        u314(.A(men_men_n170_), .B(men_men_n40_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n32_), .B(x05), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n337_), .B0(men_men_n336_), .B1(men_men_n59_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n339_), .B(x02), .Y(men_men_n340_));
  INV        u318(.A(men_men_n249_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n210_), .B(x04), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  NO3        u321(.A(men_men_n192_), .B(x13), .C(men_men_n31_), .Y(men_men_n344_));
  OAI210     u322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n98_), .Y(men_men_n345_));
  NO3        u323(.A(men_men_n210_), .B(men_men_n168_), .C(men_men_n52_), .Y(men_men_n346_));
  OAI210     u324(.A0(x12), .A1(men_men_n202_), .B0(men_men_n346_), .Y(men_men_n347_));
  NA4        u325(.A(men_men_n347_), .B(men_men_n345_), .C(men_men_n340_), .D(x06), .Y(men_men_n348_));
  NA2        u326(.A(x09), .B(x03), .Y(men_men_n349_));
  OAI220     u327(.A0(men_men_n349_), .A1(men_men_n132_), .B0(men_men_n221_), .B1(men_men_n64_), .Y(men_men_n350_));
  OAI220     u328(.A0(men_men_n169_), .A1(x09), .B0(x08), .B1(men_men_n41_), .Y(men_men_n351_));
  NO3        u329(.A(men_men_n287_), .B(men_men_n131_), .C(x08), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n351_), .A1(men_men_n237_), .B0(men_men_n352_), .Y(men_men_n353_));
  NO2        u331(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n354_));
  NO3        u332(.A(men_men_n118_), .B(men_men_n132_), .C(men_men_n38_), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n346_), .A1(men_men_n354_), .B0(men_men_n355_), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n353_), .A1(men_men_n28_), .B0(men_men_n356_), .Y(men_men_n357_));
  AO220      u335(.A0(men_men_n357_), .A1(x04), .B0(men_men_n350_), .B1(x05), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n348_), .A1(men_men_n335_), .B0(men_men_n358_), .Y(men_men_n359_));
  OAI210     u337(.A0(men_men_n325_), .A1(x12), .B0(men_men_n359_), .Y(men03));
  OR2        u338(.A(men_men_n42_), .B(men_men_n238_), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n157_), .A1(men_men_n103_), .B0(men_men_n361_), .Y(men_men_n362_));
  AO210      u340(.A0(men_men_n341_), .A1(men_men_n88_), .B0(men_men_n342_), .Y(men_men_n363_));
  NA2        u341(.A(men_men_n210_), .B(men_men_n156_), .Y(men_men_n364_));
  NA3        u342(.A(men_men_n364_), .B(men_men_n363_), .C(men_men_n214_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n362_), .B0(x05), .Y(men_men_n366_));
  NA2        u344(.A(men_men_n361_), .B(x05), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n140_), .A1(men_men_n226_), .B0(men_men_n367_), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n239_), .A1(men_men_n82_), .B0(men_men_n126_), .Y(men_men_n369_));
  OAI220     u347(.A0(men_men_n369_), .A1(men_men_n59_), .B0(men_men_n314_), .B1(men_men_n307_), .Y(men_men_n370_));
  OAI210     u348(.A0(men_men_n370_), .A1(men_men_n368_), .B0(men_men_n103_), .Y(men_men_n371_));
  AOI210     u349(.A0(men_men_n149_), .A1(men_men_n60_), .B0(men_men_n38_), .Y(men_men_n372_));
  NO2        u350(.A(men_men_n179_), .B(men_men_n135_), .Y(men_men_n373_));
  OAI220     u351(.A0(men_men_n373_), .A1(men_men_n37_), .B0(men_men_n152_), .B1(x13), .Y(men_men_n374_));
  OAI210     u352(.A0(men_men_n374_), .A1(men_men_n372_), .B0(x04), .Y(men_men_n375_));
  NO3        u353(.A(men_men_n333_), .B(men_men_n87_), .C(men_men_n59_), .Y(men_men_n376_));
  AOI210     u354(.A0(men_men_n198_), .A1(men_men_n103_), .B0(men_men_n149_), .Y(men_men_n377_));
  OA210      u355(.A0(men_men_n170_), .A1(x12), .B0(men_men_n135_), .Y(men_men_n378_));
  NO3        u356(.A(men_men_n378_), .B(men_men_n377_), .C(men_men_n376_), .Y(men_men_n379_));
  NA4        u357(.A(men_men_n379_), .B(men_men_n375_), .C(men_men_n371_), .D(men_men_n366_), .Y(men04));
  NO2        u358(.A(men_men_n91_), .B(men_men_n39_), .Y(men_men_n381_));
  XO2        u359(.A(men_men_n381_), .B(men_men_n258_), .Y(men05));
  AOI210     u360(.A0(men_men_n73_), .A1(men_men_n52_), .B0(men_men_n223_), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n383_), .A1(men_men_n313_), .B0(men_men_n25_), .Y(men_men_n384_));
  NAi41      u362(.An(men_men_n79_), .B(men_men_n145_), .C(men_men_n134_), .D(men_men_n31_), .Y(men_men_n385_));
  AOI210     u363(.A0(men_men_n240_), .A1(men_men_n57_), .B0(men_men_n92_), .Y(men_men_n386_));
  AOI210     u364(.A0(men_men_n386_), .A1(men_men_n385_), .B0(men_men_n24_), .Y(men_men_n387_));
  OAI210     u365(.A0(men_men_n387_), .A1(men_men_n384_), .B0(men_men_n103_), .Y(men_men_n388_));
  NA2        u366(.A(x11), .B(men_men_n31_), .Y(men_men_n389_));
  NA2        u367(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n390_));
  NA2        u368(.A(men_men_n263_), .B(x03), .Y(men_men_n391_));
  OAI220     u369(.A0(men_men_n391_), .A1(men_men_n390_), .B0(men_men_n389_), .B1(men_men_n83_), .Y(men_men_n392_));
  OAI210     u370(.A0(men_men_n26_), .A1(men_men_n103_), .B0(x07), .Y(men_men_n393_));
  AOI210     u371(.A0(men_men_n392_), .A1(x06), .B0(men_men_n393_), .Y(men_men_n394_));
  AOI220     u372(.A0(men_men_n83_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n395_));
  NO3        u373(.A(men_men_n395_), .B(men_men_n23_), .C(x00), .Y(men_men_n396_));
  NA2        u374(.A(men_men_n71_), .B(x02), .Y(men_men_n397_));
  AOI210     u375(.A0(men_men_n397_), .A1(men_men_n391_), .B0(men_men_n266_), .Y(men_men_n398_));
  OR2        u376(.A(men_men_n398_), .B(men_men_n248_), .Y(men_men_n399_));
  NO2        u377(.A(men_men_n23_), .B(x10), .Y(men_men_n400_));
  OAI210     u378(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n401_));
  OR3        u379(.A(men_men_n401_), .B(men_men_n400_), .C(men_men_n44_), .Y(men_men_n402_));
  NA2        u380(.A(men_men_n402_), .B(men_men_n399_), .Y(men_men_n403_));
  OAI210     u381(.A0(men_men_n403_), .A1(men_men_n396_), .B0(men_men_n103_), .Y(men_men_n404_));
  NA2        u382(.A(men_men_n33_), .B(men_men_n103_), .Y(men_men_n405_));
  AOI210     u383(.A0(men_men_n405_), .A1(men_men_n94_), .B0(x07), .Y(men_men_n406_));
  AOI220     u384(.A0(men_men_n406_), .A1(men_men_n404_), .B0(men_men_n394_), .B1(men_men_n388_), .Y(men_men_n407_));
  NA3        u385(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n408_));
  AO210      u386(.A0(men_men_n408_), .A1(men_men_n276_), .B0(men_men_n273_), .Y(men_men_n409_));
  AOI210     u387(.A0(men_men_n400_), .A1(men_men_n76_), .B0(men_men_n144_), .Y(men_men_n410_));
  OR2        u388(.A(men_men_n410_), .B(x03), .Y(men_men_n411_));
  NA2        u389(.A(men_men_n354_), .B(men_men_n61_), .Y(men_men_n412_));
  NO2        u390(.A(men_men_n412_), .B(x11), .Y(men_men_n413_));
  NO3        u391(.A(men_men_n413_), .B(men_men_n148_), .C(men_men_n28_), .Y(men_men_n414_));
  AOI220     u392(.A0(men_men_n414_), .A1(men_men_n411_), .B0(men_men_n409_), .B1(men_men_n47_), .Y(men_men_n415_));
  NO4        u393(.A(men_men_n333_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n416_));
  OAI210     u394(.A0(men_men_n416_), .A1(men_men_n415_), .B0(men_men_n104_), .Y(men_men_n417_));
  AOI210     u395(.A0(men_men_n342_), .A1(men_men_n114_), .B0(men_men_n272_), .Y(men_men_n418_));
  NOi21      u396(.An(men_men_n326_), .B(men_men_n135_), .Y(men_men_n419_));
  NO2        u397(.A(men_men_n419_), .B(men_men_n273_), .Y(men_men_n420_));
  OAI210     u398(.A0(x12), .A1(men_men_n47_), .B0(men_men_n35_), .Y(men_men_n421_));
  AOI210     u399(.A0(men_men_n258_), .A1(men_men_n47_), .B0(men_men_n421_), .Y(men_men_n422_));
  NO4        u400(.A(men_men_n422_), .B(men_men_n420_), .C(men_men_n418_), .D(x08), .Y(men_men_n423_));
  AOI210     u401(.A0(men_men_n400_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n424_));
  NA2        u402(.A(x09), .B(men_men_n41_), .Y(men_men_n425_));
  OAI220     u403(.A0(men_men_n425_), .A1(men_men_n424_), .B0(men_men_n389_), .B1(men_men_n67_), .Y(men_men_n426_));
  NO2        u404(.A(x13), .B(x12), .Y(men_men_n427_));
  NO2        u405(.A(men_men_n134_), .B(men_men_n28_), .Y(men_men_n428_));
  NO2        u406(.A(men_men_n428_), .B(men_men_n277_), .Y(men_men_n429_));
  NA3        u407(.A(men_men_n336_), .B(men_men_n127_), .C(x12), .Y(men_men_n430_));
  AO210      u408(.A0(men_men_n336_), .A1(men_men_n127_), .B0(men_men_n258_), .Y(men_men_n431_));
  NA3        u409(.A(men_men_n431_), .B(men_men_n430_), .C(x08), .Y(men_men_n432_));
  AOI210     u410(.A0(men_men_n427_), .A1(men_men_n426_), .B0(men_men_n432_), .Y(men_men_n433_));
  AOI210     u411(.A0(men_men_n423_), .A1(men_men_n417_), .B0(men_men_n433_), .Y(men_men_n434_));
  OAI210     u412(.A0(men_men_n412_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n435_));
  NA2        u413(.A(men_men_n300_), .B(x07), .Y(men_men_n436_));
  OAI220     u414(.A0(men_men_n436_), .A1(men_men_n390_), .B0(men_men_n148_), .B1(men_men_n43_), .Y(men_men_n437_));
  OAI210     u415(.A0(men_men_n437_), .A1(men_men_n435_), .B0(men_men_n197_), .Y(men_men_n438_));
  NA3        u416(.A(men_men_n429_), .B(men_men_n419_), .C(men_men_n332_), .Y(men_men_n439_));
  INV        u417(.A(x14), .Y(men_men_n440_));
  NO3        u418(.A(men_men_n326_), .B(men_men_n109_), .C(x11), .Y(men_men_n441_));
  NO3        u419(.A(men_men_n169_), .B(men_men_n76_), .C(men_men_n57_), .Y(men_men_n442_));
  NO3        u420(.A(men_men_n408_), .B(men_men_n333_), .C(men_men_n190_), .Y(men_men_n443_));
  NO4        u421(.A(men_men_n443_), .B(men_men_n442_), .C(men_men_n441_), .D(men_men_n440_), .Y(men_men_n444_));
  NA3        u422(.A(men_men_n444_), .B(men_men_n439_), .C(men_men_n438_), .Y(men_men_n445_));
  AOI220     u423(.A0(men_men_n405_), .A1(men_men_n61_), .B0(men_men_n428_), .B1(men_men_n168_), .Y(men_men_n446_));
  NOi21      u424(.An(men_men_n279_), .B(men_men_n152_), .Y(men_men_n447_));
  NO3        u425(.A(men_men_n131_), .B(men_men_n24_), .C(x06), .Y(men_men_n448_));
  AOI210     u426(.A0(men_men_n285_), .A1(men_men_n240_), .B0(men_men_n448_), .Y(men_men_n449_));
  OAI210     u427(.A0(men_men_n44_), .A1(x04), .B0(men_men_n449_), .Y(men_men_n450_));
  OAI210     u428(.A0(men_men_n450_), .A1(men_men_n447_), .B0(men_men_n103_), .Y(men_men_n451_));
  OAI210     u429(.A0(men_men_n446_), .A1(men_men_n93_), .B0(men_men_n451_), .Y(men_men_n452_));
  NO4        u430(.A(men_men_n452_), .B(men_men_n445_), .C(men_men_n434_), .D(men_men_n407_), .Y(men06));
  INV        u431(.A(x01), .Y(men_men_n456_));
  INV        u432(.A(men_men_n266_), .Y(men_men_n457_));
  INV        u433(.A(x13), .Y(men_men_n458_));
  INV        u434(.A(men_men_n86_), .Y(men_men_n459_));
  INV        u435(.A(x06), .Y(men_men_n460_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule