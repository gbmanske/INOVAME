library verilog;
use verilog.vl_types.all;
entity cla_16bits_vlg_vec_tst is
end cla_16bits_vlg_vec_tst;
