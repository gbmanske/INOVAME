//Benchmark atmr_misex3_1774_0.0156

module atmr_misex3(a, b, c, d, e, f, g, h, i, j, k, l, m, n, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13);
 input a, b, c, d, e, f, g, h, i, j, k, l, m, n;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13;
 wire ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n550_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n693_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n742_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n791_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n958_, ori_ori_n959_, ori_ori_n960_, ori_ori_n961_, ori_ori_n962_, ori_ori_n963_, ori_ori_n964_, ori_ori_n965_, ori_ori_n966_, ori_ori_n967_, ori_ori_n968_, ori_ori_n969_, ori_ori_n970_, ori_ori_n971_, ori_ori_n972_, ori_ori_n973_, ori_ori_n974_, ori_ori_n975_, ori_ori_n976_, ori_ori_n977_, ori_ori_n978_, ori_ori_n979_, ori_ori_n980_, ori_ori_n981_, ori_ori_n982_, ori_ori_n983_, ori_ori_n984_, ori_ori_n985_, ori_ori_n986_, ori_ori_n987_, ori_ori_n988_, ori_ori_n989_, ori_ori_n990_, ori_ori_n991_, ori_ori_n992_, ori_ori_n993_, ori_ori_n994_, ori_ori_n995_, ori_ori_n996_, ori_ori_n997_, ori_ori_n998_, ori_ori_n999_, ori_ori_n1000_, ori_ori_n1001_, ori_ori_n1002_, ori_ori_n1003_, ori_ori_n1004_, ori_ori_n1005_, ori_ori_n1006_, ori_ori_n1007_, ori_ori_n1008_, ori_ori_n1009_, ori_ori_n1010_, ori_ori_n1011_, ori_ori_n1012_, ori_ori_n1013_, ori_ori_n1014_, ori_ori_n1015_, ori_ori_n1016_, ori_ori_n1017_, ori_ori_n1018_, ori_ori_n1019_, ori_ori_n1020_, ori_ori_n1021_, ori_ori_n1022_, ori_ori_n1023_, ori_ori_n1024_, ori_ori_n1025_, ori_ori_n1026_, ori_ori_n1027_, ori_ori_n1028_, ori_ori_n1029_, ori_ori_n1030_, ori_ori_n1031_, ori_ori_n1032_, ori_ori_n1033_, ori_ori_n1034_, ori_ori_n1035_, ori_ori_n1036_, ori_ori_n1037_, ori_ori_n1038_, ori_ori_n1039_, ori_ori_n1040_, ori_ori_n1041_, ori_ori_n1043_, ori_ori_n1044_, ori_ori_n1045_, ori_ori_n1046_, ori_ori_n1047_, ori_ori_n1048_, ori_ori_n1049_, ori_ori_n1050_, ori_ori_n1051_, ori_ori_n1052_, ori_ori_n1053_, ori_ori_n1054_, ori_ori_n1055_, ori_ori_n1056_, ori_ori_n1057_, ori_ori_n1058_, ori_ori_n1059_, ori_ori_n1060_, ori_ori_n1062_, ori_ori_n1063_, ori_ori_n1064_, ori_ori_n1065_, ori_ori_n1066_, ori_ori_n1067_, ori_ori_n1068_, ori_ori_n1069_, ori_ori_n1070_, ori_ori_n1071_, ori_ori_n1072_, ori_ori_n1074_, ori_ori_n1075_, ori_ori_n1076_, ori_ori_n1077_, ori_ori_n1078_, ori_ori_n1079_, ori_ori_n1080_, ori_ori_n1081_, ori_ori_n1082_, ori_ori_n1083_, ori_ori_n1084_, ori_ori_n1085_, ori_ori_n1086_, ori_ori_n1087_, ori_ori_n1088_, ori_ori_n1089_, ori_ori_n1090_, ori_ori_n1091_, ori_ori_n1092_, ori_ori_n1093_, ori_ori_n1094_, ori_ori_n1095_, ori_ori_n1096_, ori_ori_n1097_, ori_ori_n1098_, ori_ori_n1099_, ori_ori_n1100_, ori_ori_n1101_, ori_ori_n1102_, ori_ori_n1103_, ori_ori_n1104_, ori_ori_n1105_, ori_ori_n1106_, ori_ori_n1107_, ori_ori_n1108_, ori_ori_n1109_, ori_ori_n1110_, ori_ori_n1111_, ori_ori_n1112_, ori_ori_n1113_, ori_ori_n1114_, ori_ori_n1115_, ori_ori_n1116_, ori_ori_n1117_, ori_ori_n1118_, ori_ori_n1119_, ori_ori_n1120_, ori_ori_n1121_, ori_ori_n1123_, ori_ori_n1124_, ori_ori_n1125_, ori_ori_n1126_, ori_ori_n1127_, ori_ori_n1128_, ori_ori_n1129_, ori_ori_n1130_, ori_ori_n1131_, ori_ori_n1132_, ori_ori_n1133_, ori_ori_n1134_, ori_ori_n1135_, ori_ori_n1136_, ori_ori_n1137_, ori_ori_n1138_, ori_ori_n1139_, ori_ori_n1140_, ori_ori_n1141_, ori_ori_n1142_, ori_ori_n1143_, ori_ori_n1144_, ori_ori_n1145_, ori_ori_n1146_, ori_ori_n1147_, ori_ori_n1148_, ori_ori_n1149_, ori_ori_n1150_, ori_ori_n1151_, ori_ori_n1152_, ori_ori_n1153_, ori_ori_n1154_, ori_ori_n1155_, ori_ori_n1156_, ori_ori_n1157_, ori_ori_n1158_, ori_ori_n1159_, ori_ori_n1160_, ori_ori_n1161_, ori_ori_n1162_, ori_ori_n1163_, ori_ori_n1164_, ori_ori_n1165_, ori_ori_n1166_, ori_ori_n1167_, ori_ori_n1168_, ori_ori_n1169_, ori_ori_n1170_, ori_ori_n1171_, ori_ori_n1173_, ori_ori_n1174_, ori_ori_n1175_, ori_ori_n1176_, ori_ori_n1177_, ori_ori_n1178_, ori_ori_n1179_, ori_ori_n1180_, ori_ori_n1181_, ori_ori_n1182_, ori_ori_n1183_, ori_ori_n1184_, ori_ori_n1185_, ori_ori_n1186_, ori_ori_n1187_, ori_ori_n1188_, ori_ori_n1189_, ori_ori_n1190_, ori_ori_n1191_, ori_ori_n1192_, ori_ori_n1193_, ori_ori_n1194_, ori_ori_n1195_, ori_ori_n1196_, ori_ori_n1197_, ori_ori_n1198_, ori_ori_n1199_, ori_ori_n1200_, ori_ori_n1201_, ori_ori_n1202_, ori_ori_n1203_, ori_ori_n1204_, ori_ori_n1205_, ori_ori_n1206_, ori_ori_n1207_, ori_ori_n1208_, ori_ori_n1209_, ori_ori_n1210_, ori_ori_n1211_, ori_ori_n1212_, ori_ori_n1213_, ori_ori_n1214_, ori_ori_n1215_, ori_ori_n1216_, ori_ori_n1217_, ori_ori_n1218_, ori_ori_n1219_, ori_ori_n1220_, ori_ori_n1221_, ori_ori_n1222_, ori_ori_n1223_, ori_ori_n1224_, ori_ori_n1225_, ori_ori_n1226_, ori_ori_n1227_, ori_ori_n1228_, ori_ori_n1229_, ori_ori_n1230_, ori_ori_n1231_, ori_ori_n1232_, ori_ori_n1233_, ori_ori_n1234_, ori_ori_n1235_, ori_ori_n1236_, ori_ori_n1237_, ori_ori_n1238_, ori_ori_n1239_, ori_ori_n1240_, ori_ori_n1241_, ori_ori_n1242_, ori_ori_n1243_, ori_ori_n1245_, ori_ori_n1246_, ori_ori_n1247_, ori_ori_n1248_, ori_ori_n1249_, ori_ori_n1250_, ori_ori_n1251_, ori_ori_n1252_, ori_ori_n1253_, ori_ori_n1254_, ori_ori_n1255_, ori_ori_n1256_, ori_ori_n1257_, ori_ori_n1258_, ori_ori_n1259_, ori_ori_n1260_, ori_ori_n1261_, ori_ori_n1262_, ori_ori_n1263_, ori_ori_n1264_, ori_ori_n1265_, ori_ori_n1266_, ori_ori_n1267_, ori_ori_n1268_, ori_ori_n1269_, ori_ori_n1270_, ori_ori_n1271_, ori_ori_n1272_, ori_ori_n1273_, ori_ori_n1274_, ori_ori_n1275_, ori_ori_n1276_, ori_ori_n1277_, ori_ori_n1278_, ori_ori_n1279_, ori_ori_n1280_, ori_ori_n1281_, ori_ori_n1282_, ori_ori_n1283_, ori_ori_n1284_, ori_ori_n1285_, ori_ori_n1286_, ori_ori_n1288_, ori_ori_n1289_, ori_ori_n1290_, ori_ori_n1291_, ori_ori_n1292_, ori_ori_n1293_, ori_ori_n1294_, ori_ori_n1295_, ori_ori_n1296_, ori_ori_n1297_, ori_ori_n1298_, ori_ori_n1299_, ori_ori_n1300_, ori_ori_n1301_, ori_ori_n1302_, ori_ori_n1303_, ori_ori_n1304_, ori_ori_n1305_, ori_ori_n1306_, ori_ori_n1307_, ori_ori_n1308_, ori_ori_n1309_, ori_ori_n1310_, ori_ori_n1311_, ori_ori_n1312_, ori_ori_n1313_, ori_ori_n1314_, ori_ori_n1315_, ori_ori_n1316_, ori_ori_n1317_, ori_ori_n1318_, ori_ori_n1319_, ori_ori_n1320_, ori_ori_n1321_, ori_ori_n1322_, ori_ori_n1323_, ori_ori_n1324_, ori_ori_n1325_, ori_ori_n1326_, ori_ori_n1327_, ori_ori_n1328_, ori_ori_n1329_, ori_ori_n1330_, ori_ori_n1331_, ori_ori_n1332_, ori_ori_n1333_, ori_ori_n1334_, ori_ori_n1335_, ori_ori_n1336_, ori_ori_n1337_, ori_ori_n1338_, ori_ori_n1339_, ori_ori_n1340_, ori_ori_n1341_, ori_ori_n1342_, ori_ori_n1343_, ori_ori_n1344_, ori_ori_n1345_, ori_ori_n1346_, ori_ori_n1347_, ori_ori_n1348_, ori_ori_n1349_, ori_ori_n1350_, ori_ori_n1351_, ori_ori_n1352_, ori_ori_n1353_, ori_ori_n1354_, ori_ori_n1355_, ori_ori_n1356_, ori_ori_n1357_, ori_ori_n1358_, ori_ori_n1359_, ori_ori_n1360_, ori_ori_n1361_, ori_ori_n1362_, ori_ori_n1363_, ori_ori_n1364_, ori_ori_n1365_, ori_ori_n1366_, ori_ori_n1367_, ori_ori_n1368_, ori_ori_n1369_, ori_ori_n1370_, ori_ori_n1371_, ori_ori_n1372_, ori_ori_n1373_, ori_ori_n1374_, ori_ori_n1375_, ori_ori_n1376_, ori_ori_n1377_, ori_ori_n1378_, ori_ori_n1379_, ori_ori_n1380_, ori_ori_n1381_, ori_ori_n1382_, ori_ori_n1383_, ori_ori_n1384_, ori_ori_n1385_, ori_ori_n1386_, ori_ori_n1387_, ori_ori_n1388_, ori_ori_n1389_, ori_ori_n1390_, ori_ori_n1391_, ori_ori_n1392_, ori_ori_n1393_, ori_ori_n1394_, ori_ori_n1395_, ori_ori_n1396_, ori_ori_n1397_, ori_ori_n1398_, ori_ori_n1399_, ori_ori_n1400_, ori_ori_n1401_, ori_ori_n1402_, ori_ori_n1403_, ori_ori_n1404_, ori_ori_n1405_, ori_ori_n1406_, ori_ori_n1407_, ori_ori_n1408_, ori_ori_n1409_, ori_ori_n1410_, ori_ori_n1411_, ori_ori_n1412_, ori_ori_n1413_, ori_ori_n1414_, ori_ori_n1415_, ori_ori_n1416_, ori_ori_n1417_, ori_ori_n1418_, ori_ori_n1419_, ori_ori_n1420_, ori_ori_n1421_, ori_ori_n1422_, ori_ori_n1424_, ori_ori_n1428_, ori_ori_n1429_, ori_ori_n1430_, ori_ori_n1431_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, mai_mai_n991_, mai_mai_n992_, mai_mai_n993_, mai_mai_n994_, mai_mai_n995_, mai_mai_n996_, mai_mai_n997_, mai_mai_n998_, mai_mai_n999_, mai_mai_n1000_, mai_mai_n1001_, mai_mai_n1002_, mai_mai_n1003_, mai_mai_n1004_, mai_mai_n1005_, mai_mai_n1006_, mai_mai_n1007_, mai_mai_n1008_, mai_mai_n1009_, mai_mai_n1010_, mai_mai_n1011_, mai_mai_n1012_, mai_mai_n1013_, mai_mai_n1014_, mai_mai_n1015_, mai_mai_n1016_, mai_mai_n1017_, mai_mai_n1018_, mai_mai_n1019_, mai_mai_n1020_, mai_mai_n1021_, mai_mai_n1022_, mai_mai_n1023_, mai_mai_n1024_, mai_mai_n1025_, mai_mai_n1026_, mai_mai_n1027_, mai_mai_n1028_, mai_mai_n1029_, mai_mai_n1030_, mai_mai_n1031_, mai_mai_n1032_, mai_mai_n1033_, mai_mai_n1034_, mai_mai_n1035_, mai_mai_n1036_, mai_mai_n1037_, mai_mai_n1038_, mai_mai_n1039_, mai_mai_n1040_, mai_mai_n1041_, mai_mai_n1042_, mai_mai_n1043_, mai_mai_n1044_, mai_mai_n1046_, mai_mai_n1047_, mai_mai_n1048_, mai_mai_n1049_, mai_mai_n1050_, mai_mai_n1051_, mai_mai_n1052_, mai_mai_n1053_, mai_mai_n1054_, mai_mai_n1055_, mai_mai_n1056_, mai_mai_n1057_, mai_mai_n1058_, mai_mai_n1059_, mai_mai_n1060_, mai_mai_n1061_, mai_mai_n1062_, mai_mai_n1063_, mai_mai_n1064_, mai_mai_n1065_, mai_mai_n1066_, mai_mai_n1067_, mai_mai_n1068_, mai_mai_n1069_, mai_mai_n1070_, mai_mai_n1071_, mai_mai_n1072_, mai_mai_n1073_, mai_mai_n1074_, mai_mai_n1075_, mai_mai_n1076_, mai_mai_n1077_, mai_mai_n1078_, mai_mai_n1079_, mai_mai_n1080_, mai_mai_n1081_, mai_mai_n1082_, mai_mai_n1083_, mai_mai_n1084_, mai_mai_n1085_, mai_mai_n1086_, mai_mai_n1087_, mai_mai_n1088_, mai_mai_n1089_, mai_mai_n1090_, mai_mai_n1091_, mai_mai_n1093_, mai_mai_n1094_, mai_mai_n1095_, mai_mai_n1096_, mai_mai_n1097_, mai_mai_n1098_, mai_mai_n1099_, mai_mai_n1100_, mai_mai_n1101_, mai_mai_n1102_, mai_mai_n1103_, mai_mai_n1104_, mai_mai_n1105_, mai_mai_n1106_, mai_mai_n1107_, mai_mai_n1108_, mai_mai_n1109_, mai_mai_n1110_, mai_mai_n1111_, mai_mai_n1112_, mai_mai_n1113_, mai_mai_n1114_, mai_mai_n1115_, mai_mai_n1116_, mai_mai_n1117_, mai_mai_n1119_, mai_mai_n1120_, mai_mai_n1121_, mai_mai_n1122_, mai_mai_n1123_, mai_mai_n1124_, mai_mai_n1125_, mai_mai_n1126_, mai_mai_n1127_, mai_mai_n1128_, mai_mai_n1129_, mai_mai_n1130_, mai_mai_n1131_, mai_mai_n1132_, mai_mai_n1133_, mai_mai_n1134_, mai_mai_n1135_, mai_mai_n1136_, mai_mai_n1137_, mai_mai_n1138_, mai_mai_n1139_, mai_mai_n1140_, mai_mai_n1141_, mai_mai_n1142_, mai_mai_n1143_, mai_mai_n1144_, mai_mai_n1145_, mai_mai_n1146_, mai_mai_n1147_, mai_mai_n1148_, mai_mai_n1149_, mai_mai_n1150_, mai_mai_n1151_, mai_mai_n1152_, mai_mai_n1153_, mai_mai_n1154_, mai_mai_n1155_, mai_mai_n1156_, mai_mai_n1157_, mai_mai_n1158_, mai_mai_n1159_, mai_mai_n1160_, mai_mai_n1162_, mai_mai_n1163_, mai_mai_n1164_, mai_mai_n1165_, mai_mai_n1166_, mai_mai_n1167_, mai_mai_n1168_, mai_mai_n1169_, mai_mai_n1170_, mai_mai_n1171_, mai_mai_n1172_, mai_mai_n1173_, mai_mai_n1174_, mai_mai_n1175_, mai_mai_n1176_, mai_mai_n1177_, mai_mai_n1178_, mai_mai_n1179_, mai_mai_n1180_, mai_mai_n1181_, mai_mai_n1182_, mai_mai_n1183_, mai_mai_n1184_, mai_mai_n1185_, mai_mai_n1186_, mai_mai_n1187_, mai_mai_n1188_, mai_mai_n1189_, mai_mai_n1190_, mai_mai_n1191_, mai_mai_n1192_, mai_mai_n1193_, mai_mai_n1194_, mai_mai_n1195_, mai_mai_n1196_, mai_mai_n1197_, mai_mai_n1198_, mai_mai_n1199_, mai_mai_n1200_, mai_mai_n1201_, mai_mai_n1202_, mai_mai_n1203_, mai_mai_n1204_, mai_mai_n1205_, mai_mai_n1206_, mai_mai_n1207_, mai_mai_n1208_, mai_mai_n1209_, mai_mai_n1210_, mai_mai_n1211_, mai_mai_n1212_, mai_mai_n1213_, mai_mai_n1214_, mai_mai_n1215_, mai_mai_n1216_, mai_mai_n1217_, mai_mai_n1218_, mai_mai_n1219_, mai_mai_n1220_, mai_mai_n1221_, mai_mai_n1222_, mai_mai_n1223_, mai_mai_n1224_, mai_mai_n1225_, mai_mai_n1227_, mai_mai_n1228_, mai_mai_n1229_, mai_mai_n1230_, mai_mai_n1231_, mai_mai_n1232_, mai_mai_n1233_, mai_mai_n1234_, mai_mai_n1235_, mai_mai_n1236_, mai_mai_n1237_, mai_mai_n1238_, mai_mai_n1239_, mai_mai_n1240_, mai_mai_n1241_, mai_mai_n1242_, mai_mai_n1243_, mai_mai_n1244_, mai_mai_n1245_, mai_mai_n1246_, mai_mai_n1247_, mai_mai_n1248_, mai_mai_n1249_, mai_mai_n1250_, mai_mai_n1251_, mai_mai_n1252_, mai_mai_n1253_, mai_mai_n1254_, mai_mai_n1255_, mai_mai_n1256_, mai_mai_n1257_, mai_mai_n1258_, mai_mai_n1259_, mai_mai_n1260_, mai_mai_n1261_, mai_mai_n1262_, mai_mai_n1263_, mai_mai_n1264_, mai_mai_n1265_, mai_mai_n1266_, mai_mai_n1267_, mai_mai_n1268_, mai_mai_n1269_, mai_mai_n1270_, mai_mai_n1271_, mai_mai_n1272_, mai_mai_n1273_, mai_mai_n1274_, mai_mai_n1275_, mai_mai_n1276_, mai_mai_n1277_, mai_mai_n1278_, mai_mai_n1279_, mai_mai_n1280_, mai_mai_n1281_, mai_mai_n1282_, mai_mai_n1283_, mai_mai_n1284_, mai_mai_n1285_, mai_mai_n1286_, mai_mai_n1287_, mai_mai_n1288_, mai_mai_n1289_, mai_mai_n1290_, mai_mai_n1292_, mai_mai_n1293_, mai_mai_n1294_, mai_mai_n1295_, mai_mai_n1296_, mai_mai_n1297_, mai_mai_n1298_, mai_mai_n1299_, mai_mai_n1300_, mai_mai_n1301_, mai_mai_n1302_, mai_mai_n1303_, mai_mai_n1304_, mai_mai_n1305_, mai_mai_n1306_, mai_mai_n1307_, mai_mai_n1308_, mai_mai_n1309_, mai_mai_n1310_, mai_mai_n1311_, mai_mai_n1312_, mai_mai_n1313_, mai_mai_n1314_, mai_mai_n1315_, mai_mai_n1316_, mai_mai_n1317_, mai_mai_n1318_, mai_mai_n1319_, mai_mai_n1320_, mai_mai_n1321_, mai_mai_n1322_, mai_mai_n1323_, mai_mai_n1324_, mai_mai_n1325_, mai_mai_n1326_, mai_mai_n1327_, mai_mai_n1328_, mai_mai_n1329_, mai_mai_n1330_, mai_mai_n1331_, mai_mai_n1332_, mai_mai_n1333_, mai_mai_n1334_, mai_mai_n1335_, mai_mai_n1336_, mai_mai_n1337_, mai_mai_n1338_, mai_mai_n1339_, mai_mai_n1341_, mai_mai_n1342_, mai_mai_n1343_, mai_mai_n1344_, mai_mai_n1345_, mai_mai_n1346_, mai_mai_n1347_, mai_mai_n1348_, mai_mai_n1349_, mai_mai_n1350_, mai_mai_n1351_, mai_mai_n1352_, mai_mai_n1353_, mai_mai_n1354_, mai_mai_n1355_, mai_mai_n1356_, mai_mai_n1357_, mai_mai_n1358_, mai_mai_n1359_, mai_mai_n1360_, mai_mai_n1361_, mai_mai_n1362_, mai_mai_n1363_, mai_mai_n1364_, mai_mai_n1365_, mai_mai_n1366_, mai_mai_n1367_, mai_mai_n1368_, mai_mai_n1369_, mai_mai_n1370_, mai_mai_n1371_, mai_mai_n1372_, mai_mai_n1373_, mai_mai_n1374_, mai_mai_n1375_, mai_mai_n1376_, mai_mai_n1377_, mai_mai_n1378_, mai_mai_n1379_, mai_mai_n1380_, mai_mai_n1381_, mai_mai_n1382_, mai_mai_n1383_, mai_mai_n1384_, mai_mai_n1385_, mai_mai_n1386_, mai_mai_n1387_, mai_mai_n1388_, mai_mai_n1389_, mai_mai_n1390_, mai_mai_n1391_, mai_mai_n1392_, mai_mai_n1393_, mai_mai_n1394_, mai_mai_n1395_, mai_mai_n1396_, mai_mai_n1397_, mai_mai_n1398_, mai_mai_n1399_, mai_mai_n1400_, mai_mai_n1401_, mai_mai_n1402_, mai_mai_n1403_, mai_mai_n1404_, mai_mai_n1405_, mai_mai_n1406_, mai_mai_n1407_, mai_mai_n1408_, mai_mai_n1409_, mai_mai_n1410_, mai_mai_n1411_, mai_mai_n1412_, mai_mai_n1413_, mai_mai_n1414_, mai_mai_n1415_, mai_mai_n1416_, mai_mai_n1417_, mai_mai_n1418_, mai_mai_n1419_, mai_mai_n1420_, mai_mai_n1421_, mai_mai_n1422_, mai_mai_n1423_, mai_mai_n1424_, mai_mai_n1425_, mai_mai_n1426_, mai_mai_n1427_, mai_mai_n1428_, mai_mai_n1429_, mai_mai_n1430_, mai_mai_n1431_, mai_mai_n1432_, mai_mai_n1433_, mai_mai_n1434_, mai_mai_n1435_, mai_mai_n1436_, mai_mai_n1437_, mai_mai_n1438_, mai_mai_n1439_, mai_mai_n1440_, mai_mai_n1441_, mai_mai_n1442_, mai_mai_n1443_, mai_mai_n1444_, mai_mai_n1445_, mai_mai_n1446_, mai_mai_n1447_, mai_mai_n1448_, mai_mai_n1449_, mai_mai_n1450_, mai_mai_n1451_, mai_mai_n1452_, mai_mai_n1453_, mai_mai_n1454_, mai_mai_n1455_, mai_mai_n1456_, mai_mai_n1457_, mai_mai_n1458_, mai_mai_n1459_, mai_mai_n1460_, mai_mai_n1461_, mai_mai_n1462_, mai_mai_n1463_, mai_mai_n1464_, mai_mai_n1465_, mai_mai_n1466_, mai_mai_n1467_, mai_mai_n1468_, mai_mai_n1469_, mai_mai_n1470_, mai_mai_n1471_, mai_mai_n1472_, mai_mai_n1473_, mai_mai_n1474_, mai_mai_n1475_, mai_mai_n1476_, mai_mai_n1477_, mai_mai_n1478_, mai_mai_n1479_, mai_mai_n1480_, mai_mai_n1481_, mai_mai_n1482_, mai_mai_n1483_, mai_mai_n1484_, mai_mai_n1485_, mai_mai_n1486_, mai_mai_n1487_, mai_mai_n1488_, mai_mai_n1489_, mai_mai_n1490_, mai_mai_n1491_, mai_mai_n1492_, mai_mai_n1493_, mai_mai_n1494_, mai_mai_n1495_, mai_mai_n1496_, mai_mai_n1497_, mai_mai_n1498_, mai_mai_n1499_, mai_mai_n1500_, mai_mai_n1501_, mai_mai_n1502_, mai_mai_n1503_, mai_mai_n1504_, mai_mai_n1505_, mai_mai_n1506_, mai_mai_n1507_, mai_mai_n1508_, mai_mai_n1509_, mai_mai_n1510_, mai_mai_n1511_, mai_mai_n1512_, mai_mai_n1513_, mai_mai_n1514_, mai_mai_n1515_, mai_mai_n1516_, mai_mai_n1517_, mai_mai_n1518_, mai_mai_n1519_, mai_mai_n1520_, mai_mai_n1521_, mai_mai_n1522_, mai_mai_n1523_, mai_mai_n1524_, mai_mai_n1525_, mai_mai_n1526_, mai_mai_n1527_, mai_mai_n1528_, mai_mai_n1529_, mai_mai_n1530_, mai_mai_n1531_, mai_mai_n1532_, mai_mai_n1533_, mai_mai_n1534_, mai_mai_n1535_, mai_mai_n1536_, mai_mai_n1537_, mai_mai_n1538_, mai_mai_n1539_, mai_mai_n1541_, mai_mai_n1542_, mai_mai_n1543_, mai_mai_n1544_, mai_mai_n1545_, mai_mai_n1546_, mai_mai_n1547_, mai_mai_n1548_, mai_mai_n1552_, mai_mai_n1553_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1039_, men_men_n1040_, men_men_n1041_, men_men_n1042_, men_men_n1043_, men_men_n1044_, men_men_n1045_, men_men_n1046_, men_men_n1047_, men_men_n1048_, men_men_n1049_, men_men_n1050_, men_men_n1051_, men_men_n1052_, men_men_n1053_, men_men_n1054_, men_men_n1055_, men_men_n1056_, men_men_n1057_, men_men_n1058_, men_men_n1060_, men_men_n1061_, men_men_n1062_, men_men_n1063_, men_men_n1064_, men_men_n1065_, men_men_n1066_, men_men_n1067_, men_men_n1068_, men_men_n1069_, men_men_n1070_, men_men_n1071_, men_men_n1072_, men_men_n1073_, men_men_n1074_, men_men_n1075_, men_men_n1076_, men_men_n1077_, men_men_n1078_, men_men_n1079_, men_men_n1080_, men_men_n1081_, men_men_n1082_, men_men_n1083_, men_men_n1084_, men_men_n1085_, men_men_n1086_, men_men_n1087_, men_men_n1088_, men_men_n1089_, men_men_n1090_, men_men_n1091_, men_men_n1092_, men_men_n1093_, men_men_n1094_, men_men_n1095_, men_men_n1096_, men_men_n1097_, men_men_n1098_, men_men_n1099_, men_men_n1100_, men_men_n1102_, men_men_n1103_, men_men_n1104_, men_men_n1105_, men_men_n1106_, men_men_n1107_, men_men_n1108_, men_men_n1109_, men_men_n1110_, men_men_n1111_, men_men_n1112_, men_men_n1113_, men_men_n1114_, men_men_n1115_, men_men_n1116_, men_men_n1117_, men_men_n1118_, men_men_n1119_, men_men_n1120_, men_men_n1121_, men_men_n1122_, men_men_n1123_, men_men_n1125_, men_men_n1126_, men_men_n1127_, men_men_n1128_, men_men_n1129_, men_men_n1130_, men_men_n1131_, men_men_n1132_, men_men_n1133_, men_men_n1134_, men_men_n1135_, men_men_n1136_, men_men_n1137_, men_men_n1138_, men_men_n1139_, men_men_n1140_, men_men_n1141_, men_men_n1142_, men_men_n1143_, men_men_n1144_, men_men_n1145_, men_men_n1146_, men_men_n1147_, men_men_n1148_, men_men_n1149_, men_men_n1150_, men_men_n1151_, men_men_n1152_, men_men_n1153_, men_men_n1154_, men_men_n1155_, men_men_n1156_, men_men_n1157_, men_men_n1158_, men_men_n1159_, men_men_n1160_, men_men_n1161_, men_men_n1162_, men_men_n1163_, men_men_n1164_, men_men_n1165_, men_men_n1166_, men_men_n1167_, men_men_n1168_, men_men_n1169_, men_men_n1170_, men_men_n1171_, men_men_n1172_, men_men_n1173_, men_men_n1174_, men_men_n1175_, men_men_n1176_, men_men_n1177_, men_men_n1179_, men_men_n1180_, men_men_n1181_, men_men_n1182_, men_men_n1183_, men_men_n1184_, men_men_n1185_, men_men_n1186_, men_men_n1187_, men_men_n1188_, men_men_n1189_, men_men_n1190_, men_men_n1191_, men_men_n1192_, men_men_n1193_, men_men_n1194_, men_men_n1195_, men_men_n1196_, men_men_n1197_, men_men_n1198_, men_men_n1199_, men_men_n1200_, men_men_n1201_, men_men_n1202_, men_men_n1203_, men_men_n1204_, men_men_n1205_, men_men_n1206_, men_men_n1207_, men_men_n1208_, men_men_n1209_, men_men_n1210_, men_men_n1211_, men_men_n1212_, men_men_n1213_, men_men_n1214_, men_men_n1215_, men_men_n1216_, men_men_n1217_, men_men_n1218_, men_men_n1219_, men_men_n1220_, men_men_n1221_, men_men_n1222_, men_men_n1223_, men_men_n1224_, men_men_n1225_, men_men_n1226_, men_men_n1227_, men_men_n1228_, men_men_n1229_, men_men_n1230_, men_men_n1231_, men_men_n1232_, men_men_n1233_, men_men_n1234_, men_men_n1235_, men_men_n1236_, men_men_n1237_, men_men_n1238_, men_men_n1239_, men_men_n1240_, men_men_n1241_, men_men_n1242_, men_men_n1243_, men_men_n1245_, men_men_n1246_, men_men_n1247_, men_men_n1248_, men_men_n1249_, men_men_n1250_, men_men_n1251_, men_men_n1252_, men_men_n1253_, men_men_n1254_, men_men_n1255_, men_men_n1256_, men_men_n1257_, men_men_n1258_, men_men_n1259_, men_men_n1260_, men_men_n1261_, men_men_n1262_, men_men_n1263_, men_men_n1264_, men_men_n1265_, men_men_n1266_, men_men_n1267_, men_men_n1268_, men_men_n1269_, men_men_n1270_, men_men_n1271_, men_men_n1272_, men_men_n1273_, men_men_n1274_, men_men_n1275_, men_men_n1276_, men_men_n1277_, men_men_n1278_, men_men_n1279_, men_men_n1280_, men_men_n1281_, men_men_n1282_, men_men_n1283_, men_men_n1284_, men_men_n1285_, men_men_n1286_, men_men_n1287_, men_men_n1288_, men_men_n1289_, men_men_n1290_, men_men_n1291_, men_men_n1292_, men_men_n1293_, men_men_n1294_, men_men_n1295_, men_men_n1296_, men_men_n1297_, men_men_n1298_, men_men_n1299_, men_men_n1300_, men_men_n1301_, men_men_n1302_, men_men_n1303_, men_men_n1304_, men_men_n1305_, men_men_n1306_, men_men_n1307_, men_men_n1308_, men_men_n1309_, men_men_n1310_, men_men_n1311_, men_men_n1312_, men_men_n1313_, men_men_n1315_, men_men_n1316_, men_men_n1317_, men_men_n1318_, men_men_n1319_, men_men_n1320_, men_men_n1321_, men_men_n1322_, men_men_n1323_, men_men_n1324_, men_men_n1325_, men_men_n1326_, men_men_n1327_, men_men_n1328_, men_men_n1329_, men_men_n1330_, men_men_n1331_, men_men_n1332_, men_men_n1333_, men_men_n1334_, men_men_n1335_, men_men_n1336_, men_men_n1337_, men_men_n1338_, men_men_n1339_, men_men_n1340_, men_men_n1341_, men_men_n1342_, men_men_n1343_, men_men_n1344_, men_men_n1345_, men_men_n1346_, men_men_n1347_, men_men_n1348_, men_men_n1349_, men_men_n1350_, men_men_n1351_, men_men_n1352_, men_men_n1353_, men_men_n1354_, men_men_n1355_, men_men_n1356_, men_men_n1357_, men_men_n1358_, men_men_n1359_, men_men_n1360_, men_men_n1361_, men_men_n1362_, men_men_n1363_, men_men_n1364_, men_men_n1365_, men_men_n1366_, men_men_n1367_, men_men_n1368_, men_men_n1369_, men_men_n1371_, men_men_n1372_, men_men_n1373_, men_men_n1374_, men_men_n1375_, men_men_n1376_, men_men_n1377_, men_men_n1378_, men_men_n1379_, men_men_n1380_, men_men_n1381_, men_men_n1382_, men_men_n1383_, men_men_n1384_, men_men_n1385_, men_men_n1386_, men_men_n1387_, men_men_n1388_, men_men_n1389_, men_men_n1390_, men_men_n1391_, men_men_n1392_, men_men_n1393_, men_men_n1394_, men_men_n1395_, men_men_n1396_, men_men_n1397_, men_men_n1398_, men_men_n1399_, men_men_n1400_, men_men_n1401_, men_men_n1402_, men_men_n1403_, men_men_n1404_, men_men_n1405_, men_men_n1406_, men_men_n1407_, men_men_n1408_, men_men_n1409_, men_men_n1410_, men_men_n1411_, men_men_n1412_, men_men_n1413_, men_men_n1414_, men_men_n1415_, men_men_n1416_, men_men_n1417_, men_men_n1418_, men_men_n1419_, men_men_n1420_, men_men_n1421_, men_men_n1422_, men_men_n1423_, men_men_n1424_, men_men_n1425_, men_men_n1426_, men_men_n1427_, men_men_n1428_, men_men_n1429_, men_men_n1430_, men_men_n1431_, men_men_n1432_, men_men_n1433_, men_men_n1434_, men_men_n1435_, men_men_n1436_, men_men_n1437_, men_men_n1438_, men_men_n1439_, men_men_n1440_, men_men_n1441_, men_men_n1442_, men_men_n1443_, men_men_n1444_, men_men_n1445_, men_men_n1446_, men_men_n1447_, men_men_n1448_, men_men_n1449_, men_men_n1450_, men_men_n1451_, men_men_n1452_, men_men_n1453_, men_men_n1454_, men_men_n1455_, men_men_n1456_, men_men_n1457_, men_men_n1458_, men_men_n1459_, men_men_n1460_, men_men_n1461_, men_men_n1462_, men_men_n1463_, men_men_n1464_, men_men_n1465_, men_men_n1466_, men_men_n1467_, men_men_n1468_, men_men_n1469_, men_men_n1470_, men_men_n1471_, men_men_n1472_, men_men_n1473_, men_men_n1474_, men_men_n1475_, men_men_n1476_, men_men_n1477_, men_men_n1478_, men_men_n1479_, men_men_n1480_, men_men_n1481_, men_men_n1482_, men_men_n1483_, men_men_n1484_, men_men_n1485_, men_men_n1486_, men_men_n1487_, men_men_n1488_, men_men_n1489_, men_men_n1490_, men_men_n1491_, men_men_n1492_, men_men_n1493_, men_men_n1494_, men_men_n1495_, men_men_n1496_, men_men_n1497_, men_men_n1498_, men_men_n1499_, men_men_n1500_, men_men_n1501_, men_men_n1502_, men_men_n1503_, men_men_n1504_, men_men_n1505_, men_men_n1506_, men_men_n1507_, men_men_n1508_, men_men_n1509_, men_men_n1510_, men_men_n1511_, men_men_n1512_, men_men_n1513_, men_men_n1514_, men_men_n1515_, men_men_n1516_, men_men_n1517_, men_men_n1518_, men_men_n1519_, men_men_n1520_, men_men_n1521_, men_men_n1522_, men_men_n1523_, men_men_n1524_, men_men_n1525_, men_men_n1526_, men_men_n1527_, men_men_n1528_, men_men_n1529_, men_men_n1530_, men_men_n1531_, men_men_n1532_, men_men_n1533_, men_men_n1534_, men_men_n1535_, men_men_n1536_, men_men_n1537_, men_men_n1538_, men_men_n1539_, men_men_n1540_, men_men_n1541_, men_men_n1542_, men_men_n1543_, men_men_n1544_, men_men_n1545_, men_men_n1546_, men_men_n1547_, men_men_n1548_, men_men_n1549_, men_men_n1550_, men_men_n1551_, men_men_n1552_, men_men_n1553_, men_men_n1554_, men_men_n1555_, men_men_n1556_, men_men_n1557_, men_men_n1558_, men_men_n1559_, men_men_n1560_, men_men_n1561_, men_men_n1562_, men_men_n1563_, men_men_n1564_, men_men_n1565_, men_men_n1566_, men_men_n1567_, men_men_n1568_, men_men_n1569_, men_men_n1570_, men_men_n1571_, men_men_n1572_, men_men_n1574_, men_men_n1575_, men_men_n1576_, men_men_n1577_, men_men_n1578_, men_men_n1579_, men_men_n1580_, men_men_n1581_, men_men_n1585_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06, ori07, mai07, men07, ori08, mai08, men08, ori09, mai09, men09, ori10, mai10, men10, ori11, mai11, men11, ori12, mai12, men12, ori13, mai13, men13;
  AN2        o0000(.A(b), .B(a), .Y(ori_ori_n29_));
  NO2        o0001(.A(d), .B(c), .Y(ori_ori_n30_));
  AN2        o0002(.A(f), .B(e), .Y(ori_ori_n31_));
  NA3        o0003(.A(ori_ori_n31_), .B(ori_ori_n30_), .C(ori_ori_n29_), .Y(ori_ori_n32_));
  NOi32      o0004(.An(m), .Bn(l), .C(n), .Y(ori_ori_n33_));
  NOi32      o0005(.An(i), .Bn(g), .C(h), .Y(ori_ori_n34_));
  NA2        o0006(.A(ori_ori_n34_), .B(ori_ori_n33_), .Y(ori_ori_n35_));
  AN2        o0007(.A(m), .B(l), .Y(ori_ori_n36_));
  NOi32      o0008(.An(j), .Bn(g), .C(k), .Y(ori_ori_n37_));
  NA2        o0009(.A(ori_ori_n37_), .B(ori_ori_n36_), .Y(ori_ori_n38_));
  NO2        o0010(.A(ori_ori_n38_), .B(n), .Y(ori_ori_n39_));
  INV        o0011(.A(h), .Y(ori_ori_n40_));
  NAi21      o0012(.An(j), .B(l), .Y(ori_ori_n41_));
  NAi32      o0013(.An(n), .Bn(g), .C(m), .Y(ori_ori_n42_));
  NO3        o0014(.A(ori_ori_n42_), .B(ori_ori_n41_), .C(ori_ori_n40_), .Y(ori_ori_n43_));
  NAi31      o0015(.An(n), .B(m), .C(l), .Y(ori_ori_n44_));
  INV        o0016(.A(i), .Y(ori_ori_n45_));
  AN2        o0017(.A(h), .B(g), .Y(ori_ori_n46_));
  NA2        o0018(.A(ori_ori_n46_), .B(ori_ori_n45_), .Y(ori_ori_n47_));
  NO2        o0019(.A(ori_ori_n47_), .B(ori_ori_n44_), .Y(ori_ori_n48_));
  NAi21      o0020(.An(n), .B(m), .Y(ori_ori_n49_));
  NOi32      o0021(.An(k), .Bn(h), .C(l), .Y(ori_ori_n50_));
  NOi32      o0022(.An(k), .Bn(h), .C(g), .Y(ori_ori_n51_));
  INV        o0023(.A(ori_ori_n51_), .Y(ori_ori_n52_));
  NO2        o0024(.A(ori_ori_n52_), .B(ori_ori_n49_), .Y(ori_ori_n53_));
  NO3        o0025(.A(ori_ori_n53_), .B(ori_ori_n48_), .C(ori_ori_n39_), .Y(ori_ori_n54_));
  AOI210     o0026(.A0(ori_ori_n54_), .A1(ori_ori_n35_), .B0(ori_ori_n32_), .Y(ori_ori_n55_));
  INV        o0027(.A(c), .Y(ori_ori_n56_));
  NA2        o0028(.A(e), .B(b), .Y(ori_ori_n57_));
  NO2        o0029(.A(ori_ori_n57_), .B(ori_ori_n56_), .Y(ori_ori_n58_));
  INV        o0030(.A(d), .Y(ori_ori_n59_));
  NA2        o0031(.A(g), .B(ori_ori_n59_), .Y(ori_ori_n60_));
  NAi21      o0032(.An(i), .B(h), .Y(ori_ori_n61_));
  NAi31      o0033(.An(i), .B(l), .C(j), .Y(ori_ori_n62_));
  OAI220     o0034(.A0(ori_ori_n62_), .A1(ori_ori_n49_), .B0(ori_ori_n61_), .B1(ori_ori_n44_), .Y(ori_ori_n63_));
  NAi31      o0035(.An(ori_ori_n60_), .B(ori_ori_n63_), .C(ori_ori_n58_), .Y(ori_ori_n64_));
  NAi41      o0036(.An(e), .B(d), .C(b), .D(a), .Y(ori_ori_n65_));
  NA2        o0037(.A(g), .B(f), .Y(ori_ori_n66_));
  NO2        o0038(.A(ori_ori_n66_), .B(ori_ori_n65_), .Y(ori_ori_n67_));
  NAi21      o0039(.An(i), .B(j), .Y(ori_ori_n68_));
  NAi32      o0040(.An(n), .Bn(k), .C(m), .Y(ori_ori_n69_));
  NAi31      o0041(.An(l), .B(m), .C(k), .Y(ori_ori_n70_));
  NAi21      o0042(.An(e), .B(h), .Y(ori_ori_n71_));
  NAi41      o0043(.An(n), .B(d), .C(b), .D(a), .Y(ori_ori_n72_));
  INV        o0044(.A(m), .Y(ori_ori_n73_));
  NOi21      o0045(.An(k), .B(l), .Y(ori_ori_n74_));
  NA2        o0046(.A(ori_ori_n74_), .B(ori_ori_n73_), .Y(ori_ori_n75_));
  AN4        o0047(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n76_));
  NOi31      o0048(.An(h), .B(g), .C(f), .Y(ori_ori_n77_));
  NA2        o0049(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n78_));
  NAi32      o0050(.An(m), .Bn(k), .C(j), .Y(ori_ori_n79_));
  NOi32      o0051(.An(h), .Bn(g), .C(f), .Y(ori_ori_n80_));
  NA2        o0052(.A(ori_ori_n80_), .B(ori_ori_n76_), .Y(ori_ori_n81_));
  OA220      o0053(.A0(ori_ori_n81_), .A1(ori_ori_n79_), .B0(ori_ori_n78_), .B1(ori_ori_n75_), .Y(ori_ori_n82_));
  NA2        o0054(.A(ori_ori_n82_), .B(ori_ori_n64_), .Y(ori_ori_n83_));
  INV        o0055(.A(n), .Y(ori_ori_n84_));
  NOi32      o0056(.An(e), .Bn(b), .C(d), .Y(ori_ori_n85_));
  NA2        o0057(.A(ori_ori_n85_), .B(ori_ori_n84_), .Y(ori_ori_n86_));
  INV        o0058(.A(j), .Y(ori_ori_n87_));
  AN3        o0059(.A(m), .B(k), .C(i), .Y(ori_ori_n88_));
  NA3        o0060(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(g), .Y(ori_ori_n89_));
  NO2        o0061(.A(ori_ori_n89_), .B(f), .Y(ori_ori_n90_));
  NAi32      o0062(.An(g), .Bn(f), .C(h), .Y(ori_ori_n91_));
  NAi31      o0063(.An(j), .B(m), .C(l), .Y(ori_ori_n92_));
  NO2        o0064(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n93_));
  NA2        o0065(.A(m), .B(l), .Y(ori_ori_n94_));
  NAi31      o0066(.An(k), .B(j), .C(g), .Y(ori_ori_n95_));
  NO3        o0067(.A(ori_ori_n95_), .B(ori_ori_n94_), .C(f), .Y(ori_ori_n96_));
  AN2        o0068(.A(j), .B(g), .Y(ori_ori_n97_));
  NOi32      o0069(.An(m), .Bn(l), .C(i), .Y(ori_ori_n98_));
  NOi21      o0070(.An(g), .B(i), .Y(ori_ori_n99_));
  NOi32      o0071(.An(m), .Bn(j), .C(k), .Y(ori_ori_n100_));
  AOI220     o0072(.A0(ori_ori_n100_), .A1(ori_ori_n99_), .B0(ori_ori_n98_), .B1(ori_ori_n97_), .Y(ori_ori_n101_));
  NO2        o0073(.A(ori_ori_n101_), .B(f), .Y(ori_ori_n102_));
  NO3        o0074(.A(ori_ori_n102_), .B(ori_ori_n93_), .C(ori_ori_n90_), .Y(ori_ori_n103_));
  NAi41      o0075(.An(m), .B(n), .C(k), .D(i), .Y(ori_ori_n104_));
  AN2        o0076(.A(e), .B(b), .Y(ori_ori_n105_));
  NOi31      o0077(.An(c), .B(h), .C(f), .Y(ori_ori_n106_));
  NA2        o0078(.A(ori_ori_n106_), .B(ori_ori_n105_), .Y(ori_ori_n107_));
  NO2        o0079(.A(ori_ori_n107_), .B(ori_ori_n104_), .Y(ori_ori_n108_));
  NOi21      o0080(.An(g), .B(f), .Y(ori_ori_n109_));
  NOi21      o0081(.An(i), .B(h), .Y(ori_ori_n110_));
  NA3        o0082(.A(ori_ori_n110_), .B(ori_ori_n109_), .C(ori_ori_n36_), .Y(ori_ori_n111_));
  INV        o0083(.A(a), .Y(ori_ori_n112_));
  NA2        o0084(.A(ori_ori_n105_), .B(ori_ori_n112_), .Y(ori_ori_n113_));
  INV        o0085(.A(l), .Y(ori_ori_n114_));
  NOi21      o0086(.An(m), .B(n), .Y(ori_ori_n115_));
  AN2        o0087(.A(k), .B(h), .Y(ori_ori_n116_));
  NO2        o0088(.A(ori_ori_n111_), .B(ori_ori_n86_), .Y(ori_ori_n117_));
  INV        o0089(.A(b), .Y(ori_ori_n118_));
  NA2        o0090(.A(l), .B(j), .Y(ori_ori_n119_));
  AN2        o0091(.A(k), .B(i), .Y(ori_ori_n120_));
  NA2        o0092(.A(ori_ori_n120_), .B(ori_ori_n119_), .Y(ori_ori_n121_));
  NA2        o0093(.A(g), .B(e), .Y(ori_ori_n122_));
  NOi32      o0094(.An(c), .Bn(a), .C(d), .Y(ori_ori_n123_));
  NA2        o0095(.A(ori_ori_n123_), .B(ori_ori_n115_), .Y(ori_ori_n124_));
  NO2        o0096(.A(ori_ori_n117_), .B(ori_ori_n108_), .Y(ori_ori_n125_));
  OAI210     o0097(.A0(ori_ori_n103_), .A1(ori_ori_n86_), .B0(ori_ori_n125_), .Y(ori_ori_n126_));
  NOi31      o0098(.An(k), .B(m), .C(j), .Y(ori_ori_n127_));
  NA3        o0099(.A(ori_ori_n127_), .B(ori_ori_n77_), .C(ori_ori_n76_), .Y(ori_ori_n128_));
  NOi31      o0100(.An(k), .B(m), .C(i), .Y(ori_ori_n129_));
  NA3        o0101(.A(ori_ori_n129_), .B(ori_ori_n80_), .C(ori_ori_n76_), .Y(ori_ori_n130_));
  NA2        o0102(.A(ori_ori_n130_), .B(ori_ori_n128_), .Y(ori_ori_n131_));
  NOi32      o0103(.An(f), .Bn(b), .C(e), .Y(ori_ori_n132_));
  NAi21      o0104(.An(g), .B(h), .Y(ori_ori_n133_));
  NAi21      o0105(.An(m), .B(n), .Y(ori_ori_n134_));
  NAi21      o0106(.An(j), .B(k), .Y(ori_ori_n135_));
  NO3        o0107(.A(ori_ori_n135_), .B(ori_ori_n134_), .C(ori_ori_n133_), .Y(ori_ori_n136_));
  NAi41      o0108(.An(e), .B(f), .C(d), .D(b), .Y(ori_ori_n137_));
  NAi31      o0109(.An(j), .B(k), .C(h), .Y(ori_ori_n138_));
  NO3        o0110(.A(ori_ori_n138_), .B(ori_ori_n137_), .C(ori_ori_n134_), .Y(ori_ori_n139_));
  AOI210     o0111(.A0(ori_ori_n136_), .A1(ori_ori_n132_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NO2        o0112(.A(k), .B(j), .Y(ori_ori_n141_));
  NO2        o0113(.A(ori_ori_n141_), .B(ori_ori_n134_), .Y(ori_ori_n142_));
  AN2        o0114(.A(k), .B(j), .Y(ori_ori_n143_));
  NAi21      o0115(.An(c), .B(b), .Y(ori_ori_n144_));
  NA2        o0116(.A(f), .B(d), .Y(ori_ori_n145_));
  NO4        o0117(.A(ori_ori_n145_), .B(ori_ori_n144_), .C(ori_ori_n143_), .D(ori_ori_n133_), .Y(ori_ori_n146_));
  NA2        o0118(.A(h), .B(c), .Y(ori_ori_n147_));
  NAi31      o0119(.An(f), .B(e), .C(b), .Y(ori_ori_n148_));
  NA2        o0120(.A(ori_ori_n146_), .B(ori_ori_n142_), .Y(ori_ori_n149_));
  NA2        o0121(.A(d), .B(b), .Y(ori_ori_n150_));
  NAi21      o0122(.An(e), .B(f), .Y(ori_ori_n151_));
  NO2        o0123(.A(ori_ori_n151_), .B(ori_ori_n150_), .Y(ori_ori_n152_));
  NA2        o0124(.A(b), .B(a), .Y(ori_ori_n153_));
  NAi21      o0125(.An(e), .B(g), .Y(ori_ori_n154_));
  NAi21      o0126(.An(c), .B(d), .Y(ori_ori_n155_));
  NAi31      o0127(.An(l), .B(k), .C(h), .Y(ori_ori_n156_));
  NO2        o0128(.A(ori_ori_n134_), .B(ori_ori_n156_), .Y(ori_ori_n157_));
  NA2        o0129(.A(ori_ori_n157_), .B(ori_ori_n152_), .Y(ori_ori_n158_));
  NAi41      o0130(.An(ori_ori_n131_), .B(ori_ori_n158_), .C(ori_ori_n149_), .D(ori_ori_n140_), .Y(ori_ori_n159_));
  NAi31      o0131(.An(e), .B(f), .C(b), .Y(ori_ori_n160_));
  NOi21      o0132(.An(g), .B(d), .Y(ori_ori_n161_));
  NO2        o0133(.A(ori_ori_n161_), .B(ori_ori_n160_), .Y(ori_ori_n162_));
  NOi21      o0134(.An(h), .B(i), .Y(ori_ori_n163_));
  NOi21      o0135(.An(k), .B(m), .Y(ori_ori_n164_));
  NA3        o0136(.A(ori_ori_n164_), .B(ori_ori_n163_), .C(n), .Y(ori_ori_n165_));
  NOi21      o0137(.An(ori_ori_n162_), .B(ori_ori_n165_), .Y(ori_ori_n166_));
  NOi21      o0138(.An(h), .B(g), .Y(ori_ori_n167_));
  NO2        o0139(.A(ori_ori_n145_), .B(ori_ori_n144_), .Y(ori_ori_n168_));
  NAi31      o0140(.An(l), .B(j), .C(h), .Y(ori_ori_n169_));
  NO2        o0141(.A(ori_ori_n169_), .B(ori_ori_n49_), .Y(ori_ori_n170_));
  NA2        o0142(.A(ori_ori_n170_), .B(ori_ori_n67_), .Y(ori_ori_n171_));
  NOi32      o0143(.An(n), .Bn(k), .C(m), .Y(ori_ori_n172_));
  NA2        o0144(.A(l), .B(i), .Y(ori_ori_n173_));
  INV        o0145(.A(ori_ori_n171_), .Y(ori_ori_n174_));
  NAi31      o0146(.An(d), .B(f), .C(c), .Y(ori_ori_n175_));
  NAi31      o0147(.An(e), .B(f), .C(c), .Y(ori_ori_n176_));
  NA2        o0148(.A(ori_ori_n176_), .B(ori_ori_n175_), .Y(ori_ori_n177_));
  NA2        o0149(.A(j), .B(h), .Y(ori_ori_n178_));
  OR3        o0150(.A(n), .B(m), .C(k), .Y(ori_ori_n179_));
  NO2        o0151(.A(ori_ori_n179_), .B(ori_ori_n178_), .Y(ori_ori_n180_));
  NAi32      o0152(.An(m), .Bn(k), .C(n), .Y(ori_ori_n181_));
  NO2        o0153(.A(ori_ori_n181_), .B(ori_ori_n178_), .Y(ori_ori_n182_));
  AOI220     o0154(.A0(ori_ori_n182_), .A1(ori_ori_n162_), .B0(ori_ori_n180_), .B1(ori_ori_n177_), .Y(ori_ori_n183_));
  NO2        o0155(.A(n), .B(m), .Y(ori_ori_n184_));
  NA2        o0156(.A(ori_ori_n184_), .B(ori_ori_n50_), .Y(ori_ori_n185_));
  NAi21      o0157(.An(f), .B(e), .Y(ori_ori_n186_));
  NA2        o0158(.A(d), .B(c), .Y(ori_ori_n187_));
  NO2        o0159(.A(ori_ori_n187_), .B(ori_ori_n186_), .Y(ori_ori_n188_));
  NOi21      o0160(.An(ori_ori_n188_), .B(ori_ori_n185_), .Y(ori_ori_n189_));
  NAi31      o0161(.An(m), .B(n), .C(b), .Y(ori_ori_n190_));
  NA2        o0162(.A(k), .B(i), .Y(ori_ori_n191_));
  NAi21      o0163(.An(h), .B(f), .Y(ori_ori_n192_));
  NO2        o0164(.A(ori_ori_n192_), .B(ori_ori_n191_), .Y(ori_ori_n193_));
  NO2        o0165(.A(ori_ori_n190_), .B(ori_ori_n155_), .Y(ori_ori_n194_));
  NA2        o0166(.A(ori_ori_n194_), .B(ori_ori_n193_), .Y(ori_ori_n195_));
  NOi32      o0167(.An(f), .Bn(c), .C(d), .Y(ori_ori_n196_));
  NOi32      o0168(.An(f), .Bn(c), .C(e), .Y(ori_ori_n197_));
  NO2        o0169(.A(ori_ori_n197_), .B(ori_ori_n196_), .Y(ori_ori_n198_));
  NO3        o0170(.A(n), .B(m), .C(j), .Y(ori_ori_n199_));
  NA2        o0171(.A(ori_ori_n199_), .B(ori_ori_n116_), .Y(ori_ori_n200_));
  AO210      o0172(.A0(ori_ori_n200_), .A1(ori_ori_n185_), .B0(ori_ori_n198_), .Y(ori_ori_n201_));
  NAi41      o0173(.An(ori_ori_n189_), .B(ori_ori_n201_), .C(ori_ori_n195_), .D(ori_ori_n183_), .Y(ori_ori_n202_));
  OR4        o0174(.A(ori_ori_n202_), .B(ori_ori_n174_), .C(ori_ori_n166_), .D(ori_ori_n159_), .Y(ori_ori_n203_));
  NO4        o0175(.A(ori_ori_n203_), .B(ori_ori_n126_), .C(ori_ori_n83_), .D(ori_ori_n55_), .Y(ori_ori_n204_));
  NA3        o0176(.A(m), .B(ori_ori_n114_), .C(j), .Y(ori_ori_n205_));
  NAi31      o0177(.An(n), .B(h), .C(g), .Y(ori_ori_n206_));
  NO2        o0178(.A(ori_ori_n206_), .B(ori_ori_n205_), .Y(ori_ori_n207_));
  NOi32      o0179(.An(m), .Bn(k), .C(l), .Y(ori_ori_n208_));
  NA3        o0180(.A(ori_ori_n208_), .B(ori_ori_n87_), .C(g), .Y(ori_ori_n209_));
  NO2        o0181(.A(ori_ori_n209_), .B(n), .Y(ori_ori_n210_));
  NOi21      o0182(.An(k), .B(j), .Y(ori_ori_n211_));
  NA4        o0183(.A(ori_ori_n211_), .B(ori_ori_n115_), .C(i), .D(g), .Y(ori_ori_n212_));
  AN2        o0184(.A(i), .B(g), .Y(ori_ori_n213_));
  NA3        o0185(.A(ori_ori_n74_), .B(ori_ori_n213_), .C(ori_ori_n115_), .Y(ori_ori_n214_));
  NO2        o0186(.A(ori_ori_n210_), .B(ori_ori_n207_), .Y(ori_ori_n215_));
  NAi41      o0187(.An(d), .B(n), .C(e), .D(b), .Y(ori_ori_n216_));
  INV        o0188(.A(ori_ori_n216_), .Y(ori_ori_n217_));
  INV        o0189(.A(f), .Y(ori_ori_n218_));
  INV        o0190(.A(g), .Y(ori_ori_n219_));
  NOi31      o0191(.An(i), .B(j), .C(h), .Y(ori_ori_n220_));
  NOi21      o0192(.An(l), .B(m), .Y(ori_ori_n221_));
  NA2        o0193(.A(ori_ori_n221_), .B(ori_ori_n220_), .Y(ori_ori_n222_));
  NO3        o0194(.A(ori_ori_n222_), .B(ori_ori_n219_), .C(ori_ori_n218_), .Y(ori_ori_n223_));
  NA2        o0195(.A(ori_ori_n223_), .B(ori_ori_n217_), .Y(ori_ori_n224_));
  OAI210     o0196(.A0(ori_ori_n215_), .A1(ori_ori_n32_), .B0(ori_ori_n224_), .Y(ori_ori_n225_));
  NOi21      o0197(.An(n), .B(m), .Y(ori_ori_n226_));
  NOi32      o0198(.An(l), .Bn(i), .C(j), .Y(ori_ori_n227_));
  NA2        o0199(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  OA220      o0200(.A0(ori_ori_n228_), .A1(ori_ori_n107_), .B0(ori_ori_n79_), .B1(ori_ori_n78_), .Y(ori_ori_n229_));
  NAi21      o0201(.An(j), .B(h), .Y(ori_ori_n230_));
  XN2        o0202(.A(i), .B(h), .Y(ori_ori_n231_));
  NA2        o0203(.A(ori_ori_n231_), .B(ori_ori_n230_), .Y(ori_ori_n232_));
  NOi31      o0204(.An(k), .B(n), .C(m), .Y(ori_ori_n233_));
  NOi31      o0205(.An(ori_ori_n233_), .B(ori_ori_n187_), .C(ori_ori_n186_), .Y(ori_ori_n234_));
  NA2        o0206(.A(ori_ori_n234_), .B(ori_ori_n232_), .Y(ori_ori_n235_));
  NAi31      o0207(.An(f), .B(e), .C(c), .Y(ori_ori_n236_));
  NO4        o0208(.A(ori_ori_n236_), .B(ori_ori_n179_), .C(ori_ori_n178_), .D(ori_ori_n59_), .Y(ori_ori_n237_));
  NA4        o0209(.A(n), .B(e), .C(c), .D(b), .Y(ori_ori_n238_));
  NAi32      o0210(.An(m), .Bn(i), .C(k), .Y(ori_ori_n239_));
  INV        o0211(.A(k), .Y(ori_ori_n240_));
  INV        o0212(.A(ori_ori_n237_), .Y(ori_ori_n241_));
  NAi21      o0213(.An(n), .B(a), .Y(ori_ori_n242_));
  NO2        o0214(.A(ori_ori_n242_), .B(ori_ori_n150_), .Y(ori_ori_n243_));
  NAi41      o0215(.An(g), .B(m), .C(k), .D(h), .Y(ori_ori_n244_));
  NO2        o0216(.A(ori_ori_n244_), .B(e), .Y(ori_ori_n245_));
  NA2        o0217(.A(ori_ori_n245_), .B(ori_ori_n243_), .Y(ori_ori_n246_));
  AN4        o0218(.A(ori_ori_n246_), .B(ori_ori_n241_), .C(ori_ori_n235_), .D(ori_ori_n229_), .Y(ori_ori_n247_));
  OR2        o0219(.A(h), .B(g), .Y(ori_ori_n248_));
  NO2        o0220(.A(ori_ori_n248_), .B(ori_ori_n104_), .Y(ori_ori_n249_));
  NA2        o0221(.A(ori_ori_n249_), .B(ori_ori_n132_), .Y(ori_ori_n250_));
  NAi41      o0222(.An(e), .B(n), .C(d), .D(b), .Y(ori_ori_n251_));
  NO2        o0223(.A(ori_ori_n251_), .B(ori_ori_n218_), .Y(ori_ori_n252_));
  NA2        o0224(.A(ori_ori_n164_), .B(ori_ori_n110_), .Y(ori_ori_n253_));
  NAi21      o0225(.An(ori_ori_n253_), .B(ori_ori_n252_), .Y(ori_ori_n254_));
  NO2        o0226(.A(n), .B(a), .Y(ori_ori_n255_));
  NAi31      o0227(.An(ori_ori_n244_), .B(ori_ori_n255_), .C(ori_ori_n105_), .Y(ori_ori_n256_));
  AN2        o0228(.A(ori_ori_n256_), .B(ori_ori_n254_), .Y(ori_ori_n257_));
  NAi21      o0229(.An(h), .B(i), .Y(ori_ori_n258_));
  NA2        o0230(.A(ori_ori_n184_), .B(k), .Y(ori_ori_n259_));
  NO2        o0231(.A(ori_ori_n259_), .B(ori_ori_n258_), .Y(ori_ori_n260_));
  NA2        o0232(.A(ori_ori_n260_), .B(ori_ori_n196_), .Y(ori_ori_n261_));
  NA3        o0233(.A(ori_ori_n261_), .B(ori_ori_n257_), .C(ori_ori_n250_), .Y(ori_ori_n262_));
  NOi21      o0234(.An(g), .B(e), .Y(ori_ori_n263_));
  NO2        o0235(.A(ori_ori_n72_), .B(ori_ori_n73_), .Y(ori_ori_n264_));
  NA2        o0236(.A(ori_ori_n264_), .B(ori_ori_n263_), .Y(ori_ori_n265_));
  NOi32      o0237(.An(l), .Bn(j), .C(i), .Y(ori_ori_n266_));
  AOI210     o0238(.A0(ori_ori_n74_), .A1(ori_ori_n87_), .B0(ori_ori_n266_), .Y(ori_ori_n267_));
  NO2        o0239(.A(ori_ori_n258_), .B(ori_ori_n44_), .Y(ori_ori_n268_));
  NAi21      o0240(.An(f), .B(g), .Y(ori_ori_n269_));
  NO2        o0241(.A(ori_ori_n269_), .B(ori_ori_n65_), .Y(ori_ori_n270_));
  NO2        o0242(.A(ori_ori_n69_), .B(ori_ori_n119_), .Y(ori_ori_n271_));
  AOI220     o0243(.A0(ori_ori_n271_), .A1(ori_ori_n270_), .B0(ori_ori_n268_), .B1(ori_ori_n67_), .Y(ori_ori_n272_));
  OAI210     o0244(.A0(ori_ori_n267_), .A1(ori_ori_n265_), .B0(ori_ori_n272_), .Y(ori_ori_n273_));
  NO2        o0245(.A(ori_ori_n135_), .B(ori_ori_n49_), .Y(ori_ori_n274_));
  NOi41      o0246(.An(ori_ori_n247_), .B(ori_ori_n273_), .C(ori_ori_n262_), .D(ori_ori_n225_), .Y(ori_ori_n275_));
  NO4        o0247(.A(ori_ori_n207_), .B(ori_ori_n48_), .C(ori_ori_n43_), .D(ori_ori_n39_), .Y(ori_ori_n276_));
  NO2        o0248(.A(ori_ori_n276_), .B(ori_ori_n113_), .Y(ori_ori_n277_));
  NA3        o0249(.A(ori_ori_n59_), .B(c), .C(b), .Y(ori_ori_n278_));
  NAi21      o0250(.An(h), .B(g), .Y(ori_ori_n279_));
  OR4        o0251(.A(ori_ori_n279_), .B(ori_ori_n278_), .C(ori_ori_n228_), .D(e), .Y(ori_ori_n280_));
  NO2        o0252(.A(ori_ori_n253_), .B(ori_ori_n269_), .Y(ori_ori_n281_));
  NAi31      o0253(.An(g), .B(k), .C(h), .Y(ori_ori_n282_));
  NAi31      o0254(.An(e), .B(d), .C(a), .Y(ori_ori_n283_));
  INV        o0255(.A(ori_ori_n280_), .Y(ori_ori_n284_));
  NA4        o0256(.A(ori_ori_n164_), .B(ori_ori_n80_), .C(ori_ori_n76_), .D(ori_ori_n119_), .Y(ori_ori_n285_));
  NA3        o0257(.A(ori_ori_n164_), .B(ori_ori_n163_), .C(ori_ori_n84_), .Y(ori_ori_n286_));
  NO2        o0258(.A(ori_ori_n286_), .B(ori_ori_n198_), .Y(ori_ori_n287_));
  NOi21      o0259(.An(ori_ori_n285_), .B(ori_ori_n287_), .Y(ori_ori_n288_));
  NA3        o0260(.A(e), .B(c), .C(b), .Y(ori_ori_n289_));
  NO2        o0261(.A(ori_ori_n60_), .B(ori_ori_n289_), .Y(ori_ori_n290_));
  NAi32      o0262(.An(k), .Bn(i), .C(j), .Y(ori_ori_n291_));
  NAi31      o0263(.An(h), .B(l), .C(i), .Y(ori_ori_n292_));
  NA3        o0264(.A(ori_ori_n292_), .B(ori_ori_n291_), .C(ori_ori_n169_), .Y(ori_ori_n293_));
  NOi21      o0265(.An(ori_ori_n293_), .B(ori_ori_n49_), .Y(ori_ori_n294_));
  OAI210     o0266(.A0(ori_ori_n270_), .A1(ori_ori_n290_), .B0(ori_ori_n294_), .Y(ori_ori_n295_));
  NAi21      o0267(.An(l), .B(k), .Y(ori_ori_n296_));
  NO2        o0268(.A(ori_ori_n296_), .B(ori_ori_n49_), .Y(ori_ori_n297_));
  NOi21      o0269(.An(l), .B(j), .Y(ori_ori_n298_));
  NA2        o0270(.A(ori_ori_n167_), .B(ori_ori_n298_), .Y(ori_ori_n299_));
  NA3        o0271(.A(ori_ori_n120_), .B(ori_ori_n119_), .C(g), .Y(ori_ori_n300_));
  OR3        o0272(.A(ori_ori_n72_), .B(ori_ori_n73_), .C(e), .Y(ori_ori_n301_));
  AOI210     o0273(.A0(ori_ori_n300_), .A1(ori_ori_n299_), .B0(ori_ori_n301_), .Y(ori_ori_n302_));
  INV        o0274(.A(ori_ori_n302_), .Y(ori_ori_n303_));
  NAi32      o0275(.An(j), .Bn(h), .C(i), .Y(ori_ori_n304_));
  NAi21      o0276(.An(m), .B(l), .Y(ori_ori_n305_));
  NO3        o0277(.A(ori_ori_n305_), .B(ori_ori_n304_), .C(ori_ori_n84_), .Y(ori_ori_n306_));
  NA2        o0278(.A(h), .B(g), .Y(ori_ori_n307_));
  NA2        o0279(.A(ori_ori_n172_), .B(ori_ori_n45_), .Y(ori_ori_n308_));
  NO2        o0280(.A(ori_ori_n308_), .B(ori_ori_n307_), .Y(ori_ori_n309_));
  NA2        o0281(.A(ori_ori_n309_), .B(ori_ori_n168_), .Y(ori_ori_n310_));
  NA4        o0282(.A(ori_ori_n310_), .B(ori_ori_n303_), .C(ori_ori_n295_), .D(ori_ori_n288_), .Y(ori_ori_n311_));
  NO2        o0283(.A(ori_ori_n148_), .B(d), .Y(ori_ori_n312_));
  NA2        o0284(.A(ori_ori_n312_), .B(ori_ori_n53_), .Y(ori_ori_n313_));
  NO2        o0285(.A(ori_ori_n107_), .B(ori_ori_n104_), .Y(ori_ori_n314_));
  NAi32      o0286(.An(n), .Bn(m), .C(l), .Y(ori_ori_n315_));
  NO2        o0287(.A(ori_ori_n315_), .B(ori_ori_n304_), .Y(ori_ori_n316_));
  NA2        o0288(.A(ori_ori_n316_), .B(ori_ori_n188_), .Y(ori_ori_n317_));
  NO2        o0289(.A(ori_ori_n124_), .B(ori_ori_n118_), .Y(ori_ori_n318_));
  NAi31      o0290(.An(k), .B(l), .C(j), .Y(ori_ori_n319_));
  OAI210     o0291(.A0(ori_ori_n296_), .A1(j), .B0(ori_ori_n319_), .Y(ori_ori_n320_));
  NOi21      o0292(.An(ori_ori_n320_), .B(ori_ori_n122_), .Y(ori_ori_n321_));
  NA2        o0293(.A(ori_ori_n321_), .B(ori_ori_n318_), .Y(ori_ori_n322_));
  NA3        o0294(.A(ori_ori_n322_), .B(ori_ori_n317_), .C(ori_ori_n313_), .Y(ori_ori_n323_));
  NO4        o0295(.A(ori_ori_n323_), .B(ori_ori_n311_), .C(ori_ori_n284_), .D(ori_ori_n277_), .Y(ori_ori_n324_));
  NA2        o0296(.A(ori_ori_n260_), .B(ori_ori_n197_), .Y(ori_ori_n325_));
  NAi21      o0297(.An(m), .B(k), .Y(ori_ori_n326_));
  NO2        o0298(.A(ori_ori_n231_), .B(ori_ori_n326_), .Y(ori_ori_n327_));
  NAi41      o0299(.An(d), .B(n), .C(c), .D(b), .Y(ori_ori_n328_));
  NO2        o0300(.A(ori_ori_n328_), .B(ori_ori_n154_), .Y(ori_ori_n329_));
  NA2        o0301(.A(ori_ori_n329_), .B(ori_ori_n327_), .Y(ori_ori_n330_));
  NA2        o0302(.A(e), .B(c), .Y(ori_ori_n331_));
  NO3        o0303(.A(ori_ori_n331_), .B(n), .C(d), .Y(ori_ori_n332_));
  NOi21      o0304(.An(f), .B(h), .Y(ori_ori_n333_));
  NA2        o0305(.A(ori_ori_n333_), .B(ori_ori_n120_), .Y(ori_ori_n334_));
  NO2        o0306(.A(ori_ori_n334_), .B(ori_ori_n219_), .Y(ori_ori_n335_));
  NAi31      o0307(.An(d), .B(e), .C(b), .Y(ori_ori_n336_));
  NO2        o0308(.A(ori_ori_n134_), .B(ori_ori_n336_), .Y(ori_ori_n337_));
  NA2        o0309(.A(ori_ori_n337_), .B(ori_ori_n335_), .Y(ori_ori_n338_));
  NA3        o0310(.A(ori_ori_n338_), .B(ori_ori_n330_), .C(ori_ori_n325_), .Y(ori_ori_n339_));
  NO4        o0311(.A(ori_ori_n328_), .B(ori_ori_n79_), .C(ori_ori_n71_), .D(ori_ori_n219_), .Y(ori_ori_n340_));
  NA2        o0312(.A(ori_ori_n255_), .B(ori_ori_n105_), .Y(ori_ori_n341_));
  OR2        o0313(.A(ori_ori_n341_), .B(ori_ori_n209_), .Y(ori_ori_n342_));
  NOi31      o0314(.An(l), .B(n), .C(m), .Y(ori_ori_n343_));
  NA2        o0315(.A(ori_ori_n343_), .B(ori_ori_n220_), .Y(ori_ori_n344_));
  NO2        o0316(.A(ori_ori_n344_), .B(ori_ori_n198_), .Y(ori_ori_n345_));
  NAi32      o0317(.An(ori_ori_n345_), .Bn(ori_ori_n340_), .C(ori_ori_n342_), .Y(ori_ori_n346_));
  NAi32      o0318(.An(m), .Bn(j), .C(k), .Y(ori_ori_n347_));
  NAi41      o0319(.An(c), .B(n), .C(d), .D(b), .Y(ori_ori_n348_));
  OAI210     o0320(.A0(ori_ori_n216_), .A1(ori_ori_n347_), .B0(ori_ori_n348_), .Y(ori_ori_n349_));
  NOi31      o0321(.An(j), .B(m), .C(k), .Y(ori_ori_n350_));
  NO2        o0322(.A(ori_ori_n127_), .B(ori_ori_n350_), .Y(ori_ori_n351_));
  AN3        o0323(.A(h), .B(g), .C(f), .Y(ori_ori_n352_));
  NAi31      o0324(.An(ori_ori_n351_), .B(ori_ori_n352_), .C(ori_ori_n349_), .Y(ori_ori_n353_));
  NOi32      o0325(.An(m), .Bn(j), .C(l), .Y(ori_ori_n354_));
  NO2        o0326(.A(ori_ori_n354_), .B(ori_ori_n98_), .Y(ori_ori_n355_));
  NO2        o0327(.A(ori_ori_n305_), .B(ori_ori_n304_), .Y(ori_ori_n356_));
  NO2        o0328(.A(ori_ori_n222_), .B(g), .Y(ori_ori_n357_));
  NO2        o0329(.A(ori_ori_n160_), .B(ori_ori_n84_), .Y(ori_ori_n358_));
  AOI220     o0330(.A0(ori_ori_n358_), .A1(ori_ori_n357_), .B0(ori_ori_n252_), .B1(ori_ori_n356_), .Y(ori_ori_n359_));
  NA2        o0331(.A(ori_ori_n239_), .B(ori_ori_n79_), .Y(ori_ori_n360_));
  NA3        o0332(.A(ori_ori_n360_), .B(ori_ori_n352_), .C(ori_ori_n217_), .Y(ori_ori_n361_));
  NA3        o0333(.A(ori_ori_n361_), .B(ori_ori_n359_), .C(ori_ori_n353_), .Y(ori_ori_n362_));
  NA3        o0334(.A(h), .B(g), .C(f), .Y(ori_ori_n363_));
  NO2        o0335(.A(ori_ori_n363_), .B(ori_ori_n75_), .Y(ori_ori_n364_));
  NA2        o0336(.A(ori_ori_n348_), .B(ori_ori_n216_), .Y(ori_ori_n365_));
  NA2        o0337(.A(ori_ori_n167_), .B(e), .Y(ori_ori_n366_));
  NO2        o0338(.A(ori_ori_n366_), .B(ori_ori_n41_), .Y(ori_ori_n367_));
  AOI220     o0339(.A0(ori_ori_n367_), .A1(ori_ori_n318_), .B0(ori_ori_n365_), .B1(ori_ori_n364_), .Y(ori_ori_n368_));
  NOi32      o0340(.An(j), .Bn(g), .C(i), .Y(ori_ori_n369_));
  NA3        o0341(.A(ori_ori_n369_), .B(ori_ori_n296_), .C(ori_ori_n115_), .Y(ori_ori_n370_));
  AO210      o0342(.A0(ori_ori_n113_), .A1(ori_ori_n32_), .B0(ori_ori_n370_), .Y(ori_ori_n371_));
  NOi32      o0343(.An(e), .Bn(b), .C(a), .Y(ori_ori_n372_));
  AN2        o0344(.A(l), .B(j), .Y(ori_ori_n373_));
  NO2        o0345(.A(ori_ori_n326_), .B(ori_ori_n373_), .Y(ori_ori_n374_));
  NO3        o0346(.A(ori_ori_n328_), .B(ori_ori_n71_), .C(ori_ori_n219_), .Y(ori_ori_n375_));
  NA3        o0347(.A(ori_ori_n214_), .B(ori_ori_n212_), .C(ori_ori_n35_), .Y(ori_ori_n376_));
  AOI220     o0348(.A0(ori_ori_n376_), .A1(ori_ori_n372_), .B0(ori_ori_n375_), .B1(ori_ori_n374_), .Y(ori_ori_n377_));
  NO2        o0349(.A(ori_ori_n336_), .B(n), .Y(ori_ori_n378_));
  NA2        o0350(.A(ori_ori_n213_), .B(k), .Y(ori_ori_n379_));
  NA3        o0351(.A(m), .B(ori_ori_n114_), .C(ori_ori_n218_), .Y(ori_ori_n380_));
  NA4        o0352(.A(ori_ori_n208_), .B(ori_ori_n87_), .C(g), .D(ori_ori_n218_), .Y(ori_ori_n381_));
  OAI210     o0353(.A0(ori_ori_n380_), .A1(ori_ori_n379_), .B0(ori_ori_n381_), .Y(ori_ori_n382_));
  NAi41      o0354(.An(d), .B(e), .C(c), .D(a), .Y(ori_ori_n383_));
  NA2        o0355(.A(ori_ori_n51_), .B(ori_ori_n115_), .Y(ori_ori_n384_));
  NO2        o0356(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n385_));
  AOI220     o0357(.A0(ori_ori_n385_), .A1(b), .B0(ori_ori_n382_), .B1(ori_ori_n378_), .Y(ori_ori_n386_));
  NA4        o0358(.A(ori_ori_n386_), .B(ori_ori_n377_), .C(ori_ori_n371_), .D(ori_ori_n368_), .Y(ori_ori_n387_));
  NO4        o0359(.A(ori_ori_n387_), .B(ori_ori_n362_), .C(ori_ori_n346_), .D(ori_ori_n339_), .Y(ori_ori_n388_));
  NA4        o0360(.A(ori_ori_n388_), .B(ori_ori_n324_), .C(ori_ori_n275_), .D(ori_ori_n204_), .Y(ori10));
  NA3        o0361(.A(m), .B(k), .C(i), .Y(ori_ori_n390_));
  NO3        o0362(.A(ori_ori_n390_), .B(j), .C(ori_ori_n219_), .Y(ori_ori_n391_));
  NOi21      o0363(.An(e), .B(f), .Y(ori_ori_n392_));
  NO4        o0364(.A(ori_ori_n155_), .B(ori_ori_n392_), .C(n), .D(ori_ori_n112_), .Y(ori_ori_n393_));
  NAi31      o0365(.An(b), .B(f), .C(c), .Y(ori_ori_n394_));
  INV        o0366(.A(ori_ori_n394_), .Y(ori_ori_n395_));
  NOi32      o0367(.An(k), .Bn(h), .C(j), .Y(ori_ori_n396_));
  NA2        o0368(.A(ori_ori_n396_), .B(ori_ori_n226_), .Y(ori_ori_n397_));
  NA2        o0369(.A(ori_ori_n165_), .B(ori_ori_n397_), .Y(ori_ori_n398_));
  AOI220     o0370(.A0(ori_ori_n398_), .A1(ori_ori_n395_), .B0(ori_ori_n393_), .B1(ori_ori_n391_), .Y(ori_ori_n399_));
  AN2        o0371(.A(j), .B(h), .Y(ori_ori_n400_));
  NO3        o0372(.A(n), .B(m), .C(k), .Y(ori_ori_n401_));
  NA2        o0373(.A(ori_ori_n401_), .B(ori_ori_n400_), .Y(ori_ori_n402_));
  NO3        o0374(.A(ori_ori_n402_), .B(ori_ori_n155_), .C(ori_ori_n218_), .Y(ori_ori_n403_));
  OR2        o0375(.A(m), .B(k), .Y(ori_ori_n404_));
  NO2        o0376(.A(ori_ori_n178_), .B(ori_ori_n404_), .Y(ori_ori_n405_));
  NA4        o0377(.A(n), .B(f), .C(c), .D(ori_ori_n118_), .Y(ori_ori_n406_));
  NOi21      o0378(.An(ori_ori_n405_), .B(ori_ori_n406_), .Y(ori_ori_n407_));
  NOi32      o0379(.An(d), .Bn(a), .C(c), .Y(ori_ori_n408_));
  NA2        o0380(.A(ori_ori_n408_), .B(ori_ori_n186_), .Y(ori_ori_n409_));
  NAi21      o0381(.An(i), .B(g), .Y(ori_ori_n410_));
  NAi31      o0382(.An(k), .B(m), .C(j), .Y(ori_ori_n411_));
  NO3        o0383(.A(ori_ori_n411_), .B(ori_ori_n410_), .C(n), .Y(ori_ori_n412_));
  NOi21      o0384(.An(ori_ori_n412_), .B(ori_ori_n409_), .Y(ori_ori_n413_));
  NO3        o0385(.A(ori_ori_n413_), .B(ori_ori_n407_), .C(ori_ori_n403_), .Y(ori_ori_n414_));
  NO2        o0386(.A(ori_ori_n406_), .B(ori_ori_n305_), .Y(ori_ori_n415_));
  NOi32      o0387(.An(f), .Bn(d), .C(c), .Y(ori_ori_n416_));
  AOI220     o0388(.A0(ori_ori_n416_), .A1(ori_ori_n316_), .B0(ori_ori_n415_), .B1(ori_ori_n220_), .Y(ori_ori_n417_));
  NA3        o0389(.A(ori_ori_n417_), .B(ori_ori_n414_), .C(ori_ori_n399_), .Y(ori_ori_n418_));
  NO2        o0390(.A(ori_ori_n59_), .B(ori_ori_n118_), .Y(ori_ori_n419_));
  NA2        o0391(.A(ori_ori_n255_), .B(ori_ori_n419_), .Y(ori_ori_n420_));
  INV        o0392(.A(e), .Y(ori_ori_n421_));
  NA2        o0393(.A(ori_ori_n46_), .B(e), .Y(ori_ori_n422_));
  OAI220     o0394(.A0(ori_ori_n422_), .A1(ori_ori_n205_), .B0(ori_ori_n209_), .B1(ori_ori_n421_), .Y(ori_ori_n423_));
  AN2        o0395(.A(g), .B(e), .Y(ori_ori_n424_));
  NA3        o0396(.A(ori_ori_n424_), .B(ori_ori_n208_), .C(i), .Y(ori_ori_n425_));
  OAI210     o0397(.A0(ori_ori_n89_), .A1(ori_ori_n421_), .B0(ori_ori_n425_), .Y(ori_ori_n426_));
  NO2        o0398(.A(ori_ori_n101_), .B(ori_ori_n421_), .Y(ori_ori_n427_));
  NO3        o0399(.A(ori_ori_n427_), .B(ori_ori_n426_), .C(ori_ori_n423_), .Y(ori_ori_n428_));
  NOi32      o0400(.An(h), .Bn(e), .C(g), .Y(ori_ori_n429_));
  NA3        o0401(.A(ori_ori_n429_), .B(ori_ori_n298_), .C(m), .Y(ori_ori_n430_));
  NOi21      o0402(.An(g), .B(h), .Y(ori_ori_n431_));
  AN3        o0403(.A(m), .B(l), .C(i), .Y(ori_ori_n432_));
  NA3        o0404(.A(ori_ori_n432_), .B(ori_ori_n431_), .C(e), .Y(ori_ori_n433_));
  AN3        o0405(.A(h), .B(g), .C(e), .Y(ori_ori_n434_));
  NA2        o0406(.A(ori_ori_n434_), .B(ori_ori_n98_), .Y(ori_ori_n435_));
  AN3        o0407(.A(ori_ori_n435_), .B(ori_ori_n433_), .C(ori_ori_n430_), .Y(ori_ori_n436_));
  AOI210     o0408(.A0(ori_ori_n436_), .A1(ori_ori_n428_), .B0(ori_ori_n420_), .Y(ori_ori_n437_));
  NA3        o0409(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(e), .Y(ori_ori_n438_));
  NO2        o0410(.A(ori_ori_n438_), .B(ori_ori_n420_), .Y(ori_ori_n439_));
  NA3        o0411(.A(ori_ori_n408_), .B(ori_ori_n186_), .C(ori_ori_n84_), .Y(ori_ori_n440_));
  NAi31      o0412(.An(b), .B(c), .C(a), .Y(ori_ori_n441_));
  NO2        o0413(.A(ori_ori_n441_), .B(n), .Y(ori_ori_n442_));
  NA2        o0414(.A(ori_ori_n51_), .B(m), .Y(ori_ori_n443_));
  NO2        o0415(.A(ori_ori_n443_), .B(ori_ori_n151_), .Y(ori_ori_n444_));
  NA2        o0416(.A(ori_ori_n444_), .B(ori_ori_n442_), .Y(ori_ori_n445_));
  INV        o0417(.A(ori_ori_n445_), .Y(ori_ori_n446_));
  NO4        o0418(.A(ori_ori_n446_), .B(ori_ori_n439_), .C(ori_ori_n437_), .D(ori_ori_n418_), .Y(ori_ori_n447_));
  NA2        o0419(.A(i), .B(g), .Y(ori_ori_n448_));
  NOi21      o0420(.An(a), .B(n), .Y(ori_ori_n449_));
  NOi21      o0421(.An(d), .B(c), .Y(ori_ori_n450_));
  NA2        o0422(.A(ori_ori_n450_), .B(ori_ori_n449_), .Y(ori_ori_n451_));
  NA3        o0423(.A(i), .B(g), .C(f), .Y(ori_ori_n452_));
  OR2        o0424(.A(ori_ori_n452_), .B(ori_ori_n70_), .Y(ori_ori_n453_));
  NA3        o0425(.A(ori_ori_n432_), .B(ori_ori_n431_), .C(ori_ori_n186_), .Y(ori_ori_n454_));
  AOI210     o0426(.A0(ori_ori_n454_), .A1(ori_ori_n453_), .B0(ori_ori_n451_), .Y(ori_ori_n455_));
  INV        o0427(.A(ori_ori_n455_), .Y(ori_ori_n456_));
  OR2        o0428(.A(n), .B(m), .Y(ori_ori_n457_));
  NO2        o0429(.A(ori_ori_n457_), .B(ori_ori_n156_), .Y(ori_ori_n458_));
  NO2        o0430(.A(ori_ori_n187_), .B(ori_ori_n151_), .Y(ori_ori_n459_));
  OAI210     o0431(.A0(ori_ori_n458_), .A1(ori_ori_n180_), .B0(ori_ori_n459_), .Y(ori_ori_n460_));
  INV        o0432(.A(ori_ori_n384_), .Y(ori_ori_n461_));
  NA3        o0433(.A(ori_ori_n461_), .B(ori_ori_n372_), .C(d), .Y(ori_ori_n462_));
  NO2        o0434(.A(ori_ori_n441_), .B(ori_ori_n49_), .Y(ori_ori_n463_));
  NO3        o0435(.A(ori_ori_n66_), .B(ori_ori_n114_), .C(e), .Y(ori_ori_n464_));
  NAi21      o0436(.An(k), .B(j), .Y(ori_ori_n465_));
  NA2        o0437(.A(ori_ori_n258_), .B(ori_ori_n465_), .Y(ori_ori_n466_));
  NA3        o0438(.A(ori_ori_n466_), .B(ori_ori_n464_), .C(ori_ori_n463_), .Y(ori_ori_n467_));
  NAi21      o0439(.An(e), .B(d), .Y(ori_ori_n468_));
  INV        o0440(.A(ori_ori_n468_), .Y(ori_ori_n469_));
  NO2        o0441(.A(ori_ori_n259_), .B(ori_ori_n218_), .Y(ori_ori_n470_));
  NA3        o0442(.A(ori_ori_n470_), .B(ori_ori_n469_), .C(ori_ori_n232_), .Y(ori_ori_n471_));
  NA4        o0443(.A(ori_ori_n471_), .B(ori_ori_n467_), .C(ori_ori_n462_), .D(ori_ori_n460_), .Y(ori_ori_n472_));
  NO2        o0444(.A(ori_ori_n344_), .B(ori_ori_n218_), .Y(ori_ori_n473_));
  NA2        o0445(.A(ori_ori_n473_), .B(ori_ori_n469_), .Y(ori_ori_n474_));
  NOi31      o0446(.An(n), .B(m), .C(k), .Y(ori_ori_n475_));
  AOI220     o0447(.A0(ori_ori_n475_), .A1(ori_ori_n400_), .B0(ori_ori_n226_), .B1(ori_ori_n50_), .Y(ori_ori_n476_));
  NAi31      o0448(.An(g), .B(f), .C(c), .Y(ori_ori_n477_));
  OR3        o0449(.A(ori_ori_n477_), .B(ori_ori_n476_), .C(e), .Y(ori_ori_n478_));
  NA3        o0450(.A(ori_ori_n478_), .B(ori_ori_n474_), .C(ori_ori_n317_), .Y(ori_ori_n479_));
  NOi41      o0451(.An(ori_ori_n456_), .B(ori_ori_n479_), .C(ori_ori_n472_), .D(ori_ori_n273_), .Y(ori_ori_n480_));
  NOi32      o0452(.An(c), .Bn(a), .C(b), .Y(ori_ori_n481_));
  NA2        o0453(.A(ori_ori_n481_), .B(ori_ori_n115_), .Y(ori_ori_n482_));
  INV        o0454(.A(ori_ori_n282_), .Y(ori_ori_n483_));
  AN2        o0455(.A(e), .B(d), .Y(ori_ori_n484_));
  NA2        o0456(.A(ori_ori_n484_), .B(ori_ori_n483_), .Y(ori_ori_n485_));
  INV        o0457(.A(ori_ori_n151_), .Y(ori_ori_n486_));
  NO2        o0458(.A(ori_ori_n133_), .B(ori_ori_n41_), .Y(ori_ori_n487_));
  NO2        o0459(.A(ori_ori_n66_), .B(e), .Y(ori_ori_n488_));
  NOi31      o0460(.An(j), .B(k), .C(i), .Y(ori_ori_n489_));
  NOi21      o0461(.An(ori_ori_n169_), .B(ori_ori_n489_), .Y(ori_ori_n490_));
  NA3        o0462(.A(ori_ori_n490_), .B(ori_ori_n267_), .C(ori_ori_n121_), .Y(ori_ori_n491_));
  AOI220     o0463(.A0(ori_ori_n491_), .A1(ori_ori_n488_), .B0(ori_ori_n487_), .B1(ori_ori_n486_), .Y(ori_ori_n492_));
  AOI210     o0464(.A0(ori_ori_n492_), .A1(ori_ori_n485_), .B0(ori_ori_n482_), .Y(ori_ori_n493_));
  INV        o0465(.A(ori_ori_n210_), .Y(ori_ori_n494_));
  NOi21      o0466(.An(a), .B(b), .Y(ori_ori_n495_));
  NA3        o0467(.A(e), .B(d), .C(c), .Y(ori_ori_n496_));
  NAi21      o0468(.An(ori_ori_n496_), .B(ori_ori_n495_), .Y(ori_ori_n497_));
  NO2        o0469(.A(ori_ori_n440_), .B(ori_ori_n209_), .Y(ori_ori_n498_));
  NOi21      o0470(.An(ori_ori_n497_), .B(ori_ori_n498_), .Y(ori_ori_n499_));
  AOI210     o0471(.A0(ori_ori_n276_), .A1(ori_ori_n494_), .B0(ori_ori_n499_), .Y(ori_ori_n500_));
  NO4        o0472(.A(ori_ori_n192_), .B(ori_ori_n104_), .C(ori_ori_n56_), .D(b), .Y(ori_ori_n501_));
  NA2        o0473(.A(ori_ori_n395_), .B(ori_ori_n157_), .Y(ori_ori_n502_));
  OR2        o0474(.A(k), .B(j), .Y(ori_ori_n503_));
  NA2        o0475(.A(l), .B(k), .Y(ori_ori_n504_));
  NA3        o0476(.A(ori_ori_n504_), .B(ori_ori_n503_), .C(ori_ori_n226_), .Y(ori_ori_n505_));
  AOI210     o0477(.A0(ori_ori_n239_), .A1(ori_ori_n347_), .B0(ori_ori_n84_), .Y(ori_ori_n506_));
  NOi21      o0478(.An(ori_ori_n505_), .B(ori_ori_n506_), .Y(ori_ori_n507_));
  OR3        o0479(.A(ori_ori_n507_), .B(ori_ori_n147_), .C(ori_ori_n137_), .Y(ori_ori_n508_));
  NA3        o0480(.A(ori_ori_n285_), .B(ori_ori_n130_), .C(ori_ori_n128_), .Y(ori_ori_n509_));
  NO3        o0481(.A(ori_ori_n440_), .B(ori_ori_n92_), .C(ori_ori_n133_), .Y(ori_ori_n510_));
  NO2        o0482(.A(ori_ori_n510_), .B(ori_ori_n509_), .Y(ori_ori_n511_));
  NA3        o0483(.A(ori_ori_n511_), .B(ori_ori_n508_), .C(ori_ori_n502_), .Y(ori_ori_n512_));
  NO4        o0484(.A(ori_ori_n512_), .B(ori_ori_n501_), .C(ori_ori_n500_), .D(ori_ori_n493_), .Y(ori_ori_n513_));
  INV        o0485(.A(e), .Y(ori_ori_n514_));
  NO2        o0486(.A(ori_ori_n192_), .B(ori_ori_n56_), .Y(ori_ori_n515_));
  NAi31      o0487(.An(j), .B(l), .C(i), .Y(ori_ori_n516_));
  OAI210     o0488(.A0(ori_ori_n516_), .A1(ori_ori_n134_), .B0(ori_ori_n104_), .Y(ori_ori_n517_));
  NA4        o0489(.A(ori_ori_n517_), .B(ori_ori_n515_), .C(ori_ori_n514_), .D(b), .Y(ori_ori_n518_));
  NO3        o0490(.A(ori_ori_n409_), .B(ori_ori_n355_), .C(ori_ori_n206_), .Y(ori_ori_n519_));
  NO2        o0491(.A(ori_ori_n409_), .B(ori_ori_n384_), .Y(ori_ori_n520_));
  NO4        o0492(.A(ori_ori_n520_), .B(ori_ori_n519_), .C(ori_ori_n189_), .D(ori_ori_n314_), .Y(ori_ori_n521_));
  NA3        o0493(.A(ori_ori_n521_), .B(ori_ori_n518_), .C(ori_ori_n247_), .Y(ori_ori_n522_));
  OAI210     o0494(.A0(ori_ori_n129_), .A1(ori_ori_n127_), .B0(n), .Y(ori_ori_n523_));
  NO2        o0495(.A(ori_ori_n523_), .B(ori_ori_n133_), .Y(ori_ori_n524_));
  AN2        o0496(.A(ori_ori_n524_), .B(ori_ori_n197_), .Y(ori_ori_n525_));
  XO2        o0497(.A(i), .B(h), .Y(ori_ori_n526_));
  NA3        o0498(.A(ori_ori_n526_), .B(ori_ori_n164_), .C(n), .Y(ori_ori_n527_));
  NAi41      o0499(.An(ori_ori_n306_), .B(ori_ori_n527_), .C(ori_ori_n476_), .D(ori_ori_n397_), .Y(ori_ori_n528_));
  NOi32      o0500(.An(ori_ori_n528_), .Bn(ori_ori_n488_), .C(ori_ori_n278_), .Y(ori_ori_n529_));
  NAi31      o0501(.An(c), .B(f), .C(d), .Y(ori_ori_n530_));
  AOI210     o0502(.A0(ori_ori_n286_), .A1(ori_ori_n200_), .B0(ori_ori_n530_), .Y(ori_ori_n531_));
  NOi21      o0503(.An(ori_ori_n82_), .B(ori_ori_n531_), .Y(ori_ori_n532_));
  NA3        o0504(.A(ori_ori_n393_), .B(ori_ori_n98_), .C(ori_ori_n97_), .Y(ori_ori_n533_));
  NA2        o0505(.A(ori_ori_n233_), .B(ori_ori_n110_), .Y(ori_ori_n534_));
  AOI210     o0506(.A0(ori_ori_n534_), .A1(ori_ori_n185_), .B0(ori_ori_n530_), .Y(ori_ori_n535_));
  AOI210     o0507(.A0(ori_ori_n370_), .A1(ori_ori_n35_), .B0(ori_ori_n497_), .Y(ori_ori_n536_));
  NOi31      o0508(.An(ori_ori_n533_), .B(ori_ori_n536_), .C(ori_ori_n535_), .Y(ori_ori_n537_));
  AO220      o0509(.A0(ori_ori_n294_), .A1(ori_ori_n270_), .B0(ori_ori_n170_), .B1(ori_ori_n67_), .Y(ori_ori_n538_));
  NA3        o0510(.A(ori_ori_n37_), .B(ori_ori_n36_), .C(f), .Y(ori_ori_n539_));
  INV        o0511(.A(ori_ori_n302_), .Y(ori_ori_n540_));
  NAi41      o0512(.An(ori_ori_n538_), .B(ori_ori_n540_), .C(ori_ori_n537_), .D(ori_ori_n532_), .Y(ori_ori_n541_));
  NO4        o0513(.A(ori_ori_n541_), .B(ori_ori_n529_), .C(ori_ori_n525_), .D(ori_ori_n522_), .Y(ori_ori_n542_));
  NA4        o0514(.A(ori_ori_n542_), .B(ori_ori_n513_), .C(ori_ori_n480_), .D(ori_ori_n447_), .Y(ori11));
  NO2        o0515(.A(ori_ori_n72_), .B(f), .Y(ori_ori_n544_));
  NA2        o0516(.A(j), .B(g), .Y(ori_ori_n545_));
  NAi31      o0517(.An(i), .B(m), .C(l), .Y(ori_ori_n546_));
  NA3        o0518(.A(m), .B(k), .C(j), .Y(ori_ori_n547_));
  OAI220     o0519(.A0(ori_ori_n547_), .A1(ori_ori_n133_), .B0(ori_ori_n546_), .B1(ori_ori_n545_), .Y(ori_ori_n548_));
  NA2        o0520(.A(ori_ori_n548_), .B(ori_ori_n544_), .Y(ori_ori_n549_));
  NOi32      o0521(.An(e), .Bn(b), .C(f), .Y(ori_ori_n550_));
  NA2        o0522(.A(ori_ori_n46_), .B(j), .Y(ori_ori_n551_));
  NO2        o0523(.A(ori_ori_n551_), .B(ori_ori_n308_), .Y(ori_ori_n552_));
  NAi31      o0524(.An(d), .B(e), .C(a), .Y(ori_ori_n553_));
  NO2        o0525(.A(ori_ori_n553_), .B(n), .Y(ori_ori_n554_));
  AOI220     o0526(.A0(ori_ori_n554_), .A1(ori_ori_n102_), .B0(ori_ori_n552_), .B1(ori_ori_n550_), .Y(ori_ori_n555_));
  NAi41      o0527(.An(f), .B(e), .C(c), .D(a), .Y(ori_ori_n556_));
  AN2        o0528(.A(ori_ori_n556_), .B(ori_ori_n383_), .Y(ori_ori_n557_));
  NA2        o0529(.A(j), .B(i), .Y(ori_ori_n558_));
  NAi31      o0530(.An(n), .B(m), .C(k), .Y(ori_ori_n559_));
  NO3        o0531(.A(ori_ori_n559_), .B(ori_ori_n558_), .C(ori_ori_n114_), .Y(ori_ori_n560_));
  NO4        o0532(.A(n), .B(d), .C(ori_ori_n118_), .D(a), .Y(ori_ori_n561_));
  OR2        o0533(.A(n), .B(c), .Y(ori_ori_n562_));
  NO2        o0534(.A(ori_ori_n562_), .B(ori_ori_n153_), .Y(ori_ori_n563_));
  NO2        o0535(.A(ori_ori_n563_), .B(ori_ori_n561_), .Y(ori_ori_n564_));
  NOi32      o0536(.An(g), .Bn(f), .C(i), .Y(ori_ori_n565_));
  AOI220     o0537(.A0(ori_ori_n565_), .A1(ori_ori_n100_), .B0(ori_ori_n548_), .B1(f), .Y(ori_ori_n566_));
  NO2        o0538(.A(ori_ori_n282_), .B(ori_ori_n49_), .Y(ori_ori_n567_));
  NO2        o0539(.A(ori_ori_n566_), .B(ori_ori_n564_), .Y(ori_ori_n568_));
  INV        o0540(.A(ori_ori_n568_), .Y(ori_ori_n569_));
  NA2        o0541(.A(ori_ori_n143_), .B(ori_ori_n34_), .Y(ori_ori_n570_));
  OAI220     o0542(.A0(ori_ori_n570_), .A1(m), .B0(ori_ori_n551_), .B1(ori_ori_n239_), .Y(ori_ori_n571_));
  NOi41      o0543(.An(d), .B(n), .C(e), .D(c), .Y(ori_ori_n572_));
  NAi32      o0544(.An(e), .Bn(b), .C(c), .Y(ori_ori_n573_));
  OR2        o0545(.A(ori_ori_n573_), .B(ori_ori_n84_), .Y(ori_ori_n574_));
  AN2        o0546(.A(ori_ori_n348_), .B(ori_ori_n328_), .Y(ori_ori_n575_));
  NA2        o0547(.A(ori_ori_n575_), .B(ori_ori_n574_), .Y(ori_ori_n576_));
  OA210      o0548(.A0(ori_ori_n576_), .A1(ori_ori_n572_), .B0(ori_ori_n571_), .Y(ori_ori_n577_));
  OAI220     o0549(.A0(ori_ori_n411_), .A1(ori_ori_n410_), .B0(ori_ori_n546_), .B1(ori_ori_n545_), .Y(ori_ori_n578_));
  NAi31      o0550(.An(d), .B(c), .C(a), .Y(ori_ori_n579_));
  NO2        o0551(.A(ori_ori_n579_), .B(n), .Y(ori_ori_n580_));
  NA3        o0552(.A(ori_ori_n580_), .B(ori_ori_n578_), .C(e), .Y(ori_ori_n581_));
  NO3        o0553(.A(ori_ori_n62_), .B(ori_ori_n49_), .C(ori_ori_n219_), .Y(ori_ori_n582_));
  NO2        o0554(.A(ori_ori_n236_), .B(ori_ori_n112_), .Y(ori_ori_n583_));
  OAI210     o0555(.A0(ori_ori_n582_), .A1(ori_ori_n412_), .B0(ori_ori_n583_), .Y(ori_ori_n584_));
  NA2        o0556(.A(ori_ori_n584_), .B(ori_ori_n581_), .Y(ori_ori_n585_));
  NO2        o0557(.A(ori_ori_n283_), .B(n), .Y(ori_ori_n586_));
  NO2        o0558(.A(ori_ori_n442_), .B(ori_ori_n586_), .Y(ori_ori_n587_));
  NA2        o0559(.A(ori_ori_n578_), .B(f), .Y(ori_ori_n588_));
  NAi32      o0560(.An(d), .Bn(a), .C(b), .Y(ori_ori_n589_));
  NO2        o0561(.A(ori_ori_n589_), .B(ori_ori_n49_), .Y(ori_ori_n590_));
  NA2        o0562(.A(h), .B(f), .Y(ori_ori_n591_));
  NO2        o0563(.A(ori_ori_n591_), .B(ori_ori_n95_), .Y(ori_ori_n592_));
  NO3        o0564(.A(ori_ori_n181_), .B(ori_ori_n178_), .C(g), .Y(ori_ori_n593_));
  AOI220     o0565(.A0(ori_ori_n593_), .A1(ori_ori_n58_), .B0(ori_ori_n592_), .B1(ori_ori_n590_), .Y(ori_ori_n594_));
  OAI210     o0566(.A0(ori_ori_n588_), .A1(ori_ori_n587_), .B0(ori_ori_n594_), .Y(ori_ori_n595_));
  AN3        o0567(.A(j), .B(h), .C(g), .Y(ori_ori_n596_));
  NO2        o0568(.A(ori_ori_n150_), .B(c), .Y(ori_ori_n597_));
  NA3        o0569(.A(ori_ori_n597_), .B(ori_ori_n596_), .C(ori_ori_n475_), .Y(ori_ori_n598_));
  NA3        o0570(.A(f), .B(d), .C(b), .Y(ori_ori_n599_));
  NO4        o0571(.A(ori_ori_n599_), .B(ori_ori_n181_), .C(ori_ori_n178_), .D(g), .Y(ori_ori_n600_));
  NAi21      o0572(.An(ori_ori_n600_), .B(ori_ori_n598_), .Y(ori_ori_n601_));
  NO4        o0573(.A(ori_ori_n601_), .B(ori_ori_n595_), .C(ori_ori_n585_), .D(ori_ori_n577_), .Y(ori_ori_n602_));
  AN4        o0574(.A(ori_ori_n602_), .B(ori_ori_n569_), .C(ori_ori_n555_), .D(ori_ori_n549_), .Y(ori_ori_n603_));
  INV        o0575(.A(k), .Y(ori_ori_n604_));
  NA3        o0576(.A(l), .B(ori_ori_n604_), .C(i), .Y(ori_ori_n605_));
  INV        o0577(.A(ori_ori_n605_), .Y(ori_ori_n606_));
  NA4        o0578(.A(ori_ori_n408_), .B(ori_ori_n431_), .C(ori_ori_n186_), .D(ori_ori_n115_), .Y(ori_ori_n607_));
  NAi32      o0579(.An(h), .Bn(f), .C(g), .Y(ori_ori_n608_));
  NAi41      o0580(.An(n), .B(e), .C(c), .D(a), .Y(ori_ori_n609_));
  OAI210     o0581(.A0(ori_ori_n553_), .A1(n), .B0(ori_ori_n609_), .Y(ori_ori_n610_));
  NA2        o0582(.A(ori_ori_n610_), .B(m), .Y(ori_ori_n611_));
  NAi31      o0583(.An(h), .B(g), .C(f), .Y(ori_ori_n612_));
  OR3        o0584(.A(ori_ori_n612_), .B(ori_ori_n283_), .C(ori_ori_n49_), .Y(ori_ori_n613_));
  NA4        o0585(.A(ori_ori_n431_), .B(ori_ori_n123_), .C(ori_ori_n115_), .D(e), .Y(ori_ori_n614_));
  AN2        o0586(.A(ori_ori_n614_), .B(ori_ori_n613_), .Y(ori_ori_n615_));
  OA210      o0587(.A0(ori_ori_n611_), .A1(ori_ori_n608_), .B0(ori_ori_n615_), .Y(ori_ori_n616_));
  NO3        o0588(.A(ori_ori_n608_), .B(ori_ori_n72_), .C(ori_ori_n73_), .Y(ori_ori_n617_));
  NO4        o0589(.A(ori_ori_n612_), .B(ori_ori_n562_), .C(ori_ori_n153_), .D(ori_ori_n73_), .Y(ori_ori_n618_));
  OR2        o0590(.A(ori_ori_n618_), .B(ori_ori_n617_), .Y(ori_ori_n619_));
  NAi31      o0591(.An(ori_ori_n619_), .B(ori_ori_n616_), .C(ori_ori_n607_), .Y(ori_ori_n620_));
  NAi31      o0592(.An(f), .B(h), .C(g), .Y(ori_ori_n621_));
  NOi32      o0593(.An(b), .Bn(a), .C(c), .Y(ori_ori_n622_));
  NOi41      o0594(.An(ori_ori_n622_), .B(ori_ori_n363_), .C(ori_ori_n69_), .D(ori_ori_n119_), .Y(ori_ori_n623_));
  NOi32      o0595(.An(d), .Bn(a), .C(e), .Y(ori_ori_n624_));
  NA2        o0596(.A(ori_ori_n624_), .B(ori_ori_n115_), .Y(ori_ori_n625_));
  NO2        o0597(.A(n), .B(c), .Y(ori_ori_n626_));
  NA3        o0598(.A(ori_ori_n626_), .B(ori_ori_n29_), .C(m), .Y(ori_ori_n627_));
  NAi32      o0599(.An(n), .Bn(f), .C(m), .Y(ori_ori_n628_));
  NA3        o0600(.A(ori_ori_n628_), .B(ori_ori_n627_), .C(ori_ori_n625_), .Y(ori_ori_n629_));
  NOi32      o0601(.An(e), .Bn(a), .C(d), .Y(ori_ori_n630_));
  AOI210     o0602(.A0(ori_ori_n29_), .A1(d), .B0(ori_ori_n630_), .Y(ori_ori_n631_));
  AOI210     o0603(.A0(ori_ori_n631_), .A1(ori_ori_n218_), .B0(ori_ori_n570_), .Y(ori_ori_n632_));
  AOI210     o0604(.A0(ori_ori_n632_), .A1(ori_ori_n629_), .B0(ori_ori_n623_), .Y(ori_ori_n633_));
  OAI210     o0605(.A0(ori_ori_n254_), .A1(ori_ori_n87_), .B0(ori_ori_n633_), .Y(ori_ori_n634_));
  AOI210     o0606(.A0(ori_ori_n620_), .A1(ori_ori_n606_), .B0(ori_ori_n634_), .Y(ori_ori_n635_));
  NO3        o0607(.A(ori_ori_n326_), .B(ori_ori_n61_), .C(n), .Y(ori_ori_n636_));
  NA3        o0608(.A(ori_ori_n530_), .B(ori_ori_n176_), .C(ori_ori_n175_), .Y(ori_ori_n637_));
  NA2        o0609(.A(ori_ori_n477_), .B(ori_ori_n236_), .Y(ori_ori_n638_));
  OR2        o0610(.A(ori_ori_n638_), .B(ori_ori_n637_), .Y(ori_ori_n639_));
  NA2        o0611(.A(ori_ori_n639_), .B(ori_ori_n636_), .Y(ori_ori_n640_));
  NO2        o0612(.A(ori_ori_n640_), .B(ori_ori_n87_), .Y(ori_ori_n641_));
  NA3        o0613(.A(ori_ori_n572_), .B(ori_ori_n350_), .C(ori_ori_n46_), .Y(ori_ori_n642_));
  NOi32      o0614(.An(e), .Bn(c), .C(f), .Y(ori_ori_n643_));
  NOi21      o0615(.An(f), .B(g), .Y(ori_ori_n644_));
  NO2        o0616(.A(ori_ori_n644_), .B(ori_ori_n216_), .Y(ori_ori_n645_));
  AOI220     o0617(.A0(ori_ori_n645_), .A1(ori_ori_n405_), .B0(ori_ori_n643_), .B1(ori_ori_n180_), .Y(ori_ori_n646_));
  NA3        o0618(.A(ori_ori_n646_), .B(ori_ori_n642_), .C(ori_ori_n183_), .Y(ori_ori_n647_));
  AOI210     o0619(.A0(ori_ori_n557_), .A1(ori_ori_n409_), .B0(ori_ori_n307_), .Y(ori_ori_n648_));
  NA2        o0620(.A(ori_ori_n648_), .B(ori_ori_n271_), .Y(ori_ori_n649_));
  NOi21      o0621(.An(j), .B(l), .Y(ori_ori_n650_));
  NAi21      o0622(.An(k), .B(h), .Y(ori_ori_n651_));
  NO2        o0623(.A(ori_ori_n651_), .B(ori_ori_n269_), .Y(ori_ori_n652_));
  NA2        o0624(.A(ori_ori_n652_), .B(ori_ori_n650_), .Y(ori_ori_n653_));
  NOi31      o0625(.An(m), .B(n), .C(k), .Y(ori_ori_n654_));
  NA2        o0626(.A(ori_ori_n650_), .B(ori_ori_n654_), .Y(ori_ori_n655_));
  AOI210     o0627(.A0(ori_ori_n409_), .A1(ori_ori_n383_), .B0(ori_ori_n307_), .Y(ori_ori_n656_));
  NAi21      o0628(.An(ori_ori_n655_), .B(ori_ori_n656_), .Y(ori_ori_n657_));
  NO2        o0629(.A(ori_ori_n283_), .B(ori_ori_n49_), .Y(ori_ori_n658_));
  NO2        o0630(.A(ori_ori_n553_), .B(ori_ori_n49_), .Y(ori_ori_n659_));
  NA2        o0631(.A(ori_ori_n657_), .B(ori_ori_n649_), .Y(ori_ori_n660_));
  NA2        o0632(.A(ori_ori_n110_), .B(ori_ori_n36_), .Y(ori_ori_n661_));
  NO2        o0633(.A(k), .B(ori_ori_n219_), .Y(ori_ori_n662_));
  INV        o0634(.A(ori_ori_n372_), .Y(ori_ori_n663_));
  NO2        o0635(.A(ori_ori_n663_), .B(n), .Y(ori_ori_n664_));
  NAi31      o0636(.An(ori_ori_n661_), .B(ori_ori_n664_), .C(ori_ori_n662_), .Y(ori_ori_n665_));
  NO2        o0637(.A(ori_ori_n551_), .B(ori_ori_n181_), .Y(ori_ori_n666_));
  NA3        o0638(.A(ori_ori_n573_), .B(ori_ori_n278_), .C(ori_ori_n148_), .Y(ori_ori_n667_));
  NA2        o0639(.A(ori_ori_n526_), .B(ori_ori_n164_), .Y(ori_ori_n668_));
  NO3        o0640(.A(ori_ori_n406_), .B(ori_ori_n668_), .C(ori_ori_n87_), .Y(ori_ori_n669_));
  AOI210     o0641(.A0(ori_ori_n667_), .A1(ori_ori_n666_), .B0(ori_ori_n669_), .Y(ori_ori_n670_));
  AN3        o0642(.A(f), .B(d), .C(b), .Y(ori_ori_n671_));
  OAI210     o0643(.A0(ori_ori_n671_), .A1(ori_ori_n132_), .B0(n), .Y(ori_ori_n672_));
  NA3        o0644(.A(ori_ori_n526_), .B(ori_ori_n164_), .C(ori_ori_n219_), .Y(ori_ori_n673_));
  AOI210     o0645(.A0(ori_ori_n672_), .A1(ori_ori_n238_), .B0(ori_ori_n673_), .Y(ori_ori_n674_));
  NAi31      o0646(.An(m), .B(n), .C(k), .Y(ori_ori_n675_));
  INV        o0647(.A(ori_ori_n256_), .Y(ori_ori_n676_));
  OAI210     o0648(.A0(ori_ori_n676_), .A1(ori_ori_n674_), .B0(j), .Y(ori_ori_n677_));
  NA3        o0649(.A(ori_ori_n677_), .B(ori_ori_n670_), .C(ori_ori_n665_), .Y(ori_ori_n678_));
  NO4        o0650(.A(ori_ori_n678_), .B(ori_ori_n660_), .C(ori_ori_n647_), .D(ori_ori_n641_), .Y(ori_ori_n679_));
  NA2        o0651(.A(ori_ori_n393_), .B(ori_ori_n167_), .Y(ori_ori_n680_));
  NAi31      o0652(.An(g), .B(h), .C(f), .Y(ori_ori_n681_));
  OR3        o0653(.A(ori_ori_n681_), .B(ori_ori_n283_), .C(n), .Y(ori_ori_n682_));
  OA210      o0654(.A0(ori_ori_n553_), .A1(n), .B0(ori_ori_n609_), .Y(ori_ori_n683_));
  NA3        o0655(.A(ori_ori_n429_), .B(ori_ori_n123_), .C(ori_ori_n84_), .Y(ori_ori_n684_));
  OAI210     o0656(.A0(ori_ori_n683_), .A1(ori_ori_n91_), .B0(ori_ori_n684_), .Y(ori_ori_n685_));
  NOi21      o0657(.An(ori_ori_n682_), .B(ori_ori_n685_), .Y(ori_ori_n686_));
  AOI210     o0658(.A0(ori_ori_n686_), .A1(ori_ori_n680_), .B0(ori_ori_n547_), .Y(ori_ori_n687_));
  NO3        o0659(.A(g), .B(ori_ori_n218_), .C(ori_ori_n56_), .Y(ori_ori_n688_));
  NAi21      o0660(.An(h), .B(j), .Y(ori_ori_n689_));
  NO2        o0661(.A(ori_ori_n534_), .B(ori_ori_n87_), .Y(ori_ori_n690_));
  OAI210     o0662(.A0(ori_ori_n690_), .A1(ori_ori_n405_), .B0(ori_ori_n688_), .Y(ori_ori_n691_));
  OR2        o0663(.A(ori_ori_n72_), .B(ori_ori_n73_), .Y(ori_ori_n692_));
  NA2        o0664(.A(ori_ori_n622_), .B(ori_ori_n352_), .Y(ori_ori_n693_));
  OA220      o0665(.A0(ori_ori_n655_), .A1(ori_ori_n693_), .B0(ori_ori_n653_), .B1(ori_ori_n692_), .Y(ori_ori_n694_));
  NA3        o0666(.A(ori_ori_n544_), .B(ori_ori_n100_), .C(ori_ori_n99_), .Y(ori_ori_n695_));
  AN2        o0667(.A(h), .B(f), .Y(ori_ori_n696_));
  NA2        o0668(.A(ori_ori_n696_), .B(ori_ori_n37_), .Y(ori_ori_n697_));
  NA2        o0669(.A(ori_ori_n100_), .B(ori_ori_n46_), .Y(ori_ori_n698_));
  OAI220     o0670(.A0(ori_ori_n698_), .A1(ori_ori_n341_), .B0(ori_ori_n697_), .B1(ori_ori_n482_), .Y(ori_ori_n699_));
  AOI210     o0671(.A0(ori_ori_n589_), .A1(ori_ori_n441_), .B0(ori_ori_n49_), .Y(ori_ori_n700_));
  OAI220     o0672(.A0(ori_ori_n612_), .A1(ori_ori_n605_), .B0(ori_ori_n334_), .B1(ori_ori_n545_), .Y(ori_ori_n701_));
  AOI210     o0673(.A0(ori_ori_n701_), .A1(ori_ori_n700_), .B0(ori_ori_n699_), .Y(ori_ori_n702_));
  NA4        o0674(.A(ori_ori_n702_), .B(ori_ori_n695_), .C(ori_ori_n694_), .D(ori_ori_n691_), .Y(ori_ori_n703_));
  NO2        o0675(.A(ori_ori_n644_), .B(ori_ori_n61_), .Y(ori_ori_n704_));
  NO2        o0676(.A(ori_ori_n704_), .B(ori_ori_n34_), .Y(ori_ori_n705_));
  NA2        o0677(.A(ori_ori_n337_), .B(ori_ori_n143_), .Y(ori_ori_n706_));
  NA2        o0678(.A(ori_ori_n134_), .B(ori_ori_n49_), .Y(ori_ori_n707_));
  AOI220     o0679(.A0(ori_ori_n707_), .A1(ori_ori_n550_), .B0(ori_ori_n372_), .B1(ori_ori_n115_), .Y(ori_ori_n708_));
  OA220      o0680(.A0(ori_ori_n708_), .A1(ori_ori_n570_), .B0(ori_ori_n370_), .B1(ori_ori_n113_), .Y(ori_ori_n709_));
  OAI210     o0681(.A0(ori_ori_n706_), .A1(ori_ori_n705_), .B0(ori_ori_n709_), .Y(ori_ori_n710_));
  NO3        o0682(.A(ori_ori_n416_), .B(ori_ori_n197_), .C(ori_ori_n196_), .Y(ori_ori_n711_));
  NA2        o0683(.A(ori_ori_n711_), .B(ori_ori_n236_), .Y(ori_ori_n712_));
  NA3        o0684(.A(ori_ori_n712_), .B(ori_ori_n260_), .C(j), .Y(ori_ori_n713_));
  NO3        o0685(.A(ori_ori_n477_), .B(ori_ori_n178_), .C(i), .Y(ori_ori_n714_));
  NA2        o0686(.A(ori_ori_n481_), .B(ori_ori_n84_), .Y(ori_ori_n715_));
  NA3        o0687(.A(ori_ori_n713_), .B(ori_ori_n533_), .C(ori_ori_n414_), .Y(ori_ori_n716_));
  NO4        o0688(.A(ori_ori_n716_), .B(ori_ori_n710_), .C(ori_ori_n703_), .D(ori_ori_n687_), .Y(ori_ori_n717_));
  NA4        o0689(.A(ori_ori_n717_), .B(ori_ori_n679_), .C(ori_ori_n635_), .D(ori_ori_n603_), .Y(ori08));
  NO2        o0690(.A(k), .B(h), .Y(ori_ori_n719_));
  AO210      o0691(.A0(ori_ori_n258_), .A1(ori_ori_n465_), .B0(ori_ori_n719_), .Y(ori_ori_n720_));
  NO2        o0692(.A(ori_ori_n720_), .B(ori_ori_n305_), .Y(ori_ori_n721_));
  NA2        o0693(.A(ori_ori_n643_), .B(ori_ori_n84_), .Y(ori_ori_n722_));
  NA2        o0694(.A(ori_ori_n722_), .B(ori_ori_n477_), .Y(ori_ori_n723_));
  AOI210     o0695(.A0(ori_ori_n723_), .A1(ori_ori_n721_), .B0(ori_ori_n510_), .Y(ori_ori_n724_));
  NA2        o0696(.A(ori_ori_n84_), .B(ori_ori_n112_), .Y(ori_ori_n725_));
  NO2        o0697(.A(ori_ori_n725_), .B(ori_ori_n57_), .Y(ori_ori_n726_));
  NO4        o0698(.A(ori_ori_n390_), .B(ori_ori_n114_), .C(j), .D(ori_ori_n219_), .Y(ori_ori_n727_));
  NA2        o0699(.A(ori_ori_n599_), .B(ori_ori_n238_), .Y(ori_ori_n728_));
  AOI220     o0700(.A0(ori_ori_n728_), .A1(ori_ori_n357_), .B0(ori_ori_n727_), .B1(ori_ori_n726_), .Y(ori_ori_n729_));
  AOI210     o0701(.A0(ori_ori_n599_), .A1(ori_ori_n160_), .B0(ori_ori_n84_), .Y(ori_ori_n730_));
  NA4        o0702(.A(ori_ori_n221_), .B(ori_ori_n143_), .C(ori_ori_n45_), .D(h), .Y(ori_ori_n731_));
  AN2        o0703(.A(l), .B(k), .Y(ori_ori_n732_));
  NA4        o0704(.A(ori_ori_n732_), .B(ori_ori_n110_), .C(ori_ori_n73_), .D(ori_ori_n219_), .Y(ori_ori_n733_));
  OAI210     o0705(.A0(ori_ori_n731_), .A1(g), .B0(ori_ori_n733_), .Y(ori_ori_n734_));
  NA2        o0706(.A(ori_ori_n734_), .B(ori_ori_n730_), .Y(ori_ori_n735_));
  NA4        o0707(.A(ori_ori_n735_), .B(ori_ori_n729_), .C(ori_ori_n724_), .D(ori_ori_n359_), .Y(ori_ori_n736_));
  NO4        o0708(.A(ori_ori_n178_), .B(ori_ori_n404_), .C(ori_ori_n114_), .D(g), .Y(ori_ori_n737_));
  NA2        o0709(.A(ori_ori_n737_), .B(ori_ori_n728_), .Y(ori_ori_n738_));
  NO2        o0710(.A(ori_ori_n38_), .B(ori_ori_n218_), .Y(ori_ori_n739_));
  AOI220     o0711(.A0(ori_ori_n645_), .A1(ori_ori_n356_), .B0(ori_ori_n739_), .B1(ori_ori_n586_), .Y(ori_ori_n740_));
  NA2        o0712(.A(ori_ori_n740_), .B(ori_ori_n738_), .Y(ori_ori_n741_));
  NO2        o0713(.A(ori_ori_n557_), .B(ori_ori_n35_), .Y(ori_ori_n742_));
  INV        o0714(.A(ori_ori_n742_), .Y(ori_ori_n743_));
  NO3        o0715(.A(ori_ori_n326_), .B(ori_ori_n133_), .C(ori_ori_n41_), .Y(ori_ori_n744_));
  NAi21      o0716(.An(ori_ori_n744_), .B(ori_ori_n733_), .Y(ori_ori_n745_));
  NA2        o0717(.A(ori_ori_n720_), .B(ori_ori_n138_), .Y(ori_ori_n746_));
  AOI220     o0718(.A0(ori_ori_n746_), .A1(ori_ori_n415_), .B0(ori_ori_n745_), .B1(ori_ori_n76_), .Y(ori_ori_n747_));
  OAI210     o0719(.A0(ori_ori_n743_), .A1(ori_ori_n87_), .B0(ori_ori_n747_), .Y(ori_ori_n748_));
  NA2        o0720(.A(ori_ori_n372_), .B(ori_ori_n43_), .Y(ori_ori_n749_));
  NA3        o0721(.A(ori_ori_n712_), .B(ori_ori_n343_), .C(ori_ori_n396_), .Y(ori_ori_n750_));
  NA3        o0722(.A(m), .B(l), .C(k), .Y(ori_ori_n751_));
  AOI210     o0723(.A0(ori_ori_n684_), .A1(ori_ori_n682_), .B0(ori_ori_n751_), .Y(ori_ori_n752_));
  NA3        o0724(.A(ori_ori_n115_), .B(k), .C(ori_ori_n87_), .Y(ori_ori_n753_));
  INV        o0725(.A(ori_ori_n752_), .Y(ori_ori_n754_));
  NA3        o0726(.A(ori_ori_n754_), .B(ori_ori_n750_), .C(ori_ori_n749_), .Y(ori_ori_n755_));
  NO4        o0727(.A(ori_ori_n755_), .B(ori_ori_n748_), .C(ori_ori_n741_), .D(ori_ori_n736_), .Y(ori_ori_n756_));
  NA2        o0728(.A(ori_ori_n645_), .B(ori_ori_n405_), .Y(ori_ori_n757_));
  NOi31      o0729(.An(g), .B(h), .C(f), .Y(ori_ori_n758_));
  NA2        o0730(.A(ori_ori_n659_), .B(ori_ori_n758_), .Y(ori_ori_n759_));
  AO210      o0731(.A0(ori_ori_n759_), .A1(ori_ori_n613_), .B0(ori_ori_n558_), .Y(ori_ori_n760_));
  NO3        o0732(.A(ori_ori_n409_), .B(ori_ori_n545_), .C(h), .Y(ori_ori_n761_));
  AOI210     o0733(.A0(ori_ori_n761_), .A1(ori_ori_n115_), .B0(ori_ori_n520_), .Y(ori_ori_n762_));
  NA4        o0734(.A(ori_ori_n762_), .B(ori_ori_n760_), .C(ori_ori_n757_), .D(ori_ori_n257_), .Y(ori_ori_n763_));
  NA2        o0735(.A(ori_ori_n732_), .B(ori_ori_n73_), .Y(ori_ori_n764_));
  NO4        o0736(.A(ori_ori_n711_), .B(ori_ori_n178_), .C(n), .D(i), .Y(ori_ori_n765_));
  NOi21      o0737(.An(h), .B(j), .Y(ori_ori_n766_));
  NA2        o0738(.A(ori_ori_n766_), .B(f), .Y(ori_ori_n767_));
  NO2        o0739(.A(ori_ori_n767_), .B(ori_ori_n251_), .Y(ori_ori_n768_));
  NO3        o0740(.A(ori_ori_n768_), .B(ori_ori_n765_), .C(ori_ori_n714_), .Y(ori_ori_n769_));
  OAI220     o0741(.A0(ori_ori_n769_), .A1(ori_ori_n764_), .B0(ori_ori_n615_), .B1(ori_ori_n62_), .Y(ori_ori_n770_));
  AOI210     o0742(.A0(ori_ori_n763_), .A1(l), .B0(ori_ori_n770_), .Y(ori_ori_n771_));
  NO2        o0743(.A(j), .B(i), .Y(ori_ori_n772_));
  NA2        o0744(.A(ori_ori_n772_), .B(ori_ori_n33_), .Y(ori_ori_n773_));
  NA2        o0745(.A(ori_ori_n434_), .B(ori_ori_n123_), .Y(ori_ori_n774_));
  OR2        o0746(.A(ori_ori_n774_), .B(ori_ori_n773_), .Y(ori_ori_n775_));
  NO3        o0747(.A(ori_ori_n155_), .B(ori_ori_n49_), .C(ori_ori_n112_), .Y(ori_ori_n776_));
  NO3        o0748(.A(ori_ori_n562_), .B(ori_ori_n153_), .C(ori_ori_n73_), .Y(ori_ori_n777_));
  NO3        o0749(.A(ori_ori_n504_), .B(ori_ori_n452_), .C(j), .Y(ori_ori_n778_));
  OAI210     o0750(.A0(ori_ori_n777_), .A1(ori_ori_n776_), .B0(ori_ori_n778_), .Y(ori_ori_n779_));
  OAI210     o0751(.A0(ori_ori_n759_), .A1(ori_ori_n62_), .B0(ori_ori_n779_), .Y(ori_ori_n780_));
  INV        o0752(.A(j), .Y(ori_ori_n781_));
  NO3        o0753(.A(ori_ori_n305_), .B(ori_ori_n781_), .C(ori_ori_n40_), .Y(ori_ori_n782_));
  AOI210     o0754(.A0(ori_ori_n550_), .A1(n), .B0(ori_ori_n572_), .Y(ori_ori_n783_));
  NA2        o0755(.A(ori_ori_n783_), .B(ori_ori_n575_), .Y(ori_ori_n784_));
  AN3        o0756(.A(ori_ori_n784_), .B(ori_ori_n782_), .C(ori_ori_n99_), .Y(ori_ori_n785_));
  NO3        o0757(.A(ori_ori_n178_), .B(ori_ori_n404_), .C(ori_ori_n114_), .Y(ori_ori_n786_));
  AOI220     o0758(.A0(ori_ori_n786_), .A1(ori_ori_n252_), .B0(ori_ori_n638_), .B1(ori_ori_n316_), .Y(ori_ori_n787_));
  NAi31      o0759(.An(ori_ori_n631_), .B(ori_ori_n93_), .C(ori_ori_n84_), .Y(ori_ori_n788_));
  NA2        o0760(.A(ori_ori_n788_), .B(ori_ori_n787_), .Y(ori_ori_n789_));
  NO2        o0761(.A(ori_ori_n305_), .B(ori_ori_n138_), .Y(ori_ori_n790_));
  AOI220     o0762(.A0(ori_ori_n790_), .A1(ori_ori_n645_), .B0(ori_ori_n744_), .B1(ori_ori_n730_), .Y(ori_ori_n791_));
  NO2        o0763(.A(ori_ori_n751_), .B(ori_ori_n91_), .Y(ori_ori_n792_));
  NA2        o0764(.A(ori_ori_n792_), .B(ori_ori_n610_), .Y(ori_ori_n793_));
  NO2        o0765(.A(ori_ori_n612_), .B(ori_ori_n119_), .Y(ori_ori_n794_));
  OAI210     o0766(.A0(ori_ori_n794_), .A1(ori_ori_n778_), .B0(ori_ori_n700_), .Y(ori_ori_n795_));
  NA3        o0767(.A(ori_ori_n795_), .B(ori_ori_n793_), .C(ori_ori_n791_), .Y(ori_ori_n796_));
  OR4        o0768(.A(ori_ori_n796_), .B(ori_ori_n789_), .C(ori_ori_n785_), .D(ori_ori_n780_), .Y(ori_ori_n797_));
  NA3        o0769(.A(ori_ori_n783_), .B(ori_ori_n575_), .C(ori_ori_n574_), .Y(ori_ori_n798_));
  NA4        o0770(.A(ori_ori_n798_), .B(ori_ori_n221_), .C(ori_ori_n465_), .D(ori_ori_n34_), .Y(ori_ori_n799_));
  NO4        o0771(.A(ori_ori_n504_), .B(ori_ori_n448_), .C(j), .D(f), .Y(ori_ori_n800_));
  OAI220     o0772(.A0(ori_ori_n731_), .A1(ori_ori_n722_), .B0(ori_ori_n341_), .B1(ori_ori_n38_), .Y(ori_ori_n801_));
  AOI210     o0773(.A0(ori_ori_n800_), .A1(ori_ori_n264_), .B0(ori_ori_n801_), .Y(ori_ori_n802_));
  NA3        o0774(.A(ori_ori_n565_), .B(ori_ori_n298_), .C(h), .Y(ori_ori_n803_));
  NO2        o0775(.A(ori_ori_n92_), .B(ori_ori_n47_), .Y(ori_ori_n804_));
  NO2        o0776(.A(ori_ori_n803_), .B(ori_ori_n627_), .Y(ori_ori_n805_));
  AOI210     o0777(.A0(ori_ori_n804_), .A1(ori_ori_n664_), .B0(ori_ori_n805_), .Y(ori_ori_n806_));
  NA3        o0778(.A(ori_ori_n806_), .B(ori_ori_n802_), .C(ori_ori_n799_), .Y(ori_ori_n807_));
  NA2        o0779(.A(ori_ori_n792_), .B(ori_ori_n243_), .Y(ori_ori_n808_));
  NO2        o0780(.A(ori_ori_n683_), .B(ori_ori_n73_), .Y(ori_ori_n809_));
  AOI210     o0781(.A0(ori_ori_n800_), .A1(ori_ori_n809_), .B0(ori_ori_n345_), .Y(ori_ori_n810_));
  OAI210     o0782(.A0(ori_ori_n751_), .A1(ori_ori_n681_), .B0(ori_ori_n539_), .Y(ori_ori_n811_));
  NA3        o0783(.A(ori_ori_n255_), .B(ori_ori_n59_), .C(b), .Y(ori_ori_n812_));
  AOI220     o0784(.A0(ori_ori_n626_), .A1(ori_ori_n29_), .B0(ori_ori_n481_), .B1(ori_ori_n84_), .Y(ori_ori_n813_));
  NA2        o0785(.A(ori_ori_n813_), .B(ori_ori_n812_), .Y(ori_ori_n814_));
  NA2        o0786(.A(ori_ori_n814_), .B(ori_ori_n811_), .Y(ori_ori_n815_));
  NA3        o0787(.A(ori_ori_n815_), .B(ori_ori_n810_), .C(ori_ori_n808_), .Y(ori_ori_n816_));
  NOi41      o0788(.An(ori_ori_n775_), .B(ori_ori_n816_), .C(ori_ori_n807_), .D(ori_ori_n797_), .Y(ori_ori_n817_));
  NO3        o0789(.A(ori_ori_n351_), .B(ori_ori_n307_), .C(ori_ori_n114_), .Y(ori_ori_n818_));
  NA2        o0790(.A(ori_ori_n818_), .B(ori_ori_n784_), .Y(ori_ori_n819_));
  NO3        o0791(.A(ori_ori_n545_), .B(ori_ori_n94_), .C(h), .Y(ori_ori_n820_));
  NA2        o0792(.A(ori_ori_n820_), .B(ori_ori_n726_), .Y(ori_ori_n821_));
  NA3        o0793(.A(ori_ori_n821_), .B(ori_ori_n819_), .C(ori_ori_n417_), .Y(ori_ori_n822_));
  OR2        o0794(.A(ori_ori_n681_), .B(ori_ori_n92_), .Y(ori_ori_n823_));
  NOi31      o0795(.An(b), .B(d), .C(a), .Y(ori_ori_n824_));
  NO2        o0796(.A(ori_ori_n824_), .B(ori_ori_n624_), .Y(ori_ori_n825_));
  NO2        o0797(.A(ori_ori_n825_), .B(n), .Y(ori_ori_n826_));
  NOi21      o0798(.An(ori_ori_n813_), .B(ori_ori_n826_), .Y(ori_ori_n827_));
  OAI220     o0799(.A0(ori_ori_n827_), .A1(ori_ori_n823_), .B0(ori_ori_n803_), .B1(ori_ori_n625_), .Y(ori_ori_n828_));
  NO2        o0800(.A(ori_ori_n573_), .B(ori_ori_n84_), .Y(ori_ori_n829_));
  NO3        o0801(.A(ori_ori_n644_), .B(ori_ori_n336_), .C(ori_ori_n119_), .Y(ori_ori_n830_));
  NOi21      o0802(.An(ori_ori_n830_), .B(ori_ori_n165_), .Y(ori_ori_n831_));
  AOI210     o0803(.A0(ori_ori_n818_), .A1(ori_ori_n829_), .B0(ori_ori_n831_), .Y(ori_ori_n832_));
  OAI210     o0804(.A0(ori_ori_n731_), .A1(ori_ori_n406_), .B0(ori_ori_n832_), .Y(ori_ori_n833_));
  NO2        o0805(.A(ori_ori_n711_), .B(n), .Y(ori_ori_n834_));
  AOI220     o0806(.A0(ori_ori_n790_), .A1(ori_ori_n688_), .B0(ori_ori_n834_), .B1(ori_ori_n721_), .Y(ori_ori_n835_));
  NO2        o0807(.A(ori_ori_n331_), .B(ori_ori_n242_), .Y(ori_ori_n836_));
  OAI210     o0808(.A0(ori_ori_n96_), .A1(ori_ori_n93_), .B0(ori_ori_n836_), .Y(ori_ori_n837_));
  NA2        o0809(.A(ori_ori_n123_), .B(ori_ori_n84_), .Y(ori_ori_n838_));
  AOI210     o0810(.A0(ori_ori_n438_), .A1(ori_ori_n430_), .B0(ori_ori_n838_), .Y(ori_ori_n839_));
  NAi21      o0811(.An(ori_ori_n839_), .B(ori_ori_n837_), .Y(ori_ori_n840_));
  OAI210     o0812(.A0(ori_ori_n618_), .A1(ori_ori_n617_), .B0(ori_ori_n373_), .Y(ori_ori_n841_));
  NAi31      o0813(.An(ori_ori_n840_), .B(ori_ori_n841_), .C(ori_ori_n835_), .Y(ori_ori_n842_));
  NO4        o0814(.A(ori_ori_n842_), .B(ori_ori_n833_), .C(ori_ori_n828_), .D(ori_ori_n822_), .Y(ori_ori_n843_));
  NA4        o0815(.A(ori_ori_n843_), .B(ori_ori_n817_), .C(ori_ori_n771_), .D(ori_ori_n756_), .Y(ori09));
  INV        o0816(.A(ori_ori_n124_), .Y(ori_ori_n845_));
  NA2        o0817(.A(f), .B(e), .Y(ori_ori_n846_));
  NO2        o0818(.A(ori_ori_n231_), .B(ori_ori_n114_), .Y(ori_ori_n847_));
  NA2        o0819(.A(ori_ori_n847_), .B(g), .Y(ori_ori_n848_));
  NA4        o0820(.A(ori_ori_n319_), .B(ori_ori_n490_), .C(ori_ori_n267_), .D(ori_ori_n121_), .Y(ori_ori_n849_));
  AOI210     o0821(.A0(ori_ori_n849_), .A1(g), .B0(ori_ori_n487_), .Y(ori_ori_n850_));
  AOI210     o0822(.A0(ori_ori_n850_), .A1(ori_ori_n848_), .B0(ori_ori_n846_), .Y(ori_ori_n851_));
  NA2        o0823(.A(ori_ori_n458_), .B(e), .Y(ori_ori_n852_));
  NO2        o0824(.A(ori_ori_n852_), .B(ori_ori_n530_), .Y(ori_ori_n853_));
  AOI210     o0825(.A0(ori_ori_n851_), .A1(ori_ori_n845_), .B0(ori_ori_n853_), .Y(ori_ori_n854_));
  NO2        o0826(.A(ori_ori_n209_), .B(ori_ori_n218_), .Y(ori_ori_n855_));
  NA3        o0827(.A(m), .B(l), .C(i), .Y(ori_ori_n856_));
  OAI220     o0828(.A0(ori_ori_n612_), .A1(ori_ori_n856_), .B0(ori_ori_n363_), .B1(ori_ori_n546_), .Y(ori_ori_n857_));
  NA4        o0829(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(g), .D(f), .Y(ori_ori_n858_));
  NAi31      o0830(.An(ori_ori_n857_), .B(ori_ori_n858_), .C(ori_ori_n453_), .Y(ori_ori_n859_));
  OR2        o0831(.A(ori_ori_n859_), .B(ori_ori_n855_), .Y(ori_ori_n860_));
  NA3        o0832(.A(ori_ori_n823_), .B(ori_ori_n588_), .C(ori_ori_n539_), .Y(ori_ori_n861_));
  OA210      o0833(.A0(ori_ori_n861_), .A1(ori_ori_n860_), .B0(ori_ori_n826_), .Y(ori_ori_n862_));
  INV        o0834(.A(ori_ori_n348_), .Y(ori_ori_n863_));
  NO2        o0835(.A(ori_ori_n129_), .B(ori_ori_n127_), .Y(ori_ori_n864_));
  NOi31      o0836(.An(k), .B(m), .C(l), .Y(ori_ori_n865_));
  NO2        o0837(.A(ori_ori_n350_), .B(ori_ori_n865_), .Y(ori_ori_n866_));
  AOI210     o0838(.A0(ori_ori_n866_), .A1(ori_ori_n864_), .B0(ori_ori_n621_), .Y(ori_ori_n867_));
  NA2        o0839(.A(ori_ori_n812_), .B(ori_ori_n341_), .Y(ori_ori_n868_));
  NA2        o0840(.A(ori_ori_n352_), .B(ori_ori_n354_), .Y(ori_ori_n869_));
  OAI210     o0841(.A0(ori_ori_n209_), .A1(ori_ori_n218_), .B0(ori_ori_n869_), .Y(ori_ori_n870_));
  AOI220     o0842(.A0(ori_ori_n870_), .A1(ori_ori_n868_), .B0(ori_ori_n867_), .B1(ori_ori_n863_), .Y(ori_ori_n871_));
  NA2        o0843(.A(ori_ori_n173_), .B(ori_ori_n116_), .Y(ori_ori_n872_));
  NA3        o0844(.A(ori_ori_n872_), .B(ori_ori_n720_), .C(ori_ori_n138_), .Y(ori_ori_n873_));
  NA3        o0845(.A(ori_ori_n873_), .B(ori_ori_n194_), .C(ori_ori_n31_), .Y(ori_ori_n874_));
  NA4        o0846(.A(ori_ori_n874_), .B(ori_ori_n871_), .C(ori_ori_n646_), .D(ori_ori_n82_), .Y(ori_ori_n875_));
  NO2        o0847(.A(ori_ori_n608_), .B(ori_ori_n516_), .Y(ori_ori_n876_));
  NOi21      o0848(.An(f), .B(d), .Y(ori_ori_n877_));
  NA2        o0849(.A(ori_ori_n877_), .B(m), .Y(ori_ori_n878_));
  NO2        o0850(.A(ori_ori_n878_), .B(ori_ori_n52_), .Y(ori_ori_n879_));
  NOi32      o0851(.An(g), .Bn(f), .C(d), .Y(ori_ori_n880_));
  NA4        o0852(.A(ori_ori_n880_), .B(ori_ori_n626_), .C(ori_ori_n29_), .D(m), .Y(ori_ori_n881_));
  NOi21      o0853(.An(ori_ori_n320_), .B(ori_ori_n881_), .Y(ori_ori_n882_));
  AOI210     o0854(.A0(ori_ori_n879_), .A1(ori_ori_n563_), .B0(ori_ori_n882_), .Y(ori_ori_n883_));
  NA3        o0855(.A(ori_ori_n319_), .B(ori_ori_n267_), .C(ori_ori_n121_), .Y(ori_ori_n884_));
  AN2        o0856(.A(f), .B(d), .Y(ori_ori_n885_));
  NA3        o0857(.A(ori_ori_n495_), .B(ori_ori_n885_), .C(ori_ori_n84_), .Y(ori_ori_n886_));
  NO3        o0858(.A(ori_ori_n886_), .B(ori_ori_n73_), .C(ori_ori_n219_), .Y(ori_ori_n887_));
  NA2        o0859(.A(ori_ori_n884_), .B(ori_ori_n887_), .Y(ori_ori_n888_));
  NAi31      o0860(.An(ori_ori_n509_), .B(ori_ori_n888_), .C(ori_ori_n883_), .Y(ori_ori_n889_));
  NO4        o0861(.A(ori_ori_n644_), .B(ori_ori_n134_), .C(ori_ori_n336_), .D(ori_ori_n156_), .Y(ori_ori_n890_));
  NO2        o0862(.A(ori_ori_n675_), .B(ori_ori_n336_), .Y(ori_ori_n891_));
  INV        o0863(.A(ori_ori_n890_), .Y(ori_ori_n892_));
  NA2        o0864(.A(ori_ori_n624_), .B(ori_ori_n84_), .Y(ori_ori_n893_));
  NO2        o0865(.A(ori_ori_n869_), .B(ori_ori_n893_), .Y(ori_ori_n894_));
  NA3        o0866(.A(ori_ori_n164_), .B(ori_ori_n110_), .C(ori_ori_n109_), .Y(ori_ori_n895_));
  OAI220     o0867(.A0(ori_ori_n886_), .A1(ori_ori_n443_), .B0(ori_ori_n348_), .B1(ori_ori_n895_), .Y(ori_ori_n896_));
  NOi41      o0868(.An(ori_ori_n229_), .B(ori_ori_n896_), .C(ori_ori_n894_), .D(ori_ori_n314_), .Y(ori_ori_n897_));
  NA2        o0869(.A(c), .B(ori_ori_n118_), .Y(ori_ori_n898_));
  NO2        o0870(.A(ori_ori_n898_), .B(ori_ori_n421_), .Y(ori_ori_n899_));
  NA3        o0871(.A(ori_ori_n899_), .B(ori_ori_n528_), .C(f), .Y(ori_ori_n900_));
  OR2        o0872(.A(ori_ori_n681_), .B(ori_ori_n559_), .Y(ori_ori_n901_));
  INV        o0873(.A(ori_ori_n901_), .Y(ori_ori_n902_));
  NA2        o0874(.A(ori_ori_n825_), .B(ori_ori_n113_), .Y(ori_ori_n903_));
  NA2        o0875(.A(ori_ori_n903_), .B(ori_ori_n902_), .Y(ori_ori_n904_));
  NA4        o0876(.A(ori_ori_n904_), .B(ori_ori_n900_), .C(ori_ori_n897_), .D(ori_ori_n892_), .Y(ori_ori_n905_));
  NO4        o0877(.A(ori_ori_n905_), .B(ori_ori_n889_), .C(ori_ori_n875_), .D(ori_ori_n862_), .Y(ori_ori_n906_));
  NA2        o0878(.A(ori_ori_n114_), .B(j), .Y(ori_ori_n907_));
  NO2        o0879(.A(ori_ori_n341_), .B(ori_ori_n858_), .Y(ori_ori_n908_));
  NO2        o0880(.A(ori_ori_n138_), .B(ori_ori_n134_), .Y(ori_ori_n909_));
  NO2        o0881(.A(ori_ori_n236_), .B(ori_ori_n230_), .Y(ori_ori_n910_));
  AOI220     o0882(.A0(ori_ori_n910_), .A1(ori_ori_n233_), .B0(ori_ori_n312_), .B1(ori_ori_n909_), .Y(ori_ori_n911_));
  NO2        o0883(.A(ori_ori_n443_), .B(ori_ori_n846_), .Y(ori_ori_n912_));
  NA2        o0884(.A(ori_ori_n912_), .B(ori_ori_n580_), .Y(ori_ori_n913_));
  NA2        o0885(.A(ori_ori_n913_), .B(ori_ori_n911_), .Y(ori_ori_n914_));
  NA2        o0886(.A(e), .B(d), .Y(ori_ori_n915_));
  OAI220     o0887(.A0(ori_ori_n915_), .A1(c), .B0(ori_ori_n331_), .B1(d), .Y(ori_ori_n916_));
  NA3        o0888(.A(ori_ori_n916_), .B(ori_ori_n470_), .C(ori_ori_n526_), .Y(ori_ori_n917_));
  AOI210     o0889(.A0(ori_ori_n534_), .A1(ori_ori_n185_), .B0(ori_ori_n236_), .Y(ori_ori_n918_));
  AOI210     o0890(.A0(ori_ori_n645_), .A1(ori_ori_n356_), .B0(ori_ori_n918_), .Y(ori_ori_n919_));
  NA2        o0891(.A(ori_ori_n291_), .B(ori_ori_n169_), .Y(ori_ori_n920_));
  NA2        o0892(.A(ori_ori_n887_), .B(ori_ori_n920_), .Y(ori_ori_n921_));
  NA3        o0893(.A(ori_ori_n172_), .B(ori_ori_n85_), .C(ori_ori_n34_), .Y(ori_ori_n922_));
  NA4        o0894(.A(ori_ori_n922_), .B(ori_ori_n921_), .C(ori_ori_n919_), .D(ori_ori_n917_), .Y(ori_ori_n923_));
  NO3        o0895(.A(ori_ori_n923_), .B(ori_ori_n914_), .C(ori_ori_n908_), .Y(ori_ori_n924_));
  OR2        o0896(.A(ori_ori_n722_), .B(ori_ori_n222_), .Y(ori_ori_n925_));
  OAI220     o0897(.A0(ori_ori_n644_), .A1(ori_ori_n61_), .B0(ori_ori_n307_), .B1(j), .Y(ori_ori_n926_));
  AOI220     o0898(.A0(ori_ori_n926_), .A1(ori_ori_n891_), .B0(ori_ori_n636_), .B1(ori_ori_n643_), .Y(ori_ori_n927_));
  OAI210     o0899(.A0(ori_ori_n852_), .A1(ori_ori_n175_), .B0(ori_ori_n927_), .Y(ori_ori_n928_));
  OAI210     o0900(.A0(ori_ori_n847_), .A1(ori_ori_n920_), .B0(ori_ori_n880_), .Y(ori_ori_n929_));
  NO2        o0901(.A(ori_ori_n929_), .B(ori_ori_n627_), .Y(ori_ori_n930_));
  AOI210     o0902(.A0(ori_ori_n120_), .A1(ori_ori_n119_), .B0(ori_ori_n266_), .Y(ori_ori_n931_));
  NO2        o0903(.A(ori_ori_n931_), .B(ori_ori_n881_), .Y(ori_ori_n932_));
  AO210      o0904(.A0(ori_ori_n868_), .A1(ori_ori_n857_), .B0(ori_ori_n932_), .Y(ori_ori_n933_));
  NO3        o0905(.A(ori_ori_n933_), .B(ori_ori_n930_), .C(ori_ori_n928_), .Y(ori_ori_n934_));
  AO220      o0906(.A0(ori_ori_n470_), .A1(ori_ori_n766_), .B0(ori_ori_n180_), .B1(f), .Y(ori_ori_n935_));
  OAI210     o0907(.A0(ori_ori_n935_), .A1(ori_ori_n473_), .B0(ori_ori_n916_), .Y(ori_ori_n936_));
  NO2        o0908(.A(ori_ori_n452_), .B(ori_ori_n70_), .Y(ori_ori_n937_));
  OAI210     o0909(.A0(ori_ori_n861_), .A1(ori_ori_n937_), .B0(ori_ori_n726_), .Y(ori_ori_n938_));
  AN4        o0910(.A(ori_ori_n938_), .B(ori_ori_n936_), .C(ori_ori_n934_), .D(ori_ori_n925_), .Y(ori_ori_n939_));
  NA4        o0911(.A(ori_ori_n939_), .B(ori_ori_n924_), .C(ori_ori_n906_), .D(ori_ori_n854_), .Y(ori12));
  NO2        o0912(.A(ori_ori_n468_), .B(c), .Y(ori_ori_n941_));
  NO4        o0913(.A(ori_ori_n457_), .B(ori_ori_n258_), .C(ori_ori_n604_), .D(ori_ori_n219_), .Y(ori_ori_n942_));
  NA2        o0914(.A(ori_ori_n942_), .B(ori_ori_n941_), .Y(ori_ori_n943_));
  NA2        o0915(.A(ori_ori_n563_), .B(ori_ori_n937_), .Y(ori_ori_n944_));
  NO2        o0916(.A(ori_ori_n468_), .B(ori_ori_n118_), .Y(ori_ori_n945_));
  NO2        o0917(.A(ori_ori_n864_), .B(ori_ori_n363_), .Y(ori_ori_n946_));
  NO2        o0918(.A(ori_ori_n681_), .B(ori_ori_n390_), .Y(ori_ori_n947_));
  AOI220     o0919(.A0(ori_ori_n947_), .A1(ori_ori_n561_), .B0(ori_ori_n946_), .B1(ori_ori_n945_), .Y(ori_ori_n948_));
  NA4        o0920(.A(ori_ori_n948_), .B(ori_ori_n944_), .C(ori_ori_n943_), .D(ori_ori_n456_), .Y(ori_ori_n949_));
  AOI210     o0921(.A0(ori_ori_n239_), .A1(ori_ori_n347_), .B0(ori_ori_n206_), .Y(ori_ori_n950_));
  OR2        o0922(.A(ori_ori_n950_), .B(ori_ori_n942_), .Y(ori_ori_n951_));
  AOI210     o0923(.A0(ori_ori_n344_), .A1(ori_ori_n402_), .B0(ori_ori_n219_), .Y(ori_ori_n952_));
  OAI210     o0924(.A0(ori_ori_n952_), .A1(ori_ori_n951_), .B0(ori_ori_n416_), .Y(ori_ori_n953_));
  NO2        o0925(.A(ori_ori_n661_), .B(ori_ori_n269_), .Y(ori_ori_n954_));
  NO2        o0926(.A(ori_ori_n612_), .B(ori_ori_n856_), .Y(ori_ori_n955_));
  AOI220     o0927(.A0(ori_ori_n955_), .A1(ori_ori_n586_), .B0(ori_ori_n836_), .B1(ori_ori_n954_), .Y(ori_ori_n956_));
  NO2        o0928(.A(ori_ori_n155_), .B(ori_ori_n242_), .Y(ori_ori_n957_));
  NA3        o0929(.A(ori_ori_n957_), .B(ori_ori_n245_), .C(i), .Y(ori_ori_n958_));
  NA3        o0930(.A(ori_ori_n958_), .B(ori_ori_n956_), .C(ori_ori_n953_), .Y(ori_ori_n959_));
  OR2        o0931(.A(ori_ori_n332_), .B(ori_ori_n945_), .Y(ori_ori_n960_));
  NA2        o0932(.A(ori_ori_n960_), .B(ori_ori_n364_), .Y(ori_ori_n961_));
  NO3        o0933(.A(ori_ori_n134_), .B(ori_ori_n156_), .C(ori_ori_n219_), .Y(ori_ori_n962_));
  NA2        o0934(.A(ori_ori_n962_), .B(ori_ori_n550_), .Y(ori_ori_n963_));
  NA4        o0935(.A(ori_ori_n458_), .B(ori_ori_n450_), .C(ori_ori_n186_), .D(g), .Y(ori_ori_n964_));
  NA3        o0936(.A(ori_ori_n964_), .B(ori_ori_n963_), .C(ori_ori_n961_), .Y(ori_ori_n965_));
  NO3        o0937(.A(ori_ori_n686_), .B(ori_ori_n92_), .C(ori_ori_n45_), .Y(ori_ori_n966_));
  NO4        o0938(.A(ori_ori_n966_), .B(ori_ori_n965_), .C(ori_ori_n959_), .D(ori_ori_n949_), .Y(ori_ori_n967_));
  NO2        o0939(.A(ori_ori_n380_), .B(ori_ori_n379_), .Y(ori_ori_n968_));
  INV        o0940(.A(ori_ori_n72_), .Y(ori_ori_n969_));
  NA2        o0941(.A(ori_ori_n573_), .B(ori_ori_n148_), .Y(ori_ori_n970_));
  NOi21      o0942(.An(ori_ori_n34_), .B(ori_ori_n675_), .Y(ori_ori_n971_));
  AOI220     o0943(.A0(ori_ori_n971_), .A1(ori_ori_n970_), .B0(ori_ori_n969_), .B1(ori_ori_n968_), .Y(ori_ori_n972_));
  OAI210     o0944(.A0(ori_ori_n256_), .A1(ori_ori_n45_), .B0(ori_ori_n972_), .Y(ori_ori_n973_));
  INV        o0945(.A(ori_ori_n330_), .Y(ori_ori_n974_));
  NO2        o0946(.A(ori_ori_n49_), .B(ori_ori_n45_), .Y(ori_ori_n975_));
  NO2        o0947(.A(ori_ori_n523_), .B(ori_ori_n307_), .Y(ori_ori_n976_));
  INV        o0948(.A(ori_ori_n976_), .Y(ori_ori_n977_));
  NO2        o0949(.A(ori_ori_n977_), .B(ori_ori_n148_), .Y(ori_ori_n978_));
  INV        o0950(.A(ori_ori_n377_), .Y(ori_ori_n979_));
  NO4        o0951(.A(ori_ori_n979_), .B(ori_ori_n978_), .C(ori_ori_n974_), .D(ori_ori_n973_), .Y(ori_ori_n980_));
  NA2        o0952(.A(ori_ori_n356_), .B(g), .Y(ori_ori_n981_));
  NA2        o0953(.A(ori_ori_n167_), .B(i), .Y(ori_ori_n982_));
  NA2        o0954(.A(ori_ori_n46_), .B(i), .Y(ori_ori_n983_));
  OAI220     o0955(.A0(ori_ori_n983_), .A1(ori_ori_n205_), .B0(ori_ori_n982_), .B1(ori_ori_n92_), .Y(ori_ori_n984_));
  AOI210     o0956(.A0(ori_ori_n432_), .A1(ori_ori_n37_), .B0(ori_ori_n984_), .Y(ori_ori_n985_));
  NO2        o0957(.A(ori_ori_n148_), .B(ori_ori_n84_), .Y(ori_ori_n986_));
  OR2        o0958(.A(ori_ori_n986_), .B(ori_ori_n572_), .Y(ori_ori_n987_));
  NA2        o0959(.A(ori_ori_n573_), .B(ori_ori_n394_), .Y(ori_ori_n988_));
  AOI210     o0960(.A0(ori_ori_n988_), .A1(n), .B0(ori_ori_n987_), .Y(ori_ori_n989_));
  OAI220     o0961(.A0(ori_ori_n989_), .A1(ori_ori_n981_), .B0(ori_ori_n985_), .B1(ori_ori_n341_), .Y(ori_ori_n990_));
  NO2        o0962(.A(ori_ori_n681_), .B(ori_ori_n516_), .Y(ori_ori_n991_));
  NA3        o0963(.A(ori_ori_n352_), .B(ori_ori_n650_), .C(i), .Y(ori_ori_n992_));
  OAI210     o0964(.A0(ori_ori_n452_), .A1(ori_ori_n319_), .B0(ori_ori_n992_), .Y(ori_ori_n993_));
  OAI220     o0965(.A0(ori_ori_n993_), .A1(ori_ori_n991_), .B0(ori_ori_n700_), .B1(ori_ori_n777_), .Y(ori_ori_n994_));
  NA3        o0966(.A(ori_ori_n333_), .B(ori_ori_n120_), .C(g), .Y(ori_ori_n995_));
  AOI210     o0967(.A0(ori_ori_n697_), .A1(ori_ori_n995_), .B0(m), .Y(ori_ori_n996_));
  OAI210     o0968(.A0(ori_ori_n996_), .A1(ori_ori_n946_), .B0(ori_ori_n332_), .Y(ori_ori_n997_));
  NA2        o0969(.A(ori_ori_n715_), .B(ori_ori_n893_), .Y(ori_ori_n998_));
  NA2        o0970(.A(ori_ori_n858_), .B(ori_ori_n453_), .Y(ori_ori_n999_));
  NA2        o0971(.A(ori_ori_n999_), .B(ori_ori_n998_), .Y(ori_ori_n1000_));
  NA3        o0972(.A(ori_ori_n1000_), .B(ori_ori_n997_), .C(ori_ori_n994_), .Y(ori_ori_n1001_));
  NO2        o0973(.A(ori_ori_n390_), .B(ori_ori_n91_), .Y(ori_ori_n1002_));
  OAI210     o0974(.A0(ori_ori_n1002_), .A1(ori_ori_n954_), .B0(ori_ori_n243_), .Y(ori_ori_n1003_));
  NA2        o0975(.A(ori_ori_n685_), .B(ori_ori_n88_), .Y(ori_ori_n1004_));
  NO2        o0976(.A(ori_ori_n476_), .B(ori_ori_n219_), .Y(ori_ori_n1005_));
  AOI220     o0977(.A0(ori_ori_n1005_), .A1(ori_ori_n395_), .B0(ori_ori_n960_), .B1(ori_ori_n223_), .Y(ori_ori_n1006_));
  AOI220     o0978(.A0(ori_ori_n947_), .A1(ori_ori_n957_), .B0(ori_ori_n610_), .B1(ori_ori_n90_), .Y(ori_ori_n1007_));
  NA4        o0979(.A(ori_ori_n1007_), .B(ori_ori_n1006_), .C(ori_ori_n1004_), .D(ori_ori_n1003_), .Y(ori_ori_n1008_));
  OAI210     o0980(.A0(ori_ori_n999_), .A1(ori_ori_n955_), .B0(ori_ori_n561_), .Y(ori_ori_n1009_));
  AOI210     o0981(.A0(ori_ori_n433_), .A1(ori_ori_n425_), .B0(ori_ori_n838_), .Y(ori_ori_n1010_));
  OAI210     o0982(.A0(ori_ori_n380_), .A1(ori_ori_n379_), .B0(ori_ori_n111_), .Y(ori_ori_n1011_));
  AOI210     o0983(.A0(ori_ori_n1011_), .A1(ori_ori_n554_), .B0(ori_ori_n1010_), .Y(ori_ori_n1012_));
  NA2        o0984(.A(ori_ori_n996_), .B(ori_ori_n945_), .Y(ori_ori_n1013_));
  NO3        o0985(.A(ori_ori_n907_), .B(ori_ori_n49_), .C(ori_ori_n45_), .Y(ori_ori_n1014_));
  AOI220     o0986(.A0(ori_ori_n1014_), .A1(ori_ori_n648_), .B0(ori_ori_n666_), .B1(ori_ori_n550_), .Y(ori_ori_n1015_));
  NA4        o0987(.A(ori_ori_n1015_), .B(ori_ori_n1013_), .C(ori_ori_n1012_), .D(ori_ori_n1009_), .Y(ori_ori_n1016_));
  NO4        o0988(.A(ori_ori_n1016_), .B(ori_ori_n1008_), .C(ori_ori_n1001_), .D(ori_ori_n990_), .Y(ori_ori_n1017_));
  NAi31      o0989(.An(ori_ori_n144_), .B(ori_ori_n434_), .C(n), .Y(ori_ori_n1018_));
  NO3        o0990(.A(ori_ori_n127_), .B(ori_ori_n350_), .C(ori_ori_n865_), .Y(ori_ori_n1019_));
  NO2        o0991(.A(ori_ori_n1019_), .B(ori_ori_n1018_), .Y(ori_ori_n1020_));
  NO3        o0992(.A(ori_ori_n279_), .B(ori_ori_n144_), .C(ori_ori_n421_), .Y(ori_ori_n1021_));
  AOI210     o0993(.A0(ori_ori_n1021_), .A1(ori_ori_n517_), .B0(ori_ori_n1020_), .Y(ori_ori_n1022_));
  NA2        o0994(.A(ori_ori_n510_), .B(i), .Y(ori_ori_n1023_));
  NA2        o0995(.A(ori_ori_n1023_), .B(ori_ori_n1022_), .Y(ori_ori_n1024_));
  NA2        o0996(.A(ori_ori_n236_), .B(ori_ori_n176_), .Y(ori_ori_n1025_));
  NO3        o0997(.A(ori_ori_n316_), .B(ori_ori_n458_), .C(ori_ori_n180_), .Y(ori_ori_n1026_));
  NOi31      o0998(.An(ori_ori_n1025_), .B(ori_ori_n1026_), .C(ori_ori_n219_), .Y(ori_ori_n1027_));
  NAi21      o0999(.An(ori_ori_n573_), .B(ori_ori_n1005_), .Y(ori_ori_n1028_));
  NA2        o1000(.A(ori_ori_n501_), .B(g), .Y(ori_ori_n1029_));
  NA2        o1001(.A(ori_ori_n1029_), .B(ori_ori_n1028_), .Y(ori_ori_n1030_));
  OAI220     o1002(.A0(ori_ori_n1018_), .A1(ori_ori_n239_), .B0(ori_ori_n992_), .B1(ori_ori_n625_), .Y(ori_ori_n1031_));
  NO2        o1003(.A(ori_ori_n682_), .B(ori_ori_n390_), .Y(ori_ori_n1032_));
  NA2        o1004(.A(ori_ori_n950_), .B(ori_ori_n941_), .Y(ori_ori_n1033_));
  OAI220     o1005(.A0(ori_ori_n947_), .A1(ori_ori_n955_), .B0(ori_ori_n563_), .B1(ori_ori_n442_), .Y(ori_ori_n1034_));
  NA3        o1006(.A(ori_ori_n1034_), .B(ori_ori_n1033_), .C(ori_ori_n642_), .Y(ori_ori_n1035_));
  OAI210     o1007(.A0(ori_ori_n950_), .A1(ori_ori_n942_), .B0(ori_ori_n1025_), .Y(ori_ori_n1036_));
  NA3        o1008(.A(ori_ori_n988_), .B(ori_ori_n506_), .C(ori_ori_n46_), .Y(ori_ori_n1037_));
  AOI210     o1009(.A0(ori_ori_n393_), .A1(ori_ori_n391_), .B0(ori_ori_n340_), .Y(ori_ori_n1038_));
  NA4        o1010(.A(ori_ori_n1038_), .B(ori_ori_n1037_), .C(ori_ori_n1036_), .D(ori_ori_n280_), .Y(ori_ori_n1039_));
  OR4        o1011(.A(ori_ori_n1039_), .B(ori_ori_n1035_), .C(ori_ori_n1032_), .D(ori_ori_n1031_), .Y(ori_ori_n1040_));
  NO4        o1012(.A(ori_ori_n1040_), .B(ori_ori_n1030_), .C(ori_ori_n1027_), .D(ori_ori_n1024_), .Y(ori_ori_n1041_));
  NA4        o1013(.A(ori_ori_n1041_), .B(ori_ori_n1017_), .C(ori_ori_n980_), .D(ori_ori_n967_), .Y(ori13));
  AN2        o1014(.A(c), .B(b), .Y(ori_ori_n1043_));
  NAi32      o1015(.An(d), .Bn(c), .C(e), .Y(ori_ori_n1044_));
  NA2        o1016(.A(ori_ori_n143_), .B(ori_ori_n45_), .Y(ori_ori_n1045_));
  NO4        o1017(.A(ori_ori_n1045_), .B(ori_ori_n1044_), .C(ori_ori_n612_), .D(ori_ori_n315_), .Y(ori_ori_n1046_));
  AN2        o1018(.A(d), .B(c), .Y(ori_ori_n1047_));
  NA2        o1019(.A(ori_ori_n1047_), .B(ori_ori_n118_), .Y(ori_ori_n1048_));
  NAi32      o1020(.An(f), .Bn(e), .C(c), .Y(ori_ori_n1049_));
  NOi41      o1021(.An(n), .B(m), .C(i), .D(h), .Y(ori_ori_n1050_));
  OR3        o1022(.A(e), .B(d), .C(c), .Y(ori_ori_n1051_));
  NA3        o1023(.A(k), .B(j), .C(i), .Y(ori_ori_n1052_));
  NO3        o1024(.A(ori_ori_n1052_), .B(ori_ori_n315_), .C(ori_ori_n91_), .Y(ori_ori_n1053_));
  NOi21      o1025(.An(ori_ori_n1053_), .B(ori_ori_n1051_), .Y(ori_ori_n1054_));
  NO2        o1026(.A(f), .B(c), .Y(ori_ori_n1055_));
  NOi21      o1027(.An(ori_ori_n1055_), .B(ori_ori_n457_), .Y(ori_ori_n1056_));
  NA2        o1028(.A(ori_ori_n1056_), .B(ori_ori_n59_), .Y(ori_ori_n1057_));
  OR2        o1029(.A(k), .B(i), .Y(ori_ori_n1058_));
  NO3        o1030(.A(ori_ori_n1058_), .B(ori_ori_n248_), .C(l), .Y(ori_ori_n1059_));
  NOi31      o1031(.An(ori_ori_n1059_), .B(ori_ori_n1057_), .C(j), .Y(ori_ori_n1060_));
  OR3        o1032(.A(ori_ori_n1060_), .B(ori_ori_n1054_), .C(ori_ori_n1046_), .Y(ori02));
  OR2        o1033(.A(l), .B(k), .Y(ori_ori_n1062_));
  OR3        o1034(.A(h), .B(g), .C(f), .Y(ori_ori_n1063_));
  OR3        o1035(.A(n), .B(m), .C(i), .Y(ori_ori_n1064_));
  NO4        o1036(.A(ori_ori_n1064_), .B(ori_ori_n1063_), .C(ori_ori_n1062_), .D(ori_ori_n1051_), .Y(ori_ori_n1065_));
  INV        o1037(.A(ori_ori_n1046_), .Y(ori_ori_n1066_));
  AN3        o1038(.A(g), .B(f), .C(c), .Y(ori_ori_n1067_));
  NA3        o1039(.A(l), .B(k), .C(j), .Y(ori_ori_n1068_));
  NA2        o1040(.A(i), .B(h), .Y(ori_ori_n1069_));
  NO3        o1041(.A(ori_ori_n1069_), .B(ori_ori_n1068_), .C(ori_ori_n134_), .Y(ori_ori_n1070_));
  NO3        o1042(.A(ori_ori_n145_), .B(ori_ori_n289_), .C(ori_ori_n219_), .Y(ori_ori_n1071_));
  NA3        o1043(.A(c), .B(b), .C(a), .Y(ori_ori_n1072_));
  NAi21      o1044(.An(ori_ori_n1065_), .B(ori_ori_n1066_), .Y(ori03));
  NO2        o1045(.A(ori_ori_n546_), .B(ori_ori_n621_), .Y(ori_ori_n1074_));
  NA4        o1046(.A(ori_ori_n88_), .B(ori_ori_n87_), .C(g), .D(ori_ori_n218_), .Y(ori_ori_n1075_));
  NA2        o1047(.A(ori_ori_n381_), .B(ori_ori_n1075_), .Y(ori_ori_n1076_));
  NO3        o1048(.A(ori_ori_n1076_), .B(ori_ori_n1074_), .C(ori_ori_n1011_), .Y(ori_ori_n1077_));
  NOi41      o1049(.An(ori_ori_n823_), .B(ori_ori_n870_), .C(ori_ori_n859_), .D(ori_ori_n739_), .Y(ori_ori_n1078_));
  OAI220     o1050(.A0(ori_ori_n1078_), .A1(ori_ori_n715_), .B0(ori_ori_n1077_), .B1(ori_ori_n609_), .Y(ori_ori_n1079_));
  NO2        o1051(.A(ori_ori_n838_), .B(ori_ori_n435_), .Y(ori_ori_n1080_));
  NOi31      o1052(.An(m), .B(n), .C(f), .Y(ori_ori_n1081_));
  NA2        o1053(.A(ori_ori_n1081_), .B(ori_ori_n51_), .Y(ori_ori_n1082_));
  AN2        o1054(.A(e), .B(c), .Y(ori_ori_n1083_));
  NA2        o1055(.A(ori_ori_n1083_), .B(a), .Y(ori_ori_n1084_));
  OAI220     o1056(.A0(ori_ori_n1084_), .A1(ori_ori_n1082_), .B0(ori_ori_n901_), .B1(ori_ori_n441_), .Y(ori_ori_n1085_));
  NA2        o1057(.A(ori_ori_n526_), .B(l), .Y(ori_ori_n1086_));
  NO3        o1058(.A(ori_ori_n1085_), .B(ori_ori_n1080_), .C(ori_ori_n1010_), .Y(ori_ori_n1087_));
  NO2        o1059(.A(ori_ori_n289_), .B(a), .Y(ori_ori_n1088_));
  INV        o1060(.A(ori_ori_n1046_), .Y(ori_ori_n1089_));
  NO2        o1061(.A(ori_ori_n87_), .B(g), .Y(ori_ori_n1090_));
  INV        o1062(.A(ori_ori_n1059_), .Y(ori_ori_n1091_));
  OR2        o1063(.A(ori_ori_n1091_), .B(ori_ori_n1057_), .Y(ori_ori_n1092_));
  NA3        o1064(.A(ori_ori_n1092_), .B(ori_ori_n1089_), .C(ori_ori_n1087_), .Y(ori_ori_n1093_));
  NO4        o1065(.A(ori_ori_n1093_), .B(ori_ori_n1079_), .C(ori_ori_n840_), .D(ori_ori_n585_), .Y(ori_ori_n1094_));
  NA2        o1066(.A(c), .B(b), .Y(ori_ori_n1095_));
  NO2        o1067(.A(ori_ori_n725_), .B(ori_ori_n1095_), .Y(ori_ori_n1096_));
  OAI210     o1068(.A0(ori_ori_n878_), .A1(ori_ori_n850_), .B0(ori_ori_n428_), .Y(ori_ori_n1097_));
  OAI210     o1069(.A0(ori_ori_n1097_), .A1(ori_ori_n879_), .B0(ori_ori_n1096_), .Y(ori_ori_n1098_));
  NAi21      o1070(.An(ori_ori_n436_), .B(ori_ori_n1096_), .Y(ori_ori_n1099_));
  NA3        o1071(.A(ori_ori_n442_), .B(ori_ori_n578_), .C(f), .Y(ori_ori_n1100_));
  OAI210     o1072(.A0(ori_ori_n567_), .A1(ori_ori_n39_), .B0(ori_ori_n1088_), .Y(ori_ori_n1101_));
  NA3        o1073(.A(ori_ori_n1101_), .B(ori_ori_n1100_), .C(ori_ori_n1099_), .Y(ori_ori_n1102_));
  NA2        o1074(.A(ori_ori_n267_), .B(ori_ori_n121_), .Y(ori_ori_n1103_));
  OAI210     o1075(.A0(ori_ori_n1103_), .A1(ori_ori_n293_), .B0(g), .Y(ori_ori_n1104_));
  NAi21      o1076(.An(f), .B(d), .Y(ori_ori_n1105_));
  NO2        o1077(.A(ori_ori_n1105_), .B(ori_ori_n1072_), .Y(ori_ori_n1106_));
  INV        o1078(.A(ori_ori_n1106_), .Y(ori_ori_n1107_));
  AOI210     o1079(.A0(ori_ori_n1104_), .A1(ori_ori_n299_), .B0(ori_ori_n1107_), .Y(ori_ori_n1108_));
  AOI210     o1080(.A0(ori_ori_n1108_), .A1(ori_ori_n115_), .B0(ori_ori_n1102_), .Y(ori_ori_n1109_));
  NA2        o1081(.A(ori_ori_n487_), .B(ori_ori_n486_), .Y(ori_ori_n1110_));
  NO2        o1082(.A(ori_ori_n187_), .B(ori_ori_n242_), .Y(ori_ori_n1111_));
  NA2        o1083(.A(ori_ori_n1111_), .B(m), .Y(ori_ori_n1112_));
  NA3        o1084(.A(ori_ori_n931_), .B(ori_ori_n1086_), .C(ori_ori_n490_), .Y(ori_ori_n1113_));
  OAI210     o1085(.A0(ori_ori_n1113_), .A1(ori_ori_n320_), .B0(ori_ori_n488_), .Y(ori_ori_n1114_));
  AOI210     o1086(.A0(ori_ori_n1114_), .A1(ori_ori_n1110_), .B0(ori_ori_n1112_), .Y(ori_ori_n1115_));
  NA2        o1087(.A(ori_ori_n580_), .B(ori_ori_n423_), .Y(ori_ori_n1116_));
  NA2        o1088(.A(ori_ori_n461_), .B(ori_ori_n1106_), .Y(ori_ori_n1117_));
  NO2        o1089(.A(ori_ori_n384_), .B(ori_ori_n383_), .Y(ori_ori_n1118_));
  NA2        o1090(.A(ori_ori_n1111_), .B(ori_ori_n444_), .Y(ori_ori_n1119_));
  NAi41      o1091(.An(ori_ori_n1118_), .B(ori_ori_n1119_), .C(ori_ori_n1117_), .D(ori_ori_n1116_), .Y(ori_ori_n1120_));
  NO2        o1092(.A(ori_ori_n1120_), .B(ori_ori_n1115_), .Y(ori_ori_n1121_));
  NA4        o1093(.A(ori_ori_n1121_), .B(ori_ori_n1109_), .C(ori_ori_n1098_), .D(ori_ori_n1094_), .Y(ori00));
  AOI210     o1094(.A0(ori_ori_n912_), .A1(ori_ori_n957_), .B0(ori_ori_n1080_), .Y(ori_ori_n1123_));
  NA2        o1095(.A(ori_ori_n1123_), .B(ori_ori_n1012_), .Y(ori_ori_n1124_));
  NA2        o1096(.A(ori_ori_n528_), .B(f), .Y(ori_ori_n1125_));
  OAI210     o1097(.A0(ori_ori_n1019_), .A1(ori_ori_n40_), .B0(ori_ori_n668_), .Y(ori_ori_n1126_));
  NA3        o1098(.A(ori_ori_n1126_), .B(ori_ori_n263_), .C(n), .Y(ori_ori_n1127_));
  AOI210     o1099(.A0(ori_ori_n1127_), .A1(ori_ori_n1125_), .B0(ori_ori_n1048_), .Y(ori_ori_n1128_));
  NO3        o1100(.A(ori_ori_n1128_), .B(ori_ori_n1124_), .C(ori_ori_n1054_), .Y(ori_ori_n1129_));
  NA3        o1101(.A(ori_ori_n172_), .B(ori_ori_n46_), .C(ori_ori_n45_), .Y(ori_ori_n1130_));
  NA3        o1102(.A(d), .B(ori_ori_n56_), .C(b), .Y(ori_ori_n1131_));
  NO2        o1103(.A(ori_ori_n1131_), .B(ori_ori_n1130_), .Y(ori_ori_n1132_));
  INV        o1104(.A(ori_ori_n598_), .Y(ori_ori_n1133_));
  NO3        o1105(.A(ori_ori_n1133_), .B(ori_ori_n1132_), .C(ori_ori_n1118_), .Y(ori_ori_n1134_));
  NO4        o1106(.A(ori_ori_n507_), .B(ori_ori_n366_), .C(ori_ori_n1095_), .D(ori_ori_n59_), .Y(ori_ori_n1135_));
  NA3        o1107(.A(ori_ori_n396_), .B(ori_ori_n226_), .C(g), .Y(ori_ori_n1136_));
  OA220      o1108(.A0(ori_ori_n1136_), .A1(ori_ori_n1131_), .B0(ori_ori_n397_), .B1(ori_ori_n137_), .Y(ori_ori_n1137_));
  NO2        o1109(.A(h), .B(g), .Y(ori_ori_n1138_));
  NA4        o1110(.A(ori_ori_n517_), .B(ori_ori_n484_), .C(ori_ori_n1138_), .D(ori_ori_n1043_), .Y(ori_ori_n1139_));
  NO2        o1111(.A(ori_ori_n92_), .B(ori_ori_n91_), .Y(ori_ori_n1140_));
  AOI220     o1112(.A0(ori_ori_n1140_), .A1(ori_ori_n554_), .B0(ori_ori_n962_), .B1(ori_ori_n597_), .Y(ori_ori_n1141_));
  AOI220     o1113(.A0(ori_ori_n327_), .A1(ori_ori_n252_), .B0(ori_ori_n182_), .B1(ori_ori_n152_), .Y(ori_ori_n1142_));
  NA4        o1114(.A(ori_ori_n1142_), .B(ori_ori_n1141_), .C(ori_ori_n1139_), .D(ori_ori_n1137_), .Y(ori_ori_n1143_));
  NO3        o1115(.A(ori_ori_n1143_), .B(ori_ori_n1135_), .C(ori_ori_n273_), .Y(ori_ori_n1144_));
  AOI210     o1116(.A0(ori_ori_n252_), .A1(ori_ori_n356_), .B0(ori_ori_n600_), .Y(ori_ori_n1145_));
  NA2        o1117(.A(ori_ori_n1145_), .B(ori_ori_n158_), .Y(ori_ori_n1146_));
  NO2        o1118(.A(ori_ori_n244_), .B(ori_ori_n186_), .Y(ori_ori_n1147_));
  NA2        o1119(.A(ori_ori_n1147_), .B(ori_ori_n442_), .Y(ori_ori_n1148_));
  NAi31      o1120(.An(ori_ori_n190_), .B(ori_ori_n876_), .C(ori_ori_n484_), .Y(ori_ori_n1149_));
  NA2        o1121(.A(ori_ori_n1149_), .B(ori_ori_n1148_), .Y(ori_ori_n1150_));
  NO4        o1122(.A(ori_ori_n1065_), .B(ori_ori_n1150_), .C(ori_ori_n1146_), .D(ori_ori_n538_), .Y(ori_ori_n1151_));
  AN3        o1123(.A(ori_ori_n1151_), .B(ori_ori_n1144_), .C(ori_ori_n1134_), .Y(ori_ori_n1152_));
  NA2        o1124(.A(ori_ori_n554_), .B(ori_ori_n102_), .Y(ori_ori_n1153_));
  NA3        o1125(.A(ori_ori_n1081_), .B(ori_ori_n630_), .C(ori_ori_n483_), .Y(ori_ori_n1154_));
  NA4        o1126(.A(ori_ori_n1154_), .B(ori_ori_n581_), .C(ori_ori_n1153_), .D(ori_ori_n246_), .Y(ori_ori_n1155_));
  NA2        o1127(.A(ori_ori_n1076_), .B(ori_ori_n554_), .Y(ori_ori_n1156_));
  NA4        o1128(.A(ori_ori_n671_), .B(ori_ori_n211_), .C(ori_ori_n226_), .D(ori_ori_n167_), .Y(ori_ori_n1157_));
  NA3        o1129(.A(ori_ori_n1157_), .B(ori_ori_n1156_), .C(ori_ori_n303_), .Y(ori_ori_n1158_));
  OAI210     o1130(.A0(ori_ori_n482_), .A1(ori_ori_n122_), .B0(ori_ori_n881_), .Y(ori_ori_n1159_));
  AOI220     o1131(.A0(ori_ori_n1159_), .A1(ori_ori_n1113_), .B0(ori_ori_n580_), .B1(ori_ori_n423_), .Y(ori_ori_n1160_));
  NA2        o1132(.A(n), .B(e), .Y(ori_ori_n1161_));
  NO2        o1133(.A(ori_ori_n1161_), .B(ori_ori_n150_), .Y(ori_ori_n1162_));
  NA2        o1134(.A(ori_ori_n1162_), .B(ori_ori_n281_), .Y(ori_ori_n1163_));
  OAI210     o1135(.A0(ori_ori_n367_), .A1(ori_ori_n321_), .B0(ori_ori_n463_), .Y(ori_ori_n1164_));
  NA3        o1136(.A(ori_ori_n1164_), .B(ori_ori_n1163_), .C(ori_ori_n1160_), .Y(ori_ori_n1165_));
  AOI210     o1137(.A0(ori_ori_n1162_), .A1(ori_ori_n867_), .B0(ori_ori_n839_), .Y(ori_ori_n1166_));
  AOI220     o1138(.A0(ori_ori_n971_), .A1(ori_ori_n597_), .B0(ori_ori_n671_), .B1(ori_ori_n249_), .Y(ori_ori_n1167_));
  NO2        o1139(.A(ori_ori_n68_), .B(h), .Y(ori_ori_n1168_));
  NA3        o1140(.A(ori_ori_n1167_), .B(ori_ori_n1166_), .C(ori_ori_n883_), .Y(ori_ori_n1169_));
  NO4        o1141(.A(ori_ori_n1169_), .B(ori_ori_n1165_), .C(ori_ori_n1158_), .D(ori_ori_n1155_), .Y(ori_ori_n1170_));
  NA2        o1142(.A(ori_ori_n851_), .B(ori_ori_n776_), .Y(ori_ori_n1171_));
  NA4        o1143(.A(ori_ori_n1171_), .B(ori_ori_n1170_), .C(ori_ori_n1152_), .D(ori_ori_n1129_), .Y(ori01));
  NO2        o1144(.A(ori_ori_n498_), .B(ori_ori_n287_), .Y(ori_ori_n1173_));
  NA2        o1145(.A(ori_ori_n407_), .B(i), .Y(ori_ori_n1174_));
  NA3        o1146(.A(ori_ori_n1174_), .B(ori_ori_n1173_), .C(ori_ori_n1033_), .Y(ori_ori_n1175_));
  NA2        o1147(.A(ori_ori_n610_), .B(ori_ori_n90_), .Y(ori_ori_n1176_));
  NA2        o1148(.A(ori_ori_n573_), .B(ori_ori_n278_), .Y(ori_ori_n1177_));
  NA2        o1149(.A(ori_ori_n976_), .B(ori_ori_n1177_), .Y(ori_ori_n1178_));
  NA4        o1150(.A(ori_ori_n1178_), .B(ori_ori_n1176_), .C(ori_ori_n927_), .D(ori_ori_n342_), .Y(ori_ori_n1179_));
  NA2        o1151(.A(ori_ori_n45_), .B(f), .Y(ori_ori_n1180_));
  NA2        o1152(.A(ori_ori_n732_), .B(ori_ori_n97_), .Y(ori_ori_n1181_));
  NO2        o1153(.A(ori_ori_n1181_), .B(ori_ori_n1180_), .Y(ori_ori_n1182_));
  OAI210     o1154(.A0(ori_ori_n803_), .A1(ori_ori_n625_), .B0(ori_ori_n1157_), .Y(ori_ori_n1183_));
  AOI210     o1155(.A0(ori_ori_n1182_), .A1(ori_ori_n658_), .B0(ori_ori_n1183_), .Y(ori_ori_n1184_));
  INV        o1156(.A(ori_ori_n120_), .Y(ori_ori_n1185_));
  OA220      o1157(.A0(ori_ori_n1185_), .A1(ori_ori_n607_), .B0(ori_ori_n683_), .B1(ori_ori_n381_), .Y(ori_ori_n1186_));
  NAi41      o1158(.An(ori_ori_n166_), .B(ori_ori_n1186_), .C(ori_ori_n1184_), .D(ori_ori_n911_), .Y(ori_ori_n1187_));
  NO2        o1159(.A(ori_ori_n699_), .B(ori_ori_n531_), .Y(ori_ori_n1188_));
  OR2        o1160(.A(ori_ori_n200_), .B(ori_ori_n198_), .Y(ori_ori_n1189_));
  NA3        o1161(.A(ori_ori_n1189_), .B(ori_ori_n1188_), .C(ori_ori_n140_), .Y(ori_ori_n1190_));
  NO4        o1162(.A(ori_ori_n1190_), .B(ori_ori_n1187_), .C(ori_ori_n1179_), .D(ori_ori_n1175_), .Y(ori_ori_n1191_));
  INV        o1163(.A(ori_ori_n1136_), .Y(ori_ori_n1192_));
  OAI210     o1164(.A0(ori_ori_n1192_), .A1(ori_ori_n309_), .B0(ori_ori_n550_), .Y(ori_ori_n1193_));
  NA2        o1165(.A(ori_ori_n557_), .B(ori_ori_n409_), .Y(ori_ori_n1194_));
  NOi21      o1166(.An(ori_ori_n582_), .B(ori_ori_n604_), .Y(ori_ori_n1195_));
  NA2        o1167(.A(ori_ori_n1195_), .B(ori_ori_n1194_), .Y(ori_ori_n1196_));
  AOI210     o1168(.A0(ori_ori_n209_), .A1(ori_ori_n89_), .B0(ori_ori_n218_), .Y(ori_ori_n1197_));
  OAI210     o1169(.A0(ori_ori_n826_), .A1(ori_ori_n442_), .B0(ori_ori_n1197_), .Y(ori_ori_n1198_));
  AN3        o1170(.A(m), .B(l), .C(k), .Y(ori_ori_n1199_));
  OAI210     o1171(.A0(ori_ori_n369_), .A1(ori_ori_n34_), .B0(ori_ori_n1199_), .Y(ori_ori_n1200_));
  NA2        o1172(.A(ori_ori_n208_), .B(ori_ori_n34_), .Y(ori_ori_n1201_));
  AO210      o1173(.A0(ori_ori_n1201_), .A1(ori_ori_n1200_), .B0(ori_ori_n341_), .Y(ori_ori_n1202_));
  NA4        o1174(.A(ori_ori_n1202_), .B(ori_ori_n1198_), .C(ori_ori_n1196_), .D(ori_ori_n1193_), .Y(ori_ori_n1203_));
  AOI210     o1175(.A0(ori_ori_n619_), .A1(ori_ori_n120_), .B0(ori_ori_n623_), .Y(ori_ori_n1204_));
  OAI210     o1176(.A0(ori_ori_n1185_), .A1(ori_ori_n616_), .B0(ori_ori_n1204_), .Y(ori_ori_n1205_));
  NA2        o1177(.A(ori_ori_n286_), .B(ori_ori_n200_), .Y(ori_ori_n1206_));
  NA2        o1178(.A(ori_ori_n1206_), .B(ori_ori_n688_), .Y(ori_ori_n1207_));
  NO3        o1179(.A(ori_ori_n838_), .B(ori_ori_n209_), .C(ori_ori_n421_), .Y(ori_ori_n1208_));
  INV        o1180(.A(ori_ori_n1208_), .Y(ori_ori_n1209_));
  OAI210     o1181(.A0(ori_ori_n1182_), .A1(ori_ori_n335_), .B0(ori_ori_n700_), .Y(ori_ori_n1210_));
  NA4        o1182(.A(ori_ori_n1210_), .B(ori_ori_n1209_), .C(ori_ori_n1207_), .D(ori_ori_n806_), .Y(ori_ori_n1211_));
  NO3        o1183(.A(ori_ori_n1211_), .B(ori_ori_n1205_), .C(ori_ori_n1203_), .Y(ori_ori_n1212_));
  NA3        o1184(.A(ori_ori_n626_), .B(ori_ori_n29_), .C(f), .Y(ori_ori_n1213_));
  NO2        o1185(.A(ori_ori_n1213_), .B(ori_ori_n209_), .Y(ori_ori_n1214_));
  AOI210     o1186(.A0(ori_ori_n524_), .A1(ori_ori_n58_), .B0(ori_ori_n1214_), .Y(ori_ori_n1215_));
  OR3        o1187(.A(ori_ori_n1181_), .B(ori_ori_n627_), .C(ori_ori_n1180_), .Y(ori_ori_n1216_));
  NO2        o1188(.A(ori_ori_n212_), .B(ori_ori_n113_), .Y(ori_ori_n1217_));
  NO2        o1189(.A(ori_ori_n1217_), .B(ori_ori_n1132_), .Y(ori_ori_n1218_));
  NA4        o1190(.A(ori_ori_n1218_), .B(ori_ori_n1216_), .C(ori_ori_n1215_), .D(ori_ori_n775_), .Y(ori_ori_n1219_));
  NO2        o1191(.A(ori_ori_n982_), .B(ori_ori_n238_), .Y(ori_ori_n1220_));
  NO2        o1192(.A(ori_ori_n983_), .B(ori_ori_n575_), .Y(ori_ori_n1221_));
  OAI210     o1193(.A0(ori_ori_n1221_), .A1(ori_ori_n1220_), .B0(ori_ori_n350_), .Y(ori_ori_n1222_));
  NA2        o1194(.A(ori_ori_n592_), .B(ori_ori_n590_), .Y(ori_ori_n1223_));
  NO3        o1195(.A(ori_ori_n79_), .B(ori_ori_n307_), .C(ori_ori_n45_), .Y(ori_ori_n1224_));
  NA2        o1196(.A(ori_ori_n1224_), .B(ori_ori_n572_), .Y(ori_ori_n1225_));
  NA3        o1197(.A(ori_ori_n1225_), .B(ori_ori_n1223_), .C(ori_ori_n694_), .Y(ori_ori_n1226_));
  OR2        o1198(.A(ori_ori_n1136_), .B(ori_ori_n1131_), .Y(ori_ori_n1227_));
  NO2        o1199(.A(ori_ori_n381_), .B(ori_ori_n72_), .Y(ori_ori_n1228_));
  INV        o1200(.A(ori_ori_n1228_), .Y(ori_ori_n1229_));
  NA2        o1201(.A(ori_ori_n1224_), .B(ori_ori_n829_), .Y(ori_ori_n1230_));
  NA4        o1202(.A(ori_ori_n1230_), .B(ori_ori_n1229_), .C(ori_ori_n1227_), .D(ori_ori_n399_), .Y(ori_ori_n1231_));
  NOi41      o1203(.An(ori_ori_n1222_), .B(ori_ori_n1231_), .C(ori_ori_n1226_), .D(ori_ori_n1219_), .Y(ori_ori_n1232_));
  NO2        o1204(.A(ori_ori_n133_), .B(ori_ori_n45_), .Y(ori_ori_n1233_));
  NO2        o1205(.A(ori_ori_n45_), .B(ori_ori_n40_), .Y(ori_ori_n1234_));
  AO220      o1206(.A0(ori_ori_n1234_), .A1(ori_ori_n645_), .B0(ori_ori_n1233_), .B1(ori_ori_n730_), .Y(ori_ori_n1235_));
  NA2        o1207(.A(ori_ori_n1235_), .B(ori_ori_n350_), .Y(ori_ori_n1236_));
  INV        o1208(.A(ori_ori_n137_), .Y(ori_ori_n1237_));
  NO3        o1209(.A(ori_ori_n1069_), .B(ori_ori_n181_), .C(ori_ori_n87_), .Y(ori_ori_n1238_));
  AOI220     o1210(.A0(ori_ori_n1238_), .A1(ori_ori_n1237_), .B0(ori_ori_n1224_), .B1(ori_ori_n986_), .Y(ori_ori_n1239_));
  NA2        o1211(.A(ori_ori_n1239_), .B(ori_ori_n1236_), .Y(ori_ori_n1240_));
  NO2        o1212(.A(ori_ori_n638_), .B(ori_ori_n637_), .Y(ori_ori_n1241_));
  NO4        o1213(.A(ori_ori_n1069_), .B(ori_ori_n1241_), .C(ori_ori_n179_), .D(ori_ori_n87_), .Y(ori_ori_n1242_));
  NO3        o1214(.A(ori_ori_n1242_), .B(ori_ori_n1240_), .C(ori_ori_n660_), .Y(ori_ori_n1243_));
  NA4        o1215(.A(ori_ori_n1243_), .B(ori_ori_n1232_), .C(ori_ori_n1212_), .D(ori_ori_n1191_), .Y(ori06));
  NO2        o1216(.A(ori_ori_n422_), .B(ori_ori_n579_), .Y(ori_ori_n1245_));
  NA2        o1217(.A(ori_ori_n274_), .B(ori_ori_n1245_), .Y(ori_ori_n1246_));
  NO2        o1218(.A(ori_ori_n230_), .B(ori_ori_n104_), .Y(ori_ori_n1247_));
  OAI210     o1219(.A0(ori_ori_n1247_), .A1(ori_ori_n1238_), .B0(ori_ori_n395_), .Y(ori_ori_n1248_));
  NO3        o1220(.A(ori_ori_n622_), .B(ori_ori_n824_), .C(ori_ori_n624_), .Y(ori_ori_n1249_));
  OR2        o1221(.A(ori_ori_n1249_), .B(ori_ori_n901_), .Y(ori_ori_n1250_));
  NA4        o1222(.A(ori_ori_n1250_), .B(ori_ori_n1248_), .C(ori_ori_n1246_), .D(ori_ori_n1222_), .Y(ori_ori_n1251_));
  NO3        o1223(.A(ori_ori_n1251_), .B(ori_ori_n1226_), .C(ori_ori_n262_), .Y(ori_ori_n1252_));
  NO2        o1224(.A(ori_ori_n307_), .B(ori_ori_n45_), .Y(ori_ori_n1253_));
  AOI210     o1225(.A0(ori_ori_n1253_), .A1(ori_ori_n987_), .B0(ori_ori_n1220_), .Y(ori_ori_n1254_));
  AOI210     o1226(.A0(ori_ori_n1253_), .A1(ori_ori_n576_), .B0(ori_ori_n1235_), .Y(ori_ori_n1255_));
  AOI210     o1227(.A0(ori_ori_n1255_), .A1(ori_ori_n1254_), .B0(ori_ori_n347_), .Y(ori_ori_n1256_));
  OAI210     o1228(.A0(ori_ori_n89_), .A1(ori_ori_n40_), .B0(ori_ori_n698_), .Y(ori_ori_n1257_));
  NA2        o1229(.A(ori_ori_n1257_), .B(ori_ori_n664_), .Y(ori_ori_n1258_));
  NO2        o1230(.A(ori_ori_n534_), .B(ori_ori_n176_), .Y(ori_ori_n1259_));
  NOi21      o1231(.An(ori_ori_n139_), .B(ori_ori_n45_), .Y(ori_ori_n1260_));
  NO2        o1232(.A(ori_ori_n631_), .B(ori_ori_n1082_), .Y(ori_ori_n1261_));
  OAI210     o1233(.A0(ori_ori_n477_), .A1(ori_ori_n253_), .B0(ori_ori_n922_), .Y(ori_ori_n1262_));
  NO4        o1234(.A(ori_ori_n1262_), .B(ori_ori_n1261_), .C(ori_ori_n1260_), .D(ori_ori_n1259_), .Y(ori_ori_n1263_));
  NO2        o1235(.A(ori_ori_n380_), .B(ori_ori_n138_), .Y(ori_ori_n1264_));
  AOI210     o1236(.A0(ori_ori_n1264_), .A1(ori_ori_n610_), .B0(ori_ori_n623_), .Y(ori_ori_n1265_));
  NA3        o1237(.A(ori_ori_n1265_), .B(ori_ori_n1263_), .C(ori_ori_n1258_), .Y(ori_ori_n1266_));
  NO2        o1238(.A(ori_ori_n767_), .B(ori_ori_n379_), .Y(ori_ori_n1267_));
  AN2        o1239(.A(ori_ori_n971_), .B(ori_ori_n667_), .Y(ori_ori_n1268_));
  NO3        o1240(.A(ori_ori_n1268_), .B(ori_ori_n1266_), .C(ori_ori_n1256_), .Y(ori_ori_n1269_));
  NO2        o1241(.A(ori_ori_n753_), .B(ori_ori_n47_), .Y(ori_ori_n1270_));
  NA2        o1242(.A(ori_ori_n372_), .B(ori_ori_n1270_), .Y(ori_ori_n1271_));
  NO3        o1243(.A(ori_ori_n248_), .B(ori_ori_n104_), .C(ori_ori_n289_), .Y(ori_ori_n1272_));
  OAI220     o1244(.A0(ori_ori_n722_), .A1(ori_ori_n253_), .B0(ori_ori_n530_), .B1(ori_ori_n534_), .Y(ori_ori_n1273_));
  NO3        o1245(.A(ori_ori_n1273_), .B(ori_ori_n1272_), .C(ori_ori_n1085_), .Y(ori_ori_n1274_));
  NA4        o1246(.A(ori_ori_n813_), .B(ori_ori_n812_), .C(ori_ori_n451_), .D(ori_ori_n893_), .Y(ori_ori_n1275_));
  NAi31      o1247(.An(ori_ori_n767_), .B(ori_ori_n1275_), .C(ori_ori_n208_), .Y(ori_ori_n1276_));
  NA4        o1248(.A(ori_ori_n1276_), .B(ori_ori_n1274_), .C(ori_ori_n1271_), .D(ori_ori_n1167_), .Y(ori_ori_n1277_));
  AOI210     o1249(.A0(ori_ori_n592_), .A1(ori_ori_n463_), .B0(ori_ori_n385_), .Y(ori_ori_n1278_));
  INV        o1250(.A(ori_ori_n1278_), .Y(ori_ori_n1279_));
  AOI220     o1251(.A0(ori_ori_n1267_), .A1(ori_ori_n776_), .B0(ori_ori_n1264_), .B1(ori_ori_n243_), .Y(ori_ori_n1280_));
  AN2        o1252(.A(ori_ori_n942_), .B(ori_ori_n941_), .Y(ori_ori_n1281_));
  NO3        o1253(.A(ori_ori_n1281_), .B(ori_ori_n520_), .C(ori_ori_n501_), .Y(ori_ori_n1282_));
  NA3        o1254(.A(ori_ori_n1282_), .B(ori_ori_n1280_), .C(ori_ori_n1230_), .Y(ori_ori_n1283_));
  NAi21      o1255(.An(j), .B(i), .Y(ori_ori_n1284_));
  NO4        o1256(.A(ori_ori_n1241_), .B(ori_ori_n1284_), .C(ori_ori_n457_), .D(ori_ori_n240_), .Y(ori_ori_n1285_));
  NO4        o1257(.A(ori_ori_n1285_), .B(ori_ori_n1283_), .C(ori_ori_n1279_), .D(ori_ori_n1277_), .Y(ori_ori_n1286_));
  NA4        o1258(.A(ori_ori_n1286_), .B(ori_ori_n1269_), .C(ori_ori_n1252_), .D(ori_ori_n1243_), .Y(ori07));
  NAi32      o1259(.An(m), .Bn(b), .C(n), .Y(ori_ori_n1288_));
  NO3        o1260(.A(ori_ori_n1288_), .B(g), .C(f), .Y(ori_ori_n1289_));
  NAi21      o1261(.An(f), .B(c), .Y(ori_ori_n1290_));
  OR2        o1262(.A(e), .B(d), .Y(ori_ori_n1291_));
  NOi31      o1263(.An(n), .B(m), .C(b), .Y(ori_ori_n1292_));
  NOi41      o1264(.An(i), .B(n), .C(m), .D(h), .Y(ori_ori_n1293_));
  NO2        o1265(.A(ori_ori_n1049_), .B(ori_ori_n457_), .Y(ori_ori_n1294_));
  NA2        o1266(.A(ori_ori_n1294_), .B(ori_ori_n219_), .Y(ori_ori_n1295_));
  NO2        o1267(.A(ori_ori_n1052_), .B(ori_ori_n315_), .Y(ori_ori_n1296_));
  NA2        o1268(.A(ori_ori_n560_), .B(ori_ori_n80_), .Y(ori_ori_n1297_));
  NA2        o1269(.A(ori_ori_n1168_), .B(ori_ori_n297_), .Y(ori_ori_n1298_));
  NA3        o1270(.A(ori_ori_n1298_), .B(ori_ori_n1297_), .C(ori_ori_n1295_), .Y(ori_ori_n1299_));
  NO2        o1271(.A(ori_ori_n1299_), .B(ori_ori_n1289_), .Y(ori_ori_n1300_));
  NO3        o1272(.A(e), .B(d), .C(c), .Y(ori_ori_n1301_));
  NO2        o1273(.A(ori_ori_n134_), .B(ori_ori_n219_), .Y(ori_ori_n1302_));
  NA2        o1274(.A(ori_ori_n1302_), .B(ori_ori_n1301_), .Y(ori_ori_n1303_));
  INV        o1275(.A(ori_ori_n1303_), .Y(ori_ori_n1304_));
  OR2        o1276(.A(h), .B(f), .Y(ori_ori_n1305_));
  NO3        o1277(.A(n), .B(m), .C(i), .Y(ori_ori_n1306_));
  NA2        o1278(.A(ori_ori_n161_), .B(ori_ori_n1306_), .Y(ori_ori_n1307_));
  NO2        o1279(.A(ori_ori_n1307_), .B(ori_ori_n1305_), .Y(ori_ori_n1308_));
  NA3        o1280(.A(ori_ori_n719_), .B(ori_ori_n707_), .C(ori_ori_n114_), .Y(ori_ori_n1309_));
  NO2        o1281(.A(ori_ori_n1309_), .B(ori_ori_n45_), .Y(ori_ori_n1310_));
  NO2        o1282(.A(l), .B(k), .Y(ori_ori_n1311_));
  NO3        o1283(.A(ori_ori_n457_), .B(d), .C(c), .Y(ori_ori_n1312_));
  NO3        o1284(.A(ori_ori_n1310_), .B(ori_ori_n1308_), .C(ori_ori_n1304_), .Y(ori_ori_n1313_));
  NO2        o1285(.A(ori_ori_n151_), .B(h), .Y(ori_ori_n1314_));
  NO2        o1286(.A(ori_ori_n1058_), .B(l), .Y(ori_ori_n1315_));
  NO2        o1287(.A(g), .B(c), .Y(ori_ori_n1316_));
  NA2        o1288(.A(ori_ori_n1316_), .B(ori_ori_n145_), .Y(ori_ori_n1317_));
  NO2        o1289(.A(ori_ori_n1317_), .B(ori_ori_n1315_), .Y(ori_ori_n1318_));
  NA2        o1290(.A(ori_ori_n1318_), .B(ori_ori_n184_), .Y(ori_ori_n1319_));
  NO2        o1291(.A(ori_ori_n468_), .B(a), .Y(ori_ori_n1320_));
  NA2        o1292(.A(ori_ori_n1320_), .B(ori_ori_n115_), .Y(ori_ori_n1321_));
  NO2        o1293(.A(i), .B(h), .Y(ori_ori_n1322_));
  NA2        o1294(.A(ori_ori_n141_), .B(ori_ori_n226_), .Y(ori_ori_n1323_));
  NO2        o1295(.A(ori_ori_n1323_), .B(ori_ori_n1430_), .Y(ori_ori_n1324_));
  NO2        o1296(.A(ori_ori_n773_), .B(ori_ori_n192_), .Y(ori_ori_n1325_));
  NOi31      o1297(.An(m), .B(n), .C(b), .Y(ori_ori_n1326_));
  NOi31      o1298(.An(f), .B(d), .C(c), .Y(ori_ori_n1327_));
  NA2        o1299(.A(ori_ori_n1327_), .B(ori_ori_n1326_), .Y(ori_ori_n1328_));
  INV        o1300(.A(ori_ori_n1328_), .Y(ori_ori_n1329_));
  NO3        o1301(.A(ori_ori_n1329_), .B(ori_ori_n1325_), .C(ori_ori_n1324_), .Y(ori_ori_n1330_));
  NA2        o1302(.A(ori_ori_n1067_), .B(ori_ori_n484_), .Y(ori_ori_n1331_));
  NO2        o1303(.A(ori_ori_n1331_), .B(ori_ori_n457_), .Y(ori_ori_n1332_));
  NO3        o1304(.A(ori_ori_n41_), .B(i), .C(h), .Y(ori_ori_n1333_));
  NO2        o1305(.A(ori_ori_n1050_), .B(ori_ori_n1332_), .Y(ori_ori_n1334_));
  AN4        o1306(.A(ori_ori_n1334_), .B(ori_ori_n1330_), .C(ori_ori_n1321_), .D(ori_ori_n1319_), .Y(ori_ori_n1335_));
  NA2        o1307(.A(ori_ori_n1292_), .B(ori_ori_n392_), .Y(ori_ori_n1336_));
  INV        o1308(.A(ori_ori_n1336_), .Y(ori_ori_n1337_));
  INV        o1309(.A(ori_ori_n1070_), .Y(ori_ori_n1338_));
  NAi21      o1310(.An(ori_ori_n1337_), .B(ori_ori_n1338_), .Y(ori_ori_n1339_));
  NO4        o1311(.A(ori_ori_n134_), .B(g), .C(f), .D(e), .Y(ori_ori_n1340_));
  NA2        o1312(.A(ori_ori_n199_), .B(ori_ori_n99_), .Y(ori_ori_n1341_));
  NA2        o1313(.A(ori_ori_n30_), .B(h), .Y(ori_ori_n1342_));
  NO2        o1314(.A(ori_ori_n1342_), .B(ori_ori_n1064_), .Y(ori_ori_n1343_));
  NA2        o1315(.A(ori_ori_n1293_), .B(ori_ori_n1311_), .Y(ori_ori_n1344_));
  INV        o1316(.A(ori_ori_n1344_), .Y(ori_ori_n1345_));
  OR3        o1317(.A(ori_ori_n559_), .B(ori_ori_n558_), .C(ori_ori_n114_), .Y(ori_ori_n1346_));
  NA2        o1318(.A(ori_ori_n1081_), .B(ori_ori_n421_), .Y(ori_ori_n1347_));
  NO2        o1319(.A(ori_ori_n1347_), .B(ori_ori_n450_), .Y(ori_ori_n1348_));
  AO210      o1320(.A0(ori_ori_n1348_), .A1(ori_ori_n118_), .B0(ori_ori_n1345_), .Y(ori_ori_n1349_));
  NO3        o1321(.A(ori_ori_n1349_), .B(ori_ori_n1343_), .C(ori_ori_n1339_), .Y(ori_ori_n1350_));
  NA4        o1322(.A(ori_ori_n1350_), .B(ori_ori_n1335_), .C(ori_ori_n1313_), .D(ori_ori_n1300_), .Y(ori_ori_n1351_));
  NO2        o1323(.A(ori_ori_n1095_), .B(ori_ori_n112_), .Y(ori_ori_n1352_));
  NA2        o1324(.A(ori_ori_n220_), .B(ori_ori_n184_), .Y(ori_ori_n1353_));
  NO2        o1325(.A(ori_ori_n404_), .B(j), .Y(ori_ori_n1354_));
  NA2        o1326(.A(ori_ori_n1333_), .B(ori_ori_n1081_), .Y(ori_ori_n1355_));
  NAi31      o1327(.An(ori_ori_n1322_), .B(ori_ori_n1056_), .C(ori_ori_n154_), .Y(ori_ori_n1356_));
  NA2        o1328(.A(ori_ori_n1356_), .B(ori_ori_n1355_), .Y(ori_ori_n1357_));
  NA2        o1329(.A(ori_ori_n1354_), .B(ori_ori_n163_), .Y(ori_ori_n1358_));
  INV        o1330(.A(ori_ori_n1358_), .Y(ori_ori_n1359_));
  NO2        o1331(.A(ori_ori_n1359_), .B(ori_ori_n1357_), .Y(ori_ori_n1360_));
  AOI210     o1332(.A0(ori_ori_n1353_), .A1(ori_ori_n1341_), .B0(ori_ori_n1049_), .Y(ori_ori_n1361_));
  OR2        o1333(.A(n), .B(i), .Y(ori_ori_n1362_));
  OAI210     o1334(.A0(ori_ori_n1362_), .A1(ori_ori_n1055_), .B0(ori_ori_n49_), .Y(ori_ori_n1363_));
  NA2        o1335(.A(ori_ori_n1363_), .B(ori_ori_n1138_), .Y(ori_ori_n1364_));
  INV        o1336(.A(ori_ori_n1364_), .Y(ori_ori_n1365_));
  NO2        o1337(.A(ori_ori_n689_), .B(ori_ori_n181_), .Y(ori_ori_n1366_));
  NO3        o1338(.A(ori_ori_n1366_), .B(ori_ori_n1365_), .C(ori_ori_n1361_), .Y(ori_ori_n1367_));
  NO3        o1339(.A(ori_ori_n1072_), .B(ori_ori_n1291_), .C(ori_ori_n49_), .Y(ori_ori_n1368_));
  NO2        o1340(.A(ori_ori_n1064_), .B(h), .Y(ori_ori_n1369_));
  NA2        o1341(.A(ori_ori_n1369_), .B(d), .Y(ori_ori_n1370_));
  INV        o1342(.A(ori_ori_n1370_), .Y(ori_ori_n1371_));
  NA3        o1343(.A(ori_ori_n1352_), .B(ori_ori_n484_), .C(f), .Y(ori_ori_n1372_));
  NO2        o1344(.A(ori_ori_n1428_), .B(ori_ori_n1372_), .Y(ori_ori_n1373_));
  NO2        o1345(.A(ori_ori_n1284_), .B(ori_ori_n179_), .Y(ori_ori_n1374_));
  NOi21      o1346(.An(d), .B(f), .Y(ori_ori_n1375_));
  NO2        o1347(.A(ori_ori_n1373_), .B(ori_ori_n1371_), .Y(ori_ori_n1376_));
  NA3        o1348(.A(ori_ori_n1376_), .B(ori_ori_n1367_), .C(ori_ori_n1360_), .Y(ori_ori_n1377_));
  NA2        o1349(.A(h), .B(ori_ori_n1296_), .Y(ori_ori_n1378_));
  OAI210     o1350(.A0(ori_ori_n1340_), .A1(ori_ori_n1292_), .B0(ori_ori_n898_), .Y(ori_ori_n1379_));
  NO2        o1351(.A(ori_ori_n1044_), .B(ori_ori_n134_), .Y(ori_ori_n1380_));
  NA2        o1352(.A(ori_ori_n1380_), .B(ori_ori_n644_), .Y(ori_ori_n1381_));
  NA3        o1353(.A(ori_ori_n1381_), .B(ori_ori_n1379_), .C(ori_ori_n1378_), .Y(ori_ori_n1382_));
  NA2        o1354(.A(ori_ori_n1316_), .B(ori_ori_n1375_), .Y(ori_ori_n1383_));
  NO2        o1355(.A(ori_ori_n1383_), .B(m), .Y(ori_ori_n1384_));
  NO2        o1356(.A(ori_ori_n155_), .B(ori_ori_n186_), .Y(ori_ori_n1385_));
  OAI210     o1357(.A0(ori_ori_n1385_), .A1(ori_ori_n112_), .B0(ori_ori_n1326_), .Y(ori_ori_n1386_));
  INV        o1358(.A(ori_ori_n1386_), .Y(ori_ori_n1387_));
  NO3        o1359(.A(ori_ori_n1387_), .B(ori_ori_n1384_), .C(ori_ori_n1382_), .Y(ori_ori_n1388_));
  NO2        o1360(.A(ori_ori_n1290_), .B(e), .Y(ori_ori_n1389_));
  NA2        o1361(.A(ori_ori_n1389_), .B(ori_ori_n419_), .Y(ori_ori_n1390_));
  BUFFER     o1362(.A(ori_ori_n134_), .Y(ori_ori_n1391_));
  NO2        o1363(.A(ori_ori_n1391_), .B(ori_ori_n1390_), .Y(ori_ori_n1392_));
  NO2        o1364(.A(ori_ori_n1346_), .B(ori_ori_n363_), .Y(ori_ori_n1393_));
  NO2        o1365(.A(ori_ori_n1393_), .B(ori_ori_n1392_), .Y(ori_ori_n1394_));
  NA2        o1366(.A(ori_ori_n1389_), .B(ori_ori_n184_), .Y(ori_ori_n1395_));
  AOI220     o1367(.A0(ori_ori_n1395_), .A1(ori_ori_n1057_), .B0(ori_ori_n551_), .B1(ori_ori_n379_), .Y(ori_ori_n1396_));
  AOI210     o1368(.A0(i), .A1(ori_ori_n1312_), .B0(ori_ori_n1368_), .Y(ori_ori_n1397_));
  INV        o1369(.A(ori_ori_n1090_), .Y(ori_ori_n1398_));
  OAI210     o1370(.A0(ori_ori_n1398_), .A1(ori_ori_n69_), .B0(ori_ori_n1397_), .Y(ori_ori_n1399_));
  OR2        o1371(.A(h), .B(ori_ori_n558_), .Y(ori_ori_n1400_));
  NO2        o1372(.A(ori_ori_n1400_), .B(ori_ori_n179_), .Y(ori_ori_n1401_));
  NA2        o1373(.A(ori_ori_n1071_), .B(ori_ori_n226_), .Y(ori_ori_n1402_));
  NO2        o1374(.A(ori_ori_n49_), .B(l), .Y(ori_ori_n1403_));
  INV        o1375(.A(ori_ori_n503_), .Y(ori_ori_n1404_));
  NA2        o1376(.A(ori_ori_n1404_), .B(ori_ori_n1403_), .Y(ori_ori_n1405_));
  NO2        o1377(.A(m), .B(i), .Y(ori_ori_n1406_));
  BUFFER     o1378(.A(ori_ori_n1406_), .Y(ori_ori_n1407_));
  NA2        o1379(.A(ori_ori_n1407_), .B(ori_ori_n1314_), .Y(ori_ori_n1408_));
  NA3        o1380(.A(ori_ori_n1408_), .B(ori_ori_n1405_), .C(ori_ori_n1402_), .Y(ori_ori_n1409_));
  NO4        o1381(.A(ori_ori_n1409_), .B(ori_ori_n1401_), .C(ori_ori_n1399_), .D(ori_ori_n1396_), .Y(ori_ori_n1410_));
  NA3        o1382(.A(ori_ori_n1410_), .B(ori_ori_n1394_), .C(ori_ori_n1388_), .Y(ori_ori_n1411_));
  NA3        o1383(.A(ori_ori_n975_), .B(ori_ori_n141_), .C(ori_ori_n46_), .Y(ori_ori_n1412_));
  INV        o1384(.A(ori_ori_n1412_), .Y(ori_ori_n1413_));
  NA2        o1385(.A(c), .B(ori_ori_n1369_), .Y(ori_ori_n1414_));
  NA2        o1386(.A(ori_ori_n1374_), .B(h), .Y(ori_ori_n1415_));
  NA2        o1387(.A(ori_ori_n1415_), .B(ori_ori_n1414_), .Y(ori_ori_n1416_));
  NO2        o1388(.A(ori_ori_n1416_), .B(ori_ori_n1413_), .Y(ori_ori_n1417_));
  AOI220     o1389(.A0(ori_ori_n1406_), .A1(ori_ori_n662_), .B0(ori_ori_n1431_), .B1(ori_ori_n164_), .Y(ori_ori_n1418_));
  NOi31      o1390(.An(ori_ori_n30_), .B(ori_ori_n1418_), .C(n), .Y(ori_ori_n1419_));
  INV        o1391(.A(ori_ori_n1419_), .Y(ori_ori_n1420_));
  NO2        o1392(.A(ori_ori_n1347_), .B(d), .Y(ori_ori_n1421_));
  NA3        o1393(.A(ori_ori_n1429_), .B(ori_ori_n1420_), .C(ori_ori_n1417_), .Y(ori_ori_n1422_));
  OR4        o1394(.A(ori_ori_n1422_), .B(ori_ori_n1411_), .C(ori_ori_n1377_), .D(ori_ori_n1351_), .Y(ori04));
  INV        o1395(.A(ori_ori_n1046_), .Y(ori_ori_n1424_));
  NA2        o1396(.A(ori_ori_n1424_), .B(ori_ori_n1092_), .Y(ori05));
  INV        o1397(.A(ori_ori_n115_), .Y(ori_ori_n1428_));
  INV        o1398(.A(ori_ori_n1421_), .Y(ori_ori_n1429_));
  INV        o1399(.A(h), .Y(ori_ori_n1430_));
  INV        o1400(.A(j), .Y(ori_ori_n1431_));
  AN2        m0000(.A(b), .B(a), .Y(mai_mai_n29_));
  NO2        m0001(.A(d), .B(c), .Y(mai_mai_n30_));
  AN2        m0002(.A(f), .B(e), .Y(mai_mai_n31_));
  NA3        m0003(.A(mai_mai_n31_), .B(mai_mai_n30_), .C(mai_mai_n29_), .Y(mai_mai_n32_));
  NOi32      m0004(.An(m), .Bn(l), .C(n), .Y(mai_mai_n33_));
  NOi32      m0005(.An(i), .Bn(g), .C(h), .Y(mai_mai_n34_));
  NA2        m0006(.A(mai_mai_n34_), .B(mai_mai_n33_), .Y(mai_mai_n35_));
  AN2        m0007(.A(m), .B(l), .Y(mai_mai_n36_));
  NOi32      m0008(.An(j), .Bn(g), .C(k), .Y(mai_mai_n37_));
  NA2        m0009(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n38_));
  NO2        m0010(.A(mai_mai_n38_), .B(n), .Y(mai_mai_n39_));
  INV        m0011(.A(h), .Y(mai_mai_n40_));
  NAi21      m0012(.An(j), .B(l), .Y(mai_mai_n41_));
  NAi32      m0013(.An(n), .Bn(g), .C(m), .Y(mai_mai_n42_));
  NO3        m0014(.A(mai_mai_n42_), .B(mai_mai_n41_), .C(mai_mai_n40_), .Y(mai_mai_n43_));
  NAi31      m0015(.An(n), .B(m), .C(l), .Y(mai_mai_n44_));
  INV        m0016(.A(i), .Y(mai_mai_n45_));
  AN2        m0017(.A(h), .B(g), .Y(mai_mai_n46_));
  NA2        m0018(.A(mai_mai_n46_), .B(mai_mai_n45_), .Y(mai_mai_n47_));
  NO2        m0019(.A(mai_mai_n47_), .B(mai_mai_n44_), .Y(mai_mai_n48_));
  NAi21      m0020(.An(n), .B(m), .Y(mai_mai_n49_));
  NOi32      m0021(.An(k), .Bn(h), .C(l), .Y(mai_mai_n50_));
  NOi32      m0022(.An(k), .Bn(h), .C(g), .Y(mai_mai_n51_));
  INV        m0023(.A(mai_mai_n51_), .Y(mai_mai_n52_));
  NO2        m0024(.A(mai_mai_n52_), .B(mai_mai_n49_), .Y(mai_mai_n53_));
  NO2        m0025(.A(mai_mai_n53_), .B(mai_mai_n43_), .Y(mai_mai_n54_));
  NO2        m0026(.A(mai_mai_n54_), .B(mai_mai_n32_), .Y(mai_mai_n55_));
  INV        m0027(.A(c), .Y(mai_mai_n56_));
  NA2        m0028(.A(e), .B(b), .Y(mai_mai_n57_));
  NO2        m0029(.A(mai_mai_n57_), .B(mai_mai_n56_), .Y(mai_mai_n58_));
  INV        m0030(.A(d), .Y(mai_mai_n59_));
  NAi21      m0031(.An(i), .B(h), .Y(mai_mai_n60_));
  NAi31      m0032(.An(i), .B(l), .C(j), .Y(mai_mai_n61_));
  NAi41      m0033(.An(e), .B(d), .C(b), .D(a), .Y(mai_mai_n62_));
  NA2        m0034(.A(g), .B(f), .Y(mai_mai_n63_));
  NO2        m0035(.A(mai_mai_n63_), .B(mai_mai_n62_), .Y(mai_mai_n64_));
  NAi21      m0036(.An(i), .B(j), .Y(mai_mai_n65_));
  NAi32      m0037(.An(n), .Bn(k), .C(m), .Y(mai_mai_n66_));
  NO2        m0038(.A(mai_mai_n66_), .B(mai_mai_n65_), .Y(mai_mai_n67_));
  NAi31      m0039(.An(l), .B(m), .C(k), .Y(mai_mai_n68_));
  NAi21      m0040(.An(e), .B(h), .Y(mai_mai_n69_));
  NAi41      m0041(.An(n), .B(d), .C(b), .D(a), .Y(mai_mai_n70_));
  NA2        m0042(.A(mai_mai_n67_), .B(mai_mai_n64_), .Y(mai_mai_n71_));
  INV        m0043(.A(m), .Y(mai_mai_n72_));
  NOi21      m0044(.An(k), .B(l), .Y(mai_mai_n73_));
  NA2        m0045(.A(mai_mai_n73_), .B(mai_mai_n72_), .Y(mai_mai_n74_));
  AN4        m0046(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n75_));
  NOi31      m0047(.An(h), .B(g), .C(f), .Y(mai_mai_n76_));
  NA2        m0048(.A(mai_mai_n76_), .B(mai_mai_n75_), .Y(mai_mai_n77_));
  NAi32      m0049(.An(m), .Bn(k), .C(j), .Y(mai_mai_n78_));
  NOi32      m0050(.An(h), .Bn(g), .C(f), .Y(mai_mai_n79_));
  NA2        m0051(.A(mai_mai_n79_), .B(mai_mai_n75_), .Y(mai_mai_n80_));
  OA220      m0052(.A0(mai_mai_n80_), .A1(mai_mai_n78_), .B0(mai_mai_n77_), .B1(mai_mai_n74_), .Y(mai_mai_n81_));
  NA2        m0053(.A(mai_mai_n81_), .B(mai_mai_n71_), .Y(mai_mai_n82_));
  INV        m0054(.A(n), .Y(mai_mai_n83_));
  NOi32      m0055(.An(e), .Bn(b), .C(d), .Y(mai_mai_n84_));
  NA2        m0056(.A(mai_mai_n84_), .B(mai_mai_n83_), .Y(mai_mai_n85_));
  INV        m0057(.A(j), .Y(mai_mai_n86_));
  AN3        m0058(.A(m), .B(k), .C(i), .Y(mai_mai_n87_));
  NA3        m0059(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(g), .Y(mai_mai_n88_));
  NAi32      m0060(.An(g), .Bn(f), .C(h), .Y(mai_mai_n89_));
  NAi31      m0061(.An(j), .B(m), .C(l), .Y(mai_mai_n90_));
  NO2        m0062(.A(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  NA2        m0063(.A(m), .B(l), .Y(mai_mai_n92_));
  NAi31      m0064(.An(k), .B(j), .C(g), .Y(mai_mai_n93_));
  NO3        m0065(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(f), .Y(mai_mai_n94_));
  AN2        m0066(.A(j), .B(g), .Y(mai_mai_n95_));
  NOi32      m0067(.An(m), .Bn(l), .C(i), .Y(mai_mai_n96_));
  NOi21      m0068(.An(g), .B(i), .Y(mai_mai_n97_));
  NOi32      m0069(.An(m), .Bn(j), .C(k), .Y(mai_mai_n98_));
  AOI220     m0070(.A0(mai_mai_n98_), .A1(mai_mai_n97_), .B0(mai_mai_n96_), .B1(mai_mai_n95_), .Y(mai_mai_n99_));
  NO2        m0071(.A(mai_mai_n99_), .B(f), .Y(mai_mai_n100_));
  NO3        m0072(.A(mai_mai_n100_), .B(mai_mai_n94_), .C(mai_mai_n91_), .Y(mai_mai_n101_));
  NAi41      m0073(.An(m), .B(n), .C(k), .D(i), .Y(mai_mai_n102_));
  AN2        m0074(.A(e), .B(b), .Y(mai_mai_n103_));
  NOi31      m0075(.An(c), .B(h), .C(f), .Y(mai_mai_n104_));
  NA2        m0076(.A(mai_mai_n104_), .B(mai_mai_n103_), .Y(mai_mai_n105_));
  NO2        m0077(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n106_));
  NOi21      m0078(.An(g), .B(f), .Y(mai_mai_n107_));
  NOi21      m0079(.An(i), .B(h), .Y(mai_mai_n108_));
  NA3        m0080(.A(mai_mai_n108_), .B(mai_mai_n107_), .C(mai_mai_n36_), .Y(mai_mai_n109_));
  INV        m0081(.A(a), .Y(mai_mai_n110_));
  NA2        m0082(.A(mai_mai_n103_), .B(mai_mai_n110_), .Y(mai_mai_n111_));
  INV        m0083(.A(l), .Y(mai_mai_n112_));
  NOi21      m0084(.An(m), .B(n), .Y(mai_mai_n113_));
  AN2        m0085(.A(k), .B(h), .Y(mai_mai_n114_));
  NO2        m0086(.A(mai_mai_n109_), .B(mai_mai_n85_), .Y(mai_mai_n115_));
  INV        m0087(.A(b), .Y(mai_mai_n116_));
  NA2        m0088(.A(l), .B(j), .Y(mai_mai_n117_));
  AN2        m0089(.A(k), .B(i), .Y(mai_mai_n118_));
  NA2        m0090(.A(mai_mai_n118_), .B(mai_mai_n117_), .Y(mai_mai_n119_));
  NA2        m0091(.A(g), .B(e), .Y(mai_mai_n120_));
  NOi32      m0092(.An(c), .Bn(a), .C(d), .Y(mai_mai_n121_));
  NA2        m0093(.A(mai_mai_n121_), .B(mai_mai_n113_), .Y(mai_mai_n122_));
  NO4        m0094(.A(mai_mai_n122_), .B(mai_mai_n120_), .C(mai_mai_n119_), .D(mai_mai_n116_), .Y(mai_mai_n123_));
  NO3        m0095(.A(mai_mai_n123_), .B(mai_mai_n115_), .C(mai_mai_n106_), .Y(mai_mai_n124_));
  OAI210     m0096(.A0(mai_mai_n101_), .A1(mai_mai_n85_), .B0(mai_mai_n124_), .Y(mai_mai_n125_));
  NOi31      m0097(.An(k), .B(m), .C(j), .Y(mai_mai_n126_));
  NA3        m0098(.A(mai_mai_n126_), .B(mai_mai_n76_), .C(mai_mai_n75_), .Y(mai_mai_n127_));
  NOi31      m0099(.An(k), .B(m), .C(i), .Y(mai_mai_n128_));
  NA3        m0100(.A(mai_mai_n128_), .B(mai_mai_n79_), .C(mai_mai_n75_), .Y(mai_mai_n129_));
  NA2        m0101(.A(mai_mai_n129_), .B(mai_mai_n127_), .Y(mai_mai_n130_));
  NOi32      m0102(.An(f), .Bn(b), .C(e), .Y(mai_mai_n131_));
  NAi21      m0103(.An(g), .B(h), .Y(mai_mai_n132_));
  NAi21      m0104(.An(m), .B(n), .Y(mai_mai_n133_));
  NAi21      m0105(.An(j), .B(k), .Y(mai_mai_n134_));
  NO3        m0106(.A(mai_mai_n134_), .B(mai_mai_n133_), .C(mai_mai_n132_), .Y(mai_mai_n135_));
  NAi41      m0107(.An(e), .B(f), .C(d), .D(b), .Y(mai_mai_n136_));
  NAi31      m0108(.An(j), .B(k), .C(h), .Y(mai_mai_n137_));
  NA2        m0109(.A(mai_mai_n135_), .B(mai_mai_n131_), .Y(mai_mai_n138_));
  NO2        m0110(.A(k), .B(j), .Y(mai_mai_n139_));
  NO2        m0111(.A(mai_mai_n139_), .B(mai_mai_n133_), .Y(mai_mai_n140_));
  AN2        m0112(.A(k), .B(j), .Y(mai_mai_n141_));
  NAi21      m0113(.An(c), .B(b), .Y(mai_mai_n142_));
  NA2        m0114(.A(f), .B(d), .Y(mai_mai_n143_));
  NO4        m0115(.A(mai_mai_n143_), .B(mai_mai_n142_), .C(mai_mai_n141_), .D(mai_mai_n132_), .Y(mai_mai_n144_));
  NA2        m0116(.A(h), .B(c), .Y(mai_mai_n145_));
  NAi31      m0117(.An(f), .B(e), .C(b), .Y(mai_mai_n146_));
  NA2        m0118(.A(mai_mai_n144_), .B(mai_mai_n140_), .Y(mai_mai_n147_));
  NA2        m0119(.A(d), .B(b), .Y(mai_mai_n148_));
  NAi21      m0120(.An(e), .B(f), .Y(mai_mai_n149_));
  NO2        m0121(.A(mai_mai_n149_), .B(mai_mai_n148_), .Y(mai_mai_n150_));
  NA2        m0122(.A(b), .B(a), .Y(mai_mai_n151_));
  NAi21      m0123(.An(e), .B(g), .Y(mai_mai_n152_));
  NAi21      m0124(.An(c), .B(d), .Y(mai_mai_n153_));
  NAi31      m0125(.An(l), .B(k), .C(h), .Y(mai_mai_n154_));
  NO2        m0126(.A(mai_mai_n133_), .B(mai_mai_n154_), .Y(mai_mai_n155_));
  NAi31      m0127(.An(mai_mai_n130_), .B(mai_mai_n147_), .C(mai_mai_n138_), .Y(mai_mai_n156_));
  NAi31      m0128(.An(e), .B(f), .C(b), .Y(mai_mai_n157_));
  NOi21      m0129(.An(g), .B(d), .Y(mai_mai_n158_));
  NO2        m0130(.A(mai_mai_n158_), .B(mai_mai_n157_), .Y(mai_mai_n159_));
  NOi21      m0131(.An(h), .B(i), .Y(mai_mai_n160_));
  NOi21      m0132(.An(k), .B(m), .Y(mai_mai_n161_));
  NA3        m0133(.A(mai_mai_n161_), .B(mai_mai_n160_), .C(n), .Y(mai_mai_n162_));
  NOi21      m0134(.An(mai_mai_n159_), .B(mai_mai_n162_), .Y(mai_mai_n163_));
  NOi21      m0135(.An(h), .B(g), .Y(mai_mai_n164_));
  NO2        m0136(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n165_));
  NA2        m0137(.A(mai_mai_n165_), .B(mai_mai_n164_), .Y(mai_mai_n166_));
  NAi31      m0138(.An(l), .B(j), .C(h), .Y(mai_mai_n167_));
  NOi32      m0139(.An(n), .Bn(k), .C(m), .Y(mai_mai_n168_));
  NA2        m0140(.A(l), .B(i), .Y(mai_mai_n169_));
  NA2        m0141(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  NO2        m0142(.A(mai_mai_n170_), .B(mai_mai_n166_), .Y(mai_mai_n171_));
  NAi31      m0143(.An(d), .B(f), .C(c), .Y(mai_mai_n172_));
  NAi31      m0144(.An(e), .B(f), .C(c), .Y(mai_mai_n173_));
  NA2        m0145(.A(mai_mai_n173_), .B(mai_mai_n172_), .Y(mai_mai_n174_));
  NA2        m0146(.A(j), .B(h), .Y(mai_mai_n175_));
  OR3        m0147(.A(n), .B(m), .C(k), .Y(mai_mai_n176_));
  NO2        m0148(.A(mai_mai_n176_), .B(mai_mai_n175_), .Y(mai_mai_n177_));
  NAi32      m0149(.An(m), .Bn(k), .C(n), .Y(mai_mai_n178_));
  NO2        m0150(.A(mai_mai_n178_), .B(mai_mai_n175_), .Y(mai_mai_n179_));
  AOI220     m0151(.A0(mai_mai_n179_), .A1(mai_mai_n159_), .B0(mai_mai_n177_), .B1(mai_mai_n174_), .Y(mai_mai_n180_));
  NO2        m0152(.A(n), .B(m), .Y(mai_mai_n181_));
  NA2        m0153(.A(mai_mai_n181_), .B(mai_mai_n50_), .Y(mai_mai_n182_));
  NAi21      m0154(.An(f), .B(e), .Y(mai_mai_n183_));
  NA2        m0155(.A(d), .B(c), .Y(mai_mai_n184_));
  NO2        m0156(.A(mai_mai_n184_), .B(mai_mai_n183_), .Y(mai_mai_n185_));
  NOi21      m0157(.An(mai_mai_n185_), .B(mai_mai_n182_), .Y(mai_mai_n186_));
  NAi21      m0158(.An(d), .B(c), .Y(mai_mai_n187_));
  NAi31      m0159(.An(m), .B(n), .C(b), .Y(mai_mai_n188_));
  NA2        m0160(.A(k), .B(i), .Y(mai_mai_n189_));
  NAi21      m0161(.An(h), .B(f), .Y(mai_mai_n190_));
  NO2        m0162(.A(mai_mai_n190_), .B(mai_mai_n189_), .Y(mai_mai_n191_));
  NO2        m0163(.A(mai_mai_n188_), .B(mai_mai_n153_), .Y(mai_mai_n192_));
  NA2        m0164(.A(mai_mai_n192_), .B(mai_mai_n191_), .Y(mai_mai_n193_));
  NOi32      m0165(.An(f), .Bn(c), .C(d), .Y(mai_mai_n194_));
  NOi32      m0166(.An(f), .Bn(c), .C(e), .Y(mai_mai_n195_));
  NO2        m0167(.A(mai_mai_n195_), .B(mai_mai_n194_), .Y(mai_mai_n196_));
  NO3        m0168(.A(n), .B(m), .C(j), .Y(mai_mai_n197_));
  NA2        m0169(.A(mai_mai_n197_), .B(mai_mai_n114_), .Y(mai_mai_n198_));
  AO210      m0170(.A0(mai_mai_n198_), .A1(mai_mai_n182_), .B0(mai_mai_n196_), .Y(mai_mai_n199_));
  NAi41      m0171(.An(mai_mai_n186_), .B(mai_mai_n199_), .C(mai_mai_n193_), .D(mai_mai_n180_), .Y(mai_mai_n200_));
  OR4        m0172(.A(mai_mai_n200_), .B(mai_mai_n171_), .C(mai_mai_n163_), .D(mai_mai_n156_), .Y(mai_mai_n201_));
  NO4        m0173(.A(mai_mai_n201_), .B(mai_mai_n125_), .C(mai_mai_n82_), .D(mai_mai_n55_), .Y(mai_mai_n202_));
  NA3        m0174(.A(m), .B(mai_mai_n112_), .C(j), .Y(mai_mai_n203_));
  NAi31      m0175(.An(n), .B(h), .C(g), .Y(mai_mai_n204_));
  NO2        m0176(.A(mai_mai_n204_), .B(mai_mai_n203_), .Y(mai_mai_n205_));
  NOi32      m0177(.An(m), .Bn(k), .C(l), .Y(mai_mai_n206_));
  NA3        m0178(.A(mai_mai_n206_), .B(mai_mai_n86_), .C(g), .Y(mai_mai_n207_));
  NO2        m0179(.A(mai_mai_n207_), .B(n), .Y(mai_mai_n208_));
  NOi21      m0180(.An(k), .B(j), .Y(mai_mai_n209_));
  NA4        m0181(.A(mai_mai_n209_), .B(mai_mai_n113_), .C(i), .D(g), .Y(mai_mai_n210_));
  AN2        m0182(.A(i), .B(g), .Y(mai_mai_n211_));
  NA3        m0183(.A(mai_mai_n73_), .B(mai_mai_n211_), .C(mai_mai_n113_), .Y(mai_mai_n212_));
  NA2        m0184(.A(mai_mai_n212_), .B(mai_mai_n210_), .Y(mai_mai_n213_));
  NO2        m0185(.A(mai_mai_n213_), .B(mai_mai_n205_), .Y(mai_mai_n214_));
  NAi41      m0186(.An(d), .B(n), .C(e), .D(b), .Y(mai_mai_n215_));
  INV        m0187(.A(mai_mai_n215_), .Y(mai_mai_n216_));
  INV        m0188(.A(f), .Y(mai_mai_n217_));
  INV        m0189(.A(g), .Y(mai_mai_n218_));
  NOi31      m0190(.An(i), .B(j), .C(h), .Y(mai_mai_n219_));
  NOi21      m0191(.An(l), .B(m), .Y(mai_mai_n220_));
  NA2        m0192(.A(mai_mai_n220_), .B(mai_mai_n219_), .Y(mai_mai_n221_));
  NO3        m0193(.A(mai_mai_n221_), .B(mai_mai_n218_), .C(mai_mai_n217_), .Y(mai_mai_n222_));
  NA2        m0194(.A(mai_mai_n222_), .B(mai_mai_n216_), .Y(mai_mai_n223_));
  OAI210     m0195(.A0(mai_mai_n214_), .A1(mai_mai_n32_), .B0(mai_mai_n223_), .Y(mai_mai_n224_));
  NOi21      m0196(.An(n), .B(m), .Y(mai_mai_n225_));
  NOi32      m0197(.An(l), .Bn(i), .C(j), .Y(mai_mai_n226_));
  NA2        m0198(.A(mai_mai_n226_), .B(mai_mai_n225_), .Y(mai_mai_n227_));
  OA220      m0199(.A0(mai_mai_n227_), .A1(mai_mai_n105_), .B0(mai_mai_n78_), .B1(mai_mai_n77_), .Y(mai_mai_n228_));
  NAi21      m0200(.An(j), .B(h), .Y(mai_mai_n229_));
  XN2        m0201(.A(i), .B(h), .Y(mai_mai_n230_));
  NA2        m0202(.A(mai_mai_n230_), .B(mai_mai_n229_), .Y(mai_mai_n231_));
  NOi31      m0203(.An(k), .B(n), .C(m), .Y(mai_mai_n232_));
  NOi31      m0204(.An(mai_mai_n232_), .B(mai_mai_n184_), .C(mai_mai_n183_), .Y(mai_mai_n233_));
  NA2        m0205(.A(mai_mai_n233_), .B(mai_mai_n231_), .Y(mai_mai_n234_));
  NAi31      m0206(.An(f), .B(e), .C(c), .Y(mai_mai_n235_));
  NO4        m0207(.A(mai_mai_n235_), .B(mai_mai_n176_), .C(mai_mai_n175_), .D(mai_mai_n59_), .Y(mai_mai_n236_));
  NA4        m0208(.A(n), .B(e), .C(c), .D(b), .Y(mai_mai_n237_));
  NAi32      m0209(.An(m), .Bn(i), .C(k), .Y(mai_mai_n238_));
  NO3        m0210(.A(mai_mai_n238_), .B(mai_mai_n89_), .C(mai_mai_n237_), .Y(mai_mai_n239_));
  INV        m0211(.A(k), .Y(mai_mai_n240_));
  NO2        m0212(.A(mai_mai_n239_), .B(mai_mai_n236_), .Y(mai_mai_n241_));
  NAi21      m0213(.An(n), .B(a), .Y(mai_mai_n242_));
  NO2        m0214(.A(mai_mai_n242_), .B(mai_mai_n148_), .Y(mai_mai_n243_));
  NAi41      m0215(.An(g), .B(m), .C(k), .D(h), .Y(mai_mai_n244_));
  NO2        m0216(.A(mai_mai_n244_), .B(e), .Y(mai_mai_n245_));
  NO3        m0217(.A(mai_mai_n149_), .B(mai_mai_n93_), .C(mai_mai_n92_), .Y(mai_mai_n246_));
  OAI210     m0218(.A0(mai_mai_n246_), .A1(mai_mai_n245_), .B0(mai_mai_n243_), .Y(mai_mai_n247_));
  AN4        m0219(.A(mai_mai_n247_), .B(mai_mai_n241_), .C(mai_mai_n234_), .D(mai_mai_n228_), .Y(mai_mai_n248_));
  OR2        m0220(.A(h), .B(g), .Y(mai_mai_n249_));
  NO2        m0221(.A(mai_mai_n249_), .B(mai_mai_n102_), .Y(mai_mai_n250_));
  NA2        m0222(.A(mai_mai_n250_), .B(mai_mai_n131_), .Y(mai_mai_n251_));
  NAi41      m0223(.An(e), .B(n), .C(d), .D(b), .Y(mai_mai_n252_));
  NO2        m0224(.A(mai_mai_n252_), .B(mai_mai_n217_), .Y(mai_mai_n253_));
  NA2        m0225(.A(mai_mai_n161_), .B(mai_mai_n108_), .Y(mai_mai_n254_));
  NAi21      m0226(.An(mai_mai_n254_), .B(mai_mai_n253_), .Y(mai_mai_n255_));
  NO2        m0227(.A(n), .B(a), .Y(mai_mai_n256_));
  NAi31      m0228(.An(mai_mai_n244_), .B(mai_mai_n256_), .C(mai_mai_n103_), .Y(mai_mai_n257_));
  AN2        m0229(.A(mai_mai_n257_), .B(mai_mai_n255_), .Y(mai_mai_n258_));
  NAi21      m0230(.An(h), .B(i), .Y(mai_mai_n259_));
  NA2        m0231(.A(mai_mai_n181_), .B(k), .Y(mai_mai_n260_));
  NO2        m0232(.A(mai_mai_n260_), .B(mai_mai_n259_), .Y(mai_mai_n261_));
  NA2        m0233(.A(mai_mai_n261_), .B(mai_mai_n194_), .Y(mai_mai_n262_));
  NA3        m0234(.A(mai_mai_n262_), .B(mai_mai_n258_), .C(mai_mai_n251_), .Y(mai_mai_n263_));
  NOi21      m0235(.An(g), .B(e), .Y(mai_mai_n264_));
  NO2        m0236(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n265_));
  NA2        m0237(.A(mai_mai_n265_), .B(mai_mai_n264_), .Y(mai_mai_n266_));
  NOi32      m0238(.An(l), .Bn(j), .C(i), .Y(mai_mai_n267_));
  AOI210     m0239(.A0(mai_mai_n73_), .A1(mai_mai_n86_), .B0(mai_mai_n267_), .Y(mai_mai_n268_));
  NO2        m0240(.A(mai_mai_n259_), .B(mai_mai_n44_), .Y(mai_mai_n269_));
  NAi21      m0241(.An(f), .B(g), .Y(mai_mai_n270_));
  NO2        m0242(.A(mai_mai_n270_), .B(mai_mai_n62_), .Y(mai_mai_n271_));
  NO2        m0243(.A(mai_mai_n66_), .B(mai_mai_n117_), .Y(mai_mai_n272_));
  AOI220     m0244(.A0(mai_mai_n272_), .A1(mai_mai_n271_), .B0(mai_mai_n269_), .B1(mai_mai_n64_), .Y(mai_mai_n273_));
  OAI210     m0245(.A0(mai_mai_n268_), .A1(mai_mai_n266_), .B0(mai_mai_n273_), .Y(mai_mai_n274_));
  NO3        m0246(.A(mai_mai_n134_), .B(mai_mai_n49_), .C(mai_mai_n45_), .Y(mai_mai_n275_));
  NOi41      m0247(.An(mai_mai_n248_), .B(mai_mai_n274_), .C(mai_mai_n263_), .D(mai_mai_n224_), .Y(mai_mai_n276_));
  NO4        m0248(.A(mai_mai_n205_), .B(mai_mai_n48_), .C(mai_mai_n43_), .D(mai_mai_n39_), .Y(mai_mai_n277_));
  NO2        m0249(.A(mai_mai_n277_), .B(mai_mai_n111_), .Y(mai_mai_n278_));
  NA3        m0250(.A(mai_mai_n59_), .B(c), .C(b), .Y(mai_mai_n279_));
  NAi21      m0251(.An(h), .B(g), .Y(mai_mai_n280_));
  OR4        m0252(.A(mai_mai_n280_), .B(mai_mai_n279_), .C(mai_mai_n227_), .D(e), .Y(mai_mai_n281_));
  NO2        m0253(.A(mai_mai_n254_), .B(mai_mai_n270_), .Y(mai_mai_n282_));
  NAi31      m0254(.An(g), .B(k), .C(h), .Y(mai_mai_n283_));
  NO3        m0255(.A(mai_mai_n133_), .B(mai_mai_n283_), .C(l), .Y(mai_mai_n284_));
  NAi31      m0256(.An(e), .B(d), .C(a), .Y(mai_mai_n285_));
  NA2        m0257(.A(mai_mai_n284_), .B(mai_mai_n131_), .Y(mai_mai_n286_));
  NA2        m0258(.A(mai_mai_n286_), .B(mai_mai_n281_), .Y(mai_mai_n287_));
  NA4        m0259(.A(mai_mai_n161_), .B(mai_mai_n79_), .C(mai_mai_n75_), .D(mai_mai_n117_), .Y(mai_mai_n288_));
  NA3        m0260(.A(mai_mai_n161_), .B(mai_mai_n160_), .C(mai_mai_n83_), .Y(mai_mai_n289_));
  NO2        m0261(.A(mai_mai_n289_), .B(mai_mai_n196_), .Y(mai_mai_n290_));
  NOi21      m0262(.An(mai_mai_n288_), .B(mai_mai_n290_), .Y(mai_mai_n291_));
  NA3        m0263(.A(e), .B(c), .C(b), .Y(mai_mai_n292_));
  NAi32      m0264(.An(k), .Bn(i), .C(j), .Y(mai_mai_n293_));
  NAi21      m0265(.An(l), .B(k), .Y(mai_mai_n294_));
  NO2        m0266(.A(mai_mai_n294_), .B(mai_mai_n49_), .Y(mai_mai_n295_));
  NOi21      m0267(.An(l), .B(j), .Y(mai_mai_n296_));
  NA2        m0268(.A(mai_mai_n164_), .B(mai_mai_n296_), .Y(mai_mai_n297_));
  NAi32      m0269(.An(j), .Bn(h), .C(i), .Y(mai_mai_n298_));
  NAi21      m0270(.An(m), .B(l), .Y(mai_mai_n299_));
  NO3        m0271(.A(mai_mai_n299_), .B(mai_mai_n298_), .C(mai_mai_n83_), .Y(mai_mai_n300_));
  NA2        m0272(.A(h), .B(g), .Y(mai_mai_n301_));
  NA2        m0273(.A(mai_mai_n168_), .B(mai_mai_n45_), .Y(mai_mai_n302_));
  NO2        m0274(.A(mai_mai_n302_), .B(mai_mai_n301_), .Y(mai_mai_n303_));
  OAI210     m0275(.A0(mai_mai_n303_), .A1(mai_mai_n300_), .B0(mai_mai_n165_), .Y(mai_mai_n304_));
  NA2        m0276(.A(mai_mai_n304_), .B(mai_mai_n291_), .Y(mai_mai_n305_));
  NO2        m0277(.A(mai_mai_n146_), .B(d), .Y(mai_mai_n306_));
  NA2        m0278(.A(mai_mai_n306_), .B(mai_mai_n53_), .Y(mai_mai_n307_));
  NO2        m0279(.A(mai_mai_n105_), .B(mai_mai_n102_), .Y(mai_mai_n308_));
  NAi32      m0280(.An(n), .Bn(m), .C(l), .Y(mai_mai_n309_));
  NO2        m0281(.A(mai_mai_n309_), .B(mai_mai_n298_), .Y(mai_mai_n310_));
  NA2        m0282(.A(mai_mai_n310_), .B(mai_mai_n185_), .Y(mai_mai_n311_));
  NAi31      m0283(.An(k), .B(l), .C(j), .Y(mai_mai_n312_));
  OAI210     m0284(.A0(mai_mai_n294_), .A1(j), .B0(mai_mai_n312_), .Y(mai_mai_n313_));
  NOi21      m0285(.An(mai_mai_n313_), .B(mai_mai_n120_), .Y(mai_mai_n314_));
  NA2        m0286(.A(mai_mai_n311_), .B(mai_mai_n307_), .Y(mai_mai_n315_));
  NO4        m0287(.A(mai_mai_n315_), .B(mai_mai_n305_), .C(mai_mai_n287_), .D(mai_mai_n278_), .Y(mai_mai_n316_));
  NA2        m0288(.A(mai_mai_n261_), .B(mai_mai_n195_), .Y(mai_mai_n317_));
  NAi21      m0289(.An(m), .B(k), .Y(mai_mai_n318_));
  NO2        m0290(.A(mai_mai_n230_), .B(mai_mai_n318_), .Y(mai_mai_n319_));
  NAi41      m0291(.An(d), .B(n), .C(c), .D(b), .Y(mai_mai_n320_));
  NO2        m0292(.A(mai_mai_n320_), .B(mai_mai_n152_), .Y(mai_mai_n321_));
  NA2        m0293(.A(mai_mai_n321_), .B(mai_mai_n319_), .Y(mai_mai_n322_));
  NAi31      m0294(.An(i), .B(l), .C(h), .Y(mai_mai_n323_));
  NO4        m0295(.A(mai_mai_n323_), .B(mai_mai_n152_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n324_));
  NA2        m0296(.A(e), .B(c), .Y(mai_mai_n325_));
  NO3        m0297(.A(mai_mai_n325_), .B(n), .C(d), .Y(mai_mai_n326_));
  NOi21      m0298(.An(f), .B(h), .Y(mai_mai_n327_));
  NA2        m0299(.A(mai_mai_n327_), .B(mai_mai_n118_), .Y(mai_mai_n328_));
  NO2        m0300(.A(mai_mai_n328_), .B(mai_mai_n218_), .Y(mai_mai_n329_));
  NAi31      m0301(.An(d), .B(e), .C(b), .Y(mai_mai_n330_));
  NO2        m0302(.A(mai_mai_n133_), .B(mai_mai_n330_), .Y(mai_mai_n331_));
  NA2        m0303(.A(mai_mai_n331_), .B(mai_mai_n329_), .Y(mai_mai_n332_));
  NAi41      m0304(.An(mai_mai_n324_), .B(mai_mai_n332_), .C(mai_mai_n322_), .D(mai_mai_n317_), .Y(mai_mai_n333_));
  NO4        m0305(.A(mai_mai_n320_), .B(mai_mai_n78_), .C(mai_mai_n69_), .D(mai_mai_n218_), .Y(mai_mai_n334_));
  NA2        m0306(.A(mai_mai_n256_), .B(mai_mai_n103_), .Y(mai_mai_n335_));
  OR2        m0307(.A(mai_mai_n335_), .B(mai_mai_n207_), .Y(mai_mai_n336_));
  NOi31      m0308(.An(l), .B(n), .C(m), .Y(mai_mai_n337_));
  NA2        m0309(.A(mai_mai_n337_), .B(mai_mai_n219_), .Y(mai_mai_n338_));
  NO2        m0310(.A(mai_mai_n338_), .B(mai_mai_n196_), .Y(mai_mai_n339_));
  NAi32      m0311(.An(mai_mai_n339_), .Bn(mai_mai_n334_), .C(mai_mai_n336_), .Y(mai_mai_n340_));
  NAi32      m0312(.An(m), .Bn(j), .C(k), .Y(mai_mai_n341_));
  NAi41      m0313(.An(c), .B(n), .C(d), .D(b), .Y(mai_mai_n342_));
  OAI210     m0314(.A0(mai_mai_n215_), .A1(mai_mai_n341_), .B0(mai_mai_n342_), .Y(mai_mai_n343_));
  NOi31      m0315(.An(j), .B(m), .C(k), .Y(mai_mai_n344_));
  NO2        m0316(.A(mai_mai_n126_), .B(mai_mai_n344_), .Y(mai_mai_n345_));
  AN3        m0317(.A(h), .B(g), .C(f), .Y(mai_mai_n346_));
  NAi31      m0318(.An(mai_mai_n345_), .B(mai_mai_n346_), .C(mai_mai_n343_), .Y(mai_mai_n347_));
  NOi32      m0319(.An(m), .Bn(j), .C(l), .Y(mai_mai_n348_));
  NO2        m0320(.A(mai_mai_n348_), .B(mai_mai_n96_), .Y(mai_mai_n349_));
  NAi32      m0321(.An(mai_mai_n349_), .Bn(mai_mai_n204_), .C(mai_mai_n306_), .Y(mai_mai_n350_));
  NO2        m0322(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n351_));
  NO2        m0323(.A(mai_mai_n221_), .B(g), .Y(mai_mai_n352_));
  NO2        m0324(.A(mai_mai_n157_), .B(mai_mai_n83_), .Y(mai_mai_n353_));
  AOI220     m0325(.A0(mai_mai_n353_), .A1(mai_mai_n352_), .B0(mai_mai_n253_), .B1(mai_mai_n351_), .Y(mai_mai_n354_));
  NA2        m0326(.A(mai_mai_n238_), .B(mai_mai_n78_), .Y(mai_mai_n355_));
  NA3        m0327(.A(mai_mai_n355_), .B(mai_mai_n346_), .C(mai_mai_n216_), .Y(mai_mai_n356_));
  NA4        m0328(.A(mai_mai_n356_), .B(mai_mai_n354_), .C(mai_mai_n350_), .D(mai_mai_n347_), .Y(mai_mai_n357_));
  NA3        m0329(.A(h), .B(g), .C(f), .Y(mai_mai_n358_));
  NO2        m0330(.A(mai_mai_n358_), .B(mai_mai_n74_), .Y(mai_mai_n359_));
  NA2        m0331(.A(mai_mai_n342_), .B(mai_mai_n215_), .Y(mai_mai_n360_));
  NA2        m0332(.A(mai_mai_n164_), .B(e), .Y(mai_mai_n361_));
  NO2        m0333(.A(mai_mai_n361_), .B(mai_mai_n41_), .Y(mai_mai_n362_));
  NA2        m0334(.A(mai_mai_n360_), .B(mai_mai_n359_), .Y(mai_mai_n363_));
  NOi32      m0335(.An(j), .Bn(g), .C(i), .Y(mai_mai_n364_));
  NA3        m0336(.A(mai_mai_n364_), .B(mai_mai_n294_), .C(mai_mai_n113_), .Y(mai_mai_n365_));
  AO210      m0337(.A0(mai_mai_n111_), .A1(mai_mai_n32_), .B0(mai_mai_n365_), .Y(mai_mai_n366_));
  NOi32      m0338(.An(e), .Bn(b), .C(a), .Y(mai_mai_n367_));
  AN2        m0339(.A(l), .B(j), .Y(mai_mai_n368_));
  NO2        m0340(.A(mai_mai_n318_), .B(mai_mai_n368_), .Y(mai_mai_n369_));
  NO3        m0341(.A(mai_mai_n320_), .B(mai_mai_n69_), .C(mai_mai_n218_), .Y(mai_mai_n370_));
  NA3        m0342(.A(mai_mai_n212_), .B(mai_mai_n210_), .C(mai_mai_n35_), .Y(mai_mai_n371_));
  AOI220     m0343(.A0(mai_mai_n371_), .A1(mai_mai_n367_), .B0(mai_mai_n370_), .B1(mai_mai_n369_), .Y(mai_mai_n372_));
  NA2        m0344(.A(mai_mai_n211_), .B(k), .Y(mai_mai_n373_));
  NA3        m0345(.A(m), .B(mai_mai_n112_), .C(mai_mai_n217_), .Y(mai_mai_n374_));
  NA4        m0346(.A(mai_mai_n206_), .B(mai_mai_n86_), .C(g), .D(mai_mai_n217_), .Y(mai_mai_n375_));
  NAi41      m0347(.An(d), .B(e), .C(c), .D(a), .Y(mai_mai_n376_));
  NA2        m0348(.A(mai_mai_n51_), .B(mai_mai_n113_), .Y(mai_mai_n377_));
  NA3        m0349(.A(mai_mai_n372_), .B(mai_mai_n366_), .C(mai_mai_n363_), .Y(mai_mai_n378_));
  NO4        m0350(.A(mai_mai_n378_), .B(mai_mai_n357_), .C(mai_mai_n340_), .D(mai_mai_n333_), .Y(mai_mai_n379_));
  NA4        m0351(.A(mai_mai_n379_), .B(mai_mai_n316_), .C(mai_mai_n276_), .D(mai_mai_n202_), .Y(mai10));
  NA3        m0352(.A(m), .B(k), .C(i), .Y(mai_mai_n381_));
  NO3        m0353(.A(mai_mai_n381_), .B(j), .C(mai_mai_n218_), .Y(mai_mai_n382_));
  NOi21      m0354(.An(e), .B(f), .Y(mai_mai_n383_));
  NO4        m0355(.A(mai_mai_n153_), .B(mai_mai_n383_), .C(n), .D(mai_mai_n110_), .Y(mai_mai_n384_));
  NAi31      m0356(.An(b), .B(f), .C(c), .Y(mai_mai_n385_));
  INV        m0357(.A(mai_mai_n385_), .Y(mai_mai_n386_));
  NOi32      m0358(.An(k), .Bn(h), .C(j), .Y(mai_mai_n387_));
  NA2        m0359(.A(mai_mai_n387_), .B(mai_mai_n225_), .Y(mai_mai_n388_));
  NA2        m0360(.A(mai_mai_n162_), .B(mai_mai_n388_), .Y(mai_mai_n389_));
  AOI220     m0361(.A0(mai_mai_n389_), .A1(mai_mai_n386_), .B0(mai_mai_n384_), .B1(mai_mai_n382_), .Y(mai_mai_n390_));
  AN2        m0362(.A(j), .B(h), .Y(mai_mai_n391_));
  NO3        m0363(.A(n), .B(m), .C(k), .Y(mai_mai_n392_));
  NA2        m0364(.A(mai_mai_n392_), .B(mai_mai_n391_), .Y(mai_mai_n393_));
  NO3        m0365(.A(mai_mai_n393_), .B(mai_mai_n153_), .C(mai_mai_n217_), .Y(mai_mai_n394_));
  OR2        m0366(.A(m), .B(k), .Y(mai_mai_n395_));
  NO2        m0367(.A(mai_mai_n175_), .B(mai_mai_n395_), .Y(mai_mai_n396_));
  NA4        m0368(.A(n), .B(f), .C(c), .D(mai_mai_n116_), .Y(mai_mai_n397_));
  NOi21      m0369(.An(mai_mai_n396_), .B(mai_mai_n397_), .Y(mai_mai_n398_));
  NOi32      m0370(.An(d), .Bn(a), .C(c), .Y(mai_mai_n399_));
  NA2        m0371(.A(mai_mai_n399_), .B(mai_mai_n183_), .Y(mai_mai_n400_));
  NAi21      m0372(.An(i), .B(g), .Y(mai_mai_n401_));
  NAi31      m0373(.An(k), .B(m), .C(j), .Y(mai_mai_n402_));
  NO3        m0374(.A(mai_mai_n402_), .B(mai_mai_n401_), .C(n), .Y(mai_mai_n403_));
  NOi21      m0375(.An(mai_mai_n403_), .B(mai_mai_n400_), .Y(mai_mai_n404_));
  NO3        m0376(.A(mai_mai_n404_), .B(mai_mai_n398_), .C(mai_mai_n394_), .Y(mai_mai_n405_));
  NO2        m0377(.A(mai_mai_n397_), .B(mai_mai_n299_), .Y(mai_mai_n406_));
  NOi32      m0378(.An(f), .Bn(d), .C(c), .Y(mai_mai_n407_));
  AOI220     m0379(.A0(mai_mai_n407_), .A1(mai_mai_n310_), .B0(mai_mai_n406_), .B1(mai_mai_n219_), .Y(mai_mai_n408_));
  NA3        m0380(.A(mai_mai_n408_), .B(mai_mai_n405_), .C(mai_mai_n390_), .Y(mai_mai_n409_));
  NO2        m0381(.A(mai_mai_n59_), .B(mai_mai_n116_), .Y(mai_mai_n410_));
  NA2        m0382(.A(mai_mai_n256_), .B(mai_mai_n410_), .Y(mai_mai_n411_));
  INV        m0383(.A(e), .Y(mai_mai_n412_));
  NA2        m0384(.A(mai_mai_n46_), .B(e), .Y(mai_mai_n413_));
  OAI220     m0385(.A0(mai_mai_n413_), .A1(mai_mai_n203_), .B0(mai_mai_n207_), .B1(mai_mai_n412_), .Y(mai_mai_n414_));
  AN2        m0386(.A(g), .B(e), .Y(mai_mai_n415_));
  NO2        m0387(.A(mai_mai_n88_), .B(mai_mai_n412_), .Y(mai_mai_n416_));
  NO2        m0388(.A(mai_mai_n99_), .B(mai_mai_n412_), .Y(mai_mai_n417_));
  NO3        m0389(.A(mai_mai_n417_), .B(mai_mai_n416_), .C(mai_mai_n414_), .Y(mai_mai_n418_));
  NOi32      m0390(.An(h), .Bn(e), .C(g), .Y(mai_mai_n419_));
  NA3        m0391(.A(mai_mai_n419_), .B(mai_mai_n296_), .C(m), .Y(mai_mai_n420_));
  NOi21      m0392(.An(g), .B(h), .Y(mai_mai_n421_));
  AN3        m0393(.A(m), .B(l), .C(i), .Y(mai_mai_n422_));
  NA3        m0394(.A(mai_mai_n422_), .B(mai_mai_n421_), .C(e), .Y(mai_mai_n423_));
  AN3        m0395(.A(h), .B(g), .C(e), .Y(mai_mai_n424_));
  NA2        m0396(.A(mai_mai_n424_), .B(mai_mai_n96_), .Y(mai_mai_n425_));
  AN3        m0397(.A(mai_mai_n425_), .B(mai_mai_n423_), .C(mai_mai_n420_), .Y(mai_mai_n426_));
  AOI210     m0398(.A0(mai_mai_n426_), .A1(mai_mai_n418_), .B0(mai_mai_n411_), .Y(mai_mai_n427_));
  NA3        m0399(.A(mai_mai_n399_), .B(mai_mai_n183_), .C(mai_mai_n83_), .Y(mai_mai_n428_));
  NAi31      m0400(.An(b), .B(c), .C(a), .Y(mai_mai_n429_));
  NO2        m0401(.A(mai_mai_n429_), .B(n), .Y(mai_mai_n430_));
  NA2        m0402(.A(mai_mai_n51_), .B(m), .Y(mai_mai_n431_));
  NO2        m0403(.A(mai_mai_n431_), .B(mai_mai_n149_), .Y(mai_mai_n432_));
  NA2        m0404(.A(mai_mai_n432_), .B(mai_mai_n430_), .Y(mai_mai_n433_));
  INV        m0405(.A(mai_mai_n433_), .Y(mai_mai_n434_));
  NO3        m0406(.A(mai_mai_n434_), .B(mai_mai_n427_), .C(mai_mai_n409_), .Y(mai_mai_n435_));
  NA2        m0407(.A(i), .B(g), .Y(mai_mai_n436_));
  NO3        m0408(.A(mai_mai_n285_), .B(mai_mai_n436_), .C(c), .Y(mai_mai_n437_));
  NOi21      m0409(.An(a), .B(n), .Y(mai_mai_n438_));
  NOi21      m0410(.An(d), .B(c), .Y(mai_mai_n439_));
  NA2        m0411(.A(mai_mai_n439_), .B(mai_mai_n438_), .Y(mai_mai_n440_));
  NA3        m0412(.A(i), .B(g), .C(f), .Y(mai_mai_n441_));
  OR2        m0413(.A(mai_mai_n441_), .B(mai_mai_n68_), .Y(mai_mai_n442_));
  NA3        m0414(.A(mai_mai_n422_), .B(mai_mai_n421_), .C(mai_mai_n183_), .Y(mai_mai_n443_));
  AOI210     m0415(.A0(mai_mai_n443_), .A1(mai_mai_n442_), .B0(mai_mai_n440_), .Y(mai_mai_n444_));
  AOI210     m0416(.A0(mai_mai_n437_), .A1(mai_mai_n295_), .B0(mai_mai_n444_), .Y(mai_mai_n445_));
  OR2        m0417(.A(n), .B(m), .Y(mai_mai_n446_));
  NO2        m0418(.A(mai_mai_n446_), .B(mai_mai_n154_), .Y(mai_mai_n447_));
  NO2        m0419(.A(mai_mai_n184_), .B(mai_mai_n149_), .Y(mai_mai_n448_));
  OAI210     m0420(.A0(mai_mai_n447_), .A1(mai_mai_n177_), .B0(mai_mai_n448_), .Y(mai_mai_n449_));
  INV        m0421(.A(mai_mai_n377_), .Y(mai_mai_n450_));
  NA3        m0422(.A(mai_mai_n450_), .B(mai_mai_n367_), .C(d), .Y(mai_mai_n451_));
  NO2        m0423(.A(mai_mai_n429_), .B(mai_mai_n49_), .Y(mai_mai_n452_));
  NO3        m0424(.A(mai_mai_n63_), .B(mai_mai_n112_), .C(e), .Y(mai_mai_n453_));
  NAi21      m0425(.An(k), .B(j), .Y(mai_mai_n454_));
  NA2        m0426(.A(mai_mai_n259_), .B(mai_mai_n454_), .Y(mai_mai_n455_));
  NA3        m0427(.A(mai_mai_n455_), .B(mai_mai_n453_), .C(mai_mai_n452_), .Y(mai_mai_n456_));
  NAi21      m0428(.An(e), .B(d), .Y(mai_mai_n457_));
  INV        m0429(.A(mai_mai_n457_), .Y(mai_mai_n458_));
  NO2        m0430(.A(mai_mai_n260_), .B(mai_mai_n217_), .Y(mai_mai_n459_));
  NA3        m0431(.A(mai_mai_n459_), .B(mai_mai_n458_), .C(mai_mai_n231_), .Y(mai_mai_n460_));
  NA4        m0432(.A(mai_mai_n460_), .B(mai_mai_n456_), .C(mai_mai_n451_), .D(mai_mai_n449_), .Y(mai_mai_n461_));
  NO2        m0433(.A(mai_mai_n338_), .B(mai_mai_n217_), .Y(mai_mai_n462_));
  NA2        m0434(.A(mai_mai_n462_), .B(mai_mai_n458_), .Y(mai_mai_n463_));
  NOi31      m0435(.An(n), .B(m), .C(k), .Y(mai_mai_n464_));
  AOI220     m0436(.A0(mai_mai_n464_), .A1(mai_mai_n391_), .B0(mai_mai_n225_), .B1(mai_mai_n50_), .Y(mai_mai_n465_));
  NAi31      m0437(.An(g), .B(f), .C(c), .Y(mai_mai_n466_));
  OR3        m0438(.A(mai_mai_n466_), .B(mai_mai_n465_), .C(e), .Y(mai_mai_n467_));
  NA3        m0439(.A(mai_mai_n467_), .B(mai_mai_n463_), .C(mai_mai_n311_), .Y(mai_mai_n468_));
  NOi41      m0440(.An(mai_mai_n445_), .B(mai_mai_n468_), .C(mai_mai_n461_), .D(mai_mai_n274_), .Y(mai_mai_n469_));
  NOi32      m0441(.An(c), .Bn(a), .C(b), .Y(mai_mai_n470_));
  NA2        m0442(.A(mai_mai_n470_), .B(mai_mai_n113_), .Y(mai_mai_n471_));
  INV        m0443(.A(mai_mai_n283_), .Y(mai_mai_n472_));
  AN2        m0444(.A(e), .B(d), .Y(mai_mai_n473_));
  NA2        m0445(.A(mai_mai_n473_), .B(mai_mai_n472_), .Y(mai_mai_n474_));
  INV        m0446(.A(mai_mai_n149_), .Y(mai_mai_n475_));
  NO2        m0447(.A(mai_mai_n132_), .B(mai_mai_n41_), .Y(mai_mai_n476_));
  NO2        m0448(.A(mai_mai_n63_), .B(e), .Y(mai_mai_n477_));
  NOi31      m0449(.An(j), .B(k), .C(i), .Y(mai_mai_n478_));
  NOi21      m0450(.An(mai_mai_n167_), .B(mai_mai_n478_), .Y(mai_mai_n479_));
  NA4        m0451(.A(mai_mai_n323_), .B(mai_mai_n479_), .C(mai_mai_n268_), .D(mai_mai_n119_), .Y(mai_mai_n480_));
  AOI220     m0452(.A0(mai_mai_n480_), .A1(mai_mai_n477_), .B0(mai_mai_n476_), .B1(mai_mai_n475_), .Y(mai_mai_n481_));
  AOI210     m0453(.A0(mai_mai_n481_), .A1(mai_mai_n474_), .B0(mai_mai_n471_), .Y(mai_mai_n482_));
  NO2        m0454(.A(mai_mai_n213_), .B(mai_mai_n208_), .Y(mai_mai_n483_));
  NOi21      m0455(.An(a), .B(b), .Y(mai_mai_n484_));
  NA3        m0456(.A(e), .B(d), .C(c), .Y(mai_mai_n485_));
  NAi21      m0457(.An(mai_mai_n485_), .B(mai_mai_n484_), .Y(mai_mai_n486_));
  NO2        m0458(.A(mai_mai_n428_), .B(mai_mai_n207_), .Y(mai_mai_n487_));
  NOi21      m0459(.An(mai_mai_n486_), .B(mai_mai_n487_), .Y(mai_mai_n488_));
  AOI210     m0460(.A0(mai_mai_n277_), .A1(mai_mai_n483_), .B0(mai_mai_n488_), .Y(mai_mai_n489_));
  NO4        m0461(.A(mai_mai_n190_), .B(mai_mai_n102_), .C(mai_mai_n56_), .D(b), .Y(mai_mai_n490_));
  NA2        m0462(.A(mai_mai_n386_), .B(mai_mai_n155_), .Y(mai_mai_n491_));
  OR2        m0463(.A(k), .B(j), .Y(mai_mai_n492_));
  NA2        m0464(.A(l), .B(k), .Y(mai_mai_n493_));
  NA3        m0465(.A(mai_mai_n493_), .B(mai_mai_n492_), .C(mai_mai_n225_), .Y(mai_mai_n494_));
  AOI210     m0466(.A0(mai_mai_n238_), .A1(mai_mai_n341_), .B0(mai_mai_n83_), .Y(mai_mai_n495_));
  NOi21      m0467(.An(mai_mai_n494_), .B(mai_mai_n495_), .Y(mai_mai_n496_));
  OR3        m0468(.A(mai_mai_n496_), .B(mai_mai_n145_), .C(mai_mai_n136_), .Y(mai_mai_n497_));
  NA3        m0469(.A(mai_mai_n288_), .B(mai_mai_n129_), .C(mai_mai_n127_), .Y(mai_mai_n498_));
  NA2        m0470(.A(mai_mai_n399_), .B(mai_mai_n113_), .Y(mai_mai_n499_));
  NO4        m0471(.A(mai_mai_n499_), .B(mai_mai_n93_), .C(mai_mai_n112_), .D(e), .Y(mai_mai_n500_));
  NO3        m0472(.A(mai_mai_n428_), .B(mai_mai_n90_), .C(mai_mai_n132_), .Y(mai_mai_n501_));
  NO4        m0473(.A(mai_mai_n501_), .B(mai_mai_n500_), .C(mai_mai_n498_), .D(mai_mai_n324_), .Y(mai_mai_n502_));
  NA3        m0474(.A(mai_mai_n502_), .B(mai_mai_n497_), .C(mai_mai_n491_), .Y(mai_mai_n503_));
  NO4        m0475(.A(mai_mai_n503_), .B(mai_mai_n490_), .C(mai_mai_n489_), .D(mai_mai_n482_), .Y(mai_mai_n504_));
  NA2        m0476(.A(mai_mai_n67_), .B(mai_mai_n64_), .Y(mai_mai_n505_));
  NOi21      m0477(.An(d), .B(e), .Y(mai_mai_n506_));
  NO2        m0478(.A(mai_mai_n190_), .B(mai_mai_n56_), .Y(mai_mai_n507_));
  NAi31      m0479(.An(j), .B(l), .C(i), .Y(mai_mai_n508_));
  OAI210     m0480(.A0(mai_mai_n508_), .A1(mai_mai_n133_), .B0(mai_mai_n102_), .Y(mai_mai_n509_));
  NA3        m0481(.A(mai_mai_n509_), .B(mai_mai_n507_), .C(mai_mai_n506_), .Y(mai_mai_n510_));
  NO3        m0482(.A(mai_mai_n400_), .B(mai_mai_n349_), .C(mai_mai_n204_), .Y(mai_mai_n511_));
  NO2        m0483(.A(mai_mai_n400_), .B(mai_mai_n377_), .Y(mai_mai_n512_));
  NO4        m0484(.A(mai_mai_n512_), .B(mai_mai_n511_), .C(mai_mai_n186_), .D(mai_mai_n308_), .Y(mai_mai_n513_));
  NA4        m0485(.A(mai_mai_n513_), .B(mai_mai_n510_), .C(mai_mai_n505_), .D(mai_mai_n248_), .Y(mai_mai_n514_));
  OAI210     m0486(.A0(mai_mai_n128_), .A1(mai_mai_n126_), .B0(n), .Y(mai_mai_n515_));
  NO2        m0487(.A(mai_mai_n515_), .B(mai_mai_n132_), .Y(mai_mai_n516_));
  BUFFER     m0488(.A(mai_mai_n250_), .Y(mai_mai_n517_));
  OA210      m0489(.A0(mai_mai_n517_), .A1(mai_mai_n516_), .B0(mai_mai_n195_), .Y(mai_mai_n518_));
  XO2        m0490(.A(i), .B(h), .Y(mai_mai_n519_));
  NA3        m0491(.A(mai_mai_n519_), .B(mai_mai_n161_), .C(n), .Y(mai_mai_n520_));
  NAi41      m0492(.An(mai_mai_n300_), .B(mai_mai_n520_), .C(mai_mai_n465_), .D(mai_mai_n388_), .Y(mai_mai_n521_));
  NOi32      m0493(.An(mai_mai_n521_), .Bn(mai_mai_n477_), .C(mai_mai_n279_), .Y(mai_mai_n522_));
  NAi31      m0494(.An(c), .B(f), .C(d), .Y(mai_mai_n523_));
  AOI210     m0495(.A0(mai_mai_n289_), .A1(mai_mai_n198_), .B0(mai_mai_n523_), .Y(mai_mai_n524_));
  NOi21      m0496(.An(mai_mai_n81_), .B(mai_mai_n524_), .Y(mai_mai_n525_));
  NA3        m0497(.A(mai_mai_n384_), .B(mai_mai_n96_), .C(mai_mai_n95_), .Y(mai_mai_n526_));
  NA2        m0498(.A(mai_mai_n232_), .B(mai_mai_n108_), .Y(mai_mai_n527_));
  AOI210     m0499(.A0(mai_mai_n527_), .A1(mai_mai_n182_), .B0(mai_mai_n523_), .Y(mai_mai_n528_));
  AOI210     m0500(.A0(mai_mai_n365_), .A1(mai_mai_n35_), .B0(mai_mai_n486_), .Y(mai_mai_n529_));
  NOi31      m0501(.An(mai_mai_n526_), .B(mai_mai_n529_), .C(mai_mai_n528_), .Y(mai_mai_n530_));
  NA3        m0502(.A(mai_mai_n37_), .B(mai_mai_n36_), .C(f), .Y(mai_mai_n531_));
  NO2        m0503(.A(mai_mai_n531_), .B(mai_mai_n440_), .Y(mai_mai_n532_));
  INV        m0504(.A(mai_mai_n532_), .Y(mai_mai_n533_));
  NA3        m0505(.A(mai_mai_n533_), .B(mai_mai_n530_), .C(mai_mai_n525_), .Y(mai_mai_n534_));
  NO4        m0506(.A(mai_mai_n534_), .B(mai_mai_n522_), .C(mai_mai_n518_), .D(mai_mai_n514_), .Y(mai_mai_n535_));
  NA4        m0507(.A(mai_mai_n535_), .B(mai_mai_n504_), .C(mai_mai_n469_), .D(mai_mai_n435_), .Y(mai11));
  NO2        m0508(.A(mai_mai_n70_), .B(f), .Y(mai_mai_n537_));
  NA2        m0509(.A(j), .B(g), .Y(mai_mai_n538_));
  NAi31      m0510(.An(i), .B(m), .C(l), .Y(mai_mai_n539_));
  NA3        m0511(.A(m), .B(k), .C(j), .Y(mai_mai_n540_));
  OAI220     m0512(.A0(mai_mai_n540_), .A1(mai_mai_n132_), .B0(mai_mai_n539_), .B1(mai_mai_n538_), .Y(mai_mai_n541_));
  NA2        m0513(.A(mai_mai_n541_), .B(mai_mai_n537_), .Y(mai_mai_n542_));
  NOi32      m0514(.An(e), .Bn(b), .C(f), .Y(mai_mai_n543_));
  NA2        m0515(.A(mai_mai_n267_), .B(mai_mai_n113_), .Y(mai_mai_n544_));
  NA2        m0516(.A(mai_mai_n46_), .B(j), .Y(mai_mai_n545_));
  NO2        m0517(.A(mai_mai_n545_), .B(mai_mai_n302_), .Y(mai_mai_n546_));
  NAi31      m0518(.An(d), .B(e), .C(a), .Y(mai_mai_n547_));
  NO2        m0519(.A(mai_mai_n547_), .B(n), .Y(mai_mai_n548_));
  AOI220     m0520(.A0(mai_mai_n548_), .A1(mai_mai_n100_), .B0(mai_mai_n546_), .B1(mai_mai_n543_), .Y(mai_mai_n549_));
  NAi41      m0521(.An(f), .B(e), .C(c), .D(a), .Y(mai_mai_n550_));
  AN2        m0522(.A(mai_mai_n550_), .B(mai_mai_n376_), .Y(mai_mai_n551_));
  AOI210     m0523(.A0(mai_mai_n551_), .A1(mai_mai_n400_), .B0(mai_mai_n280_), .Y(mai_mai_n552_));
  NA2        m0524(.A(j), .B(i), .Y(mai_mai_n553_));
  NAi31      m0525(.An(n), .B(m), .C(k), .Y(mai_mai_n554_));
  NO3        m0526(.A(mai_mai_n554_), .B(mai_mai_n553_), .C(mai_mai_n112_), .Y(mai_mai_n555_));
  NO4        m0527(.A(n), .B(d), .C(mai_mai_n116_), .D(a), .Y(mai_mai_n556_));
  OR2        m0528(.A(n), .B(c), .Y(mai_mai_n557_));
  NO2        m0529(.A(mai_mai_n557_), .B(mai_mai_n151_), .Y(mai_mai_n558_));
  NO2        m0530(.A(mai_mai_n558_), .B(mai_mai_n556_), .Y(mai_mai_n559_));
  NOi32      m0531(.An(g), .Bn(f), .C(i), .Y(mai_mai_n560_));
  AOI220     m0532(.A0(mai_mai_n560_), .A1(mai_mai_n98_), .B0(mai_mai_n541_), .B1(f), .Y(mai_mai_n561_));
  NO2        m0533(.A(mai_mai_n283_), .B(mai_mai_n49_), .Y(mai_mai_n562_));
  NO2        m0534(.A(mai_mai_n561_), .B(mai_mai_n559_), .Y(mai_mai_n563_));
  AOI210     m0535(.A0(mai_mai_n555_), .A1(mai_mai_n552_), .B0(mai_mai_n563_), .Y(mai_mai_n564_));
  NA2        m0536(.A(mai_mai_n141_), .B(mai_mai_n34_), .Y(mai_mai_n565_));
  OAI220     m0537(.A0(mai_mai_n565_), .A1(m), .B0(mai_mai_n545_), .B1(mai_mai_n238_), .Y(mai_mai_n566_));
  NOi41      m0538(.An(d), .B(n), .C(e), .D(c), .Y(mai_mai_n567_));
  NAi32      m0539(.An(e), .Bn(b), .C(c), .Y(mai_mai_n568_));
  OR2        m0540(.A(mai_mai_n568_), .B(mai_mai_n83_), .Y(mai_mai_n569_));
  AN2        m0541(.A(mai_mai_n342_), .B(mai_mai_n320_), .Y(mai_mai_n570_));
  NA2        m0542(.A(mai_mai_n570_), .B(mai_mai_n569_), .Y(mai_mai_n571_));
  OA210      m0543(.A0(mai_mai_n571_), .A1(mai_mai_n567_), .B0(mai_mai_n566_), .Y(mai_mai_n572_));
  OAI220     m0544(.A0(mai_mai_n402_), .A1(mai_mai_n401_), .B0(mai_mai_n539_), .B1(mai_mai_n538_), .Y(mai_mai_n573_));
  NO3        m0545(.A(mai_mai_n61_), .B(mai_mai_n49_), .C(mai_mai_n218_), .Y(mai_mai_n574_));
  NO2        m0546(.A(mai_mai_n235_), .B(mai_mai_n110_), .Y(mai_mai_n575_));
  OAI210     m0547(.A0(mai_mai_n574_), .A1(mai_mai_n403_), .B0(mai_mai_n575_), .Y(mai_mai_n576_));
  INV        m0548(.A(mai_mai_n576_), .Y(mai_mai_n577_));
  NO2        m0549(.A(mai_mai_n285_), .B(n), .Y(mai_mai_n578_));
  NO2        m0550(.A(mai_mai_n430_), .B(mai_mai_n578_), .Y(mai_mai_n579_));
  NA2        m0551(.A(mai_mai_n573_), .B(f), .Y(mai_mai_n580_));
  NAi32      m0552(.An(d), .Bn(a), .C(b), .Y(mai_mai_n581_));
  NO2        m0553(.A(mai_mai_n581_), .B(mai_mai_n49_), .Y(mai_mai_n582_));
  NA2        m0554(.A(h), .B(f), .Y(mai_mai_n583_));
  NO2        m0555(.A(mai_mai_n583_), .B(mai_mai_n93_), .Y(mai_mai_n584_));
  NO3        m0556(.A(mai_mai_n178_), .B(mai_mai_n175_), .C(g), .Y(mai_mai_n585_));
  AOI220     m0557(.A0(mai_mai_n585_), .A1(mai_mai_n58_), .B0(mai_mai_n584_), .B1(mai_mai_n582_), .Y(mai_mai_n586_));
  OAI210     m0558(.A0(mai_mai_n580_), .A1(mai_mai_n579_), .B0(mai_mai_n586_), .Y(mai_mai_n587_));
  AN3        m0559(.A(j), .B(h), .C(g), .Y(mai_mai_n588_));
  NO2        m0560(.A(mai_mai_n148_), .B(c), .Y(mai_mai_n589_));
  NA3        m0561(.A(mai_mai_n589_), .B(mai_mai_n588_), .C(mai_mai_n464_), .Y(mai_mai_n590_));
  NA3        m0562(.A(f), .B(d), .C(b), .Y(mai_mai_n591_));
  NO4        m0563(.A(mai_mai_n591_), .B(mai_mai_n178_), .C(mai_mai_n175_), .D(g), .Y(mai_mai_n592_));
  NAi21      m0564(.An(mai_mai_n592_), .B(mai_mai_n590_), .Y(mai_mai_n593_));
  NO4        m0565(.A(mai_mai_n593_), .B(mai_mai_n587_), .C(mai_mai_n577_), .D(mai_mai_n572_), .Y(mai_mai_n594_));
  AN4        m0566(.A(mai_mai_n594_), .B(mai_mai_n564_), .C(mai_mai_n549_), .D(mai_mai_n542_), .Y(mai_mai_n595_));
  INV        m0567(.A(k), .Y(mai_mai_n596_));
  NA3        m0568(.A(l), .B(mai_mai_n596_), .C(i), .Y(mai_mai_n597_));
  INV        m0569(.A(mai_mai_n597_), .Y(mai_mai_n598_));
  NA4        m0570(.A(mai_mai_n399_), .B(mai_mai_n421_), .C(mai_mai_n183_), .D(mai_mai_n113_), .Y(mai_mai_n599_));
  NAi32      m0571(.An(h), .Bn(f), .C(g), .Y(mai_mai_n600_));
  NAi41      m0572(.An(n), .B(e), .C(c), .D(a), .Y(mai_mai_n601_));
  OAI210     m0573(.A0(mai_mai_n547_), .A1(n), .B0(mai_mai_n601_), .Y(mai_mai_n602_));
  NA2        m0574(.A(mai_mai_n602_), .B(m), .Y(mai_mai_n603_));
  NAi31      m0575(.An(h), .B(g), .C(f), .Y(mai_mai_n604_));
  OR2        m0576(.A(mai_mai_n603_), .B(mai_mai_n600_), .Y(mai_mai_n605_));
  NA2        m0577(.A(mai_mai_n605_), .B(mai_mai_n599_), .Y(mai_mai_n606_));
  NAi31      m0578(.An(f), .B(h), .C(g), .Y(mai_mai_n607_));
  NO4        m0579(.A(mai_mai_n312_), .B(mai_mai_n607_), .C(mai_mai_n70_), .D(mai_mai_n72_), .Y(mai_mai_n608_));
  NOi32      m0580(.An(b), .Bn(a), .C(c), .Y(mai_mai_n609_));
  NOi32      m0581(.An(d), .Bn(a), .C(e), .Y(mai_mai_n610_));
  NO2        m0582(.A(n), .B(c), .Y(mai_mai_n611_));
  NAi32      m0583(.An(n), .Bn(f), .C(m), .Y(mai_mai_n612_));
  NOi32      m0584(.An(e), .Bn(a), .C(d), .Y(mai_mai_n613_));
  AOI210     m0585(.A0(mai_mai_n29_), .A1(d), .B0(mai_mai_n613_), .Y(mai_mai_n614_));
  AOI210     m0586(.A0(mai_mai_n614_), .A1(mai_mai_n217_), .B0(mai_mai_n565_), .Y(mai_mai_n615_));
  AOI210     m0587(.A0(mai_mai_n615_), .A1(mai_mai_n1552_), .B0(mai_mai_n608_), .Y(mai_mai_n616_));
  OAI210     m0588(.A0(mai_mai_n255_), .A1(mai_mai_n86_), .B0(mai_mai_n616_), .Y(mai_mai_n617_));
  AOI210     m0589(.A0(mai_mai_n606_), .A1(mai_mai_n598_), .B0(mai_mai_n617_), .Y(mai_mai_n618_));
  NO3        m0590(.A(mai_mai_n318_), .B(mai_mai_n60_), .C(n), .Y(mai_mai_n619_));
  NA3        m0591(.A(mai_mai_n523_), .B(mai_mai_n173_), .C(mai_mai_n172_), .Y(mai_mai_n620_));
  NA2        m0592(.A(mai_mai_n466_), .B(mai_mai_n235_), .Y(mai_mai_n621_));
  OR2        m0593(.A(mai_mai_n621_), .B(mai_mai_n620_), .Y(mai_mai_n622_));
  NA2        m0594(.A(mai_mai_n73_), .B(mai_mai_n113_), .Y(mai_mai_n623_));
  NO2        m0595(.A(mai_mai_n623_), .B(mai_mai_n45_), .Y(mai_mai_n624_));
  AOI220     m0596(.A0(mai_mai_n624_), .A1(mai_mai_n552_), .B0(mai_mai_n622_), .B1(mai_mai_n619_), .Y(mai_mai_n625_));
  NO2        m0597(.A(mai_mai_n625_), .B(mai_mai_n86_), .Y(mai_mai_n626_));
  NA3        m0598(.A(mai_mai_n567_), .B(mai_mai_n344_), .C(mai_mai_n46_), .Y(mai_mai_n627_));
  NOi32      m0599(.An(e), .Bn(c), .C(f), .Y(mai_mai_n628_));
  NOi21      m0600(.An(f), .B(g), .Y(mai_mai_n629_));
  NO2        m0601(.A(mai_mai_n629_), .B(mai_mai_n215_), .Y(mai_mai_n630_));
  AOI220     m0602(.A0(mai_mai_n630_), .A1(mai_mai_n396_), .B0(mai_mai_n628_), .B1(mai_mai_n177_), .Y(mai_mai_n631_));
  NA3        m0603(.A(mai_mai_n631_), .B(mai_mai_n627_), .C(mai_mai_n180_), .Y(mai_mai_n632_));
  AOI210     m0604(.A0(mai_mai_n551_), .A1(mai_mai_n400_), .B0(mai_mai_n301_), .Y(mai_mai_n633_));
  NA2        m0605(.A(mai_mai_n633_), .B(mai_mai_n272_), .Y(mai_mai_n634_));
  NOi21      m0606(.An(j), .B(l), .Y(mai_mai_n635_));
  NAi21      m0607(.An(k), .B(h), .Y(mai_mai_n636_));
  NO2        m0608(.A(mai_mai_n636_), .B(mai_mai_n270_), .Y(mai_mai_n637_));
  NA2        m0609(.A(mai_mai_n637_), .B(mai_mai_n635_), .Y(mai_mai_n638_));
  OR2        m0610(.A(mai_mai_n638_), .B(mai_mai_n603_), .Y(mai_mai_n639_));
  NOi31      m0611(.An(m), .B(n), .C(k), .Y(mai_mai_n640_));
  NO2        m0612(.A(mai_mai_n285_), .B(mai_mai_n49_), .Y(mai_mai_n641_));
  NO2        m0613(.A(mai_mai_n312_), .B(mai_mai_n607_), .Y(mai_mai_n642_));
  NO2        m0614(.A(mai_mai_n547_), .B(mai_mai_n49_), .Y(mai_mai_n643_));
  AOI220     m0615(.A0(mai_mai_n643_), .A1(mai_mai_n642_), .B0(mai_mai_n641_), .B1(mai_mai_n584_), .Y(mai_mai_n644_));
  NA3        m0616(.A(mai_mai_n644_), .B(mai_mai_n639_), .C(mai_mai_n634_), .Y(mai_mai_n645_));
  NA2        m0617(.A(mai_mai_n108_), .B(mai_mai_n36_), .Y(mai_mai_n646_));
  NO2        m0618(.A(k), .B(mai_mai_n218_), .Y(mai_mai_n647_));
  INV        m0619(.A(mai_mai_n367_), .Y(mai_mai_n648_));
  NO2        m0620(.A(mai_mai_n648_), .B(n), .Y(mai_mai_n649_));
  NAi31      m0621(.An(mai_mai_n646_), .B(mai_mai_n649_), .C(mai_mai_n647_), .Y(mai_mai_n650_));
  NO2        m0622(.A(mai_mai_n545_), .B(mai_mai_n178_), .Y(mai_mai_n651_));
  NA3        m0623(.A(mai_mai_n568_), .B(mai_mai_n279_), .C(mai_mai_n146_), .Y(mai_mai_n652_));
  NA2        m0624(.A(mai_mai_n519_), .B(mai_mai_n161_), .Y(mai_mai_n653_));
  NO3        m0625(.A(mai_mai_n397_), .B(mai_mai_n653_), .C(mai_mai_n86_), .Y(mai_mai_n654_));
  AOI210     m0626(.A0(mai_mai_n652_), .A1(mai_mai_n651_), .B0(mai_mai_n654_), .Y(mai_mai_n655_));
  AN3        m0627(.A(f), .B(d), .C(b), .Y(mai_mai_n656_));
  OAI210     m0628(.A0(mai_mai_n656_), .A1(mai_mai_n131_), .B0(n), .Y(mai_mai_n657_));
  NA3        m0629(.A(mai_mai_n519_), .B(mai_mai_n161_), .C(mai_mai_n218_), .Y(mai_mai_n658_));
  AOI210     m0630(.A0(mai_mai_n657_), .A1(mai_mai_n237_), .B0(mai_mai_n658_), .Y(mai_mai_n659_));
  NAi31      m0631(.An(m), .B(n), .C(k), .Y(mai_mai_n660_));
  OR2        m0632(.A(mai_mai_n136_), .B(mai_mai_n60_), .Y(mai_mai_n661_));
  OAI210     m0633(.A0(mai_mai_n661_), .A1(mai_mai_n660_), .B0(mai_mai_n257_), .Y(mai_mai_n662_));
  OAI210     m0634(.A0(mai_mai_n662_), .A1(mai_mai_n659_), .B0(j), .Y(mai_mai_n663_));
  NA3        m0635(.A(mai_mai_n663_), .B(mai_mai_n655_), .C(mai_mai_n650_), .Y(mai_mai_n664_));
  NO4        m0636(.A(mai_mai_n664_), .B(mai_mai_n645_), .C(mai_mai_n632_), .D(mai_mai_n626_), .Y(mai_mai_n665_));
  NA2        m0637(.A(mai_mai_n384_), .B(mai_mai_n164_), .Y(mai_mai_n666_));
  NAi31      m0638(.An(g), .B(h), .C(f), .Y(mai_mai_n667_));
  OA210      m0639(.A0(mai_mai_n547_), .A1(n), .B0(mai_mai_n601_), .Y(mai_mai_n668_));
  NO2        m0640(.A(mai_mai_n668_), .B(mai_mai_n89_), .Y(mai_mai_n669_));
  INV        m0641(.A(mai_mai_n669_), .Y(mai_mai_n670_));
  AOI210     m0642(.A0(mai_mai_n670_), .A1(mai_mai_n666_), .B0(mai_mai_n540_), .Y(mai_mai_n671_));
  NO3        m0643(.A(g), .B(mai_mai_n217_), .C(mai_mai_n56_), .Y(mai_mai_n672_));
  NAi21      m0644(.An(h), .B(j), .Y(mai_mai_n673_));
  NO2        m0645(.A(mai_mai_n527_), .B(mai_mai_n86_), .Y(mai_mai_n674_));
  OAI210     m0646(.A0(mai_mai_n674_), .A1(mai_mai_n396_), .B0(mai_mai_n672_), .Y(mai_mai_n675_));
  OR2        m0647(.A(mai_mai_n70_), .B(mai_mai_n72_), .Y(mai_mai_n676_));
  AN2        m0648(.A(h), .B(f), .Y(mai_mai_n677_));
  NA2        m0649(.A(mai_mai_n677_), .B(mai_mai_n37_), .Y(mai_mai_n678_));
  NA2        m0650(.A(mai_mai_n98_), .B(mai_mai_n46_), .Y(mai_mai_n679_));
  OAI220     m0651(.A0(mai_mai_n679_), .A1(mai_mai_n335_), .B0(mai_mai_n678_), .B1(mai_mai_n471_), .Y(mai_mai_n680_));
  AOI210     m0652(.A0(mai_mai_n581_), .A1(mai_mai_n429_), .B0(mai_mai_n49_), .Y(mai_mai_n681_));
  OAI220     m0653(.A0(mai_mai_n604_), .A1(mai_mai_n597_), .B0(mai_mai_n328_), .B1(mai_mai_n538_), .Y(mai_mai_n682_));
  AOI210     m0654(.A0(mai_mai_n682_), .A1(mai_mai_n681_), .B0(mai_mai_n680_), .Y(mai_mai_n683_));
  NA2        m0655(.A(mai_mai_n683_), .B(mai_mai_n675_), .Y(mai_mai_n684_));
  NO2        m0656(.A(mai_mai_n259_), .B(f), .Y(mai_mai_n685_));
  NO2        m0657(.A(mai_mai_n629_), .B(mai_mai_n60_), .Y(mai_mai_n686_));
  NO3        m0658(.A(mai_mai_n686_), .B(mai_mai_n685_), .C(mai_mai_n34_), .Y(mai_mai_n687_));
  NA2        m0659(.A(mai_mai_n331_), .B(mai_mai_n141_), .Y(mai_mai_n688_));
  NA2        m0660(.A(mai_mai_n133_), .B(mai_mai_n49_), .Y(mai_mai_n689_));
  AOI220     m0661(.A0(mai_mai_n689_), .A1(mai_mai_n543_), .B0(mai_mai_n367_), .B1(mai_mai_n113_), .Y(mai_mai_n690_));
  OA220      m0662(.A0(mai_mai_n690_), .A1(mai_mai_n565_), .B0(mai_mai_n365_), .B1(mai_mai_n111_), .Y(mai_mai_n691_));
  OAI210     m0663(.A0(mai_mai_n688_), .A1(mai_mai_n687_), .B0(mai_mai_n691_), .Y(mai_mai_n692_));
  NO3        m0664(.A(mai_mai_n407_), .B(mai_mai_n195_), .C(mai_mai_n194_), .Y(mai_mai_n693_));
  NA2        m0665(.A(mai_mai_n693_), .B(mai_mai_n235_), .Y(mai_mai_n694_));
  NA3        m0666(.A(mai_mai_n694_), .B(mai_mai_n261_), .C(j), .Y(mai_mai_n695_));
  NO3        m0667(.A(mai_mai_n466_), .B(mai_mai_n175_), .C(i), .Y(mai_mai_n696_));
  NA2        m0668(.A(mai_mai_n470_), .B(mai_mai_n83_), .Y(mai_mai_n697_));
  NO4        m0669(.A(mai_mai_n540_), .B(mai_mai_n697_), .C(mai_mai_n132_), .D(mai_mai_n217_), .Y(mai_mai_n698_));
  INV        m0670(.A(mai_mai_n698_), .Y(mai_mai_n699_));
  NA4        m0671(.A(mai_mai_n699_), .B(mai_mai_n695_), .C(mai_mai_n526_), .D(mai_mai_n405_), .Y(mai_mai_n700_));
  NO4        m0672(.A(mai_mai_n700_), .B(mai_mai_n692_), .C(mai_mai_n684_), .D(mai_mai_n671_), .Y(mai_mai_n701_));
  NA4        m0673(.A(mai_mai_n701_), .B(mai_mai_n665_), .C(mai_mai_n618_), .D(mai_mai_n595_), .Y(mai08));
  NO2        m0674(.A(k), .B(h), .Y(mai_mai_n703_));
  AO210      m0675(.A0(mai_mai_n259_), .A1(mai_mai_n454_), .B0(mai_mai_n703_), .Y(mai_mai_n704_));
  NO2        m0676(.A(mai_mai_n704_), .B(mai_mai_n299_), .Y(mai_mai_n705_));
  NA2        m0677(.A(mai_mai_n628_), .B(mai_mai_n83_), .Y(mai_mai_n706_));
  NA2        m0678(.A(mai_mai_n706_), .B(mai_mai_n466_), .Y(mai_mai_n707_));
  AOI210     m0679(.A0(mai_mai_n707_), .A1(mai_mai_n705_), .B0(mai_mai_n501_), .Y(mai_mai_n708_));
  NA2        m0680(.A(mai_mai_n83_), .B(mai_mai_n110_), .Y(mai_mai_n709_));
  NO2        m0681(.A(mai_mai_n709_), .B(mai_mai_n57_), .Y(mai_mai_n710_));
  NO4        m0682(.A(mai_mai_n381_), .B(mai_mai_n112_), .C(j), .D(mai_mai_n218_), .Y(mai_mai_n711_));
  NA2        m0683(.A(mai_mai_n591_), .B(mai_mai_n237_), .Y(mai_mai_n712_));
  AOI220     m0684(.A0(mai_mai_n712_), .A1(mai_mai_n352_), .B0(mai_mai_n711_), .B1(mai_mai_n710_), .Y(mai_mai_n713_));
  AOI210     m0685(.A0(mai_mai_n591_), .A1(mai_mai_n157_), .B0(mai_mai_n83_), .Y(mai_mai_n714_));
  NA4        m0686(.A(mai_mai_n220_), .B(mai_mai_n141_), .C(mai_mai_n45_), .D(h), .Y(mai_mai_n715_));
  AN2        m0687(.A(l), .B(k), .Y(mai_mai_n716_));
  NA3        m0688(.A(mai_mai_n713_), .B(mai_mai_n708_), .C(mai_mai_n354_), .Y(mai_mai_n717_));
  AN2        m0689(.A(mai_mai_n548_), .B(mai_mai_n94_), .Y(mai_mai_n718_));
  NO4        m0690(.A(mai_mai_n175_), .B(mai_mai_n395_), .C(mai_mai_n112_), .D(g), .Y(mai_mai_n719_));
  AOI210     m0691(.A0(mai_mai_n719_), .A1(mai_mai_n712_), .B0(mai_mai_n532_), .Y(mai_mai_n720_));
  NO2        m0692(.A(mai_mai_n38_), .B(mai_mai_n217_), .Y(mai_mai_n721_));
  AOI220     m0693(.A0(mai_mai_n630_), .A1(mai_mai_n351_), .B0(mai_mai_n721_), .B1(mai_mai_n578_), .Y(mai_mai_n722_));
  NAi31      m0694(.An(mai_mai_n718_), .B(mai_mai_n722_), .C(mai_mai_n720_), .Y(mai_mai_n723_));
  OAI210     m0695(.A0(mai_mai_n568_), .A1(mai_mai_n47_), .B0(mai_mai_n661_), .Y(mai_mai_n724_));
  NO2        m0696(.A(mai_mai_n493_), .B(mai_mai_n133_), .Y(mai_mai_n725_));
  NA2        m0697(.A(mai_mai_n725_), .B(mai_mai_n724_), .Y(mai_mai_n726_));
  NO3        m0698(.A(mai_mai_n318_), .B(mai_mai_n132_), .C(mai_mai_n41_), .Y(mai_mai_n727_));
  BUFFER     m0699(.A(mai_mai_n727_), .Y(mai_mai_n728_));
  NA2        m0700(.A(mai_mai_n704_), .B(mai_mai_n137_), .Y(mai_mai_n729_));
  AOI220     m0701(.A0(mai_mai_n729_), .A1(mai_mai_n406_), .B0(mai_mai_n728_), .B1(mai_mai_n75_), .Y(mai_mai_n730_));
  NA2        m0702(.A(mai_mai_n726_), .B(mai_mai_n730_), .Y(mai_mai_n731_));
  NA2        m0703(.A(mai_mai_n367_), .B(mai_mai_n43_), .Y(mai_mai_n732_));
  NA3        m0704(.A(mai_mai_n694_), .B(mai_mai_n337_), .C(mai_mai_n387_), .Y(mai_mai_n733_));
  NA2        m0705(.A(mai_mai_n716_), .B(mai_mai_n225_), .Y(mai_mai_n734_));
  NO2        m0706(.A(mai_mai_n734_), .B(mai_mai_n330_), .Y(mai_mai_n735_));
  AOI210     m0707(.A0(mai_mai_n735_), .A1(mai_mai_n685_), .B0(mai_mai_n500_), .Y(mai_mai_n736_));
  NA3        m0708(.A(m), .B(l), .C(k), .Y(mai_mai_n737_));
  NO2        m0709(.A(mai_mai_n550_), .B(mai_mai_n280_), .Y(mai_mai_n738_));
  NOi21      m0710(.An(mai_mai_n738_), .B(mai_mai_n544_), .Y(mai_mai_n739_));
  NA4        m0711(.A(mai_mai_n113_), .B(l), .C(k), .D(mai_mai_n86_), .Y(mai_mai_n740_));
  NA3        m0712(.A(mai_mai_n121_), .B(mai_mai_n415_), .C(i), .Y(mai_mai_n741_));
  NO2        m0713(.A(mai_mai_n741_), .B(mai_mai_n740_), .Y(mai_mai_n742_));
  NO2        m0714(.A(mai_mai_n742_), .B(mai_mai_n739_), .Y(mai_mai_n743_));
  NA4        m0715(.A(mai_mai_n743_), .B(mai_mai_n736_), .C(mai_mai_n733_), .D(mai_mai_n732_), .Y(mai_mai_n744_));
  NO4        m0716(.A(mai_mai_n744_), .B(mai_mai_n731_), .C(mai_mai_n723_), .D(mai_mai_n717_), .Y(mai_mai_n745_));
  NA2        m0717(.A(mai_mai_n630_), .B(mai_mai_n396_), .Y(mai_mai_n746_));
  NOi31      m0718(.An(g), .B(h), .C(f), .Y(mai_mai_n747_));
  NA2        m0719(.A(mai_mai_n643_), .B(mai_mai_n747_), .Y(mai_mai_n748_));
  OR2        m0720(.A(mai_mai_n748_), .B(mai_mai_n553_), .Y(mai_mai_n749_));
  NO3        m0721(.A(mai_mai_n400_), .B(mai_mai_n538_), .C(h), .Y(mai_mai_n750_));
  AOI210     m0722(.A0(mai_mai_n750_), .A1(mai_mai_n113_), .B0(mai_mai_n512_), .Y(mai_mai_n751_));
  NA4        m0723(.A(mai_mai_n751_), .B(mai_mai_n749_), .C(mai_mai_n746_), .D(mai_mai_n258_), .Y(mai_mai_n752_));
  NA2        m0724(.A(mai_mai_n716_), .B(mai_mai_n72_), .Y(mai_mai_n753_));
  NO4        m0725(.A(mai_mai_n693_), .B(mai_mai_n175_), .C(n), .D(i), .Y(mai_mai_n754_));
  NOi21      m0726(.An(h), .B(j), .Y(mai_mai_n755_));
  NA2        m0727(.A(mai_mai_n755_), .B(f), .Y(mai_mai_n756_));
  NO2        m0728(.A(mai_mai_n754_), .B(mai_mai_n696_), .Y(mai_mai_n757_));
  NO2        m0729(.A(mai_mai_n757_), .B(mai_mai_n753_), .Y(mai_mai_n758_));
  AOI210     m0730(.A0(mai_mai_n752_), .A1(l), .B0(mai_mai_n758_), .Y(mai_mai_n759_));
  NO2        m0731(.A(j), .B(i), .Y(mai_mai_n760_));
  NA3        m0732(.A(mai_mai_n760_), .B(mai_mai_n79_), .C(l), .Y(mai_mai_n761_));
  NA2        m0733(.A(mai_mai_n760_), .B(mai_mai_n33_), .Y(mai_mai_n762_));
  OR2        m0734(.A(mai_mai_n761_), .B(mai_mai_n603_), .Y(mai_mai_n763_));
  NO3        m0735(.A(mai_mai_n153_), .B(mai_mai_n49_), .C(mai_mai_n110_), .Y(mai_mai_n764_));
  NO3        m0736(.A(mai_mai_n557_), .B(mai_mai_n151_), .C(mai_mai_n72_), .Y(mai_mai_n765_));
  NO3        m0737(.A(mai_mai_n493_), .B(mai_mai_n441_), .C(j), .Y(mai_mai_n766_));
  OAI210     m0738(.A0(mai_mai_n765_), .A1(mai_mai_n764_), .B0(mai_mai_n766_), .Y(mai_mai_n767_));
  OAI210     m0739(.A0(mai_mai_n748_), .A1(mai_mai_n61_), .B0(mai_mai_n767_), .Y(mai_mai_n768_));
  NA2        m0740(.A(k), .B(j), .Y(mai_mai_n769_));
  NO3        m0741(.A(mai_mai_n299_), .B(mai_mai_n769_), .C(mai_mai_n40_), .Y(mai_mai_n770_));
  AOI210     m0742(.A0(mai_mai_n543_), .A1(n), .B0(mai_mai_n567_), .Y(mai_mai_n771_));
  NA2        m0743(.A(mai_mai_n771_), .B(mai_mai_n570_), .Y(mai_mai_n772_));
  AN3        m0744(.A(mai_mai_n772_), .B(mai_mai_n770_), .C(mai_mai_n97_), .Y(mai_mai_n773_));
  NO3        m0745(.A(mai_mai_n175_), .B(mai_mai_n395_), .C(mai_mai_n112_), .Y(mai_mai_n774_));
  AOI220     m0746(.A0(mai_mai_n774_), .A1(mai_mai_n253_), .B0(mai_mai_n621_), .B1(mai_mai_n310_), .Y(mai_mai_n775_));
  NAi31      m0747(.An(mai_mai_n614_), .B(mai_mai_n91_), .C(mai_mai_n83_), .Y(mai_mai_n776_));
  NA2        m0748(.A(mai_mai_n776_), .B(mai_mai_n775_), .Y(mai_mai_n777_));
  NO2        m0749(.A(mai_mai_n299_), .B(mai_mai_n137_), .Y(mai_mai_n778_));
  AOI220     m0750(.A0(mai_mai_n778_), .A1(mai_mai_n630_), .B0(mai_mai_n727_), .B1(mai_mai_n714_), .Y(mai_mai_n779_));
  NO2        m0751(.A(mai_mai_n737_), .B(mai_mai_n89_), .Y(mai_mai_n780_));
  NA2        m0752(.A(mai_mai_n780_), .B(mai_mai_n602_), .Y(mai_mai_n781_));
  NO2        m0753(.A(mai_mai_n604_), .B(mai_mai_n117_), .Y(mai_mai_n782_));
  OAI210     m0754(.A0(mai_mai_n782_), .A1(mai_mai_n766_), .B0(mai_mai_n681_), .Y(mai_mai_n783_));
  NA3        m0755(.A(mai_mai_n783_), .B(mai_mai_n781_), .C(mai_mai_n779_), .Y(mai_mai_n784_));
  OR4        m0756(.A(mai_mai_n784_), .B(mai_mai_n777_), .C(mai_mai_n773_), .D(mai_mai_n768_), .Y(mai_mai_n785_));
  NA3        m0757(.A(mai_mai_n771_), .B(mai_mai_n570_), .C(mai_mai_n569_), .Y(mai_mai_n786_));
  NA4        m0758(.A(mai_mai_n786_), .B(mai_mai_n220_), .C(mai_mai_n454_), .D(mai_mai_n34_), .Y(mai_mai_n787_));
  OAI220     m0759(.A0(mai_mai_n715_), .A1(mai_mai_n706_), .B0(mai_mai_n335_), .B1(mai_mai_n38_), .Y(mai_mai_n788_));
  INV        m0760(.A(mai_mai_n788_), .Y(mai_mai_n789_));
  NA3        m0761(.A(mai_mai_n560_), .B(mai_mai_n296_), .C(h), .Y(mai_mai_n790_));
  NOi21      m0762(.An(mai_mai_n681_), .B(mai_mai_n790_), .Y(mai_mai_n791_));
  NO2        m0763(.A(mai_mai_n90_), .B(mai_mai_n47_), .Y(mai_mai_n792_));
  NO2        m0764(.A(mai_mai_n761_), .B(mai_mai_n676_), .Y(mai_mai_n793_));
  AOI210     m0765(.A0(mai_mai_n792_), .A1(mai_mai_n649_), .B0(mai_mai_n793_), .Y(mai_mai_n794_));
  NAi41      m0766(.An(mai_mai_n791_), .B(mai_mai_n794_), .C(mai_mai_n789_), .D(mai_mai_n787_), .Y(mai_mai_n795_));
  OR2        m0767(.A(mai_mai_n780_), .B(mai_mai_n94_), .Y(mai_mai_n796_));
  AOI220     m0768(.A0(mai_mai_n796_), .A1(mai_mai_n243_), .B0(mai_mai_n766_), .B1(mai_mai_n641_), .Y(mai_mai_n797_));
  NO2        m0769(.A(mai_mai_n668_), .B(mai_mai_n72_), .Y(mai_mai_n798_));
  INV        m0770(.A(mai_mai_n339_), .Y(mai_mai_n799_));
  OAI210     m0771(.A0(mai_mai_n737_), .A1(mai_mai_n667_), .B0(mai_mai_n531_), .Y(mai_mai_n800_));
  NA3        m0772(.A(mai_mai_n256_), .B(mai_mai_n59_), .C(b), .Y(mai_mai_n801_));
  AOI220     m0773(.A0(mai_mai_n611_), .A1(mai_mai_n29_), .B0(mai_mai_n470_), .B1(mai_mai_n83_), .Y(mai_mai_n802_));
  NA2        m0774(.A(mai_mai_n802_), .B(mai_mai_n801_), .Y(mai_mai_n803_));
  NO2        m0775(.A(mai_mai_n790_), .B(mai_mai_n499_), .Y(mai_mai_n804_));
  AOI210     m0776(.A0(mai_mai_n803_), .A1(mai_mai_n800_), .B0(mai_mai_n804_), .Y(mai_mai_n805_));
  NA3        m0777(.A(mai_mai_n805_), .B(mai_mai_n799_), .C(mai_mai_n797_), .Y(mai_mai_n806_));
  NOi41      m0778(.An(mai_mai_n763_), .B(mai_mai_n806_), .C(mai_mai_n795_), .D(mai_mai_n785_), .Y(mai_mai_n807_));
  OR3        m0779(.A(mai_mai_n715_), .B(mai_mai_n237_), .C(g), .Y(mai_mai_n808_));
  NO3        m0780(.A(mai_mai_n345_), .B(mai_mai_n301_), .C(mai_mai_n112_), .Y(mai_mai_n809_));
  NA2        m0781(.A(mai_mai_n809_), .B(mai_mai_n772_), .Y(mai_mai_n810_));
  NA2        m0782(.A(mai_mai_n46_), .B(mai_mai_n56_), .Y(mai_mai_n811_));
  NO3        m0783(.A(mai_mai_n811_), .B(mai_mai_n762_), .C(mai_mai_n285_), .Y(mai_mai_n812_));
  NO3        m0784(.A(mai_mai_n538_), .B(mai_mai_n92_), .C(h), .Y(mai_mai_n813_));
  AOI210     m0785(.A0(mai_mai_n813_), .A1(mai_mai_n710_), .B0(mai_mai_n812_), .Y(mai_mai_n814_));
  NA4        m0786(.A(mai_mai_n814_), .B(mai_mai_n810_), .C(mai_mai_n808_), .D(mai_mai_n408_), .Y(mai_mai_n815_));
  OR2        m0787(.A(mai_mai_n667_), .B(mai_mai_n90_), .Y(mai_mai_n816_));
  NOi31      m0788(.An(b), .B(d), .C(a), .Y(mai_mai_n817_));
  NO2        m0789(.A(mai_mai_n817_), .B(mai_mai_n610_), .Y(mai_mai_n818_));
  NO2        m0790(.A(mai_mai_n818_), .B(n), .Y(mai_mai_n819_));
  NOi21      m0791(.An(mai_mai_n802_), .B(mai_mai_n819_), .Y(mai_mai_n820_));
  NO2        m0792(.A(mai_mai_n820_), .B(mai_mai_n816_), .Y(mai_mai_n821_));
  NO2        m0793(.A(mai_mai_n568_), .B(mai_mai_n83_), .Y(mai_mai_n822_));
  NO3        m0794(.A(mai_mai_n629_), .B(mai_mai_n330_), .C(mai_mai_n117_), .Y(mai_mai_n823_));
  NOi21      m0795(.An(mai_mai_n823_), .B(mai_mai_n162_), .Y(mai_mai_n824_));
  AOI210     m0796(.A0(mai_mai_n809_), .A1(mai_mai_n822_), .B0(mai_mai_n824_), .Y(mai_mai_n825_));
  OAI210     m0797(.A0(mai_mai_n715_), .A1(mai_mai_n397_), .B0(mai_mai_n825_), .Y(mai_mai_n826_));
  NO2        m0798(.A(mai_mai_n693_), .B(n), .Y(mai_mai_n827_));
  AOI220     m0799(.A0(mai_mai_n778_), .A1(mai_mai_n672_), .B0(mai_mai_n827_), .B1(mai_mai_n705_), .Y(mai_mai_n828_));
  NO2        m0800(.A(mai_mai_n325_), .B(mai_mai_n242_), .Y(mai_mai_n829_));
  OAI210     m0801(.A0(mai_mai_n94_), .A1(mai_mai_n91_), .B0(mai_mai_n829_), .Y(mai_mai_n830_));
  NA2        m0802(.A(mai_mai_n121_), .B(mai_mai_n83_), .Y(mai_mai_n831_));
  INV        m0803(.A(mai_mai_n830_), .Y(mai_mai_n832_));
  NA2        m0804(.A(mai_mai_n735_), .B(mai_mai_n34_), .Y(mai_mai_n833_));
  NAi21      m0805(.An(mai_mai_n740_), .B(mai_mai_n437_), .Y(mai_mai_n834_));
  NO2        m0806(.A(mai_mai_n280_), .B(i), .Y(mai_mai_n835_));
  NA2        m0807(.A(mai_mai_n719_), .B(mai_mai_n353_), .Y(mai_mai_n836_));
  AN2        m0808(.A(mai_mai_n836_), .B(mai_mai_n834_), .Y(mai_mai_n837_));
  NAi41      m0809(.An(mai_mai_n832_), .B(mai_mai_n837_), .C(mai_mai_n833_), .D(mai_mai_n828_), .Y(mai_mai_n838_));
  NO4        m0810(.A(mai_mai_n838_), .B(mai_mai_n826_), .C(mai_mai_n821_), .D(mai_mai_n815_), .Y(mai_mai_n839_));
  NA4        m0811(.A(mai_mai_n839_), .B(mai_mai_n807_), .C(mai_mai_n759_), .D(mai_mai_n745_), .Y(mai09));
  INV        m0812(.A(mai_mai_n122_), .Y(mai_mai_n841_));
  NA2        m0813(.A(f), .B(e), .Y(mai_mai_n842_));
  NO2        m0814(.A(mai_mai_n230_), .B(mai_mai_n112_), .Y(mai_mai_n843_));
  NA2        m0815(.A(mai_mai_n843_), .B(g), .Y(mai_mai_n844_));
  NA4        m0816(.A(mai_mai_n312_), .B(mai_mai_n479_), .C(mai_mai_n268_), .D(mai_mai_n119_), .Y(mai_mai_n845_));
  AOI210     m0817(.A0(mai_mai_n845_), .A1(g), .B0(mai_mai_n476_), .Y(mai_mai_n846_));
  AOI210     m0818(.A0(mai_mai_n846_), .A1(mai_mai_n844_), .B0(mai_mai_n842_), .Y(mai_mai_n847_));
  NA2        m0819(.A(mai_mai_n447_), .B(e), .Y(mai_mai_n848_));
  NO2        m0820(.A(mai_mai_n848_), .B(mai_mai_n523_), .Y(mai_mai_n849_));
  AOI210     m0821(.A0(mai_mai_n847_), .A1(mai_mai_n841_), .B0(mai_mai_n849_), .Y(mai_mai_n850_));
  NO2        m0822(.A(mai_mai_n207_), .B(mai_mai_n217_), .Y(mai_mai_n851_));
  NA3        m0823(.A(m), .B(l), .C(i), .Y(mai_mai_n852_));
  OAI220     m0824(.A0(mai_mai_n604_), .A1(mai_mai_n852_), .B0(mai_mai_n358_), .B1(mai_mai_n539_), .Y(mai_mai_n853_));
  NA4        m0825(.A(mai_mai_n87_), .B(mai_mai_n86_), .C(g), .D(f), .Y(mai_mai_n854_));
  NAi31      m0826(.An(mai_mai_n853_), .B(mai_mai_n854_), .C(mai_mai_n442_), .Y(mai_mai_n855_));
  OR2        m0827(.A(mai_mai_n855_), .B(mai_mai_n851_), .Y(mai_mai_n856_));
  NA3        m0828(.A(mai_mai_n816_), .B(mai_mai_n580_), .C(mai_mai_n531_), .Y(mai_mai_n857_));
  OA210      m0829(.A0(mai_mai_n857_), .A1(mai_mai_n856_), .B0(mai_mai_n819_), .Y(mai_mai_n858_));
  INV        m0830(.A(mai_mai_n342_), .Y(mai_mai_n859_));
  NO2        m0831(.A(mai_mai_n128_), .B(mai_mai_n126_), .Y(mai_mai_n860_));
  NOi31      m0832(.An(k), .B(m), .C(l), .Y(mai_mai_n861_));
  NO2        m0833(.A(mai_mai_n344_), .B(mai_mai_n861_), .Y(mai_mai_n862_));
  AOI210     m0834(.A0(mai_mai_n862_), .A1(mai_mai_n860_), .B0(mai_mai_n607_), .Y(mai_mai_n863_));
  NA2        m0835(.A(mai_mai_n801_), .B(mai_mai_n335_), .Y(mai_mai_n864_));
  NA2        m0836(.A(mai_mai_n346_), .B(mai_mai_n348_), .Y(mai_mai_n865_));
  OAI210     m0837(.A0(mai_mai_n207_), .A1(mai_mai_n217_), .B0(mai_mai_n865_), .Y(mai_mai_n866_));
  AOI220     m0838(.A0(mai_mai_n866_), .A1(mai_mai_n864_), .B0(mai_mai_n863_), .B1(mai_mai_n859_), .Y(mai_mai_n867_));
  NA2        m0839(.A(mai_mai_n169_), .B(mai_mai_n114_), .Y(mai_mai_n868_));
  NA3        m0840(.A(mai_mai_n868_), .B(mai_mai_n704_), .C(mai_mai_n137_), .Y(mai_mai_n869_));
  NA3        m0841(.A(mai_mai_n869_), .B(mai_mai_n192_), .C(mai_mai_n31_), .Y(mai_mai_n870_));
  NA4        m0842(.A(mai_mai_n870_), .B(mai_mai_n867_), .C(mai_mai_n631_), .D(mai_mai_n81_), .Y(mai_mai_n871_));
  NO2        m0843(.A(mai_mai_n600_), .B(mai_mai_n508_), .Y(mai_mai_n872_));
  NA2        m0844(.A(mai_mai_n872_), .B(mai_mai_n192_), .Y(mai_mai_n873_));
  NOi21      m0845(.An(f), .B(d), .Y(mai_mai_n874_));
  NA2        m0846(.A(mai_mai_n874_), .B(m), .Y(mai_mai_n875_));
  NO2        m0847(.A(mai_mai_n875_), .B(mai_mai_n52_), .Y(mai_mai_n876_));
  NOi32      m0848(.An(g), .Bn(f), .C(d), .Y(mai_mai_n877_));
  NA4        m0849(.A(mai_mai_n877_), .B(mai_mai_n611_), .C(mai_mai_n29_), .D(m), .Y(mai_mai_n878_));
  NA2        m0850(.A(mai_mai_n876_), .B(mai_mai_n558_), .Y(mai_mai_n879_));
  NA3        m0851(.A(mai_mai_n312_), .B(mai_mai_n268_), .C(mai_mai_n119_), .Y(mai_mai_n880_));
  AN2        m0852(.A(f), .B(d), .Y(mai_mai_n881_));
  NA3        m0853(.A(mai_mai_n484_), .B(mai_mai_n881_), .C(mai_mai_n83_), .Y(mai_mai_n882_));
  NO3        m0854(.A(mai_mai_n882_), .B(mai_mai_n72_), .C(mai_mai_n218_), .Y(mai_mai_n883_));
  NO2        m0855(.A(mai_mai_n293_), .B(mai_mai_n56_), .Y(mai_mai_n884_));
  NA2        m0856(.A(mai_mai_n880_), .B(mai_mai_n883_), .Y(mai_mai_n885_));
  NAi41      m0857(.An(mai_mai_n498_), .B(mai_mai_n885_), .C(mai_mai_n879_), .D(mai_mai_n873_), .Y(mai_mai_n886_));
  NO4        m0858(.A(mai_mai_n629_), .B(mai_mai_n133_), .C(mai_mai_n330_), .D(mai_mai_n154_), .Y(mai_mai_n887_));
  NO2        m0859(.A(mai_mai_n660_), .B(mai_mai_n330_), .Y(mai_mai_n888_));
  AN2        m0860(.A(mai_mai_n888_), .B(mai_mai_n685_), .Y(mai_mai_n889_));
  NO3        m0861(.A(mai_mai_n889_), .B(mai_mai_n887_), .C(mai_mai_n239_), .Y(mai_mai_n890_));
  NA2        m0862(.A(mai_mai_n610_), .B(mai_mai_n83_), .Y(mai_mai_n891_));
  NA3        m0863(.A(mai_mai_n161_), .B(mai_mai_n108_), .C(mai_mai_n107_), .Y(mai_mai_n892_));
  OAI220     m0864(.A0(mai_mai_n882_), .A1(mai_mai_n431_), .B0(mai_mai_n342_), .B1(mai_mai_n892_), .Y(mai_mai_n893_));
  NOi31      m0865(.An(mai_mai_n228_), .B(mai_mai_n893_), .C(mai_mai_n308_), .Y(mai_mai_n894_));
  NA2        m0866(.A(c), .B(mai_mai_n116_), .Y(mai_mai_n895_));
  NO2        m0867(.A(mai_mai_n895_), .B(mai_mai_n412_), .Y(mai_mai_n896_));
  NA3        m0868(.A(mai_mai_n896_), .B(mai_mai_n521_), .C(f), .Y(mai_mai_n897_));
  OR2        m0869(.A(mai_mai_n667_), .B(mai_mai_n554_), .Y(mai_mai_n898_));
  INV        m0870(.A(mai_mai_n898_), .Y(mai_mai_n899_));
  NA2        m0871(.A(mai_mai_n818_), .B(mai_mai_n111_), .Y(mai_mai_n900_));
  NA2        m0872(.A(mai_mai_n900_), .B(mai_mai_n899_), .Y(mai_mai_n901_));
  NA4        m0873(.A(mai_mai_n901_), .B(mai_mai_n897_), .C(mai_mai_n894_), .D(mai_mai_n890_), .Y(mai_mai_n902_));
  NO4        m0874(.A(mai_mai_n902_), .B(mai_mai_n886_), .C(mai_mai_n871_), .D(mai_mai_n858_), .Y(mai_mai_n903_));
  OR2        m0875(.A(mai_mai_n882_), .B(mai_mai_n72_), .Y(mai_mai_n904_));
  NA2        m0876(.A(mai_mai_n843_), .B(g), .Y(mai_mai_n905_));
  AOI210     m0877(.A0(mai_mai_n905_), .A1(mai_mai_n297_), .B0(mai_mai_n904_), .Y(mai_mai_n906_));
  NO2        m0878(.A(mai_mai_n137_), .B(mai_mai_n133_), .Y(mai_mai_n907_));
  NO2        m0879(.A(mai_mai_n235_), .B(mai_mai_n229_), .Y(mai_mai_n908_));
  AOI220     m0880(.A0(mai_mai_n908_), .A1(mai_mai_n232_), .B0(mai_mai_n306_), .B1(mai_mai_n907_), .Y(mai_mai_n909_));
  NO2        m0881(.A(mai_mai_n431_), .B(mai_mai_n842_), .Y(mai_mai_n910_));
  NA2        m0882(.A(e), .B(d), .Y(mai_mai_n911_));
  OAI220     m0883(.A0(mai_mai_n911_), .A1(c), .B0(mai_mai_n325_), .B1(d), .Y(mai_mai_n912_));
  NA3        m0884(.A(mai_mai_n912_), .B(mai_mai_n459_), .C(mai_mai_n519_), .Y(mai_mai_n913_));
  AOI210     m0885(.A0(mai_mai_n527_), .A1(mai_mai_n182_), .B0(mai_mai_n235_), .Y(mai_mai_n914_));
  AOI210     m0886(.A0(mai_mai_n630_), .A1(mai_mai_n351_), .B0(mai_mai_n914_), .Y(mai_mai_n915_));
  NA2        m0887(.A(mai_mai_n293_), .B(mai_mai_n167_), .Y(mai_mai_n916_));
  NA2        m0888(.A(mai_mai_n883_), .B(mai_mai_n916_), .Y(mai_mai_n917_));
  NA3        m0889(.A(mai_mai_n168_), .B(mai_mai_n84_), .C(mai_mai_n34_), .Y(mai_mai_n918_));
  NA4        m0890(.A(mai_mai_n918_), .B(mai_mai_n917_), .C(mai_mai_n915_), .D(mai_mai_n913_), .Y(mai_mai_n919_));
  NO3        m0891(.A(mai_mai_n919_), .B(mai_mai_n1553_), .C(mai_mai_n906_), .Y(mai_mai_n920_));
  NA2        m0892(.A(mai_mai_n859_), .B(mai_mai_n31_), .Y(mai_mai_n921_));
  AO210      m0893(.A0(mai_mai_n921_), .A1(mai_mai_n706_), .B0(mai_mai_n221_), .Y(mai_mai_n922_));
  OAI220     m0894(.A0(mai_mai_n629_), .A1(mai_mai_n60_), .B0(mai_mai_n301_), .B1(j), .Y(mai_mai_n923_));
  AOI220     m0895(.A0(mai_mai_n923_), .A1(mai_mai_n888_), .B0(mai_mai_n619_), .B1(mai_mai_n628_), .Y(mai_mai_n924_));
  OAI210     m0896(.A0(mai_mai_n848_), .A1(mai_mai_n172_), .B0(mai_mai_n924_), .Y(mai_mai_n925_));
  AOI210     m0897(.A0(mai_mai_n118_), .A1(mai_mai_n117_), .B0(mai_mai_n267_), .Y(mai_mai_n926_));
  NO2        m0898(.A(mai_mai_n926_), .B(mai_mai_n878_), .Y(mai_mai_n927_));
  AO210      m0899(.A0(mai_mai_n864_), .A1(mai_mai_n853_), .B0(mai_mai_n927_), .Y(mai_mai_n928_));
  NOi31      m0900(.An(mai_mai_n558_), .B(mai_mai_n875_), .C(mai_mai_n297_), .Y(mai_mai_n929_));
  NO3        m0901(.A(mai_mai_n929_), .B(mai_mai_n928_), .C(mai_mai_n925_), .Y(mai_mai_n930_));
  AO220      m0902(.A0(mai_mai_n459_), .A1(mai_mai_n755_), .B0(mai_mai_n177_), .B1(f), .Y(mai_mai_n931_));
  OAI210     m0903(.A0(mai_mai_n931_), .A1(mai_mai_n462_), .B0(mai_mai_n912_), .Y(mai_mai_n932_));
  NA2        m0904(.A(mai_mai_n857_), .B(mai_mai_n710_), .Y(mai_mai_n933_));
  AN4        m0905(.A(mai_mai_n933_), .B(mai_mai_n932_), .C(mai_mai_n930_), .D(mai_mai_n922_), .Y(mai_mai_n934_));
  NA4        m0906(.A(mai_mai_n934_), .B(mai_mai_n920_), .C(mai_mai_n903_), .D(mai_mai_n850_), .Y(mai12));
  NO2        m0907(.A(mai_mai_n457_), .B(c), .Y(mai_mai_n936_));
  NO4        m0908(.A(mai_mai_n446_), .B(mai_mai_n259_), .C(mai_mai_n596_), .D(mai_mai_n218_), .Y(mai_mai_n937_));
  NA2        m0909(.A(mai_mai_n937_), .B(mai_mai_n936_), .Y(mai_mai_n938_));
  NO2        m0910(.A(mai_mai_n457_), .B(mai_mai_n116_), .Y(mai_mai_n939_));
  NO2        m0911(.A(mai_mai_n860_), .B(mai_mai_n358_), .Y(mai_mai_n940_));
  NO2        m0912(.A(mai_mai_n667_), .B(mai_mai_n381_), .Y(mai_mai_n941_));
  AOI220     m0913(.A0(mai_mai_n941_), .A1(mai_mai_n556_), .B0(mai_mai_n940_), .B1(mai_mai_n939_), .Y(mai_mai_n942_));
  NA3        m0914(.A(mai_mai_n942_), .B(mai_mai_n938_), .C(mai_mai_n445_), .Y(mai_mai_n943_));
  AOI210     m0915(.A0(mai_mai_n238_), .A1(mai_mai_n341_), .B0(mai_mai_n204_), .Y(mai_mai_n944_));
  OR2        m0916(.A(mai_mai_n944_), .B(mai_mai_n937_), .Y(mai_mai_n945_));
  AOI210     m0917(.A0(mai_mai_n338_), .A1(mai_mai_n393_), .B0(mai_mai_n218_), .Y(mai_mai_n946_));
  OAI210     m0918(.A0(mai_mai_n946_), .A1(mai_mai_n945_), .B0(mai_mai_n407_), .Y(mai_mai_n947_));
  NO2        m0919(.A(mai_mai_n646_), .B(mai_mai_n270_), .Y(mai_mai_n948_));
  NO2        m0920(.A(mai_mai_n604_), .B(mai_mai_n852_), .Y(mai_mai_n949_));
  AOI220     m0921(.A0(mai_mai_n949_), .A1(mai_mai_n578_), .B0(mai_mai_n829_), .B1(mai_mai_n948_), .Y(mai_mai_n950_));
  NO2        m0922(.A(mai_mai_n153_), .B(mai_mai_n242_), .Y(mai_mai_n951_));
  NA3        m0923(.A(mai_mai_n951_), .B(mai_mai_n245_), .C(i), .Y(mai_mai_n952_));
  NA3        m0924(.A(mai_mai_n952_), .B(mai_mai_n950_), .C(mai_mai_n947_), .Y(mai_mai_n953_));
  OR2        m0925(.A(mai_mai_n326_), .B(mai_mai_n939_), .Y(mai_mai_n954_));
  NA2        m0926(.A(mai_mai_n954_), .B(mai_mai_n359_), .Y(mai_mai_n955_));
  NO3        m0927(.A(mai_mai_n133_), .B(mai_mai_n154_), .C(mai_mai_n218_), .Y(mai_mai_n956_));
  NA2        m0928(.A(mai_mai_n956_), .B(mai_mai_n543_), .Y(mai_mai_n957_));
  NA4        m0929(.A(mai_mai_n447_), .B(mai_mai_n439_), .C(mai_mai_n183_), .D(g), .Y(mai_mai_n958_));
  NA3        m0930(.A(mai_mai_n958_), .B(mai_mai_n957_), .C(mai_mai_n955_), .Y(mai_mai_n959_));
  NO3        m0931(.A(mai_mai_n670_), .B(mai_mai_n90_), .C(mai_mai_n45_), .Y(mai_mai_n960_));
  NO4        m0932(.A(mai_mai_n960_), .B(mai_mai_n959_), .C(mai_mai_n953_), .D(mai_mai_n943_), .Y(mai_mai_n961_));
  NO2        m0933(.A(mai_mai_n374_), .B(mai_mai_n373_), .Y(mai_mai_n962_));
  INV        m0934(.A(mai_mai_n601_), .Y(mai_mai_n963_));
  NA2        m0935(.A(mai_mai_n568_), .B(mai_mai_n146_), .Y(mai_mai_n964_));
  NOi21      m0936(.An(mai_mai_n34_), .B(mai_mai_n660_), .Y(mai_mai_n965_));
  AOI220     m0937(.A0(mai_mai_n965_), .A1(mai_mai_n964_), .B0(mai_mai_n963_), .B1(mai_mai_n962_), .Y(mai_mai_n966_));
  OAI210     m0938(.A0(mai_mai_n257_), .A1(mai_mai_n45_), .B0(mai_mai_n966_), .Y(mai_mai_n967_));
  NA2        m0939(.A(mai_mai_n437_), .B(mai_mai_n272_), .Y(mai_mai_n968_));
  NO3        m0940(.A(mai_mai_n831_), .B(mai_mai_n88_), .C(mai_mai_n412_), .Y(mai_mai_n969_));
  NAi31      m0941(.An(mai_mai_n969_), .B(mai_mai_n968_), .C(mai_mai_n322_), .Y(mai_mai_n970_));
  NO2        m0942(.A(mai_mai_n49_), .B(mai_mai_n45_), .Y(mai_mai_n971_));
  NO2        m0943(.A(mai_mai_n515_), .B(mai_mai_n301_), .Y(mai_mai_n972_));
  INV        m0944(.A(mai_mai_n972_), .Y(mai_mai_n973_));
  NO2        m0945(.A(mai_mai_n973_), .B(mai_mai_n146_), .Y(mai_mai_n974_));
  NA2        m0946(.A(mai_mai_n640_), .B(mai_mai_n368_), .Y(mai_mai_n975_));
  OAI210     m0947(.A0(mai_mai_n741_), .A1(mai_mai_n975_), .B0(mai_mai_n372_), .Y(mai_mai_n976_));
  NO4        m0948(.A(mai_mai_n976_), .B(mai_mai_n974_), .C(mai_mai_n970_), .D(mai_mai_n967_), .Y(mai_mai_n977_));
  NA2        m0949(.A(mai_mai_n351_), .B(g), .Y(mai_mai_n978_));
  NA2        m0950(.A(mai_mai_n164_), .B(i), .Y(mai_mai_n979_));
  NA2        m0951(.A(mai_mai_n46_), .B(i), .Y(mai_mai_n980_));
  OAI220     m0952(.A0(mai_mai_n980_), .A1(mai_mai_n203_), .B0(mai_mai_n979_), .B1(mai_mai_n90_), .Y(mai_mai_n981_));
  AOI210     m0953(.A0(mai_mai_n422_), .A1(mai_mai_n37_), .B0(mai_mai_n981_), .Y(mai_mai_n982_));
  NO2        m0954(.A(mai_mai_n146_), .B(mai_mai_n83_), .Y(mai_mai_n983_));
  OR2        m0955(.A(mai_mai_n983_), .B(mai_mai_n567_), .Y(mai_mai_n984_));
  NA2        m0956(.A(mai_mai_n568_), .B(mai_mai_n385_), .Y(mai_mai_n985_));
  AOI210     m0957(.A0(mai_mai_n985_), .A1(n), .B0(mai_mai_n984_), .Y(mai_mai_n986_));
  OAI220     m0958(.A0(mai_mai_n986_), .A1(mai_mai_n978_), .B0(mai_mai_n982_), .B1(mai_mai_n335_), .Y(mai_mai_n987_));
  NO2        m0959(.A(mai_mai_n667_), .B(mai_mai_n508_), .Y(mai_mai_n988_));
  NA3        m0960(.A(mai_mai_n346_), .B(mai_mai_n635_), .C(i), .Y(mai_mai_n989_));
  OAI210     m0961(.A0(mai_mai_n441_), .A1(mai_mai_n312_), .B0(mai_mai_n989_), .Y(mai_mai_n990_));
  OAI220     m0962(.A0(mai_mai_n990_), .A1(mai_mai_n988_), .B0(mai_mai_n681_), .B1(mai_mai_n765_), .Y(mai_mai_n991_));
  NA2        m0963(.A(mai_mai_n613_), .B(mai_mai_n113_), .Y(mai_mai_n992_));
  OR3        m0964(.A(mai_mai_n312_), .B(mai_mai_n436_), .C(f), .Y(mai_mai_n993_));
  NA3        m0965(.A(mai_mai_n635_), .B(mai_mai_n79_), .C(i), .Y(mai_mai_n994_));
  OA220      m0966(.A0(mai_mai_n994_), .A1(mai_mai_n992_), .B0(mai_mai_n993_), .B1(mai_mai_n603_), .Y(mai_mai_n995_));
  NA3        m0967(.A(mai_mai_n327_), .B(mai_mai_n118_), .C(g), .Y(mai_mai_n996_));
  AOI210     m0968(.A0(mai_mai_n678_), .A1(mai_mai_n996_), .B0(m), .Y(mai_mai_n997_));
  OAI210     m0969(.A0(mai_mai_n997_), .A1(mai_mai_n940_), .B0(mai_mai_n326_), .Y(mai_mai_n998_));
  NA2        m0970(.A(mai_mai_n697_), .B(mai_mai_n891_), .Y(mai_mai_n999_));
  NA2        m0971(.A(mai_mai_n854_), .B(mai_mai_n442_), .Y(mai_mai_n1000_));
  NA2        m0972(.A(mai_mai_n226_), .B(mai_mai_n76_), .Y(mai_mai_n1001_));
  NA3        m0973(.A(mai_mai_n1001_), .B(mai_mai_n994_), .C(mai_mai_n993_), .Y(mai_mai_n1002_));
  AOI220     m0974(.A0(mai_mai_n1002_), .A1(mai_mai_n265_), .B0(mai_mai_n1000_), .B1(mai_mai_n999_), .Y(mai_mai_n1003_));
  NA4        m0975(.A(mai_mai_n1003_), .B(mai_mai_n998_), .C(mai_mai_n995_), .D(mai_mai_n991_), .Y(mai_mai_n1004_));
  NO2        m0976(.A(mai_mai_n381_), .B(mai_mai_n89_), .Y(mai_mai_n1005_));
  NA2        m0977(.A(mai_mai_n1005_), .B(mai_mai_n243_), .Y(mai_mai_n1006_));
  NA2        m0978(.A(mai_mai_n669_), .B(mai_mai_n87_), .Y(mai_mai_n1007_));
  NO2        m0979(.A(mai_mai_n465_), .B(mai_mai_n218_), .Y(mai_mai_n1008_));
  AOI220     m0980(.A0(mai_mai_n1008_), .A1(mai_mai_n386_), .B0(mai_mai_n954_), .B1(mai_mai_n222_), .Y(mai_mai_n1009_));
  NA2        m0981(.A(mai_mai_n941_), .B(mai_mai_n951_), .Y(mai_mai_n1010_));
  NA4        m0982(.A(mai_mai_n1010_), .B(mai_mai_n1009_), .C(mai_mai_n1007_), .D(mai_mai_n1006_), .Y(mai_mai_n1011_));
  OAI210     m0983(.A0(mai_mai_n1000_), .A1(mai_mai_n949_), .B0(mai_mai_n556_), .Y(mai_mai_n1012_));
  OAI210     m0984(.A0(mai_mai_n374_), .A1(mai_mai_n373_), .B0(mai_mai_n109_), .Y(mai_mai_n1013_));
  NA2        m0985(.A(mai_mai_n1013_), .B(mai_mai_n548_), .Y(mai_mai_n1014_));
  NA2        m0986(.A(mai_mai_n997_), .B(mai_mai_n939_), .Y(mai_mai_n1015_));
  NA2        m0987(.A(mai_mai_n651_), .B(mai_mai_n543_), .Y(mai_mai_n1016_));
  NA4        m0988(.A(mai_mai_n1016_), .B(mai_mai_n1015_), .C(mai_mai_n1014_), .D(mai_mai_n1012_), .Y(mai_mai_n1017_));
  NO4        m0989(.A(mai_mai_n1017_), .B(mai_mai_n1011_), .C(mai_mai_n1004_), .D(mai_mai_n987_), .Y(mai_mai_n1018_));
  NAi31      m0990(.An(mai_mai_n142_), .B(mai_mai_n424_), .C(n), .Y(mai_mai_n1019_));
  NO3        m0991(.A(mai_mai_n126_), .B(mai_mai_n344_), .C(mai_mai_n861_), .Y(mai_mai_n1020_));
  NO2        m0992(.A(mai_mai_n1020_), .B(mai_mai_n1019_), .Y(mai_mai_n1021_));
  NO3        m0993(.A(mai_mai_n280_), .B(mai_mai_n142_), .C(mai_mai_n412_), .Y(mai_mai_n1022_));
  AOI210     m0994(.A0(mai_mai_n1022_), .A1(mai_mai_n509_), .B0(mai_mai_n1021_), .Y(mai_mai_n1023_));
  INV        m0995(.A(mai_mai_n1023_), .Y(mai_mai_n1024_));
  NA2        m0996(.A(mai_mai_n235_), .B(mai_mai_n173_), .Y(mai_mai_n1025_));
  NO3        m0997(.A(mai_mai_n310_), .B(mai_mai_n447_), .C(mai_mai_n177_), .Y(mai_mai_n1026_));
  NOi31      m0998(.An(mai_mai_n1025_), .B(mai_mai_n1026_), .C(mai_mai_n218_), .Y(mai_mai_n1027_));
  NAi21      m0999(.An(mai_mai_n568_), .B(mai_mai_n1008_), .Y(mai_mai_n1028_));
  NA2        m1000(.A(mai_mai_n440_), .B(mai_mai_n891_), .Y(mai_mai_n1029_));
  NO3        m1001(.A(mai_mai_n441_), .B(mai_mai_n312_), .C(mai_mai_n72_), .Y(mai_mai_n1030_));
  AOI220     m1002(.A0(mai_mai_n1030_), .A1(mai_mai_n1029_), .B0(mai_mai_n490_), .B1(g), .Y(mai_mai_n1031_));
  NA2        m1003(.A(mai_mai_n1031_), .B(mai_mai_n1028_), .Y(mai_mai_n1032_));
  NO2        m1004(.A(mai_mai_n1019_), .B(mai_mai_n238_), .Y(mai_mai_n1033_));
  NA2        m1005(.A(mai_mai_n944_), .B(mai_mai_n936_), .Y(mai_mai_n1034_));
  NO3        m1006(.A(mai_mai_n557_), .B(mai_mai_n151_), .C(mai_mai_n217_), .Y(mai_mai_n1035_));
  OAI210     m1007(.A0(mai_mai_n1035_), .A1(mai_mai_n537_), .B0(mai_mai_n382_), .Y(mai_mai_n1036_));
  OAI220     m1008(.A0(mai_mai_n941_), .A1(mai_mai_n949_), .B0(mai_mai_n558_), .B1(mai_mai_n430_), .Y(mai_mai_n1037_));
  NA4        m1009(.A(mai_mai_n1037_), .B(mai_mai_n1036_), .C(mai_mai_n1034_), .D(mai_mai_n627_), .Y(mai_mai_n1038_));
  OAI210     m1010(.A0(mai_mai_n944_), .A1(mai_mai_n937_), .B0(mai_mai_n1025_), .Y(mai_mai_n1039_));
  NA3        m1011(.A(mai_mai_n985_), .B(mai_mai_n495_), .C(mai_mai_n46_), .Y(mai_mai_n1040_));
  INV        m1012(.A(mai_mai_n334_), .Y(mai_mai_n1041_));
  NA4        m1013(.A(mai_mai_n1041_), .B(mai_mai_n1040_), .C(mai_mai_n1039_), .D(mai_mai_n281_), .Y(mai_mai_n1042_));
  OR3        m1014(.A(mai_mai_n1042_), .B(mai_mai_n1038_), .C(mai_mai_n1033_), .Y(mai_mai_n1043_));
  NO4        m1015(.A(mai_mai_n1043_), .B(mai_mai_n1032_), .C(mai_mai_n1027_), .D(mai_mai_n1024_), .Y(mai_mai_n1044_));
  NA4        m1016(.A(mai_mai_n1044_), .B(mai_mai_n1018_), .C(mai_mai_n977_), .D(mai_mai_n961_), .Y(mai13));
  INV        m1017(.A(mai_mai_n46_), .Y(mai_mai_n1046_));
  AN2        m1018(.A(c), .B(b), .Y(mai_mai_n1047_));
  NA3        m1019(.A(mai_mai_n256_), .B(mai_mai_n1047_), .C(m), .Y(mai_mai_n1048_));
  NA2        m1020(.A(mai_mai_n506_), .B(f), .Y(mai_mai_n1049_));
  NO4        m1021(.A(mai_mai_n1049_), .B(mai_mai_n1048_), .C(mai_mai_n1046_), .D(mai_mai_n597_), .Y(mai_mai_n1050_));
  NA2        m1022(.A(mai_mai_n272_), .B(mai_mai_n1047_), .Y(mai_mai_n1051_));
  NO3        m1023(.A(mai_mai_n1051_), .B(mai_mai_n1049_), .C(mai_mai_n979_), .Y(mai_mai_n1052_));
  NAi32      m1024(.An(d), .Bn(c), .C(e), .Y(mai_mai_n1053_));
  NA2        m1025(.A(mai_mai_n141_), .B(mai_mai_n45_), .Y(mai_mai_n1054_));
  NA2        m1026(.A(mai_mai_n673_), .B(mai_mai_n229_), .Y(mai_mai_n1055_));
  NA2        m1027(.A(mai_mai_n415_), .B(mai_mai_n217_), .Y(mai_mai_n1056_));
  AN2        m1028(.A(d), .B(c), .Y(mai_mai_n1057_));
  NA2        m1029(.A(mai_mai_n1057_), .B(mai_mai_n116_), .Y(mai_mai_n1058_));
  NO4        m1030(.A(mai_mai_n1058_), .B(mai_mai_n1056_), .C(mai_mai_n178_), .D(mai_mai_n169_), .Y(mai_mai_n1059_));
  NA2        m1031(.A(mai_mai_n506_), .B(c), .Y(mai_mai_n1060_));
  NO4        m1032(.A(mai_mai_n1054_), .B(mai_mai_n600_), .C(mai_mai_n1060_), .D(mai_mai_n309_), .Y(mai_mai_n1061_));
  AO210      m1033(.A0(mai_mai_n1059_), .A1(mai_mai_n1055_), .B0(mai_mai_n1061_), .Y(mai_mai_n1062_));
  OR3        m1034(.A(mai_mai_n1062_), .B(mai_mai_n1052_), .C(mai_mai_n1050_), .Y(mai_mai_n1063_));
  NAi32      m1035(.An(f), .Bn(e), .C(c), .Y(mai_mai_n1064_));
  NO2        m1036(.A(mai_mai_n1064_), .B(mai_mai_n148_), .Y(mai_mai_n1065_));
  NA2        m1037(.A(mai_mai_n1065_), .B(g), .Y(mai_mai_n1066_));
  OR3        m1038(.A(mai_mai_n229_), .B(mai_mai_n178_), .C(mai_mai_n169_), .Y(mai_mai_n1067_));
  NO2        m1039(.A(mai_mai_n1067_), .B(mai_mai_n1066_), .Y(mai_mai_n1068_));
  NO2        m1040(.A(mai_mai_n1060_), .B(mai_mai_n309_), .Y(mai_mai_n1069_));
  NO2        m1041(.A(j), .B(mai_mai_n45_), .Y(mai_mai_n1070_));
  NA2        m1042(.A(mai_mai_n637_), .B(mai_mai_n1070_), .Y(mai_mai_n1071_));
  NOi21      m1043(.An(mai_mai_n1069_), .B(mai_mai_n1071_), .Y(mai_mai_n1072_));
  NO2        m1044(.A(mai_mai_n769_), .B(mai_mai_n112_), .Y(mai_mai_n1073_));
  NOi41      m1045(.An(n), .B(m), .C(i), .D(h), .Y(mai_mai_n1074_));
  NA2        m1046(.A(mai_mai_n1074_), .B(mai_mai_n1073_), .Y(mai_mai_n1075_));
  NO2        m1047(.A(mai_mai_n1075_), .B(mai_mai_n1066_), .Y(mai_mai_n1076_));
  OR3        m1048(.A(e), .B(d), .C(c), .Y(mai_mai_n1077_));
  NA3        m1049(.A(k), .B(j), .C(i), .Y(mai_mai_n1078_));
  NO3        m1050(.A(mai_mai_n1078_), .B(mai_mai_n309_), .C(mai_mai_n89_), .Y(mai_mai_n1079_));
  NOi21      m1051(.An(mai_mai_n1079_), .B(mai_mai_n1077_), .Y(mai_mai_n1080_));
  OR4        m1052(.A(mai_mai_n1080_), .B(mai_mai_n1076_), .C(mai_mai_n1072_), .D(mai_mai_n1068_), .Y(mai_mai_n1081_));
  NA3        m1053(.A(mai_mai_n473_), .B(mai_mai_n337_), .C(mai_mai_n56_), .Y(mai_mai_n1082_));
  NO2        m1054(.A(mai_mai_n1082_), .B(mai_mai_n1071_), .Y(mai_mai_n1083_));
  NO4        m1055(.A(mai_mai_n1082_), .B(mai_mai_n600_), .C(mai_mai_n454_), .D(mai_mai_n45_), .Y(mai_mai_n1084_));
  NO2        m1056(.A(f), .B(c), .Y(mai_mai_n1085_));
  NOi21      m1057(.An(mai_mai_n1085_), .B(mai_mai_n446_), .Y(mai_mai_n1086_));
  NA2        m1058(.A(mai_mai_n1086_), .B(mai_mai_n59_), .Y(mai_mai_n1087_));
  OR2        m1059(.A(k), .B(i), .Y(mai_mai_n1088_));
  NO3        m1060(.A(mai_mai_n1088_), .B(mai_mai_n249_), .C(l), .Y(mai_mai_n1089_));
  NOi31      m1061(.An(mai_mai_n1089_), .B(mai_mai_n1087_), .C(j), .Y(mai_mai_n1090_));
  OR3        m1062(.A(mai_mai_n1090_), .B(mai_mai_n1084_), .C(mai_mai_n1083_), .Y(mai_mai_n1091_));
  OR3        m1063(.A(mai_mai_n1091_), .B(mai_mai_n1081_), .C(mai_mai_n1063_), .Y(mai02));
  OR2        m1064(.A(l), .B(k), .Y(mai_mai_n1093_));
  OR3        m1065(.A(h), .B(g), .C(f), .Y(mai_mai_n1094_));
  OR3        m1066(.A(n), .B(m), .C(i), .Y(mai_mai_n1095_));
  NO4        m1067(.A(mai_mai_n1095_), .B(mai_mai_n1094_), .C(mai_mai_n1093_), .D(mai_mai_n1077_), .Y(mai_mai_n1096_));
  NOi31      m1068(.An(e), .B(d), .C(c), .Y(mai_mai_n1097_));
  NA2        m1069(.A(mai_mai_n1079_), .B(mai_mai_n1097_), .Y(mai_mai_n1098_));
  AN3        m1070(.A(g), .B(f), .C(c), .Y(mai_mai_n1099_));
  NA3        m1071(.A(mai_mai_n1099_), .B(mai_mai_n473_), .C(h), .Y(mai_mai_n1100_));
  OR2        m1072(.A(mai_mai_n1078_), .B(mai_mai_n309_), .Y(mai_mai_n1101_));
  OR2        m1073(.A(mai_mai_n1101_), .B(mai_mai_n1100_), .Y(mai_mai_n1102_));
  NO3        m1074(.A(mai_mai_n1082_), .B(mai_mai_n1054_), .C(mai_mai_n600_), .Y(mai_mai_n1103_));
  NO2        m1075(.A(mai_mai_n1103_), .B(mai_mai_n1068_), .Y(mai_mai_n1104_));
  NA3        m1076(.A(l), .B(k), .C(j), .Y(mai_mai_n1105_));
  NA2        m1077(.A(i), .B(h), .Y(mai_mai_n1106_));
  NO3        m1078(.A(mai_mai_n1106_), .B(mai_mai_n1105_), .C(mai_mai_n133_), .Y(mai_mai_n1107_));
  NO3        m1079(.A(mai_mai_n143_), .B(mai_mai_n292_), .C(mai_mai_n218_), .Y(mai_mai_n1108_));
  AOI210     m1080(.A0(mai_mai_n1108_), .A1(mai_mai_n1107_), .B0(mai_mai_n1072_), .Y(mai_mai_n1109_));
  NA3        m1081(.A(c), .B(b), .C(a), .Y(mai_mai_n1110_));
  NO3        m1082(.A(mai_mai_n1110_), .B(mai_mai_n911_), .C(mai_mai_n217_), .Y(mai_mai_n1111_));
  NO4        m1083(.A(mai_mai_n1078_), .B(mai_mai_n301_), .C(mai_mai_n49_), .D(mai_mai_n112_), .Y(mai_mai_n1112_));
  AOI210     m1084(.A0(mai_mai_n1112_), .A1(mai_mai_n1111_), .B0(mai_mai_n1083_), .Y(mai_mai_n1113_));
  AN4        m1085(.A(mai_mai_n1113_), .B(mai_mai_n1109_), .C(mai_mai_n1104_), .D(mai_mai_n1102_), .Y(mai_mai_n1114_));
  NO2        m1086(.A(mai_mai_n1058_), .B(mai_mai_n1056_), .Y(mai_mai_n1115_));
  NA2        m1087(.A(mai_mai_n1075_), .B(mai_mai_n1067_), .Y(mai_mai_n1116_));
  AOI210     m1088(.A0(mai_mai_n1116_), .A1(mai_mai_n1115_), .B0(mai_mai_n1050_), .Y(mai_mai_n1117_));
  NAi41      m1089(.An(mai_mai_n1096_), .B(mai_mai_n1117_), .C(mai_mai_n1114_), .D(mai_mai_n1098_), .Y(mai03));
  NO2        m1090(.A(mai_mai_n539_), .B(mai_mai_n607_), .Y(mai_mai_n1119_));
  NA4        m1091(.A(mai_mai_n588_), .B(m), .C(mai_mai_n112_), .D(mai_mai_n217_), .Y(mai_mai_n1120_));
  NA2        m1092(.A(mai_mai_n1120_), .B(mai_mai_n375_), .Y(mai_mai_n1121_));
  NO3        m1093(.A(mai_mai_n1121_), .B(mai_mai_n1119_), .C(mai_mai_n1013_), .Y(mai_mai_n1122_));
  NOi41      m1094(.An(mai_mai_n816_), .B(mai_mai_n866_), .C(mai_mai_n855_), .D(mai_mai_n721_), .Y(mai_mai_n1123_));
  OAI220     m1095(.A0(mai_mai_n1123_), .A1(mai_mai_n697_), .B0(mai_mai_n1122_), .B1(mai_mai_n601_), .Y(mai_mai_n1124_));
  NOi31      m1096(.An(i), .B(k), .C(j), .Y(mai_mai_n1125_));
  NA4        m1097(.A(mai_mai_n1125_), .B(mai_mai_n1097_), .C(mai_mai_n346_), .D(mai_mai_n337_), .Y(mai_mai_n1126_));
  INV        m1098(.A(mai_mai_n1126_), .Y(mai_mai_n1127_));
  NOi31      m1099(.An(m), .B(n), .C(f), .Y(mai_mai_n1128_));
  NA2        m1100(.A(mai_mai_n1128_), .B(mai_mai_n51_), .Y(mai_mai_n1129_));
  AN2        m1101(.A(e), .B(c), .Y(mai_mai_n1130_));
  NO2        m1102(.A(mai_mai_n898_), .B(mai_mai_n429_), .Y(mai_mai_n1131_));
  NA2        m1103(.A(mai_mai_n519_), .B(l), .Y(mai_mai_n1132_));
  NOi31      m1104(.An(mai_mai_n877_), .B(mai_mai_n1048_), .C(mai_mai_n1132_), .Y(mai_mai_n1133_));
  NO3        m1105(.A(mai_mai_n1133_), .B(mai_mai_n1131_), .C(mai_mai_n1127_), .Y(mai_mai_n1134_));
  NO2        m1106(.A(mai_mai_n292_), .B(a), .Y(mai_mai_n1135_));
  NO2        m1107(.A(mai_mai_n1106_), .B(mai_mai_n493_), .Y(mai_mai_n1136_));
  NO2        m1108(.A(mai_mai_n86_), .B(g), .Y(mai_mai_n1137_));
  AOI210     m1109(.A0(mai_mai_n1137_), .A1(mai_mai_n1136_), .B0(mai_mai_n1089_), .Y(mai_mai_n1138_));
  OR2        m1110(.A(mai_mai_n1138_), .B(mai_mai_n1087_), .Y(mai_mai_n1139_));
  NA2        m1111(.A(mai_mai_n1139_), .B(mai_mai_n1134_), .Y(mai_mai_n1140_));
  NO4        m1112(.A(mai_mai_n1140_), .B(mai_mai_n1124_), .C(mai_mai_n832_), .D(mai_mai_n577_), .Y(mai_mai_n1141_));
  NA2        m1113(.A(c), .B(b), .Y(mai_mai_n1142_));
  NO2        m1114(.A(mai_mai_n709_), .B(mai_mai_n1142_), .Y(mai_mai_n1143_));
  OAI210     m1115(.A0(mai_mai_n875_), .A1(mai_mai_n846_), .B0(mai_mai_n418_), .Y(mai_mai_n1144_));
  OAI210     m1116(.A0(mai_mai_n1144_), .A1(mai_mai_n876_), .B0(mai_mai_n1143_), .Y(mai_mai_n1145_));
  NAi21      m1117(.An(mai_mai_n426_), .B(mai_mai_n1143_), .Y(mai_mai_n1146_));
  NA3        m1118(.A(mai_mai_n430_), .B(mai_mai_n573_), .C(f), .Y(mai_mai_n1147_));
  OAI210     m1119(.A0(mai_mai_n562_), .A1(mai_mai_n39_), .B0(mai_mai_n1135_), .Y(mai_mai_n1148_));
  NA3        m1120(.A(mai_mai_n1148_), .B(mai_mai_n1147_), .C(mai_mai_n1146_), .Y(mai_mai_n1149_));
  NAi21      m1121(.An(f), .B(d), .Y(mai_mai_n1150_));
  NO2        m1122(.A(mai_mai_n1150_), .B(mai_mai_n1110_), .Y(mai_mai_n1151_));
  INV        m1123(.A(mai_mai_n1149_), .Y(mai_mai_n1152_));
  NA3        m1124(.A(mai_mai_n926_), .B(mai_mai_n1132_), .C(mai_mai_n479_), .Y(mai_mai_n1153_));
  NA2        m1125(.A(mai_mai_n160_), .B(mai_mai_n33_), .Y(mai_mai_n1154_));
  AOI210     m1126(.A0(mai_mai_n975_), .A1(mai_mai_n1154_), .B0(mai_mai_n218_), .Y(mai_mai_n1155_));
  OAI210     m1127(.A0(mai_mai_n1155_), .A1(mai_mai_n450_), .B0(mai_mai_n1151_), .Y(mai_mai_n1156_));
  NO2        m1128(.A(mai_mai_n377_), .B(mai_mai_n376_), .Y(mai_mai_n1157_));
  INV        m1129(.A(mai_mai_n969_), .Y(mai_mai_n1158_));
  NAi31      m1130(.An(mai_mai_n1157_), .B(mai_mai_n1158_), .C(mai_mai_n1156_), .Y(mai_mai_n1159_));
  INV        m1131(.A(mai_mai_n1159_), .Y(mai_mai_n1160_));
  NA4        m1132(.A(mai_mai_n1160_), .B(mai_mai_n1152_), .C(mai_mai_n1145_), .D(mai_mai_n1141_), .Y(mai00));
  AOI210     m1133(.A0(mai_mai_n300_), .A1(mai_mai_n218_), .B0(mai_mai_n284_), .Y(mai_mai_n1162_));
  NO2        m1134(.A(mai_mai_n1162_), .B(mai_mai_n591_), .Y(mai_mai_n1163_));
  AOI210     m1135(.A0(mai_mai_n910_), .A1(mai_mai_n951_), .B0(mai_mai_n1127_), .Y(mai_mai_n1164_));
  NO3        m1136(.A(mai_mai_n1103_), .B(mai_mai_n969_), .C(mai_mai_n718_), .Y(mai_mai_n1165_));
  NA3        m1137(.A(mai_mai_n1165_), .B(mai_mai_n1164_), .C(mai_mai_n1014_), .Y(mai_mai_n1166_));
  NA2        m1138(.A(mai_mai_n521_), .B(f), .Y(mai_mai_n1167_));
  OAI210     m1139(.A0(mai_mai_n1020_), .A1(mai_mai_n40_), .B0(mai_mai_n653_), .Y(mai_mai_n1168_));
  NA3        m1140(.A(mai_mai_n1168_), .B(mai_mai_n264_), .C(n), .Y(mai_mai_n1169_));
  AOI210     m1141(.A0(mai_mai_n1169_), .A1(mai_mai_n1167_), .B0(mai_mai_n1058_), .Y(mai_mai_n1170_));
  NO4        m1142(.A(mai_mai_n1170_), .B(mai_mai_n1166_), .C(mai_mai_n1163_), .D(mai_mai_n1081_), .Y(mai_mai_n1171_));
  NA3        m1143(.A(mai_mai_n168_), .B(mai_mai_n46_), .C(mai_mai_n45_), .Y(mai_mai_n1172_));
  NA3        m1144(.A(d), .B(mai_mai_n56_), .C(b), .Y(mai_mai_n1173_));
  NOi31      m1145(.An(n), .B(m), .C(i), .Y(mai_mai_n1174_));
  NA3        m1146(.A(mai_mai_n1174_), .B(mai_mai_n656_), .C(mai_mai_n51_), .Y(mai_mai_n1175_));
  OAI210     m1147(.A0(mai_mai_n1173_), .A1(mai_mai_n1172_), .B0(mai_mai_n1175_), .Y(mai_mai_n1176_));
  INV        m1148(.A(mai_mai_n590_), .Y(mai_mai_n1177_));
  NO3        m1149(.A(mai_mai_n1177_), .B(mai_mai_n1176_), .C(mai_mai_n929_), .Y(mai_mai_n1178_));
  NO4        m1150(.A(mai_mai_n496_), .B(mai_mai_n361_), .C(mai_mai_n1142_), .D(mai_mai_n59_), .Y(mai_mai_n1179_));
  NA3        m1151(.A(mai_mai_n387_), .B(mai_mai_n225_), .C(g), .Y(mai_mai_n1180_));
  OR2        m1152(.A(mai_mai_n1180_), .B(mai_mai_n1173_), .Y(mai_mai_n1181_));
  NO2        m1153(.A(h), .B(g), .Y(mai_mai_n1182_));
  NA4        m1154(.A(mai_mai_n509_), .B(mai_mai_n473_), .C(mai_mai_n1182_), .D(mai_mai_n1047_), .Y(mai_mai_n1183_));
  OAI220     m1155(.A0(mai_mai_n539_), .A1(mai_mai_n607_), .B0(mai_mai_n90_), .B1(mai_mai_n89_), .Y(mai_mai_n1184_));
  AOI220     m1156(.A0(mai_mai_n1184_), .A1(mai_mai_n548_), .B0(mai_mai_n956_), .B1(mai_mai_n589_), .Y(mai_mai_n1185_));
  AOI220     m1157(.A0(mai_mai_n319_), .A1(mai_mai_n253_), .B0(mai_mai_n179_), .B1(mai_mai_n150_), .Y(mai_mai_n1186_));
  NA4        m1158(.A(mai_mai_n1186_), .B(mai_mai_n1185_), .C(mai_mai_n1183_), .D(mai_mai_n1181_), .Y(mai_mai_n1187_));
  NO3        m1159(.A(mai_mai_n1187_), .B(mai_mai_n1179_), .C(mai_mai_n274_), .Y(mai_mai_n1188_));
  INV        m1160(.A(mai_mai_n324_), .Y(mai_mai_n1189_));
  AOI210     m1161(.A0(mai_mai_n253_), .A1(mai_mai_n351_), .B0(mai_mai_n592_), .Y(mai_mai_n1190_));
  NA2        m1162(.A(mai_mai_n1190_), .B(mai_mai_n1189_), .Y(mai_mai_n1191_));
  NA3        m1163(.A(mai_mai_n181_), .B(mai_mai_n112_), .C(g), .Y(mai_mai_n1192_));
  NA3        m1164(.A(mai_mai_n473_), .B(mai_mai_n40_), .C(f), .Y(mai_mai_n1193_));
  NOi31      m1165(.An(mai_mai_n884_), .B(mai_mai_n1193_), .C(mai_mai_n1192_), .Y(mai_mai_n1194_));
  NO2        m1166(.A(mai_mai_n283_), .B(mai_mai_n72_), .Y(mai_mai_n1195_));
  NO3        m1167(.A(mai_mai_n429_), .B(mai_mai_n842_), .C(n), .Y(mai_mai_n1196_));
  AOI210     m1168(.A0(mai_mai_n1196_), .A1(mai_mai_n1195_), .B0(mai_mai_n1096_), .Y(mai_mai_n1197_));
  NAi31      m1169(.An(mai_mai_n1061_), .B(mai_mai_n1197_), .C(mai_mai_n71_), .Y(mai_mai_n1198_));
  NO3        m1170(.A(mai_mai_n1198_), .B(mai_mai_n1194_), .C(mai_mai_n1191_), .Y(mai_mai_n1199_));
  AN3        m1171(.A(mai_mai_n1199_), .B(mai_mai_n1188_), .C(mai_mai_n1178_), .Y(mai_mai_n1200_));
  NA2        m1172(.A(mai_mai_n548_), .B(mai_mai_n100_), .Y(mai_mai_n1201_));
  NA3        m1173(.A(mai_mai_n1128_), .B(mai_mai_n613_), .C(mai_mai_n472_), .Y(mai_mai_n1202_));
  NA3        m1174(.A(mai_mai_n1202_), .B(mai_mai_n1201_), .C(mai_mai_n247_), .Y(mai_mai_n1203_));
  NA2        m1175(.A(mai_mai_n1121_), .B(mai_mai_n548_), .Y(mai_mai_n1204_));
  NA4        m1176(.A(mai_mai_n656_), .B(mai_mai_n209_), .C(mai_mai_n225_), .D(mai_mai_n164_), .Y(mai_mai_n1205_));
  NA2        m1177(.A(mai_mai_n1205_), .B(mai_mai_n1204_), .Y(mai_mai_n1206_));
  OAI210     m1178(.A0(mai_mai_n471_), .A1(mai_mai_n120_), .B0(mai_mai_n878_), .Y(mai_mai_n1207_));
  NA2        m1179(.A(mai_mai_n1207_), .B(mai_mai_n1153_), .Y(mai_mai_n1208_));
  OR4        m1180(.A(mai_mai_n1058_), .B(mai_mai_n280_), .C(mai_mai_n227_), .D(e), .Y(mai_mai_n1209_));
  NO2        m1181(.A(mai_mai_n221_), .B(mai_mai_n218_), .Y(mai_mai_n1210_));
  NA2        m1182(.A(n), .B(e), .Y(mai_mai_n1211_));
  NO2        m1183(.A(mai_mai_n1211_), .B(mai_mai_n148_), .Y(mai_mai_n1212_));
  AOI220     m1184(.A0(mai_mai_n1212_), .A1(mai_mai_n282_), .B0(mai_mai_n859_), .B1(mai_mai_n1210_), .Y(mai_mai_n1213_));
  OAI210     m1185(.A0(mai_mai_n362_), .A1(mai_mai_n314_), .B0(mai_mai_n452_), .Y(mai_mai_n1214_));
  NA4        m1186(.A(mai_mai_n1214_), .B(mai_mai_n1213_), .C(mai_mai_n1209_), .D(mai_mai_n1208_), .Y(mai_mai_n1215_));
  NA2        m1187(.A(mai_mai_n1212_), .B(mai_mai_n863_), .Y(mai_mai_n1216_));
  AOI220     m1188(.A0(mai_mai_n965_), .A1(mai_mai_n589_), .B0(mai_mai_n656_), .B1(mai_mai_n250_), .Y(mai_mai_n1217_));
  NO2        m1189(.A(mai_mai_n65_), .B(h), .Y(mai_mai_n1218_));
  NO3        m1190(.A(mai_mai_n1058_), .B(mai_mai_n1056_), .C(mai_mai_n734_), .Y(mai_mai_n1219_));
  NO2        m1191(.A(mai_mai_n1093_), .B(mai_mai_n133_), .Y(mai_mai_n1220_));
  AN2        m1192(.A(mai_mai_n1220_), .B(mai_mai_n1108_), .Y(mai_mai_n1221_));
  OAI210     m1193(.A0(mai_mai_n1221_), .A1(mai_mai_n1219_), .B0(mai_mai_n1218_), .Y(mai_mai_n1222_));
  NA4        m1194(.A(mai_mai_n1222_), .B(mai_mai_n1217_), .C(mai_mai_n1216_), .D(mai_mai_n879_), .Y(mai_mai_n1223_));
  NO4        m1195(.A(mai_mai_n1223_), .B(mai_mai_n1215_), .C(mai_mai_n1206_), .D(mai_mai_n1203_), .Y(mai_mai_n1224_));
  NA2        m1196(.A(mai_mai_n847_), .B(mai_mai_n764_), .Y(mai_mai_n1225_));
  NA4        m1197(.A(mai_mai_n1225_), .B(mai_mai_n1224_), .C(mai_mai_n1200_), .D(mai_mai_n1171_), .Y(mai01));
  AN2        m1198(.A(mai_mai_n1036_), .B(mai_mai_n1034_), .Y(mai_mai_n1227_));
  NO4        m1199(.A(mai_mai_n812_), .B(mai_mai_n804_), .C(mai_mai_n487_), .D(mai_mai_n290_), .Y(mai_mai_n1228_));
  NA2        m1200(.A(mai_mai_n398_), .B(i), .Y(mai_mai_n1229_));
  NA3        m1201(.A(mai_mai_n1229_), .B(mai_mai_n1228_), .C(mai_mai_n1227_), .Y(mai_mai_n1230_));
  NA2        m1202(.A(mai_mai_n568_), .B(mai_mai_n279_), .Y(mai_mai_n1231_));
  NA2        m1203(.A(mai_mai_n972_), .B(mai_mai_n1231_), .Y(mai_mai_n1232_));
  NA3        m1204(.A(mai_mai_n1232_), .B(mai_mai_n924_), .C(mai_mai_n336_), .Y(mai_mai_n1233_));
  NA2        m1205(.A(mai_mai_n45_), .B(f), .Y(mai_mai_n1234_));
  NA2        m1206(.A(mai_mai_n716_), .B(mai_mai_n95_), .Y(mai_mai_n1235_));
  NO2        m1207(.A(mai_mai_n1235_), .B(mai_mai_n1234_), .Y(mai_mai_n1236_));
  INV        m1208(.A(mai_mai_n118_), .Y(mai_mai_n1237_));
  OA220      m1209(.A0(mai_mai_n1237_), .A1(mai_mai_n599_), .B0(mai_mai_n668_), .B1(mai_mai_n375_), .Y(mai_mai_n1238_));
  NAi41      m1210(.An(mai_mai_n163_), .B(mai_mai_n1238_), .C(mai_mai_n1205_), .D(mai_mai_n909_), .Y(mai_mai_n1239_));
  NO3        m1211(.A(mai_mai_n791_), .B(mai_mai_n680_), .C(mai_mai_n524_), .Y(mai_mai_n1240_));
  NA4        m1212(.A(mai_mai_n716_), .B(mai_mai_n95_), .C(mai_mai_n45_), .D(mai_mai_n217_), .Y(mai_mai_n1241_));
  OA220      m1213(.A0(mai_mai_n1241_), .A1(mai_mai_n676_), .B0(mai_mai_n198_), .B1(mai_mai_n196_), .Y(mai_mai_n1242_));
  NA3        m1214(.A(mai_mai_n1242_), .B(mai_mai_n1240_), .C(mai_mai_n138_), .Y(mai_mai_n1243_));
  NO4        m1215(.A(mai_mai_n1243_), .B(mai_mai_n1239_), .C(mai_mai_n1233_), .D(mai_mai_n1230_), .Y(mai_mai_n1244_));
  INV        m1216(.A(mai_mai_n1180_), .Y(mai_mai_n1245_));
  OAI210     m1217(.A0(mai_mai_n1245_), .A1(mai_mai_n303_), .B0(mai_mai_n543_), .Y(mai_mai_n1246_));
  NA2        m1218(.A(mai_mai_n551_), .B(mai_mai_n400_), .Y(mai_mai_n1247_));
  NOi21      m1219(.An(mai_mai_n574_), .B(mai_mai_n596_), .Y(mai_mai_n1248_));
  NA2        m1220(.A(mai_mai_n1248_), .B(mai_mai_n1247_), .Y(mai_mai_n1249_));
  AOI210     m1221(.A0(mai_mai_n207_), .A1(mai_mai_n88_), .B0(mai_mai_n217_), .Y(mai_mai_n1250_));
  OAI210     m1222(.A0(mai_mai_n819_), .A1(mai_mai_n430_), .B0(mai_mai_n1250_), .Y(mai_mai_n1251_));
  AN3        m1223(.A(m), .B(l), .C(k), .Y(mai_mai_n1252_));
  OAI210     m1224(.A0(mai_mai_n364_), .A1(mai_mai_n34_), .B0(mai_mai_n1252_), .Y(mai_mai_n1253_));
  OR2        m1225(.A(mai_mai_n1253_), .B(mai_mai_n335_), .Y(mai_mai_n1254_));
  NA4        m1226(.A(mai_mai_n1254_), .B(mai_mai_n1251_), .C(mai_mai_n1249_), .D(mai_mai_n1246_), .Y(mai_mai_n1255_));
  INV        m1227(.A(mai_mai_n608_), .Y(mai_mai_n1256_));
  OAI210     m1228(.A0(mai_mai_n1237_), .A1(mai_mai_n605_), .B0(mai_mai_n1256_), .Y(mai_mai_n1257_));
  NA2        m1229(.A(mai_mai_n289_), .B(mai_mai_n198_), .Y(mai_mai_n1258_));
  NA2        m1230(.A(mai_mai_n1258_), .B(mai_mai_n672_), .Y(mai_mai_n1259_));
  INV        m1231(.A(mai_mai_n969_), .Y(mai_mai_n1260_));
  OAI210     m1232(.A0(mai_mai_n1236_), .A1(mai_mai_n329_), .B0(mai_mai_n681_), .Y(mai_mai_n1261_));
  NA4        m1233(.A(mai_mai_n1261_), .B(mai_mai_n1260_), .C(mai_mai_n1259_), .D(mai_mai_n794_), .Y(mai_mai_n1262_));
  NO3        m1234(.A(mai_mai_n1262_), .B(mai_mai_n1257_), .C(mai_mai_n1255_), .Y(mai_mai_n1263_));
  NA2        m1235(.A(mai_mai_n516_), .B(mai_mai_n58_), .Y(mai_mai_n1264_));
  NO2        m1236(.A(mai_mai_n1241_), .B(mai_mai_n992_), .Y(mai_mai_n1265_));
  NO2        m1237(.A(mai_mai_n210_), .B(mai_mai_n111_), .Y(mai_mai_n1266_));
  NO3        m1238(.A(mai_mai_n1266_), .B(mai_mai_n1265_), .C(mai_mai_n1176_), .Y(mai_mai_n1267_));
  NA3        m1239(.A(mai_mai_n1267_), .B(mai_mai_n1264_), .C(mai_mai_n763_), .Y(mai_mai_n1268_));
  NO2        m1240(.A(mai_mai_n979_), .B(mai_mai_n237_), .Y(mai_mai_n1269_));
  NO2        m1241(.A(mai_mai_n980_), .B(mai_mai_n570_), .Y(mai_mai_n1270_));
  OAI210     m1242(.A0(mai_mai_n1270_), .A1(mai_mai_n1269_), .B0(mai_mai_n344_), .Y(mai_mai_n1271_));
  NA2        m1243(.A(mai_mai_n584_), .B(mai_mai_n582_), .Y(mai_mai_n1272_));
  NO3        m1244(.A(mai_mai_n78_), .B(mai_mai_n301_), .C(mai_mai_n45_), .Y(mai_mai_n1273_));
  NA2        m1245(.A(mai_mai_n1273_), .B(mai_mai_n567_), .Y(mai_mai_n1274_));
  NA2        m1246(.A(mai_mai_n1274_), .B(mai_mai_n1272_), .Y(mai_mai_n1275_));
  OR2        m1247(.A(mai_mai_n1180_), .B(mai_mai_n1173_), .Y(mai_mai_n1276_));
  NA2        m1248(.A(mai_mai_n1273_), .B(mai_mai_n822_), .Y(mai_mai_n1277_));
  NA3        m1249(.A(mai_mai_n1277_), .B(mai_mai_n1276_), .C(mai_mai_n390_), .Y(mai_mai_n1278_));
  NOi41      m1250(.An(mai_mai_n1271_), .B(mai_mai_n1278_), .C(mai_mai_n1275_), .D(mai_mai_n1268_), .Y(mai_mai_n1279_));
  NO2        m1251(.A(mai_mai_n132_), .B(mai_mai_n45_), .Y(mai_mai_n1280_));
  NO2        m1252(.A(mai_mai_n45_), .B(mai_mai_n40_), .Y(mai_mai_n1281_));
  AO220      m1253(.A0(mai_mai_n1281_), .A1(mai_mai_n630_), .B0(mai_mai_n1280_), .B1(mai_mai_n714_), .Y(mai_mai_n1282_));
  NA2        m1254(.A(mai_mai_n1282_), .B(mai_mai_n344_), .Y(mai_mai_n1283_));
  INV        m1255(.A(mai_mai_n136_), .Y(mai_mai_n1284_));
  NO3        m1256(.A(mai_mai_n1106_), .B(mai_mai_n178_), .C(mai_mai_n86_), .Y(mai_mai_n1285_));
  AOI220     m1257(.A0(mai_mai_n1285_), .A1(mai_mai_n1284_), .B0(mai_mai_n1273_), .B1(mai_mai_n983_), .Y(mai_mai_n1286_));
  NA2        m1258(.A(mai_mai_n1286_), .B(mai_mai_n1283_), .Y(mai_mai_n1287_));
  NO2        m1259(.A(mai_mai_n621_), .B(mai_mai_n620_), .Y(mai_mai_n1288_));
  NO4        m1260(.A(mai_mai_n1106_), .B(mai_mai_n1288_), .C(mai_mai_n176_), .D(mai_mai_n86_), .Y(mai_mai_n1289_));
  NO3        m1261(.A(mai_mai_n1289_), .B(mai_mai_n1287_), .C(mai_mai_n645_), .Y(mai_mai_n1290_));
  NA4        m1262(.A(mai_mai_n1290_), .B(mai_mai_n1279_), .C(mai_mai_n1263_), .D(mai_mai_n1244_), .Y(mai06));
  NO2        m1263(.A(mai_mai_n229_), .B(mai_mai_n102_), .Y(mai_mai_n1292_));
  OAI210     m1264(.A0(mai_mai_n1292_), .A1(mai_mai_n1285_), .B0(mai_mai_n386_), .Y(mai_mai_n1293_));
  NO3        m1265(.A(mai_mai_n609_), .B(mai_mai_n817_), .C(mai_mai_n610_), .Y(mai_mai_n1294_));
  OR2        m1266(.A(mai_mai_n1294_), .B(mai_mai_n898_), .Y(mai_mai_n1295_));
  NA3        m1267(.A(mai_mai_n1295_), .B(mai_mai_n1293_), .C(mai_mai_n1271_), .Y(mai_mai_n1296_));
  NO3        m1268(.A(mai_mai_n1296_), .B(mai_mai_n1275_), .C(mai_mai_n263_), .Y(mai_mai_n1297_));
  NO2        m1269(.A(mai_mai_n301_), .B(mai_mai_n45_), .Y(mai_mai_n1298_));
  AOI210     m1270(.A0(mai_mai_n1298_), .A1(mai_mai_n984_), .B0(mai_mai_n1269_), .Y(mai_mai_n1299_));
  AOI210     m1271(.A0(mai_mai_n1298_), .A1(mai_mai_n571_), .B0(mai_mai_n1282_), .Y(mai_mai_n1300_));
  AOI210     m1272(.A0(mai_mai_n1300_), .A1(mai_mai_n1299_), .B0(mai_mai_n341_), .Y(mai_mai_n1301_));
  OAI210     m1273(.A0(mai_mai_n88_), .A1(mai_mai_n40_), .B0(mai_mai_n679_), .Y(mai_mai_n1302_));
  NA2        m1274(.A(mai_mai_n1302_), .B(mai_mai_n649_), .Y(mai_mai_n1303_));
  NO2        m1275(.A(mai_mai_n527_), .B(mai_mai_n173_), .Y(mai_mai_n1304_));
  NO2        m1276(.A(mai_mai_n614_), .B(mai_mai_n1129_), .Y(mai_mai_n1305_));
  OAI210     m1277(.A0(mai_mai_n466_), .A1(mai_mai_n254_), .B0(mai_mai_n918_), .Y(mai_mai_n1306_));
  NO3        m1278(.A(mai_mai_n1306_), .B(mai_mai_n1305_), .C(mai_mai_n1304_), .Y(mai_mai_n1307_));
  NO2        m1279(.A(mai_mai_n374_), .B(mai_mai_n137_), .Y(mai_mai_n1308_));
  AOI210     m1280(.A0(mai_mai_n1308_), .A1(mai_mai_n602_), .B0(mai_mai_n608_), .Y(mai_mai_n1309_));
  NA3        m1281(.A(mai_mai_n1309_), .B(mai_mai_n1307_), .C(mai_mai_n1303_), .Y(mai_mai_n1310_));
  NO2        m1282(.A(mai_mai_n756_), .B(mai_mai_n373_), .Y(mai_mai_n1311_));
  NO3        m1283(.A(mai_mai_n681_), .B(mai_mai_n765_), .C(mai_mai_n641_), .Y(mai_mai_n1312_));
  NOi21      m1284(.An(mai_mai_n1311_), .B(mai_mai_n1312_), .Y(mai_mai_n1313_));
  AN2        m1285(.A(mai_mai_n965_), .B(mai_mai_n652_), .Y(mai_mai_n1314_));
  NO4        m1286(.A(mai_mai_n1314_), .B(mai_mai_n1313_), .C(mai_mai_n1310_), .D(mai_mai_n1301_), .Y(mai_mai_n1315_));
  NO2        m1287(.A(mai_mai_n811_), .B(mai_mai_n285_), .Y(mai_mai_n1316_));
  OAI220     m1288(.A0(mai_mai_n740_), .A1(mai_mai_n47_), .B0(mai_mai_n229_), .B1(mai_mai_n623_), .Y(mai_mai_n1317_));
  OAI210     m1289(.A0(mai_mai_n285_), .A1(c), .B0(mai_mai_n648_), .Y(mai_mai_n1318_));
  AOI220     m1290(.A0(mai_mai_n1318_), .A1(mai_mai_n1317_), .B0(mai_mai_n1316_), .B1(mai_mai_n275_), .Y(mai_mai_n1319_));
  NO3        m1291(.A(mai_mai_n249_), .B(mai_mai_n102_), .C(mai_mai_n292_), .Y(mai_mai_n1320_));
  OAI220     m1292(.A0(mai_mai_n706_), .A1(mai_mai_n254_), .B0(mai_mai_n523_), .B1(mai_mai_n527_), .Y(mai_mai_n1321_));
  OAI210     m1293(.A0(l), .A1(i), .B0(k), .Y(mai_mai_n1322_));
  NO3        m1294(.A(mai_mai_n1322_), .B(mai_mai_n607_), .C(j), .Y(mai_mai_n1323_));
  NOi21      m1295(.An(mai_mai_n1323_), .B(mai_mai_n676_), .Y(mai_mai_n1324_));
  NO4        m1296(.A(mai_mai_n1324_), .B(mai_mai_n1321_), .C(mai_mai_n1320_), .D(mai_mai_n1131_), .Y(mai_mai_n1325_));
  NA3        m1297(.A(mai_mai_n802_), .B(mai_mai_n801_), .C(mai_mai_n440_), .Y(mai_mai_n1326_));
  NAi31      m1298(.An(mai_mai_n756_), .B(mai_mai_n1326_), .C(mai_mai_n206_), .Y(mai_mai_n1327_));
  NA4        m1299(.A(mai_mai_n1327_), .B(mai_mai_n1325_), .C(mai_mai_n1319_), .D(mai_mai_n1217_), .Y(mai_mai_n1328_));
  NOi31      m1300(.An(mai_mai_n1294_), .B(mai_mai_n470_), .C(mai_mai_n399_), .Y(mai_mai_n1329_));
  OR3        m1301(.A(mai_mai_n1329_), .B(mai_mai_n790_), .C(mai_mai_n554_), .Y(mai_mai_n1330_));
  NA2        m1302(.A(mai_mai_n584_), .B(mai_mai_n452_), .Y(mai_mai_n1331_));
  NA2        m1303(.A(mai_mai_n1323_), .B(mai_mai_n798_), .Y(mai_mai_n1332_));
  NA3        m1304(.A(mai_mai_n1332_), .B(mai_mai_n1331_), .C(mai_mai_n1330_), .Y(mai_mai_n1333_));
  AN2        m1305(.A(mai_mai_n937_), .B(mai_mai_n936_), .Y(mai_mai_n1334_));
  NO4        m1306(.A(mai_mai_n1334_), .B(mai_mai_n889_), .C(mai_mai_n512_), .D(mai_mai_n490_), .Y(mai_mai_n1335_));
  NA2        m1307(.A(mai_mai_n1335_), .B(mai_mai_n1277_), .Y(mai_mai_n1336_));
  NAi21      m1308(.An(j), .B(i), .Y(mai_mai_n1337_));
  NO4        m1309(.A(mai_mai_n1288_), .B(mai_mai_n1337_), .C(mai_mai_n446_), .D(mai_mai_n240_), .Y(mai_mai_n1338_));
  NO4        m1310(.A(mai_mai_n1338_), .B(mai_mai_n1336_), .C(mai_mai_n1333_), .D(mai_mai_n1328_), .Y(mai_mai_n1339_));
  NA4        m1311(.A(mai_mai_n1339_), .B(mai_mai_n1315_), .C(mai_mai_n1297_), .D(mai_mai_n1290_), .Y(mai07));
  NOi21      m1312(.An(j), .B(k), .Y(mai_mai_n1341_));
  NA4        m1313(.A(mai_mai_n181_), .B(mai_mai_n108_), .C(mai_mai_n1341_), .D(f), .Y(mai_mai_n1342_));
  NAi32      m1314(.An(m), .Bn(b), .C(n), .Y(mai_mai_n1343_));
  NO3        m1315(.A(mai_mai_n1343_), .B(g), .C(f), .Y(mai_mai_n1344_));
  OAI210     m1316(.A0(mai_mai_n323_), .A1(mai_mai_n492_), .B0(mai_mai_n1344_), .Y(mai_mai_n1345_));
  NAi21      m1317(.An(f), .B(c), .Y(mai_mai_n1346_));
  OR2        m1318(.A(e), .B(d), .Y(mai_mai_n1347_));
  OAI220     m1319(.A0(mai_mai_n1347_), .A1(mai_mai_n1346_), .B0(mai_mai_n636_), .B1(mai_mai_n325_), .Y(mai_mai_n1348_));
  NA3        m1320(.A(mai_mai_n1348_), .B(mai_mai_n1070_), .C(mai_mai_n181_), .Y(mai_mai_n1349_));
  NOi31      m1321(.An(n), .B(m), .C(b), .Y(mai_mai_n1350_));
  NO3        m1322(.A(mai_mai_n133_), .B(mai_mai_n454_), .C(h), .Y(mai_mai_n1351_));
  NA3        m1323(.A(mai_mai_n1349_), .B(mai_mai_n1345_), .C(mai_mai_n1342_), .Y(mai_mai_n1352_));
  NOi41      m1324(.An(i), .B(n), .C(m), .D(h), .Y(mai_mai_n1353_));
  NOi21      m1325(.An(h), .B(k), .Y(mai_mai_n1354_));
  NO2        m1326(.A(k), .B(i), .Y(mai_mai_n1355_));
  NA3        m1327(.A(mai_mai_n1355_), .B(mai_mai_n908_), .C(mai_mai_n181_), .Y(mai_mai_n1356_));
  NA2        m1328(.A(mai_mai_n86_), .B(mai_mai_n45_), .Y(mai_mai_n1357_));
  NO2        m1329(.A(mai_mai_n1064_), .B(mai_mai_n446_), .Y(mai_mai_n1358_));
  NA3        m1330(.A(mai_mai_n1358_), .B(mai_mai_n1357_), .C(mai_mai_n218_), .Y(mai_mai_n1359_));
  NO2        m1331(.A(mai_mai_n1078_), .B(mai_mai_n309_), .Y(mai_mai_n1360_));
  NA2        m1332(.A(mai_mai_n555_), .B(mai_mai_n79_), .Y(mai_mai_n1361_));
  NA2        m1333(.A(mai_mai_n1218_), .B(mai_mai_n295_), .Y(mai_mai_n1362_));
  NA4        m1334(.A(mai_mai_n1362_), .B(mai_mai_n1361_), .C(mai_mai_n1359_), .D(mai_mai_n1356_), .Y(mai_mai_n1363_));
  NO2        m1335(.A(mai_mai_n1363_), .B(mai_mai_n1352_), .Y(mai_mai_n1364_));
  NO3        m1336(.A(e), .B(d), .C(c), .Y(mai_mai_n1365_));
  OAI210     m1337(.A0(mai_mai_n133_), .A1(mai_mai_n218_), .B0(mai_mai_n612_), .Y(mai_mai_n1366_));
  NA2        m1338(.A(mai_mai_n1366_), .B(mai_mai_n1365_), .Y(mai_mai_n1367_));
  NO2        m1339(.A(mai_mai_n1367_), .B(c), .Y(mai_mai_n1368_));
  OR2        m1340(.A(h), .B(f), .Y(mai_mai_n1369_));
  NO3        m1341(.A(n), .B(m), .C(i), .Y(mai_mai_n1370_));
  OAI210     m1342(.A0(mai_mai_n1130_), .A1(mai_mai_n158_), .B0(mai_mai_n1370_), .Y(mai_mai_n1371_));
  NO2        m1343(.A(mai_mai_n1371_), .B(mai_mai_n1369_), .Y(mai_mai_n1372_));
  NA3        m1344(.A(mai_mai_n703_), .B(mai_mai_n689_), .C(mai_mai_n112_), .Y(mai_mai_n1373_));
  NO2        m1345(.A(mai_mai_n1373_), .B(mai_mai_n45_), .Y(mai_mai_n1374_));
  NA2        m1346(.A(mai_mai_n1370_), .B(mai_mai_n647_), .Y(mai_mai_n1375_));
  NO2        m1347(.A(l), .B(k), .Y(mai_mai_n1376_));
  NOi41      m1348(.An(mai_mai_n560_), .B(mai_mai_n1376_), .C(mai_mai_n485_), .D(mai_mai_n446_), .Y(mai_mai_n1377_));
  NO3        m1349(.A(mai_mai_n446_), .B(d), .C(c), .Y(mai_mai_n1378_));
  NO4        m1350(.A(mai_mai_n1377_), .B(mai_mai_n1374_), .C(mai_mai_n1372_), .D(mai_mai_n1368_), .Y(mai_mai_n1379_));
  NO2        m1351(.A(mai_mai_n149_), .B(h), .Y(mai_mai_n1380_));
  NO2        m1352(.A(mai_mai_n1088_), .B(l), .Y(mai_mai_n1381_));
  NO2        m1353(.A(g), .B(c), .Y(mai_mai_n1382_));
  NA3        m1354(.A(mai_mai_n1382_), .B(mai_mai_n143_), .C(mai_mai_n189_), .Y(mai_mai_n1383_));
  NO2        m1355(.A(mai_mai_n1383_), .B(mai_mai_n1381_), .Y(mai_mai_n1384_));
  NA2        m1356(.A(mai_mai_n1384_), .B(mai_mai_n181_), .Y(mai_mai_n1385_));
  NA2        m1357(.A(mai_mai_n1354_), .B(mai_mai_n1088_), .Y(mai_mai_n1386_));
  NO2        m1358(.A(mai_mai_n457_), .B(a), .Y(mai_mai_n1387_));
  NA3        m1359(.A(mai_mai_n1387_), .B(mai_mai_n1386_), .C(mai_mai_n113_), .Y(mai_mai_n1388_));
  NO2        m1360(.A(i), .B(h), .Y(mai_mai_n1389_));
  NA2        m1361(.A(mai_mai_n1389_), .B(mai_mai_n225_), .Y(mai_mai_n1390_));
  AOI210     m1362(.A0(mai_mai_n1150_), .A1(h), .B0(mai_mai_n419_), .Y(mai_mai_n1391_));
  NA2        m1363(.A(mai_mai_n139_), .B(mai_mai_n225_), .Y(mai_mai_n1392_));
  AOI210     m1364(.A0(mai_mai_n264_), .A1(mai_mai_n116_), .B0(mai_mai_n543_), .Y(mai_mai_n1393_));
  OAI220     m1365(.A0(mai_mai_n1393_), .A1(mai_mai_n1390_), .B0(mai_mai_n1392_), .B1(mai_mai_n1391_), .Y(mai_mai_n1394_));
  NO2        m1366(.A(mai_mai_n762_), .B(mai_mai_n190_), .Y(mai_mai_n1395_));
  NOi31      m1367(.An(m), .B(n), .C(b), .Y(mai_mai_n1396_));
  NOi31      m1368(.An(f), .B(d), .C(c), .Y(mai_mai_n1397_));
  NA2        m1369(.A(mai_mai_n1397_), .B(mai_mai_n1396_), .Y(mai_mai_n1398_));
  INV        m1370(.A(mai_mai_n1398_), .Y(mai_mai_n1399_));
  NO3        m1371(.A(mai_mai_n1399_), .B(mai_mai_n1395_), .C(mai_mai_n1394_), .Y(mai_mai_n1400_));
  NA2        m1372(.A(mai_mai_n1099_), .B(mai_mai_n473_), .Y(mai_mai_n1401_));
  NO4        m1373(.A(mai_mai_n1401_), .B(mai_mai_n1073_), .C(mai_mai_n446_), .D(mai_mai_n45_), .Y(mai_mai_n1402_));
  OAI210     m1374(.A0(mai_mai_n184_), .A1(mai_mai_n538_), .B0(mai_mai_n1074_), .Y(mai_mai_n1403_));
  NO3        m1375(.A(mai_mai_n41_), .B(i), .C(h), .Y(mai_mai_n1404_));
  INV        m1376(.A(mai_mai_n1403_), .Y(mai_mai_n1405_));
  NO2        m1377(.A(mai_mai_n1405_), .B(mai_mai_n1402_), .Y(mai_mai_n1406_));
  AN4        m1378(.A(mai_mai_n1406_), .B(mai_mai_n1400_), .C(mai_mai_n1388_), .D(mai_mai_n1385_), .Y(mai_mai_n1407_));
  NA2        m1379(.A(mai_mai_n1350_), .B(mai_mai_n383_), .Y(mai_mai_n1408_));
  NO2        m1380(.A(mai_mai_n1408_), .B(mai_mai_n1055_), .Y(mai_mai_n1409_));
  NA2        m1381(.A(mai_mai_n1378_), .B(mai_mai_n219_), .Y(mai_mai_n1410_));
  NO2        m1382(.A(mai_mai_n190_), .B(b), .Y(mai_mai_n1411_));
  AOI220     m1383(.A0(mai_mai_n1174_), .A1(mai_mai_n1411_), .B0(mai_mai_n1107_), .B1(mai_mai_n1401_), .Y(mai_mai_n1412_));
  NAi31      m1384(.An(mai_mai_n1409_), .B(mai_mai_n1412_), .C(mai_mai_n1410_), .Y(mai_mai_n1413_));
  NO4        m1385(.A(mai_mai_n133_), .B(g), .C(f), .D(e), .Y(mai_mai_n1414_));
  NA3        m1386(.A(mai_mai_n1355_), .B(mai_mai_n296_), .C(h), .Y(mai_mai_n1415_));
  NA2        m1387(.A(mai_mai_n197_), .B(mai_mai_n97_), .Y(mai_mai_n1416_));
  OR2        m1388(.A(e), .B(a), .Y(mai_mai_n1417_));
  NO2        m1389(.A(mai_mai_n1347_), .B(mai_mai_n1346_), .Y(mai_mai_n1418_));
  AOI210     m1390(.A0(mai_mai_n30_), .A1(h), .B0(mai_mai_n1418_), .Y(mai_mai_n1419_));
  NO2        m1391(.A(mai_mai_n1419_), .B(mai_mai_n1095_), .Y(mai_mai_n1420_));
  NA2        m1392(.A(mai_mai_n1353_), .B(mai_mai_n1376_), .Y(mai_mai_n1421_));
  INV        m1393(.A(mai_mai_n1421_), .Y(mai_mai_n1422_));
  OR3        m1394(.A(mai_mai_n554_), .B(mai_mai_n553_), .C(mai_mai_n112_), .Y(mai_mai_n1423_));
  NA2        m1395(.A(mai_mai_n1128_), .B(mai_mai_n412_), .Y(mai_mai_n1424_));
  OAI220     m1396(.A0(mai_mai_n1424_), .A1(mai_mai_n439_), .B0(mai_mai_n1423_), .B1(mai_mai_n301_), .Y(mai_mai_n1425_));
  AO210      m1397(.A0(mai_mai_n1425_), .A1(mai_mai_n116_), .B0(mai_mai_n1422_), .Y(mai_mai_n1426_));
  NO3        m1398(.A(mai_mai_n1426_), .B(mai_mai_n1420_), .C(mai_mai_n1413_), .Y(mai_mai_n1427_));
  NA4        m1399(.A(mai_mai_n1427_), .B(mai_mai_n1407_), .C(mai_mai_n1379_), .D(mai_mai_n1364_), .Y(mai_mai_n1428_));
  NO2        m1400(.A(mai_mai_n1142_), .B(mai_mai_n110_), .Y(mai_mai_n1429_));
  NA2        m1401(.A(mai_mai_n383_), .B(mai_mai_n56_), .Y(mai_mai_n1430_));
  AOI210     m1402(.A0(mai_mai_n1430_), .A1(mai_mai_n1064_), .B0(mai_mai_n1375_), .Y(mai_mai_n1431_));
  NA2        m1403(.A(mai_mai_n219_), .B(mai_mai_n181_), .Y(mai_mai_n1432_));
  AOI210     m1404(.A0(mai_mai_n1432_), .A1(mai_mai_n1192_), .B0(mai_mai_n1430_), .Y(mai_mai_n1433_));
  NO2        m1405(.A(mai_mai_n1100_), .B(mai_mai_n1095_), .Y(mai_mai_n1434_));
  NO3        m1406(.A(mai_mai_n1434_), .B(mai_mai_n1433_), .C(mai_mai_n1431_), .Y(mai_mai_n1435_));
  NO2        m1407(.A(mai_mai_n395_), .B(j), .Y(mai_mai_n1436_));
  NA3        m1408(.A(mai_mai_n1404_), .B(mai_mai_n1347_), .C(mai_mai_n1128_), .Y(mai_mai_n1437_));
  NAi41      m1409(.An(mai_mai_n1389_), .B(mai_mai_n1086_), .C(mai_mai_n169_), .D(mai_mai_n152_), .Y(mai_mai_n1438_));
  NA2        m1410(.A(mai_mai_n1438_), .B(mai_mai_n1437_), .Y(mai_mai_n1439_));
  NA3        m1411(.A(g), .B(mai_mai_n1436_), .C(mai_mai_n160_), .Y(mai_mai_n1440_));
  INV        m1412(.A(mai_mai_n1440_), .Y(mai_mai_n1441_));
  NO3        m1413(.A(mai_mai_n756_), .B(mai_mai_n176_), .C(mai_mai_n415_), .Y(mai_mai_n1442_));
  NO3        m1414(.A(mai_mai_n1442_), .B(mai_mai_n1441_), .C(mai_mai_n1439_), .Y(mai_mai_n1443_));
  AOI210     m1415(.A0(mai_mai_n1432_), .A1(mai_mai_n1416_), .B0(mai_mai_n1064_), .Y(mai_mai_n1444_));
  OR2        m1416(.A(n), .B(i), .Y(mai_mai_n1445_));
  OAI210     m1417(.A0(mai_mai_n1445_), .A1(mai_mai_n1085_), .B0(mai_mai_n49_), .Y(mai_mai_n1446_));
  AOI220     m1418(.A0(mai_mai_n1446_), .A1(mai_mai_n1182_), .B0(mai_mai_n835_), .B1(mai_mai_n197_), .Y(mai_mai_n1447_));
  INV        m1419(.A(mai_mai_n1447_), .Y(mai_mai_n1448_));
  OAI220     m1420(.A0(mai_mai_n673_), .A1(g), .B0(mai_mai_n229_), .B1(c), .Y(mai_mai_n1449_));
  AOI210     m1421(.A0(mai_mai_n1411_), .A1(mai_mai_n41_), .B0(mai_mai_n1449_), .Y(mai_mai_n1450_));
  NO2        m1422(.A(mai_mai_n133_), .B(l), .Y(mai_mai_n1451_));
  NO2        m1423(.A(mai_mai_n229_), .B(k), .Y(mai_mai_n1452_));
  OAI210     m1424(.A0(mai_mai_n1452_), .A1(mai_mai_n1389_), .B0(mai_mai_n1451_), .Y(mai_mai_n1453_));
  OAI220     m1425(.A0(mai_mai_n1453_), .A1(mai_mai_n31_), .B0(mai_mai_n1450_), .B1(mai_mai_n178_), .Y(mai_mai_n1454_));
  NO3        m1426(.A(mai_mai_n1423_), .B(mai_mai_n473_), .C(mai_mai_n358_), .Y(mai_mai_n1455_));
  NO4        m1427(.A(mai_mai_n1455_), .B(mai_mai_n1454_), .C(mai_mai_n1448_), .D(mai_mai_n1444_), .Y(mai_mai_n1456_));
  NO3        m1428(.A(mai_mai_n1110_), .B(mai_mai_n1347_), .C(mai_mai_n49_), .Y(mai_mai_n1457_));
  NO2        m1429(.A(mai_mai_n1095_), .B(h), .Y(mai_mai_n1458_));
  NA3        m1430(.A(mai_mai_n1458_), .B(d), .C(mai_mai_n1056_), .Y(mai_mai_n1459_));
  NO2        m1431(.A(mai_mai_n1459_), .B(c), .Y(mai_mai_n1460_));
  NA3        m1432(.A(mai_mai_n1429_), .B(mai_mai_n473_), .C(f), .Y(mai_mai_n1461_));
  NA2        m1433(.A(mai_mai_n181_), .B(mai_mai_n112_), .Y(mai_mai_n1462_));
  NO2        m1434(.A(mai_mai_n1341_), .B(mai_mai_n42_), .Y(mai_mai_n1463_));
  AOI210     m1435(.A0(mai_mai_n113_), .A1(mai_mai_n40_), .B0(mai_mai_n1463_), .Y(mai_mai_n1464_));
  NO2        m1436(.A(mai_mai_n1464_), .B(mai_mai_n1461_), .Y(mai_mai_n1465_));
  NO2        m1437(.A(mai_mai_n1337_), .B(mai_mai_n176_), .Y(mai_mai_n1466_));
  NOi21      m1438(.An(d), .B(f), .Y(mai_mai_n1467_));
  NO3        m1439(.A(mai_mai_n1397_), .B(mai_mai_n1467_), .C(mai_mai_n40_), .Y(mai_mai_n1468_));
  NA2        m1440(.A(mai_mai_n1468_), .B(mai_mai_n1466_), .Y(mai_mai_n1469_));
  NO2        m1441(.A(mai_mai_n1347_), .B(f), .Y(mai_mai_n1470_));
  NA2        m1442(.A(mai_mai_n1387_), .B(mai_mai_n1463_), .Y(mai_mai_n1471_));
  NA2        m1443(.A(mai_mai_n1471_), .B(mai_mai_n1469_), .Y(mai_mai_n1472_));
  NO3        m1444(.A(mai_mai_n1472_), .B(mai_mai_n1465_), .C(mai_mai_n1460_), .Y(mai_mai_n1473_));
  NA4        m1445(.A(mai_mai_n1473_), .B(mai_mai_n1456_), .C(mai_mai_n1443_), .D(mai_mai_n1435_), .Y(mai_mai_n1474_));
  NO3        m1446(.A(mai_mai_n1099_), .B(mai_mai_n1085_), .C(mai_mai_n40_), .Y(mai_mai_n1475_));
  NO2        m1447(.A(mai_mai_n473_), .B(mai_mai_n301_), .Y(mai_mai_n1476_));
  OAI210     m1448(.A0(mai_mai_n1476_), .A1(mai_mai_n1475_), .B0(mai_mai_n1360_), .Y(mai_mai_n1477_));
  OAI210     m1449(.A0(mai_mai_n1414_), .A1(mai_mai_n1350_), .B0(mai_mai_n895_), .Y(mai_mai_n1478_));
  NO2        m1450(.A(mai_mai_n1053_), .B(mai_mai_n133_), .Y(mai_mai_n1479_));
  NA2        m1451(.A(mai_mai_n1479_), .B(mai_mai_n629_), .Y(mai_mai_n1480_));
  NA3        m1452(.A(mai_mai_n1480_), .B(mai_mai_n1478_), .C(mai_mai_n1477_), .Y(mai_mai_n1481_));
  NA2        m1453(.A(mai_mai_n1382_), .B(mai_mai_n1467_), .Y(mai_mai_n1482_));
  NO2        m1454(.A(mai_mai_n1482_), .B(m), .Y(mai_mai_n1483_));
  NO2        m1455(.A(mai_mai_n153_), .B(mai_mai_n183_), .Y(mai_mai_n1484_));
  OAI210     m1456(.A0(mai_mai_n1484_), .A1(mai_mai_n110_), .B0(mai_mai_n1396_), .Y(mai_mai_n1485_));
  INV        m1457(.A(mai_mai_n1485_), .Y(mai_mai_n1486_));
  NO3        m1458(.A(mai_mai_n1486_), .B(mai_mai_n1483_), .C(mai_mai_n1481_), .Y(mai_mai_n1487_));
  NO2        m1459(.A(mai_mai_n1346_), .B(e), .Y(mai_mai_n1488_));
  NA2        m1460(.A(mai_mai_n1488_), .B(mai_mai_n410_), .Y(mai_mai_n1489_));
  OAI210     m1461(.A0(mai_mai_n1470_), .A1(mai_mai_n1137_), .B0(mai_mai_n640_), .Y(mai_mai_n1490_));
  OR3        m1462(.A(mai_mai_n1452_), .B(mai_mai_n1218_), .C(mai_mai_n133_), .Y(mai_mai_n1491_));
  OAI220     m1463(.A0(mai_mai_n1491_), .A1(mai_mai_n1489_), .B0(mai_mai_n1490_), .B1(mai_mai_n448_), .Y(mai_mai_n1492_));
  INV        m1464(.A(mai_mai_n1492_), .Y(mai_mai_n1493_));
  NO2        m1465(.A(mai_mai_n183_), .B(c), .Y(mai_mai_n1494_));
  OAI210     m1466(.A0(mai_mai_n1494_), .A1(mai_mai_n1488_), .B0(mai_mai_n181_), .Y(mai_mai_n1495_));
  AOI220     m1467(.A0(mai_mai_n1495_), .A1(mai_mai_n1087_), .B0(mai_mai_n545_), .B1(mai_mai_n373_), .Y(mai_mai_n1496_));
  AOI210     m1468(.A0(j), .A1(mai_mai_n1378_), .B0(mai_mai_n1457_), .Y(mai_mai_n1497_));
  NO2        m1469(.A(mai_mai_n1417_), .B(f), .Y(mai_mai_n1498_));
  NA2        m1470(.A(mai_mai_n1137_), .B(a), .Y(mai_mai_n1499_));
  OAI220     m1471(.A0(mai_mai_n1499_), .A1(mai_mai_n66_), .B0(mai_mai_n1497_), .B1(mai_mai_n217_), .Y(mai_mai_n1500_));
  AOI210     m1472(.A0(mai_mai_n911_), .A1(mai_mai_n421_), .B0(mai_mai_n104_), .Y(mai_mai_n1501_));
  OR2        m1473(.A(mai_mai_n1501_), .B(mai_mai_n553_), .Y(mai_mai_n1502_));
  NA2        m1474(.A(mai_mai_n1498_), .B(mai_mai_n1357_), .Y(mai_mai_n1503_));
  OAI220     m1475(.A0(mai_mai_n1503_), .A1(mai_mai_n49_), .B0(mai_mai_n1502_), .B1(mai_mai_n176_), .Y(mai_mai_n1504_));
  NA4        m1476(.A(mai_mai_n1108_), .B(mai_mai_n1105_), .C(mai_mai_n225_), .D(mai_mai_n65_), .Y(mai_mai_n1505_));
  NA2        m1477(.A(mai_mai_n1351_), .B(mai_mai_n184_), .Y(mai_mai_n1506_));
  NO2        m1478(.A(mai_mai_n49_), .B(l), .Y(mai_mai_n1507_));
  OAI210     m1479(.A0(mai_mai_n1417_), .A1(mai_mai_n874_), .B0(mai_mai_n492_), .Y(mai_mai_n1508_));
  OAI210     m1480(.A0(mai_mai_n1508_), .A1(mai_mai_n1111_), .B0(mai_mai_n1507_), .Y(mai_mai_n1509_));
  NO2        m1481(.A(mai_mai_n259_), .B(g), .Y(mai_mai_n1510_));
  NO2        m1482(.A(m), .B(i), .Y(mai_mai_n1511_));
  BUFFER     m1483(.A(mai_mai_n1511_), .Y(mai_mai_n1512_));
  AOI220     m1484(.A0(mai_mai_n1512_), .A1(mai_mai_n1380_), .B0(mai_mai_n1086_), .B1(mai_mai_n1510_), .Y(mai_mai_n1513_));
  NA4        m1485(.A(mai_mai_n1513_), .B(mai_mai_n1509_), .C(mai_mai_n1506_), .D(mai_mai_n1505_), .Y(mai_mai_n1514_));
  NO4        m1486(.A(mai_mai_n1514_), .B(mai_mai_n1504_), .C(mai_mai_n1500_), .D(mai_mai_n1496_), .Y(mai_mai_n1515_));
  NA3        m1487(.A(mai_mai_n1515_), .B(mai_mai_n1493_), .C(mai_mai_n1487_), .Y(mai_mai_n1516_));
  NA3        m1488(.A(mai_mai_n971_), .B(mai_mai_n139_), .C(mai_mai_n46_), .Y(mai_mai_n1517_));
  AOI210     m1489(.A0(mai_mai_n150_), .A1(c), .B0(mai_mai_n1517_), .Y(mai_mai_n1518_));
  INV        m1490(.A(mai_mai_n187_), .Y(mai_mai_n1519_));
  NA2        m1491(.A(mai_mai_n1519_), .B(mai_mai_n1458_), .Y(mai_mai_n1520_));
  OR2        m1492(.A(mai_mai_n134_), .B(mai_mai_n1408_), .Y(mai_mai_n1521_));
  NO2        m1493(.A(mai_mai_n69_), .B(c), .Y(mai_mai_n1522_));
  NA2        m1494(.A(mai_mai_n1466_), .B(mai_mai_n1522_), .Y(mai_mai_n1523_));
  NA3        m1495(.A(mai_mai_n1523_), .B(mai_mai_n1521_), .C(mai_mai_n1520_), .Y(mai_mai_n1524_));
  NO2        m1496(.A(mai_mai_n1524_), .B(mai_mai_n1518_), .Y(mai_mai_n1525_));
  AOI210     m1497(.A0(mai_mai_n158_), .A1(mai_mai_n56_), .B0(mai_mai_n1488_), .Y(mai_mai_n1526_));
  NO2        m1498(.A(mai_mai_n1526_), .B(mai_mai_n1462_), .Y(mai_mai_n1527_));
  NOi21      m1499(.An(mai_mai_n1351_), .B(e), .Y(mai_mai_n1528_));
  NO2        m1500(.A(mai_mai_n1528_), .B(mai_mai_n1527_), .Y(mai_mai_n1529_));
  AN2        m1501(.A(mai_mai_n1108_), .B(mai_mai_n1093_), .Y(mai_mai_n1530_));
  NA2        m1502(.A(mai_mai_n1070_), .B(mai_mai_n161_), .Y(mai_mai_n1531_));
  NOi31      m1503(.An(mai_mai_n30_), .B(mai_mai_n1531_), .C(n), .Y(mai_mai_n1532_));
  AOI210     m1504(.A0(mai_mai_n1530_), .A1(mai_mai_n1174_), .B0(mai_mai_n1532_), .Y(mai_mai_n1533_));
  NO2        m1505(.A(mai_mai_n1461_), .B(mai_mai_n66_), .Y(mai_mai_n1534_));
  NA2        m1506(.A(mai_mai_n59_), .B(a), .Y(mai_mai_n1535_));
  NO2        m1507(.A(mai_mai_n1355_), .B(mai_mai_n118_), .Y(mai_mai_n1536_));
  OAI220     m1508(.A0(mai_mai_n1536_), .A1(mai_mai_n1408_), .B0(mai_mai_n1424_), .B1(mai_mai_n1535_), .Y(mai_mai_n1537_));
  NO2        m1509(.A(mai_mai_n1537_), .B(mai_mai_n1534_), .Y(mai_mai_n1538_));
  NA4        m1510(.A(mai_mai_n1538_), .B(mai_mai_n1533_), .C(mai_mai_n1529_), .D(mai_mai_n1525_), .Y(mai_mai_n1539_));
  OR4        m1511(.A(mai_mai_n1539_), .B(mai_mai_n1516_), .C(mai_mai_n1474_), .D(mai_mai_n1428_), .Y(mai04));
  NOi31      m1512(.An(mai_mai_n1414_), .B(mai_mai_n1415_), .C(mai_mai_n1058_), .Y(mai_mai_n1541_));
  NA2        m1513(.A(mai_mai_n1470_), .B(mai_mai_n835_), .Y(mai_mai_n1542_));
  NO4        m1514(.A(mai_mai_n1542_), .B(mai_mai_n1048_), .C(mai_mai_n493_), .D(j), .Y(mai_mai_n1543_));
  OR3        m1515(.A(mai_mai_n1543_), .B(mai_mai_n1541_), .C(mai_mai_n1076_), .Y(mai_mai_n1544_));
  NO2        m1516(.A(mai_mai_n1357_), .B(mai_mai_n89_), .Y(mai_mai_n1545_));
  AOI210     m1517(.A0(mai_mai_n1545_), .A1(mai_mai_n1069_), .B0(mai_mai_n1194_), .Y(mai_mai_n1546_));
  NA2        m1518(.A(mai_mai_n1546_), .B(mai_mai_n1222_), .Y(mai_mai_n1547_));
  NO4        m1519(.A(mai_mai_n1547_), .B(mai_mai_n1544_), .C(mai_mai_n1084_), .D(mai_mai_n1063_), .Y(mai_mai_n1548_));
  NA4        m1520(.A(mai_mai_n1548_), .B(mai_mai_n1139_), .C(mai_mai_n1126_), .D(mai_mai_n1114_), .Y(mai05));
  INV        m1521(.A(mai_mai_n612_), .Y(mai_mai_n1552_));
  INV        m1522(.A(mai_mai_n909_), .Y(mai_mai_n1553_));
  AN2        u0000(.A(b), .B(a), .Y(men_men_n29_));
  NO2        u0001(.A(d), .B(c), .Y(men_men_n30_));
  AN2        u0002(.A(f), .B(e), .Y(men_men_n31_));
  NA3        u0003(.A(men_men_n31_), .B(men_men_n30_), .C(men_men_n29_), .Y(men_men_n32_));
  NOi32      u0004(.An(m), .Bn(l), .C(n), .Y(men_men_n33_));
  NOi32      u0005(.An(i), .Bn(g), .C(h), .Y(men_men_n34_));
  NA2        u0006(.A(men_men_n34_), .B(men_men_n33_), .Y(men_men_n35_));
  AN2        u0007(.A(m), .B(l), .Y(men_men_n36_));
  NOi32      u0008(.An(j), .Bn(g), .C(k), .Y(men_men_n37_));
  NA2        u0009(.A(men_men_n37_), .B(men_men_n36_), .Y(men_men_n38_));
  NO2        u0010(.A(men_men_n38_), .B(n), .Y(men_men_n39_));
  INV        u0011(.A(h), .Y(men_men_n40_));
  NAi21      u0012(.An(j), .B(l), .Y(men_men_n41_));
  NAi32      u0013(.An(n), .Bn(g), .C(m), .Y(men_men_n42_));
  NO3        u0014(.A(men_men_n42_), .B(men_men_n41_), .C(men_men_n40_), .Y(men_men_n43_));
  NAi31      u0015(.An(n), .B(m), .C(l), .Y(men_men_n44_));
  INV        u0016(.A(i), .Y(men_men_n45_));
  AN2        u0017(.A(h), .B(g), .Y(men_men_n46_));
  NA2        u0018(.A(men_men_n46_), .B(men_men_n45_), .Y(men_men_n47_));
  NO2        u0019(.A(men_men_n47_), .B(men_men_n44_), .Y(men_men_n48_));
  NAi21      u0020(.An(n), .B(m), .Y(men_men_n49_));
  NOi32      u0021(.An(k), .Bn(h), .C(l), .Y(men_men_n50_));
  NOi32      u0022(.An(k), .Bn(h), .C(g), .Y(men_men_n51_));
  INV        u0023(.A(men_men_n51_), .Y(men_men_n52_));
  NO2        u0024(.A(men_men_n52_), .B(men_men_n49_), .Y(men_men_n53_));
  NO4        u0025(.A(men_men_n53_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n54_));
  AOI210     u0026(.A0(men_men_n54_), .A1(men_men_n35_), .B0(men_men_n32_), .Y(men_men_n55_));
  INV        u0027(.A(c), .Y(men_men_n56_));
  NA2        u0028(.A(e), .B(b), .Y(men_men_n57_));
  NO2        u0029(.A(men_men_n57_), .B(men_men_n56_), .Y(men_men_n58_));
  INV        u0030(.A(d), .Y(men_men_n59_));
  NA3        u0031(.A(g), .B(men_men_n59_), .C(a), .Y(men_men_n60_));
  NAi21      u0032(.An(i), .B(h), .Y(men_men_n61_));
  NA2        u0033(.A(l), .B(j), .Y(men_men_n62_));
  OAI220     u0034(.A0(men_men_n62_), .A1(men_men_n49_), .B0(men_men_n61_), .B1(men_men_n44_), .Y(men_men_n63_));
  NAi31      u0035(.An(men_men_n60_), .B(men_men_n63_), .C(men_men_n58_), .Y(men_men_n64_));
  NAi41      u0036(.An(e), .B(d), .C(b), .D(a), .Y(men_men_n65_));
  NA2        u0037(.A(g), .B(f), .Y(men_men_n66_));
  NO2        u0038(.A(men_men_n66_), .B(men_men_n65_), .Y(men_men_n67_));
  NAi21      u0039(.An(i), .B(j), .Y(men_men_n68_));
  NAi32      u0040(.An(n), .Bn(k), .C(m), .Y(men_men_n69_));
  NO2        u0041(.A(men_men_n69_), .B(men_men_n68_), .Y(men_men_n70_));
  NAi31      u0042(.An(l), .B(m), .C(k), .Y(men_men_n71_));
  NAi21      u0043(.An(e), .B(h), .Y(men_men_n72_));
  NAi41      u0044(.An(n), .B(d), .C(b), .D(a), .Y(men_men_n73_));
  NA2        u0045(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n74_));
  INV        u0046(.A(m), .Y(men_men_n75_));
  NOi21      u0047(.An(k), .B(l), .Y(men_men_n76_));
  NA2        u0048(.A(men_men_n76_), .B(men_men_n75_), .Y(men_men_n77_));
  AN4        u0049(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n78_));
  NOi31      u0050(.An(h), .B(g), .C(f), .Y(men_men_n79_));
  NA2        u0051(.A(men_men_n79_), .B(men_men_n78_), .Y(men_men_n80_));
  NAi32      u0052(.An(m), .Bn(k), .C(j), .Y(men_men_n81_));
  NOi32      u0053(.An(h), .Bn(g), .C(f), .Y(men_men_n82_));
  NA2        u0054(.A(men_men_n82_), .B(men_men_n78_), .Y(men_men_n83_));
  OA220      u0055(.A0(men_men_n83_), .A1(men_men_n81_), .B0(men_men_n80_), .B1(men_men_n77_), .Y(men_men_n84_));
  NA3        u0056(.A(men_men_n84_), .B(men_men_n74_), .C(men_men_n64_), .Y(men_men_n85_));
  INV        u0057(.A(n), .Y(men_men_n86_));
  NOi32      u0058(.An(e), .Bn(b), .C(d), .Y(men_men_n87_));
  NA2        u0059(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n88_));
  INV        u0060(.A(j), .Y(men_men_n89_));
  AN3        u0061(.A(m), .B(k), .C(i), .Y(men_men_n90_));
  NA3        u0062(.A(men_men_n90_), .B(men_men_n89_), .C(g), .Y(men_men_n91_));
  NO2        u0063(.A(men_men_n91_), .B(f), .Y(men_men_n92_));
  NAi32      u0064(.An(g), .Bn(f), .C(h), .Y(men_men_n93_));
  NAi31      u0065(.An(j), .B(m), .C(l), .Y(men_men_n94_));
  NO2        u0066(.A(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u0067(.A(m), .B(l), .Y(men_men_n96_));
  NAi31      u0068(.An(k), .B(j), .C(g), .Y(men_men_n97_));
  NO3        u0069(.A(men_men_n97_), .B(men_men_n96_), .C(f), .Y(men_men_n98_));
  AN2        u0070(.A(j), .B(g), .Y(men_men_n99_));
  NOi32      u0071(.An(m), .Bn(l), .C(i), .Y(men_men_n100_));
  NOi21      u0072(.An(g), .B(i), .Y(men_men_n101_));
  NOi32      u0073(.An(m), .Bn(j), .C(k), .Y(men_men_n102_));
  AOI220     u0074(.A0(men_men_n102_), .A1(men_men_n101_), .B0(men_men_n100_), .B1(men_men_n99_), .Y(men_men_n103_));
  NO2        u0075(.A(men_men_n98_), .B(men_men_n92_), .Y(men_men_n104_));
  NAi41      u0076(.An(m), .B(n), .C(k), .D(i), .Y(men_men_n105_));
  AN2        u0077(.A(e), .B(b), .Y(men_men_n106_));
  NOi31      u0078(.An(c), .B(h), .C(f), .Y(men_men_n107_));
  NA2        u0079(.A(men_men_n107_), .B(men_men_n106_), .Y(men_men_n108_));
  NO2        u0080(.A(men_men_n108_), .B(men_men_n105_), .Y(men_men_n109_));
  NOi21      u0081(.An(g), .B(f), .Y(men_men_n110_));
  NOi21      u0082(.An(i), .B(h), .Y(men_men_n111_));
  INV        u0083(.A(a), .Y(men_men_n112_));
  NA2        u0084(.A(men_men_n106_), .B(men_men_n112_), .Y(men_men_n113_));
  INV        u0085(.A(l), .Y(men_men_n114_));
  NOi21      u0086(.An(m), .B(n), .Y(men_men_n115_));
  AN2        u0087(.A(k), .B(h), .Y(men_men_n116_));
  INV        u0088(.A(b), .Y(men_men_n117_));
  NA2        u0089(.A(l), .B(j), .Y(men_men_n118_));
  AN2        u0090(.A(k), .B(i), .Y(men_men_n119_));
  NA2        u0091(.A(men_men_n119_), .B(men_men_n118_), .Y(men_men_n120_));
  NA2        u0092(.A(g), .B(e), .Y(men_men_n121_));
  NOi32      u0093(.An(c), .Bn(a), .C(d), .Y(men_men_n122_));
  NA2        u0094(.A(men_men_n122_), .B(men_men_n115_), .Y(men_men_n123_));
  NO4        u0095(.A(men_men_n123_), .B(men_men_n121_), .C(men_men_n120_), .D(men_men_n117_), .Y(men_men_n124_));
  NO2        u0096(.A(men_men_n124_), .B(men_men_n109_), .Y(men_men_n125_));
  OAI210     u0097(.A0(men_men_n104_), .A1(men_men_n88_), .B0(men_men_n125_), .Y(men_men_n126_));
  NOi31      u0098(.An(k), .B(m), .C(j), .Y(men_men_n127_));
  NOi31      u0099(.An(k), .B(m), .C(i), .Y(men_men_n128_));
  NOi32      u0100(.An(f), .Bn(b), .C(e), .Y(men_men_n129_));
  NAi21      u0101(.An(g), .B(h), .Y(men_men_n130_));
  NAi21      u0102(.An(m), .B(n), .Y(men_men_n131_));
  NAi21      u0103(.An(j), .B(k), .Y(men_men_n132_));
  NO3        u0104(.A(men_men_n132_), .B(men_men_n131_), .C(men_men_n130_), .Y(men_men_n133_));
  NAi41      u0105(.An(e), .B(f), .C(d), .D(b), .Y(men_men_n134_));
  NAi31      u0106(.An(j), .B(k), .C(h), .Y(men_men_n135_));
  NO3        u0107(.A(men_men_n135_), .B(men_men_n134_), .C(men_men_n131_), .Y(men_men_n136_));
  AOI210     u0108(.A0(men_men_n133_), .A1(men_men_n129_), .B0(men_men_n136_), .Y(men_men_n137_));
  NO2        u0109(.A(k), .B(j), .Y(men_men_n138_));
  AN2        u0110(.A(k), .B(j), .Y(men_men_n139_));
  NAi21      u0111(.An(c), .B(b), .Y(men_men_n140_));
  NA2        u0112(.A(f), .B(d), .Y(men_men_n141_));
  NA2        u0113(.A(h), .B(c), .Y(men_men_n142_));
  NAi31      u0114(.An(f), .B(e), .C(b), .Y(men_men_n143_));
  NA2        u0115(.A(d), .B(b), .Y(men_men_n144_));
  NAi21      u0116(.An(e), .B(f), .Y(men_men_n145_));
  NO2        u0117(.A(men_men_n145_), .B(men_men_n144_), .Y(men_men_n146_));
  NA2        u0118(.A(b), .B(a), .Y(men_men_n147_));
  NAi21      u0119(.An(e), .B(g), .Y(men_men_n148_));
  NAi21      u0120(.An(c), .B(d), .Y(men_men_n149_));
  NAi31      u0121(.An(l), .B(k), .C(h), .Y(men_men_n150_));
  NO2        u0122(.A(men_men_n131_), .B(men_men_n150_), .Y(men_men_n151_));
  NA2        u0123(.A(men_men_n151_), .B(men_men_n146_), .Y(men_men_n152_));
  NA2        u0124(.A(men_men_n152_), .B(men_men_n137_), .Y(men_men_n153_));
  NAi31      u0125(.An(e), .B(f), .C(b), .Y(men_men_n154_));
  NOi21      u0126(.An(g), .B(d), .Y(men_men_n155_));
  NO2        u0127(.A(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  NOi21      u0128(.An(h), .B(i), .Y(men_men_n157_));
  NOi21      u0129(.An(k), .B(m), .Y(men_men_n158_));
  NA3        u0130(.A(men_men_n158_), .B(men_men_n157_), .C(n), .Y(men_men_n159_));
  NOi21      u0131(.An(men_men_n156_), .B(men_men_n159_), .Y(men_men_n160_));
  NOi21      u0132(.An(h), .B(g), .Y(men_men_n161_));
  NO2        u0133(.A(men_men_n141_), .B(men_men_n140_), .Y(men_men_n162_));
  NA2        u0134(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  NAi31      u0135(.An(l), .B(j), .C(h), .Y(men_men_n164_));
  NO2        u0136(.A(men_men_n164_), .B(men_men_n49_), .Y(men_men_n165_));
  NA2        u0137(.A(men_men_n165_), .B(men_men_n67_), .Y(men_men_n166_));
  NOi32      u0138(.An(n), .Bn(k), .C(m), .Y(men_men_n167_));
  NA2        u0139(.A(l), .B(i), .Y(men_men_n168_));
  NA2        u0140(.A(men_men_n168_), .B(men_men_n167_), .Y(men_men_n169_));
  OAI210     u0141(.A0(men_men_n169_), .A1(men_men_n163_), .B0(men_men_n166_), .Y(men_men_n170_));
  NAi31      u0142(.An(d), .B(f), .C(c), .Y(men_men_n171_));
  NAi31      u0143(.An(e), .B(f), .C(c), .Y(men_men_n172_));
  NA2        u0144(.A(men_men_n172_), .B(men_men_n171_), .Y(men_men_n173_));
  NA2        u0145(.A(j), .B(h), .Y(men_men_n174_));
  OR3        u0146(.A(n), .B(m), .C(k), .Y(men_men_n175_));
  NO2        u0147(.A(men_men_n175_), .B(men_men_n174_), .Y(men_men_n176_));
  NAi32      u0148(.An(m), .Bn(k), .C(n), .Y(men_men_n177_));
  NO2        u0149(.A(men_men_n177_), .B(men_men_n174_), .Y(men_men_n178_));
  AOI220     u0150(.A0(men_men_n178_), .A1(men_men_n156_), .B0(men_men_n176_), .B1(men_men_n173_), .Y(men_men_n179_));
  NO2        u0151(.A(n), .B(m), .Y(men_men_n180_));
  NA2        u0152(.A(men_men_n180_), .B(men_men_n50_), .Y(men_men_n181_));
  NAi21      u0153(.An(f), .B(e), .Y(men_men_n182_));
  NA2        u0154(.A(d), .B(c), .Y(men_men_n183_));
  NO2        u0155(.A(men_men_n183_), .B(men_men_n182_), .Y(men_men_n184_));
  NOi21      u0156(.An(men_men_n184_), .B(men_men_n181_), .Y(men_men_n185_));
  NAi21      u0157(.An(d), .B(c), .Y(men_men_n186_));
  NAi31      u0158(.An(m), .B(n), .C(b), .Y(men_men_n187_));
  NA2        u0159(.A(k), .B(i), .Y(men_men_n188_));
  NAi21      u0160(.An(h), .B(f), .Y(men_men_n189_));
  NO2        u0161(.A(men_men_n189_), .B(men_men_n188_), .Y(men_men_n190_));
  NO2        u0162(.A(men_men_n187_), .B(men_men_n149_), .Y(men_men_n191_));
  NA2        u0163(.A(men_men_n191_), .B(men_men_n190_), .Y(men_men_n192_));
  NOi32      u0164(.An(f), .Bn(c), .C(d), .Y(men_men_n193_));
  NOi32      u0165(.An(f), .Bn(c), .C(e), .Y(men_men_n194_));
  NO2        u0166(.A(men_men_n194_), .B(men_men_n193_), .Y(men_men_n195_));
  NO3        u0167(.A(n), .B(m), .C(j), .Y(men_men_n196_));
  NA2        u0168(.A(men_men_n196_), .B(men_men_n116_), .Y(men_men_n197_));
  AO210      u0169(.A0(men_men_n197_), .A1(men_men_n181_), .B0(men_men_n195_), .Y(men_men_n198_));
  NAi41      u0170(.An(men_men_n185_), .B(men_men_n198_), .C(men_men_n192_), .D(men_men_n179_), .Y(men_men_n199_));
  OR4        u0171(.A(men_men_n199_), .B(men_men_n170_), .C(men_men_n160_), .D(men_men_n153_), .Y(men_men_n200_));
  NO4        u0172(.A(men_men_n200_), .B(men_men_n126_), .C(men_men_n85_), .D(men_men_n55_), .Y(men_men_n201_));
  NA3        u0173(.A(m), .B(men_men_n114_), .C(j), .Y(men_men_n202_));
  NAi31      u0174(.An(n), .B(h), .C(g), .Y(men_men_n203_));
  NO2        u0175(.A(men_men_n203_), .B(men_men_n202_), .Y(men_men_n204_));
  NOi32      u0176(.An(m), .Bn(k), .C(l), .Y(men_men_n205_));
  NA3        u0177(.A(men_men_n205_), .B(men_men_n89_), .C(g), .Y(men_men_n206_));
  NO2        u0178(.A(men_men_n206_), .B(n), .Y(men_men_n207_));
  NOi21      u0179(.An(k), .B(j), .Y(men_men_n208_));
  NA4        u0180(.A(men_men_n208_), .B(men_men_n115_), .C(i), .D(g), .Y(men_men_n209_));
  AN2        u0181(.A(i), .B(g), .Y(men_men_n210_));
  NA3        u0182(.A(men_men_n76_), .B(men_men_n210_), .C(men_men_n115_), .Y(men_men_n211_));
  NA2        u0183(.A(men_men_n211_), .B(men_men_n209_), .Y(men_men_n212_));
  NO3        u0184(.A(men_men_n212_), .B(men_men_n207_), .C(men_men_n204_), .Y(men_men_n213_));
  NAi41      u0185(.An(d), .B(n), .C(e), .D(b), .Y(men_men_n214_));
  INV        u0186(.A(men_men_n214_), .Y(men_men_n215_));
  INV        u0187(.A(f), .Y(men_men_n216_));
  INV        u0188(.A(g), .Y(men_men_n217_));
  NOi31      u0189(.An(i), .B(j), .C(h), .Y(men_men_n218_));
  NOi21      u0190(.An(l), .B(m), .Y(men_men_n219_));
  NA2        u0191(.A(men_men_n219_), .B(men_men_n218_), .Y(men_men_n220_));
  NO3        u0192(.A(men_men_n220_), .B(men_men_n217_), .C(men_men_n216_), .Y(men_men_n221_));
  NA2        u0193(.A(men_men_n221_), .B(men_men_n215_), .Y(men_men_n222_));
  OAI210     u0194(.A0(men_men_n213_), .A1(men_men_n32_), .B0(men_men_n222_), .Y(men_men_n223_));
  NOi21      u0195(.An(n), .B(m), .Y(men_men_n224_));
  NOi32      u0196(.An(l), .Bn(i), .C(j), .Y(men_men_n225_));
  NA2        u0197(.A(men_men_n225_), .B(men_men_n224_), .Y(men_men_n226_));
  OA220      u0198(.A0(men_men_n226_), .A1(men_men_n108_), .B0(men_men_n81_), .B1(men_men_n80_), .Y(men_men_n227_));
  NAi21      u0199(.An(j), .B(h), .Y(men_men_n228_));
  XN2        u0200(.A(i), .B(h), .Y(men_men_n229_));
  NA2        u0201(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  NOi31      u0202(.An(k), .B(n), .C(m), .Y(men_men_n231_));
  NOi31      u0203(.An(men_men_n231_), .B(men_men_n183_), .C(men_men_n182_), .Y(men_men_n232_));
  NA2        u0204(.A(men_men_n232_), .B(men_men_n230_), .Y(men_men_n233_));
  NAi31      u0205(.An(f), .B(e), .C(c), .Y(men_men_n234_));
  NO4        u0206(.A(men_men_n234_), .B(men_men_n175_), .C(men_men_n174_), .D(men_men_n59_), .Y(men_men_n235_));
  NA4        u0207(.A(n), .B(e), .C(c), .D(b), .Y(men_men_n236_));
  NAi32      u0208(.An(m), .Bn(i), .C(k), .Y(men_men_n237_));
  NO3        u0209(.A(men_men_n237_), .B(men_men_n93_), .C(men_men_n236_), .Y(men_men_n238_));
  INV        u0210(.A(k), .Y(men_men_n239_));
  NO2        u0211(.A(men_men_n238_), .B(men_men_n235_), .Y(men_men_n240_));
  NAi21      u0212(.An(n), .B(a), .Y(men_men_n241_));
  NO2        u0213(.A(men_men_n241_), .B(men_men_n144_), .Y(men_men_n242_));
  NAi41      u0214(.An(g), .B(m), .C(k), .D(h), .Y(men_men_n243_));
  NO2        u0215(.A(men_men_n243_), .B(e), .Y(men_men_n244_));
  NO3        u0216(.A(men_men_n145_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n245_));
  OAI210     u0217(.A0(men_men_n245_), .A1(men_men_n244_), .B0(men_men_n242_), .Y(men_men_n246_));
  AN4        u0218(.A(men_men_n246_), .B(men_men_n240_), .C(men_men_n233_), .D(men_men_n227_), .Y(men_men_n247_));
  OR2        u0219(.A(h), .B(g), .Y(men_men_n248_));
  NO2        u0220(.A(men_men_n248_), .B(men_men_n105_), .Y(men_men_n249_));
  NA2        u0221(.A(men_men_n249_), .B(men_men_n129_), .Y(men_men_n250_));
  NAi31      u0222(.An(e), .B(d), .C(b), .Y(men_men_n251_));
  NA2        u0223(.A(men_men_n158_), .B(men_men_n111_), .Y(men_men_n252_));
  NO2        u0224(.A(n), .B(a), .Y(men_men_n253_));
  NAi31      u0225(.An(men_men_n243_), .B(men_men_n253_), .C(men_men_n106_), .Y(men_men_n254_));
  NAi21      u0226(.An(h), .B(i), .Y(men_men_n255_));
  NA2        u0227(.A(men_men_n180_), .B(k), .Y(men_men_n256_));
  NO2        u0228(.A(men_men_n256_), .B(men_men_n255_), .Y(men_men_n257_));
  NA2        u0229(.A(men_men_n257_), .B(men_men_n193_), .Y(men_men_n258_));
  NA3        u0230(.A(men_men_n258_), .B(men_men_n254_), .C(men_men_n250_), .Y(men_men_n259_));
  NOi21      u0231(.An(g), .B(e), .Y(men_men_n260_));
  NO2        u0232(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n261_));
  NOi32      u0233(.An(l), .Bn(j), .C(i), .Y(men_men_n262_));
  AOI210     u0234(.A0(men_men_n76_), .A1(men_men_n89_), .B0(men_men_n262_), .Y(men_men_n263_));
  NAi21      u0235(.An(f), .B(g), .Y(men_men_n264_));
  NO2        u0236(.A(men_men_n264_), .B(men_men_n65_), .Y(men_men_n265_));
  NO2        u0237(.A(men_men_n69_), .B(men_men_n118_), .Y(men_men_n266_));
  NO3        u0238(.A(men_men_n132_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n267_));
  NOi31      u0239(.An(men_men_n247_), .B(men_men_n259_), .C(men_men_n223_), .Y(men_men_n268_));
  NO4        u0240(.A(men_men_n204_), .B(men_men_n48_), .C(men_men_n43_), .D(men_men_n39_), .Y(men_men_n269_));
  NO2        u0241(.A(men_men_n269_), .B(men_men_n113_), .Y(men_men_n270_));
  NA3        u0242(.A(men_men_n59_), .B(c), .C(b), .Y(men_men_n271_));
  NAi21      u0243(.An(h), .B(g), .Y(men_men_n272_));
  NO2        u0244(.A(men_men_n252_), .B(men_men_n264_), .Y(men_men_n273_));
  NAi31      u0245(.An(g), .B(k), .C(h), .Y(men_men_n274_));
  NO3        u0246(.A(men_men_n131_), .B(men_men_n274_), .C(l), .Y(men_men_n275_));
  NAi31      u0247(.An(e), .B(d), .C(a), .Y(men_men_n276_));
  NA2        u0248(.A(men_men_n275_), .B(men_men_n129_), .Y(men_men_n277_));
  INV        u0249(.A(men_men_n277_), .Y(men_men_n278_));
  NA4        u0250(.A(men_men_n158_), .B(men_men_n82_), .C(men_men_n78_), .D(men_men_n118_), .Y(men_men_n279_));
  NA3        u0251(.A(men_men_n158_), .B(men_men_n157_), .C(men_men_n86_), .Y(men_men_n280_));
  NO2        u0252(.A(men_men_n280_), .B(men_men_n195_), .Y(men_men_n281_));
  NOi21      u0253(.An(men_men_n279_), .B(men_men_n281_), .Y(men_men_n282_));
  NA3        u0254(.A(e), .B(c), .C(b), .Y(men_men_n283_));
  NO2        u0255(.A(men_men_n60_), .B(men_men_n283_), .Y(men_men_n284_));
  NAi32      u0256(.An(k), .Bn(i), .C(j), .Y(men_men_n285_));
  NAi31      u0257(.An(h), .B(l), .C(i), .Y(men_men_n286_));
  NA3        u0258(.A(men_men_n286_), .B(men_men_n285_), .C(men_men_n164_), .Y(men_men_n287_));
  NOi21      u0259(.An(men_men_n287_), .B(men_men_n49_), .Y(men_men_n288_));
  OAI210     u0260(.A0(men_men_n265_), .A1(men_men_n284_), .B0(men_men_n288_), .Y(men_men_n289_));
  NAi21      u0261(.An(l), .B(k), .Y(men_men_n290_));
  NO2        u0262(.A(men_men_n290_), .B(men_men_n49_), .Y(men_men_n291_));
  NOi21      u0263(.An(l), .B(j), .Y(men_men_n292_));
  NA2        u0264(.A(men_men_n161_), .B(men_men_n292_), .Y(men_men_n293_));
  NA3        u0265(.A(men_men_n119_), .B(men_men_n118_), .C(g), .Y(men_men_n294_));
  OR3        u0266(.A(men_men_n73_), .B(men_men_n75_), .C(e), .Y(men_men_n295_));
  AOI210     u0267(.A0(men_men_n294_), .A1(men_men_n293_), .B0(men_men_n295_), .Y(men_men_n296_));
  INV        u0268(.A(men_men_n296_), .Y(men_men_n297_));
  NAi32      u0269(.An(j), .Bn(h), .C(i), .Y(men_men_n298_));
  NAi21      u0270(.An(m), .B(l), .Y(men_men_n299_));
  NO3        u0271(.A(men_men_n299_), .B(men_men_n298_), .C(men_men_n86_), .Y(men_men_n300_));
  NA2        u0272(.A(h), .B(g), .Y(men_men_n301_));
  NA2        u0273(.A(men_men_n300_), .B(men_men_n162_), .Y(men_men_n302_));
  NA4        u0274(.A(men_men_n302_), .B(men_men_n297_), .C(men_men_n289_), .D(men_men_n282_), .Y(men_men_n303_));
  NO2        u0275(.A(men_men_n143_), .B(d), .Y(men_men_n304_));
  NA2        u0276(.A(men_men_n304_), .B(men_men_n53_), .Y(men_men_n305_));
  NO2        u0277(.A(men_men_n108_), .B(men_men_n105_), .Y(men_men_n306_));
  NAi32      u0278(.An(n), .Bn(m), .C(l), .Y(men_men_n307_));
  NO2        u0279(.A(men_men_n307_), .B(men_men_n298_), .Y(men_men_n308_));
  NA2        u0280(.A(men_men_n308_), .B(men_men_n184_), .Y(men_men_n309_));
  NO2        u0281(.A(men_men_n123_), .B(men_men_n117_), .Y(men_men_n310_));
  NAi31      u0282(.An(k), .B(l), .C(j), .Y(men_men_n311_));
  OAI210     u0283(.A0(men_men_n290_), .A1(j), .B0(men_men_n311_), .Y(men_men_n312_));
  NOi21      u0284(.An(men_men_n312_), .B(men_men_n121_), .Y(men_men_n313_));
  NA2        u0285(.A(men_men_n313_), .B(men_men_n310_), .Y(men_men_n314_));
  NA3        u0286(.A(men_men_n314_), .B(men_men_n309_), .C(men_men_n305_), .Y(men_men_n315_));
  NO4        u0287(.A(men_men_n315_), .B(men_men_n303_), .C(men_men_n278_), .D(men_men_n270_), .Y(men_men_n316_));
  NA2        u0288(.A(men_men_n257_), .B(men_men_n194_), .Y(men_men_n317_));
  NAi21      u0289(.An(m), .B(k), .Y(men_men_n318_));
  NO2        u0290(.A(men_men_n229_), .B(men_men_n318_), .Y(men_men_n319_));
  NAi41      u0291(.An(d), .B(n), .C(c), .D(b), .Y(men_men_n320_));
  NO2        u0292(.A(men_men_n320_), .B(men_men_n148_), .Y(men_men_n321_));
  NA2        u0293(.A(men_men_n321_), .B(men_men_n319_), .Y(men_men_n322_));
  NAi31      u0294(.An(i), .B(l), .C(h), .Y(men_men_n323_));
  NO4        u0295(.A(men_men_n323_), .B(men_men_n148_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n324_));
  NA2        u0296(.A(e), .B(c), .Y(men_men_n325_));
  NO3        u0297(.A(men_men_n325_), .B(n), .C(d), .Y(men_men_n326_));
  NOi21      u0298(.An(f), .B(h), .Y(men_men_n327_));
  NA2        u0299(.A(men_men_n327_), .B(men_men_n119_), .Y(men_men_n328_));
  NO2        u0300(.A(men_men_n328_), .B(men_men_n217_), .Y(men_men_n329_));
  NAi31      u0301(.An(d), .B(e), .C(b), .Y(men_men_n330_));
  NO2        u0302(.A(men_men_n131_), .B(men_men_n330_), .Y(men_men_n331_));
  NA2        u0303(.A(men_men_n331_), .B(men_men_n329_), .Y(men_men_n332_));
  NAi41      u0304(.An(men_men_n324_), .B(men_men_n332_), .C(men_men_n322_), .D(men_men_n317_), .Y(men_men_n333_));
  NO4        u0305(.A(men_men_n320_), .B(men_men_n81_), .C(men_men_n72_), .D(men_men_n217_), .Y(men_men_n334_));
  NA2        u0306(.A(men_men_n253_), .B(men_men_n106_), .Y(men_men_n335_));
  OR2        u0307(.A(men_men_n335_), .B(men_men_n206_), .Y(men_men_n336_));
  NOi31      u0308(.An(l), .B(n), .C(m), .Y(men_men_n337_));
  NA2        u0309(.A(men_men_n337_), .B(men_men_n218_), .Y(men_men_n338_));
  NO2        u0310(.A(men_men_n338_), .B(men_men_n195_), .Y(men_men_n339_));
  NAi32      u0311(.An(men_men_n339_), .Bn(men_men_n334_), .C(men_men_n336_), .Y(men_men_n340_));
  NAi32      u0312(.An(m), .Bn(j), .C(k), .Y(men_men_n341_));
  NAi41      u0313(.An(c), .B(n), .C(d), .D(b), .Y(men_men_n342_));
  OAI210     u0314(.A0(men_men_n214_), .A1(men_men_n341_), .B0(men_men_n342_), .Y(men_men_n343_));
  NOi31      u0315(.An(j), .B(m), .C(k), .Y(men_men_n344_));
  NO2        u0316(.A(men_men_n127_), .B(men_men_n344_), .Y(men_men_n345_));
  AN3        u0317(.A(h), .B(g), .C(f), .Y(men_men_n346_));
  NAi31      u0318(.An(men_men_n345_), .B(men_men_n346_), .C(men_men_n343_), .Y(men_men_n347_));
  NOi32      u0319(.An(m), .Bn(j), .C(l), .Y(men_men_n348_));
  NO2        u0320(.A(men_men_n348_), .B(men_men_n100_), .Y(men_men_n349_));
  NAi32      u0321(.An(men_men_n349_), .Bn(men_men_n203_), .C(men_men_n304_), .Y(men_men_n350_));
  NO2        u0322(.A(men_men_n299_), .B(men_men_n298_), .Y(men_men_n351_));
  NO2        u0323(.A(men_men_n220_), .B(g), .Y(men_men_n352_));
  NO2        u0324(.A(men_men_n154_), .B(men_men_n86_), .Y(men_men_n353_));
  NA2        u0325(.A(men_men_n353_), .B(men_men_n352_), .Y(men_men_n354_));
  NA2        u0326(.A(men_men_n237_), .B(men_men_n81_), .Y(men_men_n355_));
  NA3        u0327(.A(men_men_n355_), .B(men_men_n346_), .C(men_men_n215_), .Y(men_men_n356_));
  NA4        u0328(.A(men_men_n356_), .B(men_men_n354_), .C(men_men_n350_), .D(men_men_n347_), .Y(men_men_n357_));
  NA3        u0329(.A(h), .B(g), .C(f), .Y(men_men_n358_));
  NO2        u0330(.A(men_men_n358_), .B(men_men_n77_), .Y(men_men_n359_));
  NA2        u0331(.A(men_men_n342_), .B(men_men_n214_), .Y(men_men_n360_));
  NA2        u0332(.A(men_men_n161_), .B(e), .Y(men_men_n361_));
  NO2        u0333(.A(men_men_n361_), .B(men_men_n41_), .Y(men_men_n362_));
  AOI220     u0334(.A0(men_men_n362_), .A1(men_men_n310_), .B0(men_men_n360_), .B1(men_men_n359_), .Y(men_men_n363_));
  NOi32      u0335(.An(j), .Bn(g), .C(i), .Y(men_men_n364_));
  NA3        u0336(.A(men_men_n364_), .B(men_men_n290_), .C(men_men_n115_), .Y(men_men_n365_));
  AO210      u0337(.A0(men_men_n113_), .A1(men_men_n32_), .B0(men_men_n365_), .Y(men_men_n366_));
  NOi32      u0338(.An(e), .Bn(b), .C(a), .Y(men_men_n367_));
  AN2        u0339(.A(l), .B(j), .Y(men_men_n368_));
  NO2        u0340(.A(men_men_n318_), .B(men_men_n368_), .Y(men_men_n369_));
  NO3        u0341(.A(men_men_n320_), .B(men_men_n72_), .C(men_men_n217_), .Y(men_men_n370_));
  NA3        u0342(.A(men_men_n211_), .B(men_men_n209_), .C(men_men_n35_), .Y(men_men_n371_));
  AOI220     u0343(.A0(men_men_n371_), .A1(men_men_n367_), .B0(men_men_n370_), .B1(men_men_n369_), .Y(men_men_n372_));
  NO2        u0344(.A(men_men_n330_), .B(n), .Y(men_men_n373_));
  NA2        u0345(.A(men_men_n210_), .B(k), .Y(men_men_n374_));
  NA3        u0346(.A(m), .B(men_men_n114_), .C(men_men_n216_), .Y(men_men_n375_));
  NA4        u0347(.A(men_men_n205_), .B(men_men_n89_), .C(g), .D(men_men_n216_), .Y(men_men_n376_));
  OAI210     u0348(.A0(men_men_n375_), .A1(men_men_n374_), .B0(men_men_n376_), .Y(men_men_n377_));
  NAi41      u0349(.An(d), .B(e), .C(c), .D(a), .Y(men_men_n378_));
  NA2        u0350(.A(men_men_n51_), .B(men_men_n115_), .Y(men_men_n379_));
  NO2        u0351(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n380_));
  AOI220     u0352(.A0(men_men_n380_), .A1(b), .B0(men_men_n377_), .B1(men_men_n373_), .Y(men_men_n381_));
  NA4        u0353(.A(men_men_n381_), .B(men_men_n372_), .C(men_men_n366_), .D(men_men_n363_), .Y(men_men_n382_));
  NO4        u0354(.A(men_men_n382_), .B(men_men_n357_), .C(men_men_n340_), .D(men_men_n333_), .Y(men_men_n383_));
  NA4        u0355(.A(men_men_n383_), .B(men_men_n316_), .C(men_men_n268_), .D(men_men_n201_), .Y(men10));
  NA3        u0356(.A(m), .B(k), .C(i), .Y(men_men_n385_));
  NO3        u0357(.A(men_men_n385_), .B(j), .C(men_men_n217_), .Y(men_men_n386_));
  NOi21      u0358(.An(e), .B(f), .Y(men_men_n387_));
  NO4        u0359(.A(men_men_n149_), .B(men_men_n387_), .C(n), .D(men_men_n112_), .Y(men_men_n388_));
  NAi31      u0360(.An(b), .B(f), .C(c), .Y(men_men_n389_));
  INV        u0361(.A(men_men_n389_), .Y(men_men_n390_));
  NOi32      u0362(.An(k), .Bn(h), .C(j), .Y(men_men_n391_));
  NA2        u0363(.A(men_men_n391_), .B(men_men_n224_), .Y(men_men_n392_));
  NA2        u0364(.A(men_men_n159_), .B(men_men_n392_), .Y(men_men_n393_));
  AOI220     u0365(.A0(men_men_n393_), .A1(men_men_n390_), .B0(men_men_n388_), .B1(men_men_n386_), .Y(men_men_n394_));
  AN2        u0366(.A(j), .B(h), .Y(men_men_n395_));
  NO3        u0367(.A(n), .B(m), .C(k), .Y(men_men_n396_));
  NA2        u0368(.A(men_men_n396_), .B(men_men_n395_), .Y(men_men_n397_));
  NO3        u0369(.A(men_men_n397_), .B(men_men_n149_), .C(men_men_n216_), .Y(men_men_n398_));
  OR2        u0370(.A(m), .B(k), .Y(men_men_n399_));
  NO2        u0371(.A(men_men_n174_), .B(men_men_n399_), .Y(men_men_n400_));
  NA4        u0372(.A(n), .B(f), .C(c), .D(men_men_n117_), .Y(men_men_n401_));
  NOi21      u0373(.An(men_men_n400_), .B(men_men_n401_), .Y(men_men_n402_));
  NOi32      u0374(.An(d), .Bn(a), .C(c), .Y(men_men_n403_));
  NA2        u0375(.A(men_men_n403_), .B(men_men_n182_), .Y(men_men_n404_));
  NAi21      u0376(.An(i), .B(g), .Y(men_men_n405_));
  NAi31      u0377(.An(k), .B(m), .C(j), .Y(men_men_n406_));
  NO2        u0378(.A(men_men_n402_), .B(men_men_n398_), .Y(men_men_n407_));
  NO2        u0379(.A(men_men_n401_), .B(men_men_n299_), .Y(men_men_n408_));
  NOi32      u0380(.An(f), .Bn(d), .C(c), .Y(men_men_n409_));
  AOI220     u0381(.A0(men_men_n409_), .A1(men_men_n308_), .B0(men_men_n408_), .B1(men_men_n218_), .Y(men_men_n410_));
  NA3        u0382(.A(men_men_n410_), .B(men_men_n407_), .C(men_men_n394_), .Y(men_men_n411_));
  NO2        u0383(.A(men_men_n59_), .B(men_men_n117_), .Y(men_men_n412_));
  NA2        u0384(.A(men_men_n253_), .B(men_men_n412_), .Y(men_men_n413_));
  INV        u0385(.A(e), .Y(men_men_n414_));
  NA2        u0386(.A(men_men_n46_), .B(e), .Y(men_men_n415_));
  OAI220     u0387(.A0(men_men_n415_), .A1(men_men_n202_), .B0(men_men_n206_), .B1(men_men_n414_), .Y(men_men_n416_));
  AN2        u0388(.A(g), .B(e), .Y(men_men_n417_));
  NA3        u0389(.A(men_men_n417_), .B(men_men_n205_), .C(i), .Y(men_men_n418_));
  OAI210     u0390(.A0(men_men_n91_), .A1(men_men_n414_), .B0(men_men_n418_), .Y(men_men_n419_));
  NO2        u0391(.A(men_men_n103_), .B(men_men_n414_), .Y(men_men_n420_));
  NO3        u0392(.A(men_men_n420_), .B(men_men_n419_), .C(men_men_n416_), .Y(men_men_n421_));
  NOi32      u0393(.An(h), .Bn(e), .C(g), .Y(men_men_n422_));
  NA3        u0394(.A(men_men_n422_), .B(men_men_n292_), .C(m), .Y(men_men_n423_));
  NOi21      u0395(.An(g), .B(h), .Y(men_men_n424_));
  AN3        u0396(.A(m), .B(l), .C(i), .Y(men_men_n425_));
  NA3        u0397(.A(men_men_n425_), .B(men_men_n424_), .C(e), .Y(men_men_n426_));
  AN3        u0398(.A(h), .B(g), .C(e), .Y(men_men_n427_));
  NA2        u0399(.A(men_men_n427_), .B(men_men_n100_), .Y(men_men_n428_));
  AN3        u0400(.A(men_men_n428_), .B(men_men_n426_), .C(men_men_n423_), .Y(men_men_n429_));
  AOI210     u0401(.A0(men_men_n429_), .A1(men_men_n421_), .B0(men_men_n413_), .Y(men_men_n430_));
  NA3        u0402(.A(men_men_n37_), .B(men_men_n36_), .C(e), .Y(men_men_n431_));
  NO2        u0403(.A(men_men_n431_), .B(men_men_n413_), .Y(men_men_n432_));
  NA3        u0404(.A(men_men_n403_), .B(men_men_n182_), .C(men_men_n86_), .Y(men_men_n433_));
  NAi31      u0405(.An(b), .B(c), .C(a), .Y(men_men_n434_));
  NO2        u0406(.A(men_men_n434_), .B(n), .Y(men_men_n435_));
  NA2        u0407(.A(men_men_n51_), .B(m), .Y(men_men_n436_));
  NO2        u0408(.A(men_men_n436_), .B(men_men_n145_), .Y(men_men_n437_));
  NA2        u0409(.A(men_men_n437_), .B(men_men_n435_), .Y(men_men_n438_));
  INV        u0410(.A(men_men_n438_), .Y(men_men_n439_));
  NO4        u0411(.A(men_men_n439_), .B(men_men_n432_), .C(men_men_n430_), .D(men_men_n411_), .Y(men_men_n440_));
  NA2        u0412(.A(i), .B(g), .Y(men_men_n441_));
  NO3        u0413(.A(men_men_n276_), .B(men_men_n441_), .C(c), .Y(men_men_n442_));
  NOi21      u0414(.An(a), .B(n), .Y(men_men_n443_));
  NOi21      u0415(.An(d), .B(c), .Y(men_men_n444_));
  NA2        u0416(.A(men_men_n444_), .B(men_men_n443_), .Y(men_men_n445_));
  NA3        u0417(.A(i), .B(g), .C(f), .Y(men_men_n446_));
  OR2        u0418(.A(men_men_n446_), .B(men_men_n71_), .Y(men_men_n447_));
  NA2        u0419(.A(men_men_n442_), .B(men_men_n291_), .Y(men_men_n448_));
  OR2        u0420(.A(n), .B(m), .Y(men_men_n449_));
  NO2        u0421(.A(men_men_n449_), .B(men_men_n150_), .Y(men_men_n450_));
  NO2        u0422(.A(men_men_n183_), .B(men_men_n145_), .Y(men_men_n451_));
  OAI210     u0423(.A0(men_men_n450_), .A1(men_men_n176_), .B0(men_men_n451_), .Y(men_men_n452_));
  INV        u0424(.A(men_men_n379_), .Y(men_men_n453_));
  NA3        u0425(.A(men_men_n453_), .B(men_men_n367_), .C(d), .Y(men_men_n454_));
  NO2        u0426(.A(men_men_n434_), .B(men_men_n49_), .Y(men_men_n455_));
  NAi21      u0427(.An(k), .B(j), .Y(men_men_n456_));
  NAi21      u0428(.An(e), .B(d), .Y(men_men_n457_));
  INV        u0429(.A(men_men_n457_), .Y(men_men_n458_));
  NO2        u0430(.A(men_men_n256_), .B(men_men_n216_), .Y(men_men_n459_));
  NA3        u0431(.A(men_men_n459_), .B(men_men_n458_), .C(men_men_n230_), .Y(men_men_n460_));
  NA3        u0432(.A(men_men_n460_), .B(men_men_n454_), .C(men_men_n452_), .Y(men_men_n461_));
  NO2        u0433(.A(men_men_n338_), .B(men_men_n216_), .Y(men_men_n462_));
  NA2        u0434(.A(men_men_n462_), .B(men_men_n458_), .Y(men_men_n463_));
  NOi31      u0435(.An(n), .B(m), .C(k), .Y(men_men_n464_));
  AOI220     u0436(.A0(men_men_n464_), .A1(men_men_n395_), .B0(men_men_n224_), .B1(men_men_n50_), .Y(men_men_n465_));
  NAi31      u0437(.An(g), .B(f), .C(c), .Y(men_men_n466_));
  OR3        u0438(.A(men_men_n466_), .B(men_men_n465_), .C(e), .Y(men_men_n467_));
  NA3        u0439(.A(men_men_n467_), .B(men_men_n463_), .C(men_men_n309_), .Y(men_men_n468_));
  NOi31      u0440(.An(men_men_n448_), .B(men_men_n468_), .C(men_men_n461_), .Y(men_men_n469_));
  NOi32      u0441(.An(c), .Bn(a), .C(b), .Y(men_men_n470_));
  NA2        u0442(.A(men_men_n470_), .B(men_men_n115_), .Y(men_men_n471_));
  INV        u0443(.A(men_men_n274_), .Y(men_men_n472_));
  AN2        u0444(.A(e), .B(d), .Y(men_men_n473_));
  NA2        u0445(.A(men_men_n473_), .B(men_men_n472_), .Y(men_men_n474_));
  INV        u0446(.A(men_men_n145_), .Y(men_men_n475_));
  NO2        u0447(.A(men_men_n130_), .B(men_men_n41_), .Y(men_men_n476_));
  NO2        u0448(.A(men_men_n66_), .B(e), .Y(men_men_n477_));
  NOi31      u0449(.An(j), .B(k), .C(i), .Y(men_men_n478_));
  NOi21      u0450(.An(men_men_n164_), .B(men_men_n478_), .Y(men_men_n479_));
  NA4        u0451(.A(men_men_n323_), .B(men_men_n479_), .C(men_men_n263_), .D(men_men_n120_), .Y(men_men_n480_));
  AOI220     u0452(.A0(men_men_n480_), .A1(men_men_n477_), .B0(men_men_n476_), .B1(men_men_n475_), .Y(men_men_n481_));
  AOI210     u0453(.A0(men_men_n481_), .A1(men_men_n474_), .B0(men_men_n471_), .Y(men_men_n482_));
  NO2        u0454(.A(men_men_n212_), .B(men_men_n207_), .Y(men_men_n483_));
  NOi21      u0455(.An(a), .B(b), .Y(men_men_n484_));
  NA3        u0456(.A(e), .B(d), .C(c), .Y(men_men_n485_));
  NAi21      u0457(.An(men_men_n485_), .B(men_men_n484_), .Y(men_men_n486_));
  NO2        u0458(.A(men_men_n433_), .B(men_men_n206_), .Y(men_men_n487_));
  NOi21      u0459(.An(men_men_n486_), .B(men_men_n487_), .Y(men_men_n488_));
  AOI210     u0460(.A0(men_men_n269_), .A1(men_men_n483_), .B0(men_men_n488_), .Y(men_men_n489_));
  NO4        u0461(.A(men_men_n189_), .B(men_men_n105_), .C(men_men_n56_), .D(b), .Y(men_men_n490_));
  NA2        u0462(.A(men_men_n390_), .B(men_men_n151_), .Y(men_men_n491_));
  OR2        u0463(.A(k), .B(j), .Y(men_men_n492_));
  NA2        u0464(.A(l), .B(k), .Y(men_men_n493_));
  NA3        u0465(.A(men_men_n493_), .B(men_men_n492_), .C(men_men_n224_), .Y(men_men_n494_));
  AOI210     u0466(.A0(men_men_n237_), .A1(men_men_n341_), .B0(men_men_n86_), .Y(men_men_n495_));
  NOi21      u0467(.An(men_men_n494_), .B(men_men_n495_), .Y(men_men_n496_));
  OR3        u0468(.A(men_men_n496_), .B(men_men_n142_), .C(men_men_n134_), .Y(men_men_n497_));
  INV        u0469(.A(men_men_n279_), .Y(men_men_n498_));
  NA2        u0470(.A(men_men_n403_), .B(men_men_n115_), .Y(men_men_n499_));
  NO4        u0471(.A(men_men_n499_), .B(men_men_n97_), .C(men_men_n114_), .D(e), .Y(men_men_n500_));
  NO3        u0472(.A(men_men_n433_), .B(men_men_n94_), .C(men_men_n130_), .Y(men_men_n501_));
  NO4        u0473(.A(men_men_n501_), .B(men_men_n500_), .C(men_men_n498_), .D(men_men_n324_), .Y(men_men_n502_));
  NA3        u0474(.A(men_men_n502_), .B(men_men_n497_), .C(men_men_n491_), .Y(men_men_n503_));
  NO4        u0475(.A(men_men_n503_), .B(men_men_n490_), .C(men_men_n489_), .D(men_men_n482_), .Y(men_men_n504_));
  NA2        u0476(.A(men_men_n70_), .B(men_men_n67_), .Y(men_men_n505_));
  NOi21      u0477(.An(d), .B(e), .Y(men_men_n506_));
  NAi31      u0478(.An(j), .B(l), .C(i), .Y(men_men_n507_));
  OAI210     u0479(.A0(men_men_n507_), .A1(men_men_n131_), .B0(men_men_n105_), .Y(men_men_n508_));
  NO3        u0480(.A(men_men_n404_), .B(men_men_n349_), .C(men_men_n203_), .Y(men_men_n509_));
  NO2        u0481(.A(men_men_n404_), .B(men_men_n379_), .Y(men_men_n510_));
  NO4        u0482(.A(men_men_n510_), .B(men_men_n509_), .C(men_men_n185_), .D(men_men_n306_), .Y(men_men_n511_));
  NA3        u0483(.A(men_men_n511_), .B(men_men_n505_), .C(men_men_n247_), .Y(men_men_n512_));
  OAI210     u0484(.A0(men_men_n128_), .A1(men_men_n127_), .B0(n), .Y(men_men_n513_));
  NO2        u0485(.A(men_men_n513_), .B(men_men_n130_), .Y(men_men_n514_));
  OR2        u0486(.A(men_men_n300_), .B(men_men_n249_), .Y(men_men_n515_));
  OA210      u0487(.A0(men_men_n515_), .A1(men_men_n514_), .B0(men_men_n194_), .Y(men_men_n516_));
  XO2        u0488(.A(i), .B(h), .Y(men_men_n517_));
  NA3        u0489(.A(men_men_n517_), .B(men_men_n158_), .C(n), .Y(men_men_n518_));
  NAi41      u0490(.An(men_men_n300_), .B(men_men_n518_), .C(men_men_n465_), .D(men_men_n392_), .Y(men_men_n519_));
  NOi32      u0491(.An(men_men_n519_), .Bn(men_men_n477_), .C(men_men_n271_), .Y(men_men_n520_));
  NAi31      u0492(.An(c), .B(f), .C(d), .Y(men_men_n521_));
  AOI210     u0493(.A0(men_men_n280_), .A1(men_men_n197_), .B0(men_men_n521_), .Y(men_men_n522_));
  NOi21      u0494(.An(men_men_n84_), .B(men_men_n522_), .Y(men_men_n523_));
  NA2        u0495(.A(men_men_n231_), .B(men_men_n111_), .Y(men_men_n524_));
  AOI210     u0496(.A0(men_men_n524_), .A1(men_men_n181_), .B0(men_men_n521_), .Y(men_men_n525_));
  INV        u0497(.A(men_men_n525_), .Y(men_men_n526_));
  AO220      u0498(.A0(men_men_n288_), .A1(men_men_n265_), .B0(men_men_n165_), .B1(men_men_n67_), .Y(men_men_n527_));
  NA3        u0499(.A(men_men_n37_), .B(men_men_n36_), .C(f), .Y(men_men_n528_));
  NO2        u0500(.A(men_men_n528_), .B(men_men_n445_), .Y(men_men_n529_));
  NO2        u0501(.A(men_men_n529_), .B(men_men_n296_), .Y(men_men_n530_));
  NAi41      u0502(.An(men_men_n527_), .B(men_men_n530_), .C(men_men_n526_), .D(men_men_n523_), .Y(men_men_n531_));
  NO4        u0503(.A(men_men_n531_), .B(men_men_n520_), .C(men_men_n516_), .D(men_men_n512_), .Y(men_men_n532_));
  NA4        u0504(.A(men_men_n532_), .B(men_men_n504_), .C(men_men_n469_), .D(men_men_n440_), .Y(men11));
  NO2        u0505(.A(men_men_n73_), .B(f), .Y(men_men_n534_));
  NA2        u0506(.A(j), .B(g), .Y(men_men_n535_));
  NAi31      u0507(.An(i), .B(m), .C(l), .Y(men_men_n536_));
  NA3        u0508(.A(m), .B(k), .C(j), .Y(men_men_n537_));
  OAI220     u0509(.A0(men_men_n537_), .A1(men_men_n130_), .B0(men_men_n536_), .B1(men_men_n535_), .Y(men_men_n538_));
  NA2        u0510(.A(men_men_n538_), .B(men_men_n534_), .Y(men_men_n539_));
  NOi32      u0511(.An(e), .Bn(b), .C(f), .Y(men_men_n540_));
  NA2        u0512(.A(men_men_n262_), .B(men_men_n115_), .Y(men_men_n541_));
  NA2        u0513(.A(men_men_n46_), .B(j), .Y(men_men_n542_));
  NAi31      u0514(.An(d), .B(e), .C(a), .Y(men_men_n543_));
  NO2        u0515(.A(men_men_n543_), .B(n), .Y(men_men_n544_));
  NAi41      u0516(.An(f), .B(e), .C(c), .D(a), .Y(men_men_n545_));
  AN2        u0517(.A(men_men_n545_), .B(men_men_n378_), .Y(men_men_n546_));
  AOI210     u0518(.A0(men_men_n546_), .A1(men_men_n404_), .B0(men_men_n272_), .Y(men_men_n547_));
  NA2        u0519(.A(j), .B(i), .Y(men_men_n548_));
  NAi31      u0520(.An(n), .B(m), .C(k), .Y(men_men_n549_));
  NO3        u0521(.A(men_men_n549_), .B(men_men_n548_), .C(men_men_n114_), .Y(men_men_n550_));
  NO4        u0522(.A(n), .B(d), .C(men_men_n117_), .D(a), .Y(men_men_n551_));
  OR2        u0523(.A(n), .B(c), .Y(men_men_n552_));
  NO2        u0524(.A(men_men_n552_), .B(men_men_n147_), .Y(men_men_n553_));
  NO2        u0525(.A(men_men_n553_), .B(men_men_n551_), .Y(men_men_n554_));
  NOi32      u0526(.An(g), .Bn(f), .C(i), .Y(men_men_n555_));
  AOI220     u0527(.A0(men_men_n555_), .A1(men_men_n102_), .B0(men_men_n538_), .B1(f), .Y(men_men_n556_));
  NO2        u0528(.A(men_men_n274_), .B(men_men_n49_), .Y(men_men_n557_));
  NO2        u0529(.A(men_men_n556_), .B(men_men_n554_), .Y(men_men_n558_));
  AOI210     u0530(.A0(men_men_n550_), .A1(men_men_n547_), .B0(men_men_n558_), .Y(men_men_n559_));
  NA2        u0531(.A(men_men_n139_), .B(men_men_n34_), .Y(men_men_n560_));
  OAI220     u0532(.A0(men_men_n560_), .A1(m), .B0(men_men_n542_), .B1(men_men_n237_), .Y(men_men_n561_));
  NOi41      u0533(.An(d), .B(n), .C(e), .D(c), .Y(men_men_n562_));
  NAi32      u0534(.An(e), .Bn(b), .C(c), .Y(men_men_n563_));
  OR2        u0535(.A(men_men_n563_), .B(men_men_n86_), .Y(men_men_n564_));
  AN2        u0536(.A(men_men_n342_), .B(men_men_n320_), .Y(men_men_n565_));
  NA2        u0537(.A(men_men_n565_), .B(men_men_n564_), .Y(men_men_n566_));
  OA210      u0538(.A0(men_men_n566_), .A1(men_men_n562_), .B0(men_men_n561_), .Y(men_men_n567_));
  OAI220     u0539(.A0(men_men_n406_), .A1(men_men_n405_), .B0(men_men_n536_), .B1(men_men_n535_), .Y(men_men_n568_));
  NAi31      u0540(.An(d), .B(c), .C(a), .Y(men_men_n569_));
  NO2        u0541(.A(men_men_n569_), .B(n), .Y(men_men_n570_));
  NA3        u0542(.A(men_men_n570_), .B(men_men_n568_), .C(e), .Y(men_men_n571_));
  INV        u0543(.A(men_men_n571_), .Y(men_men_n572_));
  NO2        u0544(.A(men_men_n276_), .B(n), .Y(men_men_n573_));
  NO2        u0545(.A(men_men_n435_), .B(men_men_n573_), .Y(men_men_n574_));
  NA2        u0546(.A(men_men_n568_), .B(f), .Y(men_men_n575_));
  NAi32      u0547(.An(d), .Bn(a), .C(b), .Y(men_men_n576_));
  NA2        u0548(.A(h), .B(f), .Y(men_men_n577_));
  NO2        u0549(.A(men_men_n577_), .B(men_men_n97_), .Y(men_men_n578_));
  NO3        u0550(.A(men_men_n177_), .B(men_men_n174_), .C(g), .Y(men_men_n579_));
  NA2        u0551(.A(men_men_n579_), .B(men_men_n58_), .Y(men_men_n580_));
  OAI210     u0552(.A0(men_men_n575_), .A1(men_men_n574_), .B0(men_men_n580_), .Y(men_men_n581_));
  AN3        u0553(.A(j), .B(h), .C(g), .Y(men_men_n582_));
  NO2        u0554(.A(men_men_n144_), .B(c), .Y(men_men_n583_));
  NA3        u0555(.A(men_men_n583_), .B(men_men_n582_), .C(men_men_n464_), .Y(men_men_n584_));
  NA3        u0556(.A(f), .B(d), .C(b), .Y(men_men_n585_));
  NO4        u0557(.A(men_men_n585_), .B(men_men_n177_), .C(men_men_n174_), .D(g), .Y(men_men_n586_));
  INV        u0558(.A(men_men_n584_), .Y(men_men_n587_));
  NO4        u0559(.A(men_men_n587_), .B(men_men_n581_), .C(men_men_n572_), .D(men_men_n567_), .Y(men_men_n588_));
  AN3        u0560(.A(men_men_n588_), .B(men_men_n559_), .C(men_men_n539_), .Y(men_men_n589_));
  INV        u0561(.A(k), .Y(men_men_n590_));
  NA3        u0562(.A(l), .B(men_men_n590_), .C(i), .Y(men_men_n591_));
  INV        u0563(.A(men_men_n591_), .Y(men_men_n592_));
  NAi32      u0564(.An(h), .Bn(f), .C(g), .Y(men_men_n593_));
  NAi41      u0565(.An(n), .B(e), .C(c), .D(a), .Y(men_men_n594_));
  OAI210     u0566(.A0(men_men_n543_), .A1(n), .B0(men_men_n594_), .Y(men_men_n595_));
  NA2        u0567(.A(men_men_n595_), .B(m), .Y(men_men_n596_));
  NAi31      u0568(.An(h), .B(g), .C(f), .Y(men_men_n597_));
  OR3        u0569(.A(men_men_n597_), .B(men_men_n276_), .C(men_men_n49_), .Y(men_men_n598_));
  NA4        u0570(.A(men_men_n424_), .B(men_men_n122_), .C(men_men_n115_), .D(e), .Y(men_men_n599_));
  AN2        u0571(.A(men_men_n599_), .B(men_men_n598_), .Y(men_men_n600_));
  NO3        u0572(.A(men_men_n593_), .B(men_men_n73_), .C(men_men_n75_), .Y(men_men_n601_));
  NO4        u0573(.A(men_men_n597_), .B(men_men_n552_), .C(men_men_n147_), .D(men_men_n75_), .Y(men_men_n602_));
  OR2        u0574(.A(men_men_n602_), .B(men_men_n601_), .Y(men_men_n603_));
  NAi21      u0575(.An(men_men_n603_), .B(men_men_n600_), .Y(men_men_n604_));
  NAi31      u0576(.An(f), .B(h), .C(g), .Y(men_men_n605_));
  NO4        u0577(.A(men_men_n311_), .B(men_men_n605_), .C(men_men_n73_), .D(men_men_n75_), .Y(men_men_n606_));
  NOi32      u0578(.An(b), .Bn(a), .C(c), .Y(men_men_n607_));
  NOi41      u0579(.An(men_men_n607_), .B(men_men_n358_), .C(men_men_n69_), .D(men_men_n118_), .Y(men_men_n608_));
  OR2        u0580(.A(men_men_n608_), .B(men_men_n606_), .Y(men_men_n609_));
  NOi32      u0581(.An(d), .Bn(a), .C(e), .Y(men_men_n610_));
  NA2        u0582(.A(men_men_n610_), .B(men_men_n115_), .Y(men_men_n611_));
  NO2        u0583(.A(n), .B(c), .Y(men_men_n612_));
  NA3        u0584(.A(men_men_n612_), .B(men_men_n29_), .C(m), .Y(men_men_n613_));
  NA2        u0585(.A(men_men_n613_), .B(men_men_n611_), .Y(men_men_n614_));
  NOi32      u0586(.An(e), .Bn(a), .C(d), .Y(men_men_n615_));
  AOI210     u0587(.A0(men_men_n29_), .A1(d), .B0(men_men_n615_), .Y(men_men_n616_));
  AOI210     u0588(.A0(men_men_n616_), .A1(men_men_n216_), .B0(men_men_n560_), .Y(men_men_n617_));
  AOI210     u0589(.A0(men_men_n617_), .A1(men_men_n614_), .B0(men_men_n609_), .Y(men_men_n618_));
  INV        u0590(.A(men_men_n618_), .Y(men_men_n619_));
  AOI210     u0591(.A0(men_men_n604_), .A1(men_men_n592_), .B0(men_men_n619_), .Y(men_men_n620_));
  NO3        u0592(.A(men_men_n318_), .B(men_men_n61_), .C(n), .Y(men_men_n621_));
  NA3        u0593(.A(men_men_n521_), .B(men_men_n172_), .C(men_men_n171_), .Y(men_men_n622_));
  NA2        u0594(.A(men_men_n466_), .B(men_men_n234_), .Y(men_men_n623_));
  OR2        u0595(.A(men_men_n623_), .B(men_men_n622_), .Y(men_men_n624_));
  NA2        u0596(.A(men_men_n76_), .B(men_men_n115_), .Y(men_men_n625_));
  NO2        u0597(.A(men_men_n625_), .B(men_men_n45_), .Y(men_men_n626_));
  AOI220     u0598(.A0(men_men_n626_), .A1(men_men_n547_), .B0(men_men_n624_), .B1(men_men_n621_), .Y(men_men_n627_));
  NO2        u0599(.A(men_men_n627_), .B(men_men_n89_), .Y(men_men_n628_));
  NA3        u0600(.A(men_men_n562_), .B(men_men_n344_), .C(men_men_n46_), .Y(men_men_n629_));
  NOi32      u0601(.An(e), .Bn(c), .C(f), .Y(men_men_n630_));
  NOi21      u0602(.An(f), .B(g), .Y(men_men_n631_));
  NO2        u0603(.A(men_men_n631_), .B(men_men_n214_), .Y(men_men_n632_));
  AOI220     u0604(.A0(men_men_n632_), .A1(men_men_n400_), .B0(men_men_n630_), .B1(men_men_n176_), .Y(men_men_n633_));
  NA3        u0605(.A(men_men_n633_), .B(men_men_n629_), .C(men_men_n179_), .Y(men_men_n634_));
  AOI210     u0606(.A0(men_men_n546_), .A1(men_men_n404_), .B0(men_men_n301_), .Y(men_men_n635_));
  NA2        u0607(.A(men_men_n635_), .B(men_men_n266_), .Y(men_men_n636_));
  NOi21      u0608(.An(j), .B(l), .Y(men_men_n637_));
  NAi21      u0609(.An(k), .B(h), .Y(men_men_n638_));
  NO2        u0610(.A(men_men_n638_), .B(men_men_n264_), .Y(men_men_n639_));
  NA2        u0611(.A(men_men_n639_), .B(men_men_n637_), .Y(men_men_n640_));
  OR2        u0612(.A(men_men_n640_), .B(men_men_n596_), .Y(men_men_n641_));
  NOi31      u0613(.An(m), .B(n), .C(k), .Y(men_men_n642_));
  NA2        u0614(.A(men_men_n637_), .B(men_men_n642_), .Y(men_men_n643_));
  AOI210     u0615(.A0(men_men_n404_), .A1(men_men_n378_), .B0(men_men_n301_), .Y(men_men_n644_));
  NAi21      u0616(.An(men_men_n643_), .B(men_men_n644_), .Y(men_men_n645_));
  NO2        u0617(.A(men_men_n276_), .B(men_men_n49_), .Y(men_men_n646_));
  NO2        u0618(.A(men_men_n311_), .B(men_men_n605_), .Y(men_men_n647_));
  NO2        u0619(.A(men_men_n543_), .B(men_men_n49_), .Y(men_men_n648_));
  AOI220     u0620(.A0(men_men_n648_), .A1(men_men_n647_), .B0(men_men_n646_), .B1(men_men_n578_), .Y(men_men_n649_));
  NA4        u0621(.A(men_men_n649_), .B(men_men_n645_), .C(men_men_n641_), .D(men_men_n636_), .Y(men_men_n650_));
  NA2        u0622(.A(men_men_n111_), .B(men_men_n36_), .Y(men_men_n651_));
  NO2        u0623(.A(k), .B(men_men_n217_), .Y(men_men_n652_));
  INV        u0624(.A(men_men_n367_), .Y(men_men_n653_));
  NO2        u0625(.A(men_men_n653_), .B(n), .Y(men_men_n654_));
  NAi31      u0626(.An(men_men_n651_), .B(men_men_n654_), .C(men_men_n652_), .Y(men_men_n655_));
  NO2        u0627(.A(men_men_n542_), .B(men_men_n177_), .Y(men_men_n656_));
  NA3        u0628(.A(men_men_n563_), .B(men_men_n271_), .C(men_men_n143_), .Y(men_men_n657_));
  NA2        u0629(.A(men_men_n517_), .B(men_men_n158_), .Y(men_men_n658_));
  NO3        u0630(.A(men_men_n401_), .B(men_men_n658_), .C(men_men_n89_), .Y(men_men_n659_));
  AOI210     u0631(.A0(men_men_n657_), .A1(men_men_n656_), .B0(men_men_n659_), .Y(men_men_n660_));
  AN3        u0632(.A(f), .B(d), .C(b), .Y(men_men_n661_));
  OAI210     u0633(.A0(men_men_n661_), .A1(men_men_n129_), .B0(n), .Y(men_men_n662_));
  NA3        u0634(.A(men_men_n517_), .B(men_men_n158_), .C(men_men_n217_), .Y(men_men_n663_));
  AOI210     u0635(.A0(men_men_n662_), .A1(men_men_n236_), .B0(men_men_n663_), .Y(men_men_n664_));
  NAi31      u0636(.An(m), .B(n), .C(k), .Y(men_men_n665_));
  OR2        u0637(.A(men_men_n134_), .B(men_men_n61_), .Y(men_men_n666_));
  OAI210     u0638(.A0(men_men_n666_), .A1(men_men_n665_), .B0(men_men_n254_), .Y(men_men_n667_));
  OAI210     u0639(.A0(men_men_n667_), .A1(men_men_n664_), .B0(j), .Y(men_men_n668_));
  NA3        u0640(.A(men_men_n668_), .B(men_men_n660_), .C(men_men_n655_), .Y(men_men_n669_));
  NO4        u0641(.A(men_men_n669_), .B(men_men_n650_), .C(men_men_n634_), .D(men_men_n628_), .Y(men_men_n670_));
  NA2        u0642(.A(men_men_n388_), .B(men_men_n161_), .Y(men_men_n671_));
  NAi31      u0643(.An(g), .B(h), .C(f), .Y(men_men_n672_));
  OR3        u0644(.A(men_men_n672_), .B(men_men_n276_), .C(n), .Y(men_men_n673_));
  OA210      u0645(.A0(men_men_n543_), .A1(n), .B0(men_men_n594_), .Y(men_men_n674_));
  NA3        u0646(.A(men_men_n422_), .B(men_men_n122_), .C(men_men_n86_), .Y(men_men_n675_));
  OAI210     u0647(.A0(men_men_n674_), .A1(men_men_n93_), .B0(men_men_n675_), .Y(men_men_n676_));
  NOi21      u0648(.An(men_men_n673_), .B(men_men_n676_), .Y(men_men_n677_));
  AOI210     u0649(.A0(men_men_n677_), .A1(men_men_n671_), .B0(men_men_n537_), .Y(men_men_n678_));
  NO3        u0650(.A(g), .B(men_men_n216_), .C(men_men_n56_), .Y(men_men_n679_));
  NAi21      u0651(.An(h), .B(j), .Y(men_men_n680_));
  NO2        u0652(.A(men_men_n524_), .B(men_men_n89_), .Y(men_men_n681_));
  OAI210     u0653(.A0(men_men_n681_), .A1(men_men_n400_), .B0(men_men_n679_), .Y(men_men_n682_));
  OR2        u0654(.A(men_men_n73_), .B(men_men_n75_), .Y(men_men_n683_));
  NA2        u0655(.A(men_men_n607_), .B(men_men_n346_), .Y(men_men_n684_));
  OA220      u0656(.A0(men_men_n643_), .A1(men_men_n684_), .B0(men_men_n640_), .B1(men_men_n683_), .Y(men_men_n685_));
  NA3        u0657(.A(men_men_n534_), .B(men_men_n102_), .C(men_men_n101_), .Y(men_men_n686_));
  AN2        u0658(.A(h), .B(f), .Y(men_men_n687_));
  NA2        u0659(.A(men_men_n687_), .B(men_men_n37_), .Y(men_men_n688_));
  NA2        u0660(.A(men_men_n102_), .B(men_men_n46_), .Y(men_men_n689_));
  OAI220     u0661(.A0(men_men_n689_), .A1(men_men_n335_), .B0(men_men_n688_), .B1(men_men_n471_), .Y(men_men_n690_));
  AOI210     u0662(.A0(men_men_n576_), .A1(men_men_n434_), .B0(men_men_n49_), .Y(men_men_n691_));
  OAI220     u0663(.A0(men_men_n597_), .A1(men_men_n591_), .B0(men_men_n328_), .B1(men_men_n535_), .Y(men_men_n692_));
  AOI210     u0664(.A0(men_men_n692_), .A1(men_men_n691_), .B0(men_men_n690_), .Y(men_men_n693_));
  NA4        u0665(.A(men_men_n693_), .B(men_men_n686_), .C(men_men_n685_), .D(men_men_n682_), .Y(men_men_n694_));
  NO2        u0666(.A(men_men_n255_), .B(f), .Y(men_men_n695_));
  NO2        u0667(.A(men_men_n631_), .B(men_men_n61_), .Y(men_men_n696_));
  NO3        u0668(.A(men_men_n696_), .B(men_men_n695_), .C(men_men_n34_), .Y(men_men_n697_));
  NA2        u0669(.A(men_men_n331_), .B(men_men_n139_), .Y(men_men_n698_));
  NA2        u0670(.A(men_men_n131_), .B(men_men_n49_), .Y(men_men_n699_));
  AOI220     u0671(.A0(men_men_n699_), .A1(men_men_n540_), .B0(men_men_n367_), .B1(men_men_n115_), .Y(men_men_n700_));
  OA220      u0672(.A0(men_men_n700_), .A1(men_men_n560_), .B0(men_men_n365_), .B1(men_men_n113_), .Y(men_men_n701_));
  OAI210     u0673(.A0(men_men_n698_), .A1(men_men_n697_), .B0(men_men_n701_), .Y(men_men_n702_));
  NO3        u0674(.A(men_men_n409_), .B(men_men_n194_), .C(men_men_n193_), .Y(men_men_n703_));
  NA2        u0675(.A(men_men_n703_), .B(men_men_n234_), .Y(men_men_n704_));
  NA3        u0676(.A(men_men_n704_), .B(men_men_n257_), .C(j), .Y(men_men_n705_));
  NA2        u0677(.A(men_men_n470_), .B(men_men_n86_), .Y(men_men_n706_));
  NO4        u0678(.A(men_men_n537_), .B(men_men_n706_), .C(men_men_n130_), .D(men_men_n216_), .Y(men_men_n707_));
  INV        u0679(.A(men_men_n707_), .Y(men_men_n708_));
  NA3        u0680(.A(men_men_n708_), .B(men_men_n705_), .C(men_men_n407_), .Y(men_men_n709_));
  NO4        u0681(.A(men_men_n709_), .B(men_men_n702_), .C(men_men_n694_), .D(men_men_n678_), .Y(men_men_n710_));
  NA4        u0682(.A(men_men_n710_), .B(men_men_n670_), .C(men_men_n620_), .D(men_men_n589_), .Y(men08));
  NO2        u0683(.A(k), .B(h), .Y(men_men_n712_));
  AO210      u0684(.A0(men_men_n255_), .A1(men_men_n456_), .B0(men_men_n712_), .Y(men_men_n713_));
  NO2        u0685(.A(men_men_n713_), .B(men_men_n299_), .Y(men_men_n714_));
  NA2        u0686(.A(men_men_n630_), .B(men_men_n86_), .Y(men_men_n715_));
  NA2        u0687(.A(men_men_n715_), .B(men_men_n466_), .Y(men_men_n716_));
  AOI210     u0688(.A0(men_men_n716_), .A1(men_men_n714_), .B0(men_men_n501_), .Y(men_men_n717_));
  NA2        u0689(.A(men_men_n86_), .B(men_men_n112_), .Y(men_men_n718_));
  NO2        u0690(.A(men_men_n718_), .B(men_men_n57_), .Y(men_men_n719_));
  NO4        u0691(.A(men_men_n385_), .B(men_men_n114_), .C(j), .D(men_men_n217_), .Y(men_men_n720_));
  NA2        u0692(.A(men_men_n585_), .B(men_men_n236_), .Y(men_men_n721_));
  AOI220     u0693(.A0(men_men_n721_), .A1(men_men_n352_), .B0(men_men_n720_), .B1(men_men_n719_), .Y(men_men_n722_));
  AOI210     u0694(.A0(men_men_n585_), .A1(men_men_n154_), .B0(men_men_n86_), .Y(men_men_n723_));
  NA4        u0695(.A(men_men_n219_), .B(men_men_n139_), .C(men_men_n45_), .D(h), .Y(men_men_n724_));
  AN2        u0696(.A(l), .B(k), .Y(men_men_n725_));
  NA4        u0697(.A(men_men_n725_), .B(men_men_n111_), .C(men_men_n75_), .D(men_men_n217_), .Y(men_men_n726_));
  OAI210     u0698(.A0(men_men_n724_), .A1(g), .B0(men_men_n726_), .Y(men_men_n727_));
  NA2        u0699(.A(men_men_n727_), .B(men_men_n723_), .Y(men_men_n728_));
  NA4        u0700(.A(men_men_n728_), .B(men_men_n722_), .C(men_men_n717_), .D(men_men_n354_), .Y(men_men_n729_));
  AN2        u0701(.A(men_men_n544_), .B(men_men_n98_), .Y(men_men_n730_));
  NO4        u0702(.A(men_men_n174_), .B(men_men_n399_), .C(men_men_n114_), .D(g), .Y(men_men_n731_));
  AOI210     u0703(.A0(men_men_n731_), .A1(men_men_n721_), .B0(men_men_n529_), .Y(men_men_n732_));
  NA2        u0704(.A(men_men_n632_), .B(men_men_n351_), .Y(men_men_n733_));
  NAi31      u0705(.An(men_men_n730_), .B(men_men_n733_), .C(men_men_n732_), .Y(men_men_n734_));
  NO2        u0706(.A(men_men_n546_), .B(men_men_n35_), .Y(men_men_n735_));
  OAI210     u0707(.A0(men_men_n563_), .A1(men_men_n47_), .B0(men_men_n666_), .Y(men_men_n736_));
  NO2        u0708(.A(men_men_n493_), .B(men_men_n131_), .Y(men_men_n737_));
  AOI210     u0709(.A0(men_men_n737_), .A1(men_men_n736_), .B0(men_men_n735_), .Y(men_men_n738_));
  NO3        u0710(.A(men_men_n318_), .B(men_men_n130_), .C(men_men_n41_), .Y(men_men_n739_));
  INV        u0711(.A(men_men_n726_), .Y(men_men_n740_));
  NA2        u0712(.A(men_men_n713_), .B(men_men_n135_), .Y(men_men_n741_));
  AOI220     u0713(.A0(men_men_n741_), .A1(men_men_n408_), .B0(men_men_n740_), .B1(men_men_n78_), .Y(men_men_n742_));
  OAI210     u0714(.A0(men_men_n738_), .A1(men_men_n89_), .B0(men_men_n742_), .Y(men_men_n743_));
  NA2        u0715(.A(men_men_n367_), .B(men_men_n43_), .Y(men_men_n744_));
  NA3        u0716(.A(men_men_n704_), .B(men_men_n337_), .C(men_men_n391_), .Y(men_men_n745_));
  NA2        u0717(.A(men_men_n725_), .B(men_men_n224_), .Y(men_men_n746_));
  NO2        u0718(.A(men_men_n746_), .B(men_men_n330_), .Y(men_men_n747_));
  AOI210     u0719(.A0(men_men_n747_), .A1(men_men_n695_), .B0(men_men_n500_), .Y(men_men_n748_));
  NA3        u0720(.A(m), .B(l), .C(k), .Y(men_men_n749_));
  AOI210     u0721(.A0(men_men_n675_), .A1(men_men_n673_), .B0(men_men_n749_), .Y(men_men_n750_));
  NO2        u0722(.A(men_men_n545_), .B(men_men_n272_), .Y(men_men_n751_));
  NOi21      u0723(.An(men_men_n751_), .B(men_men_n541_), .Y(men_men_n752_));
  NA4        u0724(.A(men_men_n115_), .B(l), .C(k), .D(men_men_n89_), .Y(men_men_n753_));
  NA3        u0725(.A(men_men_n122_), .B(men_men_n417_), .C(i), .Y(men_men_n754_));
  NO2        u0726(.A(men_men_n754_), .B(men_men_n753_), .Y(men_men_n755_));
  NO3        u0727(.A(men_men_n755_), .B(men_men_n752_), .C(men_men_n750_), .Y(men_men_n756_));
  NA4        u0728(.A(men_men_n756_), .B(men_men_n748_), .C(men_men_n745_), .D(men_men_n744_), .Y(men_men_n757_));
  NO4        u0729(.A(men_men_n757_), .B(men_men_n743_), .C(men_men_n734_), .D(men_men_n729_), .Y(men_men_n758_));
  NA2        u0730(.A(men_men_n632_), .B(men_men_n400_), .Y(men_men_n759_));
  INV        u0731(.A(men_men_n510_), .Y(men_men_n760_));
  NA3        u0732(.A(men_men_n760_), .B(men_men_n759_), .C(men_men_n254_), .Y(men_men_n761_));
  NA2        u0733(.A(men_men_n725_), .B(men_men_n75_), .Y(men_men_n762_));
  NO4        u0734(.A(men_men_n703_), .B(men_men_n174_), .C(n), .D(i), .Y(men_men_n763_));
  NOi21      u0735(.An(h), .B(j), .Y(men_men_n764_));
  NA2        u0736(.A(men_men_n764_), .B(f), .Y(men_men_n765_));
  NO2        u0737(.A(men_men_n765_), .B(men_men_n251_), .Y(men_men_n766_));
  NO2        u0738(.A(men_men_n766_), .B(men_men_n763_), .Y(men_men_n767_));
  OAI220     u0739(.A0(men_men_n767_), .A1(men_men_n762_), .B0(men_men_n600_), .B1(men_men_n62_), .Y(men_men_n768_));
  AOI210     u0740(.A0(men_men_n761_), .A1(l), .B0(men_men_n768_), .Y(men_men_n769_));
  NO2        u0741(.A(j), .B(i), .Y(men_men_n770_));
  NA3        u0742(.A(men_men_n770_), .B(men_men_n82_), .C(l), .Y(men_men_n771_));
  NA2        u0743(.A(men_men_n770_), .B(men_men_n33_), .Y(men_men_n772_));
  NA2        u0744(.A(men_men_n427_), .B(men_men_n122_), .Y(men_men_n773_));
  OA220      u0745(.A0(men_men_n773_), .A1(men_men_n772_), .B0(men_men_n771_), .B1(men_men_n596_), .Y(men_men_n774_));
  NO3        u0746(.A(men_men_n149_), .B(men_men_n49_), .C(men_men_n112_), .Y(men_men_n775_));
  NO3        u0747(.A(men_men_n552_), .B(men_men_n147_), .C(men_men_n75_), .Y(men_men_n776_));
  NO3        u0748(.A(men_men_n493_), .B(men_men_n446_), .C(j), .Y(men_men_n777_));
  OAI210     u0749(.A0(men_men_n776_), .A1(men_men_n775_), .B0(men_men_n777_), .Y(men_men_n778_));
  INV        u0750(.A(men_men_n778_), .Y(men_men_n779_));
  NA2        u0751(.A(k), .B(j), .Y(men_men_n780_));
  NO3        u0752(.A(men_men_n299_), .B(men_men_n780_), .C(men_men_n40_), .Y(men_men_n781_));
  AOI210     u0753(.A0(men_men_n540_), .A1(n), .B0(men_men_n562_), .Y(men_men_n782_));
  NA2        u0754(.A(men_men_n782_), .B(men_men_n565_), .Y(men_men_n783_));
  AN3        u0755(.A(men_men_n783_), .B(men_men_n781_), .C(men_men_n101_), .Y(men_men_n784_));
  NA2        u0756(.A(men_men_n623_), .B(men_men_n308_), .Y(men_men_n785_));
  NAi31      u0757(.An(men_men_n616_), .B(men_men_n95_), .C(men_men_n86_), .Y(men_men_n786_));
  NA2        u0758(.A(men_men_n786_), .B(men_men_n785_), .Y(men_men_n787_));
  NO2        u0759(.A(men_men_n299_), .B(men_men_n135_), .Y(men_men_n788_));
  AOI220     u0760(.A0(men_men_n788_), .A1(men_men_n632_), .B0(men_men_n739_), .B1(men_men_n723_), .Y(men_men_n789_));
  NO2        u0761(.A(men_men_n749_), .B(men_men_n93_), .Y(men_men_n790_));
  NA2        u0762(.A(men_men_n790_), .B(men_men_n595_), .Y(men_men_n791_));
  NO2        u0763(.A(men_men_n597_), .B(men_men_n118_), .Y(men_men_n792_));
  OAI210     u0764(.A0(men_men_n792_), .A1(men_men_n777_), .B0(men_men_n691_), .Y(men_men_n793_));
  NA3        u0765(.A(men_men_n793_), .B(men_men_n791_), .C(men_men_n789_), .Y(men_men_n794_));
  OR4        u0766(.A(men_men_n794_), .B(men_men_n787_), .C(men_men_n784_), .D(men_men_n779_), .Y(men_men_n795_));
  NA3        u0767(.A(men_men_n782_), .B(men_men_n565_), .C(men_men_n564_), .Y(men_men_n796_));
  NA4        u0768(.A(men_men_n796_), .B(men_men_n219_), .C(men_men_n456_), .D(men_men_n34_), .Y(men_men_n797_));
  NO4        u0769(.A(men_men_n493_), .B(men_men_n441_), .C(j), .D(f), .Y(men_men_n798_));
  OAI220     u0770(.A0(men_men_n724_), .A1(men_men_n715_), .B0(men_men_n335_), .B1(men_men_n38_), .Y(men_men_n799_));
  AOI210     u0771(.A0(men_men_n798_), .A1(men_men_n261_), .B0(men_men_n799_), .Y(men_men_n800_));
  NA3        u0772(.A(men_men_n555_), .B(men_men_n292_), .C(h), .Y(men_men_n801_));
  NOi21      u0773(.An(men_men_n691_), .B(men_men_n801_), .Y(men_men_n802_));
  NO2        u0774(.A(men_men_n94_), .B(men_men_n47_), .Y(men_men_n803_));
  OAI220     u0775(.A0(men_men_n801_), .A1(men_men_n613_), .B0(men_men_n771_), .B1(men_men_n683_), .Y(men_men_n804_));
  AOI210     u0776(.A0(men_men_n803_), .A1(men_men_n654_), .B0(men_men_n804_), .Y(men_men_n805_));
  NAi41      u0777(.An(men_men_n802_), .B(men_men_n805_), .C(men_men_n800_), .D(men_men_n797_), .Y(men_men_n806_));
  OR2        u0778(.A(men_men_n790_), .B(men_men_n98_), .Y(men_men_n807_));
  AOI220     u0779(.A0(men_men_n807_), .A1(men_men_n242_), .B0(men_men_n777_), .B1(men_men_n646_), .Y(men_men_n808_));
  NO2        u0780(.A(men_men_n674_), .B(men_men_n75_), .Y(men_men_n809_));
  AOI210     u0781(.A0(men_men_n798_), .A1(men_men_n809_), .B0(men_men_n339_), .Y(men_men_n810_));
  OAI210     u0782(.A0(men_men_n749_), .A1(men_men_n672_), .B0(men_men_n528_), .Y(men_men_n811_));
  NA3        u0783(.A(men_men_n253_), .B(men_men_n59_), .C(b), .Y(men_men_n812_));
  AOI220     u0784(.A0(men_men_n612_), .A1(men_men_n29_), .B0(men_men_n470_), .B1(men_men_n86_), .Y(men_men_n813_));
  NA2        u0785(.A(men_men_n813_), .B(men_men_n812_), .Y(men_men_n814_));
  NO2        u0786(.A(men_men_n801_), .B(men_men_n499_), .Y(men_men_n815_));
  AOI210     u0787(.A0(men_men_n814_), .A1(men_men_n811_), .B0(men_men_n815_), .Y(men_men_n816_));
  NA3        u0788(.A(men_men_n816_), .B(men_men_n810_), .C(men_men_n808_), .Y(men_men_n817_));
  NOi41      u0789(.An(men_men_n774_), .B(men_men_n817_), .C(men_men_n806_), .D(men_men_n795_), .Y(men_men_n818_));
  OR3        u0790(.A(men_men_n724_), .B(men_men_n236_), .C(g), .Y(men_men_n819_));
  NO3        u0791(.A(men_men_n345_), .B(men_men_n301_), .C(men_men_n114_), .Y(men_men_n820_));
  NA2        u0792(.A(men_men_n820_), .B(men_men_n783_), .Y(men_men_n821_));
  NA2        u0793(.A(men_men_n46_), .B(men_men_n56_), .Y(men_men_n822_));
  NO3        u0794(.A(men_men_n822_), .B(men_men_n772_), .C(men_men_n276_), .Y(men_men_n823_));
  NO3        u0795(.A(men_men_n535_), .B(men_men_n96_), .C(h), .Y(men_men_n824_));
  AOI210     u0796(.A0(men_men_n824_), .A1(men_men_n719_), .B0(men_men_n823_), .Y(men_men_n825_));
  NA4        u0797(.A(men_men_n825_), .B(men_men_n821_), .C(men_men_n819_), .D(men_men_n410_), .Y(men_men_n826_));
  OR2        u0798(.A(men_men_n672_), .B(men_men_n94_), .Y(men_men_n827_));
  NOi31      u0799(.An(b), .B(d), .C(a), .Y(men_men_n828_));
  NO2        u0800(.A(men_men_n828_), .B(men_men_n610_), .Y(men_men_n829_));
  NO2        u0801(.A(men_men_n829_), .B(n), .Y(men_men_n830_));
  NOi21      u0802(.An(men_men_n813_), .B(men_men_n830_), .Y(men_men_n831_));
  OAI220     u0803(.A0(men_men_n831_), .A1(men_men_n827_), .B0(men_men_n801_), .B1(men_men_n611_), .Y(men_men_n832_));
  NO2        u0804(.A(men_men_n563_), .B(men_men_n86_), .Y(men_men_n833_));
  NA2        u0805(.A(men_men_n820_), .B(men_men_n833_), .Y(men_men_n834_));
  OAI210     u0806(.A0(men_men_n724_), .A1(men_men_n401_), .B0(men_men_n834_), .Y(men_men_n835_));
  NO2        u0807(.A(men_men_n703_), .B(n), .Y(men_men_n836_));
  AOI220     u0808(.A0(men_men_n788_), .A1(men_men_n679_), .B0(men_men_n836_), .B1(men_men_n714_), .Y(men_men_n837_));
  NA2        u0809(.A(men_men_n122_), .B(men_men_n86_), .Y(men_men_n838_));
  AOI210     u0810(.A0(men_men_n431_), .A1(men_men_n423_), .B0(men_men_n838_), .Y(men_men_n839_));
  NA2        u0811(.A(men_men_n747_), .B(men_men_n34_), .Y(men_men_n840_));
  NAi21      u0812(.An(men_men_n753_), .B(men_men_n442_), .Y(men_men_n841_));
  NO2        u0813(.A(men_men_n272_), .B(i), .Y(men_men_n842_));
  NA2        u0814(.A(men_men_n731_), .B(men_men_n353_), .Y(men_men_n843_));
  OAI210     u0815(.A0(men_men_n602_), .A1(men_men_n601_), .B0(men_men_n368_), .Y(men_men_n844_));
  AN3        u0816(.A(men_men_n844_), .B(men_men_n843_), .C(men_men_n841_), .Y(men_men_n845_));
  NAi41      u0817(.An(men_men_n839_), .B(men_men_n845_), .C(men_men_n840_), .D(men_men_n837_), .Y(men_men_n846_));
  NO4        u0818(.A(men_men_n846_), .B(men_men_n835_), .C(men_men_n832_), .D(men_men_n826_), .Y(men_men_n847_));
  NA4        u0819(.A(men_men_n847_), .B(men_men_n818_), .C(men_men_n769_), .D(men_men_n758_), .Y(men09));
  INV        u0820(.A(men_men_n123_), .Y(men_men_n849_));
  NA2        u0821(.A(f), .B(e), .Y(men_men_n850_));
  NO2        u0822(.A(men_men_n229_), .B(men_men_n114_), .Y(men_men_n851_));
  NA2        u0823(.A(men_men_n851_), .B(g), .Y(men_men_n852_));
  NA4        u0824(.A(men_men_n311_), .B(men_men_n479_), .C(men_men_n263_), .D(men_men_n120_), .Y(men_men_n853_));
  AOI210     u0825(.A0(men_men_n853_), .A1(g), .B0(men_men_n476_), .Y(men_men_n854_));
  AOI210     u0826(.A0(men_men_n854_), .A1(men_men_n852_), .B0(men_men_n850_), .Y(men_men_n855_));
  NA2        u0827(.A(men_men_n450_), .B(e), .Y(men_men_n856_));
  NO2        u0828(.A(men_men_n856_), .B(men_men_n521_), .Y(men_men_n857_));
  AOI210     u0829(.A0(men_men_n855_), .A1(men_men_n849_), .B0(men_men_n857_), .Y(men_men_n858_));
  NA3        u0830(.A(m), .B(l), .C(i), .Y(men_men_n859_));
  OAI220     u0831(.A0(men_men_n597_), .A1(men_men_n859_), .B0(men_men_n358_), .B1(men_men_n536_), .Y(men_men_n860_));
  NA4        u0832(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(f), .Y(men_men_n861_));
  NAi31      u0833(.An(men_men_n860_), .B(men_men_n861_), .C(men_men_n447_), .Y(men_men_n862_));
  NA3        u0834(.A(men_men_n827_), .B(men_men_n575_), .C(men_men_n528_), .Y(men_men_n863_));
  OA210      u0835(.A0(men_men_n863_), .A1(men_men_n862_), .B0(men_men_n830_), .Y(men_men_n864_));
  INV        u0836(.A(men_men_n342_), .Y(men_men_n865_));
  NO2        u0837(.A(men_men_n128_), .B(men_men_n127_), .Y(men_men_n866_));
  NOi31      u0838(.An(k), .B(m), .C(l), .Y(men_men_n867_));
  NO2        u0839(.A(men_men_n344_), .B(men_men_n867_), .Y(men_men_n868_));
  AOI210     u0840(.A0(men_men_n868_), .A1(men_men_n866_), .B0(men_men_n605_), .Y(men_men_n869_));
  NA2        u0841(.A(men_men_n812_), .B(men_men_n335_), .Y(men_men_n870_));
  NA2        u0842(.A(men_men_n346_), .B(men_men_n348_), .Y(men_men_n871_));
  OAI210     u0843(.A0(men_men_n206_), .A1(men_men_n216_), .B0(men_men_n871_), .Y(men_men_n872_));
  AOI220     u0844(.A0(men_men_n872_), .A1(men_men_n870_), .B0(men_men_n869_), .B1(men_men_n865_), .Y(men_men_n873_));
  NA2        u0845(.A(men_men_n168_), .B(men_men_n116_), .Y(men_men_n874_));
  NA3        u0846(.A(men_men_n874_), .B(men_men_n713_), .C(men_men_n135_), .Y(men_men_n875_));
  NA3        u0847(.A(men_men_n875_), .B(men_men_n191_), .C(men_men_n31_), .Y(men_men_n876_));
  NA4        u0848(.A(men_men_n876_), .B(men_men_n873_), .C(men_men_n633_), .D(men_men_n84_), .Y(men_men_n877_));
  NO2        u0849(.A(men_men_n593_), .B(men_men_n507_), .Y(men_men_n878_));
  NA2        u0850(.A(men_men_n878_), .B(men_men_n191_), .Y(men_men_n879_));
  NOi21      u0851(.An(f), .B(d), .Y(men_men_n880_));
  NA2        u0852(.A(men_men_n880_), .B(m), .Y(men_men_n881_));
  NO2        u0853(.A(men_men_n881_), .B(men_men_n52_), .Y(men_men_n882_));
  NOi32      u0854(.An(g), .Bn(f), .C(d), .Y(men_men_n883_));
  NA4        u0855(.A(men_men_n883_), .B(men_men_n612_), .C(men_men_n29_), .D(m), .Y(men_men_n884_));
  NOi21      u0856(.An(men_men_n312_), .B(men_men_n884_), .Y(men_men_n885_));
  AOI210     u0857(.A0(men_men_n882_), .A1(men_men_n553_), .B0(men_men_n885_), .Y(men_men_n886_));
  NA2        u0858(.A(men_men_n263_), .B(men_men_n120_), .Y(men_men_n887_));
  AN2        u0859(.A(f), .B(d), .Y(men_men_n888_));
  NA3        u0860(.A(men_men_n484_), .B(men_men_n888_), .C(men_men_n86_), .Y(men_men_n889_));
  NO3        u0861(.A(men_men_n889_), .B(men_men_n75_), .C(men_men_n217_), .Y(men_men_n890_));
  NO2        u0862(.A(men_men_n285_), .B(men_men_n56_), .Y(men_men_n891_));
  NA2        u0863(.A(men_men_n887_), .B(men_men_n890_), .Y(men_men_n892_));
  NAi41      u0864(.An(men_men_n498_), .B(men_men_n892_), .C(men_men_n886_), .D(men_men_n879_), .Y(men_men_n893_));
  NO4        u0865(.A(men_men_n631_), .B(men_men_n131_), .C(men_men_n330_), .D(men_men_n150_), .Y(men_men_n894_));
  NO2        u0866(.A(men_men_n665_), .B(men_men_n330_), .Y(men_men_n895_));
  AN2        u0867(.A(men_men_n895_), .B(men_men_n695_), .Y(men_men_n896_));
  NO3        u0868(.A(men_men_n896_), .B(men_men_n894_), .C(men_men_n238_), .Y(men_men_n897_));
  NA2        u0869(.A(men_men_n610_), .B(men_men_n86_), .Y(men_men_n898_));
  NO2        u0870(.A(men_men_n871_), .B(men_men_n898_), .Y(men_men_n899_));
  NA3        u0871(.A(men_men_n158_), .B(men_men_n111_), .C(men_men_n110_), .Y(men_men_n900_));
  OAI220     u0872(.A0(men_men_n889_), .A1(men_men_n436_), .B0(men_men_n342_), .B1(men_men_n900_), .Y(men_men_n901_));
  NOi41      u0873(.An(men_men_n227_), .B(men_men_n901_), .C(men_men_n899_), .D(men_men_n306_), .Y(men_men_n902_));
  NA2        u0874(.A(c), .B(men_men_n117_), .Y(men_men_n903_));
  NO2        u0875(.A(men_men_n903_), .B(men_men_n414_), .Y(men_men_n904_));
  NA3        u0876(.A(men_men_n904_), .B(men_men_n519_), .C(f), .Y(men_men_n905_));
  OR2        u0877(.A(men_men_n672_), .B(men_men_n549_), .Y(men_men_n906_));
  INV        u0878(.A(men_men_n906_), .Y(men_men_n907_));
  NA2        u0879(.A(men_men_n829_), .B(men_men_n113_), .Y(men_men_n908_));
  NA2        u0880(.A(men_men_n908_), .B(men_men_n907_), .Y(men_men_n909_));
  NA4        u0881(.A(men_men_n909_), .B(men_men_n905_), .C(men_men_n902_), .D(men_men_n897_), .Y(men_men_n910_));
  NO4        u0882(.A(men_men_n910_), .B(men_men_n893_), .C(men_men_n877_), .D(men_men_n864_), .Y(men_men_n911_));
  OR2        u0883(.A(men_men_n889_), .B(men_men_n75_), .Y(men_men_n912_));
  NA2        u0884(.A(men_men_n114_), .B(j), .Y(men_men_n913_));
  NA2        u0885(.A(men_men_n851_), .B(g), .Y(men_men_n914_));
  AOI210     u0886(.A0(men_men_n914_), .A1(men_men_n293_), .B0(men_men_n912_), .Y(men_men_n915_));
  NO2        u0887(.A(men_men_n335_), .B(men_men_n861_), .Y(men_men_n916_));
  NO2        u0888(.A(men_men_n234_), .B(men_men_n228_), .Y(men_men_n917_));
  NA2        u0889(.A(men_men_n917_), .B(men_men_n231_), .Y(men_men_n918_));
  NO2        u0890(.A(men_men_n436_), .B(men_men_n850_), .Y(men_men_n919_));
  NA2        u0891(.A(men_men_n919_), .B(men_men_n570_), .Y(men_men_n920_));
  NA2        u0892(.A(men_men_n920_), .B(men_men_n918_), .Y(men_men_n921_));
  NA2        u0893(.A(e), .B(d), .Y(men_men_n922_));
  OAI220     u0894(.A0(men_men_n922_), .A1(c), .B0(men_men_n325_), .B1(d), .Y(men_men_n923_));
  NA3        u0895(.A(men_men_n923_), .B(men_men_n459_), .C(men_men_n517_), .Y(men_men_n924_));
  AOI210     u0896(.A0(men_men_n524_), .A1(men_men_n181_), .B0(men_men_n234_), .Y(men_men_n925_));
  AOI210     u0897(.A0(men_men_n632_), .A1(men_men_n351_), .B0(men_men_n925_), .Y(men_men_n926_));
  NA2        u0898(.A(men_men_n285_), .B(men_men_n164_), .Y(men_men_n927_));
  NA2        u0899(.A(men_men_n890_), .B(men_men_n927_), .Y(men_men_n928_));
  NA3        u0900(.A(men_men_n167_), .B(men_men_n87_), .C(men_men_n34_), .Y(men_men_n929_));
  NA4        u0901(.A(men_men_n929_), .B(men_men_n928_), .C(men_men_n926_), .D(men_men_n924_), .Y(men_men_n930_));
  NO4        u0902(.A(men_men_n930_), .B(men_men_n921_), .C(men_men_n916_), .D(men_men_n915_), .Y(men_men_n931_));
  NA2        u0903(.A(men_men_n865_), .B(men_men_n31_), .Y(men_men_n932_));
  AO210      u0904(.A0(men_men_n932_), .A1(men_men_n715_), .B0(men_men_n220_), .Y(men_men_n933_));
  OAI220     u0905(.A0(men_men_n631_), .A1(men_men_n61_), .B0(men_men_n301_), .B1(j), .Y(men_men_n934_));
  AOI220     u0906(.A0(men_men_n934_), .A1(men_men_n895_), .B0(men_men_n621_), .B1(men_men_n630_), .Y(men_men_n935_));
  OAI210     u0907(.A0(men_men_n856_), .A1(men_men_n171_), .B0(men_men_n935_), .Y(men_men_n936_));
  OAI210     u0908(.A0(men_men_n851_), .A1(men_men_n927_), .B0(men_men_n883_), .Y(men_men_n937_));
  NO2        u0909(.A(men_men_n937_), .B(men_men_n613_), .Y(men_men_n938_));
  AOI210     u0910(.A0(men_men_n119_), .A1(men_men_n118_), .B0(men_men_n262_), .Y(men_men_n939_));
  NO2        u0911(.A(men_men_n939_), .B(men_men_n884_), .Y(men_men_n940_));
  AO210      u0912(.A0(men_men_n870_), .A1(men_men_n860_), .B0(men_men_n940_), .Y(men_men_n941_));
  NOi31      u0913(.An(men_men_n553_), .B(men_men_n881_), .C(men_men_n293_), .Y(men_men_n942_));
  NO4        u0914(.A(men_men_n942_), .B(men_men_n941_), .C(men_men_n938_), .D(men_men_n936_), .Y(men_men_n943_));
  AO220      u0915(.A0(men_men_n459_), .A1(men_men_n764_), .B0(men_men_n176_), .B1(f), .Y(men_men_n944_));
  OAI210     u0916(.A0(men_men_n944_), .A1(men_men_n462_), .B0(men_men_n923_), .Y(men_men_n945_));
  NO2        u0917(.A(men_men_n446_), .B(men_men_n71_), .Y(men_men_n946_));
  OAI210     u0918(.A0(men_men_n863_), .A1(men_men_n946_), .B0(men_men_n719_), .Y(men_men_n947_));
  AN4        u0919(.A(men_men_n947_), .B(men_men_n945_), .C(men_men_n943_), .D(men_men_n933_), .Y(men_men_n948_));
  NA4        u0920(.A(men_men_n948_), .B(men_men_n931_), .C(men_men_n911_), .D(men_men_n858_), .Y(men12));
  NO2        u0921(.A(men_men_n457_), .B(c), .Y(men_men_n950_));
  NO4        u0922(.A(men_men_n449_), .B(men_men_n255_), .C(men_men_n590_), .D(men_men_n217_), .Y(men_men_n951_));
  NA2        u0923(.A(men_men_n951_), .B(men_men_n950_), .Y(men_men_n952_));
  NA2        u0924(.A(men_men_n553_), .B(men_men_n946_), .Y(men_men_n953_));
  NO2        u0925(.A(men_men_n457_), .B(men_men_n117_), .Y(men_men_n954_));
  NO2        u0926(.A(men_men_n866_), .B(men_men_n358_), .Y(men_men_n955_));
  NO2        u0927(.A(men_men_n672_), .B(men_men_n385_), .Y(men_men_n956_));
  AOI220     u0928(.A0(men_men_n956_), .A1(men_men_n551_), .B0(men_men_n955_), .B1(men_men_n954_), .Y(men_men_n957_));
  NA4        u0929(.A(men_men_n957_), .B(men_men_n953_), .C(men_men_n952_), .D(men_men_n448_), .Y(men_men_n958_));
  AOI210     u0930(.A0(men_men_n237_), .A1(men_men_n341_), .B0(men_men_n203_), .Y(men_men_n959_));
  OR2        u0931(.A(men_men_n959_), .B(men_men_n951_), .Y(men_men_n960_));
  AOI210     u0932(.A0(men_men_n338_), .A1(men_men_n397_), .B0(men_men_n217_), .Y(men_men_n961_));
  OAI210     u0933(.A0(men_men_n961_), .A1(men_men_n960_), .B0(men_men_n409_), .Y(men_men_n962_));
  NO2        u0934(.A(men_men_n651_), .B(men_men_n264_), .Y(men_men_n963_));
  NO2        u0935(.A(men_men_n597_), .B(men_men_n859_), .Y(men_men_n964_));
  NO2        u0936(.A(men_men_n149_), .B(men_men_n241_), .Y(men_men_n965_));
  INV        u0937(.A(men_men_n962_), .Y(men_men_n966_));
  OR2        u0938(.A(men_men_n326_), .B(men_men_n954_), .Y(men_men_n967_));
  NA2        u0939(.A(men_men_n967_), .B(men_men_n359_), .Y(men_men_n968_));
  NA4        u0940(.A(men_men_n450_), .B(men_men_n444_), .C(men_men_n182_), .D(g), .Y(men_men_n969_));
  NA2        u0941(.A(men_men_n969_), .B(men_men_n968_), .Y(men_men_n970_));
  NO3        u0942(.A(men_men_n677_), .B(men_men_n94_), .C(men_men_n45_), .Y(men_men_n971_));
  NO4        u0943(.A(men_men_n971_), .B(men_men_n970_), .C(men_men_n966_), .D(men_men_n958_), .Y(men_men_n972_));
  NO2        u0944(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n973_));
  NA2        u0945(.A(men_men_n594_), .B(men_men_n73_), .Y(men_men_n974_));
  NA2        u0946(.A(men_men_n563_), .B(men_men_n143_), .Y(men_men_n975_));
  NOi21      u0947(.An(men_men_n34_), .B(men_men_n665_), .Y(men_men_n976_));
  AOI220     u0948(.A0(men_men_n976_), .A1(men_men_n975_), .B0(men_men_n974_), .B1(men_men_n973_), .Y(men_men_n977_));
  OAI210     u0949(.A0(men_men_n254_), .A1(men_men_n45_), .B0(men_men_n977_), .Y(men_men_n978_));
  NA2        u0950(.A(men_men_n442_), .B(men_men_n266_), .Y(men_men_n979_));
  NO3        u0951(.A(men_men_n838_), .B(men_men_n91_), .C(men_men_n414_), .Y(men_men_n980_));
  NAi31      u0952(.An(men_men_n980_), .B(men_men_n979_), .C(men_men_n322_), .Y(men_men_n981_));
  NO2        u0953(.A(men_men_n49_), .B(men_men_n45_), .Y(men_men_n982_));
  NO2        u0954(.A(men_men_n513_), .B(men_men_n301_), .Y(men_men_n983_));
  INV        u0955(.A(men_men_n983_), .Y(men_men_n984_));
  NO2        u0956(.A(men_men_n984_), .B(men_men_n143_), .Y(men_men_n985_));
  NA2        u0957(.A(men_men_n642_), .B(men_men_n368_), .Y(men_men_n986_));
  OAI210     u0958(.A0(men_men_n754_), .A1(men_men_n986_), .B0(men_men_n372_), .Y(men_men_n987_));
  NO4        u0959(.A(men_men_n987_), .B(men_men_n985_), .C(men_men_n981_), .D(men_men_n978_), .Y(men_men_n988_));
  NA2        u0960(.A(men_men_n351_), .B(g), .Y(men_men_n989_));
  NA2        u0961(.A(men_men_n161_), .B(i), .Y(men_men_n990_));
  NA2        u0962(.A(men_men_n46_), .B(i), .Y(men_men_n991_));
  OAI220     u0963(.A0(men_men_n991_), .A1(men_men_n202_), .B0(men_men_n990_), .B1(men_men_n94_), .Y(men_men_n992_));
  AOI210     u0964(.A0(men_men_n425_), .A1(men_men_n37_), .B0(men_men_n992_), .Y(men_men_n993_));
  NO2        u0965(.A(men_men_n143_), .B(men_men_n86_), .Y(men_men_n994_));
  OR2        u0966(.A(men_men_n994_), .B(men_men_n562_), .Y(men_men_n995_));
  NA2        u0967(.A(men_men_n563_), .B(men_men_n389_), .Y(men_men_n996_));
  AOI210     u0968(.A0(men_men_n996_), .A1(n), .B0(men_men_n995_), .Y(men_men_n997_));
  OAI220     u0969(.A0(men_men_n997_), .A1(men_men_n989_), .B0(men_men_n993_), .B1(men_men_n335_), .Y(men_men_n998_));
  NO2        u0970(.A(men_men_n672_), .B(men_men_n507_), .Y(men_men_n999_));
  NA3        u0971(.A(men_men_n346_), .B(men_men_n637_), .C(i), .Y(men_men_n1000_));
  OAI210     u0972(.A0(men_men_n446_), .A1(men_men_n311_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  OAI220     u0973(.A0(men_men_n1001_), .A1(men_men_n999_), .B0(men_men_n691_), .B1(men_men_n776_), .Y(men_men_n1002_));
  NA2        u0974(.A(men_men_n615_), .B(men_men_n115_), .Y(men_men_n1003_));
  OR3        u0975(.A(men_men_n311_), .B(men_men_n441_), .C(f), .Y(men_men_n1004_));
  NA3        u0976(.A(men_men_n637_), .B(men_men_n82_), .C(i), .Y(men_men_n1005_));
  OA220      u0977(.A0(men_men_n1005_), .A1(men_men_n1003_), .B0(men_men_n1004_), .B1(men_men_n596_), .Y(men_men_n1006_));
  NA3        u0978(.A(men_men_n327_), .B(men_men_n119_), .C(g), .Y(men_men_n1007_));
  AOI210     u0979(.A0(men_men_n688_), .A1(men_men_n1007_), .B0(m), .Y(men_men_n1008_));
  OAI210     u0980(.A0(men_men_n1008_), .A1(men_men_n955_), .B0(men_men_n326_), .Y(men_men_n1009_));
  NA2        u0981(.A(men_men_n706_), .B(men_men_n898_), .Y(men_men_n1010_));
  NA2        u0982(.A(men_men_n861_), .B(men_men_n447_), .Y(men_men_n1011_));
  NA2        u0983(.A(men_men_n225_), .B(men_men_n79_), .Y(men_men_n1012_));
  NA3        u0984(.A(men_men_n1012_), .B(men_men_n1005_), .C(men_men_n1004_), .Y(men_men_n1013_));
  AOI220     u0985(.A0(men_men_n1013_), .A1(men_men_n261_), .B0(men_men_n1011_), .B1(men_men_n1010_), .Y(men_men_n1014_));
  NA4        u0986(.A(men_men_n1014_), .B(men_men_n1009_), .C(men_men_n1006_), .D(men_men_n1002_), .Y(men_men_n1015_));
  NO2        u0987(.A(men_men_n385_), .B(men_men_n93_), .Y(men_men_n1016_));
  OAI210     u0988(.A0(men_men_n1016_), .A1(men_men_n963_), .B0(men_men_n242_), .Y(men_men_n1017_));
  NA2        u0989(.A(men_men_n676_), .B(men_men_n90_), .Y(men_men_n1018_));
  NO2        u0990(.A(men_men_n465_), .B(men_men_n217_), .Y(men_men_n1019_));
  AOI220     u0991(.A0(men_men_n1019_), .A1(men_men_n390_), .B0(men_men_n967_), .B1(men_men_n221_), .Y(men_men_n1020_));
  AOI220     u0992(.A0(men_men_n956_), .A1(men_men_n965_), .B0(men_men_n595_), .B1(men_men_n92_), .Y(men_men_n1021_));
  NA4        u0993(.A(men_men_n1021_), .B(men_men_n1020_), .C(men_men_n1018_), .D(men_men_n1017_), .Y(men_men_n1022_));
  OAI210     u0994(.A0(men_men_n1011_), .A1(men_men_n964_), .B0(men_men_n551_), .Y(men_men_n1023_));
  AOI210     u0995(.A0(men_men_n426_), .A1(men_men_n418_), .B0(men_men_n838_), .Y(men_men_n1024_));
  INV        u0996(.A(men_men_n1024_), .Y(men_men_n1025_));
  NA2        u0997(.A(men_men_n1008_), .B(men_men_n954_), .Y(men_men_n1026_));
  NO3        u0998(.A(men_men_n913_), .B(men_men_n49_), .C(men_men_n45_), .Y(men_men_n1027_));
  AOI220     u0999(.A0(men_men_n1027_), .A1(men_men_n635_), .B0(men_men_n656_), .B1(men_men_n540_), .Y(men_men_n1028_));
  NA4        u1000(.A(men_men_n1028_), .B(men_men_n1026_), .C(men_men_n1025_), .D(men_men_n1023_), .Y(men_men_n1029_));
  NO4        u1001(.A(men_men_n1029_), .B(men_men_n1022_), .C(men_men_n1015_), .D(men_men_n998_), .Y(men_men_n1030_));
  NAi31      u1002(.An(men_men_n140_), .B(men_men_n427_), .C(n), .Y(men_men_n1031_));
  NO3        u1003(.A(men_men_n127_), .B(men_men_n344_), .C(men_men_n867_), .Y(men_men_n1032_));
  NO2        u1004(.A(men_men_n1032_), .B(men_men_n1031_), .Y(men_men_n1033_));
  NO3        u1005(.A(men_men_n272_), .B(men_men_n140_), .C(men_men_n414_), .Y(men_men_n1034_));
  AOI210     u1006(.A0(men_men_n1034_), .A1(men_men_n508_), .B0(men_men_n1033_), .Y(men_men_n1035_));
  NA2        u1007(.A(men_men_n501_), .B(i), .Y(men_men_n1036_));
  NA2        u1008(.A(men_men_n1036_), .B(men_men_n1035_), .Y(men_men_n1037_));
  NA2        u1009(.A(men_men_n234_), .B(men_men_n172_), .Y(men_men_n1038_));
  NO3        u1010(.A(men_men_n308_), .B(men_men_n450_), .C(men_men_n176_), .Y(men_men_n1039_));
  NOi31      u1011(.An(men_men_n1038_), .B(men_men_n1039_), .C(men_men_n217_), .Y(men_men_n1040_));
  NAi21      u1012(.An(men_men_n563_), .B(men_men_n1019_), .Y(men_men_n1041_));
  NA2        u1013(.A(men_men_n445_), .B(men_men_n898_), .Y(men_men_n1042_));
  NO3        u1014(.A(men_men_n446_), .B(men_men_n311_), .C(men_men_n75_), .Y(men_men_n1043_));
  AOI220     u1015(.A0(men_men_n1043_), .A1(men_men_n1042_), .B0(men_men_n490_), .B1(g), .Y(men_men_n1044_));
  NA2        u1016(.A(men_men_n1044_), .B(men_men_n1041_), .Y(men_men_n1045_));
  NO2        u1017(.A(men_men_n1000_), .B(men_men_n611_), .Y(men_men_n1046_));
  NO2        u1018(.A(men_men_n673_), .B(men_men_n385_), .Y(men_men_n1047_));
  NA2        u1019(.A(men_men_n959_), .B(men_men_n950_), .Y(men_men_n1048_));
  NO3        u1020(.A(men_men_n552_), .B(men_men_n147_), .C(men_men_n216_), .Y(men_men_n1049_));
  OAI210     u1021(.A0(men_men_n1049_), .A1(men_men_n534_), .B0(men_men_n386_), .Y(men_men_n1050_));
  OAI220     u1022(.A0(men_men_n956_), .A1(men_men_n964_), .B0(men_men_n553_), .B1(men_men_n435_), .Y(men_men_n1051_));
  NA4        u1023(.A(men_men_n1051_), .B(men_men_n1050_), .C(men_men_n1048_), .D(men_men_n629_), .Y(men_men_n1052_));
  OAI210     u1024(.A0(men_men_n959_), .A1(men_men_n951_), .B0(men_men_n1038_), .Y(men_men_n1053_));
  NA3        u1025(.A(men_men_n996_), .B(men_men_n495_), .C(men_men_n46_), .Y(men_men_n1054_));
  AOI210     u1026(.A0(men_men_n388_), .A1(men_men_n386_), .B0(men_men_n334_), .Y(men_men_n1055_));
  NA3        u1027(.A(men_men_n1055_), .B(men_men_n1054_), .C(men_men_n1053_), .Y(men_men_n1056_));
  OR4        u1028(.A(men_men_n1056_), .B(men_men_n1052_), .C(men_men_n1047_), .D(men_men_n1046_), .Y(men_men_n1057_));
  NO4        u1029(.A(men_men_n1057_), .B(men_men_n1045_), .C(men_men_n1040_), .D(men_men_n1037_), .Y(men_men_n1058_));
  NA4        u1030(.A(men_men_n1058_), .B(men_men_n1030_), .C(men_men_n988_), .D(men_men_n972_), .Y(men13));
  AN2        u1031(.A(c), .B(b), .Y(men_men_n1060_));
  NA3        u1032(.A(men_men_n253_), .B(men_men_n1060_), .C(m), .Y(men_men_n1061_));
  NA2        u1033(.A(men_men_n506_), .B(f), .Y(men_men_n1062_));
  NO4        u1034(.A(men_men_n1062_), .B(men_men_n1061_), .C(j), .D(men_men_n591_), .Y(men_men_n1063_));
  NA2        u1035(.A(men_men_n266_), .B(men_men_n1060_), .Y(men_men_n1064_));
  NO4        u1036(.A(men_men_n1064_), .B(men_men_n1062_), .C(men_men_n990_), .D(a), .Y(men_men_n1065_));
  NAi32      u1037(.An(d), .Bn(c), .C(e), .Y(men_men_n1066_));
  NA2        u1038(.A(men_men_n139_), .B(men_men_n45_), .Y(men_men_n1067_));
  NO4        u1039(.A(men_men_n1067_), .B(men_men_n1066_), .C(men_men_n597_), .D(men_men_n307_), .Y(men_men_n1068_));
  NA2        u1040(.A(men_men_n680_), .B(men_men_n228_), .Y(men_men_n1069_));
  NA2        u1041(.A(men_men_n417_), .B(men_men_n216_), .Y(men_men_n1070_));
  AN2        u1042(.A(d), .B(c), .Y(men_men_n1071_));
  NA2        u1043(.A(men_men_n1071_), .B(men_men_n117_), .Y(men_men_n1072_));
  NO4        u1044(.A(men_men_n1072_), .B(men_men_n1070_), .C(men_men_n177_), .D(men_men_n168_), .Y(men_men_n1073_));
  NA2        u1045(.A(men_men_n506_), .B(c), .Y(men_men_n1074_));
  NO4        u1046(.A(men_men_n1067_), .B(men_men_n593_), .C(men_men_n1074_), .D(men_men_n307_), .Y(men_men_n1075_));
  AO210      u1047(.A0(men_men_n1073_), .A1(men_men_n1069_), .B0(men_men_n1075_), .Y(men_men_n1076_));
  OR4        u1048(.A(men_men_n1076_), .B(men_men_n1068_), .C(men_men_n1065_), .D(men_men_n1063_), .Y(men_men_n1077_));
  NAi32      u1049(.An(f), .Bn(e), .C(c), .Y(men_men_n1078_));
  NO2        u1050(.A(men_men_n1078_), .B(men_men_n144_), .Y(men_men_n1079_));
  NA2        u1051(.A(men_men_n1079_), .B(g), .Y(men_men_n1080_));
  OR3        u1052(.A(men_men_n228_), .B(men_men_n177_), .C(men_men_n168_), .Y(men_men_n1081_));
  NO2        u1053(.A(men_men_n1081_), .B(men_men_n1080_), .Y(men_men_n1082_));
  NO2        u1054(.A(men_men_n1074_), .B(men_men_n307_), .Y(men_men_n1083_));
  NO2        u1055(.A(j), .B(men_men_n45_), .Y(men_men_n1084_));
  NA2        u1056(.A(men_men_n639_), .B(men_men_n1084_), .Y(men_men_n1085_));
  NOi21      u1057(.An(men_men_n1083_), .B(men_men_n1085_), .Y(men_men_n1086_));
  NO2        u1058(.A(men_men_n780_), .B(men_men_n114_), .Y(men_men_n1087_));
  NOi41      u1059(.An(n), .B(m), .C(i), .D(h), .Y(men_men_n1088_));
  NA2        u1060(.A(men_men_n1088_), .B(men_men_n1087_), .Y(men_men_n1089_));
  NO2        u1061(.A(men_men_n1089_), .B(men_men_n1080_), .Y(men_men_n1090_));
  NA3        u1062(.A(k), .B(j), .C(i), .Y(men_men_n1091_));
  NO3        u1063(.A(men_men_n1091_), .B(men_men_n307_), .C(men_men_n93_), .Y(men_men_n1092_));
  OR3        u1064(.A(men_men_n1090_), .B(men_men_n1086_), .C(men_men_n1082_), .Y(men_men_n1093_));
  NA3        u1065(.A(men_men_n473_), .B(men_men_n337_), .C(men_men_n56_), .Y(men_men_n1094_));
  NO2        u1066(.A(men_men_n1094_), .B(men_men_n1085_), .Y(men_men_n1095_));
  NO4        u1067(.A(men_men_n1094_), .B(men_men_n593_), .C(men_men_n456_), .D(men_men_n45_), .Y(men_men_n1096_));
  NO2        u1068(.A(f), .B(c), .Y(men_men_n1097_));
  NOi21      u1069(.An(men_men_n1097_), .B(men_men_n449_), .Y(men_men_n1098_));
  NA2        u1070(.A(men_men_n1098_), .B(men_men_n59_), .Y(men_men_n1099_));
  OR2        u1071(.A(men_men_n1096_), .B(men_men_n1095_), .Y(men_men_n1100_));
  OR3        u1072(.A(men_men_n1100_), .B(men_men_n1093_), .C(men_men_n1077_), .Y(men02));
  OR3        u1073(.A(n), .B(m), .C(i), .Y(men_men_n1102_));
  NOi31      u1074(.An(e), .B(d), .C(c), .Y(men_men_n1103_));
  AOI210     u1075(.A0(men_men_n1092_), .A1(men_men_n1103_), .B0(men_men_n1068_), .Y(men_men_n1104_));
  AN3        u1076(.A(g), .B(f), .C(c), .Y(men_men_n1105_));
  NA3        u1077(.A(men_men_n1105_), .B(men_men_n473_), .C(h), .Y(men_men_n1106_));
  OR2        u1078(.A(men_men_n1091_), .B(men_men_n307_), .Y(men_men_n1107_));
  OR2        u1079(.A(men_men_n1107_), .B(men_men_n1106_), .Y(men_men_n1108_));
  NO3        u1080(.A(men_men_n1094_), .B(men_men_n1067_), .C(men_men_n593_), .Y(men_men_n1109_));
  NO2        u1081(.A(men_men_n1109_), .B(men_men_n1082_), .Y(men_men_n1110_));
  NA3        u1082(.A(l), .B(k), .C(j), .Y(men_men_n1111_));
  NA2        u1083(.A(i), .B(h), .Y(men_men_n1112_));
  NO3        u1084(.A(men_men_n1112_), .B(men_men_n1111_), .C(men_men_n131_), .Y(men_men_n1113_));
  NO3        u1085(.A(men_men_n141_), .B(men_men_n283_), .C(men_men_n217_), .Y(men_men_n1114_));
  AOI210     u1086(.A0(men_men_n1114_), .A1(men_men_n1113_), .B0(men_men_n1086_), .Y(men_men_n1115_));
  NA3        u1087(.A(c), .B(b), .C(a), .Y(men_men_n1116_));
  NO3        u1088(.A(men_men_n1116_), .B(men_men_n922_), .C(men_men_n216_), .Y(men_men_n1117_));
  NO3        u1089(.A(men_men_n1091_), .B(men_men_n49_), .C(men_men_n114_), .Y(men_men_n1118_));
  AOI210     u1090(.A0(men_men_n1118_), .A1(men_men_n1117_), .B0(men_men_n1095_), .Y(men_men_n1119_));
  AN4        u1091(.A(men_men_n1119_), .B(men_men_n1115_), .C(men_men_n1110_), .D(men_men_n1108_), .Y(men_men_n1120_));
  NO2        u1092(.A(men_men_n1072_), .B(men_men_n1070_), .Y(men_men_n1121_));
  NA2        u1093(.A(men_men_n1089_), .B(men_men_n1081_), .Y(men_men_n1122_));
  AOI210     u1094(.A0(men_men_n1122_), .A1(men_men_n1121_), .B0(men_men_n1063_), .Y(men_men_n1123_));
  NA3        u1095(.A(men_men_n1123_), .B(men_men_n1120_), .C(men_men_n1104_), .Y(men03));
  NA4        u1096(.A(men_men_n90_), .B(men_men_n89_), .C(g), .D(men_men_n216_), .Y(men_men_n1125_));
  NA4        u1097(.A(men_men_n582_), .B(m), .C(men_men_n114_), .D(men_men_n216_), .Y(men_men_n1126_));
  NA3        u1098(.A(men_men_n1126_), .B(men_men_n376_), .C(men_men_n1125_), .Y(men_men_n1127_));
  INV        u1099(.A(men_men_n1127_), .Y(men_men_n1128_));
  NOi31      u1100(.An(men_men_n827_), .B(men_men_n872_), .C(men_men_n862_), .Y(men_men_n1129_));
  OAI220     u1101(.A0(men_men_n1129_), .A1(men_men_n706_), .B0(men_men_n1128_), .B1(men_men_n594_), .Y(men_men_n1130_));
  NOi31      u1102(.An(i), .B(k), .C(j), .Y(men_men_n1131_));
  NA4        u1103(.A(men_men_n1131_), .B(men_men_n1103_), .C(men_men_n346_), .D(men_men_n337_), .Y(men_men_n1132_));
  OAI210     u1104(.A0(men_men_n838_), .A1(men_men_n428_), .B0(men_men_n1132_), .Y(men_men_n1133_));
  NOi31      u1105(.An(m), .B(n), .C(f), .Y(men_men_n1134_));
  NA2        u1106(.A(men_men_n1134_), .B(men_men_n51_), .Y(men_men_n1135_));
  AN2        u1107(.A(e), .B(c), .Y(men_men_n1136_));
  NA2        u1108(.A(men_men_n1136_), .B(a), .Y(men_men_n1137_));
  OAI220     u1109(.A0(men_men_n1137_), .A1(men_men_n1135_), .B0(men_men_n906_), .B1(men_men_n434_), .Y(men_men_n1138_));
  NA2        u1110(.A(men_men_n517_), .B(l), .Y(men_men_n1139_));
  NOi31      u1111(.An(men_men_n883_), .B(men_men_n1061_), .C(men_men_n1139_), .Y(men_men_n1140_));
  NO4        u1112(.A(men_men_n1140_), .B(men_men_n1138_), .C(men_men_n1133_), .D(men_men_n1024_), .Y(men_men_n1141_));
  NO2        u1113(.A(men_men_n283_), .B(a), .Y(men_men_n1142_));
  INV        u1114(.A(men_men_n1068_), .Y(men_men_n1143_));
  NO2        u1115(.A(men_men_n1112_), .B(men_men_n493_), .Y(men_men_n1144_));
  NO2        u1116(.A(men_men_n89_), .B(g), .Y(men_men_n1145_));
  NA2        u1117(.A(men_men_n1145_), .B(men_men_n1144_), .Y(men_men_n1146_));
  OR2        u1118(.A(men_men_n1146_), .B(men_men_n1099_), .Y(men_men_n1147_));
  NA3        u1119(.A(men_men_n1147_), .B(men_men_n1143_), .C(men_men_n1141_), .Y(men_men_n1148_));
  NO4        u1120(.A(men_men_n1148_), .B(men_men_n1130_), .C(men_men_n839_), .D(men_men_n572_), .Y(men_men_n1149_));
  NA2        u1121(.A(c), .B(b), .Y(men_men_n1150_));
  NO2        u1122(.A(men_men_n718_), .B(men_men_n1150_), .Y(men_men_n1151_));
  OAI210     u1123(.A0(men_men_n881_), .A1(men_men_n854_), .B0(men_men_n421_), .Y(men_men_n1152_));
  OAI210     u1124(.A0(men_men_n1152_), .A1(men_men_n882_), .B0(men_men_n1151_), .Y(men_men_n1153_));
  NAi21      u1125(.An(men_men_n429_), .B(men_men_n1151_), .Y(men_men_n1154_));
  OAI210     u1126(.A0(men_men_n557_), .A1(men_men_n39_), .B0(men_men_n1142_), .Y(men_men_n1155_));
  NA2        u1127(.A(men_men_n1155_), .B(men_men_n1154_), .Y(men_men_n1156_));
  NA2        u1128(.A(men_men_n263_), .B(men_men_n120_), .Y(men_men_n1157_));
  OAI210     u1129(.A0(men_men_n1157_), .A1(men_men_n287_), .B0(g), .Y(men_men_n1158_));
  NAi21      u1130(.An(f), .B(d), .Y(men_men_n1159_));
  NO2        u1131(.A(men_men_n1159_), .B(men_men_n1116_), .Y(men_men_n1160_));
  INV        u1132(.A(men_men_n1160_), .Y(men_men_n1161_));
  AOI210     u1133(.A0(men_men_n1158_), .A1(men_men_n293_), .B0(men_men_n1161_), .Y(men_men_n1162_));
  AOI210     u1134(.A0(men_men_n1162_), .A1(men_men_n115_), .B0(men_men_n1156_), .Y(men_men_n1163_));
  NA2        u1135(.A(men_men_n476_), .B(men_men_n475_), .Y(men_men_n1164_));
  NO2        u1136(.A(men_men_n183_), .B(men_men_n241_), .Y(men_men_n1165_));
  NA2        u1137(.A(men_men_n1165_), .B(m), .Y(men_men_n1166_));
  NA3        u1138(.A(men_men_n939_), .B(men_men_n1139_), .C(men_men_n479_), .Y(men_men_n1167_));
  OAI210     u1139(.A0(men_men_n1167_), .A1(men_men_n312_), .B0(men_men_n477_), .Y(men_men_n1168_));
  AOI210     u1140(.A0(men_men_n1168_), .A1(men_men_n1164_), .B0(men_men_n1166_), .Y(men_men_n1169_));
  NA2        u1141(.A(men_men_n570_), .B(men_men_n416_), .Y(men_men_n1170_));
  NA2        u1142(.A(men_men_n157_), .B(men_men_n33_), .Y(men_men_n1171_));
  AOI210     u1143(.A0(men_men_n986_), .A1(men_men_n1171_), .B0(men_men_n217_), .Y(men_men_n1172_));
  OAI210     u1144(.A0(men_men_n1172_), .A1(men_men_n453_), .B0(men_men_n1160_), .Y(men_men_n1173_));
  NO2        u1145(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n1174_));
  AOI210     u1146(.A0(men_men_n1165_), .A1(men_men_n437_), .B0(men_men_n980_), .Y(men_men_n1175_));
  NAi41      u1147(.An(men_men_n1174_), .B(men_men_n1175_), .C(men_men_n1173_), .D(men_men_n1170_), .Y(men_men_n1176_));
  NO2        u1148(.A(men_men_n1176_), .B(men_men_n1169_), .Y(men_men_n1177_));
  NA4        u1149(.A(men_men_n1177_), .B(men_men_n1163_), .C(men_men_n1153_), .D(men_men_n1149_), .Y(men00));
  AOI210     u1150(.A0(men_men_n300_), .A1(men_men_n217_), .B0(men_men_n275_), .Y(men_men_n1179_));
  NO2        u1151(.A(men_men_n1179_), .B(men_men_n585_), .Y(men_men_n1180_));
  AOI210     u1152(.A0(men_men_n919_), .A1(men_men_n965_), .B0(men_men_n1133_), .Y(men_men_n1181_));
  NO3        u1153(.A(men_men_n1109_), .B(men_men_n980_), .C(men_men_n730_), .Y(men_men_n1182_));
  NA3        u1154(.A(men_men_n1182_), .B(men_men_n1181_), .C(men_men_n1025_), .Y(men_men_n1183_));
  NA2        u1155(.A(men_men_n519_), .B(f), .Y(men_men_n1184_));
  OAI210     u1156(.A0(men_men_n1032_), .A1(men_men_n40_), .B0(men_men_n658_), .Y(men_men_n1185_));
  NA3        u1157(.A(men_men_n1185_), .B(men_men_n260_), .C(n), .Y(men_men_n1186_));
  AOI210     u1158(.A0(men_men_n1186_), .A1(men_men_n1184_), .B0(men_men_n1072_), .Y(men_men_n1187_));
  NO4        u1159(.A(men_men_n1187_), .B(men_men_n1183_), .C(men_men_n1180_), .D(men_men_n1093_), .Y(men_men_n1188_));
  NA3        u1160(.A(men_men_n167_), .B(men_men_n46_), .C(men_men_n45_), .Y(men_men_n1189_));
  NA3        u1161(.A(d), .B(men_men_n56_), .C(b), .Y(men_men_n1190_));
  NOi31      u1162(.An(n), .B(m), .C(i), .Y(men_men_n1191_));
  NA3        u1163(.A(men_men_n1191_), .B(men_men_n661_), .C(men_men_n51_), .Y(men_men_n1192_));
  OAI210     u1164(.A0(men_men_n1190_), .A1(men_men_n1189_), .B0(men_men_n1192_), .Y(men_men_n1193_));
  INV        u1165(.A(men_men_n584_), .Y(men_men_n1194_));
  NO4        u1166(.A(men_men_n1194_), .B(men_men_n1193_), .C(men_men_n1174_), .D(men_men_n942_), .Y(men_men_n1195_));
  NO4        u1167(.A(men_men_n496_), .B(men_men_n361_), .C(men_men_n1150_), .D(men_men_n59_), .Y(men_men_n1196_));
  NA3        u1168(.A(men_men_n391_), .B(men_men_n224_), .C(g), .Y(men_men_n1197_));
  OA220      u1169(.A0(men_men_n1197_), .A1(men_men_n1190_), .B0(men_men_n392_), .B1(men_men_n134_), .Y(men_men_n1198_));
  NO2        u1170(.A(h), .B(g), .Y(men_men_n1199_));
  NA4        u1171(.A(men_men_n508_), .B(men_men_n473_), .C(men_men_n1199_), .D(men_men_n1060_), .Y(men_men_n1200_));
  OAI220     u1172(.A0(men_men_n536_), .A1(men_men_n605_), .B0(men_men_n94_), .B1(men_men_n93_), .Y(men_men_n1201_));
  NA2        u1173(.A(men_men_n1201_), .B(men_men_n544_), .Y(men_men_n1202_));
  NA3        u1174(.A(men_men_n1202_), .B(men_men_n1200_), .C(men_men_n1198_), .Y(men_men_n1203_));
  NO2        u1175(.A(men_men_n1203_), .B(men_men_n1196_), .Y(men_men_n1204_));
  INV        u1176(.A(men_men_n324_), .Y(men_men_n1205_));
  INV        u1177(.A(men_men_n586_), .Y(men_men_n1206_));
  NA3        u1178(.A(men_men_n1206_), .B(men_men_n1205_), .C(men_men_n152_), .Y(men_men_n1207_));
  NO2        u1179(.A(men_men_n243_), .B(men_men_n182_), .Y(men_men_n1208_));
  NA2        u1180(.A(men_men_n1208_), .B(men_men_n435_), .Y(men_men_n1209_));
  NA3        u1181(.A(men_men_n180_), .B(men_men_n114_), .C(g), .Y(men_men_n1210_));
  NA2        u1182(.A(men_men_n473_), .B(f), .Y(men_men_n1211_));
  NOi31      u1183(.An(men_men_n891_), .B(men_men_n1211_), .C(men_men_n1210_), .Y(men_men_n1212_));
  NAi31      u1184(.An(men_men_n187_), .B(men_men_n878_), .C(men_men_n473_), .Y(men_men_n1213_));
  NAi31      u1185(.An(men_men_n1212_), .B(men_men_n1213_), .C(men_men_n1209_), .Y(men_men_n1214_));
  NO2        u1186(.A(men_men_n274_), .B(men_men_n75_), .Y(men_men_n1215_));
  NO3        u1187(.A(men_men_n434_), .B(men_men_n850_), .C(n), .Y(men_men_n1216_));
  NA2        u1188(.A(men_men_n1216_), .B(men_men_n1215_), .Y(men_men_n1217_));
  NAi31      u1189(.An(men_men_n1075_), .B(men_men_n1217_), .C(men_men_n74_), .Y(men_men_n1218_));
  NO4        u1190(.A(men_men_n1218_), .B(men_men_n1214_), .C(men_men_n1207_), .D(men_men_n527_), .Y(men_men_n1219_));
  AN3        u1191(.A(men_men_n1219_), .B(men_men_n1204_), .C(men_men_n1195_), .Y(men_men_n1220_));
  NA3        u1192(.A(men_men_n1134_), .B(men_men_n615_), .C(men_men_n472_), .Y(men_men_n1221_));
  NA3        u1193(.A(men_men_n1221_), .B(men_men_n571_), .C(men_men_n246_), .Y(men_men_n1222_));
  NA2        u1194(.A(men_men_n1127_), .B(men_men_n544_), .Y(men_men_n1223_));
  NA2        u1195(.A(men_men_n1223_), .B(men_men_n297_), .Y(men_men_n1224_));
  OAI210     u1196(.A0(men_men_n471_), .A1(men_men_n121_), .B0(men_men_n884_), .Y(men_men_n1225_));
  AOI220     u1197(.A0(men_men_n1225_), .A1(men_men_n1167_), .B0(men_men_n570_), .B1(men_men_n416_), .Y(men_men_n1226_));
  OR4        u1198(.A(men_men_n1072_), .B(men_men_n272_), .C(men_men_n226_), .D(e), .Y(men_men_n1227_));
  NO2        u1199(.A(men_men_n220_), .B(men_men_n217_), .Y(men_men_n1228_));
  NA2        u1200(.A(n), .B(e), .Y(men_men_n1229_));
  NO2        u1201(.A(men_men_n1229_), .B(men_men_n144_), .Y(men_men_n1230_));
  AOI220     u1202(.A0(men_men_n1230_), .A1(men_men_n273_), .B0(men_men_n865_), .B1(men_men_n1228_), .Y(men_men_n1231_));
  OAI210     u1203(.A0(men_men_n362_), .A1(men_men_n313_), .B0(men_men_n455_), .Y(men_men_n1232_));
  NA4        u1204(.A(men_men_n1232_), .B(men_men_n1231_), .C(men_men_n1227_), .D(men_men_n1226_), .Y(men_men_n1233_));
  AOI210     u1205(.A0(men_men_n1230_), .A1(men_men_n869_), .B0(men_men_n839_), .Y(men_men_n1234_));
  AOI220     u1206(.A0(men_men_n976_), .A1(men_men_n583_), .B0(men_men_n661_), .B1(men_men_n249_), .Y(men_men_n1235_));
  NO2        u1207(.A(men_men_n68_), .B(h), .Y(men_men_n1236_));
  NO3        u1208(.A(men_men_n1072_), .B(men_men_n1070_), .C(men_men_n746_), .Y(men_men_n1237_));
  INV        u1209(.A(men_men_n131_), .Y(men_men_n1238_));
  AN2        u1210(.A(men_men_n1238_), .B(men_men_n1114_), .Y(men_men_n1239_));
  OAI210     u1211(.A0(men_men_n1239_), .A1(men_men_n1237_), .B0(men_men_n1236_), .Y(men_men_n1240_));
  NA4        u1212(.A(men_men_n1240_), .B(men_men_n1235_), .C(men_men_n1234_), .D(men_men_n886_), .Y(men_men_n1241_));
  NO4        u1213(.A(men_men_n1241_), .B(men_men_n1233_), .C(men_men_n1224_), .D(men_men_n1222_), .Y(men_men_n1242_));
  NA2        u1214(.A(men_men_n855_), .B(men_men_n775_), .Y(men_men_n1243_));
  NA4        u1215(.A(men_men_n1243_), .B(men_men_n1242_), .C(men_men_n1220_), .D(men_men_n1188_), .Y(men01));
  AN2        u1216(.A(men_men_n1050_), .B(men_men_n1048_), .Y(men_men_n1245_));
  NO4        u1217(.A(men_men_n823_), .B(men_men_n815_), .C(men_men_n487_), .D(men_men_n281_), .Y(men_men_n1246_));
  NA2        u1218(.A(men_men_n402_), .B(i), .Y(men_men_n1247_));
  NA3        u1219(.A(men_men_n1247_), .B(men_men_n1246_), .C(men_men_n1245_), .Y(men_men_n1248_));
  NA2        u1220(.A(men_men_n595_), .B(men_men_n92_), .Y(men_men_n1249_));
  NA2        u1221(.A(men_men_n563_), .B(men_men_n271_), .Y(men_men_n1250_));
  NA2        u1222(.A(men_men_n983_), .B(men_men_n1250_), .Y(men_men_n1251_));
  NA4        u1223(.A(men_men_n1251_), .B(men_men_n1249_), .C(men_men_n935_), .D(men_men_n336_), .Y(men_men_n1252_));
  NA2        u1224(.A(men_men_n45_), .B(f), .Y(men_men_n1253_));
  NA2        u1225(.A(men_men_n725_), .B(men_men_n99_), .Y(men_men_n1254_));
  NO2        u1226(.A(men_men_n1254_), .B(men_men_n1253_), .Y(men_men_n1255_));
  NO2        u1227(.A(men_men_n801_), .B(men_men_n611_), .Y(men_men_n1256_));
  AOI210     u1228(.A0(men_men_n1255_), .A1(men_men_n646_), .B0(men_men_n1256_), .Y(men_men_n1257_));
  INV        u1229(.A(men_men_n119_), .Y(men_men_n1258_));
  OR2        u1230(.A(men_men_n674_), .B(men_men_n376_), .Y(men_men_n1259_));
  NAi41      u1231(.An(men_men_n160_), .B(men_men_n1259_), .C(men_men_n1257_), .D(men_men_n918_), .Y(men_men_n1260_));
  NO3        u1232(.A(men_men_n802_), .B(men_men_n690_), .C(men_men_n522_), .Y(men_men_n1261_));
  NA4        u1233(.A(men_men_n725_), .B(men_men_n99_), .C(men_men_n45_), .D(men_men_n216_), .Y(men_men_n1262_));
  OA220      u1234(.A0(men_men_n1262_), .A1(men_men_n683_), .B0(men_men_n197_), .B1(men_men_n195_), .Y(men_men_n1263_));
  NA3        u1235(.A(men_men_n1263_), .B(men_men_n1261_), .C(men_men_n137_), .Y(men_men_n1264_));
  NO4        u1236(.A(men_men_n1264_), .B(men_men_n1260_), .C(men_men_n1252_), .D(men_men_n1248_), .Y(men_men_n1265_));
  INV        u1237(.A(men_men_n1197_), .Y(men_men_n1266_));
  NA2        u1238(.A(men_men_n1266_), .B(men_men_n540_), .Y(men_men_n1267_));
  AOI210     u1239(.A0(men_men_n206_), .A1(men_men_n91_), .B0(men_men_n216_), .Y(men_men_n1268_));
  OAI210     u1240(.A0(men_men_n830_), .A1(men_men_n435_), .B0(men_men_n1268_), .Y(men_men_n1269_));
  AN3        u1241(.A(m), .B(l), .C(k), .Y(men_men_n1270_));
  OAI210     u1242(.A0(men_men_n364_), .A1(men_men_n34_), .B0(men_men_n1270_), .Y(men_men_n1271_));
  NA2        u1243(.A(men_men_n205_), .B(men_men_n34_), .Y(men_men_n1272_));
  AO210      u1244(.A0(men_men_n1272_), .A1(men_men_n1271_), .B0(men_men_n335_), .Y(men_men_n1273_));
  NA3        u1245(.A(men_men_n1273_), .B(men_men_n1269_), .C(men_men_n1267_), .Y(men_men_n1274_));
  AOI210     u1246(.A0(men_men_n603_), .A1(men_men_n119_), .B0(men_men_n609_), .Y(men_men_n1275_));
  OAI210     u1247(.A0(men_men_n1258_), .A1(men_men_n600_), .B0(men_men_n1275_), .Y(men_men_n1276_));
  NA2        u1248(.A(men_men_n280_), .B(men_men_n197_), .Y(men_men_n1277_));
  NA2        u1249(.A(men_men_n1277_), .B(men_men_n679_), .Y(men_men_n1278_));
  NO3        u1250(.A(men_men_n838_), .B(men_men_n206_), .C(men_men_n414_), .Y(men_men_n1279_));
  NO2        u1251(.A(men_men_n1279_), .B(men_men_n980_), .Y(men_men_n1280_));
  OAI210     u1252(.A0(men_men_n1255_), .A1(men_men_n329_), .B0(men_men_n691_), .Y(men_men_n1281_));
  NA4        u1253(.A(men_men_n1281_), .B(men_men_n1280_), .C(men_men_n1278_), .D(men_men_n805_), .Y(men_men_n1282_));
  NO3        u1254(.A(men_men_n1282_), .B(men_men_n1276_), .C(men_men_n1274_), .Y(men_men_n1283_));
  NA3        u1255(.A(men_men_n612_), .B(men_men_n29_), .C(f), .Y(men_men_n1284_));
  NO2        u1256(.A(men_men_n1284_), .B(men_men_n206_), .Y(men_men_n1285_));
  AOI210     u1257(.A0(men_men_n514_), .A1(men_men_n58_), .B0(men_men_n1285_), .Y(men_men_n1286_));
  OR3        u1258(.A(men_men_n1254_), .B(men_men_n613_), .C(men_men_n1253_), .Y(men_men_n1287_));
  NO2        u1259(.A(men_men_n1262_), .B(men_men_n1003_), .Y(men_men_n1288_));
  NO2        u1260(.A(men_men_n209_), .B(men_men_n113_), .Y(men_men_n1289_));
  NO3        u1261(.A(men_men_n1289_), .B(men_men_n1288_), .C(men_men_n1193_), .Y(men_men_n1290_));
  NA4        u1262(.A(men_men_n1290_), .B(men_men_n1287_), .C(men_men_n1286_), .D(men_men_n774_), .Y(men_men_n1291_));
  NO2        u1263(.A(men_men_n990_), .B(men_men_n236_), .Y(men_men_n1292_));
  NO2        u1264(.A(men_men_n991_), .B(men_men_n565_), .Y(men_men_n1293_));
  OAI210     u1265(.A0(men_men_n1293_), .A1(men_men_n1292_), .B0(men_men_n344_), .Y(men_men_n1294_));
  NO3        u1266(.A(men_men_n81_), .B(men_men_n301_), .C(men_men_n45_), .Y(men_men_n1295_));
  NA2        u1267(.A(men_men_n1295_), .B(men_men_n562_), .Y(men_men_n1296_));
  NA2        u1268(.A(men_men_n1296_), .B(men_men_n685_), .Y(men_men_n1297_));
  OR2        u1269(.A(men_men_n1197_), .B(men_men_n1190_), .Y(men_men_n1298_));
  NO2        u1270(.A(men_men_n376_), .B(men_men_n73_), .Y(men_men_n1299_));
  INV        u1271(.A(men_men_n1299_), .Y(men_men_n1300_));
  NA2        u1272(.A(men_men_n1295_), .B(men_men_n833_), .Y(men_men_n1301_));
  NA4        u1273(.A(men_men_n1301_), .B(men_men_n1300_), .C(men_men_n1298_), .D(men_men_n394_), .Y(men_men_n1302_));
  NOi41      u1274(.An(men_men_n1294_), .B(men_men_n1302_), .C(men_men_n1297_), .D(men_men_n1291_), .Y(men_men_n1303_));
  NO2        u1275(.A(men_men_n130_), .B(men_men_n45_), .Y(men_men_n1304_));
  NO2        u1276(.A(men_men_n45_), .B(men_men_n40_), .Y(men_men_n1305_));
  AO220      u1277(.A0(men_men_n1305_), .A1(men_men_n632_), .B0(men_men_n1304_), .B1(men_men_n723_), .Y(men_men_n1306_));
  NA2        u1278(.A(men_men_n1306_), .B(men_men_n344_), .Y(men_men_n1307_));
  NO3        u1279(.A(men_men_n1112_), .B(men_men_n177_), .C(men_men_n89_), .Y(men_men_n1308_));
  NA2        u1280(.A(men_men_n1295_), .B(men_men_n994_), .Y(men_men_n1309_));
  NA2        u1281(.A(men_men_n1309_), .B(men_men_n1307_), .Y(men_men_n1310_));
  NO2        u1282(.A(men_men_n623_), .B(men_men_n622_), .Y(men_men_n1311_));
  NO4        u1283(.A(men_men_n1112_), .B(men_men_n1311_), .C(men_men_n175_), .D(men_men_n89_), .Y(men_men_n1312_));
  NO3        u1284(.A(men_men_n1312_), .B(men_men_n1310_), .C(men_men_n650_), .Y(men_men_n1313_));
  NA4        u1285(.A(men_men_n1313_), .B(men_men_n1303_), .C(men_men_n1283_), .D(men_men_n1265_), .Y(men06));
  NO2        u1286(.A(men_men_n415_), .B(men_men_n569_), .Y(men_men_n1315_));
  INV        u1287(.A(men_men_n753_), .Y(men_men_n1316_));
  OAI210     u1288(.A0(men_men_n1316_), .A1(men_men_n267_), .B0(men_men_n1315_), .Y(men_men_n1317_));
  NO2        u1289(.A(men_men_n228_), .B(men_men_n105_), .Y(men_men_n1318_));
  OAI210     u1290(.A0(men_men_n1318_), .A1(men_men_n1308_), .B0(men_men_n390_), .Y(men_men_n1319_));
  NO3        u1291(.A(men_men_n607_), .B(men_men_n828_), .C(men_men_n610_), .Y(men_men_n1320_));
  OR2        u1292(.A(men_men_n1320_), .B(men_men_n906_), .Y(men_men_n1321_));
  NA4        u1293(.A(men_men_n1321_), .B(men_men_n1319_), .C(men_men_n1317_), .D(men_men_n1294_), .Y(men_men_n1322_));
  NO3        u1294(.A(men_men_n1322_), .B(men_men_n1297_), .C(men_men_n259_), .Y(men_men_n1323_));
  NO2        u1295(.A(men_men_n301_), .B(men_men_n45_), .Y(men_men_n1324_));
  AOI210     u1296(.A0(men_men_n1324_), .A1(men_men_n995_), .B0(men_men_n1292_), .Y(men_men_n1325_));
  AOI210     u1297(.A0(men_men_n1324_), .A1(men_men_n566_), .B0(men_men_n1306_), .Y(men_men_n1326_));
  AOI210     u1298(.A0(men_men_n1326_), .A1(men_men_n1325_), .B0(men_men_n341_), .Y(men_men_n1327_));
  OAI210     u1299(.A0(men_men_n91_), .A1(men_men_n40_), .B0(men_men_n689_), .Y(men_men_n1328_));
  NA2        u1300(.A(men_men_n1328_), .B(men_men_n654_), .Y(men_men_n1329_));
  NO2        u1301(.A(men_men_n524_), .B(men_men_n172_), .Y(men_men_n1330_));
  NOi21      u1302(.An(men_men_n136_), .B(men_men_n45_), .Y(men_men_n1331_));
  NO2        u1303(.A(men_men_n616_), .B(men_men_n1135_), .Y(men_men_n1332_));
  OAI210     u1304(.A0(men_men_n466_), .A1(men_men_n252_), .B0(men_men_n929_), .Y(men_men_n1333_));
  NO4        u1305(.A(men_men_n1333_), .B(men_men_n1332_), .C(men_men_n1331_), .D(men_men_n1330_), .Y(men_men_n1334_));
  OR2        u1306(.A(men_men_n608_), .B(men_men_n606_), .Y(men_men_n1335_));
  NO2        u1307(.A(men_men_n375_), .B(men_men_n135_), .Y(men_men_n1336_));
  AOI210     u1308(.A0(men_men_n1336_), .A1(men_men_n595_), .B0(men_men_n1335_), .Y(men_men_n1337_));
  NA3        u1309(.A(men_men_n1337_), .B(men_men_n1334_), .C(men_men_n1329_), .Y(men_men_n1338_));
  NO2        u1310(.A(men_men_n765_), .B(men_men_n374_), .Y(men_men_n1339_));
  NO3        u1311(.A(men_men_n691_), .B(men_men_n776_), .C(men_men_n646_), .Y(men_men_n1340_));
  NOi21      u1312(.An(men_men_n1339_), .B(men_men_n1340_), .Y(men_men_n1341_));
  AN2        u1313(.A(men_men_n976_), .B(men_men_n657_), .Y(men_men_n1342_));
  NO4        u1314(.A(men_men_n1342_), .B(men_men_n1341_), .C(men_men_n1338_), .D(men_men_n1327_), .Y(men_men_n1343_));
  NO2        u1315(.A(men_men_n822_), .B(men_men_n276_), .Y(men_men_n1344_));
  OAI220     u1316(.A0(men_men_n753_), .A1(men_men_n47_), .B0(men_men_n228_), .B1(men_men_n625_), .Y(men_men_n1345_));
  OAI210     u1317(.A0(men_men_n276_), .A1(c), .B0(men_men_n653_), .Y(men_men_n1346_));
  AOI220     u1318(.A0(men_men_n1346_), .A1(men_men_n1345_), .B0(men_men_n1344_), .B1(men_men_n267_), .Y(men_men_n1347_));
  NO3        u1319(.A(men_men_n248_), .B(men_men_n105_), .C(men_men_n283_), .Y(men_men_n1348_));
  OAI220     u1320(.A0(men_men_n715_), .A1(men_men_n252_), .B0(men_men_n521_), .B1(men_men_n524_), .Y(men_men_n1349_));
  OAI210     u1321(.A0(l), .A1(i), .B0(k), .Y(men_men_n1350_));
  NO3        u1322(.A(men_men_n1350_), .B(men_men_n605_), .C(j), .Y(men_men_n1351_));
  NOi21      u1323(.An(men_men_n1351_), .B(men_men_n683_), .Y(men_men_n1352_));
  NO4        u1324(.A(men_men_n1352_), .B(men_men_n1349_), .C(men_men_n1348_), .D(men_men_n1138_), .Y(men_men_n1353_));
  NA3        u1325(.A(men_men_n813_), .B(men_men_n812_), .C(men_men_n898_), .Y(men_men_n1354_));
  NAi31      u1326(.An(men_men_n765_), .B(men_men_n1354_), .C(men_men_n205_), .Y(men_men_n1355_));
  NA4        u1327(.A(men_men_n1355_), .B(men_men_n1353_), .C(men_men_n1347_), .D(men_men_n1235_), .Y(men_men_n1356_));
  NOi31      u1328(.An(men_men_n1320_), .B(men_men_n470_), .C(men_men_n403_), .Y(men_men_n1357_));
  OR3        u1329(.A(men_men_n1357_), .B(men_men_n801_), .C(men_men_n549_), .Y(men_men_n1358_));
  OR3        u1330(.A(men_men_n378_), .B(men_men_n228_), .C(men_men_n625_), .Y(men_men_n1359_));
  AOI210     u1331(.A0(men_men_n578_), .A1(men_men_n455_), .B0(men_men_n380_), .Y(men_men_n1360_));
  NA2        u1332(.A(men_men_n1351_), .B(men_men_n809_), .Y(men_men_n1361_));
  NA4        u1333(.A(men_men_n1361_), .B(men_men_n1360_), .C(men_men_n1359_), .D(men_men_n1358_), .Y(men_men_n1362_));
  AOI220     u1334(.A0(men_men_n1339_), .A1(men_men_n775_), .B0(men_men_n1336_), .B1(men_men_n242_), .Y(men_men_n1363_));
  AN2        u1335(.A(men_men_n951_), .B(men_men_n950_), .Y(men_men_n1364_));
  NO4        u1336(.A(men_men_n1364_), .B(men_men_n896_), .C(men_men_n510_), .D(men_men_n490_), .Y(men_men_n1365_));
  NA3        u1337(.A(men_men_n1365_), .B(men_men_n1363_), .C(men_men_n1301_), .Y(men_men_n1366_));
  NAi21      u1338(.An(j), .B(i), .Y(men_men_n1367_));
  NO4        u1339(.A(men_men_n1311_), .B(men_men_n1367_), .C(men_men_n449_), .D(men_men_n239_), .Y(men_men_n1368_));
  NO4        u1340(.A(men_men_n1368_), .B(men_men_n1366_), .C(men_men_n1362_), .D(men_men_n1356_), .Y(men_men_n1369_));
  NA4        u1341(.A(men_men_n1369_), .B(men_men_n1343_), .C(men_men_n1323_), .D(men_men_n1313_), .Y(men07));
  NOi21      u1342(.An(j), .B(k), .Y(men_men_n1371_));
  NA4        u1343(.A(men_men_n180_), .B(men_men_n111_), .C(men_men_n1371_), .D(f), .Y(men_men_n1372_));
  NAi32      u1344(.An(m), .Bn(b), .C(n), .Y(men_men_n1373_));
  NO3        u1345(.A(men_men_n1373_), .B(g), .C(f), .Y(men_men_n1374_));
  OAI210     u1346(.A0(men_men_n323_), .A1(men_men_n492_), .B0(men_men_n1374_), .Y(men_men_n1375_));
  NAi21      u1347(.An(f), .B(c), .Y(men_men_n1376_));
  OR2        u1348(.A(e), .B(d), .Y(men_men_n1377_));
  OAI220     u1349(.A0(men_men_n1377_), .A1(men_men_n1376_), .B0(men_men_n638_), .B1(men_men_n325_), .Y(men_men_n1378_));
  NA3        u1350(.A(men_men_n1378_), .B(men_men_n1084_), .C(men_men_n180_), .Y(men_men_n1379_));
  NOi31      u1351(.An(n), .B(m), .C(b), .Y(men_men_n1380_));
  NO3        u1352(.A(men_men_n131_), .B(men_men_n456_), .C(h), .Y(men_men_n1381_));
  NA3        u1353(.A(men_men_n1379_), .B(men_men_n1375_), .C(men_men_n1372_), .Y(men_men_n1382_));
  NOi41      u1354(.An(i), .B(n), .C(m), .D(h), .Y(men_men_n1383_));
  NA3        u1355(.A(men_men_n1383_), .B(men_men_n888_), .C(men_men_n417_), .Y(men_men_n1384_));
  NO2        u1356(.A(men_men_n1384_), .B(men_men_n56_), .Y(men_men_n1385_));
  NA2        u1357(.A(men_men_n1114_), .B(men_men_n224_), .Y(men_men_n1386_));
  NO2        u1358(.A(men_men_n1386_), .B(men_men_n61_), .Y(men_men_n1387_));
  NO2        u1359(.A(k), .B(i), .Y(men_men_n1388_));
  NA3        u1360(.A(men_men_n1388_), .B(men_men_n917_), .C(men_men_n180_), .Y(men_men_n1389_));
  NA2        u1361(.A(men_men_n89_), .B(men_men_n45_), .Y(men_men_n1390_));
  NO2        u1362(.A(men_men_n1078_), .B(men_men_n449_), .Y(men_men_n1391_));
  NA3        u1363(.A(men_men_n1391_), .B(men_men_n1390_), .C(men_men_n217_), .Y(men_men_n1392_));
  NO2        u1364(.A(men_men_n1091_), .B(men_men_n307_), .Y(men_men_n1393_));
  NA2        u1365(.A(men_men_n550_), .B(men_men_n82_), .Y(men_men_n1394_));
  NA2        u1366(.A(men_men_n1236_), .B(men_men_n291_), .Y(men_men_n1395_));
  NA4        u1367(.A(men_men_n1395_), .B(men_men_n1394_), .C(men_men_n1392_), .D(men_men_n1389_), .Y(men_men_n1396_));
  NO4        u1368(.A(men_men_n1396_), .B(men_men_n1387_), .C(men_men_n1385_), .D(men_men_n1382_), .Y(men_men_n1397_));
  NO3        u1369(.A(e), .B(d), .C(c), .Y(men_men_n1398_));
  NO2        u1370(.A(men_men_n131_), .B(men_men_n217_), .Y(men_men_n1399_));
  NA2        u1371(.A(men_men_n1399_), .B(men_men_n1398_), .Y(men_men_n1400_));
  NO2        u1372(.A(men_men_n1400_), .B(c), .Y(men_men_n1401_));
  OR2        u1373(.A(h), .B(f), .Y(men_men_n1402_));
  NO3        u1374(.A(n), .B(m), .C(i), .Y(men_men_n1403_));
  OAI210     u1375(.A0(men_men_n1136_), .A1(men_men_n155_), .B0(men_men_n1403_), .Y(men_men_n1404_));
  NO2        u1376(.A(i), .B(g), .Y(men_men_n1405_));
  OR3        u1377(.A(men_men_n1405_), .B(men_men_n1373_), .C(men_men_n72_), .Y(men_men_n1406_));
  OAI220     u1378(.A0(men_men_n1406_), .A1(men_men_n492_), .B0(men_men_n1404_), .B1(men_men_n1402_), .Y(men_men_n1407_));
  NA3        u1379(.A(men_men_n712_), .B(men_men_n699_), .C(men_men_n114_), .Y(men_men_n1408_));
  NA3        u1380(.A(men_men_n1380_), .B(men_men_n1087_), .C(men_men_n687_), .Y(men_men_n1409_));
  AOI210     u1381(.A0(men_men_n1409_), .A1(men_men_n1408_), .B0(men_men_n45_), .Y(men_men_n1410_));
  NO2        u1382(.A(l), .B(k), .Y(men_men_n1411_));
  NOi41      u1383(.An(men_men_n555_), .B(men_men_n1411_), .C(men_men_n485_), .D(men_men_n449_), .Y(men_men_n1412_));
  NO3        u1384(.A(men_men_n449_), .B(d), .C(c), .Y(men_men_n1413_));
  NO4        u1385(.A(men_men_n1412_), .B(men_men_n1410_), .C(men_men_n1407_), .D(men_men_n1401_), .Y(men_men_n1414_));
  NO2        u1386(.A(men_men_n145_), .B(h), .Y(men_men_n1415_));
  NO2        u1387(.A(g), .B(c), .Y(men_men_n1416_));
  NA3        u1388(.A(men_men_n1416_), .B(men_men_n141_), .C(men_men_n188_), .Y(men_men_n1417_));
  INV        u1389(.A(men_men_n1417_), .Y(men_men_n1418_));
  NA2        u1390(.A(men_men_n1418_), .B(men_men_n180_), .Y(men_men_n1419_));
  NO2        u1391(.A(men_men_n457_), .B(a), .Y(men_men_n1420_));
  NA3        u1392(.A(men_men_n1420_), .B(k), .C(men_men_n115_), .Y(men_men_n1421_));
  NO2        u1393(.A(i), .B(h), .Y(men_men_n1422_));
  AOI210     u1394(.A0(men_men_n1159_), .A1(h), .B0(men_men_n422_), .Y(men_men_n1423_));
  NA2        u1395(.A(men_men_n138_), .B(men_men_n224_), .Y(men_men_n1424_));
  NO2        u1396(.A(men_men_n1424_), .B(men_men_n1423_), .Y(men_men_n1425_));
  NO2        u1397(.A(men_men_n772_), .B(men_men_n189_), .Y(men_men_n1426_));
  NOi31      u1398(.An(m), .B(n), .C(b), .Y(men_men_n1427_));
  NOi31      u1399(.An(f), .B(d), .C(c), .Y(men_men_n1428_));
  NA2        u1400(.A(men_men_n1428_), .B(men_men_n1427_), .Y(men_men_n1429_));
  INV        u1401(.A(men_men_n1429_), .Y(men_men_n1430_));
  NO3        u1402(.A(men_men_n1430_), .B(men_men_n1426_), .C(men_men_n1425_), .Y(men_men_n1431_));
  NA2        u1403(.A(men_men_n1105_), .B(men_men_n473_), .Y(men_men_n1432_));
  NO4        u1404(.A(men_men_n1432_), .B(men_men_n1087_), .C(men_men_n449_), .D(men_men_n45_), .Y(men_men_n1433_));
  OAI210     u1405(.A0(men_men_n183_), .A1(men_men_n535_), .B0(men_men_n1088_), .Y(men_men_n1434_));
  NO3        u1406(.A(men_men_n41_), .B(i), .C(h), .Y(men_men_n1435_));
  INV        u1407(.A(men_men_n1434_), .Y(men_men_n1436_));
  NO2        u1408(.A(men_men_n1436_), .B(men_men_n1433_), .Y(men_men_n1437_));
  AN4        u1409(.A(men_men_n1437_), .B(men_men_n1431_), .C(men_men_n1421_), .D(men_men_n1419_), .Y(men_men_n1438_));
  NA2        u1410(.A(men_men_n1380_), .B(men_men_n387_), .Y(men_men_n1439_));
  NO2        u1411(.A(men_men_n1439_), .B(men_men_n1069_), .Y(men_men_n1440_));
  NA2        u1412(.A(men_men_n1413_), .B(men_men_n218_), .Y(men_men_n1441_));
  NO2        u1413(.A(men_men_n189_), .B(b), .Y(men_men_n1442_));
  AOI220     u1414(.A0(men_men_n1191_), .A1(men_men_n1442_), .B0(men_men_n1113_), .B1(men_men_n1432_), .Y(men_men_n1443_));
  NO2        u1415(.A(i), .B(men_men_n216_), .Y(men_men_n1444_));
  NA4        u1416(.A(men_men_n1165_), .B(men_men_n1444_), .C(men_men_n106_), .D(m), .Y(men_men_n1445_));
  NAi41      u1417(.An(men_men_n1440_), .B(men_men_n1445_), .C(men_men_n1443_), .D(men_men_n1441_), .Y(men_men_n1446_));
  NO4        u1418(.A(men_men_n131_), .B(g), .C(f), .D(e), .Y(men_men_n1447_));
  NA3        u1419(.A(men_men_n1388_), .B(men_men_n292_), .C(h), .Y(men_men_n1448_));
  NA2        u1420(.A(men_men_n196_), .B(men_men_n101_), .Y(men_men_n1449_));
  OR2        u1421(.A(e), .B(a), .Y(men_men_n1450_));
  NO2        u1422(.A(men_men_n1377_), .B(men_men_n1376_), .Y(men_men_n1451_));
  AOI210     u1423(.A0(men_men_n30_), .A1(h), .B0(men_men_n1451_), .Y(men_men_n1452_));
  NO2        u1424(.A(men_men_n1452_), .B(men_men_n1102_), .Y(men_men_n1453_));
  NOi41      u1425(.An(h), .B(f), .C(e), .D(a), .Y(men_men_n1454_));
  NA2        u1426(.A(men_men_n1454_), .B(men_men_n115_), .Y(men_men_n1455_));
  NA2        u1427(.A(men_men_n1383_), .B(men_men_n1411_), .Y(men_men_n1456_));
  NA2        u1428(.A(men_men_n1456_), .B(men_men_n1455_), .Y(men_men_n1457_));
  OR3        u1429(.A(men_men_n549_), .B(men_men_n548_), .C(men_men_n114_), .Y(men_men_n1458_));
  NA2        u1430(.A(men_men_n1134_), .B(men_men_n414_), .Y(men_men_n1459_));
  OAI220     u1431(.A0(men_men_n1459_), .A1(men_men_n444_), .B0(men_men_n1458_), .B1(men_men_n301_), .Y(men_men_n1460_));
  AO210      u1432(.A0(men_men_n1460_), .A1(men_men_n117_), .B0(men_men_n1457_), .Y(men_men_n1461_));
  NO3        u1433(.A(men_men_n1461_), .B(men_men_n1453_), .C(men_men_n1446_), .Y(men_men_n1462_));
  NA4        u1434(.A(men_men_n1462_), .B(men_men_n1438_), .C(men_men_n1414_), .D(men_men_n1397_), .Y(men_men_n1463_));
  NA2        u1435(.A(men_men_n387_), .B(men_men_n56_), .Y(men_men_n1464_));
  NA2        u1436(.A(men_men_n218_), .B(men_men_n180_), .Y(men_men_n1465_));
  AOI210     u1437(.A0(men_men_n1465_), .A1(men_men_n1210_), .B0(men_men_n1464_), .Y(men_men_n1466_));
  NO2        u1438(.A(men_men_n399_), .B(j), .Y(men_men_n1467_));
  NA3        u1439(.A(men_men_n1435_), .B(men_men_n1377_), .C(men_men_n1134_), .Y(men_men_n1468_));
  NAi41      u1440(.An(men_men_n1422_), .B(men_men_n1098_), .C(men_men_n168_), .D(men_men_n148_), .Y(men_men_n1469_));
  NA2        u1441(.A(men_men_n1469_), .B(men_men_n1468_), .Y(men_men_n1470_));
  NA3        u1442(.A(g), .B(men_men_n1467_), .C(men_men_n157_), .Y(men_men_n1471_));
  INV        u1443(.A(men_men_n1471_), .Y(men_men_n1472_));
  NO3        u1444(.A(men_men_n765_), .B(men_men_n175_), .C(men_men_n417_), .Y(men_men_n1473_));
  NO3        u1445(.A(men_men_n1473_), .B(men_men_n1472_), .C(men_men_n1470_), .Y(men_men_n1474_));
  NO3        u1446(.A(men_men_n1102_), .B(men_men_n590_), .C(g), .Y(men_men_n1475_));
  NOi21      u1447(.An(men_men_n1465_), .B(men_men_n1475_), .Y(men_men_n1476_));
  AOI210     u1448(.A0(men_men_n1476_), .A1(men_men_n1449_), .B0(men_men_n1078_), .Y(men_men_n1477_));
  OR2        u1449(.A(n), .B(i), .Y(men_men_n1478_));
  OAI210     u1450(.A0(men_men_n1478_), .A1(men_men_n1097_), .B0(men_men_n49_), .Y(men_men_n1479_));
  AOI220     u1451(.A0(men_men_n1479_), .A1(men_men_n1199_), .B0(men_men_n842_), .B1(men_men_n196_), .Y(men_men_n1480_));
  INV        u1452(.A(men_men_n1480_), .Y(men_men_n1481_));
  NO2        u1453(.A(men_men_n131_), .B(l), .Y(men_men_n1482_));
  NO2        u1454(.A(men_men_n228_), .B(k), .Y(men_men_n1483_));
  OAI210     u1455(.A0(men_men_n1483_), .A1(men_men_n1422_), .B0(men_men_n1482_), .Y(men_men_n1484_));
  NO2        u1456(.A(men_men_n1484_), .B(men_men_n31_), .Y(men_men_n1485_));
  NO3        u1457(.A(men_men_n1485_), .B(men_men_n1481_), .C(men_men_n1477_), .Y(men_men_n1486_));
  INV        u1458(.A(men_men_n49_), .Y(men_men_n1487_));
  NO3        u1459(.A(men_men_n1116_), .B(men_men_n1377_), .C(men_men_n49_), .Y(men_men_n1488_));
  NA2        u1460(.A(men_men_n1117_), .B(men_men_n1487_), .Y(men_men_n1489_));
  NO2        u1461(.A(men_men_n1102_), .B(h), .Y(men_men_n1490_));
  NA3        u1462(.A(men_men_n1490_), .B(d), .C(men_men_n1070_), .Y(men_men_n1491_));
  OAI220     u1463(.A0(men_men_n1491_), .A1(c), .B0(men_men_n1489_), .B1(j), .Y(men_men_n1492_));
  NA2        u1464(.A(men_men_n180_), .B(men_men_n114_), .Y(men_men_n1493_));
  AOI210     u1465(.A0(men_men_n535_), .A1(h), .B0(men_men_n69_), .Y(men_men_n1494_));
  NA2        u1466(.A(men_men_n1494_), .B(men_men_n1420_), .Y(men_men_n1495_));
  NO2        u1467(.A(men_men_n1367_), .B(men_men_n175_), .Y(men_men_n1496_));
  NOi21      u1468(.An(d), .B(f), .Y(men_men_n1497_));
  NO3        u1469(.A(men_men_n1428_), .B(men_men_n1497_), .C(men_men_n40_), .Y(men_men_n1498_));
  NA2        u1470(.A(men_men_n1498_), .B(men_men_n1496_), .Y(men_men_n1499_));
  NO2        u1471(.A(men_men_n1377_), .B(f), .Y(men_men_n1500_));
  NO2        u1472(.A(men_men_n301_), .B(c), .Y(men_men_n1501_));
  NA2        u1473(.A(men_men_n1501_), .B(men_men_n550_), .Y(men_men_n1502_));
  NA3        u1474(.A(men_men_n1502_), .B(men_men_n1499_), .C(men_men_n1495_), .Y(men_men_n1503_));
  NO2        u1475(.A(men_men_n1503_), .B(men_men_n1492_), .Y(men_men_n1504_));
  NA4        u1476(.A(men_men_n1504_), .B(men_men_n1486_), .C(men_men_n1474_), .D(men_men_n1585_), .Y(men_men_n1505_));
  NO3        u1477(.A(men_men_n1105_), .B(men_men_n1097_), .C(men_men_n40_), .Y(men_men_n1506_));
  NO2        u1478(.A(men_men_n473_), .B(men_men_n301_), .Y(men_men_n1507_));
  OAI210     u1479(.A0(men_men_n1507_), .A1(men_men_n1506_), .B0(men_men_n1393_), .Y(men_men_n1508_));
  OAI210     u1480(.A0(men_men_n1447_), .A1(men_men_n1380_), .B0(men_men_n903_), .Y(men_men_n1509_));
  NO2        u1481(.A(men_men_n1066_), .B(men_men_n131_), .Y(men_men_n1510_));
  NA2        u1482(.A(men_men_n1510_), .B(men_men_n631_), .Y(men_men_n1511_));
  NA3        u1483(.A(men_men_n1511_), .B(men_men_n1509_), .C(men_men_n1508_), .Y(men_men_n1512_));
  NA2        u1484(.A(men_men_n1416_), .B(men_men_n1497_), .Y(men_men_n1513_));
  NO2        u1485(.A(men_men_n1513_), .B(m), .Y(men_men_n1514_));
  NA3        u1486(.A(men_men_n1114_), .B(men_men_n111_), .C(men_men_n224_), .Y(men_men_n1515_));
  NO2        u1487(.A(men_men_n149_), .B(men_men_n182_), .Y(men_men_n1516_));
  OAI210     u1488(.A0(men_men_n1516_), .A1(men_men_n112_), .B0(men_men_n1427_), .Y(men_men_n1517_));
  NA2        u1489(.A(men_men_n1517_), .B(men_men_n1515_), .Y(men_men_n1518_));
  NO3        u1490(.A(men_men_n1518_), .B(men_men_n1514_), .C(men_men_n1512_), .Y(men_men_n1519_));
  NO2        u1491(.A(men_men_n1376_), .B(e), .Y(men_men_n1520_));
  NA2        u1492(.A(men_men_n1520_), .B(men_men_n412_), .Y(men_men_n1521_));
  OAI210     u1493(.A0(men_men_n1500_), .A1(men_men_n1145_), .B0(men_men_n642_), .Y(men_men_n1522_));
  OR3        u1494(.A(men_men_n1483_), .B(men_men_n1236_), .C(men_men_n131_), .Y(men_men_n1523_));
  OAI220     u1495(.A0(men_men_n1523_), .A1(men_men_n1521_), .B0(men_men_n1522_), .B1(men_men_n451_), .Y(men_men_n1524_));
  NO3        u1496(.A(men_men_n1458_), .B(men_men_n358_), .C(a), .Y(men_men_n1525_));
  NO2        u1497(.A(men_men_n1525_), .B(men_men_n1524_), .Y(men_men_n1526_));
  NO2        u1498(.A(men_men_n182_), .B(c), .Y(men_men_n1527_));
  OAI210     u1499(.A0(men_men_n1527_), .A1(men_men_n1520_), .B0(men_men_n180_), .Y(men_men_n1528_));
  AOI220     u1500(.A0(men_men_n1528_), .A1(men_men_n1099_), .B0(men_men_n542_), .B1(men_men_n374_), .Y(men_men_n1529_));
  NA2        u1501(.A(men_men_n548_), .B(g), .Y(men_men_n1530_));
  AOI210     u1502(.A0(men_men_n1530_), .A1(men_men_n1413_), .B0(men_men_n1488_), .Y(men_men_n1531_));
  NA2        u1503(.A(men_men_n1145_), .B(a), .Y(men_men_n1532_));
  OAI220     u1504(.A0(men_men_n1532_), .A1(men_men_n69_), .B0(men_men_n1531_), .B1(men_men_n216_), .Y(men_men_n1533_));
  AOI210     u1505(.A0(men_men_n922_), .A1(men_men_n424_), .B0(men_men_n107_), .Y(men_men_n1534_));
  OR2        u1506(.A(men_men_n1534_), .B(men_men_n548_), .Y(men_men_n1535_));
  NO2        u1507(.A(men_men_n1535_), .B(men_men_n175_), .Y(men_men_n1536_));
  NA4        u1508(.A(men_men_n1114_), .B(men_men_n1111_), .C(men_men_n224_), .D(men_men_n68_), .Y(men_men_n1537_));
  NA2        u1509(.A(men_men_n1381_), .B(men_men_n183_), .Y(men_men_n1538_));
  NO2        u1510(.A(men_men_n49_), .B(l), .Y(men_men_n1539_));
  OAI210     u1511(.A0(men_men_n1450_), .A1(men_men_n880_), .B0(men_men_n492_), .Y(men_men_n1540_));
  OAI210     u1512(.A0(men_men_n1540_), .A1(men_men_n1117_), .B0(men_men_n1539_), .Y(men_men_n1541_));
  NO2        u1513(.A(men_men_n255_), .B(g), .Y(men_men_n1542_));
  NO2        u1514(.A(m), .B(i), .Y(men_men_n1543_));
  BUFFER     u1515(.A(men_men_n1543_), .Y(men_men_n1544_));
  AOI220     u1516(.A0(men_men_n1544_), .A1(men_men_n1415_), .B0(men_men_n1098_), .B1(men_men_n1542_), .Y(men_men_n1545_));
  NA4        u1517(.A(men_men_n1545_), .B(men_men_n1541_), .C(men_men_n1538_), .D(men_men_n1537_), .Y(men_men_n1546_));
  NO4        u1518(.A(men_men_n1546_), .B(men_men_n1536_), .C(men_men_n1533_), .D(men_men_n1529_), .Y(men_men_n1547_));
  NA3        u1519(.A(men_men_n1547_), .B(men_men_n1526_), .C(men_men_n1519_), .Y(men_men_n1548_));
  NA3        u1520(.A(men_men_n982_), .B(men_men_n138_), .C(men_men_n46_), .Y(men_men_n1549_));
  AOI210     u1521(.A0(men_men_n146_), .A1(c), .B0(men_men_n1549_), .Y(men_men_n1550_));
  INV        u1522(.A(men_men_n186_), .Y(men_men_n1551_));
  NA2        u1523(.A(men_men_n1551_), .B(men_men_n1490_), .Y(men_men_n1552_));
  OR2        u1524(.A(men_men_n132_), .B(men_men_n1439_), .Y(men_men_n1553_));
  NO2        u1525(.A(men_men_n72_), .B(c), .Y(men_men_n1554_));
  NO4        u1526(.A(men_men_n1402_), .B(men_men_n187_), .C(men_men_n456_), .D(men_men_n45_), .Y(men_men_n1555_));
  AOI210     u1527(.A0(men_men_n1496_), .A1(men_men_n1554_), .B0(men_men_n1555_), .Y(men_men_n1556_));
  NA3        u1528(.A(men_men_n1556_), .B(men_men_n1553_), .C(men_men_n1552_), .Y(men_men_n1557_));
  NO2        u1529(.A(men_men_n1557_), .B(men_men_n1550_), .Y(men_men_n1558_));
  NO4        u1530(.A(men_men_n228_), .B(men_men_n187_), .C(men_men_n260_), .D(k), .Y(men_men_n1559_));
  AOI210     u1531(.A0(men_men_n155_), .A1(men_men_n56_), .B0(men_men_n1520_), .Y(men_men_n1560_));
  NO2        u1532(.A(men_men_n1560_), .B(men_men_n1493_), .Y(men_men_n1561_));
  NO2        u1533(.A(men_men_n1549_), .B(men_men_n112_), .Y(men_men_n1562_));
  NOi21      u1534(.An(men_men_n1381_), .B(e), .Y(men_men_n1563_));
  NO4        u1535(.A(men_men_n1563_), .B(men_men_n1562_), .C(men_men_n1561_), .D(men_men_n1559_), .Y(men_men_n1564_));
  AOI220     u1536(.A0(men_men_n1543_), .A1(men_men_n652_), .B0(men_men_n1084_), .B1(men_men_n158_), .Y(men_men_n1565_));
  NOi31      u1537(.An(men_men_n30_), .B(men_men_n1565_), .C(n), .Y(men_men_n1566_));
  INV        u1538(.A(men_men_n1566_), .Y(men_men_n1567_));
  NA2        u1539(.A(men_men_n59_), .B(a), .Y(men_men_n1568_));
  NO2        u1540(.A(men_men_n1388_), .B(men_men_n119_), .Y(men_men_n1569_));
  OAI220     u1541(.A0(men_men_n1569_), .A1(men_men_n1439_), .B0(men_men_n1459_), .B1(men_men_n1568_), .Y(men_men_n1570_));
  INV        u1542(.A(men_men_n1570_), .Y(men_men_n1571_));
  NA4        u1543(.A(men_men_n1571_), .B(men_men_n1567_), .C(men_men_n1564_), .D(men_men_n1558_), .Y(men_men_n1572_));
  OR4        u1544(.A(men_men_n1572_), .B(men_men_n1548_), .C(men_men_n1505_), .D(men_men_n1463_), .Y(men04));
  NOi31      u1545(.An(men_men_n1447_), .B(men_men_n1448_), .C(men_men_n1072_), .Y(men_men_n1574_));
  NA2        u1546(.A(men_men_n1500_), .B(men_men_n842_), .Y(men_men_n1575_));
  NO4        u1547(.A(men_men_n1575_), .B(men_men_n1061_), .C(men_men_n493_), .D(j), .Y(men_men_n1576_));
  OR3        u1548(.A(men_men_n1576_), .B(men_men_n1574_), .C(men_men_n1090_), .Y(men_men_n1577_));
  NO3        u1549(.A(men_men_n1390_), .B(men_men_n93_), .C(k), .Y(men_men_n1578_));
  AOI210     u1550(.A0(men_men_n1578_), .A1(men_men_n1083_), .B0(men_men_n1212_), .Y(men_men_n1579_));
  NA2        u1551(.A(men_men_n1579_), .B(men_men_n1240_), .Y(men_men_n1580_));
  NO4        u1552(.A(men_men_n1580_), .B(men_men_n1577_), .C(men_men_n1096_), .D(men_men_n1077_), .Y(men_men_n1581_));
  NA4        u1553(.A(men_men_n1581_), .B(men_men_n1147_), .C(men_men_n1132_), .D(men_men_n1120_), .Y(men05));
  INV        u1554(.A(men_men_n1466_), .Y(men_men_n1585_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
  VOTADOR g7(.A(ori07), .B(mai07), .C(men07), .Y(z7));
  VOTADOR g8(.A(ori08), .B(mai08), .C(men08), .Y(z8));
  VOTADOR g9(.A(ori09), .B(mai09), .C(men09), .Y(z9));
  VOTADOR g10(.A(ori10), .B(mai10), .C(men10), .Y(z10));
  VOTADOR g11(.A(ori11), .B(mai11), .C(men11), .Y(z11));
  VOTADOR g12(.A(ori12), .B(mai12), .C(men12), .Y(z12));
  VOTADOR g13(.A(ori13), .B(mai13), .C(men13), .Y(z13));
endmodule