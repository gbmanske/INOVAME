// Benchmark "top" written by ABC on Fri Jun 21 17:49:28 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n129_, new_new_n130_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n409_,
    new_new_n410_, new_new_n411_, new_new_n412_, new_new_n413_,
    new_new_n414_, new_new_n415_, new_new_n416_, new_new_n417_,
    new_new_n418_, new_new_n419_, new_new_n420_, new_new_n421_,
    new_new_n422_, new_new_n423_, new_new_n424_, new_new_n425_,
    new_new_n426_, new_new_n427_, new_new_n428_, new_new_n429_,
    new_new_n430_, new_new_n431_, new_new_n432_, new_new_n433_,
    new_new_n434_, new_new_n435_, new_new_n436_, new_new_n437_,
    new_new_n438_, new_new_n439_, new_new_n440_, new_new_n441_,
    new_new_n442_, new_new_n443_, new_new_n444_, new_new_n445_,
    new_new_n446_, new_new_n447_, new_new_n448_, new_new_n449_,
    new_new_n450_, new_new_n451_, new_new_n452_, new_new_n453_,
    new_new_n454_, new_new_n455_, new_new_n456_, new_new_n457_,
    new_new_n458_, new_new_n459_, new_new_n460_, new_new_n461_,
    new_new_n462_, new_new_n463_, new_new_n464_, new_new_n465_,
    new_new_n466_, new_new_n467_, new_new_n468_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n532_, new_new_n533_, new_new_n534_,
    new_new_n535_, new_new_n536_, new_new_n537_, new_new_n538_,
    new_new_n539_, new_new_n540_, new_new_n541_, new_new_n542_,
    new_new_n543_, new_new_n544_, new_new_n545_, new_new_n546_,
    new_new_n547_, new_new_n548_, new_new_n549_, new_new_n550_,
    new_new_n551_, new_new_n552_, new_new_n553_, new_new_n554_,
    new_new_n555_, new_new_n556_, new_new_n557_, new_new_n558_,
    new_new_n559_, new_new_n560_, new_new_n561_, new_new_n562_,
    new_new_n563_, new_new_n564_, new_new_n565_, new_new_n566_,
    new_new_n567_, new_new_n568_, new_new_n569_, new_new_n570_,
    new_new_n571_, new_new_n572_, new_new_n573_, new_new_n575_,
    new_new_n576_, new_new_n577_, new_new_n578_, new_new_n579_,
    new_new_n580_, new_new_n581_, new_new_n582_, new_new_n583_,
    new_new_n584_, new_new_n585_, new_new_n586_, new_new_n587_,
    new_new_n588_, new_new_n589_, new_new_n590_, new_new_n591_,
    new_new_n592_, new_new_n593_, new_new_n594_, new_new_n595_,
    new_new_n596_, new_new_n597_, new_new_n598_, new_new_n599_,
    new_new_n600_, new_new_n601_, new_new_n602_, new_new_n603_,
    new_new_n604_, new_new_n605_, new_new_n606_, new_new_n607_,
    new_new_n608_, new_new_n609_, new_new_n610_, new_new_n611_,
    new_new_n612_, new_new_n614_, new_new_n615_, new_new_n616_,
    new_new_n617_, new_new_n618_, new_new_n619_, new_new_n620_,
    new_new_n621_, new_new_n622_, new_new_n623_, new_new_n624_,
    new_new_n625_, new_new_n626_, new_new_n627_, new_new_n628_,
    new_new_n629_, new_new_n630_, new_new_n631_, new_new_n632_,
    new_new_n633_, new_new_n634_, new_new_n635_, new_new_n636_,
    new_new_n637_, new_new_n638_, new_new_n639_, new_new_n640_,
    new_new_n641_, new_new_n642_, new_new_n643_, new_new_n644_,
    new_new_n645_, new_new_n646_, new_new_n647_, new_new_n648_,
    new_new_n649_, new_new_n650_, new_new_n651_, new_new_n652_,
    new_new_n653_, new_new_n654_, new_new_n655_, new_new_n656_,
    new_new_n657_, new_new_n658_, new_new_n659_, new_new_n660_,
    new_new_n661_, new_new_n662_, new_new_n663_, new_new_n664_,
    new_new_n665_, new_new_n666_, new_new_n667_, new_new_n668_,
    new_new_n669_, new_new_n670_, new_new_n671_, new_new_n672_,
    new_new_n673_, new_new_n674_, new_new_n675_, new_new_n676_,
    new_new_n677_, new_new_n678_, new_new_n679_, new_new_n680_,
    new_new_n681_, new_new_n682_, new_new_n683_, new_new_n684_,
    new_new_n685_, new_new_n686_, new_new_n687_, new_new_n688_,
    new_new_n689_, new_new_n690_, new_new_n691_, new_new_n692_,
    new_new_n693_, new_new_n694_, new_new_n695_, new_new_n696_,
    new_new_n697_, new_new_n698_, new_new_n699_, new_new_n700_,
    new_new_n701_, new_new_n702_, new_new_n703_, new_new_n704_,
    new_new_n705_, new_new_n706_, new_new_n707_, new_new_n708_,
    new_new_n709_, new_new_n710_, new_new_n711_, new_new_n712_,
    new_new_n713_, new_new_n714_, new_new_n715_, new_new_n716_,
    new_new_n717_, new_new_n718_, new_new_n719_, new_new_n720_,
    new_new_n721_, new_new_n722_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n764_, new_new_n765_, new_new_n766_, new_new_n767_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(ori1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  NA2        g023(.A(i_0_), .B(i_3_), .Y(new_new_n46_));
  INV        g024(.A(i_5_), .Y(new_new_n47_));
  NO2        g025(.A(i_7_), .B(i_10_), .Y(new_new_n48_));
  AOI210     g026(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n48_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_5_), .A1(new_new_n46_), .B0(new_new_n45_), .Y(new_new_n50_));
  NA2        g028(.A(i_0_), .B(i_2_), .Y(new_new_n51_));
  NA2        g029(.A(i_7_), .B(i_9_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n51_), .Y(new_new_n53_));
  NA2        g031(.A(new_new_n50_), .B(new_new_n44_), .Y(new_new_n54_));
  NO2        g032(.A(i_1_), .B(i_6_), .Y(new_new_n55_));
  NA2        g033(.A(i_8_), .B(i_7_), .Y(new_new_n56_));
  NAi21      g034(.An(i_2_), .B(i_7_), .Y(new_new_n57_));
  INV        g035(.A(i_1_), .Y(new_new_n58_));
  NA2        g036(.A(new_new_n58_), .B(i_6_), .Y(new_new_n59_));
  NA3        g037(.A(new_new_n59_), .B(new_new_n57_), .C(new_new_n31_), .Y(new_new_n60_));
  NA2        g038(.A(i_1_), .B(i_10_), .Y(new_new_n61_));
  NO2        g039(.A(new_new_n61_), .B(i_6_), .Y(new_new_n62_));
  NAi21      g040(.An(new_new_n62_), .B(new_new_n60_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n49_), .B(i_2_), .Y(new_new_n64_));
  AOI210     g042(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_6_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(new_new_n25_), .Y(new_new_n67_));
  INV        g045(.A(i_0_), .Y(new_new_n68_));
  NAi21      g046(.An(i_5_), .B(i_10_), .Y(new_new_n69_));
  NA2        g047(.A(i_5_), .B(i_9_), .Y(new_new_n70_));
  AOI210     g048(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n68_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n67_), .Y(new_new_n72_));
  INV        g050(.A(new_new_n72_), .Y(new_new_n73_));
  OAI210     g051(.A0(new_new_n73_), .A1(new_new_n63_), .B0(i_0_), .Y(new_new_n74_));
  NA2        g052(.A(i_12_), .B(i_5_), .Y(new_new_n75_));
  INV        g053(.A(i_8_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n55_), .Y(new_new_n77_));
  INV        g055(.A(i_3_), .Y(new_new_n78_));
  NO2        g056(.A(i_3_), .B(i_7_), .Y(new_new_n79_));
  NO2        g057(.A(new_new_n78_), .B(new_new_n58_), .Y(new_new_n80_));
  INV        g058(.A(i_6_), .Y(new_new_n81_));
  OR4        g059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n82_));
  INV        g060(.A(new_new_n82_), .Y(new_new_n83_));
  NO2        g061(.A(i_2_), .B(i_7_), .Y(new_new_n84_));
  INV        g062(.A(new_new_n84_), .Y(new_new_n85_));
  OAI210     g063(.A0(new_new_n80_), .A1(new_new_n77_), .B0(new_new_n85_), .Y(new_new_n86_));
  NAi21      g064(.An(i_6_), .B(i_10_), .Y(new_new_n87_));
  NA2        g065(.A(i_6_), .B(i_9_), .Y(new_new_n88_));
  AOI210     g066(.A0(new_new_n88_), .A1(new_new_n87_), .B0(new_new_n58_), .Y(new_new_n89_));
  NA2        g067(.A(i_2_), .B(i_6_), .Y(new_new_n90_));
  NO3        g068(.A(new_new_n90_), .B(new_new_n48_), .C(new_new_n25_), .Y(new_new_n91_));
  NO2        g069(.A(new_new_n91_), .B(new_new_n89_), .Y(new_new_n92_));
  AOI210     g070(.A0(new_new_n92_), .A1(new_new_n86_), .B0(new_new_n75_), .Y(new_new_n93_));
  AN3        g071(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n94_));
  NAi21      g072(.An(i_6_), .B(i_11_), .Y(new_new_n95_));
  NA2        g073(.A(new_new_n94_), .B(new_new_n32_), .Y(new_new_n96_));
  INV        g074(.A(i_7_), .Y(new_new_n97_));
  NA2        g075(.A(new_new_n45_), .B(new_new_n97_), .Y(new_new_n98_));
  NO2        g076(.A(i_0_), .B(i_5_), .Y(new_new_n99_));
  NO2        g077(.A(new_new_n99_), .B(new_new_n81_), .Y(new_new_n100_));
  NA2        g078(.A(i_12_), .B(i_3_), .Y(new_new_n101_));
  INV        g079(.A(new_new_n101_), .Y(new_new_n102_));
  NA3        g080(.A(new_new_n102_), .B(new_new_n100_), .C(new_new_n98_), .Y(new_new_n103_));
  NAi21      g081(.An(i_7_), .B(i_11_), .Y(new_new_n104_));
  NO3        g082(.A(new_new_n104_), .B(new_new_n87_), .C(new_new_n51_), .Y(new_new_n105_));
  AN2        g083(.A(i_2_), .B(i_10_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(i_7_), .Y(new_new_n107_));
  OR2        g085(.A(new_new_n75_), .B(new_new_n55_), .Y(new_new_n108_));
  NA2        g086(.A(i_12_), .B(i_7_), .Y(new_new_n109_));
  NA2        g087(.A(i_11_), .B(i_12_), .Y(new_new_n110_));
  NAi41      g088(.An(new_new_n105_), .B(new_new_n110_), .C(new_new_n103_), .D(new_new_n96_), .Y(new_new_n111_));
  NOi21      g089(.An(i_1_), .B(i_5_), .Y(new_new_n112_));
  NA2        g090(.A(new_new_n112_), .B(i_11_), .Y(new_new_n113_));
  NA2        g091(.A(new_new_n97_), .B(new_new_n37_), .Y(new_new_n114_));
  NA2        g092(.A(i_7_), .B(new_new_n25_), .Y(new_new_n115_));
  NA2        g093(.A(new_new_n115_), .B(new_new_n114_), .Y(new_new_n116_));
  NO2        g094(.A(new_new_n116_), .B(new_new_n45_), .Y(new_new_n117_));
  NA2        g095(.A(new_new_n88_), .B(new_new_n87_), .Y(new_new_n118_));
  NAi21      g096(.An(i_3_), .B(i_8_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(new_new_n57_), .Y(new_new_n120_));
  NOi31      g098(.An(new_new_n120_), .B(new_new_n118_), .C(new_new_n117_), .Y(new_new_n121_));
  NO2        g099(.A(i_1_), .B(new_new_n81_), .Y(new_new_n122_));
  NO2        g100(.A(i_6_), .B(i_5_), .Y(new_new_n123_));
  NA2        g101(.A(new_new_n123_), .B(i_3_), .Y(new_new_n124_));
  AO210      g102(.A0(new_new_n124_), .A1(new_new_n46_), .B0(new_new_n122_), .Y(new_new_n125_));
  OAI220     g103(.A0(new_new_n125_), .A1(new_new_n104_), .B0(new_new_n121_), .B1(new_new_n113_), .Y(new_new_n126_));
  NO3        g104(.A(new_new_n126_), .B(new_new_n111_), .C(new_new_n93_), .Y(new_new_n127_));
  NA3        g105(.A(new_new_n127_), .B(new_new_n74_), .C(new_new_n54_), .Y(ori2));
  NO2        g106(.A(new_new_n58_), .B(new_new_n37_), .Y(new_new_n129_));
  NA2        g107(.A(new_new_n764_), .B(new_new_n129_), .Y(new_new_n130_));
  NA4        g108(.A(new_new_n130_), .B(new_new_n72_), .C(new_new_n64_), .D(new_new_n30_), .Y(ori0));
  NO2        g109(.A(i_12_), .B(i_13_), .Y(new_new_n132_));
  NAi21      g110(.An(i_5_), .B(i_11_), .Y(new_new_n133_));
  NOi21      g111(.An(new_new_n132_), .B(new_new_n133_), .Y(new_new_n134_));
  NO2        g112(.A(i_0_), .B(i_1_), .Y(new_new_n135_));
  NA2        g113(.A(i_2_), .B(i_3_), .Y(new_new_n136_));
  NO2        g114(.A(new_new_n136_), .B(i_4_), .Y(new_new_n137_));
  NA3        g115(.A(new_new_n137_), .B(new_new_n135_), .C(new_new_n134_), .Y(new_new_n138_));
  NA2        g116(.A(i_1_), .B(i_5_), .Y(new_new_n139_));
  OR2        g117(.A(i_0_), .B(i_1_), .Y(new_new_n140_));
  NAi32      g118(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n141_));
  NOi21      g119(.An(i_4_), .B(i_10_), .Y(new_new_n142_));
  NA2        g120(.A(new_new_n142_), .B(new_new_n39_), .Y(new_new_n143_));
  NOi21      g121(.An(i_4_), .B(i_9_), .Y(new_new_n144_));
  NOi21      g122(.An(i_11_), .B(i_13_), .Y(new_new_n145_));
  NA2        g123(.A(new_new_n145_), .B(new_new_n144_), .Y(new_new_n146_));
  NO2        g124(.A(i_4_), .B(i_5_), .Y(new_new_n147_));
  NAi21      g125(.An(i_12_), .B(i_11_), .Y(new_new_n148_));
  NO2        g126(.A(new_new_n148_), .B(i_13_), .Y(new_new_n149_));
  NO2        g127(.A(new_new_n68_), .B(new_new_n58_), .Y(new_new_n150_));
  NO2        g128(.A(new_new_n68_), .B(i_5_), .Y(new_new_n151_));
  NO2        g129(.A(i_13_), .B(i_10_), .Y(new_new_n152_));
  NA3        g130(.A(new_new_n152_), .B(new_new_n151_), .C(new_new_n43_), .Y(new_new_n153_));
  NO2        g131(.A(i_2_), .B(i_1_), .Y(new_new_n154_));
  NA2        g132(.A(new_new_n154_), .B(i_3_), .Y(new_new_n155_));
  NAi21      g133(.An(i_4_), .B(i_12_), .Y(new_new_n156_));
  INV        g134(.A(i_8_), .Y(new_new_n157_));
  NO3        g135(.A(i_3_), .B(new_new_n81_), .C(new_new_n47_), .Y(new_new_n158_));
  NA2        g136(.A(new_new_n158_), .B(new_new_n766_), .Y(new_new_n159_));
  NO3        g137(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n160_));
  NO3        g138(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n161_));
  NA2        g139(.A(i_12_), .B(new_new_n161_), .Y(new_new_n162_));
  NO2        g140(.A(new_new_n162_), .B(new_new_n159_), .Y(new_new_n163_));
  NO2        g141(.A(i_3_), .B(i_8_), .Y(new_new_n164_));
  NO3        g142(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n165_));
  NA3        g143(.A(new_new_n165_), .B(new_new_n164_), .C(new_new_n39_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n99_), .B(new_new_n55_), .Y(new_new_n167_));
  NO2        g145(.A(i_13_), .B(i_9_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_3_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n43_), .B(i_5_), .Y(new_new_n170_));
  INV        g148(.A(new_new_n163_), .Y(new_new_n171_));
  NO2        g149(.A(new_new_n171_), .B(i_4_), .Y(new_new_n172_));
  NAi21      g150(.An(i_12_), .B(i_7_), .Y(new_new_n173_));
  NA3        g151(.A(i_13_), .B(new_new_n157_), .C(i_10_), .Y(new_new_n174_));
  NO2        g152(.A(new_new_n174_), .B(new_new_n173_), .Y(new_new_n175_));
  NA2        g153(.A(i_0_), .B(i_5_), .Y(new_new_n176_));
  OAI220     g154(.A0(new_new_n81_), .A1(new_new_n155_), .B0(i_2_), .B1(new_new_n124_), .Y(new_new_n177_));
  NAi31      g155(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n178_));
  NO2        g156(.A(new_new_n36_), .B(i_13_), .Y(new_new_n179_));
  NO2        g157(.A(new_new_n45_), .B(new_new_n58_), .Y(new_new_n180_));
  NA3        g158(.A(new_new_n180_), .B(i_3_), .C(new_new_n179_), .Y(new_new_n181_));
  INV        g159(.A(i_13_), .Y(new_new_n182_));
  NO2        g160(.A(i_12_), .B(new_new_n182_), .Y(new_new_n183_));
  NA3        g161(.A(new_new_n183_), .B(new_new_n160_), .C(new_new_n158_), .Y(new_new_n184_));
  OAI210     g162(.A0(new_new_n181_), .A1(new_new_n178_), .B0(new_new_n184_), .Y(new_new_n185_));
  AOI220     g163(.A0(new_new_n185_), .A1(i_7_), .B0(new_new_n177_), .B1(new_new_n175_), .Y(new_new_n186_));
  NO2        g164(.A(i_12_), .B(new_new_n37_), .Y(new_new_n187_));
  OR2        g165(.A(i_8_), .B(i_7_), .Y(new_new_n188_));
  INV        g166(.A(i_12_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n43_), .B(new_new_n189_), .Y(new_new_n190_));
  NO3        g168(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n191_));
  NA2        g169(.A(i_2_), .B(i_1_), .Y(new_new_n192_));
  NO3        g170(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n193_));
  NAi21      g171(.An(i_4_), .B(i_3_), .Y(new_new_n194_));
  NO2        g172(.A(i_0_), .B(i_6_), .Y(new_new_n195_));
  NOi41      g173(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n196_));
  NO2        g174(.A(i_11_), .B(new_new_n182_), .Y(new_new_n197_));
  NOi21      g175(.An(i_1_), .B(i_6_), .Y(new_new_n198_));
  NAi21      g176(.An(i_3_), .B(i_7_), .Y(new_new_n199_));
  NA2        g177(.A(new_new_n189_), .B(i_9_), .Y(new_new_n200_));
  OR4        g178(.A(new_new_n200_), .B(new_new_n199_), .C(new_new_n198_), .D(new_new_n151_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n68_), .B(i_5_), .Y(new_new_n202_));
  NA2        g180(.A(i_3_), .B(i_9_), .Y(new_new_n203_));
  NAi21      g181(.An(i_7_), .B(i_10_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n204_), .B(new_new_n203_), .Y(new_new_n205_));
  NA3        g183(.A(new_new_n205_), .B(new_new_n202_), .C(new_new_n59_), .Y(new_new_n206_));
  NA2        g184(.A(new_new_n206_), .B(new_new_n201_), .Y(new_new_n207_));
  NA2        g185(.A(new_new_n189_), .B(i_13_), .Y(new_new_n208_));
  NA2        g186(.A(new_new_n207_), .B(new_new_n197_), .Y(new_new_n209_));
  NO2        g187(.A(new_new_n188_), .B(new_new_n37_), .Y(new_new_n210_));
  NA2        g188(.A(i_12_), .B(i_6_), .Y(new_new_n211_));
  OR2        g189(.A(i_13_), .B(i_9_), .Y(new_new_n212_));
  NO3        g190(.A(new_new_n212_), .B(new_new_n211_), .C(new_new_n47_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n194_), .B(i_2_), .Y(new_new_n214_));
  NA3        g192(.A(new_new_n214_), .B(new_new_n213_), .C(new_new_n43_), .Y(new_new_n215_));
  NA2        g193(.A(new_new_n197_), .B(i_9_), .Y(new_new_n216_));
  NA2        g194(.A(new_new_n202_), .B(new_new_n59_), .Y(new_new_n217_));
  OAI210     g195(.A0(new_new_n217_), .A1(new_new_n216_), .B0(new_new_n215_), .Y(new_new_n218_));
  NO3        g196(.A(i_11_), .B(new_new_n182_), .C(new_new_n25_), .Y(new_new_n219_));
  NA2        g197(.A(new_new_n218_), .B(new_new_n210_), .Y(new_new_n220_));
  NA3        g198(.A(new_new_n220_), .B(new_new_n209_), .C(new_new_n186_), .Y(new_new_n221_));
  NO3        g199(.A(i_12_), .B(new_new_n182_), .C(new_new_n37_), .Y(new_new_n222_));
  NO2        g200(.A(new_new_n192_), .B(i_0_), .Y(new_new_n223_));
  NO2        g201(.A(i_3_), .B(i_10_), .Y(new_new_n224_));
  NO2        g202(.A(i_2_), .B(new_new_n97_), .Y(new_new_n225_));
  AN2        g203(.A(i_3_), .B(i_10_), .Y(new_new_n226_));
  NO2        g204(.A(i_5_), .B(new_new_n37_), .Y(new_new_n227_));
  NO2        g205(.A(new_new_n45_), .B(new_new_n26_), .Y(new_new_n228_));
  NO2        g206(.A(new_new_n221_), .B(new_new_n172_), .Y(new_new_n229_));
  NO3        g207(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n230_));
  NO2        g208(.A(i_2_), .B(i_3_), .Y(new_new_n231_));
  OR2        g209(.A(i_0_), .B(i_5_), .Y(new_new_n232_));
  NA2        g210(.A(new_new_n176_), .B(new_new_n232_), .Y(new_new_n233_));
  NO2        g211(.A(new_new_n140_), .B(new_new_n45_), .Y(new_new_n234_));
  NO2        g212(.A(i_12_), .B(i_10_), .Y(new_new_n235_));
  NOi21      g213(.An(i_5_), .B(i_0_), .Y(new_new_n236_));
  NO2        g214(.A(i_2_), .B(new_new_n97_), .Y(new_new_n237_));
  NO4        g215(.A(new_new_n237_), .B(i_4_), .C(new_new_n236_), .D(new_new_n119_), .Y(new_new_n238_));
  NA4        g216(.A(new_new_n79_), .B(new_new_n36_), .C(new_new_n81_), .D(i_8_), .Y(new_new_n239_));
  NA2        g217(.A(new_new_n238_), .B(new_new_n235_), .Y(new_new_n240_));
  NO2        g218(.A(i_6_), .B(i_8_), .Y(new_new_n241_));
  NO2        g219(.A(i_1_), .B(i_7_), .Y(new_new_n242_));
  INV        g220(.A(new_new_n240_), .Y(new_new_n243_));
  NA3        g221(.A(new_new_n198_), .B(new_new_n225_), .C(new_new_n157_), .Y(new_new_n244_));
  NO2        g222(.A(new_new_n157_), .B(i_9_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n245_), .B(new_new_n167_), .Y(new_new_n246_));
  NO2        g224(.A(new_new_n244_), .B(new_new_n143_), .Y(new_new_n247_));
  AOI210     g225(.A0(new_new_n243_), .A1(new_new_n230_), .B0(new_new_n247_), .Y(new_new_n248_));
  NOi32      g226(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n249_));
  INV        g227(.A(new_new_n249_), .Y(new_new_n250_));
  NAi21      g228(.An(i_1_), .B(i_5_), .Y(new_new_n251_));
  NAi41      g229(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n252_));
  OAI220     g230(.A0(new_new_n252_), .A1(new_new_n251_), .B0(new_new_n178_), .B1(new_new_n141_), .Y(new_new_n253_));
  AOI210     g231(.A0(new_new_n252_), .A1(new_new_n141_), .B0(new_new_n140_), .Y(new_new_n254_));
  NOi32      g232(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n255_));
  NAi21      g233(.An(i_6_), .B(i_1_), .Y(new_new_n256_));
  NA3        g234(.A(new_new_n256_), .B(new_new_n255_), .C(new_new_n45_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n257_), .B(i_0_), .Y(new_new_n258_));
  OR3        g236(.A(new_new_n258_), .B(new_new_n254_), .C(new_new_n253_), .Y(new_new_n259_));
  NO2        g237(.A(i_1_), .B(new_new_n97_), .Y(new_new_n260_));
  NAi21      g238(.An(i_3_), .B(i_4_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n261_), .B(i_9_), .Y(new_new_n262_));
  AN2        g240(.A(i_6_), .B(i_7_), .Y(new_new_n263_));
  OAI210     g241(.A0(new_new_n263_), .A1(new_new_n260_), .B0(new_new_n262_), .Y(new_new_n264_));
  NA2        g242(.A(i_2_), .B(i_7_), .Y(new_new_n265_));
  NO2        g243(.A(new_new_n261_), .B(i_10_), .Y(new_new_n266_));
  NO2        g244(.A(new_new_n264_), .B(new_new_n151_), .Y(new_new_n267_));
  AOI210     g245(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n268_));
  OAI210     g246(.A0(new_new_n268_), .A1(new_new_n154_), .B0(new_new_n266_), .Y(new_new_n269_));
  AOI220     g247(.A0(new_new_n266_), .A1(new_new_n242_), .B0(new_new_n191_), .B1(new_new_n154_), .Y(new_new_n270_));
  AOI210     g248(.A0(new_new_n270_), .A1(new_new_n269_), .B0(i_5_), .Y(new_new_n271_));
  NO3        g249(.A(new_new_n271_), .B(new_new_n267_), .C(new_new_n259_), .Y(new_new_n272_));
  NO2        g250(.A(new_new_n272_), .B(new_new_n250_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n56_), .B(new_new_n25_), .Y(new_new_n274_));
  AN2        g252(.A(i_12_), .B(i_5_), .Y(new_new_n275_));
  NO2        g253(.A(i_4_), .B(new_new_n26_), .Y(new_new_n276_));
  NA2        g254(.A(new_new_n276_), .B(new_new_n275_), .Y(new_new_n277_));
  NO2        g255(.A(i_11_), .B(i_6_), .Y(new_new_n278_));
  NA3        g256(.A(new_new_n278_), .B(new_new_n234_), .C(new_new_n182_), .Y(new_new_n279_));
  NO2        g257(.A(new_new_n279_), .B(new_new_n277_), .Y(new_new_n280_));
  NO2        g258(.A(i_5_), .B(i_10_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n281_), .B(new_new_n214_), .Y(new_new_n282_));
  NA2        g260(.A(new_new_n132_), .B(new_new_n44_), .Y(new_new_n283_));
  NO2        g261(.A(new_new_n283_), .B(new_new_n282_), .Y(new_new_n284_));
  OAI210     g262(.A0(new_new_n284_), .A1(new_new_n280_), .B0(new_new_n274_), .Y(new_new_n285_));
  NO2        g263(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n286_));
  NO2        g264(.A(new_new_n138_), .B(new_new_n81_), .Y(new_new_n287_));
  OAI210     g265(.A0(new_new_n287_), .A1(new_new_n280_), .B0(new_new_n286_), .Y(new_new_n288_));
  NA3        g266(.A(new_new_n224_), .B(new_new_n88_), .C(new_new_n70_), .Y(new_new_n289_));
  NO2        g267(.A(i_11_), .B(i_12_), .Y(new_new_n290_));
  NA2        g268(.A(new_new_n290_), .B(new_new_n36_), .Y(new_new_n291_));
  NO2        g269(.A(new_new_n289_), .B(new_new_n291_), .Y(new_new_n292_));
  NA2        g270(.A(new_new_n281_), .B(new_new_n189_), .Y(new_new_n293_));
  NAi21      g271(.An(i_13_), .B(i_0_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n294_), .B(new_new_n192_), .Y(new_new_n295_));
  NA2        g273(.A(new_new_n292_), .B(new_new_n295_), .Y(new_new_n296_));
  NA3        g274(.A(new_new_n296_), .B(new_new_n288_), .C(new_new_n285_), .Y(new_new_n297_));
  NA2        g275(.A(new_new_n43_), .B(new_new_n182_), .Y(new_new_n298_));
  NO2        g276(.A(i_0_), .B(i_11_), .Y(new_new_n299_));
  NOi21      g277(.An(i_2_), .B(i_12_), .Y(new_new_n300_));
  NAi21      g278(.An(i_9_), .B(i_4_), .Y(new_new_n301_));
  OR2        g279(.A(i_13_), .B(i_10_), .Y(new_new_n302_));
  NO2        g280(.A(new_new_n146_), .B(new_new_n114_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n97_), .B(new_new_n25_), .Y(new_new_n304_));
  NA2        g282(.A(new_new_n157_), .B(i_10_), .Y(new_new_n305_));
  NA3        g283(.A(new_new_n202_), .B(new_new_n59_), .C(i_2_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(new_new_n305_), .Y(new_new_n307_));
  NA2        g285(.A(i_8_), .B(new_new_n233_), .Y(new_new_n308_));
  NO2        g286(.A(new_new_n308_), .B(new_new_n155_), .Y(new_new_n309_));
  NO2        g287(.A(new_new_n309_), .B(new_new_n307_), .Y(new_new_n310_));
  NO2        g288(.A(new_new_n310_), .B(new_new_n216_), .Y(new_new_n311_));
  NO3        g289(.A(new_new_n311_), .B(new_new_n297_), .C(new_new_n273_), .Y(new_new_n312_));
  NO2        g290(.A(i_10_), .B(i_9_), .Y(new_new_n313_));
  NAi21      g291(.An(i_12_), .B(i_8_), .Y(new_new_n314_));
  NO2        g292(.A(new_new_n314_), .B(i_3_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n45_), .B(i_4_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n100_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n317_), .B(new_new_n166_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n228_), .B(i_0_), .Y(new_new_n319_));
  NO3        g297(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n320_));
  NA2        g298(.A(new_new_n211_), .B(new_new_n95_), .Y(new_new_n321_));
  NA2        g299(.A(new_new_n321_), .B(new_new_n320_), .Y(new_new_n322_));
  NA2        g300(.A(i_8_), .B(i_9_), .Y(new_new_n323_));
  NO2        g301(.A(i_7_), .B(i_2_), .Y(new_new_n324_));
  OR2        g302(.A(new_new_n324_), .B(new_new_n323_), .Y(new_new_n325_));
  NA2        g303(.A(new_new_n222_), .B(new_new_n167_), .Y(new_new_n326_));
  OAI220     g304(.A0(new_new_n326_), .A1(new_new_n325_), .B0(new_new_n322_), .B1(new_new_n319_), .Y(new_new_n327_));
  NO3        g305(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n327_), .B(new_new_n318_), .Y(new_new_n329_));
  BUFFER     g307(.A(new_new_n246_), .Y(new_new_n330_));
  OR2        g308(.A(new_new_n330_), .B(new_new_n143_), .Y(new_new_n331_));
  NA2        g309(.A(new_new_n94_), .B(i_13_), .Y(new_new_n332_));
  NA2        g310(.A(i_5_), .B(new_new_n274_), .Y(new_new_n333_));
  NO2        g311(.A(i_2_), .B(i_13_), .Y(new_new_n334_));
  NO2        g312(.A(new_new_n333_), .B(new_new_n332_), .Y(new_new_n335_));
  NO3        g313(.A(i_4_), .B(new_new_n47_), .C(i_8_), .Y(new_new_n336_));
  NO2        g314(.A(i_6_), .B(i_7_), .Y(new_new_n337_));
  NO2        g315(.A(i_11_), .B(i_1_), .Y(new_new_n338_));
  NO2        g316(.A(i_3_), .B(new_new_n157_), .Y(new_new_n339_));
  NO2        g317(.A(i_6_), .B(i_10_), .Y(new_new_n340_));
  NA3        g318(.A(new_new_n196_), .B(new_new_n145_), .C(new_new_n123_), .Y(new_new_n341_));
  NA3        g319(.A(new_new_n286_), .B(new_new_n150_), .C(new_new_n137_), .Y(new_new_n342_));
  NA2        g320(.A(new_new_n342_), .B(new_new_n341_), .Y(new_new_n343_));
  NO2        g321(.A(new_new_n343_), .B(new_new_n335_), .Y(new_new_n344_));
  NA2        g322(.A(new_new_n320_), .B(new_new_n275_), .Y(new_new_n345_));
  NA2        g323(.A(new_new_n328_), .B(new_new_n281_), .Y(new_new_n346_));
  NO2        g324(.A(new_new_n346_), .B(new_new_n181_), .Y(new_new_n347_));
  NAi21      g325(.An(new_new_n174_), .B(new_new_n290_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n242_), .B(new_new_n176_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(new_new_n348_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n230_), .B(new_new_n191_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n351_), .B(new_new_n306_), .Y(new_new_n352_));
  NO3        g330(.A(new_new_n352_), .B(new_new_n350_), .C(new_new_n347_), .Y(new_new_n353_));
  NA4        g331(.A(new_new_n353_), .B(new_new_n344_), .C(new_new_n331_), .D(new_new_n329_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n113_), .B(new_new_n108_), .Y(new_new_n355_));
  AN2        g333(.A(new_new_n355_), .B(new_new_n320_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n356_), .B(new_new_n228_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n275_), .B(new_new_n182_), .Y(new_new_n358_));
  NA2        g336(.A(new_new_n249_), .B(new_new_n68_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n263_), .B(new_new_n255_), .Y(new_new_n360_));
  OR2        g338(.A(new_new_n358_), .B(new_new_n360_), .Y(new_new_n361_));
  NO2        g339(.A(new_new_n36_), .B(i_8_), .Y(new_new_n362_));
  INV        g340(.A(new_new_n361_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n202_), .B(new_new_n59_), .Y(new_new_n364_));
  OAI210     g342(.A0(i_8_), .A1(new_new_n364_), .B0(new_new_n125_), .Y(new_new_n365_));
  NA2        g343(.A(new_new_n365_), .B(new_new_n303_), .Y(new_new_n366_));
  NA3        g344(.A(new_new_n366_), .B(new_new_n361_), .C(new_new_n357_), .Y(new_new_n367_));
  NO2        g345(.A(i_12_), .B(new_new_n157_), .Y(new_new_n368_));
  NO2        g346(.A(i_8_), .B(i_7_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n43_), .B(i_10_), .Y(new_new_n370_));
  NO2        g348(.A(new_new_n370_), .B(i_6_), .Y(new_new_n371_));
  AOI220     g349(.A0(i_5_), .A1(new_new_n234_), .B0(i_2_), .B1(new_new_n195_), .Y(new_new_n372_));
  OAI220     g350(.A0(new_new_n372_), .A1(new_new_n208_), .B0(new_new_n332_), .B1(new_new_n124_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n373_), .B(new_new_n210_), .Y(new_new_n374_));
  NA3        g352(.A(new_new_n226_), .B(new_new_n147_), .C(new_new_n94_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n140_), .B(i_5_), .Y(new_new_n376_));
  NA3        g354(.A(new_new_n376_), .B(new_new_n298_), .C(new_new_n231_), .Y(new_new_n377_));
  NA2        g355(.A(new_new_n377_), .B(new_new_n375_), .Y(new_new_n378_));
  NA2        g356(.A(new_new_n378_), .B(new_new_n328_), .Y(new_new_n379_));
  NA2        g357(.A(new_new_n379_), .B(new_new_n374_), .Y(new_new_n380_));
  AOI210     g358(.A0(new_new_n256_), .A1(new_new_n45_), .B0(new_new_n260_), .Y(new_new_n381_));
  NA2        g359(.A(i_0_), .B(new_new_n47_), .Y(new_new_n382_));
  NA3        g360(.A(new_new_n368_), .B(new_new_n219_), .C(new_new_n382_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n381_), .B(new_new_n383_), .Y(new_new_n384_));
  INV        g362(.A(new_new_n384_), .Y(new_new_n385_));
  NO4        g363(.A(new_new_n198_), .B(new_new_n41_), .C(i_2_), .D(new_new_n47_), .Y(new_new_n386_));
  NO3        g364(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n387_));
  NOi21      g365(.An(i_10_), .B(i_6_), .Y(new_new_n388_));
  NO2        g366(.A(new_new_n81_), .B(new_new_n25_), .Y(new_new_n389_));
  AOI220     g367(.A0(new_new_n222_), .A1(new_new_n389_), .B0(new_new_n219_), .B1(new_new_n388_), .Y(new_new_n390_));
  NO2        g368(.A(new_new_n390_), .B(new_new_n319_), .Y(new_new_n391_));
  NO2        g369(.A(new_new_n109_), .B(new_new_n23_), .Y(new_new_n392_));
  NO2        g370(.A(new_new_n160_), .B(new_new_n37_), .Y(new_new_n393_));
  NOi31      g371(.An(new_new_n134_), .B(new_new_n393_), .C(new_new_n239_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n394_), .B(new_new_n391_), .Y(new_new_n395_));
  NO2        g373(.A(new_new_n359_), .B(new_new_n270_), .Y(new_new_n396_));
  INV        g374(.A(new_new_n231_), .Y(new_new_n397_));
  NO2        g375(.A(i_12_), .B(new_new_n81_), .Y(new_new_n398_));
  NA3        g376(.A(new_new_n398_), .B(new_new_n219_), .C(new_new_n382_), .Y(new_new_n399_));
  NA3        g377(.A(new_new_n278_), .B(new_new_n222_), .C(new_new_n176_), .Y(new_new_n400_));
  AOI210     g378(.A0(new_new_n400_), .A1(new_new_n399_), .B0(new_new_n397_), .Y(new_new_n401_));
  OR2        g379(.A(i_2_), .B(i_5_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n265_), .B(new_new_n195_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n403_), .B(new_new_n348_), .Y(new_new_n404_));
  NO3        g382(.A(new_new_n404_), .B(new_new_n401_), .C(new_new_n396_), .Y(new_new_n405_));
  NA3        g383(.A(new_new_n405_), .B(new_new_n395_), .C(new_new_n385_), .Y(new_new_n406_));
  NO4        g384(.A(new_new_n406_), .B(new_new_n380_), .C(new_new_n367_), .D(new_new_n354_), .Y(new_new_n407_));
  NA4        g385(.A(new_new_n407_), .B(new_new_n312_), .C(new_new_n248_), .D(new_new_n229_), .Y(ori7));
  NO2        g386(.A(new_new_n104_), .B(new_new_n87_), .Y(new_new_n409_));
  NA2        g387(.A(new_new_n276_), .B(new_new_n409_), .Y(new_new_n410_));
  NA2        g388(.A(new_new_n340_), .B(new_new_n79_), .Y(new_new_n411_));
  NA2        g389(.A(i_11_), .B(new_new_n157_), .Y(new_new_n412_));
  NA2        g390(.A(new_new_n132_), .B(new_new_n412_), .Y(new_new_n413_));
  OAI210     g391(.A0(new_new_n413_), .A1(new_new_n411_), .B0(new_new_n410_), .Y(new_new_n414_));
  NO2        g392(.A(new_new_n189_), .B(i_4_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(i_8_), .Y(new_new_n416_));
  NA2        g394(.A(i_2_), .B(new_new_n81_), .Y(new_new_n417_));
  OAI210     g395(.A0(new_new_n84_), .A1(new_new_n164_), .B0(new_new_n165_), .Y(new_new_n418_));
  NO2        g396(.A(i_7_), .B(new_new_n37_), .Y(new_new_n419_));
  NO2        g397(.A(new_new_n418_), .B(i_13_), .Y(new_new_n420_));
  NO2        g398(.A(new_new_n420_), .B(new_new_n414_), .Y(new_new_n421_));
  AOI210     g399(.A0(new_new_n119_), .A1(new_new_n57_), .B0(i_10_), .Y(new_new_n422_));
  AOI210     g400(.A0(new_new_n422_), .A1(new_new_n189_), .B0(new_new_n142_), .Y(new_new_n423_));
  OR2        g401(.A(i_6_), .B(i_10_), .Y(new_new_n424_));
  INV        g402(.A(new_new_n161_), .Y(new_new_n425_));
  OR2        g403(.A(new_new_n423_), .B(new_new_n212_), .Y(new_new_n426_));
  AOI210     g404(.A0(new_new_n426_), .A1(new_new_n421_), .B0(new_new_n58_), .Y(new_new_n427_));
  NOi21      g405(.An(i_11_), .B(i_7_), .Y(new_new_n428_));
  AO210      g406(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n429_));
  NO2        g407(.A(new_new_n429_), .B(new_new_n428_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n430_), .B(new_new_n168_), .Y(new_new_n431_));
  NA3        g409(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n432_));
  NAi21      g410(.An(new_new_n432_), .B(i_11_), .Y(new_new_n433_));
  AOI210     g411(.A0(new_new_n433_), .A1(new_new_n431_), .B0(new_new_n58_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n83_), .B(new_new_n58_), .Y(new_new_n435_));
  AO210      g413(.A0(new_new_n435_), .A1(new_new_n270_), .B0(new_new_n40_), .Y(new_new_n436_));
  NO3        g414(.A(new_new_n204_), .B(new_new_n169_), .C(new_new_n412_), .Y(new_new_n437_));
  OAI210     g415(.A0(new_new_n437_), .A1(new_new_n183_), .B0(new_new_n58_), .Y(new_new_n438_));
  NO2        g416(.A(new_new_n58_), .B(i_9_), .Y(new_new_n439_));
  NO2        g417(.A(i_1_), .B(i_12_), .Y(new_new_n440_));
  NA3        g418(.A(new_new_n440_), .B(new_new_n106_), .C(new_new_n24_), .Y(new_new_n441_));
  BUFFER     g419(.A(new_new_n441_), .Y(new_new_n442_));
  NA3        g420(.A(new_new_n442_), .B(new_new_n438_), .C(new_new_n436_), .Y(new_new_n443_));
  OAI210     g421(.A0(new_new_n443_), .A1(new_new_n434_), .B0(i_6_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n432_), .B(new_new_n104_), .Y(new_new_n445_));
  NA2        g423(.A(new_new_n445_), .B(new_new_n398_), .Y(new_new_n446_));
  NO2        g424(.A(i_6_), .B(i_11_), .Y(new_new_n447_));
  NA2        g425(.A(new_new_n446_), .B(new_new_n322_), .Y(new_new_n448_));
  NO3        g426(.A(new_new_n424_), .B(new_new_n188_), .C(new_new_n23_), .Y(new_new_n449_));
  AOI210     g427(.A0(i_1_), .A1(new_new_n205_), .B0(new_new_n449_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n450_), .B(new_new_n43_), .Y(new_new_n451_));
  NA3        g429(.A(new_new_n369_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n452_));
  INV        g430(.A(i_2_), .Y(new_new_n453_));
  NA2        g431(.A(new_new_n129_), .B(i_9_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n45_), .B(i_1_), .Y(new_new_n455_));
  NO2        g433(.A(new_new_n454_), .B(new_new_n453_), .Y(new_new_n456_));
  NA3        g434(.A(new_new_n439_), .B(new_new_n231_), .C(i_6_), .Y(new_new_n457_));
  NO2        g435(.A(new_new_n457_), .B(new_new_n23_), .Y(new_new_n458_));
  AOI210     g436(.A0(new_new_n338_), .A1(new_new_n304_), .B0(new_new_n193_), .Y(new_new_n459_));
  NO2        g437(.A(new_new_n459_), .B(new_new_n417_), .Y(new_new_n460_));
  NAi21      g438(.An(new_new_n452_), .B(new_new_n89_), .Y(new_new_n461_));
  NA2        g439(.A(new_new_n455_), .B(new_new_n211_), .Y(new_new_n462_));
  NO2        g440(.A(i_11_), .B(new_new_n37_), .Y(new_new_n463_));
  NA2        g441(.A(new_new_n463_), .B(new_new_n24_), .Y(new_new_n464_));
  OAI210     g442(.A0(new_new_n464_), .A1(new_new_n462_), .B0(new_new_n461_), .Y(new_new_n465_));
  OR4        g443(.A(new_new_n465_), .B(new_new_n460_), .C(new_new_n458_), .D(new_new_n456_), .Y(new_new_n466_));
  NO3        g444(.A(new_new_n466_), .B(new_new_n451_), .C(new_new_n448_), .Y(new_new_n467_));
  NO2        g445(.A(i_12_), .B(new_new_n428_), .Y(new_new_n468_));
  NO2        g446(.A(new_new_n301_), .B(new_new_n81_), .Y(new_new_n469_));
  NA2        g447(.A(i_3_), .B(new_new_n157_), .Y(new_new_n470_));
  NO2        g448(.A(new_new_n470_), .B(new_new_n109_), .Y(new_new_n471_));
  AN2        g449(.A(new_new_n471_), .B(new_new_n371_), .Y(new_new_n472_));
  NO2        g450(.A(new_new_n188_), .B(new_new_n43_), .Y(new_new_n473_));
  NO3        g451(.A(new_new_n473_), .B(new_new_n228_), .C(new_new_n190_), .Y(new_new_n474_));
  NO2        g452(.A(new_new_n110_), .B(new_new_n37_), .Y(new_new_n475_));
  NO2        g453(.A(new_new_n475_), .B(i_6_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n81_), .B(i_9_), .Y(new_new_n477_));
  NO2        g455(.A(new_new_n477_), .B(new_new_n58_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n478_), .B(new_new_n440_), .Y(new_new_n479_));
  NO4        g457(.A(new_new_n479_), .B(new_new_n476_), .C(new_new_n474_), .D(i_4_), .Y(new_new_n480_));
  NA2        g458(.A(i_1_), .B(i_3_), .Y(new_new_n481_));
  NO2        g459(.A(new_new_n323_), .B(new_new_n90_), .Y(new_new_n482_));
  AOI210     g460(.A0(new_new_n473_), .A1(new_new_n388_), .B0(new_new_n482_), .Y(new_new_n483_));
  NO2        g461(.A(new_new_n483_), .B(new_new_n481_), .Y(new_new_n484_));
  NO3        g462(.A(new_new_n484_), .B(new_new_n480_), .C(new_new_n472_), .Y(new_new_n485_));
  NA3        g463(.A(new_new_n485_), .B(new_new_n467_), .C(new_new_n444_), .Y(new_new_n486_));
  NA2        g464(.A(new_new_n263_), .B(new_new_n262_), .Y(new_new_n487_));
  NA3        g465(.A(new_new_n340_), .B(new_new_n362_), .C(new_new_n45_), .Y(new_new_n488_));
  NA3        g466(.A(new_new_n142_), .B(new_new_n79_), .C(new_new_n81_), .Y(new_new_n489_));
  NA3        g467(.A(new_new_n489_), .B(new_new_n488_), .C(new_new_n487_), .Y(new_new_n490_));
  NA2        g468(.A(new_new_n490_), .B(i_1_), .Y(new_new_n491_));
  AOI210     g469(.A0(new_new_n211_), .A1(new_new_n95_), .B0(i_1_), .Y(new_new_n492_));
  NO2        g470(.A(new_new_n261_), .B(i_2_), .Y(new_new_n493_));
  NA2        g471(.A(new_new_n493_), .B(new_new_n492_), .Y(new_new_n494_));
  OAI210     g472(.A0(new_new_n457_), .A1(new_new_n314_), .B0(new_new_n494_), .Y(new_new_n495_));
  INV        g473(.A(new_new_n495_), .Y(new_new_n496_));
  AOI210     g474(.A0(new_new_n496_), .A1(new_new_n491_), .B0(i_13_), .Y(new_new_n497_));
  OR2        g475(.A(i_11_), .B(i_7_), .Y(new_new_n498_));
  NA3        g476(.A(new_new_n498_), .B(new_new_n102_), .C(new_new_n129_), .Y(new_new_n499_));
  AOI220     g477(.A0(new_new_n334_), .A1(new_new_n142_), .B0(new_new_n316_), .B1(new_new_n129_), .Y(new_new_n500_));
  OAI210     g478(.A0(new_new_n500_), .A1(new_new_n43_), .B0(new_new_n499_), .Y(new_new_n501_));
  NO2        g479(.A(new_new_n52_), .B(i_12_), .Y(new_new_n502_));
  INV        g480(.A(new_new_n502_), .Y(new_new_n503_));
  NA2        g481(.A(i_7_), .B(new_new_n469_), .Y(new_new_n504_));
  OAI220     g482(.A0(new_new_n504_), .A1(new_new_n40_), .B0(new_new_n503_), .B1(new_new_n90_), .Y(new_new_n505_));
  AOI210     g483(.A0(new_new_n501_), .A1(new_new_n241_), .B0(new_new_n505_), .Y(new_new_n506_));
  INV        g484(.A(new_new_n109_), .Y(new_new_n507_));
  AOI220     g485(.A0(new_new_n507_), .A1(new_new_n67_), .B0(new_new_n278_), .B1(new_new_n455_), .Y(new_new_n508_));
  NO2        g486(.A(new_new_n508_), .B(new_new_n194_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n118_), .B(i_13_), .Y(new_new_n510_));
  NO2        g488(.A(new_new_n510_), .B(new_new_n492_), .Y(new_new_n511_));
  NO3        g489(.A(new_new_n66_), .B(new_new_n32_), .C(new_new_n97_), .Y(new_new_n512_));
  AOI220     g490(.A0(new_new_n278_), .A1(new_new_n455_), .B0(new_new_n89_), .B1(new_new_n98_), .Y(new_new_n513_));
  OAI220     g491(.A0(new_new_n513_), .A1(new_new_n416_), .B0(new_new_n765_), .B1(new_new_n425_), .Y(new_new_n514_));
  NO3        g492(.A(new_new_n514_), .B(new_new_n511_), .C(new_new_n509_), .Y(new_new_n515_));
  NA3        g493(.A(new_new_n300_), .B(new_new_n419_), .C(new_new_n95_), .Y(new_new_n516_));
  NA2        g494(.A(new_new_n447_), .B(i_13_), .Y(new_new_n517_));
  NAi21      g495(.An(i_11_), .B(i_12_), .Y(new_new_n518_));
  NOi41      g496(.An(new_new_n107_), .B(new_new_n518_), .C(i_13_), .D(new_new_n81_), .Y(new_new_n519_));
  INV        g497(.A(new_new_n519_), .Y(new_new_n520_));
  NA3        g498(.A(new_new_n520_), .B(new_new_n517_), .C(new_new_n516_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n521_), .B(new_new_n58_), .Y(new_new_n522_));
  NO2        g500(.A(i_2_), .B(i_12_), .Y(new_new_n523_));
  NA2        g501(.A(new_new_n260_), .B(new_new_n523_), .Y(new_new_n524_));
  NA2        g502(.A(i_8_), .B(new_new_n25_), .Y(new_new_n525_));
  NO2        g503(.A(new_new_n525_), .B(new_new_n276_), .Y(new_new_n526_));
  OAI210     g504(.A0(new_new_n526_), .A1(new_new_n262_), .B0(new_new_n260_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n527_), .B(new_new_n524_), .Y(new_new_n528_));
  NA3        g506(.A(new_new_n528_), .B(new_new_n44_), .C(new_new_n182_), .Y(new_new_n529_));
  NA4        g507(.A(new_new_n529_), .B(new_new_n522_), .C(new_new_n515_), .D(new_new_n506_), .Y(new_new_n530_));
  OR4        g508(.A(new_new_n530_), .B(new_new_n497_), .C(new_new_n486_), .D(new_new_n427_), .Y(ori5));
  NA2        g509(.A(new_new_n468_), .B(new_new_n214_), .Y(new_new_n532_));
  AN2        g510(.A(new_new_n24_), .B(i_10_), .Y(new_new_n533_));
  NA3        g511(.A(new_new_n533_), .B(new_new_n523_), .C(new_new_n104_), .Y(new_new_n534_));
  NO2        g512(.A(new_new_n416_), .B(i_11_), .Y(new_new_n535_));
  NA2        g513(.A(new_new_n84_), .B(new_new_n535_), .Y(new_new_n536_));
  NA3        g514(.A(new_new_n536_), .B(new_new_n534_), .C(new_new_n532_), .Y(new_new_n537_));
  NO3        g515(.A(i_11_), .B(new_new_n189_), .C(i_13_), .Y(new_new_n538_));
  NO2        g516(.A(new_new_n115_), .B(new_new_n23_), .Y(new_new_n539_));
  NA2        g517(.A(i_12_), .B(i_8_), .Y(new_new_n540_));
  INV        g518(.A(new_new_n313_), .Y(new_new_n541_));
  AOI220     g519(.A0(new_new_n231_), .A1(new_new_n392_), .B0(i_12_), .B1(new_new_n539_), .Y(new_new_n542_));
  INV        g520(.A(new_new_n542_), .Y(new_new_n543_));
  NO2        g521(.A(new_new_n543_), .B(new_new_n537_), .Y(new_new_n544_));
  INV        g522(.A(new_new_n145_), .Y(new_new_n545_));
  INV        g523(.A(new_new_n196_), .Y(new_new_n546_));
  OAI210     g524(.A0(new_new_n493_), .A1(new_new_n315_), .B0(new_new_n107_), .Y(new_new_n547_));
  AOI210     g525(.A0(new_new_n547_), .A1(new_new_n546_), .B0(new_new_n545_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n323_), .B(new_new_n26_), .Y(new_new_n549_));
  NO2        g527(.A(new_new_n549_), .B(new_new_n304_), .Y(new_new_n550_));
  NA2        g528(.A(new_new_n550_), .B(i_2_), .Y(new_new_n551_));
  INV        g529(.A(new_new_n551_), .Y(new_new_n552_));
  AOI210     g530(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n302_), .Y(new_new_n553_));
  AOI210     g531(.A0(new_new_n553_), .A1(new_new_n552_), .B0(new_new_n548_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n156_), .B(new_new_n116_), .Y(new_new_n555_));
  OAI210     g533(.A0(new_new_n555_), .A1(new_new_n539_), .B0(i_2_), .Y(new_new_n556_));
  INV        g534(.A(new_new_n146_), .Y(new_new_n557_));
  NA2        g535(.A(new_new_n557_), .B(new_new_n84_), .Y(new_new_n558_));
  AOI210     g536(.A0(new_new_n558_), .A1(new_new_n556_), .B0(new_new_n157_), .Y(new_new_n559_));
  OA210      g537(.A0(new_new_n430_), .A1(new_new_n117_), .B0(i_13_), .Y(new_new_n560_));
  NA2        g538(.A(new_new_n161_), .B(new_new_n164_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n561_), .B(new_new_n265_), .Y(new_new_n562_));
  AOI210     g540(.A0(new_new_n169_), .A1(new_new_n136_), .B0(new_new_n362_), .Y(new_new_n563_));
  NA2        g541(.A(new_new_n563_), .B(new_new_n304_), .Y(new_new_n564_));
  NO2        g542(.A(new_new_n98_), .B(new_new_n43_), .Y(new_new_n565_));
  INV        g543(.A(new_new_n225_), .Y(new_new_n566_));
  NA4        g544(.A(new_new_n566_), .B(new_new_n226_), .C(new_new_n115_), .D(new_new_n41_), .Y(new_new_n567_));
  OAI210     g545(.A0(new_new_n567_), .A1(new_new_n565_), .B0(new_new_n564_), .Y(new_new_n568_));
  NO4        g546(.A(new_new_n568_), .B(new_new_n562_), .C(new_new_n560_), .D(new_new_n559_), .Y(new_new_n569_));
  NO2        g547(.A(new_new_n57_), .B(i_12_), .Y(new_new_n570_));
  NO2        g548(.A(new_new_n570_), .B(new_new_n117_), .Y(new_new_n571_));
  NO2        g549(.A(new_new_n571_), .B(new_new_n412_), .Y(new_new_n572_));
  NA2        g550(.A(new_new_n572_), .B(new_new_n36_), .Y(new_new_n573_));
  NA4        g551(.A(new_new_n573_), .B(new_new_n569_), .C(new_new_n554_), .D(new_new_n544_), .Y(ori6));
  NA4        g552(.A(new_new_n281_), .B(new_new_n339_), .C(new_new_n66_), .D(new_new_n97_), .Y(new_new_n575_));
  INV        g553(.A(new_new_n575_), .Y(new_new_n576_));
  NO2        g554(.A(i_11_), .B(i_9_), .Y(new_new_n577_));
  NO2        g555(.A(new_new_n576_), .B(new_new_n236_), .Y(new_new_n578_));
  OR2        g556(.A(new_new_n578_), .B(i_12_), .Y(new_new_n579_));
  NA2        g557(.A(new_new_n266_), .B(new_new_n242_), .Y(new_new_n580_));
  NA2        g558(.A(new_new_n398_), .B(new_new_n58_), .Y(new_new_n581_));
  BUFFER     g559(.A(new_new_n435_), .Y(new_new_n582_));
  NA3        g560(.A(new_new_n582_), .B(new_new_n581_), .C(new_new_n580_), .Y(new_new_n583_));
  INV        g561(.A(new_new_n159_), .Y(new_new_n584_));
  AOI220     g562(.A0(new_new_n584_), .A1(new_new_n577_), .B0(new_new_n583_), .B1(new_new_n68_), .Y(new_new_n585_));
  INV        g563(.A(new_new_n235_), .Y(new_new_n586_));
  NA2        g564(.A(new_new_n70_), .B(new_new_n122_), .Y(new_new_n587_));
  INV        g565(.A(new_new_n115_), .Y(new_new_n588_));
  NA2        g566(.A(new_new_n588_), .B(new_new_n45_), .Y(new_new_n589_));
  AOI210     g567(.A0(new_new_n589_), .A1(new_new_n587_), .B0(new_new_n586_), .Y(new_new_n590_));
  NO2        g568(.A(new_new_n198_), .B(i_9_), .Y(new_new_n591_));
  NA2        g569(.A(new_new_n591_), .B(new_new_n570_), .Y(new_new_n592_));
  AOI210     g570(.A0(new_new_n592_), .A1(new_new_n360_), .B0(new_new_n151_), .Y(new_new_n593_));
  NO2        g571(.A(new_new_n32_), .B(i_11_), .Y(new_new_n594_));
  NA3        g572(.A(new_new_n594_), .B(new_new_n337_), .C(new_new_n281_), .Y(new_new_n595_));
  INV        g573(.A(new_new_n595_), .Y(new_new_n596_));
  OR3        g574(.A(new_new_n596_), .B(new_new_n593_), .C(new_new_n590_), .Y(new_new_n597_));
  OR2        g575(.A(new_new_n430_), .B(new_new_n315_), .Y(new_new_n598_));
  NA3        g576(.A(new_new_n598_), .B(new_new_n135_), .C(new_new_n64_), .Y(new_new_n599_));
  AO210      g577(.A0(new_new_n346_), .A1(new_new_n541_), .B0(new_new_n36_), .Y(new_new_n600_));
  NA2        g578(.A(new_new_n600_), .B(new_new_n599_), .Y(new_new_n601_));
  OAI210     g579(.A0(i_6_), .A1(i_11_), .B0(new_new_n82_), .Y(new_new_n602_));
  NA2        g580(.A(new_new_n602_), .B(new_new_n387_), .Y(new_new_n603_));
  NA3        g581(.A(new_new_n265_), .B(new_new_n191_), .C(new_new_n135_), .Y(new_new_n604_));
  NA3        g582(.A(new_new_n604_), .B(new_new_n603_), .C(new_new_n418_), .Y(new_new_n605_));
  AO210      g583(.A0(new_new_n362_), .A1(new_new_n45_), .B0(new_new_n83_), .Y(new_new_n606_));
  NA3        g584(.A(new_new_n606_), .B(new_new_n340_), .C(new_new_n176_), .Y(new_new_n607_));
  AOI210     g585(.A0(new_new_n315_), .A1(new_new_n313_), .B0(new_new_n386_), .Y(new_new_n608_));
  NO2        g586(.A(new_new_n424_), .B(new_new_n98_), .Y(new_new_n609_));
  OAI210     g587(.A0(new_new_n609_), .A1(new_new_n108_), .B0(new_new_n299_), .Y(new_new_n610_));
  NA3        g588(.A(new_new_n610_), .B(new_new_n608_), .C(new_new_n607_), .Y(new_new_n611_));
  NO4        g589(.A(new_new_n611_), .B(new_new_n605_), .C(new_new_n601_), .D(new_new_n597_), .Y(new_new_n612_));
  NA4        g590(.A(new_new_n612_), .B(new_new_n585_), .C(new_new_n579_), .D(new_new_n272_), .Y(ori3));
  NA2        g591(.A(i_12_), .B(i_10_), .Y(new_new_n614_));
  NO2        g592(.A(i_11_), .B(new_new_n189_), .Y(new_new_n615_));
  NA3        g593(.A(new_new_n604_), .B(new_new_n418_), .C(new_new_n264_), .Y(new_new_n616_));
  NA2        g594(.A(new_new_n616_), .B(new_new_n39_), .Y(new_new_n617_));
  NOi21      g595(.An(new_new_n94_), .B(new_new_n550_), .Y(new_new_n618_));
  NA2        g596(.A(new_new_n300_), .B(new_new_n44_), .Y(new_new_n619_));
  AN2        g597(.A(new_new_n321_), .B(new_new_n53_), .Y(new_new_n620_));
  NO2        g598(.A(new_new_n620_), .B(new_new_n618_), .Y(new_new_n621_));
  AOI210     g599(.A0(new_new_n621_), .A1(new_new_n617_), .B0(new_new_n47_), .Y(new_new_n622_));
  NO4        g600(.A(new_new_n268_), .B(new_new_n275_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n623_));
  NA2        g601(.A(new_new_n151_), .B(new_new_n388_), .Y(new_new_n624_));
  NOi21      g602(.An(new_new_n624_), .B(new_new_n623_), .Y(new_new_n625_));
  NO2        g603(.A(new_new_n625_), .B(new_new_n58_), .Y(new_new_n626_));
  NO2        g604(.A(new_new_n626_), .B(new_new_n622_), .Y(new_new_n627_));
  NA2        g605(.A(new_new_n151_), .B(new_new_n24_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n475_), .B(new_new_n409_), .Y(new_new_n629_));
  NO2        g607(.A(new_new_n629_), .B(new_new_n628_), .Y(new_new_n630_));
  NA2        g608(.A(new_new_n230_), .B(new_new_n120_), .Y(new_new_n631_));
  NO2        g609(.A(new_new_n631_), .B(new_new_n293_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n632_), .B(new_new_n630_), .Y(new_new_n633_));
  NA2        g611(.A(new_new_n389_), .B(i_0_), .Y(new_new_n634_));
  NO3        g612(.A(new_new_n634_), .B(new_new_n277_), .C(new_new_n84_), .Y(new_new_n635_));
  NO3        g613(.A(new_new_n402_), .B(new_new_n173_), .C(new_new_n302_), .Y(new_new_n636_));
  AOI210     g614(.A0(new_new_n636_), .A1(i_11_), .B0(new_new_n635_), .Y(new_new_n637_));
  NA2        g615(.A(new_new_n538_), .B(new_new_n236_), .Y(new_new_n638_));
  AOI210     g616(.A0(new_new_n340_), .A1(new_new_n84_), .B0(new_new_n55_), .Y(new_new_n639_));
  NO2        g617(.A(new_new_n639_), .B(new_new_n638_), .Y(new_new_n640_));
  NO2        g618(.A(new_new_n200_), .B(new_new_n139_), .Y(new_new_n641_));
  NA2        g619(.A(i_0_), .B(i_10_), .Y(new_new_n642_));
  INV        g620(.A(new_new_n370_), .Y(new_new_n643_));
  NO3        g621(.A(new_new_n109_), .B(new_new_n470_), .C(i_5_), .Y(new_new_n644_));
  AO220      g622(.A0(new_new_n644_), .A1(new_new_n643_), .B0(new_new_n641_), .B1(i_6_), .Y(new_new_n645_));
  NO2        g623(.A(new_new_n645_), .B(new_new_n640_), .Y(new_new_n646_));
  NA3        g624(.A(new_new_n646_), .B(new_new_n637_), .C(new_new_n633_), .Y(new_new_n647_));
  NO2        g625(.A(new_new_n99_), .B(new_new_n37_), .Y(new_new_n648_));
  NA2        g626(.A(i_11_), .B(i_9_), .Y(new_new_n649_));
  NO3        g627(.A(i_12_), .B(new_new_n649_), .C(new_new_n417_), .Y(new_new_n650_));
  AN2        g628(.A(new_new_n650_), .B(new_new_n648_), .Y(new_new_n651_));
  NA2        g629(.A(new_new_n286_), .B(new_new_n150_), .Y(new_new_n652_));
  INV        g630(.A(new_new_n652_), .Y(new_new_n653_));
  NO2        g631(.A(new_new_n649_), .B(new_new_n68_), .Y(new_new_n654_));
  NO2        g632(.A(new_new_n148_), .B(i_0_), .Y(new_new_n655_));
  NO2        g633(.A(new_new_n653_), .B(new_new_n651_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n463_), .B(new_new_n112_), .Y(new_new_n657_));
  NO2        g635(.A(i_6_), .B(new_new_n657_), .Y(new_new_n658_));
  NA2        g636(.A(new_new_n145_), .B(new_new_n99_), .Y(new_new_n659_));
  NO2        g637(.A(new_new_n767_), .B(new_new_n619_), .Y(new_new_n660_));
  NO2        g638(.A(new_new_n660_), .B(new_new_n658_), .Y(new_new_n661_));
  NOi21      g639(.An(i_7_), .B(i_5_), .Y(new_new_n662_));
  NOi31      g640(.An(new_new_n662_), .B(i_0_), .C(new_new_n518_), .Y(new_new_n663_));
  NA3        g641(.A(new_new_n663_), .B(new_new_n276_), .C(i_6_), .Y(new_new_n664_));
  BUFFER     g642(.A(new_new_n664_), .Y(new_new_n665_));
  INV        g643(.A(new_new_n232_), .Y(new_new_n666_));
  NA3        g644(.A(new_new_n665_), .B(new_new_n661_), .C(new_new_n656_), .Y(new_new_n667_));
  NO2        g645(.A(new_new_n614_), .B(new_new_n231_), .Y(new_new_n668_));
  OA210      g646(.A0(new_new_n337_), .A1(new_new_n180_), .B0(new_new_n336_), .Y(new_new_n669_));
  NA2        g647(.A(new_new_n668_), .B(new_new_n654_), .Y(new_new_n670_));
  NA2        g648(.A(new_new_n654_), .B(new_new_n226_), .Y(new_new_n671_));
  OAI210     g649(.A0(i_3_), .A1(new_new_n153_), .B0(new_new_n671_), .Y(new_new_n672_));
  NA2        g650(.A(new_new_n672_), .B(new_new_n337_), .Y(new_new_n673_));
  NA3        g651(.A(i_5_), .B(new_new_n274_), .C(i_6_), .Y(new_new_n674_));
  NA2        g652(.A(new_new_n90_), .B(new_new_n43_), .Y(new_new_n675_));
  NO2        g653(.A(new_new_n70_), .B(new_new_n540_), .Y(new_new_n676_));
  AOI220     g654(.A0(new_new_n676_), .A1(new_new_n675_), .B0(new_new_n147_), .B1(new_new_n409_), .Y(new_new_n677_));
  AOI210     g655(.A0(new_new_n677_), .A1(new_new_n674_), .B0(new_new_n46_), .Y(new_new_n678_));
  NO3        g656(.A(new_new_n402_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n679_));
  AOI210     g657(.A0(i_7_), .A1(new_new_n376_), .B0(new_new_n679_), .Y(new_new_n680_));
  NAi21      g658(.An(i_9_), .B(i_5_), .Y(new_new_n681_));
  NO2        g659(.A(new_new_n681_), .B(new_new_n294_), .Y(new_new_n682_));
  NA2        g660(.A(new_new_n682_), .B(new_new_n430_), .Y(new_new_n683_));
  OAI220     g661(.A0(new_new_n683_), .A1(new_new_n81_), .B0(new_new_n680_), .B1(new_new_n146_), .Y(new_new_n684_));
  NO3        g662(.A(new_new_n684_), .B(new_new_n678_), .C(new_new_n363_), .Y(new_new_n685_));
  NA3        g663(.A(new_new_n685_), .B(new_new_n673_), .C(new_new_n670_), .Y(new_new_n686_));
  NO3        g664(.A(new_new_n686_), .B(new_new_n667_), .C(new_new_n647_), .Y(new_new_n687_));
  NO2        g665(.A(i_0_), .B(new_new_n518_), .Y(new_new_n688_));
  AOI210     g666(.A0(new_new_n581_), .A1(new_new_n487_), .B0(new_new_n659_), .Y(new_new_n689_));
  INV        g667(.A(new_new_n689_), .Y(new_new_n690_));
  NA2        g668(.A(new_new_n195_), .B(new_new_n187_), .Y(new_new_n691_));
  AOI210     g669(.A0(new_new_n691_), .A1(new_new_n634_), .B0(new_new_n139_), .Y(new_new_n692_));
  INV        g670(.A(new_new_n692_), .Y(new_new_n693_));
  NA2        g671(.A(new_new_n693_), .B(new_new_n690_), .Y(new_new_n694_));
  NO3        g672(.A(new_new_n642_), .B(i_5_), .C(new_new_n156_), .Y(new_new_n695_));
  NA2        g673(.A(new_new_n695_), .B(i_11_), .Y(new_new_n696_));
  NO3        g674(.A(new_new_n170_), .B(new_new_n275_), .C(i_0_), .Y(new_new_n697_));
  OAI210     g675(.A0(new_new_n697_), .A1(new_new_n71_), .B0(i_13_), .Y(new_new_n698_));
  NA2        g676(.A(new_new_n698_), .B(new_new_n696_), .Y(new_new_n699_));
  NO2        g677(.A(new_new_n194_), .B(new_new_n90_), .Y(new_new_n700_));
  AOI210     g678(.A0(new_new_n700_), .A1(new_new_n688_), .B0(new_new_n105_), .Y(new_new_n701_));
  OR2        g679(.A(new_new_n701_), .B(i_5_), .Y(new_new_n702_));
  AOI210     g680(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n148_), .Y(new_new_n703_));
  NA2        g681(.A(new_new_n703_), .B(new_new_n669_), .Y(new_new_n704_));
  NA2        g682(.A(new_new_n345_), .B(new_new_n341_), .Y(new_new_n705_));
  INV        g683(.A(new_new_n705_), .Y(new_new_n706_));
  NA3        g684(.A(new_new_n281_), .B(new_new_n145_), .C(new_new_n144_), .Y(new_new_n707_));
  NA3        g685(.A(i_5_), .B(new_new_n223_), .C(new_new_n187_), .Y(new_new_n708_));
  NA2        g686(.A(new_new_n708_), .B(new_new_n707_), .Y(new_new_n709_));
  NO3        g687(.A(new_new_n649_), .B(new_new_n176_), .C(new_new_n156_), .Y(new_new_n710_));
  NO2        g688(.A(new_new_n710_), .B(new_new_n709_), .Y(new_new_n711_));
  NA4        g689(.A(new_new_n711_), .B(new_new_n706_), .C(new_new_n704_), .D(new_new_n702_), .Y(new_new_n712_));
  NO2        g690(.A(new_new_n81_), .B(i_5_), .Y(new_new_n713_));
  NA3        g691(.A(new_new_n615_), .B(new_new_n106_), .C(new_new_n115_), .Y(new_new_n714_));
  INV        g692(.A(new_new_n714_), .Y(new_new_n715_));
  NA2        g693(.A(new_new_n715_), .B(new_new_n713_), .Y(new_new_n716_));
  NA2        g694(.A(new_new_n226_), .B(i_5_), .Y(new_new_n717_));
  NAi31      g695(.An(new_new_n193_), .B(new_new_n717_), .C(new_new_n194_), .Y(new_new_n718_));
  NO4        g696(.A(new_new_n192_), .B(new_new_n170_), .C(i_0_), .D(i_12_), .Y(new_new_n719_));
  AOI220     g697(.A0(new_new_n719_), .A1(new_new_n718_), .B0(new_new_n576_), .B1(new_new_n149_), .Y(new_new_n720_));
  AN2        g698(.A(new_new_n642_), .B(new_new_n139_), .Y(new_new_n721_));
  NO3        g699(.A(new_new_n721_), .B(i_12_), .C(new_new_n452_), .Y(new_new_n722_));
  NA2        g700(.A(new_new_n722_), .B(new_new_n176_), .Y(new_new_n723_));
  NA2        g701(.A(new_new_n662_), .B(new_new_n334_), .Y(new_new_n724_));
  NA2        g702(.A(new_new_n59_), .B(new_new_n97_), .Y(new_new_n725_));
  OAI220     g703(.A0(new_new_n725_), .A1(new_new_n717_), .B0(new_new_n724_), .B1(new_new_n478_), .Y(new_new_n726_));
  NA2        g704(.A(new_new_n726_), .B(new_new_n655_), .Y(new_new_n727_));
  NA4        g705(.A(new_new_n727_), .B(new_new_n723_), .C(new_new_n720_), .D(new_new_n716_), .Y(new_new_n728_));
  NO4        g706(.A(new_new_n728_), .B(new_new_n712_), .C(new_new_n699_), .D(new_new_n694_), .Y(new_new_n729_));
  NA2        g707(.A(new_new_n594_), .B(new_new_n37_), .Y(new_new_n730_));
  NA2        g708(.A(new_new_n730_), .B(new_new_n423_), .Y(new_new_n731_));
  NA2        g709(.A(new_new_n731_), .B(new_new_n168_), .Y(new_new_n732_));
  BUFFER     g710(.A(new_new_n498_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n152_), .B(new_new_n154_), .Y(new_new_n734_));
  AO210      g712(.A0(new_new_n733_), .A1(new_new_n33_), .B0(new_new_n734_), .Y(new_new_n735_));
  NAi31      g713(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n736_));
  NO2        g714(.A(new_new_n65_), .B(new_new_n736_), .Y(new_new_n737_));
  NO2        g715(.A(new_new_n737_), .B(new_new_n449_), .Y(new_new_n738_));
  NA2        g716(.A(new_new_n738_), .B(new_new_n735_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n739_), .A1(new_new_n47_), .B0(new_new_n636_), .Y(new_new_n740_));
  AOI210     g718(.A0(new_new_n740_), .A1(new_new_n732_), .B0(new_new_n68_), .Y(new_new_n741_));
  INV        g719(.A(new_new_n271_), .Y(new_new_n742_));
  NO2        g720(.A(new_new_n742_), .B(new_new_n545_), .Y(new_new_n743_));
  INV        g721(.A(new_new_n71_), .Y(new_new_n744_));
  AOI210     g722(.A0(new_new_n703_), .A1(i_5_), .B0(new_new_n663_), .Y(new_new_n745_));
  AOI210     g723(.A0(new_new_n745_), .A1(new_new_n744_), .B0(new_new_n481_), .Y(new_new_n746_));
  INV        g724(.A(new_new_n746_), .Y(new_new_n747_));
  NA2        g725(.A(new_new_n213_), .B(new_new_n84_), .Y(new_new_n748_));
  NA3        g726(.A(new_new_n549_), .B(new_new_n223_), .C(new_new_n75_), .Y(new_new_n749_));
  AOI210     g727(.A0(new_new_n749_), .A1(new_new_n748_), .B0(i_11_), .Y(new_new_n750_));
  NO3        g728(.A(new_new_n56_), .B(new_new_n55_), .C(i_4_), .Y(new_new_n751_));
  OAI210     g729(.A0(new_new_n666_), .A1(new_new_n227_), .B0(new_new_n751_), .Y(new_new_n752_));
  NO2        g730(.A(new_new_n752_), .B(new_new_n518_), .Y(new_new_n753_));
  NO4        g731(.A(new_new_n681_), .B(i_11_), .C(new_new_n199_), .D(new_new_n198_), .Y(new_new_n754_));
  NO2        g732(.A(new_new_n754_), .B(new_new_n386_), .Y(new_new_n755_));
  INV        g733(.A(new_new_n253_), .Y(new_new_n756_));
  AOI210     g734(.A0(new_new_n756_), .A1(new_new_n755_), .B0(new_new_n40_), .Y(new_new_n757_));
  NO3        g735(.A(new_new_n757_), .B(new_new_n753_), .C(new_new_n750_), .Y(new_new_n758_));
  OAI210     g736(.A0(new_new_n747_), .A1(i_4_), .B0(new_new_n758_), .Y(new_new_n759_));
  NO3        g737(.A(new_new_n759_), .B(new_new_n743_), .C(new_new_n741_), .Y(new_new_n760_));
  NA4        g738(.A(new_new_n760_), .B(new_new_n729_), .C(new_new_n687_), .D(new_new_n627_), .Y(ori4));
  INV        g739(.A(i_6_), .Y(new_new_n764_));
  INV        g740(.A(new_new_n512_), .Y(new_new_n765_));
  INV        g741(.A(i_8_), .Y(new_new_n766_));
  INV        g742(.A(new_new_n236_), .Y(new_new_n767_));
endmodule


