//Benchmark atmr_max1024_476_0.0156

module atmr_max1024(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, z0, z1, z2, z3, z4, z5);
 input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
 output z0, z1, z2, z3, z4, z5;
 wire ori_ori_n17_, ori_ori_n18_, ori_ori_n19_, ori_ori_n20_, ori_ori_n21_, ori_ori_n22_, ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, mai_mai_n17_, mai_mai_n18_, mai_mai_n19_, mai_mai_n20_, mai_mai_n21_, mai_mai_n22_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, men_men_n17_, men_men_n18_, men_men_n19_, men_men_n20_, men_men_n21_, men_men_n22_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05;
  INV        o000(.A(x0), .Y(ori_ori_n17_));
  INV        o001(.A(x1), .Y(ori_ori_n18_));
  NO2        o002(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n19_));
  NO2        o003(.A(x6), .B(x5), .Y(ori_ori_n20_));
  OR2        o004(.A(x8), .B(x7), .Y(ori_ori_n21_));
  NOi21      o005(.An(ori_ori_n20_), .B(ori_ori_n21_), .Y(ori_ori_n22_));
  NAi21      o006(.An(ori_ori_n22_), .B(ori_ori_n19_), .Y(ori_ori_n23_));
  NA2        o007(.A(ori_ori_n18_), .B(ori_ori_n17_), .Y(ori_ori_n24_));
  INV        o008(.A(x5), .Y(ori_ori_n25_));
  NA2        o009(.A(x7), .B(x6), .Y(ori_ori_n26_));
  NA2        o010(.A(x8), .B(x3), .Y(ori_ori_n27_));
  NA2        o011(.A(x4), .B(x2), .Y(ori_ori_n28_));
  NO4        o012(.A(ori_ori_n28_), .B(ori_ori_n27_), .C(ori_ori_n26_), .D(ori_ori_n25_), .Y(ori_ori_n29_));
  NO2        o013(.A(ori_ori_n29_), .B(ori_ori_n24_), .Y(ori_ori_n30_));
  NO2        o014(.A(x4), .B(x3), .Y(ori_ori_n31_));
  INV        o015(.A(ori_ori_n31_), .Y(ori_ori_n32_));
  OA210      o016(.A0(ori_ori_n32_), .A1(x2), .B0(ori_ori_n19_), .Y(ori_ori_n33_));
  NOi31      o017(.An(ori_ori_n23_), .B(ori_ori_n33_), .C(ori_ori_n30_), .Y(ori00));
  NO2        o018(.A(x1), .B(x0), .Y(ori_ori_n35_));
  INV        o019(.A(x6), .Y(ori_ori_n36_));
  NO2        o020(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n37_));
  AN2        o021(.A(x8), .B(x7), .Y(ori_ori_n38_));
  NA3        o022(.A(ori_ori_n38_), .B(ori_ori_n37_), .C(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o023(.A(x4), .B(x3), .Y(ori_ori_n40_));
  AOI210     o024(.A0(ori_ori_n39_), .A1(ori_ori_n23_), .B0(ori_ori_n40_), .Y(ori_ori_n41_));
  NO2        o025(.A(x2), .B(x0), .Y(ori_ori_n42_));
  INV        o026(.A(x3), .Y(ori_ori_n43_));
  NO2        o027(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n44_));
  INV        o028(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO2        o029(.A(ori_ori_n37_), .B(x4), .Y(ori_ori_n46_));
  OAI210     o030(.A0(ori_ori_n46_), .A1(ori_ori_n45_), .B0(ori_ori_n42_), .Y(ori_ori_n47_));
  INV        o031(.A(x4), .Y(ori_ori_n48_));
  NO2        o032(.A(ori_ori_n48_), .B(ori_ori_n17_), .Y(ori_ori_n49_));
  NA2        o033(.A(ori_ori_n49_), .B(x2), .Y(ori_ori_n50_));
  OAI210     o034(.A0(ori_ori_n50_), .A1(ori_ori_n20_), .B0(ori_ori_n47_), .Y(ori_ori_n51_));
  NA2        o035(.A(ori_ori_n38_), .B(ori_ori_n37_), .Y(ori_ori_n52_));
  AOI220     o036(.A0(ori_ori_n52_), .A1(ori_ori_n35_), .B0(ori_ori_n22_), .B1(ori_ori_n19_), .Y(ori_ori_n53_));
  INV        o037(.A(x2), .Y(ori_ori_n54_));
  NO2        o038(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n55_));
  NA2        o039(.A(ori_ori_n43_), .B(ori_ori_n18_), .Y(ori_ori_n56_));
  NA2        o040(.A(ori_ori_n56_), .B(ori_ori_n55_), .Y(ori_ori_n57_));
  OAI210     o041(.A0(ori_ori_n53_), .A1(ori_ori_n32_), .B0(ori_ori_n57_), .Y(ori_ori_n58_));
  NO3        o042(.A(ori_ori_n58_), .B(ori_ori_n51_), .C(ori_ori_n41_), .Y(ori01));
  NA2        o043(.A(x8), .B(x7), .Y(ori_ori_n60_));
  NA2        o044(.A(ori_ori_n43_), .B(x1), .Y(ori_ori_n61_));
  INV        o045(.A(x9), .Y(ori_ori_n62_));
  NO2        o046(.A(ori_ori_n62_), .B(ori_ori_n36_), .Y(ori_ori_n63_));
  INV        o047(.A(ori_ori_n63_), .Y(ori_ori_n64_));
  NO3        o048(.A(ori_ori_n64_), .B(ori_ori_n61_), .C(ori_ori_n60_), .Y(ori_ori_n65_));
  NO2        o049(.A(x7), .B(x6), .Y(ori_ori_n66_));
  NO2        o050(.A(ori_ori_n61_), .B(x5), .Y(ori_ori_n67_));
  NO2        o051(.A(x8), .B(x2), .Y(ori_ori_n68_));
  INV        o052(.A(ori_ori_n68_), .Y(ori_ori_n69_));
  AN2        o053(.A(ori_ori_n67_), .B(ori_ori_n66_), .Y(ori_ori_n70_));
  OAI210     o054(.A0(ori_ori_n44_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n71_));
  OAI210     o055(.A0(ori_ori_n56_), .A1(ori_ori_n20_), .B0(ori_ori_n71_), .Y(ori_ori_n72_));
  NAi31      o056(.An(x1), .B(x9), .C(x5), .Y(ori_ori_n73_));
  NO2        o057(.A(ori_ori_n72_), .B(ori_ori_n70_), .Y(ori_ori_n74_));
  OAI210     o058(.A0(ori_ori_n74_), .A1(ori_ori_n65_), .B0(x4), .Y(ori_ori_n75_));
  NA2        o059(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n76_));
  OAI210     o060(.A0(ori_ori_n76_), .A1(ori_ori_n56_), .B0(x0), .Y(ori_ori_n77_));
  NA2        o061(.A(x5), .B(x3), .Y(ori_ori_n78_));
  NO2        o062(.A(x8), .B(x6), .Y(ori_ori_n79_));
  NO4        o063(.A(ori_ori_n79_), .B(ori_ori_n78_), .C(ori_ori_n66_), .D(ori_ori_n54_), .Y(ori_ori_n80_));
  NAi21      o064(.An(x4), .B(x3), .Y(ori_ori_n81_));
  INV        o065(.A(ori_ori_n81_), .Y(ori_ori_n82_));
  NO2        o066(.A(ori_ori_n82_), .B(ori_ori_n22_), .Y(ori_ori_n83_));
  NO2        o067(.A(x4), .B(x2), .Y(ori_ori_n84_));
  NO2        o068(.A(ori_ori_n84_), .B(x3), .Y(ori_ori_n85_));
  NO3        o069(.A(ori_ori_n85_), .B(ori_ori_n83_), .C(ori_ori_n18_), .Y(ori_ori_n86_));
  NO3        o070(.A(ori_ori_n86_), .B(ori_ori_n80_), .C(ori_ori_n77_), .Y(ori_ori_n87_));
  NA2        o071(.A(x3), .B(ori_ori_n18_), .Y(ori_ori_n88_));
  NO2        o072(.A(ori_ori_n88_), .B(ori_ori_n25_), .Y(ori_ori_n89_));
  INV        o073(.A(x8), .Y(ori_ori_n90_));
  NA2        o074(.A(x2), .B(x1), .Y(ori_ori_n91_));
  NO2        o075(.A(ori_ori_n91_), .B(ori_ori_n90_), .Y(ori_ori_n92_));
  NO2        o076(.A(ori_ori_n92_), .B(ori_ori_n89_), .Y(ori_ori_n93_));
  NO2        o077(.A(ori_ori_n93_), .B(ori_ori_n26_), .Y(ori_ori_n94_));
  AOI210     o078(.A0(ori_ori_n56_), .A1(ori_ori_n25_), .B0(ori_ori_n54_), .Y(ori_ori_n95_));
  OAI210     o079(.A0(ori_ori_n45_), .A1(ori_ori_n37_), .B0(ori_ori_n48_), .Y(ori_ori_n96_));
  NO3        o080(.A(ori_ori_n96_), .B(ori_ori_n95_), .C(ori_ori_n94_), .Y(ori_ori_n97_));
  NA2        o081(.A(x4), .B(ori_ori_n43_), .Y(ori_ori_n98_));
  NO2        o082(.A(ori_ori_n48_), .B(ori_ori_n54_), .Y(ori_ori_n99_));
  OAI210     o083(.A0(ori_ori_n99_), .A1(ori_ori_n43_), .B0(ori_ori_n18_), .Y(ori_ori_n100_));
  AOI210     o084(.A0(ori_ori_n98_), .A1(ori_ori_n52_), .B0(ori_ori_n100_), .Y(ori_ori_n101_));
  NO2        o085(.A(x3), .B(x2), .Y(ori_ori_n102_));
  NA3        o086(.A(ori_ori_n102_), .B(ori_ori_n26_), .C(ori_ori_n25_), .Y(ori_ori_n103_));
  AOI210     o087(.A0(x8), .A1(x6), .B0(ori_ori_n103_), .Y(ori_ori_n104_));
  NA2        o088(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n105_));
  OAI210     o089(.A0(ori_ori_n105_), .A1(ori_ori_n40_), .B0(ori_ori_n17_), .Y(ori_ori_n106_));
  NO4        o090(.A(ori_ori_n106_), .B(ori_ori_n104_), .C(ori_ori_n101_), .D(ori_ori_n97_), .Y(ori_ori_n107_));
  AO210      o091(.A0(ori_ori_n87_), .A1(ori_ori_n75_), .B0(ori_ori_n107_), .Y(ori02));
  NO2        o092(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n109_));
  NO2        o093(.A(x8), .B(ori_ori_n18_), .Y(ori_ori_n110_));
  NA2        o094(.A(ori_ori_n54_), .B(ori_ori_n17_), .Y(ori_ori_n111_));
  NA2        o095(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n112_));
  INV        o096(.A(ori_ori_n112_), .Y(ori_ori_n113_));
  AOI220     o097(.A0(ori_ori_n113_), .A1(ori_ori_n110_), .B0(ori_ori_n109_), .B1(x4), .Y(ori_ori_n114_));
  NO3        o098(.A(ori_ori_n114_), .B(x7), .C(x5), .Y(ori_ori_n115_));
  NA2        o099(.A(x9), .B(x2), .Y(ori_ori_n116_));
  OR2        o100(.A(x8), .B(x0), .Y(ori_ori_n117_));
  INV        o101(.A(ori_ori_n117_), .Y(ori_ori_n118_));
  NAi21      o102(.An(x2), .B(x8), .Y(ori_ori_n119_));
  INV        o103(.A(ori_ori_n119_), .Y(ori_ori_n120_));
  NO2        o104(.A(x4), .B(x1), .Y(ori_ori_n121_));
  NA3        o105(.A(ori_ori_n121_), .B(x2), .C(ori_ori_n60_), .Y(ori_ori_n122_));
  NOi21      o106(.An(x0), .B(x1), .Y(ori_ori_n123_));
  NO3        o107(.A(x9), .B(x8), .C(x7), .Y(ori_ori_n124_));
  NOi21      o108(.An(x0), .B(x4), .Y(ori_ori_n125_));
  NAi21      o109(.An(x8), .B(x7), .Y(ori_ori_n126_));
  NO2        o110(.A(ori_ori_n126_), .B(ori_ori_n62_), .Y(ori_ori_n127_));
  AOI220     o111(.A0(ori_ori_n127_), .A1(ori_ori_n125_), .B0(ori_ori_n124_), .B1(ori_ori_n123_), .Y(ori_ori_n128_));
  AOI210     o112(.A0(ori_ori_n128_), .A1(ori_ori_n122_), .B0(ori_ori_n78_), .Y(ori_ori_n129_));
  NO2        o113(.A(x5), .B(ori_ori_n48_), .Y(ori_ori_n130_));
  NA2        o114(.A(x2), .B(ori_ori_n18_), .Y(ori_ori_n131_));
  AOI210     o115(.A0(ori_ori_n131_), .A1(ori_ori_n105_), .B0(ori_ori_n112_), .Y(ori_ori_n132_));
  OAI210     o116(.A0(ori_ori_n132_), .A1(ori_ori_n35_), .B0(ori_ori_n130_), .Y(ori_ori_n133_));
  NAi21      o117(.An(x0), .B(x4), .Y(ori_ori_n134_));
  NO2        o118(.A(ori_ori_n134_), .B(x1), .Y(ori_ori_n135_));
  NO2        o119(.A(x7), .B(x0), .Y(ori_ori_n136_));
  NO2        o120(.A(ori_ori_n84_), .B(ori_ori_n99_), .Y(ori_ori_n137_));
  NO2        o121(.A(ori_ori_n137_), .B(x3), .Y(ori_ori_n138_));
  OAI210     o122(.A0(ori_ori_n136_), .A1(ori_ori_n135_), .B0(ori_ori_n138_), .Y(ori_ori_n139_));
  NO2        o123(.A(ori_ori_n21_), .B(ori_ori_n43_), .Y(ori_ori_n140_));
  NA2        o124(.A(x5), .B(x0), .Y(ori_ori_n141_));
  NO2        o125(.A(ori_ori_n48_), .B(x2), .Y(ori_ori_n142_));
  NA3        o126(.A(ori_ori_n142_), .B(ori_ori_n141_), .C(ori_ori_n140_), .Y(ori_ori_n143_));
  NA4        o127(.A(ori_ori_n143_), .B(ori_ori_n139_), .C(ori_ori_n133_), .D(ori_ori_n36_), .Y(ori_ori_n144_));
  NO3        o128(.A(ori_ori_n144_), .B(ori_ori_n129_), .C(ori_ori_n115_), .Y(ori_ori_n145_));
  NO3        o129(.A(ori_ori_n78_), .B(ori_ori_n76_), .C(ori_ori_n24_), .Y(ori_ori_n146_));
  NO2        o130(.A(ori_ori_n28_), .B(ori_ori_n25_), .Y(ori_ori_n147_));
  AOI220     o131(.A0(ori_ori_n123_), .A1(ori_ori_n147_), .B0(ori_ori_n67_), .B1(ori_ori_n17_), .Y(ori_ori_n148_));
  NO3        o132(.A(ori_ori_n148_), .B(ori_ori_n60_), .C(ori_ori_n62_), .Y(ori_ori_n149_));
  NA2        o133(.A(x7), .B(x3), .Y(ori_ori_n150_));
  NO2        o134(.A(ori_ori_n98_), .B(x5), .Y(ori_ori_n151_));
  NO2        o135(.A(x9), .B(x7), .Y(ori_ori_n152_));
  NOi21      o136(.An(x8), .B(x0), .Y(ori_ori_n153_));
  OA210      o137(.A0(ori_ori_n152_), .A1(x1), .B0(ori_ori_n153_), .Y(ori_ori_n154_));
  NO2        o138(.A(ori_ori_n43_), .B(x2), .Y(ori_ori_n155_));
  INV        o139(.A(x7), .Y(ori_ori_n156_));
  NA2        o140(.A(ori_ori_n156_), .B(ori_ori_n18_), .Y(ori_ori_n157_));
  AOI220     o141(.A0(ori_ori_n157_), .A1(ori_ori_n155_), .B0(ori_ori_n109_), .B1(ori_ori_n38_), .Y(ori_ori_n158_));
  NO2        o142(.A(ori_ori_n25_), .B(x4), .Y(ori_ori_n159_));
  NO2        o143(.A(ori_ori_n159_), .B(ori_ori_n125_), .Y(ori_ori_n160_));
  NO2        o144(.A(ori_ori_n160_), .B(ori_ori_n158_), .Y(ori_ori_n161_));
  AOI210     o145(.A0(ori_ori_n154_), .A1(ori_ori_n151_), .B0(ori_ori_n161_), .Y(ori_ori_n162_));
  OAI210     o146(.A0(ori_ori_n150_), .A1(ori_ori_n50_), .B0(ori_ori_n162_), .Y(ori_ori_n163_));
  NA2        o147(.A(x5), .B(x1), .Y(ori_ori_n164_));
  INV        o148(.A(ori_ori_n164_), .Y(ori_ori_n165_));
  AOI210     o149(.A0(ori_ori_n165_), .A1(ori_ori_n125_), .B0(ori_ori_n36_), .Y(ori_ori_n166_));
  NO2        o150(.A(ori_ori_n62_), .B(ori_ori_n90_), .Y(ori_ori_n167_));
  NAi21      o151(.An(x2), .B(x7), .Y(ori_ori_n168_));
  NO3        o152(.A(ori_ori_n168_), .B(ori_ori_n167_), .C(ori_ori_n48_), .Y(ori_ori_n169_));
  NA2        o153(.A(ori_ori_n169_), .B(ori_ori_n67_), .Y(ori_ori_n170_));
  NAi31      o154(.An(ori_ori_n78_), .B(ori_ori_n38_), .C(ori_ori_n35_), .Y(ori_ori_n171_));
  NA3        o155(.A(ori_ori_n171_), .B(ori_ori_n170_), .C(ori_ori_n166_), .Y(ori_ori_n172_));
  NO4        o156(.A(ori_ori_n172_), .B(ori_ori_n163_), .C(ori_ori_n149_), .D(ori_ori_n146_), .Y(ori_ori_n173_));
  NO2        o157(.A(ori_ori_n173_), .B(ori_ori_n145_), .Y(ori_ori_n174_));
  NO2        o158(.A(ori_ori_n141_), .B(ori_ori_n137_), .Y(ori_ori_n175_));
  NA2        o159(.A(ori_ori_n25_), .B(ori_ori_n18_), .Y(ori_ori_n176_));
  NA2        o160(.A(ori_ori_n25_), .B(ori_ori_n17_), .Y(ori_ori_n177_));
  NA3        o161(.A(ori_ori_n177_), .B(ori_ori_n176_), .C(ori_ori_n24_), .Y(ori_ori_n178_));
  AN2        o162(.A(ori_ori_n178_), .B(ori_ori_n142_), .Y(ori_ori_n179_));
  NA2        o163(.A(x8), .B(x0), .Y(ori_ori_n180_));
  NO2        o164(.A(ori_ori_n156_), .B(ori_ori_n25_), .Y(ori_ori_n181_));
  NO2        o165(.A(ori_ori_n123_), .B(x4), .Y(ori_ori_n182_));
  NA2        o166(.A(ori_ori_n182_), .B(ori_ori_n181_), .Y(ori_ori_n183_));
  AOI210     o167(.A0(ori_ori_n180_), .A1(ori_ori_n131_), .B0(ori_ori_n183_), .Y(ori_ori_n184_));
  NA2        o168(.A(x2), .B(x0), .Y(ori_ori_n185_));
  NA2        o169(.A(x4), .B(x1), .Y(ori_ori_n186_));
  NAi21      o170(.An(ori_ori_n121_), .B(ori_ori_n186_), .Y(ori_ori_n187_));
  NOi31      o171(.An(ori_ori_n187_), .B(ori_ori_n159_), .C(ori_ori_n185_), .Y(ori_ori_n188_));
  NO4        o172(.A(ori_ori_n188_), .B(ori_ori_n184_), .C(ori_ori_n179_), .D(ori_ori_n175_), .Y(ori_ori_n189_));
  NO2        o173(.A(ori_ori_n189_), .B(ori_ori_n43_), .Y(ori_ori_n190_));
  NO2        o174(.A(ori_ori_n178_), .B(ori_ori_n76_), .Y(ori_ori_n191_));
  INV        o175(.A(ori_ori_n130_), .Y(ori_ori_n192_));
  NO2        o176(.A(ori_ori_n105_), .B(ori_ori_n17_), .Y(ori_ori_n193_));
  AOI210     o177(.A0(ori_ori_n35_), .A1(ori_ori_n90_), .B0(ori_ori_n193_), .Y(ori_ori_n194_));
  NO3        o178(.A(ori_ori_n194_), .B(ori_ori_n192_), .C(x7), .Y(ori_ori_n195_));
  NA3        o179(.A(ori_ori_n187_), .B(ori_ori_n192_), .C(ori_ori_n42_), .Y(ori_ori_n196_));
  OAI210     o180(.A0(ori_ori_n177_), .A1(ori_ori_n137_), .B0(ori_ori_n196_), .Y(ori_ori_n197_));
  NO3        o181(.A(ori_ori_n197_), .B(ori_ori_n195_), .C(ori_ori_n191_), .Y(ori_ori_n198_));
  NO2        o182(.A(ori_ori_n198_), .B(x3), .Y(ori_ori_n199_));
  NO3        o183(.A(ori_ori_n199_), .B(ori_ori_n190_), .C(ori_ori_n174_), .Y(ori03));
  NO2        o184(.A(ori_ori_n48_), .B(x3), .Y(ori_ori_n201_));
  NO2        o185(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n202_));
  INV        o186(.A(ori_ori_n202_), .Y(ori_ori_n203_));
  NO2        o187(.A(ori_ori_n54_), .B(x1), .Y(ori_ori_n204_));
  OAI210     o188(.A0(ori_ori_n204_), .A1(ori_ori_n25_), .B0(ori_ori_n63_), .Y(ori_ori_n205_));
  OAI220     o189(.A0(ori_ori_n205_), .A1(ori_ori_n17_), .B0(ori_ori_n203_), .B1(ori_ori_n105_), .Y(ori_ori_n206_));
  NA2        o190(.A(ori_ori_n206_), .B(ori_ori_n201_), .Y(ori_ori_n207_));
  NO2        o191(.A(ori_ori_n78_), .B(x6), .Y(ori_ori_n208_));
  NA2        o192(.A(x6), .B(ori_ori_n25_), .Y(ori_ori_n209_));
  NO2        o193(.A(ori_ori_n209_), .B(x4), .Y(ori_ori_n210_));
  NO2        o194(.A(ori_ori_n18_), .B(x0), .Y(ori_ori_n211_));
  AN2        o195(.A(ori_ori_n208_), .B(ori_ori_n55_), .Y(ori_ori_n212_));
  NA2        o196(.A(ori_ori_n212_), .B(ori_ori_n62_), .Y(ori_ori_n213_));
  NA2        o197(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n214_));
  NO2        o198(.A(ori_ori_n214_), .B(ori_ori_n209_), .Y(ori_ori_n215_));
  NA2        o199(.A(x9), .B(ori_ori_n54_), .Y(ori_ori_n216_));
  NA2        o200(.A(ori_ori_n216_), .B(x4), .Y(ori_ori_n217_));
  NA2        o201(.A(ori_ori_n209_), .B(ori_ori_n81_), .Y(ori_ori_n218_));
  AOI210     o202(.A0(ori_ori_n25_), .A1(x3), .B0(ori_ori_n185_), .Y(ori_ori_n219_));
  AOI220     o203(.A0(ori_ori_n219_), .A1(ori_ori_n218_), .B0(ori_ori_n217_), .B1(ori_ori_n215_), .Y(ori_ori_n220_));
  NO3        o204(.A(x6), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n221_));
  NO2        o205(.A(x5), .B(x1), .Y(ori_ori_n222_));
  NO2        o206(.A(ori_ori_n214_), .B(ori_ori_n176_), .Y(ori_ori_n223_));
  NO3        o207(.A(x3), .B(x2), .C(x1), .Y(ori_ori_n224_));
  NO2        o208(.A(ori_ori_n224_), .B(ori_ori_n223_), .Y(ori_ori_n225_));
  INV        o209(.A(ori_ori_n225_), .Y(ori_ori_n226_));
  AOI220     o210(.A0(ori_ori_n226_), .A1(ori_ori_n48_), .B0(ori_ori_n221_), .B1(ori_ori_n130_), .Y(ori_ori_n227_));
  NA4        o211(.A(ori_ori_n227_), .B(ori_ori_n220_), .C(ori_ori_n213_), .D(ori_ori_n207_), .Y(ori_ori_n228_));
  NO2        o212(.A(ori_ori_n48_), .B(ori_ori_n43_), .Y(ori_ori_n229_));
  NA2        o213(.A(ori_ori_n229_), .B(ori_ori_n19_), .Y(ori_ori_n230_));
  NO2        o214(.A(x3), .B(ori_ori_n17_), .Y(ori_ori_n231_));
  NO2        o215(.A(ori_ori_n231_), .B(x6), .Y(ori_ori_n232_));
  NOi21      o216(.An(ori_ori_n84_), .B(ori_ori_n232_), .Y(ori_ori_n233_));
  NA2        o217(.A(ori_ori_n62_), .B(ori_ori_n90_), .Y(ori_ori_n234_));
  NA3        o218(.A(ori_ori_n234_), .B(ori_ori_n231_), .C(x6), .Y(ori_ori_n235_));
  AOI210     o219(.A0(ori_ori_n235_), .A1(ori_ori_n233_), .B0(ori_ori_n156_), .Y(ori_ori_n236_));
  AO210      o220(.A0(ori_ori_n236_), .A1(ori_ori_n230_), .B0(ori_ori_n181_), .Y(ori_ori_n237_));
  NA2        o221(.A(ori_ori_n43_), .B(ori_ori_n54_), .Y(ori_ori_n238_));
  OAI210     o222(.A0(ori_ori_n238_), .A1(ori_ori_n25_), .B0(ori_ori_n177_), .Y(ori_ori_n239_));
  NO3        o223(.A(ori_ori_n186_), .B(ori_ori_n62_), .C(x6), .Y(ori_ori_n240_));
  AOI220     o224(.A0(ori_ori_n240_), .A1(ori_ori_n239_), .B0(ori_ori_n142_), .B1(ori_ori_n89_), .Y(ori_ori_n241_));
  NA2        o225(.A(x6), .B(ori_ori_n48_), .Y(ori_ori_n242_));
  OAI210     o226(.A0(ori_ori_n118_), .A1(ori_ori_n79_), .B0(x4), .Y(ori_ori_n243_));
  AOI210     o227(.A0(ori_ori_n243_), .A1(ori_ori_n242_), .B0(ori_ori_n78_), .Y(ori_ori_n244_));
  NO2        o228(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n245_));
  NO2        o229(.A(ori_ori_n164_), .B(ori_ori_n43_), .Y(ori_ori_n246_));
  OAI210     o230(.A0(ori_ori_n246_), .A1(ori_ori_n223_), .B0(ori_ori_n245_), .Y(ori_ori_n247_));
  NA2        o231(.A(ori_ori_n202_), .B(ori_ori_n135_), .Y(ori_ori_n248_));
  NA3        o232(.A(ori_ori_n214_), .B(ori_ori_n130_), .C(x6), .Y(ori_ori_n249_));
  OAI210     o233(.A0(ori_ori_n90_), .A1(ori_ori_n36_), .B0(ori_ori_n67_), .Y(ori_ori_n250_));
  NA4        o234(.A(ori_ori_n250_), .B(ori_ori_n249_), .C(ori_ori_n248_), .D(ori_ori_n247_), .Y(ori_ori_n251_));
  OAI210     o235(.A0(ori_ori_n251_), .A1(ori_ori_n244_), .B0(x2), .Y(ori_ori_n252_));
  NA3        o236(.A(ori_ori_n252_), .B(ori_ori_n241_), .C(ori_ori_n237_), .Y(ori_ori_n253_));
  AOI210     o237(.A0(ori_ori_n228_), .A1(x8), .B0(ori_ori_n253_), .Y(ori_ori_n254_));
  NO2        o238(.A(ori_ori_n90_), .B(x3), .Y(ori_ori_n255_));
  NA2        o239(.A(ori_ori_n255_), .B(ori_ori_n210_), .Y(ori_ori_n256_));
  NO3        o240(.A(ori_ori_n88_), .B(ori_ori_n79_), .C(ori_ori_n25_), .Y(ori_ori_n257_));
  AOI210     o241(.A0(ori_ori_n232_), .A1(ori_ori_n159_), .B0(ori_ori_n257_), .Y(ori_ori_n258_));
  AOI210     o242(.A0(ori_ori_n258_), .A1(ori_ori_n256_), .B0(x2), .Y(ori_ori_n259_));
  NO2        o243(.A(x4), .B(ori_ori_n54_), .Y(ori_ori_n260_));
  AOI220     o244(.A0(ori_ori_n210_), .A1(ori_ori_n193_), .B0(ori_ori_n260_), .B1(ori_ori_n67_), .Y(ori_ori_n261_));
  NA2        o245(.A(ori_ori_n62_), .B(x6), .Y(ori_ori_n262_));
  NA2        o246(.A(ori_ori_n43_), .B(ori_ori_n17_), .Y(ori_ori_n263_));
  NO2        o247(.A(ori_ori_n263_), .B(ori_ori_n25_), .Y(ori_ori_n264_));
  NA2        o248(.A(ori_ori_n264_), .B(ori_ori_n121_), .Y(ori_ori_n265_));
  NA2        o249(.A(ori_ori_n214_), .B(x6), .Y(ori_ori_n266_));
  NO2        o250(.A(ori_ori_n214_), .B(x6), .Y(ori_ori_n267_));
  NAi21      o251(.An(ori_ori_n167_), .B(ori_ori_n267_), .Y(ori_ori_n268_));
  NA3        o252(.A(ori_ori_n268_), .B(ori_ori_n266_), .C(ori_ori_n147_), .Y(ori_ori_n269_));
  NA4        o253(.A(ori_ori_n269_), .B(ori_ori_n265_), .C(ori_ori_n261_), .D(ori_ori_n156_), .Y(ori_ori_n270_));
  NA2        o254(.A(ori_ori_n202_), .B(ori_ori_n231_), .Y(ori_ori_n271_));
  NO2        o255(.A(ori_ori_n141_), .B(ori_ori_n18_), .Y(ori_ori_n272_));
  NAi21      o256(.An(x1), .B(x4), .Y(ori_ori_n273_));
  AOI210     o257(.A0(x3), .A1(x2), .B0(ori_ori_n48_), .Y(ori_ori_n274_));
  OAI210     o258(.A0(ori_ori_n141_), .A1(x3), .B0(ori_ori_n274_), .Y(ori_ori_n275_));
  NA2        o259(.A(ori_ori_n275_), .B(ori_ori_n273_), .Y(ori_ori_n276_));
  NA2        o260(.A(ori_ori_n276_), .B(ori_ori_n271_), .Y(ori_ori_n277_));
  NA2        o261(.A(ori_ori_n62_), .B(x2), .Y(ori_ori_n278_));
  NO2        o262(.A(ori_ori_n278_), .B(ori_ori_n271_), .Y(ori_ori_n279_));
  NA2        o263(.A(x6), .B(x2), .Y(ori_ori_n280_));
  NO2        o264(.A(ori_ori_n182_), .B(ori_ori_n46_), .Y(ori_ori_n281_));
  OAI210     o265(.A0(ori_ori_n281_), .A1(ori_ori_n279_), .B0(ori_ori_n277_), .Y(ori_ori_n282_));
  NA2        o266(.A(x9), .B(ori_ori_n43_), .Y(ori_ori_n283_));
  NO2        o267(.A(ori_ori_n283_), .B(ori_ori_n209_), .Y(ori_ori_n284_));
  OR3        o268(.A(ori_ori_n284_), .B(ori_ori_n208_), .C(ori_ori_n151_), .Y(ori_ori_n285_));
  NA2        o269(.A(x4), .B(x0), .Y(ori_ori_n286_));
  NO3        o270(.A(ori_ori_n73_), .B(ori_ori_n286_), .C(x6), .Y(ori_ori_n287_));
  AOI210     o271(.A0(ori_ori_n285_), .A1(ori_ori_n42_), .B0(ori_ori_n287_), .Y(ori_ori_n288_));
  AOI210     o272(.A0(ori_ori_n288_), .A1(ori_ori_n282_), .B0(x8), .Y(ori_ori_n289_));
  INV        o273(.A(ori_ori_n262_), .Y(ori_ori_n290_));
  OAI210     o274(.A0(ori_ori_n272_), .A1(ori_ori_n222_), .B0(ori_ori_n290_), .Y(ori_ori_n291_));
  INV        o275(.A(ori_ori_n180_), .Y(ori_ori_n292_));
  OAI210     o276(.A0(ori_ori_n292_), .A1(x4), .B0(ori_ori_n20_), .Y(ori_ori_n293_));
  AOI210     o277(.A0(ori_ori_n293_), .A1(ori_ori_n291_), .B0(ori_ori_n238_), .Y(ori_ori_n294_));
  NO4        o278(.A(ori_ori_n294_), .B(ori_ori_n289_), .C(ori_ori_n270_), .D(ori_ori_n259_), .Y(ori_ori_n295_));
  NO2        o279(.A(ori_ori_n167_), .B(x1), .Y(ori_ori_n296_));
  NO3        o280(.A(ori_ori_n296_), .B(x3), .C(ori_ori_n36_), .Y(ori_ori_n297_));
  OAI210     o281(.A0(ori_ori_n297_), .A1(ori_ori_n267_), .B0(x2), .Y(ori_ori_n298_));
  OAI210     o282(.A0(ori_ori_n292_), .A1(x6), .B0(ori_ori_n44_), .Y(ori_ori_n299_));
  AOI210     o283(.A0(ori_ori_n299_), .A1(ori_ori_n298_), .B0(ori_ori_n192_), .Y(ori_ori_n300_));
  NOi21      o284(.An(ori_ori_n280_), .B(ori_ori_n17_), .Y(ori_ori_n301_));
  NA3        o285(.A(ori_ori_n301_), .B(ori_ori_n222_), .C(ori_ori_n40_), .Y(ori_ori_n302_));
  AOI210     o286(.A0(ori_ori_n36_), .A1(ori_ori_n54_), .B0(x0), .Y(ori_ori_n303_));
  NA3        o287(.A(ori_ori_n303_), .B(ori_ori_n165_), .C(ori_ori_n32_), .Y(ori_ori_n304_));
  NA2        o288(.A(x3), .B(x2), .Y(ori_ori_n305_));
  AOI220     o289(.A0(ori_ori_n305_), .A1(ori_ori_n238_), .B0(ori_ori_n304_), .B1(ori_ori_n302_), .Y(ori_ori_n306_));
  NAi21      o290(.An(x4), .B(x0), .Y(ori_ori_n307_));
  NO3        o291(.A(ori_ori_n307_), .B(ori_ori_n44_), .C(x2), .Y(ori_ori_n308_));
  OAI210     o292(.A0(x6), .A1(ori_ori_n18_), .B0(ori_ori_n308_), .Y(ori_ori_n309_));
  OAI220     o293(.A0(ori_ori_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(ori_ori_n310_));
  NO2        o294(.A(x9), .B(x8), .Y(ori_ori_n311_));
  NA3        o295(.A(ori_ori_n311_), .B(ori_ori_n36_), .C(ori_ori_n54_), .Y(ori_ori_n312_));
  OAI210     o296(.A0(ori_ori_n303_), .A1(ori_ori_n301_), .B0(ori_ori_n312_), .Y(ori_ori_n313_));
  AOI220     o297(.A0(ori_ori_n313_), .A1(ori_ori_n82_), .B0(ori_ori_n310_), .B1(ori_ori_n31_), .Y(ori_ori_n314_));
  AOI210     o298(.A0(ori_ori_n314_), .A1(ori_ori_n309_), .B0(ori_ori_n25_), .Y(ori_ori_n315_));
  NA3        o299(.A(ori_ori_n36_), .B(x1), .C(ori_ori_n17_), .Y(ori_ori_n316_));
  OAI210     o300(.A0(ori_ori_n303_), .A1(ori_ori_n301_), .B0(ori_ori_n316_), .Y(ori_ori_n317_));
  INV        o301(.A(ori_ori_n223_), .Y(ori_ori_n318_));
  NA2        o302(.A(ori_ori_n36_), .B(ori_ori_n43_), .Y(ori_ori_n319_));
  OR2        o303(.A(ori_ori_n319_), .B(ori_ori_n286_), .Y(ori_ori_n320_));
  OAI220     o304(.A0(ori_ori_n320_), .A1(ori_ori_n164_), .B0(ori_ori_n242_), .B1(ori_ori_n318_), .Y(ori_ori_n321_));
  AO210      o305(.A0(ori_ori_n317_), .A1(ori_ori_n151_), .B0(ori_ori_n321_), .Y(ori_ori_n322_));
  NO4        o306(.A(ori_ori_n322_), .B(ori_ori_n315_), .C(ori_ori_n306_), .D(ori_ori_n300_), .Y(ori_ori_n323_));
  OAI210     o307(.A0(ori_ori_n295_), .A1(ori_ori_n254_), .B0(ori_ori_n323_), .Y(ori04));
  NO2        o308(.A(x2), .B(x1), .Y(ori_ori_n325_));
  OAI210     o309(.A0(ori_ori_n263_), .A1(ori_ori_n325_), .B0(ori_ori_n36_), .Y(ori_ori_n326_));
  NO2        o310(.A(ori_ori_n325_), .B(ori_ori_n307_), .Y(ori_ori_n327_));
  AOI210     o311(.A0(ori_ori_n62_), .A1(x4), .B0(ori_ori_n111_), .Y(ori_ori_n328_));
  OAI210     o312(.A0(ori_ori_n328_), .A1(ori_ori_n327_), .B0(ori_ori_n255_), .Y(ori_ori_n329_));
  NO2        o313(.A(ori_ori_n278_), .B(ori_ori_n88_), .Y(ori_ori_n330_));
  NO2        o314(.A(ori_ori_n330_), .B(ori_ori_n36_), .Y(ori_ori_n331_));
  NO2        o315(.A(ori_ori_n305_), .B(ori_ori_n211_), .Y(ori_ori_n332_));
  NA2        o316(.A(x9), .B(x0), .Y(ori_ori_n333_));
  AOI210     o317(.A0(ori_ori_n88_), .A1(ori_ori_n76_), .B0(ori_ori_n333_), .Y(ori_ori_n334_));
  OAI210     o318(.A0(ori_ori_n334_), .A1(ori_ori_n332_), .B0(ori_ori_n90_), .Y(ori_ori_n335_));
  NA3        o319(.A(ori_ori_n335_), .B(ori_ori_n331_), .C(ori_ori_n329_), .Y(ori_ori_n336_));
  NA2        o320(.A(ori_ori_n336_), .B(ori_ori_n326_), .Y(ori_ori_n337_));
  NO2        o321(.A(ori_ori_n216_), .B(ori_ori_n112_), .Y(ori_ori_n338_));
  NO3        o322(.A(ori_ori_n262_), .B(ori_ori_n119_), .C(ori_ori_n18_), .Y(ori_ori_n339_));
  NO2        o323(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  OAI210     o324(.A0(ori_ori_n117_), .A1(ori_ori_n105_), .B0(ori_ori_n180_), .Y(ori_ori_n341_));
  NA3        o325(.A(ori_ori_n341_), .B(x6), .C(x3), .Y(ori_ori_n342_));
  NOi21      o326(.An(ori_ori_n153_), .B(ori_ori_n131_), .Y(ori_ori_n343_));
  AOI210     o327(.A0(x8), .A1(x0), .B0(x1), .Y(ori_ori_n344_));
  OAI220     o328(.A0(ori_ori_n344_), .A1(ori_ori_n319_), .B0(ori_ori_n278_), .B1(ori_ori_n316_), .Y(ori_ori_n345_));
  AOI210     o329(.A0(ori_ori_n343_), .A1(ori_ori_n63_), .B0(ori_ori_n345_), .Y(ori_ori_n346_));
  NA2        o330(.A(x2), .B(ori_ori_n17_), .Y(ori_ori_n347_));
  OAI210     o331(.A0(ori_ori_n105_), .A1(ori_ori_n17_), .B0(ori_ori_n347_), .Y(ori_ori_n348_));
  NA2        o332(.A(ori_ori_n348_), .B(ori_ori_n79_), .Y(ori_ori_n349_));
  NA4        o333(.A(ori_ori_n349_), .B(ori_ori_n346_), .C(ori_ori_n342_), .D(ori_ori_n340_), .Y(ori_ori_n350_));
  OAI210     o334(.A0(ori_ori_n110_), .A1(x3), .B0(ori_ori_n308_), .Y(ori_ori_n351_));
  NA2        o335(.A(ori_ori_n221_), .B(ori_ori_n84_), .Y(ori_ori_n352_));
  NA3        o336(.A(ori_ori_n352_), .B(ori_ori_n351_), .C(ori_ori_n156_), .Y(ori_ori_n353_));
  AOI210     o337(.A0(ori_ori_n350_), .A1(x4), .B0(ori_ori_n353_), .Y(ori_ori_n354_));
  NA3        o338(.A(ori_ori_n327_), .B(ori_ori_n216_), .C(ori_ori_n90_), .Y(ori_ori_n355_));
  NOi21      o339(.An(x4), .B(x0), .Y(ori_ori_n356_));
  XO2        o340(.A(x4), .B(x0), .Y(ori_ori_n357_));
  OAI210     o341(.A0(ori_ori_n357_), .A1(ori_ori_n116_), .B0(ori_ori_n273_), .Y(ori_ori_n358_));
  AOI220     o342(.A0(ori_ori_n358_), .A1(x8), .B0(ori_ori_n356_), .B1(ori_ori_n91_), .Y(ori_ori_n359_));
  AOI210     o343(.A0(ori_ori_n359_), .A1(ori_ori_n355_), .B0(x3), .Y(ori_ori_n360_));
  INV        o344(.A(ori_ori_n91_), .Y(ori_ori_n361_));
  NO2        o345(.A(ori_ori_n90_), .B(x4), .Y(ori_ori_n362_));
  AOI220     o346(.A0(ori_ori_n362_), .A1(ori_ori_n44_), .B0(ori_ori_n125_), .B1(ori_ori_n361_), .Y(ori_ori_n363_));
  NO3        o347(.A(ori_ori_n357_), .B(ori_ori_n167_), .C(x2), .Y(ori_ori_n364_));
  NO3        o348(.A(ori_ori_n234_), .B(ori_ori_n28_), .C(ori_ori_n24_), .Y(ori_ori_n365_));
  NO2        o349(.A(ori_ori_n365_), .B(ori_ori_n364_), .Y(ori_ori_n366_));
  NA4        o350(.A(ori_ori_n366_), .B(ori_ori_n363_), .C(ori_ori_n230_), .D(x6), .Y(ori_ori_n367_));
  OAI220     o351(.A0(ori_ori_n307_), .A1(ori_ori_n88_), .B0(ori_ori_n185_), .B1(ori_ori_n90_), .Y(ori_ori_n368_));
  NO2        o352(.A(ori_ori_n43_), .B(x0), .Y(ori_ori_n369_));
  OR2        o353(.A(ori_ori_n362_), .B(ori_ori_n369_), .Y(ori_ori_n370_));
  NO2        o354(.A(ori_ori_n153_), .B(ori_ori_n105_), .Y(ori_ori_n371_));
  AOI220     o355(.A0(ori_ori_n371_), .A1(ori_ori_n370_), .B0(ori_ori_n368_), .B1(ori_ori_n61_), .Y(ori_ori_n372_));
  NO2        o356(.A(ori_ori_n153_), .B(ori_ori_n81_), .Y(ori_ori_n373_));
  NO2        o357(.A(ori_ori_n35_), .B(x2), .Y(ori_ori_n374_));
  NOi21      o358(.An(ori_ori_n121_), .B(ori_ori_n27_), .Y(ori_ori_n375_));
  AOI210     o359(.A0(ori_ori_n374_), .A1(ori_ori_n373_), .B0(ori_ori_n375_), .Y(ori_ori_n376_));
  OAI210     o360(.A0(ori_ori_n372_), .A1(ori_ori_n62_), .B0(ori_ori_n376_), .Y(ori_ori_n377_));
  OAI220     o361(.A0(ori_ori_n377_), .A1(x6), .B0(ori_ori_n367_), .B1(ori_ori_n360_), .Y(ori_ori_n378_));
  OAI210     o362(.A0(ori_ori_n63_), .A1(ori_ori_n48_), .B0(ori_ori_n42_), .Y(ori_ori_n379_));
  OAI210     o363(.A0(ori_ori_n379_), .A1(ori_ori_n90_), .B0(ori_ori_n320_), .Y(ori_ori_n380_));
  AOI210     o364(.A0(ori_ori_n380_), .A1(ori_ori_n18_), .B0(ori_ori_n156_), .Y(ori_ori_n381_));
  AO220      o365(.A0(ori_ori_n381_), .A1(ori_ori_n378_), .B0(ori_ori_n354_), .B1(ori_ori_n337_), .Y(ori_ori_n382_));
  NA2        o366(.A(ori_ori_n374_), .B(x6), .Y(ori_ori_n383_));
  AOI210     o367(.A0(x6), .A1(x1), .B0(ori_ori_n155_), .Y(ori_ori_n384_));
  NA2        o368(.A(ori_ori_n362_), .B(x0), .Y(ori_ori_n385_));
  NA2        o369(.A(ori_ori_n84_), .B(x6), .Y(ori_ori_n386_));
  OAI210     o370(.A0(ori_ori_n385_), .A1(ori_ori_n384_), .B0(ori_ori_n386_), .Y(ori_ori_n387_));
  AOI220     o371(.A0(ori_ori_n387_), .A1(ori_ori_n383_), .B0(ori_ori_n224_), .B1(ori_ori_n49_), .Y(ori_ori_n388_));
  NA2        o372(.A(ori_ori_n388_), .B(ori_ori_n382_), .Y(ori_ori_n389_));
  AOI210     o373(.A0(ori_ori_n204_), .A1(x8), .B0(ori_ori_n110_), .Y(ori_ori_n390_));
  NA2        o374(.A(ori_ori_n390_), .B(ori_ori_n347_), .Y(ori_ori_n391_));
  NA3        o375(.A(ori_ori_n391_), .B(ori_ori_n201_), .C(ori_ori_n156_), .Y(ori_ori_n392_));
  OAI210     o376(.A0(ori_ori_n28_), .A1(x1), .B0(ori_ori_n238_), .Y(ori_ori_n393_));
  AO220      o377(.A0(ori_ori_n393_), .A1(ori_ori_n152_), .B0(ori_ori_n109_), .B1(x4), .Y(ori_ori_n394_));
  NA3        o378(.A(x7), .B(x3), .C(x0), .Y(ori_ori_n395_));
  NA2        o379(.A(ori_ori_n229_), .B(x0), .Y(ori_ori_n396_));
  OAI220     o380(.A0(ori_ori_n396_), .A1(ori_ori_n216_), .B0(ori_ori_n395_), .B1(ori_ori_n361_), .Y(ori_ori_n397_));
  AOI210     o381(.A0(ori_ori_n394_), .A1(ori_ori_n118_), .B0(ori_ori_n397_), .Y(ori_ori_n398_));
  AOI210     o382(.A0(ori_ori_n398_), .A1(ori_ori_n392_), .B0(ori_ori_n25_), .Y(ori_ori_n399_));
  NA3        o383(.A(ori_ori_n120_), .B(ori_ori_n229_), .C(x0), .Y(ori_ori_n400_));
  OAI210     o384(.A0(ori_ori_n201_), .A1(ori_ori_n68_), .B0(ori_ori_n211_), .Y(ori_ori_n401_));
  NO2        o385(.A(ori_ori_n401_), .B(ori_ori_n25_), .Y(ori_ori_n402_));
  AOI210     o386(.A0(ori_ori_n119_), .A1(ori_ori_n117_), .B0(ori_ori_n42_), .Y(ori_ori_n403_));
  NOi31      o387(.An(ori_ori_n403_), .B(ori_ori_n369_), .C(ori_ori_n186_), .Y(ori_ori_n404_));
  OAI210     o388(.A0(ori_ori_n404_), .A1(ori_ori_n402_), .B0(ori_ori_n152_), .Y(ori_ori_n405_));
  NAi31      o389(.An(ori_ori_n50_), .B(ori_ori_n296_), .C(ori_ori_n181_), .Y(ori_ori_n406_));
  NA3        o390(.A(ori_ori_n406_), .B(ori_ori_n405_), .C(ori_ori_n400_), .Y(ori_ori_n407_));
  OAI210     o391(.A0(ori_ori_n407_), .A1(ori_ori_n399_), .B0(x6), .Y(ori_ori_n408_));
  OAI210     o392(.A0(ori_ori_n167_), .A1(ori_ori_n48_), .B0(ori_ori_n136_), .Y(ori_ori_n409_));
  NA3        o393(.A(ori_ori_n55_), .B(ori_ori_n38_), .C(ori_ori_n31_), .Y(ori_ori_n410_));
  AOI220     o394(.A0(ori_ori_n410_), .A1(ori_ori_n409_), .B0(ori_ori_n40_), .B1(ori_ori_n32_), .Y(ori_ori_n411_));
  NO2        o395(.A(ori_ori_n156_), .B(x0), .Y(ori_ori_n412_));
  AOI220     o396(.A0(ori_ori_n412_), .A1(ori_ori_n229_), .B0(ori_ori_n201_), .B1(ori_ori_n156_), .Y(ori_ori_n413_));
  AOI210     o397(.A0(ori_ori_n127_), .A1(ori_ori_n260_), .B0(x1), .Y(ori_ori_n414_));
  OAI210     o398(.A0(ori_ori_n413_), .A1(x8), .B0(ori_ori_n414_), .Y(ori_ori_n415_));
  NAi31      o399(.An(x2), .B(x8), .C(x0), .Y(ori_ori_n416_));
  OAI210     o400(.A0(ori_ori_n416_), .A1(x4), .B0(ori_ori_n168_), .Y(ori_ori_n417_));
  NA3        o401(.A(ori_ori_n417_), .B(ori_ori_n150_), .C(x9), .Y(ori_ori_n418_));
  NO4        o402(.A(ori_ori_n126_), .B(ori_ori_n307_), .C(x9), .D(x2), .Y(ori_ori_n419_));
  NOi21      o403(.An(ori_ori_n124_), .B(ori_ori_n185_), .Y(ori_ori_n420_));
  NO3        o404(.A(ori_ori_n420_), .B(ori_ori_n419_), .C(ori_ori_n18_), .Y(ori_ori_n421_));
  NO3        o405(.A(x9), .B(ori_ori_n156_), .C(x0), .Y(ori_ori_n422_));
  AOI220     o406(.A0(ori_ori_n422_), .A1(ori_ori_n255_), .B0(ori_ori_n373_), .B1(ori_ori_n156_), .Y(ori_ori_n423_));
  NA4        o407(.A(ori_ori_n423_), .B(ori_ori_n421_), .C(ori_ori_n418_), .D(ori_ori_n50_), .Y(ori_ori_n424_));
  OAI210     o408(.A0(ori_ori_n415_), .A1(ori_ori_n411_), .B0(ori_ori_n424_), .Y(ori_ori_n425_));
  NOi31      o409(.An(ori_ori_n412_), .B(ori_ori_n32_), .C(x8), .Y(ori_ori_n426_));
  AOI210     o410(.A0(ori_ori_n38_), .A1(x9), .B0(ori_ori_n134_), .Y(ori_ori_n427_));
  NO3        o411(.A(ori_ori_n427_), .B(ori_ori_n124_), .C(ori_ori_n43_), .Y(ori_ori_n428_));
  NOi31      o412(.An(x1), .B(x8), .C(x7), .Y(ori_ori_n429_));
  AOI220     o413(.A0(ori_ori_n429_), .A1(ori_ori_n356_), .B0(ori_ori_n125_), .B1(x3), .Y(ori_ori_n430_));
  AOI210     o414(.A0(ori_ori_n273_), .A1(ori_ori_n60_), .B0(ori_ori_n123_), .Y(ori_ori_n431_));
  OAI210     o415(.A0(ori_ori_n431_), .A1(x3), .B0(ori_ori_n430_), .Y(ori_ori_n432_));
  NO3        o416(.A(ori_ori_n432_), .B(ori_ori_n428_), .C(x2), .Y(ori_ori_n433_));
  OAI220     o417(.A0(ori_ori_n357_), .A1(ori_ori_n311_), .B0(ori_ori_n307_), .B1(ori_ori_n43_), .Y(ori_ori_n434_));
  AOI210     o418(.A0(x9), .A1(ori_ori_n48_), .B0(ori_ori_n395_), .Y(ori_ori_n435_));
  AOI220     o419(.A0(ori_ori_n435_), .A1(ori_ori_n90_), .B0(ori_ori_n434_), .B1(ori_ori_n156_), .Y(ori_ori_n436_));
  NO2        o420(.A(ori_ori_n436_), .B(ori_ori_n54_), .Y(ori_ori_n437_));
  NO3        o421(.A(ori_ori_n437_), .B(ori_ori_n433_), .C(ori_ori_n426_), .Y(ori_ori_n438_));
  AOI210     o422(.A0(ori_ori_n438_), .A1(ori_ori_n425_), .B0(ori_ori_n25_), .Y(ori_ori_n439_));
  NA4        o423(.A(ori_ori_n31_), .B(ori_ori_n90_), .C(x2), .D(ori_ori_n17_), .Y(ori_ori_n440_));
  NO3        o424(.A(ori_ori_n62_), .B(x4), .C(x1), .Y(ori_ori_n441_));
  NO3        o425(.A(ori_ori_n68_), .B(ori_ori_n18_), .C(x0), .Y(ori_ori_n442_));
  AOI220     o426(.A0(ori_ori_n442_), .A1(ori_ori_n274_), .B0(ori_ori_n441_), .B1(ori_ori_n403_), .Y(ori_ori_n443_));
  NO2        o427(.A(ori_ori_n443_), .B(ori_ori_n102_), .Y(ori_ori_n444_));
  NO3        o428(.A(ori_ori_n278_), .B(ori_ori_n180_), .C(ori_ori_n40_), .Y(ori_ori_n445_));
  OAI210     o429(.A0(ori_ori_n445_), .A1(ori_ori_n444_), .B0(x7), .Y(ori_ori_n446_));
  NA2        o430(.A(ori_ori_n234_), .B(x7), .Y(ori_ori_n447_));
  NA3        o431(.A(ori_ori_n447_), .B(ori_ori_n155_), .C(ori_ori_n135_), .Y(ori_ori_n448_));
  NA3        o432(.A(ori_ori_n448_), .B(ori_ori_n446_), .C(ori_ori_n440_), .Y(ori_ori_n449_));
  OAI210     o433(.A0(ori_ori_n449_), .A1(ori_ori_n439_), .B0(ori_ori_n36_), .Y(ori_ori_n450_));
  NO2        o434(.A(ori_ori_n422_), .B(ori_ori_n211_), .Y(ori_ori_n451_));
  NO4        o435(.A(ori_ori_n451_), .B(ori_ori_n78_), .C(x4), .D(ori_ori_n54_), .Y(ori_ori_n452_));
  NA2        o436(.A(ori_ori_n263_), .B(ori_ori_n21_), .Y(ori_ori_n453_));
  NO2        o437(.A(ori_ori_n164_), .B(ori_ori_n136_), .Y(ori_ori_n454_));
  NA2        o438(.A(ori_ori_n454_), .B(ori_ori_n453_), .Y(ori_ori_n455_));
  AOI210     o439(.A0(ori_ori_n455_), .A1(ori_ori_n171_), .B0(ori_ori_n28_), .Y(ori_ori_n456_));
  AOI220     o440(.A0(ori_ori_n369_), .A1(ori_ori_n90_), .B0(ori_ori_n153_), .B1(ori_ori_n204_), .Y(ori_ori_n457_));
  NA3        o441(.A(ori_ori_n457_), .B(ori_ori_n416_), .C(ori_ori_n88_), .Y(ori_ori_n458_));
  NA2        o442(.A(ori_ori_n458_), .B(ori_ori_n181_), .Y(ori_ori_n459_));
  OAI220     o443(.A0(ori_ori_n283_), .A1(ori_ori_n69_), .B0(ori_ori_n164_), .B1(ori_ori_n43_), .Y(ori_ori_n460_));
  NA2        o444(.A(x3), .B(ori_ori_n54_), .Y(ori_ori_n461_));
  AOI210     o445(.A0(ori_ori_n168_), .A1(ori_ori_n27_), .B0(ori_ori_n73_), .Y(ori_ori_n462_));
  OAI210     o446(.A0(ori_ori_n152_), .A1(ori_ori_n18_), .B0(ori_ori_n21_), .Y(ori_ori_n463_));
  NO3        o447(.A(ori_ori_n429_), .B(x3), .C(ori_ori_n54_), .Y(ori_ori_n464_));
  AOI210     o448(.A0(ori_ori_n464_), .A1(ori_ori_n463_), .B0(ori_ori_n462_), .Y(ori_ori_n465_));
  OAI210     o449(.A0(ori_ori_n157_), .A1(ori_ori_n461_), .B0(ori_ori_n465_), .Y(ori_ori_n466_));
  AOI220     o450(.A0(ori_ori_n466_), .A1(x0), .B0(ori_ori_n460_), .B1(ori_ori_n136_), .Y(ori_ori_n467_));
  AOI210     o451(.A0(ori_ori_n467_), .A1(ori_ori_n459_), .B0(ori_ori_n242_), .Y(ori_ori_n468_));
  NO3        o452(.A(ori_ori_n468_), .B(ori_ori_n456_), .C(ori_ori_n452_), .Y(ori_ori_n469_));
  NA3        o453(.A(ori_ori_n469_), .B(ori_ori_n450_), .C(ori_ori_n408_), .Y(ori_ori_n470_));
  AOI210     o454(.A0(ori_ori_n389_), .A1(ori_ori_n25_), .B0(ori_ori_n470_), .Y(ori05));
  INV        m000(.A(x0), .Y(mai_mai_n17_));
  INV        m001(.A(x1), .Y(mai_mai_n18_));
  NO2        m002(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n19_));
  NO2        m003(.A(x6), .B(x5), .Y(mai_mai_n20_));
  OR2        m004(.A(x8), .B(x7), .Y(mai_mai_n21_));
  NOi21      m005(.An(mai_mai_n20_), .B(mai_mai_n21_), .Y(mai_mai_n22_));
  NAi21      m006(.An(mai_mai_n22_), .B(mai_mai_n19_), .Y(mai_mai_n23_));
  NA2        m007(.A(mai_mai_n18_), .B(mai_mai_n17_), .Y(mai_mai_n24_));
  INV        m008(.A(x5), .Y(mai_mai_n25_));
  NA2        m009(.A(x7), .B(x6), .Y(mai_mai_n26_));
  NA2        m010(.A(x8), .B(x3), .Y(mai_mai_n27_));
  NA2        m011(.A(x4), .B(x2), .Y(mai_mai_n28_));
  INV        m012(.A(mai_mai_n24_), .Y(mai_mai_n29_));
  NO2        m013(.A(x4), .B(x3), .Y(mai_mai_n30_));
  INV        m014(.A(mai_mai_n30_), .Y(mai_mai_n31_));
  OA210      m015(.A0(mai_mai_n31_), .A1(x2), .B0(mai_mai_n19_), .Y(mai_mai_n32_));
  NOi31      m016(.An(mai_mai_n23_), .B(mai_mai_n32_), .C(mai_mai_n29_), .Y(mai00));
  NO2        m017(.A(x1), .B(x0), .Y(mai_mai_n34_));
  INV        m018(.A(x6), .Y(mai_mai_n35_));
  NO2        m019(.A(mai_mai_n35_), .B(mai_mai_n25_), .Y(mai_mai_n36_));
  AN2        m020(.A(x8), .B(x7), .Y(mai_mai_n37_));
  NA2        m021(.A(x4), .B(x3), .Y(mai_mai_n38_));
  NO2        m022(.A(mai_mai_n23_), .B(mai_mai_n38_), .Y(mai_mai_n39_));
  NO2        m023(.A(x2), .B(x0), .Y(mai_mai_n40_));
  INV        m024(.A(x3), .Y(mai_mai_n41_));
  NO2        m025(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n42_));
  INV        m026(.A(mai_mai_n42_), .Y(mai_mai_n43_));
  NO2        m027(.A(mai_mai_n36_), .B(x4), .Y(mai_mai_n44_));
  OAI210     m028(.A0(mai_mai_n44_), .A1(mai_mai_n43_), .B0(mai_mai_n40_), .Y(mai_mai_n45_));
  INV        m029(.A(x4), .Y(mai_mai_n46_));
  NO2        m030(.A(mai_mai_n46_), .B(mai_mai_n17_), .Y(mai_mai_n47_));
  NA2        m031(.A(mai_mai_n47_), .B(x2), .Y(mai_mai_n48_));
  OAI210     m032(.A0(mai_mai_n48_), .A1(mai_mai_n20_), .B0(mai_mai_n45_), .Y(mai_mai_n49_));
  NA2        m033(.A(mai_mai_n37_), .B(mai_mai_n36_), .Y(mai_mai_n50_));
  AOI220     m034(.A0(mai_mai_n50_), .A1(mai_mai_n34_), .B0(mai_mai_n22_), .B1(mai_mai_n19_), .Y(mai_mai_n51_));
  INV        m035(.A(x2), .Y(mai_mai_n52_));
  NO2        m036(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n53_));
  NA2        m037(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n54_));
  NA2        m038(.A(mai_mai_n54_), .B(mai_mai_n53_), .Y(mai_mai_n55_));
  OAI210     m039(.A0(mai_mai_n51_), .A1(mai_mai_n31_), .B0(mai_mai_n55_), .Y(mai_mai_n56_));
  NO3        m040(.A(mai_mai_n56_), .B(mai_mai_n49_), .C(mai_mai_n39_), .Y(mai01));
  NA2        m041(.A(x8), .B(x7), .Y(mai_mai_n58_));
  NA2        m042(.A(mai_mai_n41_), .B(x1), .Y(mai_mai_n59_));
  INV        m043(.A(x9), .Y(mai_mai_n60_));
  NO2        m044(.A(mai_mai_n60_), .B(mai_mai_n35_), .Y(mai_mai_n61_));
  INV        m045(.A(mai_mai_n61_), .Y(mai_mai_n62_));
  NO3        m046(.A(mai_mai_n62_), .B(mai_mai_n59_), .C(mai_mai_n58_), .Y(mai_mai_n63_));
  NO2        m047(.A(x7), .B(x6), .Y(mai_mai_n64_));
  NO2        m048(.A(mai_mai_n59_), .B(x5), .Y(mai_mai_n65_));
  NO2        m049(.A(x8), .B(x2), .Y(mai_mai_n66_));
  INV        m050(.A(mai_mai_n66_), .Y(mai_mai_n67_));
  NO2        m051(.A(mai_mai_n67_), .B(x1), .Y(mai_mai_n68_));
  OA210      m052(.A0(mai_mai_n68_), .A1(mai_mai_n65_), .B0(mai_mai_n64_), .Y(mai_mai_n69_));
  OAI210     m053(.A0(mai_mai_n42_), .A1(mai_mai_n25_), .B0(mai_mai_n52_), .Y(mai_mai_n70_));
  OAI210     m054(.A0(mai_mai_n54_), .A1(mai_mai_n20_), .B0(mai_mai_n70_), .Y(mai_mai_n71_));
  NO2        m055(.A(mai_mai_n71_), .B(mai_mai_n69_), .Y(mai_mai_n72_));
  OAI210     m056(.A0(mai_mai_n72_), .A1(mai_mai_n63_), .B0(x4), .Y(mai_mai_n73_));
  NA2        m057(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n74_));
  OAI210     m058(.A0(mai_mai_n74_), .A1(mai_mai_n54_), .B0(x0), .Y(mai_mai_n75_));
  NA2        m059(.A(x5), .B(x3), .Y(mai_mai_n76_));
  NO2        m060(.A(x8), .B(x6), .Y(mai_mai_n77_));
  NO4        m061(.A(mai_mai_n77_), .B(mai_mai_n76_), .C(mai_mai_n64_), .D(mai_mai_n52_), .Y(mai_mai_n78_));
  NAi21      m062(.An(x4), .B(x3), .Y(mai_mai_n79_));
  INV        m063(.A(mai_mai_n79_), .Y(mai_mai_n80_));
  NO2        m064(.A(mai_mai_n80_), .B(mai_mai_n22_), .Y(mai_mai_n81_));
  NO2        m065(.A(x4), .B(x2), .Y(mai_mai_n82_));
  NO2        m066(.A(mai_mai_n82_), .B(x3), .Y(mai_mai_n83_));
  NO3        m067(.A(mai_mai_n83_), .B(mai_mai_n81_), .C(mai_mai_n18_), .Y(mai_mai_n84_));
  NO3        m068(.A(mai_mai_n84_), .B(mai_mai_n78_), .C(mai_mai_n75_), .Y(mai_mai_n85_));
  NO4        m069(.A(mai_mai_n21_), .B(x6), .C(mai_mai_n41_), .D(x1), .Y(mai_mai_n86_));
  NA2        m070(.A(mai_mai_n60_), .B(mai_mai_n46_), .Y(mai_mai_n87_));
  INV        m071(.A(mai_mai_n87_), .Y(mai_mai_n88_));
  OAI210     m072(.A0(mai_mai_n86_), .A1(mai_mai_n65_), .B0(mai_mai_n88_), .Y(mai_mai_n89_));
  NA2        m073(.A(x3), .B(mai_mai_n18_), .Y(mai_mai_n90_));
  NO2        m074(.A(mai_mai_n90_), .B(mai_mai_n25_), .Y(mai_mai_n91_));
  INV        m075(.A(x8), .Y(mai_mai_n92_));
  NA2        m076(.A(x2), .B(x1), .Y(mai_mai_n93_));
  NO2        m077(.A(mai_mai_n93_), .B(mai_mai_n92_), .Y(mai_mai_n94_));
  NO2        m078(.A(mai_mai_n94_), .B(mai_mai_n91_), .Y(mai_mai_n95_));
  NO2        m079(.A(mai_mai_n95_), .B(mai_mai_n26_), .Y(mai_mai_n96_));
  AOI210     m080(.A0(mai_mai_n54_), .A1(mai_mai_n25_), .B0(mai_mai_n52_), .Y(mai_mai_n97_));
  OAI210     m081(.A0(mai_mai_n43_), .A1(mai_mai_n36_), .B0(mai_mai_n46_), .Y(mai_mai_n98_));
  NO3        m082(.A(mai_mai_n98_), .B(mai_mai_n97_), .C(mai_mai_n96_), .Y(mai_mai_n99_));
  NA2        m083(.A(x4), .B(mai_mai_n41_), .Y(mai_mai_n100_));
  NO2        m084(.A(mai_mai_n46_), .B(mai_mai_n52_), .Y(mai_mai_n101_));
  NA2        m085(.A(mai_mai_n41_), .B(mai_mai_n18_), .Y(mai_mai_n102_));
  AOI210     m086(.A0(mai_mai_n100_), .A1(mai_mai_n50_), .B0(mai_mai_n102_), .Y(mai_mai_n103_));
  NO2        m087(.A(x3), .B(x2), .Y(mai_mai_n104_));
  NA3        m088(.A(mai_mai_n104_), .B(mai_mai_n26_), .C(mai_mai_n25_), .Y(mai_mai_n105_));
  AOI210     m089(.A0(x8), .A1(x6), .B0(mai_mai_n105_), .Y(mai_mai_n106_));
  NA2        m090(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n107_));
  OAI210     m091(.A0(mai_mai_n107_), .A1(mai_mai_n38_), .B0(mai_mai_n17_), .Y(mai_mai_n108_));
  NO4        m092(.A(mai_mai_n108_), .B(mai_mai_n106_), .C(mai_mai_n103_), .D(mai_mai_n99_), .Y(mai_mai_n109_));
  AO220      m093(.A0(mai_mai_n109_), .A1(mai_mai_n89_), .B0(mai_mai_n85_), .B1(mai_mai_n73_), .Y(mai02));
  NO2        m094(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n111_));
  NO2        m095(.A(x8), .B(mai_mai_n18_), .Y(mai_mai_n112_));
  NA2        m096(.A(mai_mai_n52_), .B(mai_mai_n17_), .Y(mai_mai_n113_));
  NA2        m097(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n114_));
  OAI210     m098(.A0(mai_mai_n87_), .A1(mai_mai_n113_), .B0(mai_mai_n114_), .Y(mai_mai_n115_));
  AOI220     m099(.A0(mai_mai_n115_), .A1(mai_mai_n112_), .B0(mai_mai_n111_), .B1(x4), .Y(mai_mai_n116_));
  NO3        m100(.A(mai_mai_n116_), .B(x7), .C(x5), .Y(mai_mai_n117_));
  NA2        m101(.A(x9), .B(x2), .Y(mai_mai_n118_));
  OR2        m102(.A(x8), .B(x0), .Y(mai_mai_n119_));
  INV        m103(.A(mai_mai_n119_), .Y(mai_mai_n120_));
  NAi21      m104(.An(x2), .B(x8), .Y(mai_mai_n121_));
  INV        m105(.A(mai_mai_n121_), .Y(mai_mai_n122_));
  OAI220     m106(.A0(mai_mai_n122_), .A1(mai_mai_n120_), .B0(mai_mai_n118_), .B1(x7), .Y(mai_mai_n123_));
  NO2        m107(.A(x4), .B(x1), .Y(mai_mai_n124_));
  NA3        m108(.A(mai_mai_n124_), .B(mai_mai_n123_), .C(mai_mai_n58_), .Y(mai_mai_n125_));
  NOi21      m109(.An(x0), .B(x1), .Y(mai_mai_n126_));
  NO3        m110(.A(x9), .B(x8), .C(x7), .Y(mai_mai_n127_));
  NOi21      m111(.An(x0), .B(x4), .Y(mai_mai_n128_));
  NAi21      m112(.An(x8), .B(x7), .Y(mai_mai_n129_));
  NO2        m113(.A(mai_mai_n129_), .B(mai_mai_n60_), .Y(mai_mai_n130_));
  AOI220     m114(.A0(mai_mai_n130_), .A1(mai_mai_n128_), .B0(mai_mai_n127_), .B1(mai_mai_n126_), .Y(mai_mai_n131_));
  AOI210     m115(.A0(mai_mai_n131_), .A1(mai_mai_n125_), .B0(mai_mai_n76_), .Y(mai_mai_n132_));
  NO2        m116(.A(x5), .B(mai_mai_n46_), .Y(mai_mai_n133_));
  NA2        m117(.A(x2), .B(mai_mai_n18_), .Y(mai_mai_n134_));
  AOI210     m118(.A0(mai_mai_n134_), .A1(mai_mai_n107_), .B0(mai_mai_n114_), .Y(mai_mai_n135_));
  OAI210     m119(.A0(mai_mai_n135_), .A1(mai_mai_n34_), .B0(mai_mai_n133_), .Y(mai_mai_n136_));
  NAi21      m120(.An(x0), .B(x4), .Y(mai_mai_n137_));
  NO2        m121(.A(mai_mai_n137_), .B(x1), .Y(mai_mai_n138_));
  NO2        m122(.A(x7), .B(x0), .Y(mai_mai_n139_));
  NO2        m123(.A(mai_mai_n82_), .B(mai_mai_n101_), .Y(mai_mai_n140_));
  NO2        m124(.A(mai_mai_n140_), .B(x3), .Y(mai_mai_n141_));
  OAI210     m125(.A0(mai_mai_n139_), .A1(mai_mai_n138_), .B0(mai_mai_n141_), .Y(mai_mai_n142_));
  NO2        m126(.A(mai_mai_n21_), .B(mai_mai_n41_), .Y(mai_mai_n143_));
  NA2        m127(.A(x5), .B(x0), .Y(mai_mai_n144_));
  NO2        m128(.A(mai_mai_n46_), .B(x2), .Y(mai_mai_n145_));
  NA3        m129(.A(mai_mai_n145_), .B(mai_mai_n144_), .C(mai_mai_n143_), .Y(mai_mai_n146_));
  NA4        m130(.A(mai_mai_n146_), .B(mai_mai_n142_), .C(mai_mai_n136_), .D(mai_mai_n35_), .Y(mai_mai_n147_));
  NO3        m131(.A(mai_mai_n147_), .B(mai_mai_n132_), .C(mai_mai_n117_), .Y(mai_mai_n148_));
  NO3        m132(.A(mai_mai_n76_), .B(mai_mai_n74_), .C(mai_mai_n24_), .Y(mai_mai_n149_));
  NO2        m133(.A(mai_mai_n28_), .B(mai_mai_n25_), .Y(mai_mai_n150_));
  AOI220     m134(.A0(mai_mai_n126_), .A1(mai_mai_n150_), .B0(mai_mai_n65_), .B1(mai_mai_n17_), .Y(mai_mai_n151_));
  NO3        m135(.A(mai_mai_n151_), .B(mai_mai_n58_), .C(mai_mai_n60_), .Y(mai_mai_n152_));
  NA2        m136(.A(x7), .B(x3), .Y(mai_mai_n153_));
  NO2        m137(.A(mai_mai_n100_), .B(x5), .Y(mai_mai_n154_));
  NO2        m138(.A(x9), .B(x7), .Y(mai_mai_n155_));
  NOi21      m139(.An(x8), .B(x0), .Y(mai_mai_n156_));
  OA210      m140(.A0(mai_mai_n155_), .A1(x1), .B0(mai_mai_n156_), .Y(mai_mai_n157_));
  NO2        m141(.A(mai_mai_n41_), .B(x2), .Y(mai_mai_n158_));
  INV        m142(.A(x7), .Y(mai_mai_n159_));
  NA2        m143(.A(mai_mai_n159_), .B(mai_mai_n18_), .Y(mai_mai_n160_));
  AOI220     m144(.A0(mai_mai_n160_), .A1(mai_mai_n158_), .B0(mai_mai_n111_), .B1(mai_mai_n37_), .Y(mai_mai_n161_));
  NO2        m145(.A(mai_mai_n25_), .B(x4), .Y(mai_mai_n162_));
  NO2        m146(.A(mai_mai_n162_), .B(mai_mai_n128_), .Y(mai_mai_n163_));
  NO2        m147(.A(mai_mai_n163_), .B(mai_mai_n161_), .Y(mai_mai_n164_));
  AOI210     m148(.A0(mai_mai_n157_), .A1(mai_mai_n154_), .B0(mai_mai_n164_), .Y(mai_mai_n165_));
  OAI210     m149(.A0(mai_mai_n153_), .A1(mai_mai_n48_), .B0(mai_mai_n165_), .Y(mai_mai_n166_));
  NA2        m150(.A(x5), .B(x1), .Y(mai_mai_n167_));
  INV        m151(.A(mai_mai_n167_), .Y(mai_mai_n168_));
  AOI210     m152(.A0(mai_mai_n168_), .A1(mai_mai_n128_), .B0(mai_mai_n35_), .Y(mai_mai_n169_));
  NO2        m153(.A(mai_mai_n60_), .B(mai_mai_n92_), .Y(mai_mai_n170_));
  NAi21      m154(.An(x2), .B(x7), .Y(mai_mai_n171_));
  NO3        m155(.A(mai_mai_n171_), .B(mai_mai_n170_), .C(mai_mai_n46_), .Y(mai_mai_n172_));
  NA2        m156(.A(mai_mai_n172_), .B(mai_mai_n65_), .Y(mai_mai_n173_));
  NAi31      m157(.An(mai_mai_n76_), .B(mai_mai_n37_), .C(mai_mai_n34_), .Y(mai_mai_n174_));
  NA2        m158(.A(mai_mai_n173_), .B(mai_mai_n169_), .Y(mai_mai_n175_));
  NO4        m159(.A(mai_mai_n175_), .B(mai_mai_n166_), .C(mai_mai_n152_), .D(mai_mai_n149_), .Y(mai_mai_n176_));
  NO2        m160(.A(mai_mai_n176_), .B(mai_mai_n148_), .Y(mai_mai_n177_));
  NO2        m161(.A(mai_mai_n144_), .B(mai_mai_n140_), .Y(mai_mai_n178_));
  NA2        m162(.A(mai_mai_n25_), .B(mai_mai_n18_), .Y(mai_mai_n179_));
  NA2        m163(.A(mai_mai_n25_), .B(mai_mai_n17_), .Y(mai_mai_n180_));
  NA3        m164(.A(mai_mai_n180_), .B(mai_mai_n179_), .C(mai_mai_n24_), .Y(mai_mai_n181_));
  AN2        m165(.A(mai_mai_n181_), .B(mai_mai_n145_), .Y(mai_mai_n182_));
  NA2        m166(.A(x8), .B(x0), .Y(mai_mai_n183_));
  NO2        m167(.A(mai_mai_n159_), .B(mai_mai_n25_), .Y(mai_mai_n184_));
  NO2        m168(.A(mai_mai_n126_), .B(x4), .Y(mai_mai_n185_));
  NA2        m169(.A(mai_mai_n185_), .B(mai_mai_n184_), .Y(mai_mai_n186_));
  AOI210     m170(.A0(mai_mai_n183_), .A1(mai_mai_n134_), .B0(mai_mai_n186_), .Y(mai_mai_n187_));
  NA2        m171(.A(x2), .B(x0), .Y(mai_mai_n188_));
  NA2        m172(.A(x4), .B(x1), .Y(mai_mai_n189_));
  NAi21      m173(.An(mai_mai_n124_), .B(mai_mai_n189_), .Y(mai_mai_n190_));
  NOi31      m174(.An(mai_mai_n190_), .B(mai_mai_n162_), .C(mai_mai_n188_), .Y(mai_mai_n191_));
  NO4        m175(.A(mai_mai_n191_), .B(mai_mai_n187_), .C(mai_mai_n182_), .D(mai_mai_n178_), .Y(mai_mai_n192_));
  NO2        m176(.A(mai_mai_n192_), .B(mai_mai_n41_), .Y(mai_mai_n193_));
  NO2        m177(.A(mai_mai_n181_), .B(mai_mai_n74_), .Y(mai_mai_n194_));
  INV        m178(.A(mai_mai_n133_), .Y(mai_mai_n195_));
  NO2        m179(.A(mai_mai_n107_), .B(mai_mai_n17_), .Y(mai_mai_n196_));
  AOI210     m180(.A0(mai_mai_n34_), .A1(mai_mai_n92_), .B0(mai_mai_n196_), .Y(mai_mai_n197_));
  NO3        m181(.A(mai_mai_n197_), .B(mai_mai_n195_), .C(x7), .Y(mai_mai_n198_));
  NA3        m182(.A(mai_mai_n190_), .B(mai_mai_n195_), .C(mai_mai_n40_), .Y(mai_mai_n199_));
  OAI210     m183(.A0(mai_mai_n180_), .A1(mai_mai_n140_), .B0(mai_mai_n199_), .Y(mai_mai_n200_));
  NO3        m184(.A(mai_mai_n200_), .B(mai_mai_n198_), .C(mai_mai_n194_), .Y(mai_mai_n201_));
  NO2        m185(.A(mai_mai_n201_), .B(x3), .Y(mai_mai_n202_));
  NO3        m186(.A(mai_mai_n202_), .B(mai_mai_n193_), .C(mai_mai_n177_), .Y(mai03));
  NO2        m187(.A(mai_mai_n46_), .B(x3), .Y(mai_mai_n204_));
  NO2        m188(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n205_));
  INV        m189(.A(mai_mai_n205_), .Y(mai_mai_n206_));
  NO2        m190(.A(mai_mai_n52_), .B(x1), .Y(mai_mai_n207_));
  OAI210     m191(.A0(mai_mai_n207_), .A1(mai_mai_n25_), .B0(mai_mai_n61_), .Y(mai_mai_n208_));
  OAI220     m192(.A0(mai_mai_n208_), .A1(mai_mai_n17_), .B0(mai_mai_n206_), .B1(mai_mai_n107_), .Y(mai_mai_n209_));
  NA2        m193(.A(mai_mai_n209_), .B(mai_mai_n204_), .Y(mai_mai_n210_));
  NO2        m194(.A(mai_mai_n76_), .B(x6), .Y(mai_mai_n211_));
  NA2        m195(.A(x6), .B(mai_mai_n25_), .Y(mai_mai_n212_));
  NO2        m196(.A(mai_mai_n212_), .B(x4), .Y(mai_mai_n213_));
  NO2        m197(.A(mai_mai_n18_), .B(x0), .Y(mai_mai_n214_));
  AO220      m198(.A0(mai_mai_n214_), .A1(mai_mai_n213_), .B0(mai_mai_n211_), .B1(mai_mai_n53_), .Y(mai_mai_n215_));
  NA2        m199(.A(mai_mai_n215_), .B(mai_mai_n60_), .Y(mai_mai_n216_));
  NA2        m200(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n217_));
  NO2        m201(.A(mai_mai_n217_), .B(mai_mai_n212_), .Y(mai_mai_n218_));
  NA2        m202(.A(x9), .B(mai_mai_n52_), .Y(mai_mai_n219_));
  NA2        m203(.A(mai_mai_n219_), .B(x4), .Y(mai_mai_n220_));
  NA2        m204(.A(mai_mai_n212_), .B(mai_mai_n79_), .Y(mai_mai_n221_));
  AOI210     m205(.A0(mai_mai_n25_), .A1(x3), .B0(mai_mai_n188_), .Y(mai_mai_n222_));
  AOI220     m206(.A0(mai_mai_n222_), .A1(mai_mai_n221_), .B0(mai_mai_n220_), .B1(mai_mai_n218_), .Y(mai_mai_n223_));
  NO3        m207(.A(x6), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n224_));
  NO2        m208(.A(x5), .B(x1), .Y(mai_mai_n225_));
  AOI220     m209(.A0(mai_mai_n225_), .A1(mai_mai_n17_), .B0(mai_mai_n104_), .B1(x5), .Y(mai_mai_n226_));
  NO2        m210(.A(mai_mai_n217_), .B(mai_mai_n179_), .Y(mai_mai_n227_));
  NO3        m211(.A(x3), .B(x2), .C(x1), .Y(mai_mai_n228_));
  NO2        m212(.A(mai_mai_n228_), .B(mai_mai_n227_), .Y(mai_mai_n229_));
  OAI210     m213(.A0(mai_mai_n226_), .A1(mai_mai_n62_), .B0(mai_mai_n229_), .Y(mai_mai_n230_));
  AOI220     m214(.A0(mai_mai_n230_), .A1(mai_mai_n46_), .B0(mai_mai_n224_), .B1(mai_mai_n133_), .Y(mai_mai_n231_));
  NA4        m215(.A(mai_mai_n231_), .B(mai_mai_n223_), .C(mai_mai_n216_), .D(mai_mai_n210_), .Y(mai_mai_n232_));
  NO2        m216(.A(mai_mai_n46_), .B(mai_mai_n41_), .Y(mai_mai_n233_));
  NA2        m217(.A(mai_mai_n233_), .B(mai_mai_n19_), .Y(mai_mai_n234_));
  NO2        m218(.A(x3), .B(mai_mai_n17_), .Y(mai_mai_n235_));
  NO2        m219(.A(mai_mai_n235_), .B(x6), .Y(mai_mai_n236_));
  NOi21      m220(.An(mai_mai_n82_), .B(mai_mai_n236_), .Y(mai_mai_n237_));
  NA2        m221(.A(mai_mai_n60_), .B(mai_mai_n92_), .Y(mai_mai_n238_));
  NA3        m222(.A(mai_mai_n238_), .B(mai_mai_n235_), .C(x6), .Y(mai_mai_n239_));
  AOI210     m223(.A0(mai_mai_n239_), .A1(mai_mai_n237_), .B0(mai_mai_n159_), .Y(mai_mai_n240_));
  AO210      m224(.A0(mai_mai_n240_), .A1(mai_mai_n234_), .B0(mai_mai_n184_), .Y(mai_mai_n241_));
  NA2        m225(.A(mai_mai_n41_), .B(mai_mai_n52_), .Y(mai_mai_n242_));
  NA2        m226(.A(mai_mai_n145_), .B(mai_mai_n91_), .Y(mai_mai_n243_));
  NA2        m227(.A(x6), .B(mai_mai_n46_), .Y(mai_mai_n244_));
  OAI210     m228(.A0(mai_mai_n120_), .A1(mai_mai_n77_), .B0(x4), .Y(mai_mai_n245_));
  AOI210     m229(.A0(mai_mai_n245_), .A1(mai_mai_n244_), .B0(mai_mai_n76_), .Y(mai_mai_n246_));
  NO2        m230(.A(mai_mai_n60_), .B(x6), .Y(mai_mai_n247_));
  NO2        m231(.A(mai_mai_n167_), .B(mai_mai_n41_), .Y(mai_mai_n248_));
  OAI210     m232(.A0(mai_mai_n248_), .A1(mai_mai_n227_), .B0(mai_mai_n247_), .Y(mai_mai_n249_));
  NA2        m233(.A(mai_mai_n205_), .B(mai_mai_n138_), .Y(mai_mai_n250_));
  NA3        m234(.A(mai_mai_n217_), .B(mai_mai_n133_), .C(x6), .Y(mai_mai_n251_));
  OAI210     m235(.A0(mai_mai_n92_), .A1(mai_mai_n35_), .B0(mai_mai_n65_), .Y(mai_mai_n252_));
  NA4        m236(.A(mai_mai_n252_), .B(mai_mai_n251_), .C(mai_mai_n250_), .D(mai_mai_n249_), .Y(mai_mai_n253_));
  OAI210     m237(.A0(mai_mai_n253_), .A1(mai_mai_n246_), .B0(x2), .Y(mai_mai_n254_));
  NA3        m238(.A(mai_mai_n254_), .B(mai_mai_n243_), .C(mai_mai_n241_), .Y(mai_mai_n255_));
  AOI210     m239(.A0(mai_mai_n232_), .A1(x8), .B0(mai_mai_n255_), .Y(mai_mai_n256_));
  NO2        m240(.A(mai_mai_n92_), .B(x3), .Y(mai_mai_n257_));
  NA2        m241(.A(mai_mai_n257_), .B(mai_mai_n213_), .Y(mai_mai_n258_));
  NO3        m242(.A(mai_mai_n90_), .B(mai_mai_n77_), .C(mai_mai_n25_), .Y(mai_mai_n259_));
  AOI210     m243(.A0(mai_mai_n236_), .A1(mai_mai_n162_), .B0(mai_mai_n259_), .Y(mai_mai_n260_));
  AOI210     m244(.A0(mai_mai_n260_), .A1(mai_mai_n258_), .B0(x2), .Y(mai_mai_n261_));
  NO2        m245(.A(x4), .B(mai_mai_n52_), .Y(mai_mai_n262_));
  AOI220     m246(.A0(mai_mai_n213_), .A1(mai_mai_n196_), .B0(mai_mai_n262_), .B1(mai_mai_n65_), .Y(mai_mai_n263_));
  NA2        m247(.A(mai_mai_n60_), .B(x6), .Y(mai_mai_n264_));
  NA3        m248(.A(mai_mai_n25_), .B(x3), .C(x2), .Y(mai_mai_n265_));
  AOI210     m249(.A0(mai_mai_n265_), .A1(mai_mai_n144_), .B0(mai_mai_n264_), .Y(mai_mai_n266_));
  NA2        m250(.A(mai_mai_n41_), .B(mai_mai_n17_), .Y(mai_mai_n267_));
  NO2        m251(.A(mai_mai_n267_), .B(mai_mai_n25_), .Y(mai_mai_n268_));
  OAI210     m252(.A0(mai_mai_n268_), .A1(mai_mai_n266_), .B0(mai_mai_n124_), .Y(mai_mai_n269_));
  NA2        m253(.A(mai_mai_n217_), .B(x6), .Y(mai_mai_n270_));
  NO2        m254(.A(mai_mai_n217_), .B(x6), .Y(mai_mai_n271_));
  NAi21      m255(.An(mai_mai_n170_), .B(mai_mai_n271_), .Y(mai_mai_n272_));
  NA3        m256(.A(mai_mai_n272_), .B(mai_mai_n270_), .C(mai_mai_n150_), .Y(mai_mai_n273_));
  NA4        m257(.A(mai_mai_n273_), .B(mai_mai_n269_), .C(mai_mai_n263_), .D(mai_mai_n159_), .Y(mai_mai_n274_));
  NA2        m258(.A(mai_mai_n205_), .B(mai_mai_n235_), .Y(mai_mai_n275_));
  NO2        m259(.A(x9), .B(x6), .Y(mai_mai_n276_));
  NO2        m260(.A(mai_mai_n144_), .B(mai_mai_n18_), .Y(mai_mai_n277_));
  NAi21      m261(.An(mai_mai_n277_), .B(mai_mai_n265_), .Y(mai_mai_n278_));
  NAi21      m262(.An(x1), .B(x4), .Y(mai_mai_n279_));
  AOI210     m263(.A0(x3), .A1(x2), .B0(mai_mai_n46_), .Y(mai_mai_n280_));
  OAI210     m264(.A0(mai_mai_n144_), .A1(x3), .B0(mai_mai_n280_), .Y(mai_mai_n281_));
  AOI220     m265(.A0(mai_mai_n281_), .A1(mai_mai_n279_), .B0(mai_mai_n278_), .B1(mai_mai_n276_), .Y(mai_mai_n282_));
  NA2        m266(.A(mai_mai_n282_), .B(mai_mai_n275_), .Y(mai_mai_n283_));
  NA2        m267(.A(mai_mai_n60_), .B(x2), .Y(mai_mai_n284_));
  NO2        m268(.A(mai_mai_n284_), .B(mai_mai_n275_), .Y(mai_mai_n285_));
  NO3        m269(.A(x9), .B(x6), .C(x0), .Y(mai_mai_n286_));
  NA2        m270(.A(mai_mai_n107_), .B(mai_mai_n25_), .Y(mai_mai_n287_));
  NA2        m271(.A(x6), .B(x2), .Y(mai_mai_n288_));
  NO2        m272(.A(mai_mai_n288_), .B(mai_mai_n179_), .Y(mai_mai_n289_));
  AOI210     m273(.A0(mai_mai_n287_), .A1(mai_mai_n286_), .B0(mai_mai_n289_), .Y(mai_mai_n290_));
  OAI220     m274(.A0(mai_mai_n290_), .A1(mai_mai_n41_), .B0(mai_mai_n185_), .B1(mai_mai_n44_), .Y(mai_mai_n291_));
  OAI210     m275(.A0(mai_mai_n291_), .A1(mai_mai_n285_), .B0(mai_mai_n283_), .Y(mai_mai_n292_));
  NA2        m276(.A(x9), .B(mai_mai_n41_), .Y(mai_mai_n293_));
  NO2        m277(.A(mai_mai_n293_), .B(mai_mai_n212_), .Y(mai_mai_n294_));
  OR3        m278(.A(mai_mai_n294_), .B(mai_mai_n211_), .C(mai_mai_n154_), .Y(mai_mai_n295_));
  NA2        m279(.A(x4), .B(x0), .Y(mai_mai_n296_));
  NA2        m280(.A(mai_mai_n295_), .B(mai_mai_n40_), .Y(mai_mai_n297_));
  AOI210     m281(.A0(mai_mai_n297_), .A1(mai_mai_n292_), .B0(x8), .Y(mai_mai_n298_));
  INV        m282(.A(mai_mai_n264_), .Y(mai_mai_n299_));
  NA2        m283(.A(mai_mai_n225_), .B(mai_mai_n299_), .Y(mai_mai_n300_));
  INV        m284(.A(mai_mai_n183_), .Y(mai_mai_n301_));
  OAI210     m285(.A0(mai_mai_n301_), .A1(x4), .B0(mai_mai_n20_), .Y(mai_mai_n302_));
  AOI210     m286(.A0(mai_mai_n302_), .A1(mai_mai_n300_), .B0(mai_mai_n242_), .Y(mai_mai_n303_));
  NO4        m287(.A(mai_mai_n303_), .B(mai_mai_n298_), .C(mai_mai_n274_), .D(mai_mai_n261_), .Y(mai_mai_n304_));
  NO2        m288(.A(mai_mai_n170_), .B(x1), .Y(mai_mai_n305_));
  NO3        m289(.A(mai_mai_n305_), .B(x3), .C(mai_mai_n35_), .Y(mai_mai_n306_));
  OAI210     m290(.A0(mai_mai_n306_), .A1(mai_mai_n271_), .B0(x2), .Y(mai_mai_n307_));
  OAI210     m291(.A0(mai_mai_n301_), .A1(x6), .B0(mai_mai_n42_), .Y(mai_mai_n308_));
  AOI210     m292(.A0(mai_mai_n308_), .A1(mai_mai_n307_), .B0(mai_mai_n195_), .Y(mai_mai_n309_));
  NOi21      m293(.An(mai_mai_n288_), .B(mai_mai_n17_), .Y(mai_mai_n310_));
  NA3        m294(.A(mai_mai_n310_), .B(mai_mai_n225_), .C(mai_mai_n38_), .Y(mai_mai_n311_));
  AOI210     m295(.A0(mai_mai_n35_), .A1(mai_mai_n52_), .B0(x0), .Y(mai_mai_n312_));
  NA3        m296(.A(mai_mai_n312_), .B(mai_mai_n168_), .C(mai_mai_n31_), .Y(mai_mai_n313_));
  NA2        m297(.A(x3), .B(x2), .Y(mai_mai_n314_));
  AOI220     m298(.A0(mai_mai_n314_), .A1(mai_mai_n242_), .B0(mai_mai_n313_), .B1(mai_mai_n311_), .Y(mai_mai_n315_));
  NAi21      m299(.An(x4), .B(x0), .Y(mai_mai_n316_));
  NO3        m300(.A(mai_mai_n316_), .B(mai_mai_n42_), .C(x2), .Y(mai_mai_n317_));
  OAI210     m301(.A0(x6), .A1(mai_mai_n18_), .B0(mai_mai_n317_), .Y(mai_mai_n318_));
  OAI220     m302(.A0(mai_mai_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(mai_mai_n319_));
  NO2        m303(.A(x9), .B(x8), .Y(mai_mai_n320_));
  NA3        m304(.A(mai_mai_n320_), .B(mai_mai_n35_), .C(mai_mai_n52_), .Y(mai_mai_n321_));
  OAI210     m305(.A0(mai_mai_n312_), .A1(mai_mai_n310_), .B0(mai_mai_n321_), .Y(mai_mai_n322_));
  AOI220     m306(.A0(mai_mai_n322_), .A1(mai_mai_n80_), .B0(mai_mai_n319_), .B1(mai_mai_n30_), .Y(mai_mai_n323_));
  AOI210     m307(.A0(mai_mai_n323_), .A1(mai_mai_n318_), .B0(mai_mai_n25_), .Y(mai_mai_n324_));
  NA3        m308(.A(mai_mai_n35_), .B(x1), .C(mai_mai_n17_), .Y(mai_mai_n325_));
  OAI210     m309(.A0(mai_mai_n312_), .A1(mai_mai_n310_), .B0(mai_mai_n325_), .Y(mai_mai_n326_));
  INV        m310(.A(mai_mai_n227_), .Y(mai_mai_n327_));
  NA2        m311(.A(mai_mai_n35_), .B(mai_mai_n41_), .Y(mai_mai_n328_));
  OR2        m312(.A(mai_mai_n328_), .B(mai_mai_n296_), .Y(mai_mai_n329_));
  OAI220     m313(.A0(mai_mai_n329_), .A1(mai_mai_n167_), .B0(mai_mai_n244_), .B1(mai_mai_n327_), .Y(mai_mai_n330_));
  AO210      m314(.A0(mai_mai_n326_), .A1(mai_mai_n154_), .B0(mai_mai_n330_), .Y(mai_mai_n331_));
  NO4        m315(.A(mai_mai_n331_), .B(mai_mai_n324_), .C(mai_mai_n315_), .D(mai_mai_n309_), .Y(mai_mai_n332_));
  OAI210     m316(.A0(mai_mai_n304_), .A1(mai_mai_n256_), .B0(mai_mai_n332_), .Y(mai04));
  OAI210     m317(.A0(x8), .A1(mai_mai_n18_), .B0(x4), .Y(mai_mai_n334_));
  NA3        m318(.A(mai_mai_n334_), .B(mai_mai_n286_), .C(mai_mai_n83_), .Y(mai_mai_n335_));
  NO2        m319(.A(x2), .B(x1), .Y(mai_mai_n336_));
  OAI210     m320(.A0(mai_mai_n267_), .A1(mai_mai_n336_), .B0(mai_mai_n35_), .Y(mai_mai_n337_));
  NO2        m321(.A(mai_mai_n336_), .B(mai_mai_n316_), .Y(mai_mai_n338_));
  AOI210     m322(.A0(mai_mai_n60_), .A1(x4), .B0(mai_mai_n113_), .Y(mai_mai_n339_));
  OAI210     m323(.A0(mai_mai_n339_), .A1(mai_mai_n338_), .B0(mai_mai_n257_), .Y(mai_mai_n340_));
  NO2        m324(.A(mai_mai_n284_), .B(mai_mai_n90_), .Y(mai_mai_n341_));
  NO2        m325(.A(mai_mai_n341_), .B(mai_mai_n35_), .Y(mai_mai_n342_));
  NO2        m326(.A(mai_mai_n314_), .B(mai_mai_n214_), .Y(mai_mai_n343_));
  NA2        m327(.A(mai_mai_n343_), .B(mai_mai_n92_), .Y(mai_mai_n344_));
  NA3        m328(.A(mai_mai_n344_), .B(mai_mai_n342_), .C(mai_mai_n340_), .Y(mai_mai_n345_));
  NA2        m329(.A(mai_mai_n345_), .B(mai_mai_n337_), .Y(mai_mai_n346_));
  NO2        m330(.A(mai_mai_n219_), .B(mai_mai_n114_), .Y(mai_mai_n347_));
  NO3        m331(.A(mai_mai_n264_), .B(mai_mai_n121_), .C(mai_mai_n18_), .Y(mai_mai_n348_));
  NO2        m332(.A(mai_mai_n348_), .B(mai_mai_n347_), .Y(mai_mai_n349_));
  OAI210     m333(.A0(mai_mai_n119_), .A1(mai_mai_n107_), .B0(mai_mai_n183_), .Y(mai_mai_n350_));
  NA3        m334(.A(mai_mai_n350_), .B(x6), .C(x3), .Y(mai_mai_n351_));
  NOi21      m335(.An(mai_mai_n156_), .B(mai_mai_n134_), .Y(mai_mai_n352_));
  AOI210     m336(.A0(x8), .A1(x0), .B0(x1), .Y(mai_mai_n353_));
  OAI220     m337(.A0(mai_mai_n353_), .A1(mai_mai_n328_), .B0(mai_mai_n284_), .B1(mai_mai_n325_), .Y(mai_mai_n354_));
  AOI210     m338(.A0(mai_mai_n352_), .A1(mai_mai_n61_), .B0(mai_mai_n354_), .Y(mai_mai_n355_));
  NA2        m339(.A(x2), .B(mai_mai_n17_), .Y(mai_mai_n356_));
  OAI210     m340(.A0(mai_mai_n107_), .A1(mai_mai_n17_), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  AOI220     m341(.A0(mai_mai_n357_), .A1(mai_mai_n77_), .B0(mai_mai_n341_), .B1(mai_mai_n92_), .Y(mai_mai_n358_));
  NA4        m342(.A(mai_mai_n358_), .B(mai_mai_n355_), .C(mai_mai_n351_), .D(mai_mai_n349_), .Y(mai_mai_n359_));
  OAI210     m343(.A0(mai_mai_n112_), .A1(x3), .B0(mai_mai_n317_), .Y(mai_mai_n360_));
  NA3        m344(.A(mai_mai_n238_), .B(mai_mai_n224_), .C(mai_mai_n82_), .Y(mai_mai_n361_));
  NA3        m345(.A(mai_mai_n361_), .B(mai_mai_n360_), .C(mai_mai_n159_), .Y(mai_mai_n362_));
  AOI210     m346(.A0(mai_mai_n359_), .A1(x4), .B0(mai_mai_n362_), .Y(mai_mai_n363_));
  NA3        m347(.A(mai_mai_n338_), .B(mai_mai_n219_), .C(mai_mai_n92_), .Y(mai_mai_n364_));
  NOi21      m348(.An(x4), .B(x0), .Y(mai_mai_n365_));
  XO2        m349(.A(x4), .B(x0), .Y(mai_mai_n366_));
  OAI210     m350(.A0(mai_mai_n366_), .A1(mai_mai_n118_), .B0(mai_mai_n279_), .Y(mai_mai_n367_));
  AOI220     m351(.A0(mai_mai_n367_), .A1(x8), .B0(mai_mai_n365_), .B1(mai_mai_n93_), .Y(mai_mai_n368_));
  AOI210     m352(.A0(mai_mai_n368_), .A1(mai_mai_n364_), .B0(x3), .Y(mai_mai_n369_));
  INV        m353(.A(mai_mai_n93_), .Y(mai_mai_n370_));
  NO2        m354(.A(mai_mai_n92_), .B(x4), .Y(mai_mai_n371_));
  AOI220     m355(.A0(mai_mai_n371_), .A1(mai_mai_n42_), .B0(mai_mai_n128_), .B1(mai_mai_n370_), .Y(mai_mai_n372_));
  NO3        m356(.A(mai_mai_n366_), .B(mai_mai_n170_), .C(x2), .Y(mai_mai_n373_));
  INV        m357(.A(mai_mai_n373_), .Y(mai_mai_n374_));
  NA4        m358(.A(mai_mai_n374_), .B(mai_mai_n372_), .C(mai_mai_n234_), .D(x6), .Y(mai_mai_n375_));
  OAI220     m359(.A0(mai_mai_n316_), .A1(mai_mai_n90_), .B0(mai_mai_n188_), .B1(mai_mai_n92_), .Y(mai_mai_n376_));
  NO2        m360(.A(mai_mai_n41_), .B(x0), .Y(mai_mai_n377_));
  NA2        m361(.A(mai_mai_n376_), .B(mai_mai_n59_), .Y(mai_mai_n378_));
  NO2        m362(.A(mai_mai_n156_), .B(mai_mai_n79_), .Y(mai_mai_n379_));
  NO2        m363(.A(mai_mai_n34_), .B(x2), .Y(mai_mai_n380_));
  NOi21      m364(.An(mai_mai_n124_), .B(mai_mai_n27_), .Y(mai_mai_n381_));
  AOI210     m365(.A0(mai_mai_n380_), .A1(mai_mai_n379_), .B0(mai_mai_n381_), .Y(mai_mai_n382_));
  OAI210     m366(.A0(mai_mai_n378_), .A1(mai_mai_n60_), .B0(mai_mai_n382_), .Y(mai_mai_n383_));
  OAI220     m367(.A0(mai_mai_n383_), .A1(x6), .B0(mai_mai_n375_), .B1(mai_mai_n369_), .Y(mai_mai_n384_));
  OAI210     m368(.A0(mai_mai_n61_), .A1(mai_mai_n46_), .B0(mai_mai_n40_), .Y(mai_mai_n385_));
  OAI210     m369(.A0(mai_mai_n385_), .A1(mai_mai_n92_), .B0(mai_mai_n329_), .Y(mai_mai_n386_));
  AOI210     m370(.A0(mai_mai_n386_), .A1(mai_mai_n18_), .B0(mai_mai_n159_), .Y(mai_mai_n387_));
  AO220      m371(.A0(mai_mai_n387_), .A1(mai_mai_n384_), .B0(mai_mai_n363_), .B1(mai_mai_n346_), .Y(mai_mai_n388_));
  NA2        m372(.A(mai_mai_n380_), .B(x6), .Y(mai_mai_n389_));
  AOI210     m373(.A0(x6), .A1(x1), .B0(mai_mai_n158_), .Y(mai_mai_n390_));
  NA2        m374(.A(mai_mai_n371_), .B(x0), .Y(mai_mai_n391_));
  NA2        m375(.A(mai_mai_n82_), .B(x6), .Y(mai_mai_n392_));
  OAI210     m376(.A0(mai_mai_n391_), .A1(mai_mai_n390_), .B0(mai_mai_n392_), .Y(mai_mai_n393_));
  AOI220     m377(.A0(mai_mai_n393_), .A1(mai_mai_n389_), .B0(mai_mai_n228_), .B1(mai_mai_n47_), .Y(mai_mai_n394_));
  NA3        m378(.A(mai_mai_n394_), .B(mai_mai_n388_), .C(mai_mai_n335_), .Y(mai_mai_n395_));
  AOI210     m379(.A0(mai_mai_n207_), .A1(x8), .B0(mai_mai_n112_), .Y(mai_mai_n396_));
  NA2        m380(.A(mai_mai_n396_), .B(mai_mai_n356_), .Y(mai_mai_n397_));
  NA3        m381(.A(mai_mai_n397_), .B(mai_mai_n204_), .C(mai_mai_n159_), .Y(mai_mai_n398_));
  OAI210     m382(.A0(mai_mai_n28_), .A1(x1), .B0(mai_mai_n242_), .Y(mai_mai_n399_));
  AO220      m383(.A0(mai_mai_n399_), .A1(mai_mai_n155_), .B0(mai_mai_n111_), .B1(x4), .Y(mai_mai_n400_));
  NA3        m384(.A(x7), .B(x3), .C(x0), .Y(mai_mai_n401_));
  NA2        m385(.A(mai_mai_n233_), .B(x0), .Y(mai_mai_n402_));
  OAI220     m386(.A0(mai_mai_n402_), .A1(mai_mai_n219_), .B0(mai_mai_n401_), .B1(mai_mai_n370_), .Y(mai_mai_n403_));
  AOI210     m387(.A0(mai_mai_n400_), .A1(mai_mai_n120_), .B0(mai_mai_n403_), .Y(mai_mai_n404_));
  AOI210     m388(.A0(mai_mai_n404_), .A1(mai_mai_n398_), .B0(mai_mai_n25_), .Y(mai_mai_n405_));
  NA3        m389(.A(mai_mai_n122_), .B(mai_mai_n233_), .C(x0), .Y(mai_mai_n406_));
  OAI210     m390(.A0(mai_mai_n204_), .A1(mai_mai_n66_), .B0(mai_mai_n214_), .Y(mai_mai_n407_));
  NA3        m391(.A(mai_mai_n207_), .B(mai_mai_n235_), .C(x8), .Y(mai_mai_n408_));
  AOI210     m392(.A0(mai_mai_n408_), .A1(mai_mai_n407_), .B0(mai_mai_n25_), .Y(mai_mai_n409_));
  NA2        m393(.A(mai_mai_n409_), .B(mai_mai_n155_), .Y(mai_mai_n410_));
  NAi31      m394(.An(mai_mai_n48_), .B(mai_mai_n305_), .C(mai_mai_n184_), .Y(mai_mai_n411_));
  NA3        m395(.A(mai_mai_n411_), .B(mai_mai_n410_), .C(mai_mai_n406_), .Y(mai_mai_n412_));
  OAI210     m396(.A0(mai_mai_n412_), .A1(mai_mai_n405_), .B0(x6), .Y(mai_mai_n413_));
  OAI210     m397(.A0(mai_mai_n170_), .A1(mai_mai_n46_), .B0(mai_mai_n139_), .Y(mai_mai_n414_));
  NA3        m398(.A(mai_mai_n53_), .B(mai_mai_n37_), .C(mai_mai_n30_), .Y(mai_mai_n415_));
  AOI220     m399(.A0(mai_mai_n415_), .A1(mai_mai_n414_), .B0(mai_mai_n38_), .B1(mai_mai_n31_), .Y(mai_mai_n416_));
  NO2        m400(.A(mai_mai_n159_), .B(x0), .Y(mai_mai_n417_));
  AOI220     m401(.A0(mai_mai_n417_), .A1(mai_mai_n233_), .B0(mai_mai_n204_), .B1(mai_mai_n159_), .Y(mai_mai_n418_));
  AOI210     m402(.A0(mai_mai_n130_), .A1(mai_mai_n262_), .B0(x1), .Y(mai_mai_n419_));
  OAI210     m403(.A0(mai_mai_n418_), .A1(x8), .B0(mai_mai_n419_), .Y(mai_mai_n420_));
  NAi31      m404(.An(x2), .B(x8), .C(x0), .Y(mai_mai_n421_));
  OAI210     m405(.A0(mai_mai_n421_), .A1(x4), .B0(mai_mai_n171_), .Y(mai_mai_n422_));
  NA3        m406(.A(mai_mai_n422_), .B(mai_mai_n153_), .C(x9), .Y(mai_mai_n423_));
  NO4        m407(.A(mai_mai_n129_), .B(mai_mai_n316_), .C(x9), .D(x2), .Y(mai_mai_n424_));
  NOi21      m408(.An(mai_mai_n127_), .B(mai_mai_n188_), .Y(mai_mai_n425_));
  NO3        m409(.A(mai_mai_n425_), .B(mai_mai_n424_), .C(mai_mai_n18_), .Y(mai_mai_n426_));
  NO3        m410(.A(x9), .B(mai_mai_n159_), .C(x0), .Y(mai_mai_n427_));
  AOI220     m411(.A0(mai_mai_n427_), .A1(mai_mai_n257_), .B0(mai_mai_n379_), .B1(mai_mai_n159_), .Y(mai_mai_n428_));
  NA4        m412(.A(mai_mai_n428_), .B(mai_mai_n426_), .C(mai_mai_n423_), .D(mai_mai_n48_), .Y(mai_mai_n429_));
  OAI210     m413(.A0(mai_mai_n420_), .A1(mai_mai_n416_), .B0(mai_mai_n429_), .Y(mai_mai_n430_));
  NOi31      m414(.An(mai_mai_n417_), .B(mai_mai_n31_), .C(x8), .Y(mai_mai_n431_));
  AOI210     m415(.A0(mai_mai_n37_), .A1(x9), .B0(mai_mai_n137_), .Y(mai_mai_n432_));
  NO3        m416(.A(mai_mai_n432_), .B(mai_mai_n127_), .C(mai_mai_n41_), .Y(mai_mai_n433_));
  NOi31      m417(.An(x1), .B(x8), .C(x7), .Y(mai_mai_n434_));
  AOI220     m418(.A0(mai_mai_n434_), .A1(mai_mai_n365_), .B0(mai_mai_n128_), .B1(x3), .Y(mai_mai_n435_));
  AOI210     m419(.A0(mai_mai_n279_), .A1(mai_mai_n58_), .B0(mai_mai_n126_), .Y(mai_mai_n436_));
  OAI210     m420(.A0(mai_mai_n436_), .A1(x3), .B0(mai_mai_n435_), .Y(mai_mai_n437_));
  NO3        m421(.A(mai_mai_n437_), .B(mai_mai_n433_), .C(x2), .Y(mai_mai_n438_));
  OAI220     m422(.A0(mai_mai_n366_), .A1(mai_mai_n320_), .B0(mai_mai_n316_), .B1(mai_mai_n41_), .Y(mai_mai_n439_));
  AOI210     m423(.A0(x9), .A1(mai_mai_n46_), .B0(mai_mai_n401_), .Y(mai_mai_n440_));
  AOI220     m424(.A0(mai_mai_n440_), .A1(mai_mai_n92_), .B0(mai_mai_n439_), .B1(mai_mai_n159_), .Y(mai_mai_n441_));
  NO2        m425(.A(mai_mai_n441_), .B(mai_mai_n52_), .Y(mai_mai_n442_));
  NO3        m426(.A(mai_mai_n442_), .B(mai_mai_n438_), .C(mai_mai_n431_), .Y(mai_mai_n443_));
  AOI210     m427(.A0(mai_mai_n443_), .A1(mai_mai_n430_), .B0(mai_mai_n25_), .Y(mai_mai_n444_));
  NA4        m428(.A(mai_mai_n30_), .B(mai_mai_n92_), .C(x2), .D(mai_mai_n17_), .Y(mai_mai_n445_));
  NO3        m429(.A(mai_mai_n66_), .B(mai_mai_n18_), .C(x0), .Y(mai_mai_n446_));
  NA2        m430(.A(mai_mai_n446_), .B(mai_mai_n280_), .Y(mai_mai_n447_));
  NO2        m431(.A(mai_mai_n447_), .B(mai_mai_n104_), .Y(mai_mai_n448_));
  NO3        m432(.A(mai_mai_n284_), .B(mai_mai_n183_), .C(mai_mai_n38_), .Y(mai_mai_n449_));
  OAI210     m433(.A0(mai_mai_n449_), .A1(mai_mai_n448_), .B0(x7), .Y(mai_mai_n450_));
  NA2        m434(.A(mai_mai_n238_), .B(x7), .Y(mai_mai_n451_));
  NA3        m435(.A(mai_mai_n451_), .B(mai_mai_n158_), .C(mai_mai_n138_), .Y(mai_mai_n452_));
  NA3        m436(.A(mai_mai_n452_), .B(mai_mai_n450_), .C(mai_mai_n445_), .Y(mai_mai_n453_));
  OAI210     m437(.A0(mai_mai_n453_), .A1(mai_mai_n444_), .B0(mai_mai_n35_), .Y(mai_mai_n454_));
  NO2        m438(.A(mai_mai_n427_), .B(mai_mai_n214_), .Y(mai_mai_n455_));
  NO4        m439(.A(mai_mai_n455_), .B(mai_mai_n76_), .C(x4), .D(mai_mai_n52_), .Y(mai_mai_n456_));
  NA2        m440(.A(mai_mai_n267_), .B(mai_mai_n21_), .Y(mai_mai_n457_));
  NO2        m441(.A(mai_mai_n167_), .B(mai_mai_n139_), .Y(mai_mai_n458_));
  NA2        m442(.A(mai_mai_n458_), .B(mai_mai_n457_), .Y(mai_mai_n459_));
  AOI210     m443(.A0(mai_mai_n459_), .A1(mai_mai_n174_), .B0(mai_mai_n28_), .Y(mai_mai_n460_));
  AOI220     m444(.A0(mai_mai_n377_), .A1(mai_mai_n92_), .B0(mai_mai_n156_), .B1(mai_mai_n207_), .Y(mai_mai_n461_));
  NA3        m445(.A(mai_mai_n461_), .B(mai_mai_n421_), .C(mai_mai_n90_), .Y(mai_mai_n462_));
  NA2        m446(.A(mai_mai_n462_), .B(mai_mai_n184_), .Y(mai_mai_n463_));
  OAI220     m447(.A0(mai_mai_n293_), .A1(mai_mai_n67_), .B0(mai_mai_n167_), .B1(mai_mai_n41_), .Y(mai_mai_n464_));
  NA2        m448(.A(x3), .B(mai_mai_n52_), .Y(mai_mai_n465_));
  OAI210     m449(.A0(mai_mai_n155_), .A1(mai_mai_n18_), .B0(mai_mai_n21_), .Y(mai_mai_n466_));
  NO3        m450(.A(mai_mai_n434_), .B(x3), .C(mai_mai_n52_), .Y(mai_mai_n467_));
  NA2        m451(.A(mai_mai_n467_), .B(mai_mai_n466_), .Y(mai_mai_n468_));
  OAI210     m452(.A0(mai_mai_n160_), .A1(mai_mai_n465_), .B0(mai_mai_n468_), .Y(mai_mai_n469_));
  AOI220     m453(.A0(mai_mai_n469_), .A1(x0), .B0(mai_mai_n464_), .B1(mai_mai_n139_), .Y(mai_mai_n470_));
  AOI210     m454(.A0(mai_mai_n470_), .A1(mai_mai_n463_), .B0(mai_mai_n244_), .Y(mai_mai_n471_));
  NA2        m455(.A(x9), .B(x5), .Y(mai_mai_n472_));
  NO4        m456(.A(mai_mai_n107_), .B(mai_mai_n472_), .C(mai_mai_n58_), .D(mai_mai_n31_), .Y(mai_mai_n473_));
  NO4        m457(.A(mai_mai_n473_), .B(mai_mai_n471_), .C(mai_mai_n460_), .D(mai_mai_n456_), .Y(mai_mai_n474_));
  NA3        m458(.A(mai_mai_n474_), .B(mai_mai_n454_), .C(mai_mai_n413_), .Y(mai_mai_n475_));
  AOI210     m459(.A0(mai_mai_n395_), .A1(mai_mai_n25_), .B0(mai_mai_n475_), .Y(mai05));
  INV        u000(.A(x0), .Y(men_men_n17_));
  INV        u001(.A(x1), .Y(men_men_n18_));
  NO2        u002(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n19_));
  NO2        u003(.A(x6), .B(x5), .Y(men_men_n20_));
  OR2        u004(.A(x8), .B(x7), .Y(men_men_n21_));
  NOi21      u005(.An(men_men_n20_), .B(men_men_n21_), .Y(men_men_n22_));
  NAi21      u006(.An(men_men_n22_), .B(men_men_n19_), .Y(men_men_n23_));
  NA2        u007(.A(men_men_n18_), .B(men_men_n17_), .Y(men_men_n24_));
  INV        u008(.A(x5), .Y(men_men_n25_));
  NA2        u009(.A(x7), .B(x6), .Y(men_men_n26_));
  NA2        u010(.A(x8), .B(x3), .Y(men_men_n27_));
  NA2        u011(.A(x4), .B(x2), .Y(men_men_n28_));
  NO4        u012(.A(men_men_n28_), .B(men_men_n27_), .C(men_men_n26_), .D(men_men_n25_), .Y(men_men_n29_));
  NO2        u013(.A(men_men_n29_), .B(men_men_n24_), .Y(men_men_n30_));
  NO2        u014(.A(x4), .B(x3), .Y(men_men_n31_));
  INV        u015(.A(men_men_n31_), .Y(men_men_n32_));
  OA210      u016(.A0(men_men_n32_), .A1(x2), .B0(men_men_n19_), .Y(men_men_n33_));
  NOi31      u017(.An(men_men_n23_), .B(men_men_n33_), .C(men_men_n30_), .Y(men00));
  NO2        u018(.A(x1), .B(x0), .Y(men_men_n35_));
  INV        u019(.A(x6), .Y(men_men_n36_));
  NO2        u020(.A(men_men_n36_), .B(men_men_n25_), .Y(men_men_n37_));
  AN2        u021(.A(x8), .B(x7), .Y(men_men_n38_));
  NA3        u022(.A(men_men_n38_), .B(men_men_n37_), .C(men_men_n35_), .Y(men_men_n39_));
  NA2        u023(.A(x4), .B(x3), .Y(men_men_n40_));
  AOI210     u024(.A0(men_men_n39_), .A1(men_men_n23_), .B0(men_men_n40_), .Y(men_men_n41_));
  NO2        u025(.A(x2), .B(x0), .Y(men_men_n42_));
  INV        u026(.A(x3), .Y(men_men_n43_));
  NO2        u027(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n44_));
  INV        u028(.A(men_men_n44_), .Y(men_men_n45_));
  NO2        u029(.A(men_men_n37_), .B(x4), .Y(men_men_n46_));
  OAI210     u030(.A0(men_men_n46_), .A1(men_men_n45_), .B0(men_men_n42_), .Y(men_men_n47_));
  INV        u031(.A(x4), .Y(men_men_n48_));
  NO2        u032(.A(men_men_n48_), .B(men_men_n17_), .Y(men_men_n49_));
  NA2        u033(.A(men_men_n49_), .B(x2), .Y(men_men_n50_));
  OAI210     u034(.A0(men_men_n50_), .A1(men_men_n20_), .B0(men_men_n47_), .Y(men_men_n51_));
  NA2        u035(.A(men_men_n38_), .B(men_men_n37_), .Y(men_men_n52_));
  AOI220     u036(.A0(men_men_n52_), .A1(men_men_n35_), .B0(men_men_n22_), .B1(men_men_n19_), .Y(men_men_n53_));
  INV        u037(.A(x2), .Y(men_men_n54_));
  NO2        u038(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n55_));
  NA2        u039(.A(men_men_n43_), .B(men_men_n18_), .Y(men_men_n56_));
  NA2        u040(.A(men_men_n56_), .B(men_men_n55_), .Y(men_men_n57_));
  OAI210     u041(.A0(men_men_n53_), .A1(men_men_n32_), .B0(men_men_n57_), .Y(men_men_n58_));
  NO3        u042(.A(men_men_n58_), .B(men_men_n51_), .C(men_men_n41_), .Y(men01));
  NA2        u043(.A(x8), .B(x7), .Y(men_men_n60_));
  NA2        u044(.A(men_men_n43_), .B(x1), .Y(men_men_n61_));
  INV        u045(.A(x9), .Y(men_men_n62_));
  NO2        u046(.A(men_men_n62_), .B(men_men_n36_), .Y(men_men_n63_));
  INV        u047(.A(men_men_n63_), .Y(men_men_n64_));
  NO2        u048(.A(x7), .B(x6), .Y(men_men_n65_));
  NO2        u049(.A(men_men_n61_), .B(x5), .Y(men_men_n66_));
  NO2        u050(.A(x8), .B(x2), .Y(men_men_n67_));
  INV        u051(.A(men_men_n67_), .Y(men_men_n68_));
  NO2        u052(.A(men_men_n68_), .B(x1), .Y(men_men_n69_));
  OA210      u053(.A0(men_men_n69_), .A1(men_men_n66_), .B0(men_men_n65_), .Y(men_men_n70_));
  OAI210     u054(.A0(men_men_n44_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n71_));
  OAI210     u055(.A0(men_men_n56_), .A1(men_men_n20_), .B0(men_men_n71_), .Y(men_men_n72_));
  NAi31      u056(.An(x1), .B(x9), .C(x5), .Y(men_men_n73_));
  OAI220     u057(.A0(men_men_n73_), .A1(men_men_n43_), .B0(men_men_n72_), .B1(men_men_n70_), .Y(men_men_n74_));
  NA2        u058(.A(men_men_n74_), .B(x4), .Y(men_men_n75_));
  NA2        u059(.A(men_men_n48_), .B(x2), .Y(men_men_n76_));
  OAI210     u060(.A0(men_men_n76_), .A1(men_men_n56_), .B0(x0), .Y(men_men_n77_));
  NA2        u061(.A(x5), .B(x3), .Y(men_men_n78_));
  NO2        u062(.A(x8), .B(x6), .Y(men_men_n79_));
  NO4        u063(.A(men_men_n79_), .B(men_men_n78_), .C(men_men_n65_), .D(men_men_n54_), .Y(men_men_n80_));
  NAi21      u064(.An(x4), .B(x3), .Y(men_men_n81_));
  INV        u065(.A(men_men_n81_), .Y(men_men_n82_));
  NO2        u066(.A(men_men_n82_), .B(men_men_n22_), .Y(men_men_n83_));
  NO2        u067(.A(x4), .B(x2), .Y(men_men_n84_));
  NO2        u068(.A(men_men_n84_), .B(x3), .Y(men_men_n85_));
  NO3        u069(.A(men_men_n85_), .B(men_men_n83_), .C(men_men_n18_), .Y(men_men_n86_));
  NO3        u070(.A(men_men_n86_), .B(men_men_n80_), .C(men_men_n77_), .Y(men_men_n87_));
  NO4        u071(.A(men_men_n21_), .B(x6), .C(men_men_n43_), .D(x1), .Y(men_men_n88_));
  NA2        u072(.A(men_men_n62_), .B(men_men_n48_), .Y(men_men_n89_));
  NA2        u073(.A(men_men_n88_), .B(men_men_n48_), .Y(men_men_n90_));
  NA2        u074(.A(x3), .B(men_men_n18_), .Y(men_men_n91_));
  NO2        u075(.A(men_men_n91_), .B(men_men_n25_), .Y(men_men_n92_));
  INV        u076(.A(x8), .Y(men_men_n93_));
  NA2        u077(.A(x2), .B(x1), .Y(men_men_n94_));
  INV        u078(.A(men_men_n92_), .Y(men_men_n95_));
  NO2        u079(.A(men_men_n95_), .B(men_men_n26_), .Y(men_men_n96_));
  AOI210     u080(.A0(men_men_n56_), .A1(men_men_n25_), .B0(men_men_n54_), .Y(men_men_n97_));
  OAI210     u081(.A0(men_men_n45_), .A1(men_men_n37_), .B0(men_men_n48_), .Y(men_men_n98_));
  NO3        u082(.A(men_men_n98_), .B(men_men_n97_), .C(men_men_n96_), .Y(men_men_n99_));
  NA2        u083(.A(x4), .B(men_men_n43_), .Y(men_men_n100_));
  NO2        u084(.A(men_men_n48_), .B(men_men_n54_), .Y(men_men_n101_));
  OAI210     u085(.A0(men_men_n101_), .A1(men_men_n43_), .B0(men_men_n18_), .Y(men_men_n102_));
  AOI210     u086(.A0(men_men_n100_), .A1(men_men_n52_), .B0(men_men_n102_), .Y(men_men_n103_));
  NO2        u087(.A(x3), .B(x2), .Y(men_men_n104_));
  NA3        u088(.A(men_men_n104_), .B(men_men_n26_), .C(men_men_n25_), .Y(men_men_n105_));
  AOI210     u089(.A0(x8), .A1(x6), .B0(men_men_n105_), .Y(men_men_n106_));
  NA2        u090(.A(men_men_n54_), .B(x1), .Y(men_men_n107_));
  OAI210     u091(.A0(men_men_n107_), .A1(men_men_n40_), .B0(men_men_n17_), .Y(men_men_n108_));
  NO4        u092(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n103_), .D(men_men_n99_), .Y(men_men_n109_));
  AO220      u093(.A0(men_men_n109_), .A1(men_men_n90_), .B0(men_men_n87_), .B1(men_men_n75_), .Y(men02));
  NO2        u094(.A(x3), .B(men_men_n54_), .Y(men_men_n111_));
  NO2        u095(.A(x8), .B(men_men_n18_), .Y(men_men_n112_));
  NA2        u096(.A(men_men_n54_), .B(men_men_n17_), .Y(men_men_n113_));
  NA2        u097(.A(men_men_n43_), .B(x0), .Y(men_men_n114_));
  OAI210     u098(.A0(men_men_n89_), .A1(men_men_n113_), .B0(men_men_n114_), .Y(men_men_n115_));
  AOI220     u099(.A0(men_men_n115_), .A1(men_men_n112_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n116_));
  NO3        u100(.A(men_men_n116_), .B(x7), .C(x5), .Y(men_men_n117_));
  NA2        u101(.A(x9), .B(x2), .Y(men_men_n118_));
  OR2        u102(.A(x8), .B(x0), .Y(men_men_n119_));
  INV        u103(.A(men_men_n119_), .Y(men_men_n120_));
  NAi21      u104(.An(x2), .B(x8), .Y(men_men_n121_));
  INV        u105(.A(men_men_n121_), .Y(men_men_n122_));
  NO2        u106(.A(men_men_n122_), .B(men_men_n120_), .Y(men_men_n123_));
  NO2        u107(.A(x4), .B(x1), .Y(men_men_n124_));
  NA3        u108(.A(men_men_n124_), .B(men_men_n123_), .C(men_men_n60_), .Y(men_men_n125_));
  NOi21      u109(.An(x0), .B(x1), .Y(men_men_n126_));
  NO3        u110(.A(x9), .B(x8), .C(x7), .Y(men_men_n127_));
  NOi21      u111(.An(x0), .B(x4), .Y(men_men_n128_));
  NO2        u112(.A(men_men_n125_), .B(men_men_n78_), .Y(men_men_n129_));
  NO2        u113(.A(x5), .B(men_men_n48_), .Y(men_men_n130_));
  NA2        u114(.A(x2), .B(men_men_n18_), .Y(men_men_n131_));
  AOI210     u115(.A0(men_men_n131_), .A1(men_men_n107_), .B0(men_men_n114_), .Y(men_men_n132_));
  OAI210     u116(.A0(men_men_n132_), .A1(men_men_n35_), .B0(men_men_n130_), .Y(men_men_n133_));
  NAi21      u117(.An(x0), .B(x4), .Y(men_men_n134_));
  NO2        u118(.A(men_men_n134_), .B(x1), .Y(men_men_n135_));
  NO2        u119(.A(x7), .B(x0), .Y(men_men_n136_));
  NO2        u120(.A(men_men_n84_), .B(men_men_n101_), .Y(men_men_n137_));
  NO2        u121(.A(men_men_n137_), .B(x3), .Y(men_men_n138_));
  OAI210     u122(.A0(men_men_n136_), .A1(men_men_n135_), .B0(men_men_n138_), .Y(men_men_n139_));
  NO2        u123(.A(men_men_n21_), .B(men_men_n43_), .Y(men_men_n140_));
  NA2        u124(.A(x5), .B(x0), .Y(men_men_n141_));
  NO2        u125(.A(men_men_n48_), .B(x2), .Y(men_men_n142_));
  NA3        u126(.A(men_men_n142_), .B(men_men_n141_), .C(men_men_n140_), .Y(men_men_n143_));
  NA4        u127(.A(men_men_n143_), .B(men_men_n139_), .C(men_men_n133_), .D(men_men_n36_), .Y(men_men_n144_));
  NO3        u128(.A(men_men_n144_), .B(men_men_n129_), .C(men_men_n117_), .Y(men_men_n145_));
  NO3        u129(.A(men_men_n78_), .B(men_men_n76_), .C(men_men_n24_), .Y(men_men_n146_));
  NO2        u130(.A(men_men_n28_), .B(men_men_n25_), .Y(men_men_n147_));
  NA2        u131(.A(x7), .B(x3), .Y(men_men_n148_));
  NO2        u132(.A(men_men_n100_), .B(x5), .Y(men_men_n149_));
  NO2        u133(.A(x9), .B(x7), .Y(men_men_n150_));
  NOi21      u134(.An(x8), .B(x0), .Y(men_men_n151_));
  OA210      u135(.A0(men_men_n150_), .A1(x1), .B0(men_men_n151_), .Y(men_men_n152_));
  NO2        u136(.A(men_men_n43_), .B(x2), .Y(men_men_n153_));
  INV        u137(.A(x7), .Y(men_men_n154_));
  NA2        u138(.A(men_men_n154_), .B(men_men_n18_), .Y(men_men_n155_));
  AOI220     u139(.A0(men_men_n155_), .A1(men_men_n153_), .B0(men_men_n111_), .B1(men_men_n38_), .Y(men_men_n156_));
  NO2        u140(.A(men_men_n25_), .B(x4), .Y(men_men_n157_));
  NO2        u141(.A(men_men_n157_), .B(men_men_n128_), .Y(men_men_n158_));
  NO2        u142(.A(men_men_n158_), .B(men_men_n156_), .Y(men_men_n159_));
  AOI210     u143(.A0(men_men_n152_), .A1(men_men_n149_), .B0(men_men_n159_), .Y(men_men_n160_));
  OAI210     u144(.A0(men_men_n148_), .A1(men_men_n50_), .B0(men_men_n160_), .Y(men_men_n161_));
  NA2        u145(.A(x5), .B(x1), .Y(men_men_n162_));
  INV        u146(.A(men_men_n162_), .Y(men_men_n163_));
  AOI210     u147(.A0(men_men_n163_), .A1(men_men_n128_), .B0(men_men_n36_), .Y(men_men_n164_));
  NO2        u148(.A(men_men_n62_), .B(men_men_n93_), .Y(men_men_n165_));
  NAi21      u149(.An(x2), .B(x7), .Y(men_men_n166_));
  NO2        u150(.A(men_men_n166_), .B(men_men_n48_), .Y(men_men_n167_));
  NA2        u151(.A(men_men_n167_), .B(men_men_n66_), .Y(men_men_n168_));
  NAi31      u152(.An(men_men_n78_), .B(men_men_n38_), .C(men_men_n35_), .Y(men_men_n169_));
  NA3        u153(.A(men_men_n169_), .B(men_men_n168_), .C(men_men_n164_), .Y(men_men_n170_));
  NO3        u154(.A(men_men_n170_), .B(men_men_n161_), .C(men_men_n146_), .Y(men_men_n171_));
  NO2        u155(.A(men_men_n171_), .B(men_men_n145_), .Y(men_men_n172_));
  NO2        u156(.A(men_men_n141_), .B(men_men_n137_), .Y(men_men_n173_));
  NA2        u157(.A(men_men_n25_), .B(men_men_n18_), .Y(men_men_n174_));
  NA2        u158(.A(men_men_n25_), .B(men_men_n17_), .Y(men_men_n175_));
  NA3        u159(.A(men_men_n175_), .B(men_men_n174_), .C(men_men_n24_), .Y(men_men_n176_));
  AN2        u160(.A(men_men_n176_), .B(men_men_n142_), .Y(men_men_n177_));
  NA2        u161(.A(x8), .B(x0), .Y(men_men_n178_));
  NO2        u162(.A(men_men_n154_), .B(men_men_n25_), .Y(men_men_n179_));
  NO2        u163(.A(men_men_n126_), .B(x4), .Y(men_men_n180_));
  NA2        u164(.A(men_men_n180_), .B(men_men_n179_), .Y(men_men_n181_));
  AOI210     u165(.A0(men_men_n178_), .A1(men_men_n131_), .B0(men_men_n181_), .Y(men_men_n182_));
  NA2        u166(.A(x2), .B(x0), .Y(men_men_n183_));
  NA2        u167(.A(x4), .B(x1), .Y(men_men_n184_));
  NAi21      u168(.An(men_men_n124_), .B(men_men_n184_), .Y(men_men_n185_));
  NOi31      u169(.An(men_men_n185_), .B(men_men_n157_), .C(men_men_n183_), .Y(men_men_n186_));
  NO4        u170(.A(men_men_n186_), .B(men_men_n182_), .C(men_men_n177_), .D(men_men_n173_), .Y(men_men_n187_));
  NO2        u171(.A(men_men_n187_), .B(men_men_n43_), .Y(men_men_n188_));
  NO2        u172(.A(men_men_n176_), .B(men_men_n76_), .Y(men_men_n189_));
  INV        u173(.A(men_men_n130_), .Y(men_men_n190_));
  NO2        u174(.A(men_men_n107_), .B(men_men_n17_), .Y(men_men_n191_));
  AOI210     u175(.A0(men_men_n35_), .A1(men_men_n93_), .B0(men_men_n191_), .Y(men_men_n192_));
  NO3        u176(.A(men_men_n192_), .B(men_men_n190_), .C(x7), .Y(men_men_n193_));
  NA3        u177(.A(men_men_n185_), .B(men_men_n190_), .C(men_men_n42_), .Y(men_men_n194_));
  OAI210     u178(.A0(men_men_n175_), .A1(men_men_n137_), .B0(men_men_n194_), .Y(men_men_n195_));
  NO3        u179(.A(men_men_n195_), .B(men_men_n193_), .C(men_men_n189_), .Y(men_men_n196_));
  NO2        u180(.A(men_men_n196_), .B(x3), .Y(men_men_n197_));
  NO3        u181(.A(men_men_n197_), .B(men_men_n188_), .C(men_men_n172_), .Y(men03));
  NO2        u182(.A(men_men_n48_), .B(x3), .Y(men_men_n199_));
  NO2        u183(.A(x6), .B(men_men_n25_), .Y(men_men_n200_));
  NO2        u184(.A(men_men_n54_), .B(x1), .Y(men_men_n201_));
  NO2        u185(.A(men_men_n78_), .B(x6), .Y(men_men_n202_));
  NA2        u186(.A(x6), .B(men_men_n25_), .Y(men_men_n203_));
  NO2        u187(.A(men_men_n203_), .B(x4), .Y(men_men_n204_));
  NO2        u188(.A(men_men_n18_), .B(x0), .Y(men_men_n205_));
  AO220      u189(.A0(men_men_n205_), .A1(men_men_n204_), .B0(men_men_n202_), .B1(men_men_n55_), .Y(men_men_n206_));
  INV        u190(.A(men_men_n206_), .Y(men_men_n207_));
  NA2        u191(.A(x3), .B(men_men_n17_), .Y(men_men_n208_));
  NA2        u192(.A(x9), .B(men_men_n54_), .Y(men_men_n209_));
  NA2        u193(.A(men_men_n203_), .B(men_men_n81_), .Y(men_men_n210_));
  AOI210     u194(.A0(men_men_n25_), .A1(x3), .B0(men_men_n183_), .Y(men_men_n211_));
  NA2        u195(.A(men_men_n211_), .B(men_men_n210_), .Y(men_men_n212_));
  NO3        u196(.A(x6), .B(men_men_n18_), .C(x0), .Y(men_men_n213_));
  NO2        u197(.A(x5), .B(x1), .Y(men_men_n214_));
  AOI220     u198(.A0(men_men_n214_), .A1(men_men_n17_), .B0(men_men_n104_), .B1(x5), .Y(men_men_n215_));
  NO2        u199(.A(men_men_n208_), .B(men_men_n174_), .Y(men_men_n216_));
  NO3        u200(.A(x3), .B(x2), .C(x1), .Y(men_men_n217_));
  NO2        u201(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n218_));
  OAI210     u202(.A0(men_men_n215_), .A1(men_men_n64_), .B0(men_men_n218_), .Y(men_men_n219_));
  AOI220     u203(.A0(men_men_n219_), .A1(men_men_n48_), .B0(men_men_n213_), .B1(men_men_n130_), .Y(men_men_n220_));
  NA3        u204(.A(men_men_n220_), .B(men_men_n212_), .C(men_men_n207_), .Y(men_men_n221_));
  NO2        u205(.A(men_men_n48_), .B(men_men_n43_), .Y(men_men_n222_));
  NA2        u206(.A(men_men_n222_), .B(men_men_n19_), .Y(men_men_n223_));
  NO2        u207(.A(x3), .B(men_men_n17_), .Y(men_men_n224_));
  NO2        u208(.A(men_men_n224_), .B(x6), .Y(men_men_n225_));
  NOi21      u209(.An(men_men_n84_), .B(men_men_n225_), .Y(men_men_n226_));
  NA2        u210(.A(men_men_n62_), .B(men_men_n93_), .Y(men_men_n227_));
  NA3        u211(.A(men_men_n227_), .B(men_men_n224_), .C(x6), .Y(men_men_n228_));
  AOI210     u212(.A0(men_men_n228_), .A1(men_men_n226_), .B0(men_men_n154_), .Y(men_men_n229_));
  AO210      u213(.A0(men_men_n229_), .A1(men_men_n223_), .B0(men_men_n179_), .Y(men_men_n230_));
  NA2        u214(.A(men_men_n43_), .B(men_men_n54_), .Y(men_men_n231_));
  OAI210     u215(.A0(men_men_n231_), .A1(men_men_n25_), .B0(men_men_n175_), .Y(men_men_n232_));
  NO3        u216(.A(men_men_n184_), .B(men_men_n62_), .C(x6), .Y(men_men_n233_));
  AOI220     u217(.A0(men_men_n233_), .A1(men_men_n232_), .B0(men_men_n142_), .B1(men_men_n92_), .Y(men_men_n234_));
  NA2        u218(.A(x6), .B(men_men_n48_), .Y(men_men_n235_));
  OAI210     u219(.A0(men_men_n120_), .A1(men_men_n79_), .B0(x4), .Y(men_men_n236_));
  AOI210     u220(.A0(men_men_n236_), .A1(men_men_n235_), .B0(men_men_n78_), .Y(men_men_n237_));
  NA2        u221(.A(men_men_n200_), .B(men_men_n135_), .Y(men_men_n238_));
  NA3        u222(.A(men_men_n208_), .B(men_men_n130_), .C(x6), .Y(men_men_n239_));
  OAI210     u223(.A0(men_men_n93_), .A1(men_men_n36_), .B0(men_men_n66_), .Y(men_men_n240_));
  NA3        u224(.A(men_men_n240_), .B(men_men_n239_), .C(men_men_n238_), .Y(men_men_n241_));
  OAI210     u225(.A0(men_men_n241_), .A1(men_men_n237_), .B0(x2), .Y(men_men_n242_));
  NA3        u226(.A(men_men_n242_), .B(men_men_n234_), .C(men_men_n230_), .Y(men_men_n243_));
  AOI210     u227(.A0(men_men_n221_), .A1(x8), .B0(men_men_n243_), .Y(men_men_n244_));
  NO2        u228(.A(men_men_n93_), .B(x3), .Y(men_men_n245_));
  NA2        u229(.A(men_men_n245_), .B(men_men_n204_), .Y(men_men_n246_));
  NO3        u230(.A(men_men_n91_), .B(men_men_n79_), .C(men_men_n25_), .Y(men_men_n247_));
  AOI210     u231(.A0(men_men_n225_), .A1(men_men_n157_), .B0(men_men_n247_), .Y(men_men_n248_));
  AOI210     u232(.A0(men_men_n248_), .A1(men_men_n246_), .B0(x2), .Y(men_men_n249_));
  NO2        u233(.A(x4), .B(men_men_n54_), .Y(men_men_n250_));
  AOI220     u234(.A0(men_men_n204_), .A1(men_men_n191_), .B0(men_men_n250_), .B1(men_men_n66_), .Y(men_men_n251_));
  NA2        u235(.A(men_men_n62_), .B(x6), .Y(men_men_n252_));
  NA3        u236(.A(men_men_n25_), .B(x3), .C(x2), .Y(men_men_n253_));
  AOI210     u237(.A0(men_men_n253_), .A1(men_men_n141_), .B0(men_men_n252_), .Y(men_men_n254_));
  NA2        u238(.A(men_men_n43_), .B(men_men_n17_), .Y(men_men_n255_));
  NO2        u239(.A(men_men_n255_), .B(men_men_n25_), .Y(men_men_n256_));
  OAI210     u240(.A0(men_men_n256_), .A1(men_men_n254_), .B0(men_men_n124_), .Y(men_men_n257_));
  NA2        u241(.A(men_men_n208_), .B(x6), .Y(men_men_n258_));
  NO2        u242(.A(men_men_n208_), .B(x6), .Y(men_men_n259_));
  NAi21      u243(.An(men_men_n165_), .B(men_men_n259_), .Y(men_men_n260_));
  NA3        u244(.A(men_men_n260_), .B(men_men_n258_), .C(men_men_n147_), .Y(men_men_n261_));
  NA4        u245(.A(men_men_n261_), .B(men_men_n257_), .C(men_men_n251_), .D(men_men_n154_), .Y(men_men_n262_));
  NO2        u246(.A(x9), .B(x6), .Y(men_men_n263_));
  NO2        u247(.A(men_men_n141_), .B(men_men_n18_), .Y(men_men_n264_));
  NAi21      u248(.An(men_men_n264_), .B(men_men_n253_), .Y(men_men_n265_));
  NAi21      u249(.An(x1), .B(x4), .Y(men_men_n266_));
  AOI210     u250(.A0(x3), .A1(x2), .B0(men_men_n48_), .Y(men_men_n267_));
  OAI210     u251(.A0(men_men_n141_), .A1(x3), .B0(men_men_n267_), .Y(men_men_n268_));
  AOI220     u252(.A0(men_men_n268_), .A1(men_men_n266_), .B0(men_men_n265_), .B1(men_men_n263_), .Y(men_men_n269_));
  INV        u253(.A(men_men_n269_), .Y(men_men_n270_));
  NA2        u254(.A(men_men_n62_), .B(x2), .Y(men_men_n271_));
  NO3        u255(.A(x9), .B(x6), .C(x0), .Y(men_men_n272_));
  NA2        u256(.A(men_men_n107_), .B(men_men_n25_), .Y(men_men_n273_));
  NA2        u257(.A(x6), .B(x2), .Y(men_men_n274_));
  NO2        u258(.A(men_men_n274_), .B(men_men_n174_), .Y(men_men_n275_));
  AOI210     u259(.A0(men_men_n273_), .A1(men_men_n272_), .B0(men_men_n275_), .Y(men_men_n276_));
  OAI220     u260(.A0(men_men_n276_), .A1(men_men_n43_), .B0(men_men_n180_), .B1(men_men_n46_), .Y(men_men_n277_));
  NA2        u261(.A(men_men_n277_), .B(men_men_n270_), .Y(men_men_n278_));
  NA2        u262(.A(x9), .B(men_men_n43_), .Y(men_men_n279_));
  NO2        u263(.A(men_men_n279_), .B(men_men_n203_), .Y(men_men_n280_));
  OR3        u264(.A(men_men_n280_), .B(men_men_n202_), .C(men_men_n149_), .Y(men_men_n281_));
  NA2        u265(.A(x4), .B(x0), .Y(men_men_n282_));
  NO3        u266(.A(men_men_n73_), .B(men_men_n282_), .C(x6), .Y(men_men_n283_));
  AOI210     u267(.A0(men_men_n281_), .A1(men_men_n42_), .B0(men_men_n283_), .Y(men_men_n284_));
  AOI210     u268(.A0(men_men_n284_), .A1(men_men_n278_), .B0(x8), .Y(men_men_n285_));
  INV        u269(.A(men_men_n252_), .Y(men_men_n286_));
  OAI210     u270(.A0(men_men_n264_), .A1(men_men_n214_), .B0(men_men_n286_), .Y(men_men_n287_));
  INV        u271(.A(men_men_n178_), .Y(men_men_n288_));
  OAI210     u272(.A0(men_men_n288_), .A1(x4), .B0(men_men_n20_), .Y(men_men_n289_));
  AOI210     u273(.A0(men_men_n289_), .A1(men_men_n287_), .B0(men_men_n231_), .Y(men_men_n290_));
  NO4        u274(.A(men_men_n290_), .B(men_men_n285_), .C(men_men_n262_), .D(men_men_n249_), .Y(men_men_n291_));
  NO2        u275(.A(men_men_n165_), .B(x1), .Y(men_men_n292_));
  NO3        u276(.A(men_men_n292_), .B(x3), .C(men_men_n36_), .Y(men_men_n293_));
  OAI210     u277(.A0(men_men_n293_), .A1(men_men_n259_), .B0(x2), .Y(men_men_n294_));
  OAI210     u278(.A0(men_men_n288_), .A1(x6), .B0(men_men_n44_), .Y(men_men_n295_));
  AOI210     u279(.A0(men_men_n295_), .A1(men_men_n294_), .B0(men_men_n190_), .Y(men_men_n296_));
  NOi21      u280(.An(men_men_n274_), .B(men_men_n17_), .Y(men_men_n297_));
  NA3        u281(.A(men_men_n297_), .B(men_men_n214_), .C(men_men_n40_), .Y(men_men_n298_));
  AOI210     u282(.A0(men_men_n36_), .A1(men_men_n54_), .B0(x0), .Y(men_men_n299_));
  NA3        u283(.A(men_men_n299_), .B(men_men_n163_), .C(men_men_n32_), .Y(men_men_n300_));
  NA2        u284(.A(x3), .B(x2), .Y(men_men_n301_));
  AOI220     u285(.A0(men_men_n301_), .A1(men_men_n231_), .B0(men_men_n300_), .B1(men_men_n298_), .Y(men_men_n302_));
  NAi21      u286(.An(x4), .B(x0), .Y(men_men_n303_));
  NO3        u287(.A(men_men_n303_), .B(men_men_n44_), .C(x2), .Y(men_men_n304_));
  OAI210     u288(.A0(x6), .A1(men_men_n18_), .B0(men_men_n304_), .Y(men_men_n305_));
  OAI220     u289(.A0(men_men_n24_), .A1(x8), .B0(x6), .B1(x1), .Y(men_men_n306_));
  NO2        u290(.A(x9), .B(x8), .Y(men_men_n307_));
  NO2        u291(.A(men_men_n299_), .B(men_men_n297_), .Y(men_men_n308_));
  AOI220     u292(.A0(men_men_n308_), .A1(men_men_n82_), .B0(men_men_n306_), .B1(men_men_n31_), .Y(men_men_n309_));
  AOI210     u293(.A0(men_men_n309_), .A1(men_men_n305_), .B0(men_men_n25_), .Y(men_men_n310_));
  NA3        u294(.A(men_men_n36_), .B(x1), .C(men_men_n17_), .Y(men_men_n311_));
  OAI210     u295(.A0(men_men_n299_), .A1(men_men_n297_), .B0(men_men_n311_), .Y(men_men_n312_));
  INV        u296(.A(men_men_n216_), .Y(men_men_n313_));
  NA2        u297(.A(men_men_n36_), .B(men_men_n43_), .Y(men_men_n314_));
  OR2        u298(.A(men_men_n314_), .B(men_men_n282_), .Y(men_men_n315_));
  OAI220     u299(.A0(men_men_n315_), .A1(men_men_n162_), .B0(men_men_n235_), .B1(men_men_n313_), .Y(men_men_n316_));
  AO210      u300(.A0(men_men_n312_), .A1(men_men_n149_), .B0(men_men_n316_), .Y(men_men_n317_));
  NO4        u301(.A(men_men_n317_), .B(men_men_n310_), .C(men_men_n302_), .D(men_men_n296_), .Y(men_men_n318_));
  OAI210     u302(.A0(men_men_n291_), .A1(men_men_n244_), .B0(men_men_n318_), .Y(men04));
  OAI210     u303(.A0(x8), .A1(men_men_n18_), .B0(x4), .Y(men_men_n320_));
  NA3        u304(.A(men_men_n320_), .B(men_men_n272_), .C(men_men_n85_), .Y(men_men_n321_));
  NO2        u305(.A(x2), .B(x1), .Y(men_men_n322_));
  OAI210     u306(.A0(men_men_n255_), .A1(men_men_n322_), .B0(men_men_n36_), .Y(men_men_n323_));
  NO2        u307(.A(men_men_n322_), .B(men_men_n303_), .Y(men_men_n324_));
  AOI210     u308(.A0(men_men_n62_), .A1(x4), .B0(men_men_n113_), .Y(men_men_n325_));
  OAI210     u309(.A0(men_men_n325_), .A1(men_men_n324_), .B0(men_men_n245_), .Y(men_men_n326_));
  NO2        u310(.A(men_men_n271_), .B(men_men_n91_), .Y(men_men_n327_));
  NO2        u311(.A(men_men_n327_), .B(men_men_n36_), .Y(men_men_n328_));
  NO2        u312(.A(men_men_n301_), .B(men_men_n205_), .Y(men_men_n329_));
  NA2        u313(.A(x9), .B(x0), .Y(men_men_n330_));
  AOI210     u314(.A0(men_men_n91_), .A1(men_men_n76_), .B0(men_men_n330_), .Y(men_men_n331_));
  OAI210     u315(.A0(men_men_n331_), .A1(men_men_n329_), .B0(men_men_n93_), .Y(men_men_n332_));
  NA3        u316(.A(men_men_n332_), .B(men_men_n328_), .C(men_men_n326_), .Y(men_men_n333_));
  NA2        u317(.A(men_men_n333_), .B(men_men_n323_), .Y(men_men_n334_));
  NO2        u318(.A(men_men_n209_), .B(men_men_n114_), .Y(men_men_n335_));
  NO3        u319(.A(men_men_n252_), .B(men_men_n121_), .C(men_men_n18_), .Y(men_men_n336_));
  NO2        u320(.A(men_men_n336_), .B(men_men_n335_), .Y(men_men_n337_));
  OAI210     u321(.A0(men_men_n119_), .A1(men_men_n107_), .B0(men_men_n178_), .Y(men_men_n338_));
  NA3        u322(.A(men_men_n338_), .B(x6), .C(x3), .Y(men_men_n339_));
  NOi21      u323(.An(men_men_n151_), .B(men_men_n131_), .Y(men_men_n340_));
  AOI210     u324(.A0(x8), .A1(x0), .B0(x1), .Y(men_men_n341_));
  OAI220     u325(.A0(men_men_n341_), .A1(men_men_n314_), .B0(men_men_n271_), .B1(men_men_n311_), .Y(men_men_n342_));
  AOI210     u326(.A0(men_men_n340_), .A1(men_men_n63_), .B0(men_men_n342_), .Y(men_men_n343_));
  NA2        u327(.A(x2), .B(men_men_n17_), .Y(men_men_n344_));
  OAI210     u328(.A0(men_men_n107_), .A1(men_men_n17_), .B0(men_men_n344_), .Y(men_men_n345_));
  AOI220     u329(.A0(men_men_n345_), .A1(men_men_n79_), .B0(men_men_n327_), .B1(men_men_n93_), .Y(men_men_n346_));
  NA4        u330(.A(men_men_n346_), .B(men_men_n343_), .C(men_men_n339_), .D(men_men_n337_), .Y(men_men_n347_));
  OAI210     u331(.A0(men_men_n112_), .A1(x3), .B0(men_men_n304_), .Y(men_men_n348_));
  NA3        u332(.A(men_men_n227_), .B(men_men_n213_), .C(men_men_n84_), .Y(men_men_n349_));
  NA3        u333(.A(men_men_n349_), .B(men_men_n348_), .C(men_men_n154_), .Y(men_men_n350_));
  AOI210     u334(.A0(men_men_n347_), .A1(x4), .B0(men_men_n350_), .Y(men_men_n351_));
  NA3        u335(.A(men_men_n324_), .B(men_men_n209_), .C(men_men_n93_), .Y(men_men_n352_));
  NOi21      u336(.An(x4), .B(x0), .Y(men_men_n353_));
  XO2        u337(.A(x4), .B(x0), .Y(men_men_n354_));
  OAI210     u338(.A0(men_men_n354_), .A1(men_men_n118_), .B0(men_men_n266_), .Y(men_men_n355_));
  AOI220     u339(.A0(men_men_n355_), .A1(x8), .B0(men_men_n353_), .B1(men_men_n94_), .Y(men_men_n356_));
  AOI210     u340(.A0(men_men_n356_), .A1(men_men_n352_), .B0(x3), .Y(men_men_n357_));
  INV        u341(.A(men_men_n94_), .Y(men_men_n358_));
  NO2        u342(.A(men_men_n93_), .B(x4), .Y(men_men_n359_));
  AOI220     u343(.A0(men_men_n359_), .A1(men_men_n44_), .B0(men_men_n128_), .B1(men_men_n358_), .Y(men_men_n360_));
  NO3        u344(.A(men_men_n354_), .B(men_men_n165_), .C(x2), .Y(men_men_n361_));
  NO3        u345(.A(men_men_n227_), .B(men_men_n28_), .C(men_men_n24_), .Y(men_men_n362_));
  NO2        u346(.A(men_men_n362_), .B(men_men_n361_), .Y(men_men_n363_));
  NA4        u347(.A(men_men_n363_), .B(men_men_n360_), .C(men_men_n223_), .D(x6), .Y(men_men_n364_));
  OAI220     u348(.A0(men_men_n303_), .A1(men_men_n91_), .B0(men_men_n183_), .B1(men_men_n93_), .Y(men_men_n365_));
  NO2        u349(.A(men_men_n43_), .B(x0), .Y(men_men_n366_));
  OR2        u350(.A(men_men_n359_), .B(men_men_n366_), .Y(men_men_n367_));
  NO2        u351(.A(men_men_n151_), .B(men_men_n107_), .Y(men_men_n368_));
  AOI220     u352(.A0(men_men_n368_), .A1(men_men_n367_), .B0(men_men_n365_), .B1(men_men_n61_), .Y(men_men_n369_));
  NO2        u353(.A(men_men_n151_), .B(men_men_n81_), .Y(men_men_n370_));
  NO2        u354(.A(men_men_n35_), .B(x2), .Y(men_men_n371_));
  NOi21      u355(.An(men_men_n124_), .B(men_men_n27_), .Y(men_men_n372_));
  AOI210     u356(.A0(men_men_n371_), .A1(men_men_n370_), .B0(men_men_n372_), .Y(men_men_n373_));
  OAI210     u357(.A0(men_men_n369_), .A1(men_men_n62_), .B0(men_men_n373_), .Y(men_men_n374_));
  OAI220     u358(.A0(men_men_n374_), .A1(x6), .B0(men_men_n364_), .B1(men_men_n357_), .Y(men_men_n375_));
  OAI210     u359(.A0(men_men_n63_), .A1(men_men_n48_), .B0(men_men_n42_), .Y(men_men_n376_));
  OAI210     u360(.A0(men_men_n376_), .A1(men_men_n93_), .B0(men_men_n315_), .Y(men_men_n377_));
  AOI210     u361(.A0(men_men_n377_), .A1(men_men_n18_), .B0(men_men_n154_), .Y(men_men_n378_));
  AO220      u362(.A0(men_men_n378_), .A1(men_men_n375_), .B0(men_men_n351_), .B1(men_men_n334_), .Y(men_men_n379_));
  NA2        u363(.A(men_men_n371_), .B(x6), .Y(men_men_n380_));
  AOI210     u364(.A0(x6), .A1(x1), .B0(men_men_n153_), .Y(men_men_n381_));
  NA2        u365(.A(men_men_n359_), .B(x0), .Y(men_men_n382_));
  NA2        u366(.A(men_men_n84_), .B(x6), .Y(men_men_n383_));
  OAI210     u367(.A0(men_men_n382_), .A1(men_men_n381_), .B0(men_men_n383_), .Y(men_men_n384_));
  AOI220     u368(.A0(men_men_n384_), .A1(men_men_n380_), .B0(men_men_n217_), .B1(men_men_n49_), .Y(men_men_n385_));
  NA3        u369(.A(men_men_n385_), .B(men_men_n379_), .C(men_men_n321_), .Y(men_men_n386_));
  AOI210     u370(.A0(men_men_n201_), .A1(x8), .B0(men_men_n112_), .Y(men_men_n387_));
  NA2        u371(.A(men_men_n387_), .B(men_men_n344_), .Y(men_men_n388_));
  NA3        u372(.A(men_men_n388_), .B(men_men_n199_), .C(men_men_n154_), .Y(men_men_n389_));
  OAI210     u373(.A0(men_men_n28_), .A1(x1), .B0(men_men_n231_), .Y(men_men_n390_));
  AO220      u374(.A0(men_men_n390_), .A1(men_men_n150_), .B0(men_men_n111_), .B1(x4), .Y(men_men_n391_));
  NA3        u375(.A(x7), .B(x3), .C(x0), .Y(men_men_n392_));
  NA2        u376(.A(men_men_n222_), .B(x0), .Y(men_men_n393_));
  OAI220     u377(.A0(men_men_n393_), .A1(men_men_n209_), .B0(men_men_n392_), .B1(men_men_n358_), .Y(men_men_n394_));
  AOI210     u378(.A0(men_men_n391_), .A1(men_men_n120_), .B0(men_men_n394_), .Y(men_men_n395_));
  AOI210     u379(.A0(men_men_n395_), .A1(men_men_n389_), .B0(men_men_n25_), .Y(men_men_n396_));
  NA3        u380(.A(men_men_n122_), .B(men_men_n222_), .C(x0), .Y(men_men_n397_));
  OAI210     u381(.A0(men_men_n199_), .A1(men_men_n67_), .B0(men_men_n205_), .Y(men_men_n398_));
  NA3        u382(.A(men_men_n201_), .B(men_men_n224_), .C(x8), .Y(men_men_n399_));
  AOI210     u383(.A0(men_men_n399_), .A1(men_men_n398_), .B0(men_men_n25_), .Y(men_men_n400_));
  AOI210     u384(.A0(men_men_n121_), .A1(men_men_n119_), .B0(men_men_n42_), .Y(men_men_n401_));
  NOi31      u385(.An(men_men_n401_), .B(men_men_n366_), .C(men_men_n184_), .Y(men_men_n402_));
  OAI210     u386(.A0(men_men_n402_), .A1(men_men_n400_), .B0(men_men_n150_), .Y(men_men_n403_));
  NAi31      u387(.An(men_men_n50_), .B(men_men_n292_), .C(men_men_n179_), .Y(men_men_n404_));
  NA3        u388(.A(men_men_n404_), .B(men_men_n403_), .C(men_men_n397_), .Y(men_men_n405_));
  OAI210     u389(.A0(men_men_n405_), .A1(men_men_n396_), .B0(x6), .Y(men_men_n406_));
  OAI210     u390(.A0(men_men_n165_), .A1(men_men_n48_), .B0(men_men_n136_), .Y(men_men_n407_));
  NA3        u391(.A(men_men_n55_), .B(men_men_n38_), .C(men_men_n31_), .Y(men_men_n408_));
  AOI220     u392(.A0(men_men_n408_), .A1(men_men_n407_), .B0(men_men_n40_), .B1(men_men_n32_), .Y(men_men_n409_));
  NO2        u393(.A(men_men_n154_), .B(x0), .Y(men_men_n410_));
  AOI220     u394(.A0(men_men_n410_), .A1(men_men_n222_), .B0(men_men_n199_), .B1(men_men_n154_), .Y(men_men_n411_));
  INV        u395(.A(x1), .Y(men_men_n412_));
  OAI210     u396(.A0(men_men_n411_), .A1(x8), .B0(men_men_n412_), .Y(men_men_n413_));
  NAi31      u397(.An(x2), .B(x8), .C(x0), .Y(men_men_n414_));
  OAI210     u398(.A0(men_men_n414_), .A1(x4), .B0(men_men_n166_), .Y(men_men_n415_));
  NA3        u399(.A(men_men_n415_), .B(men_men_n148_), .C(x9), .Y(men_men_n416_));
  NO3        u400(.A(x9), .B(men_men_n154_), .C(x0), .Y(men_men_n417_));
  AOI220     u401(.A0(men_men_n417_), .A1(men_men_n245_), .B0(men_men_n370_), .B1(men_men_n154_), .Y(men_men_n418_));
  NA4        u402(.A(men_men_n418_), .B(x1), .C(men_men_n416_), .D(men_men_n50_), .Y(men_men_n419_));
  OAI210     u403(.A0(men_men_n413_), .A1(men_men_n409_), .B0(men_men_n419_), .Y(men_men_n420_));
  NOi31      u404(.An(men_men_n410_), .B(men_men_n32_), .C(x8), .Y(men_men_n421_));
  AOI210     u405(.A0(men_men_n38_), .A1(x9), .B0(men_men_n134_), .Y(men_men_n422_));
  NO3        u406(.A(men_men_n422_), .B(men_men_n127_), .C(men_men_n43_), .Y(men_men_n423_));
  NOi31      u407(.An(x1), .B(x8), .C(x7), .Y(men_men_n424_));
  AOI220     u408(.A0(men_men_n424_), .A1(men_men_n353_), .B0(men_men_n128_), .B1(x3), .Y(men_men_n425_));
  AOI210     u409(.A0(men_men_n266_), .A1(men_men_n60_), .B0(men_men_n126_), .Y(men_men_n426_));
  OAI210     u410(.A0(men_men_n426_), .A1(x3), .B0(men_men_n425_), .Y(men_men_n427_));
  NO3        u411(.A(men_men_n427_), .B(men_men_n423_), .C(x2), .Y(men_men_n428_));
  OAI220     u412(.A0(men_men_n354_), .A1(men_men_n307_), .B0(men_men_n303_), .B1(men_men_n43_), .Y(men_men_n429_));
  INV        u413(.A(men_men_n392_), .Y(men_men_n430_));
  AOI220     u414(.A0(men_men_n430_), .A1(men_men_n93_), .B0(men_men_n429_), .B1(men_men_n154_), .Y(men_men_n431_));
  NO2        u415(.A(men_men_n431_), .B(men_men_n54_), .Y(men_men_n432_));
  NO3        u416(.A(men_men_n432_), .B(men_men_n428_), .C(men_men_n421_), .Y(men_men_n433_));
  AOI210     u417(.A0(men_men_n433_), .A1(men_men_n420_), .B0(men_men_n25_), .Y(men_men_n434_));
  NA4        u418(.A(men_men_n31_), .B(men_men_n93_), .C(x2), .D(men_men_n17_), .Y(men_men_n435_));
  NO3        u419(.A(men_men_n62_), .B(x4), .C(x1), .Y(men_men_n436_));
  NO3        u420(.A(men_men_n67_), .B(men_men_n18_), .C(x0), .Y(men_men_n437_));
  AOI220     u421(.A0(men_men_n437_), .A1(men_men_n267_), .B0(men_men_n436_), .B1(men_men_n401_), .Y(men_men_n438_));
  NO2        u422(.A(men_men_n438_), .B(men_men_n104_), .Y(men_men_n439_));
  NO3        u423(.A(men_men_n271_), .B(men_men_n178_), .C(men_men_n40_), .Y(men_men_n440_));
  OAI210     u424(.A0(men_men_n440_), .A1(men_men_n439_), .B0(x7), .Y(men_men_n441_));
  NA2        u425(.A(men_men_n227_), .B(x7), .Y(men_men_n442_));
  NA3        u426(.A(men_men_n442_), .B(men_men_n153_), .C(men_men_n135_), .Y(men_men_n443_));
  NA3        u427(.A(men_men_n443_), .B(men_men_n441_), .C(men_men_n435_), .Y(men_men_n444_));
  OAI210     u428(.A0(men_men_n444_), .A1(men_men_n434_), .B0(men_men_n36_), .Y(men_men_n445_));
  NO2        u429(.A(men_men_n417_), .B(men_men_n205_), .Y(men_men_n446_));
  NO4        u430(.A(men_men_n446_), .B(men_men_n78_), .C(x4), .D(men_men_n54_), .Y(men_men_n447_));
  NA2        u431(.A(men_men_n255_), .B(men_men_n21_), .Y(men_men_n448_));
  NO2        u432(.A(men_men_n162_), .B(men_men_n136_), .Y(men_men_n449_));
  NA2        u433(.A(men_men_n449_), .B(men_men_n448_), .Y(men_men_n450_));
  AOI210     u434(.A0(men_men_n450_), .A1(men_men_n169_), .B0(men_men_n28_), .Y(men_men_n451_));
  AOI220     u435(.A0(men_men_n366_), .A1(men_men_n93_), .B0(men_men_n151_), .B1(men_men_n201_), .Y(men_men_n452_));
  NA3        u436(.A(men_men_n452_), .B(men_men_n414_), .C(men_men_n91_), .Y(men_men_n453_));
  NA2        u437(.A(men_men_n453_), .B(men_men_n179_), .Y(men_men_n454_));
  OAI220     u438(.A0(men_men_n279_), .A1(men_men_n68_), .B0(men_men_n162_), .B1(men_men_n43_), .Y(men_men_n455_));
  NA2        u439(.A(x3), .B(men_men_n54_), .Y(men_men_n456_));
  AOI210     u440(.A0(men_men_n166_), .A1(men_men_n27_), .B0(men_men_n73_), .Y(men_men_n457_));
  OAI210     u441(.A0(men_men_n150_), .A1(men_men_n18_), .B0(men_men_n21_), .Y(men_men_n458_));
  NO3        u442(.A(men_men_n424_), .B(x3), .C(men_men_n54_), .Y(men_men_n459_));
  AOI210     u443(.A0(men_men_n459_), .A1(men_men_n458_), .B0(men_men_n457_), .Y(men_men_n460_));
  OAI210     u444(.A0(men_men_n155_), .A1(men_men_n456_), .B0(men_men_n460_), .Y(men_men_n461_));
  AOI220     u445(.A0(men_men_n461_), .A1(x0), .B0(men_men_n455_), .B1(men_men_n136_), .Y(men_men_n462_));
  AOI210     u446(.A0(men_men_n462_), .A1(men_men_n454_), .B0(men_men_n235_), .Y(men_men_n463_));
  NA2        u447(.A(x9), .B(x5), .Y(men_men_n464_));
  NO4        u448(.A(men_men_n107_), .B(men_men_n464_), .C(men_men_n60_), .D(men_men_n32_), .Y(men_men_n465_));
  NO4        u449(.A(men_men_n465_), .B(men_men_n463_), .C(men_men_n451_), .D(men_men_n447_), .Y(men_men_n466_));
  NA3        u450(.A(men_men_n466_), .B(men_men_n445_), .C(men_men_n406_), .Y(men_men_n467_));
  AOI210     u451(.A0(men_men_n386_), .A1(men_men_n25_), .B0(men_men_n467_), .Y(men05));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
endmodule