// Benchmark "top" written by ABC on Thu Jun 20 14:59:13 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output mai1, mai2, mai0, mai7, mai5, mai6, mai3, mai4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n43_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n83_, new_new_n84_,
    new_new_n86_, new_new_n87_, new_new_n88_, new_new_n89_, new_new_n90_,
    new_new_n91_, new_new_n92_, new_new_n93_, new_new_n94_, new_new_n95_,
    new_new_n96_, new_new_n97_, new_new_n98_, new_new_n99_, new_new_n100_,
    new_new_n101_, new_new_n102_, new_new_n103_, new_new_n104_,
    new_new_n105_, new_new_n106_, new_new_n107_, new_new_n108_,
    new_new_n109_, new_new_n110_, new_new_n111_, new_new_n112_,
    new_new_n113_, new_new_n114_, new_new_n115_, new_new_n116_,
    new_new_n117_, new_new_n118_, new_new_n119_, new_new_n120_,
    new_new_n121_, new_new_n122_, new_new_n123_, new_new_n124_,
    new_new_n125_, new_new_n126_, new_new_n127_, new_new_n128_,
    new_new_n129_, new_new_n130_, new_new_n131_, new_new_n132_,
    new_new_n133_, new_new_n134_, new_new_n135_, new_new_n136_,
    new_new_n137_, new_new_n138_, new_new_n139_, new_new_n140_,
    new_new_n141_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n267_, new_new_n268_, new_new_n269_,
    new_new_n270_, new_new_n271_, new_new_n272_, new_new_n273_,
    new_new_n274_, new_new_n275_, new_new_n276_, new_new_n277_,
    new_new_n278_, new_new_n279_, new_new_n280_, new_new_n281_,
    new_new_n282_, new_new_n283_, new_new_n284_, new_new_n285_,
    new_new_n286_, new_new_n287_, new_new_n288_, new_new_n289_,
    new_new_n290_, new_new_n291_, new_new_n292_, new_new_n293_,
    new_new_n294_, new_new_n295_, new_new_n296_, new_new_n297_,
    new_new_n298_, new_new_n299_, new_new_n300_, new_new_n301_,
    new_new_n302_, new_new_n303_, new_new_n304_, new_new_n305_,
    new_new_n306_, new_new_n307_, new_new_n308_, new_new_n309_,
    new_new_n310_, new_new_n311_, new_new_n312_, new_new_n313_,
    new_new_n315_, new_new_n316_, new_new_n317_, new_new_n318_,
    new_new_n319_, new_new_n320_, new_new_n321_, new_new_n322_,
    new_new_n323_, new_new_n324_, new_new_n325_, new_new_n326_,
    new_new_n327_, new_new_n328_, new_new_n329_, new_new_n330_,
    new_new_n331_, new_new_n332_, new_new_n333_, new_new_n334_,
    new_new_n335_, new_new_n336_, new_new_n337_, new_new_n338_,
    new_new_n339_, new_new_n340_, new_new_n341_, new_new_n342_,
    new_new_n343_, new_new_n344_, new_new_n345_, new_new_n346_,
    new_new_n347_, new_new_n348_, new_new_n349_, new_new_n350_,
    new_new_n351_, new_new_n352_, new_new_n353_, new_new_n355_,
    new_new_n356_, new_new_n357_, new_new_n358_, new_new_n359_,
    new_new_n360_, new_new_n361_, new_new_n362_, new_new_n363_,
    new_new_n364_, new_new_n365_, new_new_n366_, new_new_n367_,
    new_new_n368_, new_new_n369_, new_new_n370_, new_new_n371_,
    new_new_n372_, new_new_n373_, new_new_n374_, new_new_n375_,
    new_new_n376_, new_new_n377_, new_new_n378_, new_new_n379_,
    new_new_n380_, new_new_n381_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n429_, new_new_n430_, new_new_n431_,
    new_new_n432_, new_new_n433_, new_new_n434_, new_new_n435_,
    new_new_n436_, new_new_n437_, new_new_n438_, new_new_n439_,
    new_new_n440_, new_new_n441_, new_new_n442_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NOi21      g016(.An(i_12_), .B(i_13_), .Y(new_new_n39_));
  INV        g017(.A(new_new_n39_), .Y(new_new_n40_));
  NAi31      g018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n41_));
  INV        g019(.A(new_new_n35_), .Y(mai1));
  INV        g020(.A(i_11_), .Y(new_new_n43_));
  NO2        g021(.A(new_new_n43_), .B(i_6_), .Y(new_new_n44_));
  INV        g022(.A(i_2_), .Y(new_new_n45_));
  INV        g023(.A(i_5_), .Y(new_new_n46_));
  NO2        g024(.A(i_7_), .B(i_10_), .Y(new_new_n47_));
  AOI210     g025(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n47_), .Y(new_new_n48_));
  INV        g026(.A(i_1_), .Y(new_new_n49_));
  NA2        g027(.A(new_new_n48_), .B(i_2_), .Y(new_new_n50_));
  AOI210     g028(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n51_));
  NA2        g029(.A(i_1_), .B(i_6_), .Y(new_new_n52_));
  NO2        g030(.A(new_new_n52_), .B(new_new_n25_), .Y(new_new_n53_));
  INV        g031(.A(i_0_), .Y(new_new_n54_));
  NAi21      g032(.An(i_5_), .B(i_10_), .Y(new_new_n55_));
  NA2        g033(.A(i_5_), .B(i_9_), .Y(new_new_n56_));
  AOI210     g034(.A0(new_new_n56_), .A1(new_new_n55_), .B0(new_new_n54_), .Y(new_new_n57_));
  NO2        g035(.A(new_new_n57_), .B(new_new_n53_), .Y(new_new_n58_));
  NA2        g036(.A(i_12_), .B(i_5_), .Y(new_new_n59_));
  NO2        g037(.A(i_3_), .B(i_9_), .Y(new_new_n60_));
  INV        g038(.A(i_6_), .Y(new_new_n61_));
  INV        g039(.A(i_11_), .Y(new_new_n62_));
  NO2        g040(.A(i_2_), .B(i_7_), .Y(new_new_n63_));
  NAi21      g041(.An(i_6_), .B(i_10_), .Y(new_new_n64_));
  NA2        g042(.A(i_6_), .B(i_9_), .Y(new_new_n65_));
  AN3        g043(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n66_));
  NAi21      g044(.An(i_6_), .B(i_11_), .Y(new_new_n67_));
  NA2        g045(.A(new_new_n66_), .B(new_new_n32_), .Y(new_new_n68_));
  INV        g046(.A(i_7_), .Y(new_new_n69_));
  NO2        g047(.A(i_0_), .B(i_5_), .Y(new_new_n70_));
  NO2        g048(.A(i_2_), .B(i_7_), .Y(new_new_n71_));
  NA2        g049(.A(i_12_), .B(i_7_), .Y(new_new_n72_));
  NO2        g050(.A(new_new_n49_), .B(new_new_n26_), .Y(new_new_n73_));
  NA2        g051(.A(i_11_), .B(i_12_), .Y(new_new_n74_));
  NA2        g052(.A(new_new_n74_), .B(new_new_n68_), .Y(new_new_n75_));
  NA2        g053(.A(new_new_n69_), .B(new_new_n37_), .Y(new_new_n76_));
  NA2        g054(.A(i_7_), .B(new_new_n25_), .Y(new_new_n77_));
  NA2        g055(.A(new_new_n77_), .B(new_new_n76_), .Y(new_new_n78_));
  NO2        g056(.A(new_new_n78_), .B(new_new_n45_), .Y(new_new_n79_));
  NA2        g057(.A(new_new_n65_), .B(new_new_n64_), .Y(new_new_n80_));
  INV        g058(.A(new_new_n75_), .Y(new_new_n81_));
  NA2        g059(.A(new_new_n81_), .B(new_new_n436_), .Y(mai2));
  NO2        g060(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n83_));
  NA2        g061(.A(new_new_n432_), .B(new_new_n83_), .Y(new_new_n84_));
  NA4        g062(.A(new_new_n84_), .B(new_new_n58_), .C(new_new_n50_), .D(new_new_n30_), .Y(mai0));
  AN2        g063(.A(i_8_), .B(i_7_), .Y(new_new_n86_));
  NO2        g064(.A(i_12_), .B(i_13_), .Y(new_new_n87_));
  NAi21      g065(.An(i_5_), .B(i_11_), .Y(new_new_n88_));
  NOi21      g066(.An(new_new_n87_), .B(new_new_n88_), .Y(new_new_n89_));
  NO2        g067(.A(i_0_), .B(i_1_), .Y(new_new_n90_));
  NA2        g068(.A(i_2_), .B(i_3_), .Y(new_new_n91_));
  NO2        g069(.A(new_new_n91_), .B(i_4_), .Y(new_new_n92_));
  AN2        g070(.A(new_new_n87_), .B(new_new_n60_), .Y(new_new_n93_));
  OR2        g071(.A(i_0_), .B(i_1_), .Y(new_new_n94_));
  NO3        g072(.A(new_new_n94_), .B(new_new_n59_), .C(i_13_), .Y(new_new_n95_));
  NAi32      g073(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n96_));
  NAi21      g074(.An(new_new_n96_), .B(new_new_n95_), .Y(new_new_n97_));
  NOi21      g075(.An(i_4_), .B(i_10_), .Y(new_new_n98_));
  NA2        g076(.A(new_new_n98_), .B(new_new_n39_), .Y(new_new_n99_));
  NOi21      g077(.An(i_11_), .B(i_13_), .Y(new_new_n100_));
  NA2        g078(.A(new_new_n100_), .B(i_4_), .Y(new_new_n101_));
  NO2        g079(.A(new_new_n54_), .B(new_new_n49_), .Y(new_new_n102_));
  NA2        g080(.A(i_3_), .B(i_5_), .Y(new_new_n103_));
  NO2        g081(.A(new_new_n54_), .B(i_5_), .Y(new_new_n104_));
  NO2        g082(.A(i_13_), .B(i_10_), .Y(new_new_n105_));
  NA3        g083(.A(new_new_n105_), .B(new_new_n104_), .C(new_new_n43_), .Y(new_new_n106_));
  NAi21      g084(.An(i_4_), .B(i_12_), .Y(new_new_n107_));
  INV        g085(.A(i_8_), .Y(new_new_n108_));
  NO3        g086(.A(i_3_), .B(new_new_n61_), .C(new_new_n46_), .Y(new_new_n109_));
  INV        g087(.A(new_new_n109_), .Y(new_new_n110_));
  NO2        g088(.A(i_0_), .B(i_1_), .Y(new_new_n111_));
  NA3        g089(.A(new_new_n111_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n112_));
  NO3        g090(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n113_));
  NA2        g091(.A(i_12_), .B(new_new_n113_), .Y(new_new_n114_));
  AOI210     g092(.A0(new_new_n114_), .A1(new_new_n112_), .B0(new_new_n110_), .Y(new_new_n115_));
  NO3        g093(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n116_));
  NO2        g094(.A(i_13_), .B(i_9_), .Y(new_new_n117_));
  NAi21      g095(.An(i_12_), .B(i_3_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n43_), .B(i_5_), .Y(new_new_n119_));
  NA3        g097(.A(i_13_), .B(new_new_n108_), .C(i_10_), .Y(new_new_n120_));
  NO2        g098(.A(new_new_n120_), .B(i_12_), .Y(new_new_n121_));
  NA2        g099(.A(i_0_), .B(i_5_), .Y(new_new_n122_));
  NAi31      g100(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n123_));
  NO2        g101(.A(new_new_n45_), .B(new_new_n49_), .Y(new_new_n124_));
  INV        g102(.A(i_13_), .Y(new_new_n125_));
  NO2        g103(.A(i_12_), .B(new_new_n125_), .Y(new_new_n126_));
  NA3        g104(.A(new_new_n126_), .B(new_new_n111_), .C(new_new_n109_), .Y(new_new_n127_));
  INV        g105(.A(new_new_n127_), .Y(new_new_n128_));
  AOI220     g106(.A0(new_new_n128_), .A1(new_new_n86_), .B0(i_3_), .B1(new_new_n121_), .Y(new_new_n129_));
  INV        g107(.A(i_12_), .Y(new_new_n130_));
  NO3        g108(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n131_));
  NA2        g109(.A(i_2_), .B(i_1_), .Y(new_new_n132_));
  NO3        g110(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n133_));
  NAi21      g111(.An(i_4_), .B(i_3_), .Y(new_new_n134_));
  NOi41      g112(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n135_));
  NO2        g113(.A(i_11_), .B(new_new_n125_), .Y(new_new_n136_));
  NO2        g114(.A(i_12_), .B(i_3_), .Y(new_new_n137_));
  NA2        g115(.A(new_new_n130_), .B(i_13_), .Y(new_new_n138_));
  NO2        g116(.A(new_new_n138_), .B(new_new_n56_), .Y(new_new_n139_));
  NA2        g117(.A(new_new_n139_), .B(new_new_n86_), .Y(new_new_n140_));
  NO2        g118(.A(i_8_), .B(new_new_n37_), .Y(new_new_n141_));
  NA2        g119(.A(i_12_), .B(i_6_), .Y(new_new_n142_));
  NO2        g120(.A(new_new_n134_), .B(i_2_), .Y(new_new_n143_));
  NA3        g121(.A(new_new_n143_), .B(new_new_n434_), .C(new_new_n43_), .Y(new_new_n144_));
  NA2        g122(.A(new_new_n136_), .B(i_9_), .Y(new_new_n145_));
  INV        g123(.A(new_new_n144_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(new_new_n141_), .Y(new_new_n147_));
  NA3        g125(.A(new_new_n147_), .B(new_new_n140_), .C(new_new_n129_), .Y(new_new_n148_));
  NO3        g126(.A(i_12_), .B(new_new_n125_), .C(new_new_n37_), .Y(new_new_n149_));
  INV        g127(.A(new_new_n149_), .Y(new_new_n150_));
  NO2        g128(.A(i_3_), .B(i_10_), .Y(new_new_n151_));
  NA3        g129(.A(new_new_n151_), .B(new_new_n39_), .C(new_new_n43_), .Y(new_new_n152_));
  AN2        g130(.A(i_3_), .B(i_10_), .Y(new_new_n153_));
  NO2        g131(.A(i_5_), .B(new_new_n37_), .Y(new_new_n154_));
  OAI220     g132(.A0(new_new_n152_), .A1(i_6_), .B0(new_new_n442_), .B1(new_new_n150_), .Y(new_new_n155_));
  NO3        g133(.A(new_new_n155_), .B(new_new_n148_), .C(new_new_n115_), .Y(new_new_n156_));
  NO3        g134(.A(new_new_n43_), .B(i_13_), .C(i_9_), .Y(new_new_n157_));
  NOi21      g135(.An(i_5_), .B(i_0_), .Y(new_new_n158_));
  INV        g136(.A(new_new_n99_), .Y(new_new_n159_));
  AOI210     g137(.A0(i_4_), .A1(new_new_n157_), .B0(new_new_n159_), .Y(new_new_n160_));
  NOi32      g138(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n161_));
  INV        g139(.A(new_new_n161_), .Y(new_new_n162_));
  NO2        g140(.A(i_9_), .B(new_new_n96_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n164_));
  NOi32      g142(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n165_));
  NA2        g143(.A(new_new_n165_), .B(new_new_n45_), .Y(new_new_n166_));
  NO2        g144(.A(new_new_n166_), .B(i_0_), .Y(new_new_n167_));
  OR2        g145(.A(new_new_n167_), .B(new_new_n164_), .Y(new_new_n168_));
  NAi21      g146(.An(i_3_), .B(i_4_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_9_), .Y(new_new_n170_));
  NA2        g148(.A(i_7_), .B(new_new_n170_), .Y(new_new_n171_));
  NA2        g149(.A(i_2_), .B(i_7_), .Y(new_new_n172_));
  NO2        g150(.A(new_new_n169_), .B(i_10_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n171_), .B(new_new_n104_), .Y(new_new_n174_));
  INV        g152(.A(new_new_n173_), .Y(new_new_n175_));
  NO2        g153(.A(new_new_n175_), .B(i_5_), .Y(new_new_n176_));
  NO4        g154(.A(new_new_n176_), .B(new_new_n174_), .C(new_new_n168_), .D(new_new_n163_), .Y(new_new_n177_));
  NO2        g155(.A(new_new_n177_), .B(new_new_n162_), .Y(new_new_n178_));
  AN2        g156(.A(i_12_), .B(i_5_), .Y(new_new_n179_));
  NA2        g157(.A(i_3_), .B(new_new_n179_), .Y(new_new_n180_));
  NO2        g158(.A(i_11_), .B(i_6_), .Y(new_new_n181_));
  NA3        g159(.A(new_new_n181_), .B(i_2_), .C(new_new_n125_), .Y(new_new_n182_));
  NO2        g160(.A(new_new_n182_), .B(new_new_n180_), .Y(new_new_n183_));
  NO2        g161(.A(i_5_), .B(i_10_), .Y(new_new_n184_));
  INV        g162(.A(new_new_n183_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n186_));
  NO3        g164(.A(new_new_n61_), .B(new_new_n46_), .C(i_9_), .Y(new_new_n187_));
  INV        g165(.A(new_new_n123_), .Y(new_new_n188_));
  NAi21      g166(.An(i_13_), .B(i_0_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n189_), .B(new_new_n132_), .Y(new_new_n190_));
  NA2        g168(.A(new_new_n188_), .B(new_new_n190_), .Y(new_new_n191_));
  NA2        g169(.A(new_new_n191_), .B(new_new_n185_), .Y(new_new_n192_));
  NA2        g170(.A(new_new_n43_), .B(new_new_n125_), .Y(new_new_n193_));
  NO2        g171(.A(i_0_), .B(i_11_), .Y(new_new_n194_));
  AN2        g172(.A(i_1_), .B(i_6_), .Y(new_new_n195_));
  NA2        g173(.A(new_new_n86_), .B(i_9_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n196_), .B(i_4_), .Y(new_new_n197_));
  OR2        g175(.A(i_13_), .B(i_10_), .Y(new_new_n198_));
  NO2        g176(.A(new_new_n69_), .B(new_new_n25_), .Y(new_new_n199_));
  INV        g177(.A(new_new_n145_), .Y(new_new_n200_));
  NO3        g178(.A(new_new_n200_), .B(new_new_n192_), .C(new_new_n178_), .Y(new_new_n201_));
  NO2        g179(.A(new_new_n54_), .B(i_13_), .Y(new_new_n202_));
  NO2        g180(.A(i_10_), .B(i_9_), .Y(new_new_n203_));
  NO2        g181(.A(i_12_), .B(i_3_), .Y(new_new_n204_));
  NA2        g182(.A(i_8_), .B(i_9_), .Y(new_new_n205_));
  INV        g183(.A(new_new_n149_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n206_), .B(new_new_n205_), .Y(new_new_n207_));
  NA2        g185(.A(new_new_n136_), .B(new_new_n154_), .Y(new_new_n208_));
  NO3        g186(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n209_));
  INV        g187(.A(new_new_n209_), .Y(new_new_n210_));
  NA3        g188(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n211_));
  NA3        g189(.A(new_new_n88_), .B(new_new_n73_), .C(new_new_n23_), .Y(new_new_n212_));
  OAI220     g190(.A0(new_new_n212_), .A1(new_new_n211_), .B0(new_new_n210_), .B1(new_new_n208_), .Y(new_new_n213_));
  NO2        g191(.A(new_new_n213_), .B(new_new_n207_), .Y(new_new_n214_));
  NA2        g192(.A(new_new_n66_), .B(i_13_), .Y(new_new_n215_));
  NA2        g193(.A(i_3_), .B(i_9_), .Y(new_new_n216_));
  NO2        g194(.A(new_new_n216_), .B(new_new_n215_), .Y(new_new_n217_));
  NO2        g195(.A(i_11_), .B(i_1_), .Y(new_new_n218_));
  NA2        g196(.A(i_2_), .B(i_0_), .Y(new_new_n219_));
  NO2        g197(.A(new_new_n198_), .B(i_6_), .Y(new_new_n220_));
  NA2        g198(.A(new_new_n220_), .B(i_1_), .Y(new_new_n221_));
  NO2        g199(.A(new_new_n221_), .B(new_new_n219_), .Y(new_new_n222_));
  NO2        g200(.A(i_6_), .B(i_10_), .Y(new_new_n223_));
  NA2        g201(.A(new_new_n135_), .B(new_new_n100_), .Y(new_new_n224_));
  NO2        g202(.A(new_new_n94_), .B(i_3_), .Y(new_new_n225_));
  NAi31      g203(.An(i_11_), .B(new_new_n225_), .C(new_new_n126_), .Y(new_new_n226_));
  NA3        g204(.A(new_new_n186_), .B(new_new_n102_), .C(new_new_n92_), .Y(new_new_n227_));
  NA3        g205(.A(new_new_n227_), .B(new_new_n226_), .C(new_new_n224_), .Y(new_new_n228_));
  NO3        g206(.A(new_new_n228_), .B(new_new_n222_), .C(new_new_n217_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n229_), .B(new_new_n214_), .Y(new_new_n230_));
  INV        g208(.A(new_new_n157_), .Y(new_new_n231_));
  NO2        g209(.A(new_new_n231_), .B(i_12_), .Y(new_new_n232_));
  INV        g210(.A(new_new_n232_), .Y(new_new_n233_));
  NA3        g211(.A(new_new_n202_), .B(i_1_), .C(i_2_), .Y(new_new_n234_));
  INV        g212(.A(new_new_n234_), .Y(new_new_n235_));
  NA2        g213(.A(new_new_n179_), .B(new_new_n125_), .Y(new_new_n236_));
  NA2        g214(.A(i_7_), .B(new_new_n165_), .Y(new_new_n237_));
  OR2        g215(.A(new_new_n236_), .B(new_new_n237_), .Y(new_new_n238_));
  NO2        g216(.A(new_new_n36_), .B(i_8_), .Y(new_new_n239_));
  INV        g217(.A(new_new_n238_), .Y(new_new_n240_));
  AOI210     g218(.A0(new_new_n235_), .A1(new_new_n116_), .B0(new_new_n240_), .Y(new_new_n241_));
  NO2        g219(.A(i_7_), .B(new_new_n112_), .Y(new_new_n242_));
  NA2        g220(.A(i_5_), .B(new_new_n242_), .Y(new_new_n243_));
  NA3        g221(.A(new_new_n243_), .B(new_new_n241_), .C(new_new_n233_), .Y(new_new_n244_));
  NOi31      g222(.An(i_8_), .B(new_new_n198_), .C(new_new_n38_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n245_), .B(new_new_n437_), .Y(new_new_n246_));
  NO2        g224(.A(i_8_), .B(i_7_), .Y(new_new_n247_));
  INV        g225(.A(new_new_n124_), .Y(new_new_n248_));
  OAI220     g226(.A0(i_9_), .A1(new_new_n103_), .B0(new_new_n248_), .B1(new_new_n134_), .Y(new_new_n249_));
  NA3        g227(.A(i_10_), .B(new_new_n249_), .C(new_new_n247_), .Y(new_new_n250_));
  NO2        g228(.A(new_new_n215_), .B(i_6_), .Y(new_new_n251_));
  NA2        g229(.A(new_new_n251_), .B(new_new_n141_), .Y(new_new_n252_));
  NO2        g230(.A(new_new_n94_), .B(i_5_), .Y(new_new_n253_));
  NA2        g231(.A(new_new_n253_), .B(new_new_n193_), .Y(new_new_n254_));
  INV        g232(.A(new_new_n254_), .Y(new_new_n255_));
  NA2        g233(.A(new_new_n255_), .B(new_new_n209_), .Y(new_new_n256_));
  NA4        g234(.A(new_new_n256_), .B(new_new_n252_), .C(new_new_n250_), .D(new_new_n246_), .Y(new_new_n257_));
  NO3        g235(.A(new_new_n41_), .B(i_2_), .C(new_new_n46_), .Y(new_new_n258_));
  NO3        g236(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n259_));
  AN4        g237(.A(new_new_n435_), .B(new_new_n197_), .C(i_3_), .D(i_2_), .Y(new_new_n260_));
  INV        g238(.A(new_new_n260_), .Y(new_new_n261_));
  NO2        g239(.A(new_new_n72_), .B(new_new_n23_), .Y(new_new_n262_));
  NOi21      g240(.An(new_new_n89_), .B(i_4_), .Y(new_new_n263_));
  NA3        g241(.A(new_new_n152_), .B(new_new_n438_), .C(new_new_n261_), .Y(new_new_n264_));
  NO4        g242(.A(new_new_n264_), .B(new_new_n257_), .C(new_new_n244_), .D(new_new_n230_), .Y(new_new_n265_));
  NA4        g243(.A(new_new_n265_), .B(new_new_n201_), .C(new_new_n160_), .D(new_new_n156_), .Y(mai7));
  NA2        g244(.A(i_11_), .B(new_new_n108_), .Y(new_new_n267_));
  NA2        g245(.A(i_12_), .B(i_8_), .Y(new_new_n268_));
  INV        g246(.A(new_new_n116_), .Y(new_new_n269_));
  OR3        g247(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n270_));
  INV        g248(.A(new_new_n113_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n270_), .B(new_new_n49_), .Y(new_new_n272_));
  NOi21      g250(.An(i_11_), .B(i_7_), .Y(new_new_n273_));
  AO210      g251(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n274_));
  NO2        g252(.A(new_new_n274_), .B(new_new_n273_), .Y(new_new_n275_));
  NA2        g253(.A(new_new_n62_), .B(new_new_n49_), .Y(new_new_n276_));
  OR2        g254(.A(new_new_n276_), .B(new_new_n40_), .Y(new_new_n277_));
  NA2        g255(.A(new_new_n126_), .B(new_new_n49_), .Y(new_new_n278_));
  NO2        g256(.A(new_new_n49_), .B(i_9_), .Y(new_new_n279_));
  NO2        g257(.A(i_1_), .B(i_12_), .Y(new_new_n280_));
  NA2        g258(.A(new_new_n278_), .B(new_new_n277_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n281_), .B(i_6_), .Y(new_new_n282_));
  NO2        g260(.A(i_6_), .B(i_11_), .Y(new_new_n283_));
  NO3        g261(.A(i_12_), .B(i_13_), .C(new_new_n61_), .Y(new_new_n284_));
  NA2        g262(.A(new_new_n284_), .B(new_new_n279_), .Y(new_new_n285_));
  INV        g263(.A(new_new_n285_), .Y(new_new_n286_));
  INV        g264(.A(i_2_), .Y(new_new_n287_));
  NA2        g265(.A(new_new_n83_), .B(i_9_), .Y(new_new_n288_));
  NO2        g266(.A(new_new_n288_), .B(new_new_n287_), .Y(new_new_n289_));
  NA2        g267(.A(new_new_n279_), .B(i_6_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(new_new_n23_), .Y(new_new_n291_));
  AOI210     g269(.A0(new_new_n218_), .A1(new_new_n199_), .B0(new_new_n133_), .Y(new_new_n292_));
  NO2        g270(.A(new_new_n292_), .B(new_new_n440_), .Y(new_new_n293_));
  NO2        g271(.A(i_11_), .B(new_new_n37_), .Y(new_new_n294_));
  OR3        g272(.A(new_new_n293_), .B(new_new_n291_), .C(new_new_n289_), .Y(new_new_n295_));
  NO2        g273(.A(new_new_n295_), .B(new_new_n286_), .Y(new_new_n296_));
  NO2        g274(.A(new_new_n130_), .B(new_new_n69_), .Y(new_new_n297_));
  NO2        g275(.A(new_new_n297_), .B(new_new_n273_), .Y(new_new_n298_));
  NA2        g276(.A(new_new_n296_), .B(new_new_n282_), .Y(new_new_n299_));
  AOI210     g277(.A0(new_new_n142_), .A1(new_new_n67_), .B0(i_1_), .Y(new_new_n300_));
  NA2        g278(.A(i_4_), .B(new_new_n300_), .Y(new_new_n301_));
  NO2        g279(.A(new_new_n301_), .B(i_13_), .Y(new_new_n302_));
  NA2        g280(.A(new_new_n80_), .B(i_13_), .Y(new_new_n303_));
  NO2        g281(.A(new_new_n303_), .B(new_new_n300_), .Y(new_new_n304_));
  NO2        g282(.A(new_new_n130_), .B(new_new_n61_), .Y(new_new_n305_));
  NO2        g283(.A(new_new_n431_), .B(new_new_n271_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(new_new_n304_), .Y(new_new_n307_));
  NA2        g285(.A(new_new_n283_), .B(i_13_), .Y(new_new_n308_));
  INV        g286(.A(new_new_n308_), .Y(new_new_n309_));
  NA2        g287(.A(new_new_n309_), .B(new_new_n49_), .Y(new_new_n310_));
  NO2        g288(.A(i_2_), .B(i_12_), .Y(new_new_n311_));
  NA3        g289(.A(new_new_n280_), .B(new_new_n44_), .C(new_new_n125_), .Y(new_new_n312_));
  NA3        g290(.A(new_new_n312_), .B(new_new_n310_), .C(new_new_n307_), .Y(new_new_n313_));
  OR4        g291(.A(new_new_n313_), .B(new_new_n302_), .C(new_new_n299_), .D(new_new_n272_), .Y(mai5));
  NA2        g292(.A(new_new_n298_), .B(new_new_n143_), .Y(new_new_n315_));
  AN2        g293(.A(new_new_n24_), .B(i_10_), .Y(new_new_n316_));
  NA2        g294(.A(new_new_n316_), .B(new_new_n311_), .Y(new_new_n317_));
  NO2        g295(.A(new_new_n268_), .B(i_11_), .Y(new_new_n318_));
  NA2        g296(.A(new_new_n63_), .B(new_new_n318_), .Y(new_new_n319_));
  NA3        g297(.A(new_new_n319_), .B(new_new_n317_), .C(new_new_n315_), .Y(new_new_n320_));
  NO3        g298(.A(i_11_), .B(new_new_n130_), .C(i_13_), .Y(new_new_n321_));
  NO2        g299(.A(new_new_n77_), .B(new_new_n23_), .Y(new_new_n322_));
  INV        g300(.A(new_new_n203_), .Y(new_new_n323_));
  NA2        g301(.A(i_12_), .B(new_new_n322_), .Y(new_new_n324_));
  INV        g302(.A(new_new_n324_), .Y(new_new_n325_));
  NO2        g303(.A(new_new_n325_), .B(new_new_n320_), .Y(new_new_n326_));
  INV        g304(.A(new_new_n100_), .Y(new_new_n327_));
  OAI210     g305(.A0(i_4_), .A1(new_new_n204_), .B0(new_new_n71_), .Y(new_new_n328_));
  NO2        g306(.A(new_new_n328_), .B(new_new_n327_), .Y(new_new_n329_));
  AOI210     g307(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n198_), .Y(new_new_n330_));
  AOI210     g308(.A0(new_new_n330_), .A1(i_2_), .B0(new_new_n329_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n107_), .B(new_new_n78_), .Y(new_new_n332_));
  OAI210     g310(.A0(new_new_n332_), .A1(new_new_n322_), .B0(i_2_), .Y(new_new_n333_));
  NO3        g311(.A(new_new_n274_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n334_));
  INV        g312(.A(new_new_n334_), .Y(new_new_n335_));
  AOI210     g313(.A0(new_new_n335_), .A1(new_new_n333_), .B0(new_new_n108_), .Y(new_new_n336_));
  OA210      g314(.A0(new_new_n275_), .A1(new_new_n79_), .B0(i_13_), .Y(new_new_n337_));
  INV        g315(.A(new_new_n113_), .Y(new_new_n338_));
  INV        g316(.A(new_new_n93_), .Y(new_new_n339_));
  AOI210     g317(.A0(new_new_n339_), .A1(new_new_n338_), .B0(new_new_n172_), .Y(new_new_n340_));
  AOI210     g318(.A0(new_new_n118_), .A1(new_new_n91_), .B0(new_new_n239_), .Y(new_new_n341_));
  NA2        g319(.A(new_new_n341_), .B(new_new_n199_), .Y(new_new_n342_));
  NO2        g320(.A(i_2_), .B(new_new_n43_), .Y(new_new_n343_));
  NA3        g321(.A(new_new_n153_), .B(new_new_n77_), .C(new_new_n41_), .Y(new_new_n344_));
  OAI210     g322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(new_new_n342_), .Y(new_new_n345_));
  NO4        g323(.A(new_new_n345_), .B(new_new_n340_), .C(new_new_n337_), .D(new_new_n336_), .Y(new_new_n346_));
  INV        g324(.A(new_new_n262_), .Y(new_new_n347_));
  NA2        g325(.A(new_new_n321_), .B(i_7_), .Y(new_new_n348_));
  NA2        g326(.A(new_new_n348_), .B(new_new_n347_), .Y(new_new_n349_));
  NO2        g327(.A(i_2_), .B(i_12_), .Y(new_new_n350_));
  NO2        g328(.A(new_new_n350_), .B(new_new_n79_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n351_), .B(new_new_n267_), .Y(new_new_n352_));
  AOI220     g330(.A0(new_new_n352_), .A1(new_new_n36_), .B0(new_new_n349_), .B1(new_new_n45_), .Y(new_new_n353_));
  NA4        g331(.A(new_new_n353_), .B(new_new_n346_), .C(new_new_n331_), .D(new_new_n326_), .Y(mai6));
  NO2        g332(.A(new_new_n123_), .B(i_11_), .Y(new_new_n355_));
  NO2        g333(.A(i_11_), .B(i_9_), .Y(new_new_n356_));
  NO2        g334(.A(new_new_n184_), .B(new_new_n158_), .Y(new_new_n357_));
  OR2        g335(.A(new_new_n357_), .B(i_12_), .Y(new_new_n358_));
  AOI220     g336(.A0(new_new_n109_), .A1(new_new_n356_), .B0(new_new_n173_), .B1(new_new_n54_), .Y(new_new_n359_));
  NA2        g337(.A(new_new_n430_), .B(new_new_n350_), .Y(new_new_n360_));
  AOI210     g338(.A0(new_new_n360_), .A1(new_new_n237_), .B0(new_new_n104_), .Y(new_new_n361_));
  INV        g339(.A(i_11_), .Y(new_new_n362_));
  NA2        g340(.A(new_new_n362_), .B(new_new_n184_), .Y(new_new_n363_));
  NAi32      g341(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n364_));
  AOI210     g342(.A0(i_11_), .A1(i_11_), .B0(new_new_n364_), .Y(new_new_n365_));
  NA2        g343(.A(i_4_), .B(new_new_n259_), .Y(new_new_n366_));
  NAi31      g344(.An(new_new_n365_), .B(new_new_n366_), .C(new_new_n363_), .Y(new_new_n367_));
  OR2        g345(.A(new_new_n367_), .B(new_new_n361_), .Y(new_new_n368_));
  NA3        g346(.A(new_new_n439_), .B(new_new_n137_), .C(i_7_), .Y(new_new_n369_));
  NA2        g347(.A(new_new_n433_), .B(new_new_n90_), .Y(new_new_n370_));
  OR2        g348(.A(new_new_n323_), .B(new_new_n36_), .Y(new_new_n371_));
  NA3        g349(.A(new_new_n371_), .B(new_new_n370_), .C(new_new_n369_), .Y(new_new_n372_));
  INV        g350(.A(new_new_n355_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n131_), .B(new_new_n90_), .Y(new_new_n374_));
  OAI210     g352(.A0(new_new_n187_), .A1(new_new_n116_), .B0(new_new_n51_), .Y(new_new_n375_));
  NA4        g353(.A(new_new_n375_), .B(new_new_n374_), .C(new_new_n373_), .D(new_new_n269_), .Y(new_new_n376_));
  NA3        g354(.A(new_new_n239_), .B(new_new_n223_), .C(new_new_n122_), .Y(new_new_n377_));
  AOI210     g355(.A0(new_new_n204_), .A1(new_new_n203_), .B0(new_new_n258_), .Y(new_new_n378_));
  INV        g356(.A(new_new_n194_), .Y(new_new_n379_));
  NA3        g357(.A(new_new_n379_), .B(new_new_n378_), .C(new_new_n377_), .Y(new_new_n380_));
  NO4        g358(.A(new_new_n380_), .B(new_new_n376_), .C(new_new_n372_), .D(new_new_n368_), .Y(new_new_n381_));
  NA4        g359(.A(new_new_n381_), .B(new_new_n359_), .C(new_new_n358_), .D(new_new_n177_), .Y(mai3));
  NA2        g360(.A(new_new_n170_), .B(new_new_n39_), .Y(new_new_n383_));
  NO2        g361(.A(new_new_n383_), .B(new_new_n46_), .Y(new_new_n384_));
  NOi21      g362(.An(i_5_), .B(i_9_), .Y(new_new_n385_));
  NA2        g363(.A(new_new_n385_), .B(new_new_n202_), .Y(new_new_n386_));
  INV        g364(.A(new_new_n384_), .Y(new_new_n387_));
  NO4        g365(.A(i_5_), .B(i_12_), .C(new_new_n198_), .D(new_new_n195_), .Y(new_new_n388_));
  NA2        g366(.A(new_new_n388_), .B(i_11_), .Y(new_new_n389_));
  NA2        g367(.A(new_new_n321_), .B(new_new_n158_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n390_), .B(new_new_n389_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n186_), .B(new_new_n102_), .Y(new_new_n392_));
  NA3        g370(.A(new_new_n392_), .B(new_new_n208_), .C(new_new_n97_), .Y(new_new_n393_));
  NO2        g371(.A(i_12_), .B(new_new_n386_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n394_), .B(new_new_n393_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n294_), .B(i_1_), .Y(new_new_n396_));
  NO2        g374(.A(i_6_), .B(new_new_n396_), .Y(new_new_n397_));
  NA2        g375(.A(new_new_n100_), .B(new_new_n70_), .Y(new_new_n398_));
  INV        g376(.A(new_new_n397_), .Y(new_new_n399_));
  NA2        g377(.A(new_new_n399_), .B(new_new_n395_), .Y(new_new_n400_));
  NO3        g378(.A(i_5_), .B(i_0_), .C(new_new_n24_), .Y(new_new_n401_));
  INV        g379(.A(new_new_n401_), .Y(new_new_n402_));
  NAi21      g380(.An(i_9_), .B(i_5_), .Y(new_new_n403_));
  NO2        g381(.A(new_new_n403_), .B(new_new_n189_), .Y(new_new_n404_));
  NA2        g382(.A(new_new_n404_), .B(new_new_n275_), .Y(new_new_n405_));
  OAI220     g383(.A0(new_new_n405_), .A1(new_new_n61_), .B0(new_new_n402_), .B1(new_new_n101_), .Y(new_new_n406_));
  NO2        g384(.A(new_new_n406_), .B(new_new_n240_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n407_), .B(new_new_n106_), .Y(new_new_n408_));
  NO3        g386(.A(new_new_n408_), .B(new_new_n400_), .C(new_new_n391_), .Y(new_new_n409_));
  NO2        g387(.A(i_12_), .B(new_new_n398_), .Y(new_new_n410_));
  INV        g388(.A(new_new_n158_), .Y(new_new_n411_));
  NO2        g389(.A(new_new_n99_), .B(new_new_n411_), .Y(new_new_n412_));
  NO3        g390(.A(new_new_n119_), .B(new_new_n179_), .C(i_0_), .Y(new_new_n413_));
  OAI210     g391(.A0(new_new_n413_), .A1(new_new_n57_), .B0(i_13_), .Y(new_new_n414_));
  INV        g392(.A(new_new_n122_), .Y(new_new_n415_));
  NA3        g393(.A(new_new_n113_), .B(i_7_), .C(new_new_n415_), .Y(new_new_n416_));
  NA3        g394(.A(new_new_n416_), .B(new_new_n414_), .C(new_new_n429_), .Y(new_new_n417_));
  NA3        g395(.A(new_new_n184_), .B(new_new_n100_), .C(i_4_), .Y(new_new_n418_));
  NO3        g396(.A(new_new_n441_), .B(new_new_n417_), .C(new_new_n410_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n37_), .B(new_new_n117_), .Y(new_new_n420_));
  NO2        g398(.A(new_new_n420_), .B(new_new_n54_), .Y(new_new_n421_));
  INV        g399(.A(new_new_n258_), .Y(new_new_n422_));
  INV        g400(.A(new_new_n365_), .Y(new_new_n423_));
  AOI210     g401(.A0(new_new_n423_), .A1(new_new_n422_), .B0(new_new_n40_), .Y(new_new_n424_));
  NO2        g402(.A(new_new_n424_), .B(new_new_n421_), .Y(new_new_n425_));
  NA4        g403(.A(new_new_n425_), .B(new_new_n419_), .C(new_new_n409_), .D(new_new_n387_), .Y(mai4));
  INV        g404(.A(new_new_n412_), .Y(new_new_n429_));
  INV        g405(.A(i_9_), .Y(new_new_n430_));
  INV        g406(.A(new_new_n305_), .Y(new_new_n431_));
  INV        g407(.A(i_6_), .Y(new_new_n432_));
  INV        g408(.A(i_12_), .Y(new_new_n433_));
  INV        g409(.A(i_9_), .Y(new_new_n434_));
  INV        g410(.A(i_10_), .Y(new_new_n435_));
  INV        g411(.A(new_new_n57_), .Y(new_new_n436_));
  INV        g412(.A(new_new_n134_), .Y(new_new_n437_));
  INV        g413(.A(new_new_n263_), .Y(new_new_n438_));
  INV        g414(.A(i_9_), .Y(new_new_n439_));
  INV        g415(.A(i_2_), .Y(new_new_n440_));
  INV        g416(.A(new_new_n418_), .Y(new_new_n441_));
  INV        g417(.A(new_new_n26_), .Y(new_new_n442_));
endmodule


