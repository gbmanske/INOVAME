library verilog;
use verilog.vl_types.all;
entity ex_rca32bits_vlg_vec_tst is
end ex_rca32bits_vlg_vec_tst;
