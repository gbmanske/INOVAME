//Benchmark atmr_alu4_1266_0.0313

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n336_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n356_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n379_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n449_, ori_ori_n450_, ori_ori_n451_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, ori_ori_n455_, ori_ori_n456_, ori_ori_n457_, ori_ori_n458_, ori_ori_n459_, ori_ori_n460_, ori_ori_n461_, ori_ori_n462_, ori_ori_n463_, ori_ori_n464_, ori_ori_n465_, ori_ori_n466_, ori_ori_n467_, ori_ori_n468_, ori_ori_n469_, ori_ori_n470_, ori_ori_n471_, ori_ori_n472_, ori_ori_n473_, ori_ori_n474_, ori_ori_n475_, ori_ori_n476_, ori_ori_n477_, ori_ori_n478_, ori_ori_n479_, ori_ori_n480_, ori_ori_n481_, ori_ori_n482_, ori_ori_n483_, ori_ori_n484_, ori_ori_n485_, ori_ori_n486_, ori_ori_n487_, ori_ori_n488_, ori_ori_n489_, ori_ori_n490_, ori_ori_n491_, ori_ori_n492_, ori_ori_n493_, ori_ori_n494_, ori_ori_n495_, ori_ori_n496_, ori_ori_n497_, ori_ori_n498_, ori_ori_n499_, ori_ori_n500_, ori_ori_n501_, ori_ori_n502_, ori_ori_n503_, ori_ori_n504_, ori_ori_n505_, ori_ori_n506_, ori_ori_n507_, ori_ori_n508_, ori_ori_n509_, ori_ori_n510_, ori_ori_n511_, ori_ori_n512_, ori_ori_n513_, ori_ori_n514_, ori_ori_n515_, ori_ori_n516_, ori_ori_n517_, ori_ori_n518_, ori_ori_n519_, ori_ori_n520_, ori_ori_n521_, ori_ori_n522_, ori_ori_n523_, ori_ori_n524_, ori_ori_n525_, ori_ori_n526_, ori_ori_n527_, ori_ori_n528_, ori_ori_n529_, ori_ori_n530_, ori_ori_n531_, ori_ori_n532_, ori_ori_n533_, ori_ori_n534_, ori_ori_n535_, ori_ori_n536_, ori_ori_n537_, ori_ori_n538_, ori_ori_n539_, ori_ori_n540_, ori_ori_n541_, ori_ori_n542_, ori_ori_n543_, ori_ori_n544_, ori_ori_n545_, ori_ori_n546_, ori_ori_n547_, ori_ori_n548_, ori_ori_n549_, ori_ori_n551_, ori_ori_n552_, ori_ori_n553_, ori_ori_n554_, ori_ori_n555_, ori_ori_n556_, ori_ori_n557_, ori_ori_n558_, ori_ori_n559_, ori_ori_n560_, ori_ori_n561_, ori_ori_n562_, ori_ori_n563_, ori_ori_n564_, ori_ori_n565_, ori_ori_n566_, ori_ori_n567_, ori_ori_n568_, ori_ori_n569_, ori_ori_n570_, ori_ori_n571_, ori_ori_n572_, ori_ori_n573_, ori_ori_n574_, ori_ori_n575_, ori_ori_n576_, ori_ori_n577_, ori_ori_n578_, ori_ori_n579_, ori_ori_n580_, ori_ori_n581_, ori_ori_n582_, ori_ori_n583_, ori_ori_n584_, ori_ori_n585_, ori_ori_n586_, ori_ori_n587_, ori_ori_n588_, ori_ori_n589_, ori_ori_n590_, ori_ori_n591_, ori_ori_n592_, ori_ori_n593_, ori_ori_n594_, ori_ori_n595_, ori_ori_n596_, ori_ori_n597_, ori_ori_n598_, ori_ori_n599_, ori_ori_n600_, ori_ori_n601_, ori_ori_n602_, ori_ori_n603_, ori_ori_n604_, ori_ori_n605_, ori_ori_n606_, ori_ori_n607_, ori_ori_n608_, ori_ori_n609_, ori_ori_n610_, ori_ori_n611_, ori_ori_n612_, ori_ori_n613_, ori_ori_n614_, ori_ori_n615_, ori_ori_n616_, ori_ori_n617_, ori_ori_n618_, ori_ori_n619_, ori_ori_n620_, ori_ori_n621_, ori_ori_n622_, ori_ori_n623_, ori_ori_n624_, ori_ori_n625_, ori_ori_n626_, ori_ori_n627_, ori_ori_n628_, ori_ori_n629_, ori_ori_n630_, ori_ori_n631_, ori_ori_n632_, ori_ori_n633_, ori_ori_n634_, ori_ori_n635_, ori_ori_n636_, ori_ori_n637_, ori_ori_n638_, ori_ori_n639_, ori_ori_n640_, ori_ori_n641_, ori_ori_n642_, ori_ori_n643_, ori_ori_n644_, ori_ori_n645_, ori_ori_n646_, ori_ori_n647_, ori_ori_n648_, ori_ori_n649_, ori_ori_n650_, ori_ori_n651_, ori_ori_n652_, ori_ori_n653_, ori_ori_n654_, ori_ori_n655_, ori_ori_n656_, ori_ori_n657_, ori_ori_n658_, ori_ori_n659_, ori_ori_n660_, ori_ori_n661_, ori_ori_n662_, ori_ori_n663_, ori_ori_n664_, ori_ori_n665_, ori_ori_n666_, ori_ori_n667_, ori_ori_n668_, ori_ori_n669_, ori_ori_n670_, ori_ori_n671_, ori_ori_n672_, ori_ori_n673_, ori_ori_n674_, ori_ori_n675_, ori_ori_n676_, ori_ori_n677_, ori_ori_n678_, ori_ori_n679_, ori_ori_n680_, ori_ori_n681_, ori_ori_n682_, ori_ori_n683_, ori_ori_n684_, ori_ori_n685_, ori_ori_n686_, ori_ori_n687_, ori_ori_n688_, ori_ori_n689_, ori_ori_n690_, ori_ori_n691_, ori_ori_n692_, ori_ori_n694_, ori_ori_n695_, ori_ori_n696_, ori_ori_n697_, ori_ori_n698_, ori_ori_n699_, ori_ori_n700_, ori_ori_n701_, ori_ori_n702_, ori_ori_n703_, ori_ori_n704_, ori_ori_n705_, ori_ori_n706_, ori_ori_n707_, ori_ori_n708_, ori_ori_n709_, ori_ori_n710_, ori_ori_n711_, ori_ori_n712_, ori_ori_n713_, ori_ori_n714_, ori_ori_n715_, ori_ori_n716_, ori_ori_n717_, ori_ori_n718_, ori_ori_n719_, ori_ori_n720_, ori_ori_n721_, ori_ori_n722_, ori_ori_n723_, ori_ori_n724_, ori_ori_n725_, ori_ori_n726_, ori_ori_n727_, ori_ori_n728_, ori_ori_n729_, ori_ori_n730_, ori_ori_n731_, ori_ori_n732_, ori_ori_n733_, ori_ori_n734_, ori_ori_n735_, ori_ori_n736_, ori_ori_n737_, ori_ori_n738_, ori_ori_n739_, ori_ori_n740_, ori_ori_n741_, ori_ori_n743_, ori_ori_n744_, ori_ori_n745_, ori_ori_n746_, ori_ori_n747_, ori_ori_n748_, ori_ori_n749_, ori_ori_n750_, ori_ori_n751_, ori_ori_n752_, ori_ori_n753_, ori_ori_n754_, ori_ori_n755_, ori_ori_n756_, ori_ori_n757_, ori_ori_n758_, ori_ori_n759_, ori_ori_n760_, ori_ori_n761_, ori_ori_n762_, ori_ori_n763_, ori_ori_n764_, ori_ori_n765_, ori_ori_n766_, ori_ori_n767_, ori_ori_n768_, ori_ori_n769_, ori_ori_n770_, ori_ori_n771_, ori_ori_n772_, ori_ori_n773_, ori_ori_n774_, ori_ori_n775_, ori_ori_n776_, ori_ori_n777_, ori_ori_n778_, ori_ori_n779_, ori_ori_n780_, ori_ori_n781_, ori_ori_n782_, ori_ori_n783_, ori_ori_n784_, ori_ori_n785_, ori_ori_n786_, ori_ori_n787_, ori_ori_n788_, ori_ori_n789_, ori_ori_n790_, ori_ori_n792_, ori_ori_n793_, ori_ori_n794_, ori_ori_n795_, ori_ori_n796_, ori_ori_n797_, ori_ori_n798_, ori_ori_n799_, ori_ori_n800_, ori_ori_n801_, ori_ori_n802_, ori_ori_n803_, ori_ori_n804_, ori_ori_n805_, ori_ori_n806_, ori_ori_n807_, ori_ori_n808_, ori_ori_n809_, ori_ori_n810_, ori_ori_n811_, ori_ori_n812_, ori_ori_n813_, ori_ori_n814_, ori_ori_n815_, ori_ori_n816_, ori_ori_n817_, ori_ori_n818_, ori_ori_n819_, ori_ori_n820_, ori_ori_n821_, ori_ori_n822_, ori_ori_n823_, ori_ori_n824_, ori_ori_n825_, ori_ori_n826_, ori_ori_n827_, ori_ori_n828_, ori_ori_n829_, ori_ori_n830_, ori_ori_n831_, ori_ori_n832_, ori_ori_n833_, ori_ori_n834_, ori_ori_n835_, ori_ori_n836_, ori_ori_n837_, ori_ori_n838_, ori_ori_n839_, ori_ori_n840_, ori_ori_n841_, ori_ori_n842_, ori_ori_n843_, ori_ori_n844_, ori_ori_n845_, ori_ori_n846_, ori_ori_n847_, ori_ori_n848_, ori_ori_n849_, ori_ori_n850_, ori_ori_n851_, ori_ori_n852_, ori_ori_n853_, ori_ori_n854_, ori_ori_n855_, ori_ori_n856_, ori_ori_n857_, ori_ori_n858_, ori_ori_n859_, ori_ori_n860_, ori_ori_n861_, ori_ori_n862_, ori_ori_n863_, ori_ori_n864_, ori_ori_n865_, ori_ori_n866_, ori_ori_n867_, ori_ori_n868_, ori_ori_n869_, ori_ori_n870_, ori_ori_n871_, ori_ori_n872_, ori_ori_n873_, ori_ori_n874_, ori_ori_n875_, ori_ori_n876_, ori_ori_n877_, ori_ori_n878_, ori_ori_n879_, ori_ori_n880_, ori_ori_n881_, ori_ori_n882_, ori_ori_n883_, ori_ori_n884_, ori_ori_n885_, ori_ori_n886_, ori_ori_n887_, ori_ori_n888_, ori_ori_n889_, ori_ori_n890_, ori_ori_n891_, ori_ori_n892_, ori_ori_n893_, ori_ori_n894_, ori_ori_n895_, ori_ori_n896_, ori_ori_n897_, ori_ori_n898_, ori_ori_n899_, ori_ori_n900_, ori_ori_n901_, ori_ori_n902_, ori_ori_n903_, ori_ori_n904_, ori_ori_n905_, ori_ori_n906_, ori_ori_n907_, ori_ori_n908_, ori_ori_n909_, ori_ori_n910_, ori_ori_n911_, ori_ori_n912_, ori_ori_n913_, ori_ori_n914_, ori_ori_n915_, ori_ori_n916_, ori_ori_n917_, ori_ori_n918_, ori_ori_n919_, ori_ori_n920_, ori_ori_n921_, ori_ori_n922_, ori_ori_n923_, ori_ori_n924_, ori_ori_n925_, ori_ori_n926_, ori_ori_n927_, ori_ori_n928_, ori_ori_n929_, ori_ori_n930_, ori_ori_n931_, ori_ori_n932_, ori_ori_n933_, ori_ori_n934_, ori_ori_n935_, ori_ori_n936_, ori_ori_n937_, ori_ori_n938_, ori_ori_n939_, ori_ori_n940_, ori_ori_n941_, ori_ori_n942_, ori_ori_n943_, ori_ori_n944_, ori_ori_n945_, ori_ori_n946_, ori_ori_n947_, ori_ori_n948_, ori_ori_n949_, ori_ori_n950_, ori_ori_n951_, ori_ori_n952_, ori_ori_n953_, ori_ori_n954_, ori_ori_n955_, ori_ori_n956_, ori_ori_n957_, ori_ori_n961_, ori_ori_n962_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n509_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n639_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n678_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n723_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n898_, mai_mai_n899_, mai_mai_n900_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, mai_mai_n918_, mai_mai_n919_, mai_mai_n920_, mai_mai_n921_, mai_mai_n922_, mai_mai_n923_, mai_mai_n924_, mai_mai_n925_, mai_mai_n926_, mai_mai_n927_, mai_mai_n928_, mai_mai_n929_, mai_mai_n930_, mai_mai_n931_, mai_mai_n932_, mai_mai_n933_, mai_mai_n934_, mai_mai_n935_, mai_mai_n936_, mai_mai_n937_, mai_mai_n938_, mai_mai_n939_, mai_mai_n940_, mai_mai_n941_, mai_mai_n942_, mai_mai_n943_, mai_mai_n944_, mai_mai_n945_, mai_mai_n946_, mai_mai_n947_, mai_mai_n948_, mai_mai_n949_, mai_mai_n950_, mai_mai_n951_, mai_mai_n952_, mai_mai_n953_, mai_mai_n954_, mai_mai_n955_, mai_mai_n956_, mai_mai_n957_, mai_mai_n958_, mai_mai_n959_, mai_mai_n960_, mai_mai_n961_, mai_mai_n962_, mai_mai_n963_, mai_mai_n964_, mai_mai_n965_, mai_mai_n966_, mai_mai_n967_, mai_mai_n968_, mai_mai_n969_, mai_mai_n970_, mai_mai_n971_, mai_mai_n972_, mai_mai_n973_, mai_mai_n974_, mai_mai_n975_, mai_mai_n976_, mai_mai_n977_, mai_mai_n978_, mai_mai_n979_, mai_mai_n980_, mai_mai_n981_, mai_mai_n982_, mai_mai_n983_, mai_mai_n984_, mai_mai_n985_, mai_mai_n986_, mai_mai_n987_, mai_mai_n988_, mai_mai_n989_, mai_mai_n990_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n588_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n708_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n747_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n786_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1007_, men_men_n1008_, men_men_n1009_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, men_men_n1023_, men_men_n1024_, men_men_n1025_, men_men_n1026_, men_men_n1027_, men_men_n1028_, men_men_n1029_, men_men_n1030_, men_men_n1031_, men_men_n1032_, men_men_n1033_, men_men_n1034_, men_men_n1035_, men_men_n1036_, men_men_n1037_, men_men_n1038_, men_men_n1042_, men_men_n1043_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  NOi21      o008(.An(i_11_), .B(i_8_), .Y(ori_ori_n31_));
  AO210      o009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n32_));
  OR2        o010(.A(ori_ori_n32_), .B(ori_ori_n31_), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n30_), .Y(ori_ori_n34_));
  XO2        o012(.A(ori_ori_n34_), .B(ori_ori_n23_), .Y(ori_ori_n35_));
  INV        o013(.A(i_4_), .Y(ori_ori_n36_));
  INV        o014(.A(i_10_), .Y(ori_ori_n37_));
  NAi21      o015(.An(i_11_), .B(i_9_), .Y(ori_ori_n38_));
  NO3        o016(.A(ori_ori_n38_), .B(i_12_), .C(ori_ori_n37_), .Y(ori_ori_n39_));
  NOi21      o017(.An(i_12_), .B(i_13_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n40_), .Y(ori_ori_n41_));
  NAi31      o019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(ori_ori_n42_));
  INV        o020(.A(ori_ori_n35_), .Y(ori1));
  INV        o021(.A(i_11_), .Y(ori_ori_n44_));
  NO2        o022(.A(ori_ori_n44_), .B(i_6_), .Y(ori_ori_n45_));
  INV        o023(.A(i_2_), .Y(ori_ori_n46_));
  NA2        o024(.A(i_0_), .B(i_3_), .Y(ori_ori_n47_));
  INV        o025(.A(i_5_), .Y(ori_ori_n48_));
  NO2        o026(.A(i_7_), .B(i_10_), .Y(ori_ori_n49_));
  AOI210     o027(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n49_), .Y(ori_ori_n50_));
  OAI210     o028(.A0(ori_ori_n50_), .A1(i_3_), .B0(ori_ori_n48_), .Y(ori_ori_n51_));
  AOI210     o029(.A0(ori_ori_n51_), .A1(ori_ori_n47_), .B0(ori_ori_n46_), .Y(ori_ori_n52_));
  NA2        o030(.A(i_0_), .B(i_2_), .Y(ori_ori_n53_));
  NA2        o031(.A(i_7_), .B(i_9_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n53_), .Y(ori_ori_n55_));
  NA2        o033(.A(ori_ori_n52_), .B(ori_ori_n45_), .Y(ori_ori_n56_));
  NO2        o034(.A(i_1_), .B(i_6_), .Y(ori_ori_n57_));
  NA2        o035(.A(i_8_), .B(i_7_), .Y(ori_ori_n58_));
  NO2        o036(.A(ori_ori_n58_), .B(ori_ori_n57_), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(i_12_), .Y(ori_ori_n60_));
  NAi21      o038(.An(i_2_), .B(i_7_), .Y(ori_ori_n61_));
  INV        o039(.A(i_1_), .Y(ori_ori_n62_));
  NA2        o040(.A(ori_ori_n62_), .B(i_6_), .Y(ori_ori_n63_));
  NA3        o041(.A(ori_ori_n63_), .B(ori_ori_n61_), .C(ori_ori_n31_), .Y(ori_ori_n64_));
  NA2        o042(.A(i_1_), .B(i_10_), .Y(ori_ori_n65_));
  NO2        o043(.A(ori_ori_n65_), .B(i_6_), .Y(ori_ori_n66_));
  NAi31      o044(.An(ori_ori_n66_), .B(ori_ori_n64_), .C(ori_ori_n60_), .Y(ori_ori_n67_));
  NA2        o045(.A(ori_ori_n50_), .B(i_2_), .Y(ori_ori_n68_));
  AOI210     o046(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n69_));
  NA2        o047(.A(i_1_), .B(i_6_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n70_), .B(ori_ori_n25_), .Y(ori_ori_n71_));
  INV        o049(.A(i_0_), .Y(ori_ori_n72_));
  NAi21      o050(.An(i_5_), .B(i_10_), .Y(ori_ori_n73_));
  NA2        o051(.A(i_5_), .B(i_9_), .Y(ori_ori_n74_));
  AOI210     o052(.A0(ori_ori_n74_), .A1(ori_ori_n73_), .B0(ori_ori_n72_), .Y(ori_ori_n75_));
  NO2        o053(.A(ori_ori_n75_), .B(ori_ori_n71_), .Y(ori_ori_n76_));
  OAI210     o054(.A0(ori_ori_n69_), .A1(ori_ori_n68_), .B0(ori_ori_n76_), .Y(ori_ori_n77_));
  OAI210     o055(.A0(ori_ori_n77_), .A1(ori_ori_n67_), .B0(i_0_), .Y(ori_ori_n78_));
  NA2        o056(.A(i_12_), .B(i_5_), .Y(ori_ori_n79_));
  NA2        o057(.A(i_2_), .B(i_8_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(ori_ori_n57_), .Y(ori_ori_n81_));
  NO2        o059(.A(i_3_), .B(i_9_), .Y(ori_ori_n82_));
  NO2        o060(.A(i_3_), .B(i_7_), .Y(ori_ori_n83_));
  NO2        o061(.A(ori_ori_n82_), .B(ori_ori_n62_), .Y(ori_ori_n84_));
  INV        o062(.A(i_6_), .Y(ori_ori_n85_));
  NO2        o063(.A(i_2_), .B(i_7_), .Y(ori_ori_n86_));
  INV        o064(.A(ori_ori_n86_), .Y(ori_ori_n87_));
  OAI210     o065(.A0(ori_ori_n84_), .A1(ori_ori_n81_), .B0(ori_ori_n87_), .Y(ori_ori_n88_));
  NAi21      o066(.An(i_6_), .B(i_10_), .Y(ori_ori_n89_));
  NA2        o067(.A(i_6_), .B(i_9_), .Y(ori_ori_n90_));
  AOI210     o068(.A0(ori_ori_n90_), .A1(ori_ori_n89_), .B0(ori_ori_n62_), .Y(ori_ori_n91_));
  NA2        o069(.A(i_2_), .B(i_6_), .Y(ori_ori_n92_));
  NO3        o070(.A(ori_ori_n92_), .B(ori_ori_n49_), .C(ori_ori_n25_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(ori_ori_n91_), .Y(ori_ori_n94_));
  AOI210     o072(.A0(ori_ori_n94_), .A1(ori_ori_n88_), .B0(ori_ori_n79_), .Y(ori_ori_n95_));
  AN3        o073(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n96_));
  NAi21      o074(.An(i_6_), .B(i_11_), .Y(ori_ori_n97_));
  NO2        o075(.A(i_5_), .B(i_8_), .Y(ori_ori_n98_));
  NOi21      o076(.An(ori_ori_n98_), .B(ori_ori_n97_), .Y(ori_ori_n99_));
  AOI220     o077(.A0(ori_ori_n99_), .A1(ori_ori_n61_), .B0(ori_ori_n96_), .B1(ori_ori_n32_), .Y(ori_ori_n100_));
  INV        o078(.A(i_7_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n46_), .B(ori_ori_n101_), .Y(ori_ori_n102_));
  NO2        o080(.A(i_0_), .B(i_5_), .Y(ori_ori_n103_));
  NO2        o081(.A(ori_ori_n103_), .B(ori_ori_n85_), .Y(ori_ori_n104_));
  NA2        o082(.A(i_12_), .B(i_3_), .Y(ori_ori_n105_));
  INV        o083(.A(ori_ori_n105_), .Y(ori_ori_n106_));
  NA3        o084(.A(ori_ori_n106_), .B(ori_ori_n104_), .C(ori_ori_n102_), .Y(ori_ori_n107_));
  NAi21      o085(.An(i_7_), .B(i_11_), .Y(ori_ori_n108_));
  NO3        o086(.A(ori_ori_n108_), .B(ori_ori_n89_), .C(ori_ori_n53_), .Y(ori_ori_n109_));
  AN2        o087(.A(i_2_), .B(i_10_), .Y(ori_ori_n110_));
  NO2        o088(.A(ori_ori_n110_), .B(i_7_), .Y(ori_ori_n111_));
  OR2        o089(.A(ori_ori_n79_), .B(ori_ori_n57_), .Y(ori_ori_n112_));
  NO2        o090(.A(i_8_), .B(ori_ori_n101_), .Y(ori_ori_n113_));
  NO3        o091(.A(ori_ori_n113_), .B(ori_ori_n112_), .C(ori_ori_n111_), .Y(ori_ori_n114_));
  NA2        o092(.A(i_12_), .B(i_7_), .Y(ori_ori_n115_));
  NO2        o093(.A(ori_ori_n62_), .B(ori_ori_n26_), .Y(ori_ori_n116_));
  NA2        o094(.A(ori_ori_n116_), .B(i_0_), .Y(ori_ori_n117_));
  NA2        o095(.A(i_11_), .B(i_12_), .Y(ori_ori_n118_));
  OAI210     o096(.A0(ori_ori_n117_), .A1(ori_ori_n115_), .B0(ori_ori_n118_), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n119_), .B(ori_ori_n114_), .Y(ori_ori_n120_));
  NAi41      o098(.An(ori_ori_n109_), .B(ori_ori_n120_), .C(ori_ori_n107_), .D(ori_ori_n100_), .Y(ori_ori_n121_));
  NOi21      o099(.An(i_1_), .B(i_5_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n122_), .B(i_11_), .Y(ori_ori_n123_));
  NA2        o101(.A(ori_ori_n101_), .B(ori_ori_n37_), .Y(ori_ori_n124_));
  NA2        o102(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n125_));
  NA2        o103(.A(ori_ori_n125_), .B(ori_ori_n124_), .Y(ori_ori_n126_));
  NO2        o104(.A(ori_ori_n126_), .B(ori_ori_n46_), .Y(ori_ori_n127_));
  NA2        o105(.A(ori_ori_n90_), .B(ori_ori_n89_), .Y(ori_ori_n128_));
  NAi21      o106(.An(i_3_), .B(i_8_), .Y(ori_ori_n129_));
  NA2        o107(.A(ori_ori_n129_), .B(ori_ori_n61_), .Y(ori_ori_n130_));
  NOi31      o108(.An(ori_ori_n130_), .B(ori_ori_n128_), .C(ori_ori_n127_), .Y(ori_ori_n131_));
  NO2        o109(.A(i_1_), .B(ori_ori_n85_), .Y(ori_ori_n132_));
  NO2        o110(.A(i_6_), .B(i_5_), .Y(ori_ori_n133_));
  NA2        o111(.A(ori_ori_n133_), .B(i_3_), .Y(ori_ori_n134_));
  AO210      o112(.A0(ori_ori_n134_), .A1(ori_ori_n47_), .B0(ori_ori_n132_), .Y(ori_ori_n135_));
  OAI220     o113(.A0(ori_ori_n135_), .A1(ori_ori_n108_), .B0(ori_ori_n131_), .B1(ori_ori_n123_), .Y(ori_ori_n136_));
  NO3        o114(.A(ori_ori_n136_), .B(ori_ori_n121_), .C(ori_ori_n95_), .Y(ori_ori_n137_));
  NA3        o115(.A(ori_ori_n137_), .B(ori_ori_n78_), .C(ori_ori_n56_), .Y(ori2));
  NO2        o116(.A(ori_ori_n62_), .B(ori_ori_n37_), .Y(ori_ori_n139_));
  NA2        o117(.A(i_6_), .B(ori_ori_n25_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n140_), .B(ori_ori_n139_), .Y(ori_ori_n141_));
  NA4        o119(.A(ori_ori_n141_), .B(ori_ori_n76_), .C(ori_ori_n68_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o120(.A(i_8_), .B(i_7_), .Y(ori_ori_n143_));
  NA2        o121(.A(ori_ori_n143_), .B(i_6_), .Y(ori_ori_n144_));
  NO2        o122(.A(i_12_), .B(i_13_), .Y(ori_ori_n145_));
  NAi21      o123(.An(i_5_), .B(i_11_), .Y(ori_ori_n146_));
  NOi21      o124(.An(ori_ori_n145_), .B(ori_ori_n146_), .Y(ori_ori_n147_));
  NO2        o125(.A(i_0_), .B(i_1_), .Y(ori_ori_n148_));
  NA2        o126(.A(i_2_), .B(i_3_), .Y(ori_ori_n149_));
  NO2        o127(.A(ori_ori_n149_), .B(i_4_), .Y(ori_ori_n150_));
  NA3        o128(.A(ori_ori_n150_), .B(ori_ori_n148_), .C(ori_ori_n147_), .Y(ori_ori_n151_));
  AN2        o129(.A(ori_ori_n145_), .B(ori_ori_n82_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n152_), .B(ori_ori_n27_), .Y(ori_ori_n153_));
  NA2        o131(.A(i_1_), .B(i_5_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n72_), .B(ori_ori_n46_), .Y(ori_ori_n155_));
  NA2        o133(.A(ori_ori_n155_), .B(ori_ori_n36_), .Y(ori_ori_n156_));
  NO3        o134(.A(ori_ori_n156_), .B(ori_ori_n154_), .C(ori_ori_n153_), .Y(ori_ori_n157_));
  OR2        o135(.A(i_0_), .B(i_1_), .Y(ori_ori_n158_));
  NO3        o136(.A(ori_ori_n158_), .B(ori_ori_n79_), .C(i_13_), .Y(ori_ori_n159_));
  NAi32      o137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(ori_ori_n160_));
  NAi21      o138(.An(ori_ori_n160_), .B(ori_ori_n159_), .Y(ori_ori_n161_));
  NOi21      o139(.An(i_4_), .B(i_10_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n162_), .B(ori_ori_n40_), .Y(ori_ori_n163_));
  NO2        o141(.A(i_3_), .B(i_5_), .Y(ori_ori_n164_));
  NO3        o142(.A(ori_ori_n72_), .B(i_2_), .C(i_1_), .Y(ori_ori_n165_));
  NA2        o143(.A(ori_ori_n165_), .B(ori_ori_n164_), .Y(ori_ori_n166_));
  OAI210     o144(.A0(ori_ori_n166_), .A1(ori_ori_n163_), .B0(ori_ori_n161_), .Y(ori_ori_n167_));
  NO2        o145(.A(ori_ori_n167_), .B(ori_ori_n157_), .Y(ori_ori_n168_));
  NO2        o146(.A(ori_ori_n168_), .B(ori_ori_n144_), .Y(ori_ori_n169_));
  NOi21      o147(.An(i_4_), .B(i_9_), .Y(ori_ori_n170_));
  NOi21      o148(.An(i_11_), .B(i_13_), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n171_), .B(ori_ori_n170_), .Y(ori_ori_n172_));
  NO2        o150(.A(i_4_), .B(i_5_), .Y(ori_ori_n173_));
  NAi21      o151(.An(i_12_), .B(i_11_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n72_), .B(ori_ori_n62_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n46_), .Y(ori_ori_n176_));
  NAi31      o154(.An(i_4_), .B(ori_ori_n152_), .C(i_11_), .Y(ori_ori_n177_));
  NA2        o155(.A(i_3_), .B(i_5_), .Y(ori_ori_n178_));
  OR2        o156(.A(ori_ori_n178_), .B(ori_ori_n172_), .Y(ori_ori_n179_));
  AOI210     o157(.A0(ori_ori_n179_), .A1(ori_ori_n177_), .B0(ori_ori_n176_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n181_));
  NO2        o159(.A(i_13_), .B(i_10_), .Y(ori_ori_n182_));
  NA3        o160(.A(ori_ori_n182_), .B(ori_ori_n181_), .C(ori_ori_n44_), .Y(ori_ori_n183_));
  NO2        o161(.A(i_2_), .B(i_1_), .Y(ori_ori_n184_));
  NA2        o162(.A(ori_ori_n184_), .B(i_3_), .Y(ori_ori_n185_));
  NAi21      o163(.An(i_4_), .B(i_12_), .Y(ori_ori_n186_));
  INV        o164(.A(ori_ori_n180_), .Y(ori_ori_n187_));
  INV        o165(.A(i_8_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n188_), .B(i_7_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n189_), .B(i_6_), .Y(ori_ori_n190_));
  NO3        o168(.A(i_3_), .B(ori_ori_n85_), .C(ori_ori_n48_), .Y(ori_ori_n191_));
  NA2        o169(.A(ori_ori_n191_), .B(ori_ori_n113_), .Y(ori_ori_n192_));
  NO3        o170(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n193_));
  NA3        o171(.A(ori_ori_n193_), .B(ori_ori_n40_), .C(ori_ori_n44_), .Y(ori_ori_n194_));
  NO3        o172(.A(i_11_), .B(i_13_), .C(i_9_), .Y(ori_ori_n195_));
  OAI210     o173(.A0(ori_ori_n96_), .A1(i_12_), .B0(ori_ori_n195_), .Y(ori_ori_n196_));
  AOI210     o174(.A0(ori_ori_n196_), .A1(ori_ori_n194_), .B0(ori_ori_n192_), .Y(ori_ori_n197_));
  NO2        o175(.A(i_3_), .B(i_8_), .Y(ori_ori_n198_));
  NO3        o176(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n199_));
  NA3        o177(.A(ori_ori_n199_), .B(ori_ori_n198_), .C(ori_ori_n40_), .Y(ori_ori_n200_));
  NO2        o178(.A(ori_ori_n103_), .B(ori_ori_n57_), .Y(ori_ori_n201_));
  INV        o179(.A(ori_ori_n201_), .Y(ori_ori_n202_));
  NO2        o180(.A(i_13_), .B(i_9_), .Y(ori_ori_n203_));
  NAi21      o181(.An(i_12_), .B(i_3_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n44_), .B(i_5_), .Y(ori_ori_n205_));
  NO3        o183(.A(i_0_), .B(i_2_), .C(ori_ori_n62_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n202_), .B(ori_ori_n200_), .Y(ori_ori_n207_));
  AOI210     o185(.A0(ori_ori_n207_), .A1(i_7_), .B0(ori_ori_n197_), .Y(ori_ori_n208_));
  OAI220     o186(.A0(ori_ori_n208_), .A1(i_4_), .B0(ori_ori_n190_), .B1(ori_ori_n187_), .Y(ori_ori_n209_));
  NAi21      o187(.An(i_12_), .B(i_7_), .Y(ori_ori_n210_));
  NA3        o188(.A(i_13_), .B(ori_ori_n188_), .C(i_10_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(ori_ori_n210_), .Y(ori_ori_n212_));
  NA2        o190(.A(i_0_), .B(i_5_), .Y(ori_ori_n213_));
  NA2        o191(.A(ori_ori_n213_), .B(ori_ori_n104_), .Y(ori_ori_n214_));
  OAI220     o192(.A0(ori_ori_n214_), .A1(ori_ori_n185_), .B0(ori_ori_n176_), .B1(ori_ori_n134_), .Y(ori_ori_n215_));
  NAi31      o193(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n216_));
  NO2        o194(.A(ori_ori_n36_), .B(i_13_), .Y(ori_ori_n217_));
  NO2        o195(.A(ori_ori_n46_), .B(ori_ori_n62_), .Y(ori_ori_n218_));
  INV        o196(.A(i_13_), .Y(ori_ori_n219_));
  NO2        o197(.A(i_12_), .B(ori_ori_n219_), .Y(ori_ori_n220_));
  NA2        o198(.A(ori_ori_n215_), .B(ori_ori_n212_), .Y(ori_ori_n221_));
  NO2        o199(.A(i_12_), .B(ori_ori_n37_), .Y(ori_ori_n222_));
  NO2        o200(.A(ori_ori_n178_), .B(i_4_), .Y(ori_ori_n223_));
  NA2        o201(.A(ori_ori_n223_), .B(ori_ori_n222_), .Y(ori_ori_n224_));
  OR2        o202(.A(i_8_), .B(i_7_), .Y(ori_ori_n225_));
  NO2        o203(.A(ori_ori_n225_), .B(ori_ori_n85_), .Y(ori_ori_n226_));
  NO2        o204(.A(ori_ori_n53_), .B(i_1_), .Y(ori_ori_n227_));
  NA2        o205(.A(ori_ori_n227_), .B(ori_ori_n226_), .Y(ori_ori_n228_));
  INV        o206(.A(i_12_), .Y(ori_ori_n229_));
  NO2        o207(.A(ori_ori_n44_), .B(ori_ori_n229_), .Y(ori_ori_n230_));
  NO3        o208(.A(ori_ori_n36_), .B(i_8_), .C(i_10_), .Y(ori_ori_n231_));
  NA2        o209(.A(i_2_), .B(i_1_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n228_), .B(ori_ori_n224_), .Y(ori_ori_n233_));
  NO3        o211(.A(i_11_), .B(i_7_), .C(ori_ori_n37_), .Y(ori_ori_n234_));
  NAi21      o212(.An(i_4_), .B(i_3_), .Y(ori_ori_n235_));
  NO2        o213(.A(ori_ori_n235_), .B(ori_ori_n74_), .Y(ori_ori_n236_));
  NO2        o214(.A(i_0_), .B(i_6_), .Y(ori_ori_n237_));
  NOi41      o215(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n238_));
  NO2        o216(.A(ori_ori_n232_), .B(ori_ori_n178_), .Y(ori_ori_n239_));
  INV        o217(.A(ori_ori_n233_), .Y(ori_ori_n240_));
  NO2        o218(.A(i_11_), .B(ori_ori_n219_), .Y(ori_ori_n241_));
  NOi21      o219(.An(i_1_), .B(i_6_), .Y(ori_ori_n242_));
  NAi21      o220(.An(i_3_), .B(i_7_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n229_), .B(i_9_), .Y(ori_ori_n244_));
  NO2        o222(.A(i_12_), .B(i_3_), .Y(ori_ori_n245_));
  NA2        o223(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n246_));
  NA2        o224(.A(i_3_), .B(i_9_), .Y(ori_ori_n247_));
  NAi21      o225(.An(i_7_), .B(i_10_), .Y(ori_ori_n248_));
  NO2        o226(.A(ori_ori_n248_), .B(ori_ori_n247_), .Y(ori_ori_n249_));
  NA3        o227(.A(ori_ori_n249_), .B(ori_ori_n246_), .C(ori_ori_n63_), .Y(ori_ori_n250_));
  INV        o228(.A(ori_ori_n250_), .Y(ori_ori_n251_));
  INV        o229(.A(ori_ori_n144_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n229_), .B(i_13_), .Y(ori_ori_n253_));
  NO2        o231(.A(ori_ori_n253_), .B(ori_ori_n74_), .Y(ori_ori_n254_));
  AOI220     o232(.A0(ori_ori_n254_), .A1(ori_ori_n252_), .B0(ori_ori_n251_), .B1(ori_ori_n241_), .Y(ori_ori_n255_));
  NO2        o233(.A(ori_ori_n225_), .B(ori_ori_n37_), .Y(ori_ori_n256_));
  NA2        o234(.A(i_12_), .B(i_6_), .Y(ori_ori_n257_));
  OR2        o235(.A(i_13_), .B(i_9_), .Y(ori_ori_n258_));
  NO3        o236(.A(ori_ori_n258_), .B(ori_ori_n257_), .C(ori_ori_n48_), .Y(ori_ori_n259_));
  NO2        o237(.A(ori_ori_n235_), .B(i_2_), .Y(ori_ori_n260_));
  NA3        o238(.A(ori_ori_n260_), .B(ori_ori_n259_), .C(ori_ori_n44_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n241_), .B(i_9_), .Y(ori_ori_n262_));
  NA2        o240(.A(ori_ori_n246_), .B(ori_ori_n63_), .Y(ori_ori_n263_));
  OAI210     o241(.A0(ori_ori_n263_), .A1(ori_ori_n262_), .B0(ori_ori_n261_), .Y(ori_ori_n264_));
  NA2        o242(.A(ori_ori_n155_), .B(ori_ori_n62_), .Y(ori_ori_n265_));
  NO3        o243(.A(i_11_), .B(ori_ori_n219_), .C(ori_ori_n25_), .Y(ori_ori_n266_));
  NO2        o244(.A(ori_ori_n243_), .B(i_8_), .Y(ori_ori_n267_));
  NO2        o245(.A(i_6_), .B(ori_ori_n48_), .Y(ori_ori_n268_));
  NA3        o246(.A(ori_ori_n268_), .B(ori_ori_n267_), .C(ori_ori_n266_), .Y(ori_ori_n269_));
  NO3        o247(.A(ori_ori_n26_), .B(ori_ori_n85_), .C(i_5_), .Y(ori_ori_n270_));
  NA3        o248(.A(ori_ori_n270_), .B(ori_ori_n256_), .C(ori_ori_n220_), .Y(ori_ori_n271_));
  AOI210     o249(.A0(ori_ori_n271_), .A1(ori_ori_n269_), .B0(ori_ori_n265_), .Y(ori_ori_n272_));
  AOI210     o250(.A0(ori_ori_n264_), .A1(ori_ori_n256_), .B0(ori_ori_n272_), .Y(ori_ori_n273_));
  NA4        o251(.A(ori_ori_n273_), .B(ori_ori_n255_), .C(ori_ori_n240_), .D(ori_ori_n221_), .Y(ori_ori_n274_));
  NO3        o252(.A(i_12_), .B(ori_ori_n219_), .C(ori_ori_n37_), .Y(ori_ori_n275_));
  INV        o253(.A(ori_ori_n275_), .Y(ori_ori_n276_));
  NA2        o254(.A(i_8_), .B(ori_ori_n101_), .Y(ori_ori_n277_));
  NO3        o255(.A(i_0_), .B(ori_ori_n46_), .C(i_1_), .Y(ori_ori_n278_));
  AOI220     o256(.A0(ori_ori_n278_), .A1(ori_ori_n191_), .B0(ori_ori_n164_), .B1(ori_ori_n227_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n279_), .B(ori_ori_n277_), .Y(ori_ori_n280_));
  NO3        o258(.A(i_0_), .B(i_2_), .C(ori_ori_n62_), .Y(ori_ori_n281_));
  NO2        o259(.A(ori_ori_n232_), .B(i_0_), .Y(ori_ori_n282_));
  AOI220     o260(.A0(ori_ori_n282_), .A1(ori_ori_n189_), .B0(ori_ori_n281_), .B1(ori_ori_n143_), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n268_), .B(ori_ori_n26_), .Y(ori_ori_n284_));
  NO2        o262(.A(ori_ori_n284_), .B(ori_ori_n283_), .Y(ori_ori_n285_));
  NO2        o263(.A(ori_ori_n58_), .B(i_6_), .Y(ori_ori_n286_));
  NO2        o264(.A(ori_ori_n166_), .B(ori_ori_n144_), .Y(ori_ori_n287_));
  NO3        o265(.A(ori_ori_n287_), .B(ori_ori_n285_), .C(ori_ori_n280_), .Y(ori_ori_n288_));
  NO2        o266(.A(i_3_), .B(i_10_), .Y(ori_ori_n289_));
  NA3        o267(.A(ori_ori_n289_), .B(ori_ori_n40_), .C(ori_ori_n44_), .Y(ori_ori_n290_));
  NO2        o268(.A(i_2_), .B(ori_ori_n101_), .Y(ori_ori_n291_));
  NA2        o269(.A(i_1_), .B(ori_ori_n36_), .Y(ori_ori_n292_));
  AN2        o270(.A(i_3_), .B(i_10_), .Y(ori_ori_n293_));
  NO2        o271(.A(i_5_), .B(ori_ori_n37_), .Y(ori_ori_n294_));
  NO2        o272(.A(ori_ori_n46_), .B(ori_ori_n26_), .Y(ori_ori_n295_));
  NO2        o273(.A(ori_ori_n288_), .B(ori_ori_n276_), .Y(ori_ori_n296_));
  NO4        o274(.A(ori_ori_n296_), .B(ori_ori_n274_), .C(ori_ori_n209_), .D(ori_ori_n169_), .Y(ori_ori_n297_));
  NO3        o275(.A(ori_ori_n44_), .B(i_13_), .C(i_9_), .Y(ori_ori_n298_));
  NO3        o276(.A(i_6_), .B(ori_ori_n188_), .C(i_7_), .Y(ori_ori_n299_));
  NA2        o277(.A(ori_ori_n299_), .B(ori_ori_n193_), .Y(ori_ori_n300_));
  INV        o278(.A(ori_ori_n300_), .Y(ori_ori_n301_));
  NO2        o279(.A(i_2_), .B(i_3_), .Y(ori_ori_n302_));
  OR2        o280(.A(i_0_), .B(i_5_), .Y(ori_ori_n303_));
  NA2        o281(.A(ori_ori_n213_), .B(ori_ori_n303_), .Y(ori_ori_n304_));
  NA4        o282(.A(ori_ori_n304_), .B(ori_ori_n226_), .C(ori_ori_n302_), .D(i_1_), .Y(ori_ori_n305_));
  NA3        o283(.A(ori_ori_n282_), .B(ori_ori_n164_), .C(ori_ori_n113_), .Y(ori_ori_n306_));
  NAi21      o284(.An(i_8_), .B(i_7_), .Y(ori_ori_n307_));
  NO2        o285(.A(ori_ori_n158_), .B(ori_ori_n46_), .Y(ori_ori_n308_));
  NA2        o286(.A(ori_ori_n306_), .B(ori_ori_n305_), .Y(ori_ori_n309_));
  OAI210     o287(.A0(ori_ori_n309_), .A1(ori_ori_n301_), .B0(i_4_), .Y(ori_ori_n310_));
  NO2        o288(.A(i_12_), .B(i_10_), .Y(ori_ori_n311_));
  NOi21      o289(.An(i_5_), .B(i_0_), .Y(ori_ori_n312_));
  NO2        o290(.A(i_2_), .B(ori_ori_n101_), .Y(ori_ori_n313_));
  NO4        o291(.A(ori_ori_n313_), .B(ori_ori_n292_), .C(ori_ori_n312_), .D(ori_ori_n129_), .Y(ori_ori_n314_));
  NA4        o292(.A(ori_ori_n83_), .B(ori_ori_n36_), .C(ori_ori_n85_), .D(i_8_), .Y(ori_ori_n315_));
  NA2        o293(.A(ori_ori_n314_), .B(ori_ori_n311_), .Y(ori_ori_n316_));
  NO2        o294(.A(i_6_), .B(i_8_), .Y(ori_ori_n317_));
  NOi21      o295(.An(i_0_), .B(i_2_), .Y(ori_ori_n318_));
  AN2        o296(.A(ori_ori_n318_), .B(ori_ori_n317_), .Y(ori_ori_n319_));
  NO2        o297(.A(i_1_), .B(i_7_), .Y(ori_ori_n320_));
  NA2        o298(.A(ori_ori_n316_), .B(ori_ori_n310_), .Y(ori_ori_n321_));
  NO3        o299(.A(ori_ori_n225_), .B(ori_ori_n46_), .C(i_1_), .Y(ori_ori_n322_));
  NO3        o300(.A(ori_ori_n307_), .B(i_2_), .C(i_1_), .Y(ori_ori_n323_));
  OAI210     o301(.A0(ori_ori_n323_), .A1(ori_ori_n322_), .B0(i_6_), .Y(ori_ori_n324_));
  NA3        o302(.A(ori_ori_n242_), .B(ori_ori_n291_), .C(ori_ori_n188_), .Y(ori_ori_n325_));
  AOI210     o303(.A0(ori_ori_n325_), .A1(ori_ori_n324_), .B0(ori_ori_n304_), .Y(ori_ori_n326_));
  NOi21      o304(.An(ori_ori_n154_), .B(ori_ori_n104_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n327_), .B(ori_ori_n125_), .Y(ori_ori_n328_));
  OAI210     o306(.A0(ori_ori_n328_), .A1(ori_ori_n326_), .B0(i_3_), .Y(ori_ori_n329_));
  NO2        o307(.A(ori_ori_n188_), .B(i_9_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n330_), .B(ori_ori_n201_), .Y(ori_ori_n331_));
  NO2        o309(.A(ori_ori_n331_), .B(ori_ori_n46_), .Y(ori_ori_n332_));
  NO2        o310(.A(ori_ori_n332_), .B(ori_ori_n285_), .Y(ori_ori_n333_));
  AOI210     o311(.A0(ori_ori_n333_), .A1(ori_ori_n329_), .B0(ori_ori_n163_), .Y(ori_ori_n334_));
  AOI210     o312(.A0(ori_ori_n321_), .A1(ori_ori_n298_), .B0(ori_ori_n334_), .Y(ori_ori_n335_));
  NOi32      o313(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n336_));
  INV        o314(.A(ori_ori_n336_), .Y(ori_ori_n337_));
  NAi21      o315(.An(i_0_), .B(i_6_), .Y(ori_ori_n338_));
  NAi21      o316(.An(i_1_), .B(i_5_), .Y(ori_ori_n339_));
  NA2        o317(.A(ori_ori_n339_), .B(ori_ori_n338_), .Y(ori_ori_n340_));
  NA2        o318(.A(ori_ori_n340_), .B(ori_ori_n25_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n341_), .B(ori_ori_n160_), .Y(ori_ori_n342_));
  NAi41      o320(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(ori_ori_n343_));
  OAI220     o321(.A0(ori_ori_n343_), .A1(ori_ori_n339_), .B0(ori_ori_n216_), .B1(ori_ori_n160_), .Y(ori_ori_n344_));
  AOI210     o322(.A0(ori_ori_n343_), .A1(ori_ori_n160_), .B0(ori_ori_n158_), .Y(ori_ori_n345_));
  NOi32      o323(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n346_));
  NAi21      o324(.An(i_6_), .B(i_1_), .Y(ori_ori_n347_));
  NA3        o325(.A(ori_ori_n347_), .B(ori_ori_n346_), .C(ori_ori_n46_), .Y(ori_ori_n348_));
  NO2        o326(.A(ori_ori_n348_), .B(i_0_), .Y(ori_ori_n349_));
  OR3        o327(.A(ori_ori_n349_), .B(ori_ori_n345_), .C(ori_ori_n344_), .Y(ori_ori_n350_));
  NO2        o328(.A(i_1_), .B(ori_ori_n101_), .Y(ori_ori_n351_));
  NAi21      o329(.An(i_3_), .B(i_4_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(i_9_), .Y(ori_ori_n353_));
  AN2        o331(.A(i_6_), .B(i_7_), .Y(ori_ori_n354_));
  OAI210     o332(.A0(ori_ori_n354_), .A1(ori_ori_n351_), .B0(ori_ori_n353_), .Y(ori_ori_n355_));
  NA2        o333(.A(i_2_), .B(i_7_), .Y(ori_ori_n356_));
  NO2        o334(.A(ori_ori_n352_), .B(i_10_), .Y(ori_ori_n357_));
  NA3        o335(.A(ori_ori_n357_), .B(ori_ori_n356_), .C(ori_ori_n237_), .Y(ori_ori_n358_));
  AOI210     o336(.A0(ori_ori_n358_), .A1(ori_ori_n355_), .B0(ori_ori_n181_), .Y(ori_ori_n359_));
  AOI210     o337(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(ori_ori_n360_));
  OAI210     o338(.A0(ori_ori_n360_), .A1(ori_ori_n184_), .B0(ori_ori_n357_), .Y(ori_ori_n361_));
  AOI220     o339(.A0(ori_ori_n357_), .A1(ori_ori_n320_), .B0(ori_ori_n231_), .B1(ori_ori_n184_), .Y(ori_ori_n362_));
  AOI210     o340(.A0(ori_ori_n362_), .A1(ori_ori_n361_), .B0(i_5_), .Y(ori_ori_n363_));
  NO4        o341(.A(ori_ori_n363_), .B(ori_ori_n359_), .C(ori_ori_n350_), .D(ori_ori_n342_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n364_), .B(ori_ori_n337_), .Y(ori_ori_n365_));
  NO2        o343(.A(ori_ori_n58_), .B(ori_ori_n25_), .Y(ori_ori_n366_));
  AN2        o344(.A(i_12_), .B(i_5_), .Y(ori_ori_n367_));
  NO2        o345(.A(i_4_), .B(ori_ori_n26_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n368_), .B(ori_ori_n367_), .Y(ori_ori_n369_));
  NO2        o347(.A(i_11_), .B(i_6_), .Y(ori_ori_n370_));
  NA3        o348(.A(ori_ori_n370_), .B(ori_ori_n308_), .C(ori_ori_n219_), .Y(ori_ori_n371_));
  NO2        o349(.A(ori_ori_n371_), .B(ori_ori_n369_), .Y(ori_ori_n372_));
  NO2        o350(.A(ori_ori_n235_), .B(i_5_), .Y(ori_ori_n373_));
  NO2        o351(.A(i_5_), .B(i_10_), .Y(ori_ori_n374_));
  AOI220     o352(.A0(ori_ori_n374_), .A1(ori_ori_n260_), .B0(ori_ori_n373_), .B1(ori_ori_n193_), .Y(ori_ori_n375_));
  NA2        o353(.A(ori_ori_n145_), .B(ori_ori_n45_), .Y(ori_ori_n376_));
  NO2        o354(.A(ori_ori_n376_), .B(ori_ori_n375_), .Y(ori_ori_n377_));
  OAI210     o355(.A0(ori_ori_n377_), .A1(ori_ori_n372_), .B0(ori_ori_n366_), .Y(ori_ori_n378_));
  NO2        o356(.A(ori_ori_n37_), .B(ori_ori_n25_), .Y(ori_ori_n379_));
  NO2        o357(.A(ori_ori_n151_), .B(ori_ori_n85_), .Y(ori_ori_n380_));
  OAI210     o358(.A0(ori_ori_n380_), .A1(ori_ori_n372_), .B0(ori_ori_n379_), .Y(ori_ori_n381_));
  NO3        o359(.A(ori_ori_n85_), .B(ori_ori_n48_), .C(i_9_), .Y(ori_ori_n382_));
  NA3        o360(.A(ori_ori_n289_), .B(ori_ori_n74_), .C(ori_ori_n54_), .Y(ori_ori_n383_));
  NO2        o361(.A(i_11_), .B(i_12_), .Y(ori_ori_n384_));
  NA2        o362(.A(ori_ori_n384_), .B(ori_ori_n36_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n383_), .B(ori_ori_n385_), .Y(ori_ori_n386_));
  NA2        o364(.A(ori_ori_n374_), .B(ori_ori_n229_), .Y(ori_ori_n387_));
  NAi21      o365(.An(i_13_), .B(i_0_), .Y(ori_ori_n388_));
  NO2        o366(.A(ori_ori_n388_), .B(ori_ori_n232_), .Y(ori_ori_n389_));
  NA2        o367(.A(ori_ori_n386_), .B(ori_ori_n389_), .Y(ori_ori_n390_));
  NA3        o368(.A(ori_ori_n390_), .B(ori_ori_n381_), .C(ori_ori_n378_), .Y(ori_ori_n391_));
  NA2        o369(.A(ori_ori_n44_), .B(ori_ori_n219_), .Y(ori_ori_n392_));
  NO2        o370(.A(i_0_), .B(i_11_), .Y(ori_ori_n393_));
  AN2        o371(.A(i_1_), .B(i_6_), .Y(ori_ori_n394_));
  NOi21      o372(.An(i_2_), .B(i_12_), .Y(ori_ori_n395_));
  NAi21      o373(.An(i_9_), .B(i_4_), .Y(ori_ori_n396_));
  OR2        o374(.A(i_13_), .B(i_10_), .Y(ori_ori_n397_));
  NO3        o375(.A(ori_ori_n397_), .B(ori_ori_n118_), .C(ori_ori_n396_), .Y(ori_ori_n398_));
  NO2        o376(.A(ori_ori_n172_), .B(ori_ori_n124_), .Y(ori_ori_n399_));
  OR2        o377(.A(ori_ori_n211_), .B(ori_ori_n210_), .Y(ori_ori_n400_));
  NO2        o378(.A(ori_ori_n101_), .B(ori_ori_n25_), .Y(ori_ori_n401_));
  NA2        o379(.A(ori_ori_n275_), .B(ori_ori_n401_), .Y(ori_ori_n402_));
  NA2        o380(.A(ori_ori_n268_), .B(ori_ori_n206_), .Y(ori_ori_n403_));
  OAI220     o381(.A0(ori_ori_n403_), .A1(ori_ori_n400_), .B0(ori_ori_n402_), .B1(ori_ori_n327_), .Y(ori_ori_n404_));
  INV        o382(.A(ori_ori_n404_), .Y(ori_ori_n405_));
  NO2        o383(.A(ori_ori_n405_), .B(ori_ori_n26_), .Y(ori_ori_n406_));
  NA2        o384(.A(ori_ori_n306_), .B(ori_ori_n305_), .Y(ori_ori_n407_));
  NO2        o385(.A(ori_ori_n178_), .B(ori_ori_n85_), .Y(ori_ori_n408_));
  AOI220     o386(.A0(ori_ori_n408_), .A1(i_1_), .B0(ori_ori_n270_), .B1(ori_ori_n206_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n409_), .B(ori_ori_n277_), .Y(ori_ori_n410_));
  NO2        o388(.A(ori_ori_n410_), .B(ori_ori_n407_), .Y(ori_ori_n411_));
  NA2        o389(.A(ori_ori_n191_), .B(ori_ori_n96_), .Y(ori_ori_n412_));
  NA2        o390(.A(ori_ori_n308_), .B(ori_ori_n164_), .Y(ori_ori_n413_));
  AOI210     o391(.A0(ori_ori_n413_), .A1(ori_ori_n412_), .B0(ori_ori_n307_), .Y(ori_ori_n414_));
  NA2        o392(.A(ori_ori_n188_), .B(i_10_), .Y(ori_ori_n415_));
  NA3        o393(.A(ori_ori_n246_), .B(ori_ori_n63_), .C(i_2_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n286_), .B(ori_ori_n227_), .Y(ori_ori_n417_));
  OAI220     o395(.A0(ori_ori_n417_), .A1(ori_ori_n178_), .B0(ori_ori_n416_), .B1(ori_ori_n415_), .Y(ori_ori_n418_));
  NO2        o396(.A(i_3_), .B(ori_ori_n48_), .Y(ori_ori_n419_));
  NO2        o397(.A(ori_ori_n418_), .B(ori_ori_n414_), .Y(ori_ori_n420_));
  AOI210     o398(.A0(ori_ori_n420_), .A1(ori_ori_n411_), .B0(ori_ori_n262_), .Y(ori_ori_n421_));
  NO4        o399(.A(ori_ori_n421_), .B(ori_ori_n406_), .C(ori_ori_n391_), .D(ori_ori_n365_), .Y(ori_ori_n422_));
  NO2        o400(.A(ori_ori_n72_), .B(i_13_), .Y(ori_ori_n423_));
  NO2        o401(.A(i_10_), .B(i_9_), .Y(ori_ori_n424_));
  NAi21      o402(.An(i_12_), .B(i_8_), .Y(ori_ori_n425_));
  NO2        o403(.A(ori_ori_n425_), .B(i_3_), .Y(ori_ori_n426_));
  NO2        o404(.A(ori_ori_n46_), .B(i_4_), .Y(ori_ori_n427_));
  NA2        o405(.A(ori_ori_n427_), .B(ori_ori_n104_), .Y(ori_ori_n428_));
  NO2        o406(.A(ori_ori_n428_), .B(ori_ori_n200_), .Y(ori_ori_n429_));
  NO3        o407(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n430_));
  NA2        o408(.A(ori_ori_n257_), .B(ori_ori_n97_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n431_), .B(ori_ori_n430_), .Y(ori_ori_n432_));
  NA2        o410(.A(i_8_), .B(i_9_), .Y(ori_ori_n433_));
  AOI210     o411(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n434_));
  OR2        o412(.A(ori_ori_n434_), .B(ori_ori_n433_), .Y(ori_ori_n435_));
  NA2        o413(.A(ori_ori_n275_), .B(ori_ori_n201_), .Y(ori_ori_n436_));
  NO2        o414(.A(ori_ori_n436_), .B(ori_ori_n435_), .Y(ori_ori_n437_));
  NA2        o415(.A(ori_ori_n241_), .B(ori_ori_n294_), .Y(ori_ori_n438_));
  NO3        o416(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n439_));
  INV        o417(.A(ori_ori_n439_), .Y(ori_ori_n440_));
  NA3        o418(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n441_));
  NA4        o419(.A(ori_ori_n146_), .B(ori_ori_n116_), .C(ori_ori_n79_), .D(ori_ori_n23_), .Y(ori_ori_n442_));
  OAI220     o420(.A0(ori_ori_n442_), .A1(ori_ori_n441_), .B0(ori_ori_n440_), .B1(ori_ori_n438_), .Y(ori_ori_n443_));
  NO3        o421(.A(ori_ori_n443_), .B(ori_ori_n437_), .C(ori_ori_n429_), .Y(ori_ori_n444_));
  NA2        o422(.A(ori_ori_n96_), .B(i_13_), .Y(ori_ori_n445_));
  NA2        o423(.A(ori_ori_n408_), .B(ori_ori_n366_), .Y(ori_ori_n446_));
  NO2        o424(.A(i_2_), .B(i_13_), .Y(ori_ori_n447_));
  NO2        o425(.A(ori_ori_n446_), .B(ori_ori_n445_), .Y(ori_ori_n448_));
  NO3        o426(.A(i_4_), .B(ori_ori_n48_), .C(i_8_), .Y(ori_ori_n449_));
  NO2        o427(.A(i_6_), .B(i_7_), .Y(ori_ori_n450_));
  NO2        o428(.A(i_11_), .B(i_1_), .Y(ori_ori_n451_));
  OR2        o429(.A(i_11_), .B(i_8_), .Y(ori_ori_n452_));
  NOi21      o430(.An(i_2_), .B(i_7_), .Y(ori_ori_n453_));
  NO2        o431(.A(i_3_), .B(ori_ori_n188_), .Y(ori_ori_n454_));
  NO2        o432(.A(i_6_), .B(i_10_), .Y(ori_ori_n455_));
  NA4        o433(.A(ori_ori_n455_), .B(ori_ori_n298_), .C(ori_ori_n454_), .D(ori_ori_n229_), .Y(ori_ori_n456_));
  NO2        o434(.A(ori_ori_n456_), .B(ori_ori_n156_), .Y(ori_ori_n457_));
  NA3        o435(.A(ori_ori_n238_), .B(ori_ori_n171_), .C(ori_ori_n133_), .Y(ori_ori_n458_));
  NA2        o436(.A(ori_ori_n46_), .B(ori_ori_n44_), .Y(ori_ori_n459_));
  NO2        o437(.A(ori_ori_n158_), .B(i_3_), .Y(ori_ori_n460_));
  NAi31      o438(.An(ori_ori_n459_), .B(ori_ori_n460_), .C(ori_ori_n220_), .Y(ori_ori_n461_));
  NA3        o439(.A(ori_ori_n379_), .B(ori_ori_n175_), .C(ori_ori_n150_), .Y(ori_ori_n462_));
  NA3        o440(.A(ori_ori_n462_), .B(ori_ori_n461_), .C(ori_ori_n458_), .Y(ori_ori_n463_));
  NO3        o441(.A(ori_ori_n463_), .B(ori_ori_n457_), .C(ori_ori_n448_), .Y(ori_ori_n464_));
  NA2        o442(.A(ori_ori_n430_), .B(ori_ori_n367_), .Y(ori_ori_n465_));
  NA2        o443(.A(ori_ori_n439_), .B(ori_ori_n374_), .Y(ori_ori_n466_));
  NAi21      o444(.An(ori_ori_n211_), .B(ori_ori_n384_), .Y(ori_ori_n467_));
  NO2        o445(.A(ori_ori_n26_), .B(i_5_), .Y(ori_ori_n468_));
  NO2        o446(.A(i_0_), .B(ori_ori_n85_), .Y(ori_ori_n469_));
  NA3        o447(.A(ori_ori_n469_), .B(ori_ori_n468_), .C(ori_ori_n143_), .Y(ori_ori_n470_));
  OR3        o448(.A(ori_ori_n292_), .B(ori_ori_n38_), .C(ori_ori_n46_), .Y(ori_ori_n471_));
  NO2        o449(.A(ori_ori_n471_), .B(ori_ori_n470_), .Y(ori_ori_n472_));
  NA2        o450(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n473_));
  NA2        o451(.A(ori_ori_n298_), .B(ori_ori_n231_), .Y(ori_ori_n474_));
  OAI220     o452(.A0(ori_ori_n474_), .A1(ori_ori_n416_), .B0(ori_ori_n473_), .B1(ori_ori_n445_), .Y(ori_ori_n475_));
  NO2        o453(.A(ori_ori_n475_), .B(ori_ori_n472_), .Y(ori_ori_n476_));
  NA3        o454(.A(ori_ori_n476_), .B(ori_ori_n464_), .C(ori_ori_n444_), .Y(ori_ori_n477_));
  NA2        o455(.A(ori_ori_n123_), .B(ori_ori_n112_), .Y(ori_ori_n478_));
  AN2        o456(.A(ori_ori_n478_), .B(ori_ori_n430_), .Y(ori_ori_n479_));
  NA2        o457(.A(ori_ori_n479_), .B(ori_ori_n295_), .Y(ori_ori_n480_));
  NA2        o458(.A(ori_ori_n367_), .B(ori_ori_n219_), .Y(ori_ori_n481_));
  NA2        o459(.A(ori_ori_n336_), .B(ori_ori_n72_), .Y(ori_ori_n482_));
  NA2        o460(.A(ori_ori_n354_), .B(ori_ori_n346_), .Y(ori_ori_n483_));
  OR2        o461(.A(ori_ori_n481_), .B(ori_ori_n483_), .Y(ori_ori_n484_));
  NO2        o462(.A(ori_ori_n36_), .B(i_8_), .Y(ori_ori_n485_));
  AOI210     o463(.A0(ori_ori_n39_), .A1(i_13_), .B0(ori_ori_n398_), .Y(ori_ori_n486_));
  NA2        o464(.A(ori_ori_n486_), .B(ori_ori_n484_), .Y(ori_ori_n487_));
  INV        o465(.A(ori_ori_n487_), .Y(ori_ori_n488_));
  NA2        o466(.A(ori_ori_n246_), .B(ori_ori_n63_), .Y(ori_ori_n489_));
  OAI210     o467(.A0(i_8_), .A1(ori_ori_n489_), .B0(ori_ori_n135_), .Y(ori_ori_n490_));
  AOI210     o468(.A0(ori_ori_n189_), .A1(i_9_), .B0(ori_ori_n256_), .Y(ori_ori_n491_));
  NO2        o469(.A(ori_ori_n491_), .B(ori_ori_n194_), .Y(ori_ori_n492_));
  NO2        o470(.A(ori_ori_n178_), .B(ori_ori_n85_), .Y(ori_ori_n493_));
  AOI220     o471(.A0(ori_ori_n493_), .A1(ori_ori_n492_), .B0(ori_ori_n490_), .B1(ori_ori_n399_), .Y(ori_ori_n494_));
  NA3        o472(.A(ori_ori_n494_), .B(ori_ori_n488_), .C(ori_ori_n480_), .Y(ori_ori_n495_));
  NO2        o473(.A(i_12_), .B(ori_ori_n188_), .Y(ori_ori_n496_));
  NA2        o474(.A(ori_ori_n496_), .B(ori_ori_n219_), .Y(ori_ori_n497_));
  NO2        o475(.A(i_8_), .B(i_7_), .Y(ori_ori_n498_));
  OAI210     o476(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(ori_ori_n499_));
  NA2        o477(.A(ori_ori_n499_), .B(ori_ori_n218_), .Y(ori_ori_n500_));
  AOI220     o478(.A0(ori_ori_n308_), .A1(ori_ori_n40_), .B0(ori_ori_n227_), .B1(ori_ori_n203_), .Y(ori_ori_n501_));
  OAI220     o479(.A0(ori_ori_n501_), .A1(ori_ori_n178_), .B0(ori_ori_n500_), .B1(ori_ori_n235_), .Y(ori_ori_n502_));
  NA2        o480(.A(ori_ori_n44_), .B(i_10_), .Y(ori_ori_n503_));
  NO2        o481(.A(ori_ori_n503_), .B(i_6_), .Y(ori_ori_n504_));
  NA3        o482(.A(ori_ori_n504_), .B(ori_ori_n502_), .C(ori_ori_n498_), .Y(ori_ori_n505_));
  AOI220     o483(.A0(ori_ori_n408_), .A1(ori_ori_n308_), .B0(ori_ori_n239_), .B1(ori_ori_n237_), .Y(ori_ori_n506_));
  OAI220     o484(.A0(ori_ori_n506_), .A1(ori_ori_n253_), .B0(ori_ori_n445_), .B1(ori_ori_n134_), .Y(ori_ori_n507_));
  NA2        o485(.A(ori_ori_n507_), .B(ori_ori_n256_), .Y(ori_ori_n508_));
  NOi31      o486(.An(ori_ori_n282_), .B(ori_ori_n290_), .C(i_4_), .Y(ori_ori_n509_));
  NA3        o487(.A(ori_ori_n293_), .B(ori_ori_n173_), .C(ori_ori_n96_), .Y(ori_ori_n510_));
  NO2        o488(.A(ori_ori_n217_), .B(ori_ori_n44_), .Y(ori_ori_n511_));
  NO2        o489(.A(ori_ori_n158_), .B(i_5_), .Y(ori_ori_n512_));
  NA3        o490(.A(ori_ori_n512_), .B(ori_ori_n392_), .C(ori_ori_n302_), .Y(ori_ori_n513_));
  OAI210     o491(.A0(ori_ori_n513_), .A1(ori_ori_n511_), .B0(ori_ori_n510_), .Y(ori_ori_n514_));
  OAI210     o492(.A0(ori_ori_n514_), .A1(ori_ori_n509_), .B0(ori_ori_n439_), .Y(ori_ori_n515_));
  NA3        o493(.A(ori_ori_n515_), .B(ori_ori_n508_), .C(ori_ori_n505_), .Y(ori_ori_n516_));
  NA2        o494(.A(ori_ori_n286_), .B(ori_ori_n278_), .Y(ori_ori_n517_));
  NO2        o495(.A(ori_ori_n517_), .B(ori_ori_n172_), .Y(ori_ori_n518_));
  AOI210     o496(.A0(ori_ori_n347_), .A1(ori_ori_n46_), .B0(ori_ori_n351_), .Y(ori_ori_n519_));
  NA2        o497(.A(i_0_), .B(ori_ori_n48_), .Y(ori_ori_n520_));
  NA3        o498(.A(ori_ori_n496_), .B(ori_ori_n266_), .C(ori_ori_n520_), .Y(ori_ori_n521_));
  NO2        o499(.A(ori_ori_n519_), .B(ori_ori_n521_), .Y(ori_ori_n522_));
  NO2        o500(.A(ori_ori_n522_), .B(ori_ori_n518_), .Y(ori_ori_n523_));
  NO3        o501(.A(i_1_), .B(i_5_), .C(i_10_), .Y(ori_ori_n524_));
  NO2        o502(.A(ori_ori_n225_), .B(ori_ori_n36_), .Y(ori_ori_n525_));
  NO2        o503(.A(ori_ori_n397_), .B(i_1_), .Y(ori_ori_n526_));
  NOi31      o504(.An(ori_ori_n526_), .B(ori_ori_n431_), .C(ori_ori_n72_), .Y(ori_ori_n527_));
  NOi21      o505(.An(i_10_), .B(i_6_), .Y(ori_ori_n528_));
  NO2        o506(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n529_));
  NO2        o507(.A(ori_ori_n115_), .B(ori_ori_n23_), .Y(ori_ori_n530_));
  NA2        o508(.A(ori_ori_n299_), .B(ori_ori_n165_), .Y(ori_ori_n531_));
  AOI220     o509(.A0(ori_ori_n531_), .A1(ori_ori_n417_), .B0(ori_ori_n179_), .B1(ori_ori_n177_), .Y(ori_ori_n532_));
  NO2        o510(.A(ori_ori_n193_), .B(ori_ori_n37_), .Y(ori_ori_n533_));
  NOi31      o511(.An(ori_ori_n147_), .B(ori_ori_n533_), .C(ori_ori_n315_), .Y(ori_ori_n534_));
  NO2        o512(.A(ori_ori_n534_), .B(ori_ori_n532_), .Y(ori_ori_n535_));
  NO2        o513(.A(ori_ori_n482_), .B(ori_ori_n362_), .Y(ori_ori_n536_));
  INV        o514(.A(ori_ori_n302_), .Y(ori_ori_n537_));
  NO2        o515(.A(i_12_), .B(ori_ori_n85_), .Y(ori_ori_n538_));
  NA3        o516(.A(ori_ori_n538_), .B(ori_ori_n266_), .C(ori_ori_n520_), .Y(ori_ori_n539_));
  NA3        o517(.A(ori_ori_n370_), .B(ori_ori_n275_), .C(ori_ori_n213_), .Y(ori_ori_n540_));
  AOI210     o518(.A0(ori_ori_n540_), .A1(ori_ori_n539_), .B0(ori_ori_n537_), .Y(ori_ori_n541_));
  NO3        o519(.A(i_4_), .B(ori_ori_n324_), .C(ori_ori_n290_), .Y(ori_ori_n542_));
  OR2        o520(.A(i_2_), .B(i_5_), .Y(ori_ori_n543_));
  OR2        o521(.A(ori_ori_n543_), .B(ori_ori_n394_), .Y(ori_ori_n544_));
  AOI210     o522(.A0(ori_ori_n356_), .A1(ori_ori_n237_), .B0(ori_ori_n193_), .Y(ori_ori_n545_));
  AOI210     o523(.A0(ori_ori_n545_), .A1(ori_ori_n544_), .B0(ori_ori_n467_), .Y(ori_ori_n546_));
  NO4        o524(.A(ori_ori_n546_), .B(ori_ori_n542_), .C(ori_ori_n541_), .D(ori_ori_n536_), .Y(ori_ori_n547_));
  NA3        o525(.A(ori_ori_n547_), .B(ori_ori_n535_), .C(ori_ori_n523_), .Y(ori_ori_n548_));
  NO4        o526(.A(ori_ori_n548_), .B(ori_ori_n516_), .C(ori_ori_n495_), .D(ori_ori_n477_), .Y(ori_ori_n549_));
  NA4        o527(.A(ori_ori_n549_), .B(ori_ori_n422_), .C(ori_ori_n335_), .D(ori_ori_n297_), .Y(ori7));
  NO2        o528(.A(ori_ori_n92_), .B(ori_ori_n54_), .Y(ori_ori_n551_));
  NO2        o529(.A(ori_ori_n108_), .B(ori_ori_n89_), .Y(ori_ori_n552_));
  NA2        o530(.A(ori_ori_n368_), .B(ori_ori_n552_), .Y(ori_ori_n553_));
  NA2        o531(.A(ori_ori_n455_), .B(ori_ori_n83_), .Y(ori_ori_n554_));
  NA2        o532(.A(i_11_), .B(ori_ori_n188_), .Y(ori_ori_n555_));
  NA2        o533(.A(ori_ori_n145_), .B(ori_ori_n555_), .Y(ori_ori_n556_));
  OAI210     o534(.A0(ori_ori_n556_), .A1(ori_ori_n554_), .B0(ori_ori_n553_), .Y(ori_ori_n557_));
  NA3        o535(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n558_));
  NO2        o536(.A(ori_ori_n229_), .B(i_4_), .Y(ori_ori_n559_));
  NA2        o537(.A(ori_ori_n559_), .B(i_8_), .Y(ori_ori_n560_));
  NO2        o538(.A(ori_ori_n105_), .B(ori_ori_n558_), .Y(ori_ori_n561_));
  NA2        o539(.A(i_2_), .B(ori_ori_n85_), .Y(ori_ori_n562_));
  OAI210     o540(.A0(ori_ori_n86_), .A1(ori_ori_n198_), .B0(ori_ori_n199_), .Y(ori_ori_n563_));
  NO2        o541(.A(i_7_), .B(ori_ori_n37_), .Y(ori_ori_n564_));
  NA2        o542(.A(i_4_), .B(i_8_), .Y(ori_ori_n565_));
  AOI210     o543(.A0(ori_ori_n565_), .A1(ori_ori_n293_), .B0(ori_ori_n564_), .Y(ori_ori_n566_));
  OAI220     o544(.A0(ori_ori_n566_), .A1(ori_ori_n562_), .B0(ori_ori_n563_), .B1(i_13_), .Y(ori_ori_n567_));
  NO4        o545(.A(ori_ori_n567_), .B(ori_ori_n561_), .C(ori_ori_n557_), .D(ori_ori_n551_), .Y(ori_ori_n568_));
  AOI210     o546(.A0(ori_ori_n129_), .A1(ori_ori_n61_), .B0(i_10_), .Y(ori_ori_n569_));
  AOI210     o547(.A0(ori_ori_n569_), .A1(ori_ori_n229_), .B0(ori_ori_n162_), .Y(ori_ori_n570_));
  OR2        o548(.A(i_6_), .B(i_10_), .Y(ori_ori_n571_));
  OR3        o549(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n572_));
  INV        o550(.A(ori_ori_n195_), .Y(ori_ori_n573_));
  OR2        o551(.A(ori_ori_n570_), .B(ori_ori_n258_), .Y(ori_ori_n574_));
  AOI210     o552(.A0(ori_ori_n574_), .A1(ori_ori_n568_), .B0(ori_ori_n62_), .Y(ori_ori_n575_));
  NOi21      o553(.An(i_11_), .B(i_7_), .Y(ori_ori_n576_));
  AO210      o554(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n577_));
  NO2        o555(.A(ori_ori_n577_), .B(ori_ori_n576_), .Y(ori_ori_n578_));
  NA2        o556(.A(ori_ori_n578_), .B(ori_ori_n203_), .Y(ori_ori_n579_));
  NO2        o557(.A(ori_ori_n579_), .B(ori_ori_n62_), .Y(ori_ori_n580_));
  OR2        o558(.A(ori_ori_n362_), .B(ori_ori_n41_), .Y(ori_ori_n581_));
  NO3        o559(.A(ori_ori_n248_), .B(ori_ori_n204_), .C(ori_ori_n555_), .Y(ori_ori_n582_));
  OAI210     o560(.A0(ori_ori_n582_), .A1(ori_ori_n220_), .B0(ori_ori_n62_), .Y(ori_ori_n583_));
  NA2        o561(.A(ori_ori_n395_), .B(ori_ori_n31_), .Y(ori_ori_n584_));
  OR2        o562(.A(ori_ori_n204_), .B(ori_ori_n108_), .Y(ori_ori_n585_));
  NA2        o563(.A(ori_ori_n585_), .B(ori_ori_n584_), .Y(ori_ori_n586_));
  NO2        o564(.A(ori_ori_n62_), .B(i_9_), .Y(ori_ori_n587_));
  NO2        o565(.A(ori_ori_n587_), .B(i_4_), .Y(ori_ori_n588_));
  NA2        o566(.A(ori_ori_n588_), .B(ori_ori_n586_), .Y(ori_ori_n589_));
  NO2        o567(.A(i_1_), .B(i_12_), .Y(ori_ori_n590_));
  NA3        o568(.A(ori_ori_n590_), .B(ori_ori_n110_), .C(ori_ori_n24_), .Y(ori_ori_n591_));
  BUFFER     o569(.A(ori_ori_n591_), .Y(ori_ori_n592_));
  NA4        o570(.A(ori_ori_n592_), .B(ori_ori_n589_), .C(ori_ori_n583_), .D(ori_ori_n581_), .Y(ori_ori_n593_));
  OAI210     o571(.A0(ori_ori_n593_), .A1(ori_ori_n580_), .B0(i_6_), .Y(ori_ori_n594_));
  NO2        o572(.A(ori_ori_n229_), .B(ori_ori_n85_), .Y(ori_ori_n595_));
  NO2        o573(.A(ori_ori_n595_), .B(i_11_), .Y(ori_ori_n596_));
  INV        o574(.A(ori_ori_n432_), .Y(ori_ori_n597_));
  NA2        o575(.A(ori_ori_n229_), .B(i_6_), .Y(ori_ori_n598_));
  NO3        o576(.A(ori_ori_n571_), .B(ori_ori_n225_), .C(ori_ori_n23_), .Y(ori_ori_n599_));
  AOI210     o577(.A0(i_1_), .A1(ori_ori_n249_), .B0(ori_ori_n599_), .Y(ori_ori_n600_));
  NO2        o578(.A(ori_ori_n600_), .B(ori_ori_n44_), .Y(ori_ori_n601_));
  NA3        o579(.A(ori_ori_n498_), .B(i_11_), .C(ori_ori_n36_), .Y(ori_ori_n602_));
  INV        o580(.A(i_2_), .Y(ori_ori_n603_));
  NA2        o581(.A(ori_ori_n139_), .B(i_9_), .Y(ori_ori_n604_));
  NO2        o582(.A(ori_ori_n46_), .B(i_1_), .Y(ori_ori_n605_));
  NO2        o583(.A(ori_ori_n604_), .B(ori_ori_n603_), .Y(ori_ori_n606_));
  NA3        o584(.A(ori_ori_n587_), .B(ori_ori_n302_), .C(i_6_), .Y(ori_ori_n607_));
  NO2        o585(.A(ori_ori_n607_), .B(ori_ori_n23_), .Y(ori_ori_n608_));
  AOI210     o586(.A0(ori_ori_n451_), .A1(ori_ori_n401_), .B0(ori_ori_n234_), .Y(ori_ori_n609_));
  NO2        o587(.A(ori_ori_n609_), .B(ori_ori_n562_), .Y(ori_ori_n610_));
  NAi21      o588(.An(ori_ori_n602_), .B(ori_ori_n91_), .Y(ori_ori_n611_));
  NA2        o589(.A(ori_ori_n605_), .B(ori_ori_n257_), .Y(ori_ori_n612_));
  NO2        o590(.A(i_11_), .B(ori_ori_n37_), .Y(ori_ori_n613_));
  NA2        o591(.A(ori_ori_n613_), .B(ori_ori_n24_), .Y(ori_ori_n614_));
  OAI210     o592(.A0(ori_ori_n614_), .A1(ori_ori_n612_), .B0(ori_ori_n611_), .Y(ori_ori_n615_));
  OR4        o593(.A(ori_ori_n615_), .B(ori_ori_n610_), .C(ori_ori_n608_), .D(ori_ori_n606_), .Y(ori_ori_n616_));
  NO3        o594(.A(ori_ori_n616_), .B(ori_ori_n601_), .C(ori_ori_n597_), .Y(ori_ori_n617_));
  NO2        o595(.A(ori_ori_n229_), .B(ori_ori_n101_), .Y(ori_ori_n618_));
  NO2        o596(.A(ori_ori_n618_), .B(ori_ori_n576_), .Y(ori_ori_n619_));
  NA2        o597(.A(ori_ori_n619_), .B(i_1_), .Y(ori_ori_n620_));
  NO2        o598(.A(ori_ori_n620_), .B(ori_ori_n572_), .Y(ori_ori_n621_));
  NO2        o599(.A(ori_ori_n396_), .B(ori_ori_n85_), .Y(ori_ori_n622_));
  NA2        o600(.A(ori_ori_n621_), .B(ori_ori_n46_), .Y(ori_ori_n623_));
  NA2        o601(.A(i_3_), .B(ori_ori_n188_), .Y(ori_ori_n624_));
  NO2        o602(.A(ori_ori_n225_), .B(ori_ori_n44_), .Y(ori_ori_n625_));
  NO3        o603(.A(ori_ori_n625_), .B(ori_ori_n295_), .C(ori_ori_n230_), .Y(ori_ori_n626_));
  NO2        o604(.A(ori_ori_n118_), .B(ori_ori_n37_), .Y(ori_ori_n627_));
  NO2        o605(.A(ori_ori_n627_), .B(i_6_), .Y(ori_ori_n628_));
  NO2        o606(.A(ori_ori_n85_), .B(i_9_), .Y(ori_ori_n629_));
  NO2        o607(.A(ori_ori_n629_), .B(ori_ori_n62_), .Y(ori_ori_n630_));
  NO2        o608(.A(ori_ori_n630_), .B(ori_ori_n590_), .Y(ori_ori_n631_));
  NO4        o609(.A(ori_ori_n631_), .B(ori_ori_n628_), .C(ori_ori_n626_), .D(i_4_), .Y(ori_ori_n632_));
  NA2        o610(.A(i_1_), .B(i_3_), .Y(ori_ori_n633_));
  NO2        o611(.A(ori_ori_n433_), .B(ori_ori_n92_), .Y(ori_ori_n634_));
  AOI210     o612(.A0(ori_ori_n625_), .A1(ori_ori_n528_), .B0(ori_ori_n634_), .Y(ori_ori_n635_));
  NO2        o613(.A(ori_ori_n635_), .B(ori_ori_n633_), .Y(ori_ori_n636_));
  NO2        o614(.A(ori_ori_n636_), .B(ori_ori_n632_), .Y(ori_ori_n637_));
  NA4        o615(.A(ori_ori_n637_), .B(ori_ori_n623_), .C(ori_ori_n617_), .D(ori_ori_n594_), .Y(ori_ori_n638_));
  NO3        o616(.A(ori_ori_n452_), .B(i_3_), .C(i_7_), .Y(ori_ori_n639_));
  NA2        o617(.A(ori_ori_n354_), .B(ori_ori_n353_), .Y(ori_ori_n640_));
  NA3        o618(.A(ori_ori_n455_), .B(ori_ori_n485_), .C(ori_ori_n46_), .Y(ori_ori_n641_));
  NA3        o619(.A(ori_ori_n162_), .B(ori_ori_n83_), .C(ori_ori_n85_), .Y(ori_ori_n642_));
  NA3        o620(.A(ori_ori_n642_), .B(ori_ori_n641_), .C(ori_ori_n640_), .Y(ori_ori_n643_));
  NA2        o621(.A(ori_ori_n643_), .B(i_1_), .Y(ori_ori_n644_));
  AOI210     o622(.A0(ori_ori_n257_), .A1(ori_ori_n97_), .B0(i_1_), .Y(ori_ori_n645_));
  NO2        o623(.A(ori_ori_n352_), .B(i_2_), .Y(ori_ori_n646_));
  NA2        o624(.A(ori_ori_n646_), .B(ori_ori_n645_), .Y(ori_ori_n647_));
  OAI210     o625(.A0(ori_ori_n607_), .A1(ori_ori_n425_), .B0(ori_ori_n647_), .Y(ori_ori_n648_));
  INV        o626(.A(ori_ori_n648_), .Y(ori_ori_n649_));
  AOI210     o627(.A0(ori_ori_n649_), .A1(ori_ori_n644_), .B0(i_13_), .Y(ori_ori_n650_));
  OR2        o628(.A(i_11_), .B(i_7_), .Y(ori_ori_n651_));
  NA3        o629(.A(ori_ori_n651_), .B(ori_ori_n106_), .C(ori_ori_n139_), .Y(ori_ori_n652_));
  AOI220     o630(.A0(ori_ori_n447_), .A1(ori_ori_n162_), .B0(ori_ori_n427_), .B1(ori_ori_n139_), .Y(ori_ori_n653_));
  OAI210     o631(.A0(ori_ori_n653_), .A1(ori_ori_n44_), .B0(ori_ori_n652_), .Y(ori_ori_n654_));
  NO2        o632(.A(ori_ori_n54_), .B(i_12_), .Y(ori_ori_n655_));
  NO2        o633(.A(ori_ori_n453_), .B(ori_ori_n24_), .Y(ori_ori_n656_));
  AOI220     o634(.A0(ori_ori_n656_), .A1(ori_ori_n622_), .B0(ori_ori_n238_), .B1(ori_ori_n132_), .Y(ori_ori_n657_));
  OAI220     o635(.A0(ori_ori_n657_), .A1(ori_ori_n41_), .B0(ori_ori_n961_), .B1(ori_ori_n92_), .Y(ori_ori_n658_));
  AOI210     o636(.A0(ori_ori_n654_), .A1(ori_ori_n317_), .B0(ori_ori_n658_), .Y(ori_ori_n659_));
  INV        o637(.A(ori_ori_n115_), .Y(ori_ori_n660_));
  AOI220     o638(.A0(ori_ori_n660_), .A1(ori_ori_n71_), .B0(ori_ori_n370_), .B1(ori_ori_n605_), .Y(ori_ori_n661_));
  NO2        o639(.A(ori_ori_n661_), .B(ori_ori_n235_), .Y(ori_ori_n662_));
  AOI210     o640(.A0(ori_ori_n425_), .A1(ori_ori_n36_), .B0(i_13_), .Y(ori_ori_n663_));
  NOi31      o641(.An(ori_ori_n663_), .B(ori_ori_n554_), .C(ori_ori_n44_), .Y(ori_ori_n664_));
  NA2        o642(.A(ori_ori_n128_), .B(i_13_), .Y(ori_ori_n665_));
  NO2        o643(.A(ori_ori_n665_), .B(ori_ori_n645_), .Y(ori_ori_n666_));
  NO3        o644(.A(ori_ori_n70_), .B(ori_ori_n32_), .C(ori_ori_n101_), .Y(ori_ori_n667_));
  NA2        o645(.A(ori_ori_n26_), .B(ori_ori_n188_), .Y(ori_ori_n668_));
  NA2        o646(.A(ori_ori_n668_), .B(i_7_), .Y(ori_ori_n669_));
  NO3        o647(.A(ori_ori_n453_), .B(ori_ori_n229_), .C(ori_ori_n85_), .Y(ori_ori_n670_));
  AOI210     o648(.A0(ori_ori_n670_), .A1(ori_ori_n669_), .B0(ori_ori_n667_), .Y(ori_ori_n671_));
  AOI220     o649(.A0(ori_ori_n370_), .A1(ori_ori_n605_), .B0(ori_ori_n91_), .B1(ori_ori_n102_), .Y(ori_ori_n672_));
  OAI220     o650(.A0(ori_ori_n672_), .A1(ori_ori_n560_), .B0(ori_ori_n671_), .B1(ori_ori_n573_), .Y(ori_ori_n673_));
  NO4        o651(.A(ori_ori_n673_), .B(ori_ori_n666_), .C(ori_ori_n664_), .D(ori_ori_n662_), .Y(ori_ori_n674_));
  OR2        o652(.A(i_11_), .B(i_6_), .Y(ori_ori_n675_));
  NA3        o653(.A(ori_ori_n559_), .B(ori_ori_n668_), .C(i_7_), .Y(ori_ori_n676_));
  NO2        o654(.A(ori_ori_n676_), .B(ori_ori_n675_), .Y(ori_ori_n677_));
  NA3        o655(.A(ori_ori_n395_), .B(ori_ori_n564_), .C(ori_ori_n97_), .Y(ori_ori_n678_));
  NA2        o656(.A(ori_ori_n596_), .B(i_13_), .Y(ori_ori_n679_));
  NAi21      o657(.An(i_11_), .B(i_12_), .Y(ori_ori_n680_));
  NOi41      o658(.An(ori_ori_n111_), .B(ori_ori_n680_), .C(i_13_), .D(ori_ori_n85_), .Y(ori_ori_n681_));
  NO3        o659(.A(ori_ori_n453_), .B(ori_ori_n538_), .C(ori_ori_n565_), .Y(ori_ori_n682_));
  AOI220     o660(.A0(ori_ori_n682_), .A1(ori_ori_n298_), .B0(ori_ori_n681_), .B1(ori_ori_n46_), .Y(ori_ori_n683_));
  NA3        o661(.A(ori_ori_n683_), .B(ori_ori_n679_), .C(ori_ori_n678_), .Y(ori_ori_n684_));
  OAI210     o662(.A0(ori_ori_n684_), .A1(ori_ori_n677_), .B0(ori_ori_n62_), .Y(ori_ori_n685_));
  NO2        o663(.A(i_2_), .B(i_12_), .Y(ori_ori_n686_));
  NA2        o664(.A(ori_ori_n351_), .B(ori_ori_n686_), .Y(ori_ori_n687_));
  NO2        o665(.A(ori_ori_n129_), .B(i_2_), .Y(ori_ori_n688_));
  NA2        o666(.A(ori_ori_n688_), .B(ori_ori_n590_), .Y(ori_ori_n689_));
  NA2        o667(.A(ori_ori_n689_), .B(ori_ori_n687_), .Y(ori_ori_n690_));
  NA3        o668(.A(ori_ori_n690_), .B(ori_ori_n45_), .C(ori_ori_n219_), .Y(ori_ori_n691_));
  NA4        o669(.A(ori_ori_n691_), .B(ori_ori_n685_), .C(ori_ori_n674_), .D(ori_ori_n659_), .Y(ori_ori_n692_));
  OR4        o670(.A(ori_ori_n692_), .B(ori_ori_n650_), .C(ori_ori_n638_), .D(ori_ori_n575_), .Y(ori5));
  NA2        o671(.A(ori_ori_n619_), .B(ori_ori_n260_), .Y(ori_ori_n694_));
  AN2        o672(.A(ori_ori_n24_), .B(i_10_), .Y(ori_ori_n695_));
  NA3        o673(.A(ori_ori_n695_), .B(ori_ori_n686_), .C(ori_ori_n108_), .Y(ori_ori_n696_));
  NO2        o674(.A(ori_ori_n560_), .B(i_11_), .Y(ori_ori_n697_));
  NA2        o675(.A(ori_ori_n86_), .B(ori_ori_n697_), .Y(ori_ori_n698_));
  NA3        o676(.A(ori_ori_n698_), .B(ori_ori_n696_), .C(ori_ori_n694_), .Y(ori_ori_n699_));
  NO3        o677(.A(i_11_), .B(ori_ori_n229_), .C(i_13_), .Y(ori_ori_n700_));
  NO2        o678(.A(ori_ori_n125_), .B(ori_ori_n23_), .Y(ori_ori_n701_));
  NA2        o679(.A(i_12_), .B(i_8_), .Y(ori_ori_n702_));
  OAI210     o680(.A0(ori_ori_n46_), .A1(i_3_), .B0(ori_ori_n702_), .Y(ori_ori_n703_));
  INV        o681(.A(ori_ori_n424_), .Y(ori_ori_n704_));
  AOI220     o682(.A0(ori_ori_n302_), .A1(ori_ori_n530_), .B0(ori_ori_n703_), .B1(ori_ori_n701_), .Y(ori_ori_n705_));
  INV        o683(.A(ori_ori_n705_), .Y(ori_ori_n706_));
  NO2        o684(.A(ori_ori_n706_), .B(ori_ori_n699_), .Y(ori_ori_n707_));
  INV        o685(.A(ori_ori_n171_), .Y(ori_ori_n708_));
  INV        o686(.A(ori_ori_n238_), .Y(ori_ori_n709_));
  OAI210     o687(.A0(ori_ori_n646_), .A1(ori_ori_n426_), .B0(ori_ori_n111_), .Y(ori_ori_n710_));
  AOI210     o688(.A0(ori_ori_n710_), .A1(ori_ori_n709_), .B0(ori_ori_n708_), .Y(ori_ori_n711_));
  NO2        o689(.A(ori_ori_n433_), .B(ori_ori_n26_), .Y(ori_ori_n712_));
  NO2        o690(.A(ori_ori_n712_), .B(ori_ori_n401_), .Y(ori_ori_n713_));
  NA2        o691(.A(ori_ori_n713_), .B(i_2_), .Y(ori_ori_n714_));
  INV        o692(.A(ori_ori_n714_), .Y(ori_ori_n715_));
  AOI210     o693(.A0(ori_ori_n33_), .A1(ori_ori_n36_), .B0(ori_ori_n397_), .Y(ori_ori_n716_));
  AOI210     o694(.A0(ori_ori_n716_), .A1(ori_ori_n715_), .B0(ori_ori_n711_), .Y(ori_ori_n717_));
  NO2        o695(.A(ori_ori_n186_), .B(ori_ori_n126_), .Y(ori_ori_n718_));
  OAI210     o696(.A0(ori_ori_n718_), .A1(ori_ori_n701_), .B0(i_2_), .Y(ori_ori_n719_));
  INV        o697(.A(ori_ori_n172_), .Y(ori_ori_n720_));
  NO3        o698(.A(ori_ori_n577_), .B(ori_ori_n38_), .C(ori_ori_n26_), .Y(ori_ori_n721_));
  AOI210     o699(.A0(ori_ori_n720_), .A1(ori_ori_n86_), .B0(ori_ori_n721_), .Y(ori_ori_n722_));
  AOI210     o700(.A0(ori_ori_n722_), .A1(ori_ori_n719_), .B0(ori_ori_n188_), .Y(ori_ori_n723_));
  OA210      o701(.A0(ori_ori_n578_), .A1(ori_ori_n127_), .B0(i_13_), .Y(ori_ori_n724_));
  NA2        o702(.A(ori_ori_n195_), .B(ori_ori_n198_), .Y(ori_ori_n725_));
  NA2        o703(.A(ori_ori_n152_), .B(ori_ori_n555_), .Y(ori_ori_n726_));
  AOI210     o704(.A0(ori_ori_n726_), .A1(ori_ori_n725_), .B0(ori_ori_n356_), .Y(ori_ori_n727_));
  AOI210     o705(.A0(ori_ori_n204_), .A1(ori_ori_n149_), .B0(ori_ori_n485_), .Y(ori_ori_n728_));
  NA2        o706(.A(ori_ori_n728_), .B(ori_ori_n401_), .Y(ori_ori_n729_));
  NO2        o707(.A(ori_ori_n102_), .B(ori_ori_n44_), .Y(ori_ori_n730_));
  INV        o708(.A(ori_ori_n291_), .Y(ori_ori_n731_));
  NA4        o709(.A(ori_ori_n731_), .B(ori_ori_n293_), .C(ori_ori_n125_), .D(ori_ori_n42_), .Y(ori_ori_n732_));
  OAI210     o710(.A0(ori_ori_n732_), .A1(ori_ori_n730_), .B0(ori_ori_n729_), .Y(ori_ori_n733_));
  NO4        o711(.A(ori_ori_n733_), .B(ori_ori_n727_), .C(ori_ori_n724_), .D(ori_ori_n723_), .Y(ori_ori_n734_));
  NA2        o712(.A(ori_ori_n530_), .B(ori_ori_n28_), .Y(ori_ori_n735_));
  NA2        o713(.A(ori_ori_n700_), .B(ori_ori_n267_), .Y(ori_ori_n736_));
  NA2        o714(.A(ori_ori_n736_), .B(ori_ori_n735_), .Y(ori_ori_n737_));
  NO2        o715(.A(ori_ori_n61_), .B(i_12_), .Y(ori_ori_n738_));
  NO2        o716(.A(ori_ori_n738_), .B(ori_ori_n127_), .Y(ori_ori_n739_));
  NO2        o717(.A(ori_ori_n739_), .B(ori_ori_n555_), .Y(ori_ori_n740_));
  AOI220     o718(.A0(ori_ori_n740_), .A1(ori_ori_n36_), .B0(ori_ori_n737_), .B1(ori_ori_n46_), .Y(ori_ori_n741_));
  NA4        o719(.A(ori_ori_n741_), .B(ori_ori_n734_), .C(ori_ori_n717_), .D(ori_ori_n707_), .Y(ori6));
  NO3        o720(.A(i_9_), .B(ori_ori_n294_), .C(i_1_), .Y(ori_ori_n743_));
  NO2        o721(.A(ori_ori_n181_), .B(ori_ori_n140_), .Y(ori_ori_n744_));
  OAI210     o722(.A0(ori_ori_n744_), .A1(ori_ori_n743_), .B0(ori_ori_n688_), .Y(ori_ori_n745_));
  NO2        o723(.A(ori_ori_n216_), .B(ori_ori_n459_), .Y(ori_ori_n746_));
  NO2        o724(.A(i_11_), .B(i_9_), .Y(ori_ori_n747_));
  INV        o725(.A(ori_ori_n312_), .Y(ori_ori_n748_));
  AO210      o726(.A0(ori_ori_n748_), .A1(ori_ori_n745_), .B0(i_12_), .Y(ori_ori_n749_));
  NA2        o727(.A(ori_ori_n538_), .B(ori_ori_n62_), .Y(ori_ori_n750_));
  INV        o728(.A(ori_ori_n750_), .Y(ori_ori_n751_));
  INV        o729(.A(ori_ori_n192_), .Y(ori_ori_n752_));
  AOI220     o730(.A0(ori_ori_n752_), .A1(ori_ori_n747_), .B0(ori_ori_n751_), .B1(ori_ori_n72_), .Y(ori_ori_n753_));
  INV        o731(.A(ori_ori_n311_), .Y(ori_ori_n754_));
  NA2        o732(.A(ori_ori_n74_), .B(ori_ori_n132_), .Y(ori_ori_n755_));
  INV        o733(.A(ori_ori_n125_), .Y(ori_ori_n756_));
  NA2        o734(.A(ori_ori_n756_), .B(ori_ori_n46_), .Y(ori_ori_n757_));
  AOI210     o735(.A0(ori_ori_n757_), .A1(ori_ori_n755_), .B0(ori_ori_n754_), .Y(ori_ori_n758_));
  NO2        o736(.A(ori_ori_n242_), .B(i_9_), .Y(ori_ori_n759_));
  NA2        o737(.A(ori_ori_n759_), .B(ori_ori_n738_), .Y(ori_ori_n760_));
  AOI210     o738(.A0(ori_ori_n760_), .A1(ori_ori_n483_), .B0(ori_ori_n181_), .Y(ori_ori_n761_));
  NO2        o739(.A(ori_ori_n32_), .B(i_11_), .Y(ori_ori_n762_));
  NAi32      o740(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n763_));
  NO2        o741(.A(ori_ori_n675_), .B(ori_ori_n763_), .Y(ori_ori_n764_));
  OAI210     o742(.A0(ori_ori_n639_), .A1(ori_ori_n525_), .B0(ori_ori_n524_), .Y(ori_ori_n765_));
  NAi21      o743(.An(ori_ori_n764_), .B(ori_ori_n765_), .Y(ori_ori_n766_));
  OR3        o744(.A(ori_ori_n766_), .B(ori_ori_n761_), .C(ori_ori_n758_), .Y(ori_ori_n767_));
  NO2        o745(.A(ori_ori_n651_), .B(i_2_), .Y(ori_ori_n768_));
  NA2        o746(.A(ori_ori_n48_), .B(ori_ori_n37_), .Y(ori_ori_n769_));
  NO2        o747(.A(ori_ori_n769_), .B(ori_ori_n394_), .Y(ori_ori_n770_));
  NA2        o748(.A(ori_ori_n770_), .B(ori_ori_n768_), .Y(ori_ori_n771_));
  AO220      o749(.A0(ori_ori_n340_), .A1(ori_ori_n330_), .B0(ori_ori_n382_), .B1(ori_ori_n555_), .Y(ori_ori_n772_));
  NA3        o750(.A(ori_ori_n772_), .B(ori_ori_n245_), .C(i_7_), .Y(ori_ori_n773_));
  OR2        o751(.A(ori_ori_n578_), .B(ori_ori_n426_), .Y(ori_ori_n774_));
  NA3        o752(.A(ori_ori_n774_), .B(ori_ori_n148_), .C(ori_ori_n68_), .Y(ori_ori_n775_));
  AO210      o753(.A0(ori_ori_n466_), .A1(ori_ori_n704_), .B0(ori_ori_n36_), .Y(ori_ori_n776_));
  NA4        o754(.A(ori_ori_n776_), .B(ori_ori_n775_), .C(ori_ori_n773_), .D(ori_ori_n771_), .Y(ori_ori_n777_));
  NO2        o755(.A(ori_ori_n595_), .B(i_11_), .Y(ori_ori_n778_));
  AOI220     o756(.A0(ori_ori_n778_), .A1(ori_ori_n524_), .B0(ori_ori_n746_), .B1(ori_ori_n669_), .Y(ori_ori_n779_));
  NA3        o757(.A(ori_ori_n356_), .B(ori_ori_n231_), .C(ori_ori_n148_), .Y(ori_ori_n780_));
  NA2        o758(.A(ori_ori_n382_), .B(ori_ori_n69_), .Y(ori_ori_n781_));
  NA4        o759(.A(ori_ori_n781_), .B(ori_ori_n780_), .C(ori_ori_n779_), .D(ori_ori_n563_), .Y(ori_ori_n782_));
  NA2        o760(.A(ori_ori_n426_), .B(ori_ori_n424_), .Y(ori_ori_n783_));
  NO2        o761(.A(ori_ori_n571_), .B(ori_ori_n102_), .Y(ori_ori_n784_));
  OAI210     o762(.A0(ori_ori_n784_), .A1(ori_ori_n112_), .B0(ori_ori_n393_), .Y(ori_ori_n785_));
  NA2        o763(.A(ori_ori_n237_), .B(ori_ori_n46_), .Y(ori_ori_n786_));
  INV        o764(.A(ori_ori_n544_), .Y(ori_ori_n787_));
  NA3        o765(.A(ori_ori_n787_), .B(ori_ori_n311_), .C(i_7_), .Y(ori_ori_n788_));
  NA3        o766(.A(ori_ori_n788_), .B(ori_ori_n785_), .C(ori_ori_n783_), .Y(ori_ori_n789_));
  NO4        o767(.A(ori_ori_n789_), .B(ori_ori_n782_), .C(ori_ori_n777_), .D(ori_ori_n767_), .Y(ori_ori_n790_));
  NA4        o768(.A(ori_ori_n790_), .B(ori_ori_n753_), .C(ori_ori_n749_), .D(ori_ori_n364_), .Y(ori3));
  NA2        o769(.A(i_12_), .B(i_10_), .Y(ori_ori_n792_));
  NO2        o770(.A(i_11_), .B(ori_ori_n229_), .Y(ori_ori_n793_));
  NA2        o771(.A(ori_ori_n780_), .B(ori_ori_n563_), .Y(ori_ori_n794_));
  NA2        o772(.A(ori_ori_n794_), .B(ori_ori_n40_), .Y(ori_ori_n795_));
  NOi21      o773(.An(ori_ori_n96_), .B(ori_ori_n713_), .Y(ori_ori_n796_));
  NO3        o774(.A(ori_ori_n585_), .B(ori_ori_n433_), .C(ori_ori_n132_), .Y(ori_ori_n797_));
  NA2        o775(.A(ori_ori_n395_), .B(ori_ori_n45_), .Y(ori_ori_n798_));
  AN2        o776(.A(ori_ori_n431_), .B(ori_ori_n55_), .Y(ori_ori_n799_));
  NO3        o777(.A(ori_ori_n799_), .B(ori_ori_n797_), .C(ori_ori_n796_), .Y(ori_ori_n800_));
  AOI210     o778(.A0(ori_ori_n800_), .A1(ori_ori_n795_), .B0(ori_ori_n48_), .Y(ori_ori_n801_));
  NO4        o779(.A(ori_ori_n360_), .B(ori_ori_n367_), .C(ori_ori_n38_), .D(i_0_), .Y(ori_ori_n802_));
  NA2        o780(.A(ori_ori_n181_), .B(ori_ori_n528_), .Y(ori_ori_n803_));
  NOi21      o781(.An(ori_ori_n803_), .B(ori_ori_n802_), .Y(ori_ori_n804_));
  NA2        o782(.A(ori_ori_n663_), .B(ori_ori_n629_), .Y(ori_ori_n805_));
  NA2        o783(.A(ori_ori_n318_), .B(ori_ori_n419_), .Y(ori_ori_n806_));
  OAI220     o784(.A0(ori_ori_n806_), .A1(ori_ori_n805_), .B0(ori_ori_n804_), .B1(ori_ori_n62_), .Y(ori_ori_n807_));
  NOi21      o785(.An(i_5_), .B(i_9_), .Y(ori_ori_n808_));
  NA2        o786(.A(ori_ori_n808_), .B(ori_ori_n423_), .Y(ori_ori_n809_));
  BUFFER     o787(.A(ori_ori_n257_), .Y(ori_ori_n810_));
  NA2        o788(.A(ori_ori_n810_), .B(ori_ori_n451_), .Y(ori_ori_n811_));
  NO2        o789(.A(ori_ori_n811_), .B(ori_ori_n809_), .Y(ori_ori_n812_));
  NO3        o790(.A(ori_ori_n812_), .B(ori_ori_n807_), .C(ori_ori_n801_), .Y(ori_ori_n813_));
  NA2        o791(.A(ori_ori_n181_), .B(ori_ori_n24_), .Y(ori_ori_n814_));
  NO2        o792(.A(ori_ori_n627_), .B(ori_ori_n552_), .Y(ori_ori_n815_));
  NO2        o793(.A(ori_ori_n815_), .B(ori_ori_n814_), .Y(ori_ori_n816_));
  NA2        o794(.A(ori_ori_n298_), .B(ori_ori_n130_), .Y(ori_ori_n817_));
  NAi21      o795(.An(ori_ori_n163_), .B(ori_ori_n419_), .Y(ori_ori_n818_));
  OAI220     o796(.A0(ori_ori_n818_), .A1(ori_ori_n786_), .B0(ori_ori_n817_), .B1(ori_ori_n387_), .Y(ori_ori_n819_));
  NO2        o797(.A(ori_ori_n819_), .B(ori_ori_n816_), .Y(ori_ori_n820_));
  NA2        o798(.A(ori_ori_n529_), .B(i_0_), .Y(ori_ori_n821_));
  NO3        o799(.A(ori_ori_n821_), .B(ori_ori_n369_), .C(ori_ori_n86_), .Y(ori_ori_n822_));
  NO4        o800(.A(ori_ori_n543_), .B(ori_ori_n210_), .C(ori_ori_n397_), .D(ori_ori_n394_), .Y(ori_ori_n823_));
  AOI210     o801(.A0(ori_ori_n823_), .A1(i_11_), .B0(ori_ori_n822_), .Y(ori_ori_n824_));
  INV        o802(.A(ori_ori_n450_), .Y(ori_ori_n825_));
  AN2        o803(.A(ori_ori_n96_), .B(ori_ori_n236_), .Y(ori_ori_n826_));
  NA2        o804(.A(ori_ori_n700_), .B(ori_ori_n312_), .Y(ori_ori_n827_));
  AOI210     o805(.A0(ori_ori_n455_), .A1(ori_ori_n86_), .B0(ori_ori_n57_), .Y(ori_ori_n828_));
  OAI220     o806(.A0(ori_ori_n828_), .A1(ori_ori_n827_), .B0(ori_ori_n614_), .B1(ori_ori_n500_), .Y(ori_ori_n829_));
  NO2        o807(.A(ori_ori_n244_), .B(ori_ori_n154_), .Y(ori_ori_n830_));
  NA2        o808(.A(i_0_), .B(i_10_), .Y(ori_ori_n831_));
  INV        o809(.A(ori_ori_n503_), .Y(ori_ori_n832_));
  NO4        o810(.A(ori_ori_n115_), .B(ori_ori_n57_), .C(ori_ori_n624_), .D(i_5_), .Y(ori_ori_n833_));
  AO220      o811(.A0(ori_ori_n833_), .A1(ori_ori_n832_), .B0(ori_ori_n830_), .B1(i_6_), .Y(ori_ori_n834_));
  NO3        o812(.A(ori_ori_n834_), .B(ori_ori_n829_), .C(ori_ori_n826_), .Y(ori_ori_n835_));
  NA3        o813(.A(ori_ori_n835_), .B(ori_ori_n824_), .C(ori_ori_n820_), .Y(ori_ori_n836_));
  NA2        o814(.A(i_11_), .B(i_9_), .Y(ori_ori_n837_));
  NA2        o815(.A(ori_ori_n379_), .B(ori_ori_n175_), .Y(ori_ori_n838_));
  NA2        o816(.A(ori_ori_n838_), .B(ori_ori_n161_), .Y(ori_ori_n839_));
  NO2        o817(.A(ori_ori_n837_), .B(ori_ori_n72_), .Y(ori_ori_n840_));
  NO2        o818(.A(ori_ori_n174_), .B(i_0_), .Y(ori_ori_n841_));
  INV        o819(.A(ori_ori_n841_), .Y(ori_ori_n842_));
  NA2        o820(.A(ori_ori_n450_), .B(ori_ori_n223_), .Y(ori_ori_n843_));
  NO2        o821(.A(ori_ori_n843_), .B(ori_ori_n842_), .Y(ori_ori_n844_));
  NO2        o822(.A(ori_ori_n844_), .B(ori_ori_n839_), .Y(ori_ori_n845_));
  NA2        o823(.A(ori_ori_n613_), .B(ori_ori_n122_), .Y(ori_ori_n846_));
  NO2        o824(.A(i_6_), .B(ori_ori_n846_), .Y(ori_ori_n847_));
  AOI210     o825(.A0(ori_ori_n425_), .A1(ori_ori_n36_), .B0(i_3_), .Y(ori_ori_n848_));
  NA2        o826(.A(ori_ori_n171_), .B(ori_ori_n103_), .Y(ori_ori_n849_));
  NOi32      o827(.An(ori_ori_n848_), .Bn(ori_ori_n184_), .C(ori_ori_n849_), .Y(ori_ori_n850_));
  NA2        o828(.A(ori_ori_n564_), .B(ori_ori_n312_), .Y(ori_ori_n851_));
  NO2        o829(.A(ori_ori_n851_), .B(ori_ori_n798_), .Y(ori_ori_n852_));
  NO3        o830(.A(ori_ori_n852_), .B(ori_ori_n850_), .C(ori_ori_n847_), .Y(ori_ori_n853_));
  INV        o831(.A(ori_ori_n303_), .Y(ori_ori_n854_));
  NA2        o832(.A(ori_ori_n853_), .B(ori_ori_n845_), .Y(ori_ori_n855_));
  NO2        o833(.A(ori_ori_n792_), .B(ori_ori_n302_), .Y(ori_ori_n856_));
  NA2        o834(.A(ori_ori_n856_), .B(ori_ori_n840_), .Y(ori_ori_n857_));
  NA3        o835(.A(ori_ori_n449_), .B(ori_ori_n395_), .C(ori_ori_n45_), .Y(ori_ori_n858_));
  OAI210     o836(.A0(ori_ori_n818_), .A1(ori_ori_n825_), .B0(ori_ori_n858_), .Y(ori_ori_n859_));
  NA2        o837(.A(ori_ori_n840_), .B(ori_ori_n293_), .Y(ori_ori_n860_));
  NA2        o838(.A(ori_ori_n183_), .B(ori_ori_n860_), .Y(ori_ori_n861_));
  AOI220     o839(.A0(ori_ori_n861_), .A1(ori_ori_n450_), .B0(ori_ori_n859_), .B1(ori_ori_n72_), .Y(ori_ori_n862_));
  NA3        o840(.A(ori_ori_n769_), .B(ori_ori_n366_), .C(ori_ori_n595_), .Y(ori_ori_n863_));
  NA2        o841(.A(ori_ori_n92_), .B(ori_ori_n44_), .Y(ori_ori_n864_));
  NO2        o842(.A(ori_ori_n74_), .B(ori_ori_n702_), .Y(ori_ori_n865_));
  AOI220     o843(.A0(ori_ori_n865_), .A1(ori_ori_n864_), .B0(ori_ori_n173_), .B1(ori_ori_n552_), .Y(ori_ori_n866_));
  AOI210     o844(.A0(ori_ori_n866_), .A1(ori_ori_n863_), .B0(ori_ori_n47_), .Y(ori_ori_n867_));
  NO3        o845(.A(ori_ori_n543_), .B(ori_ori_n338_), .C(ori_ori_n24_), .Y(ori_ori_n868_));
  AOI210     o846(.A0(ori_ori_n656_), .A1(ori_ori_n512_), .B0(ori_ori_n868_), .Y(ori_ori_n869_));
  NAi21      o847(.An(i_9_), .B(i_5_), .Y(ori_ori_n870_));
  NO2        o848(.A(ori_ori_n869_), .B(ori_ori_n172_), .Y(ori_ori_n871_));
  NO3        o849(.A(ori_ori_n871_), .B(ori_ori_n867_), .C(ori_ori_n487_), .Y(ori_ori_n872_));
  NA3        o850(.A(ori_ori_n872_), .B(ori_ori_n862_), .C(ori_ori_n857_), .Y(ori_ori_n873_));
  NO3        o851(.A(ori_ori_n873_), .B(ori_ori_n855_), .C(ori_ori_n836_), .Y(ori_ori_n874_));
  NO2        o852(.A(i_0_), .B(ori_ori_n680_), .Y(ori_ori_n875_));
  NA2        o853(.A(ori_ori_n72_), .B(ori_ori_n44_), .Y(ori_ori_n876_));
  AOI210     o854(.A0(ori_ori_n750_), .A1(ori_ori_n640_), .B0(ori_ori_n849_), .Y(ori_ori_n877_));
  INV        o855(.A(ori_ori_n877_), .Y(ori_ori_n878_));
  NO2        o856(.A(ori_ori_n765_), .B(ori_ori_n388_), .Y(ori_ori_n879_));
  NA2        o857(.A(ori_ori_n793_), .B(i_9_), .Y(ori_ori_n880_));
  NO2        o858(.A(ori_ori_n470_), .B(ori_ori_n880_), .Y(ori_ori_n881_));
  NA2        o859(.A(ori_ori_n237_), .B(ori_ori_n222_), .Y(ori_ori_n882_));
  AOI210     o860(.A0(ori_ori_n882_), .A1(ori_ori_n821_), .B0(ori_ori_n154_), .Y(ori_ori_n883_));
  NO3        o861(.A(ori_ori_n883_), .B(ori_ori_n881_), .C(ori_ori_n879_), .Y(ori_ori_n884_));
  NA2        o862(.A(ori_ori_n884_), .B(ori_ori_n878_), .Y(ori_ori_n885_));
  NO3        o863(.A(ori_ori_n831_), .B(ori_ori_n808_), .C(ori_ori_n186_), .Y(ori_ori_n886_));
  AOI220     o864(.A0(ori_ori_n886_), .A1(i_11_), .B0(ori_ori_n527_), .B1(ori_ori_n74_), .Y(ori_ori_n887_));
  NO3        o865(.A(ori_ori_n205_), .B(ori_ori_n367_), .C(i_0_), .Y(ori_ori_n888_));
  OAI210     o866(.A0(ori_ori_n888_), .A1(ori_ori_n75_), .B0(i_13_), .Y(ori_ori_n889_));
  INV        o867(.A(ori_ori_n213_), .Y(ori_ori_n890_));
  OAI220     o868(.A0(ori_ori_n497_), .A1(ori_ori_n140_), .B0(ori_ori_n598_), .B1(ori_ori_n573_), .Y(ori_ori_n891_));
  NA3        o869(.A(ori_ori_n891_), .B(i_7_), .C(ori_ori_n890_), .Y(ori_ori_n892_));
  NA3        o870(.A(ori_ori_n892_), .B(ori_ori_n889_), .C(ori_ori_n887_), .Y(ori_ori_n893_));
  NO2        o871(.A(ori_ori_n235_), .B(ori_ori_n92_), .Y(ori_ori_n894_));
  AOI210     o872(.A0(ori_ori_n894_), .A1(ori_ori_n875_), .B0(ori_ori_n109_), .Y(ori_ori_n895_));
  OR2        o873(.A(ori_ori_n895_), .B(i_5_), .Y(ori_ori_n896_));
  INV        o874(.A(ori_ori_n510_), .Y(ori_ori_n897_));
  NO3        o875(.A(ori_ori_n798_), .B(ori_ori_n54_), .C(ori_ori_n48_), .Y(ori_ori_n898_));
  NA2        o876(.A(ori_ori_n465_), .B(ori_ori_n458_), .Y(ori_ori_n899_));
  NO3        o877(.A(ori_ori_n899_), .B(ori_ori_n898_), .C(ori_ori_n897_), .Y(ori_ori_n900_));
  NA3        o878(.A(ori_ori_n374_), .B(ori_ori_n171_), .C(ori_ori_n170_), .Y(ori_ori_n901_));
  INV        o879(.A(ori_ori_n901_), .Y(ori_ori_n902_));
  NA3        o880(.A(ori_ori_n374_), .B(ori_ori_n319_), .C(ori_ori_n217_), .Y(ori_ori_n903_));
  INV        o881(.A(ori_ori_n903_), .Y(ori_ori_n904_));
  NOi31      o882(.An(ori_ori_n373_), .B(ori_ori_n876_), .C(ori_ori_n232_), .Y(ori_ori_n905_));
  NO3        o883(.A(ori_ori_n837_), .B(ori_ori_n213_), .C(ori_ori_n186_), .Y(ori_ori_n906_));
  NO4        o884(.A(ori_ori_n906_), .B(ori_ori_n905_), .C(ori_ori_n904_), .D(ori_ori_n902_), .Y(ori_ori_n907_));
  NA3        o885(.A(ori_ori_n907_), .B(ori_ori_n900_), .C(ori_ori_n896_), .Y(ori_ori_n908_));
  NO2        o886(.A(ori_ori_n85_), .B(i_5_), .Y(ori_ori_n909_));
  NA3        o887(.A(ori_ori_n793_), .B(ori_ori_n110_), .C(ori_ori_n125_), .Y(ori_ori_n910_));
  INV        o888(.A(ori_ori_n910_), .Y(ori_ori_n911_));
  NA2        o889(.A(ori_ori_n911_), .B(ori_ori_n909_), .Y(ori_ori_n912_));
  NAi21      o890(.An(ori_ori_n234_), .B(ori_ori_n235_), .Y(ori_ori_n913_));
  NO4        o891(.A(ori_ori_n232_), .B(ori_ori_n205_), .C(i_0_), .D(i_12_), .Y(ori_ori_n914_));
  NA2        o892(.A(ori_ori_n914_), .B(ori_ori_n913_), .Y(ori_ori_n915_));
  AN2        o893(.A(ori_ori_n831_), .B(ori_ori_n154_), .Y(ori_ori_n916_));
  NO4        o894(.A(ori_ori_n916_), .B(i_12_), .C(ori_ori_n602_), .D(ori_ori_n132_), .Y(ori_ori_n917_));
  NA2        o895(.A(ori_ori_n917_), .B(ori_ori_n213_), .Y(ori_ori_n918_));
  NA3        o896(.A(ori_ori_n98_), .B(ori_ori_n528_), .C(i_11_), .Y(ori_ori_n919_));
  NO2        o897(.A(ori_ori_n919_), .B(ori_ori_n156_), .Y(ori_ori_n920_));
  INV        o898(.A(ori_ori_n920_), .Y(ori_ori_n921_));
  NA4        o899(.A(ori_ori_n921_), .B(ori_ori_n918_), .C(ori_ori_n915_), .D(ori_ori_n912_), .Y(ori_ori_n922_));
  NO4        o900(.A(ori_ori_n922_), .B(ori_ori_n908_), .C(ori_ori_n893_), .D(ori_ori_n885_), .Y(ori_ori_n923_));
  OAI210     o901(.A0(ori_ori_n768_), .A1(ori_ori_n762_), .B0(ori_ori_n37_), .Y(ori_ori_n924_));
  NA3        o902(.A(ori_ori_n848_), .B(ori_ori_n351_), .C(i_5_), .Y(ori_ori_n925_));
  NA3        o903(.A(ori_ori_n925_), .B(ori_ori_n924_), .C(ori_ori_n570_), .Y(ori_ori_n926_));
  NA2        o904(.A(ori_ori_n926_), .B(ori_ori_n203_), .Y(ori_ori_n927_));
  AN2        o905(.A(ori_ori_n651_), .B(ori_ori_n352_), .Y(ori_ori_n928_));
  NA2        o906(.A(ori_ori_n182_), .B(ori_ori_n184_), .Y(ori_ori_n929_));
  AO210      o907(.A0(ori_ori_n928_), .A1(ori_ori_n33_), .B0(ori_ori_n929_), .Y(ori_ori_n930_));
  INV        o908(.A(ori_ori_n930_), .Y(ori_ori_n931_));
  INV        o909(.A(ori_ori_n823_), .Y(ori_ori_n932_));
  OAI210     o910(.A0(ori_ori_n919_), .A1(ori_ori_n149_), .B0(ori_ori_n932_), .Y(ori_ori_n933_));
  AOI210     o911(.A0(ori_ori_n931_), .A1(ori_ori_n48_), .B0(ori_ori_n933_), .Y(ori_ori_n934_));
  AOI210     o912(.A0(ori_ori_n934_), .A1(ori_ori_n927_), .B0(ori_ori_n72_), .Y(ori_ori_n935_));
  INV        o913(.A(ori_ori_n363_), .Y(ori_ori_n936_));
  NO2        o914(.A(ori_ori_n936_), .B(ori_ori_n708_), .Y(ori_ori_n937_));
  OAI210     o915(.A0(ori_ori_n79_), .A1(ori_ori_n54_), .B0(ori_ori_n108_), .Y(ori_ori_n938_));
  NA2        o916(.A(ori_ori_n938_), .B(ori_ori_n75_), .Y(ori_ori_n939_));
  NO2        o917(.A(ori_ori_n939_), .B(ori_ori_n633_), .Y(ori_ori_n940_));
  INV        o918(.A(ori_ori_n940_), .Y(ori_ori_n941_));
  OAI210     o919(.A0(ori_ori_n259_), .A1(ori_ori_n159_), .B0(ori_ori_n86_), .Y(ori_ori_n942_));
  NA3        o920(.A(ori_ori_n712_), .B(ori_ori_n282_), .C(ori_ori_n79_), .Y(ori_ori_n943_));
  AOI210     o921(.A0(ori_ori_n943_), .A1(ori_ori_n942_), .B0(i_11_), .Y(ori_ori_n944_));
  OAI210     o922(.A0(ori_ori_n962_), .A1(ori_ori_n848_), .B0(ori_ori_n203_), .Y(ori_ori_n945_));
  NA2        o923(.A(ori_ori_n165_), .B(i_5_), .Y(ori_ori_n946_));
  NO2        o924(.A(ori_ori_n945_), .B(ori_ori_n946_), .Y(ori_ori_n947_));
  NO3        o925(.A(ori_ori_n58_), .B(ori_ori_n57_), .C(i_4_), .Y(ori_ori_n948_));
  OAI210     o926(.A0(ori_ori_n854_), .A1(ori_ori_n294_), .B0(ori_ori_n948_), .Y(ori_ori_n949_));
  NO2        o927(.A(ori_ori_n949_), .B(ori_ori_n680_), .Y(ori_ori_n950_));
  NO4        o928(.A(ori_ori_n870_), .B(ori_ori_n452_), .C(ori_ori_n243_), .D(ori_ori_n242_), .Y(ori_ori_n951_));
  INV        o929(.A(ori_ori_n951_), .Y(ori_ori_n952_));
  INV        o930(.A(ori_ori_n344_), .Y(ori_ori_n953_));
  AOI210     o931(.A0(ori_ori_n953_), .A1(ori_ori_n952_), .B0(ori_ori_n41_), .Y(ori_ori_n954_));
  NO4        o932(.A(ori_ori_n954_), .B(ori_ori_n950_), .C(ori_ori_n947_), .D(ori_ori_n944_), .Y(ori_ori_n955_));
  OAI210     o933(.A0(ori_ori_n941_), .A1(i_4_), .B0(ori_ori_n955_), .Y(ori_ori_n956_));
  NO3        o934(.A(ori_ori_n956_), .B(ori_ori_n937_), .C(ori_ori_n935_), .Y(ori_ori_n957_));
  NA4        o935(.A(ori_ori_n957_), .B(ori_ori_n923_), .C(ori_ori_n874_), .D(ori_ori_n813_), .Y(ori4));
  INV        o936(.A(ori_ori_n655_), .Y(ori_ori_n961_));
  INV        o937(.A(i_12_), .Y(ori_ori_n962_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NAi21      m015(.An(i_11_), .B(i_9_), .Y(mai_mai_n38_));
  NO3        m016(.A(mai_mai_n38_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n39_));
  NOi21      m017(.An(i_12_), .B(i_13_), .Y(mai_mai_n40_));
  INV        m018(.A(mai_mai_n40_), .Y(mai_mai_n41_));
  NO2        m019(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n42_));
  NAi31      m020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n43_));
  INV        m021(.A(mai_mai_n35_), .Y(mai1));
  INV        m022(.A(i_11_), .Y(mai_mai_n45_));
  NO2        m023(.A(mai_mai_n45_), .B(i_6_), .Y(mai_mai_n46_));
  INV        m024(.A(i_2_), .Y(mai_mai_n47_));
  NA2        m025(.A(i_0_), .B(i_3_), .Y(mai_mai_n48_));
  INV        m026(.A(i_5_), .Y(mai_mai_n49_));
  NO2        m027(.A(i_7_), .B(i_10_), .Y(mai_mai_n50_));
  AOI210     m028(.A0(i_7_), .A1(mai_mai_n25_), .B0(mai_mai_n50_), .Y(mai_mai_n51_));
  OAI210     m029(.A0(mai_mai_n51_), .A1(i_3_), .B0(mai_mai_n49_), .Y(mai_mai_n52_));
  AOI210     m030(.A0(mai_mai_n52_), .A1(mai_mai_n48_), .B0(mai_mai_n47_), .Y(mai_mai_n53_));
  NA2        m031(.A(i_0_), .B(i_2_), .Y(mai_mai_n54_));
  NA2        m032(.A(i_7_), .B(i_9_), .Y(mai_mai_n55_));
  NO2        m033(.A(mai_mai_n55_), .B(mai_mai_n54_), .Y(mai_mai_n56_));
  NA2        m034(.A(mai_mai_n53_), .B(mai_mai_n46_), .Y(mai_mai_n57_));
  NA3        m035(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n58_));
  NO2        m036(.A(i_1_), .B(i_6_), .Y(mai_mai_n59_));
  NA2        m037(.A(i_8_), .B(i_7_), .Y(mai_mai_n60_));
  OAI210     m038(.A0(mai_mai_n60_), .A1(mai_mai_n59_), .B0(mai_mai_n58_), .Y(mai_mai_n61_));
  NA2        m039(.A(mai_mai_n61_), .B(i_12_), .Y(mai_mai_n62_));
  NAi21      m040(.An(i_2_), .B(i_7_), .Y(mai_mai_n63_));
  INV        m041(.A(i_1_), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(i_6_), .Y(mai_mai_n65_));
  NA3        m043(.A(mai_mai_n65_), .B(mai_mai_n63_), .C(mai_mai_n31_), .Y(mai_mai_n66_));
  NA2        m044(.A(i_1_), .B(i_10_), .Y(mai_mai_n67_));
  NO2        m045(.A(mai_mai_n67_), .B(i_6_), .Y(mai_mai_n68_));
  NAi31      m046(.An(mai_mai_n68_), .B(mai_mai_n66_), .C(mai_mai_n62_), .Y(mai_mai_n69_));
  NA2        m047(.A(mai_mai_n51_), .B(i_2_), .Y(mai_mai_n70_));
  AOI210     m048(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_1_), .B(i_6_), .Y(mai_mai_n72_));
  NO2        m050(.A(mai_mai_n72_), .B(mai_mai_n25_), .Y(mai_mai_n73_));
  INV        m051(.A(i_0_), .Y(mai_mai_n74_));
  NAi21      m052(.An(i_5_), .B(i_10_), .Y(mai_mai_n75_));
  NA2        m053(.A(i_5_), .B(i_9_), .Y(mai_mai_n76_));
  AOI210     m054(.A0(mai_mai_n76_), .A1(mai_mai_n75_), .B0(mai_mai_n74_), .Y(mai_mai_n77_));
  NO2        m055(.A(mai_mai_n77_), .B(mai_mai_n73_), .Y(mai_mai_n78_));
  OAI210     m056(.A0(mai_mai_n71_), .A1(mai_mai_n70_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  OAI210     m057(.A0(mai_mai_n79_), .A1(mai_mai_n69_), .B0(i_0_), .Y(mai_mai_n80_));
  NA2        m058(.A(i_12_), .B(i_5_), .Y(mai_mai_n81_));
  NA2        m059(.A(i_2_), .B(i_8_), .Y(mai_mai_n82_));
  NO2        m060(.A(mai_mai_n82_), .B(mai_mai_n59_), .Y(mai_mai_n83_));
  NO2        m061(.A(i_3_), .B(i_9_), .Y(mai_mai_n84_));
  NO2        m062(.A(i_3_), .B(i_7_), .Y(mai_mai_n85_));
  NO3        m063(.A(mai_mai_n85_), .B(mai_mai_n84_), .C(mai_mai_n64_), .Y(mai_mai_n86_));
  INV        m064(.A(i_6_), .Y(mai_mai_n87_));
  OR4        m065(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n88_));
  INV        m066(.A(mai_mai_n88_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_2_), .B(i_7_), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n89_), .B(mai_mai_n90_), .Y(mai_mai_n91_));
  OAI210     m069(.A0(mai_mai_n86_), .A1(mai_mai_n83_), .B0(mai_mai_n91_), .Y(mai_mai_n92_));
  NAi21      m070(.An(i_6_), .B(i_10_), .Y(mai_mai_n93_));
  NA2        m071(.A(i_6_), .B(i_9_), .Y(mai_mai_n94_));
  AOI210     m072(.A0(mai_mai_n94_), .A1(mai_mai_n93_), .B0(mai_mai_n64_), .Y(mai_mai_n95_));
  NA2        m073(.A(i_2_), .B(i_6_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n50_), .C(mai_mai_n25_), .Y(mai_mai_n97_));
  NO2        m075(.A(mai_mai_n97_), .B(mai_mai_n95_), .Y(mai_mai_n98_));
  AOI210     m076(.A0(mai_mai_n98_), .A1(mai_mai_n92_), .B0(mai_mai_n81_), .Y(mai_mai_n99_));
  AN3        m077(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n100_));
  NAi21      m078(.An(i_6_), .B(i_11_), .Y(mai_mai_n101_));
  NO2        m079(.A(i_5_), .B(i_8_), .Y(mai_mai_n102_));
  NOi21      m080(.An(mai_mai_n102_), .B(mai_mai_n101_), .Y(mai_mai_n103_));
  AOI220     m081(.A0(mai_mai_n103_), .A1(mai_mai_n63_), .B0(mai_mai_n100_), .B1(mai_mai_n32_), .Y(mai_mai_n104_));
  INV        m082(.A(i_7_), .Y(mai_mai_n105_));
  NA2        m083(.A(mai_mai_n47_), .B(mai_mai_n105_), .Y(mai_mai_n106_));
  NO2        m084(.A(i_0_), .B(i_5_), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n107_), .B(mai_mai_n87_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_12_), .B(i_3_), .Y(mai_mai_n109_));
  INV        m087(.A(mai_mai_n109_), .Y(mai_mai_n110_));
  NA3        m088(.A(mai_mai_n110_), .B(mai_mai_n108_), .C(mai_mai_n106_), .Y(mai_mai_n111_));
  NAi21      m089(.An(i_7_), .B(i_11_), .Y(mai_mai_n112_));
  AN2        m090(.A(i_2_), .B(i_10_), .Y(mai_mai_n113_));
  NO2        m091(.A(mai_mai_n113_), .B(i_7_), .Y(mai_mai_n114_));
  OR2        m092(.A(mai_mai_n81_), .B(mai_mai_n59_), .Y(mai_mai_n115_));
  NO2        m093(.A(i_8_), .B(mai_mai_n105_), .Y(mai_mai_n116_));
  NO3        m094(.A(mai_mai_n116_), .B(mai_mai_n115_), .C(mai_mai_n114_), .Y(mai_mai_n117_));
  NA2        m095(.A(i_12_), .B(i_7_), .Y(mai_mai_n118_));
  NO2        m096(.A(mai_mai_n64_), .B(mai_mai_n26_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(i_0_), .Y(mai_mai_n120_));
  NA2        m098(.A(i_11_), .B(i_12_), .Y(mai_mai_n121_));
  OAI210     m099(.A0(mai_mai_n120_), .A1(mai_mai_n118_), .B0(mai_mai_n121_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n122_), .B(mai_mai_n117_), .Y(mai_mai_n123_));
  NA3        m101(.A(mai_mai_n123_), .B(mai_mai_n111_), .C(mai_mai_n104_), .Y(mai_mai_n124_));
  NOi21      m102(.An(i_1_), .B(i_5_), .Y(mai_mai_n125_));
  NA2        m103(.A(mai_mai_n125_), .B(i_11_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n105_), .B(mai_mai_n37_), .Y(mai_mai_n127_));
  NA2        m105(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n128_));
  NA2        m106(.A(mai_mai_n128_), .B(mai_mai_n127_), .Y(mai_mai_n129_));
  NO2        m107(.A(mai_mai_n129_), .B(mai_mai_n47_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n94_), .B(mai_mai_n93_), .Y(mai_mai_n131_));
  NAi21      m109(.An(i_3_), .B(i_8_), .Y(mai_mai_n132_));
  NA2        m110(.A(mai_mai_n132_), .B(mai_mai_n63_), .Y(mai_mai_n133_));
  NOi31      m111(.An(mai_mai_n133_), .B(mai_mai_n131_), .C(mai_mai_n130_), .Y(mai_mai_n134_));
  NO2        m112(.A(i_1_), .B(mai_mai_n87_), .Y(mai_mai_n135_));
  NO2        m113(.A(i_6_), .B(i_5_), .Y(mai_mai_n136_));
  NA2        m114(.A(mai_mai_n136_), .B(i_3_), .Y(mai_mai_n137_));
  AO210      m115(.A0(mai_mai_n137_), .A1(mai_mai_n48_), .B0(mai_mai_n135_), .Y(mai_mai_n138_));
  OAI220     m116(.A0(mai_mai_n138_), .A1(mai_mai_n112_), .B0(mai_mai_n134_), .B1(mai_mai_n126_), .Y(mai_mai_n139_));
  NO3        m117(.A(mai_mai_n139_), .B(mai_mai_n124_), .C(mai_mai_n99_), .Y(mai_mai_n140_));
  NA3        m118(.A(mai_mai_n140_), .B(mai_mai_n80_), .C(mai_mai_n57_), .Y(mai2));
  NO2        m119(.A(mai_mai_n64_), .B(mai_mai_n37_), .Y(mai_mai_n142_));
  INV        m120(.A(i_6_), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NA4        m122(.A(mai_mai_n144_), .B(mai_mai_n78_), .C(mai_mai_n70_), .D(mai_mai_n30_), .Y(mai0));
  AN2        m123(.A(i_8_), .B(i_7_), .Y(mai_mai_n146_));
  NA2        m124(.A(mai_mai_n146_), .B(i_6_), .Y(mai_mai_n147_));
  NO2        m125(.A(i_12_), .B(i_13_), .Y(mai_mai_n148_));
  NAi21      m126(.An(i_5_), .B(i_11_), .Y(mai_mai_n149_));
  NOi21      m127(.An(mai_mai_n148_), .B(mai_mai_n149_), .Y(mai_mai_n150_));
  NO2        m128(.A(i_0_), .B(i_1_), .Y(mai_mai_n151_));
  NA2        m129(.A(i_2_), .B(i_3_), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n152_), .B(i_4_), .Y(mai_mai_n153_));
  NA3        m131(.A(mai_mai_n153_), .B(mai_mai_n151_), .C(mai_mai_n150_), .Y(mai_mai_n154_));
  OR2        m132(.A(mai_mai_n154_), .B(mai_mai_n25_), .Y(mai_mai_n155_));
  AN2        m133(.A(mai_mai_n148_), .B(mai_mai_n84_), .Y(mai_mai_n156_));
  NA2        m134(.A(i_1_), .B(i_5_), .Y(mai_mai_n157_));
  OR2        m135(.A(i_0_), .B(i_1_), .Y(mai_mai_n158_));
  NAi32      m136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n159_));
  NOi21      m137(.An(i_4_), .B(i_10_), .Y(mai_mai_n160_));
  NA2        m138(.A(mai_mai_n160_), .B(mai_mai_n40_), .Y(mai_mai_n161_));
  NO2        m139(.A(i_3_), .B(i_5_), .Y(mai_mai_n162_));
  NO3        m140(.A(mai_mai_n74_), .B(i_2_), .C(i_1_), .Y(mai_mai_n163_));
  NA2        m141(.A(mai_mai_n163_), .B(mai_mai_n162_), .Y(mai_mai_n164_));
  NO2        m142(.A(mai_mai_n155_), .B(mai_mai_n147_), .Y(mai_mai_n165_));
  NA3        m143(.A(mai_mai_n74_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n166_));
  NA2        m144(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n167_));
  NOi21      m145(.An(i_4_), .B(i_9_), .Y(mai_mai_n168_));
  NOi21      m146(.An(i_11_), .B(i_13_), .Y(mai_mai_n169_));
  NA2        m147(.A(mai_mai_n169_), .B(mai_mai_n168_), .Y(mai_mai_n170_));
  OR2        m148(.A(mai_mai_n170_), .B(mai_mai_n167_), .Y(mai_mai_n171_));
  NO2        m149(.A(i_4_), .B(i_5_), .Y(mai_mai_n172_));
  NAi21      m150(.An(i_12_), .B(i_11_), .Y(mai_mai_n173_));
  NO2        m151(.A(mai_mai_n173_), .B(i_13_), .Y(mai_mai_n174_));
  NA3        m152(.A(mai_mai_n174_), .B(mai_mai_n172_), .C(mai_mai_n84_), .Y(mai_mai_n175_));
  AOI210     m153(.A0(mai_mai_n175_), .A1(mai_mai_n171_), .B0(mai_mai_n166_), .Y(mai_mai_n176_));
  NO2        m154(.A(mai_mai_n74_), .B(mai_mai_n64_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n177_), .B(mai_mai_n47_), .Y(mai_mai_n178_));
  NA2        m156(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n179_));
  NA2        m157(.A(i_3_), .B(i_5_), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n181_));
  NO2        m159(.A(i_2_), .B(i_1_), .Y(mai_mai_n182_));
  NA2        m160(.A(mai_mai_n182_), .B(i_3_), .Y(mai_mai_n183_));
  NAi21      m161(.An(i_4_), .B(i_12_), .Y(mai_mai_n184_));
  NO4        m162(.A(mai_mai_n184_), .B(mai_mai_n183_), .C(i_11_), .D(mai_mai_n25_), .Y(mai_mai_n185_));
  NO2        m163(.A(mai_mai_n185_), .B(mai_mai_n176_), .Y(mai_mai_n186_));
  INV        m164(.A(i_8_), .Y(mai_mai_n187_));
  NO2        m165(.A(mai_mai_n187_), .B(i_7_), .Y(mai_mai_n188_));
  NA2        m166(.A(mai_mai_n188_), .B(i_6_), .Y(mai_mai_n189_));
  NO3        m167(.A(i_3_), .B(mai_mai_n87_), .C(mai_mai_n49_), .Y(mai_mai_n190_));
  NO3        m168(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n191_));
  NO2        m169(.A(i_3_), .B(i_8_), .Y(mai_mai_n192_));
  NO3        m170(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n193_));
  NA3        m171(.A(mai_mai_n193_), .B(mai_mai_n192_), .C(mai_mai_n40_), .Y(mai_mai_n194_));
  NO2        m172(.A(mai_mai_n107_), .B(mai_mai_n59_), .Y(mai_mai_n195_));
  INV        m173(.A(mai_mai_n195_), .Y(mai_mai_n196_));
  NO2        m174(.A(i_13_), .B(i_9_), .Y(mai_mai_n197_));
  NA3        m175(.A(mai_mai_n197_), .B(i_6_), .C(mai_mai_n187_), .Y(mai_mai_n198_));
  NAi21      m176(.An(i_12_), .B(i_3_), .Y(mai_mai_n199_));
  OR2        m177(.A(mai_mai_n199_), .B(mai_mai_n198_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n45_), .B(i_5_), .Y(mai_mai_n201_));
  NA3        m179(.A(i_1_), .B(mai_mai_n201_), .C(i_10_), .Y(mai_mai_n202_));
  OAI220     m180(.A0(mai_mai_n202_), .A1(mai_mai_n200_), .B0(mai_mai_n196_), .B1(mai_mai_n194_), .Y(mai_mai_n203_));
  NA2        m181(.A(mai_mai_n203_), .B(i_7_), .Y(mai_mai_n204_));
  OAI220     m182(.A0(mai_mai_n204_), .A1(i_4_), .B0(mai_mai_n189_), .B1(mai_mai_n186_), .Y(mai_mai_n205_));
  NAi21      m183(.An(i_12_), .B(i_7_), .Y(mai_mai_n206_));
  NA3        m184(.A(i_13_), .B(mai_mai_n187_), .C(i_10_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n207_), .B(mai_mai_n206_), .Y(mai_mai_n208_));
  NA2        m186(.A(i_0_), .B(i_5_), .Y(mai_mai_n209_));
  INV        m187(.A(mai_mai_n108_), .Y(mai_mai_n210_));
  OAI220     m188(.A0(mai_mai_n210_), .A1(mai_mai_n183_), .B0(mai_mai_n178_), .B1(mai_mai_n137_), .Y(mai_mai_n211_));
  NAi31      m189(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n212_));
  NO2        m190(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n213_));
  NO2        m191(.A(mai_mai_n74_), .B(mai_mai_n26_), .Y(mai_mai_n214_));
  NO2        m192(.A(mai_mai_n47_), .B(mai_mai_n64_), .Y(mai_mai_n215_));
  NA3        m193(.A(mai_mai_n215_), .B(mai_mai_n214_), .C(mai_mai_n213_), .Y(mai_mai_n216_));
  INV        m194(.A(i_13_), .Y(mai_mai_n217_));
  NO2        m195(.A(i_12_), .B(mai_mai_n217_), .Y(mai_mai_n218_));
  NA3        m196(.A(mai_mai_n218_), .B(mai_mai_n191_), .C(mai_mai_n190_), .Y(mai_mai_n219_));
  OAI210     m197(.A0(mai_mai_n216_), .A1(mai_mai_n212_), .B0(mai_mai_n219_), .Y(mai_mai_n220_));
  AOI220     m198(.A0(mai_mai_n220_), .A1(mai_mai_n146_), .B0(mai_mai_n211_), .B1(mai_mai_n208_), .Y(mai_mai_n221_));
  NO2        m199(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n222_));
  NO2        m200(.A(mai_mai_n180_), .B(i_4_), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n223_), .B(mai_mai_n222_), .Y(mai_mai_n224_));
  OR2        m202(.A(i_8_), .B(i_7_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n225_), .B(mai_mai_n87_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n54_), .B(i_1_), .Y(mai_mai_n227_));
  INV        m205(.A(i_12_), .Y(mai_mai_n228_));
  NO2        m206(.A(mai_mai_n45_), .B(mai_mai_n228_), .Y(mai_mai_n229_));
  NO3        m207(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n230_));
  NA2        m208(.A(i_2_), .B(i_1_), .Y(mai_mai_n231_));
  NO3        m209(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n232_));
  NAi21      m210(.An(i_4_), .B(i_3_), .Y(mai_mai_n233_));
  NO2        m211(.A(i_0_), .B(i_6_), .Y(mai_mai_n234_));
  NOi41      m212(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n235_), .B(mai_mai_n234_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n231_), .B(mai_mai_n180_), .Y(mai_mai_n237_));
  NAi21      m215(.An(mai_mai_n236_), .B(mai_mai_n237_), .Y(mai_mai_n238_));
  INV        m216(.A(mai_mai_n238_), .Y(mai_mai_n239_));
  NA2        m217(.A(mai_mai_n239_), .B(mai_mai_n40_), .Y(mai_mai_n240_));
  NO2        m218(.A(i_11_), .B(mai_mai_n217_), .Y(mai_mai_n241_));
  NOi21      m219(.An(i_1_), .B(i_6_), .Y(mai_mai_n242_));
  NAi21      m220(.An(i_3_), .B(i_7_), .Y(mai_mai_n243_));
  NA2        m221(.A(mai_mai_n228_), .B(i_9_), .Y(mai_mai_n244_));
  OR4        m222(.A(mai_mai_n244_), .B(mai_mai_n243_), .C(mai_mai_n242_), .D(mai_mai_n181_), .Y(mai_mai_n245_));
  NO2        m223(.A(mai_mai_n49_), .B(mai_mai_n25_), .Y(mai_mai_n246_));
  NA2        m224(.A(mai_mai_n74_), .B(i_5_), .Y(mai_mai_n247_));
  NA2        m225(.A(i_3_), .B(i_9_), .Y(mai_mai_n248_));
  NAi21      m226(.An(i_7_), .B(i_10_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n249_), .B(mai_mai_n248_), .Y(mai_mai_n250_));
  NA3        m228(.A(mai_mai_n250_), .B(mai_mai_n247_), .C(mai_mai_n65_), .Y(mai_mai_n251_));
  NA2        m229(.A(mai_mai_n251_), .B(mai_mai_n245_), .Y(mai_mai_n252_));
  NA3        m230(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n253_));
  INV        m231(.A(mai_mai_n147_), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n228_), .B(i_13_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n255_), .B(mai_mai_n76_), .Y(mai_mai_n256_));
  AOI220     m234(.A0(mai_mai_n256_), .A1(mai_mai_n254_), .B0(mai_mai_n252_), .B1(mai_mai_n241_), .Y(mai_mai_n257_));
  NA2        m235(.A(i_12_), .B(i_6_), .Y(mai_mai_n258_));
  OR2        m236(.A(i_13_), .B(i_9_), .Y(mai_mai_n259_));
  NO2        m237(.A(mai_mai_n233_), .B(i_2_), .Y(mai_mai_n260_));
  NA2        m238(.A(mai_mai_n241_), .B(i_9_), .Y(mai_mai_n261_));
  NO3        m239(.A(i_11_), .B(mai_mai_n217_), .C(mai_mai_n25_), .Y(mai_mai_n262_));
  NO2        m240(.A(mai_mai_n243_), .B(i_8_), .Y(mai_mai_n263_));
  NO2        m241(.A(i_6_), .B(mai_mai_n49_), .Y(mai_mai_n264_));
  NA3        m242(.A(mai_mai_n257_), .B(mai_mai_n240_), .C(mai_mai_n221_), .Y(mai_mai_n265_));
  NO3        m243(.A(i_12_), .B(mai_mai_n217_), .C(mai_mai_n37_), .Y(mai_mai_n266_));
  INV        m244(.A(mai_mai_n266_), .Y(mai_mai_n267_));
  NA2        m245(.A(i_8_), .B(mai_mai_n105_), .Y(mai_mai_n268_));
  NOi21      m246(.An(mai_mai_n162_), .B(mai_mai_n87_), .Y(mai_mai_n269_));
  NO3        m247(.A(i_0_), .B(mai_mai_n47_), .C(i_1_), .Y(mai_mai_n270_));
  AOI220     m248(.A0(mai_mai_n270_), .A1(mai_mai_n190_), .B0(mai_mai_n269_), .B1(mai_mai_n227_), .Y(mai_mai_n271_));
  NO2        m249(.A(mai_mai_n271_), .B(mai_mai_n268_), .Y(mai_mai_n272_));
  NO3        m250(.A(i_0_), .B(i_2_), .C(mai_mai_n64_), .Y(mai_mai_n273_));
  NO2        m251(.A(mai_mai_n231_), .B(i_0_), .Y(mai_mai_n274_));
  AOI220     m252(.A0(mai_mai_n274_), .A1(mai_mai_n188_), .B0(mai_mai_n273_), .B1(mai_mai_n146_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n264_), .B(mai_mai_n26_), .Y(mai_mai_n276_));
  NO2        m254(.A(mai_mai_n276_), .B(mai_mai_n275_), .Y(mai_mai_n277_));
  NA2        m255(.A(i_0_), .B(i_1_), .Y(mai_mai_n278_));
  NO2        m256(.A(mai_mai_n278_), .B(i_2_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n280_));
  NA3        m258(.A(mai_mai_n280_), .B(mai_mai_n279_), .C(mai_mai_n162_), .Y(mai_mai_n281_));
  OAI210     m259(.A0(mai_mai_n164_), .A1(mai_mai_n147_), .B0(mai_mai_n281_), .Y(mai_mai_n282_));
  NO3        m260(.A(mai_mai_n282_), .B(mai_mai_n277_), .C(mai_mai_n272_), .Y(mai_mai_n283_));
  NO2        m261(.A(i_3_), .B(i_10_), .Y(mai_mai_n284_));
  NA3        m262(.A(mai_mai_n284_), .B(mai_mai_n40_), .C(mai_mai_n45_), .Y(mai_mai_n285_));
  NO2        m263(.A(i_2_), .B(mai_mai_n105_), .Y(mai_mai_n286_));
  NOi21      m264(.An(mai_mai_n209_), .B(mai_mai_n107_), .Y(mai_mai_n287_));
  NA3        m265(.A(mai_mai_n287_), .B(i_1_), .C(mai_mai_n286_), .Y(mai_mai_n288_));
  AN2        m266(.A(i_3_), .B(i_10_), .Y(mai_mai_n289_));
  NA4        m267(.A(mai_mai_n289_), .B(mai_mai_n191_), .C(mai_mai_n174_), .D(mai_mai_n172_), .Y(mai_mai_n290_));
  NO2        m268(.A(i_5_), .B(mai_mai_n37_), .Y(mai_mai_n291_));
  NO2        m269(.A(mai_mai_n47_), .B(mai_mai_n26_), .Y(mai_mai_n292_));
  OR2        m270(.A(mai_mai_n288_), .B(mai_mai_n285_), .Y(mai_mai_n293_));
  OAI220     m271(.A0(mai_mai_n293_), .A1(i_6_), .B0(mai_mai_n283_), .B1(mai_mai_n267_), .Y(mai_mai_n294_));
  NO4        m272(.A(mai_mai_n294_), .B(mai_mai_n265_), .C(mai_mai_n205_), .D(mai_mai_n165_), .Y(mai_mai_n295_));
  NO3        m273(.A(mai_mai_n45_), .B(i_13_), .C(i_9_), .Y(mai_mai_n296_));
  NO2        m274(.A(mai_mai_n60_), .B(mai_mai_n87_), .Y(mai_mai_n297_));
  NA2        m275(.A(mai_mai_n274_), .B(mai_mai_n297_), .Y(mai_mai_n298_));
  NO3        m276(.A(i_6_), .B(mai_mai_n187_), .C(i_7_), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n298_), .B(mai_mai_n167_), .Y(mai_mai_n300_));
  NO2        m278(.A(i_2_), .B(i_3_), .Y(mai_mai_n301_));
  OR2        m279(.A(i_0_), .B(i_5_), .Y(mai_mai_n302_));
  NA2        m280(.A(mai_mai_n209_), .B(mai_mai_n302_), .Y(mai_mai_n303_));
  NA4        m281(.A(mai_mai_n303_), .B(mai_mai_n226_), .C(mai_mai_n301_), .D(i_1_), .Y(mai_mai_n304_));
  NA3        m282(.A(mai_mai_n274_), .B(mai_mai_n269_), .C(mai_mai_n116_), .Y(mai_mai_n305_));
  NAi21      m283(.An(i_8_), .B(i_7_), .Y(mai_mai_n306_));
  NO2        m284(.A(mai_mai_n306_), .B(i_6_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n158_), .B(mai_mai_n47_), .Y(mai_mai_n308_));
  NA3        m286(.A(mai_mai_n308_), .B(mai_mai_n307_), .C(mai_mai_n162_), .Y(mai_mai_n309_));
  NA3        m287(.A(mai_mai_n309_), .B(mai_mai_n305_), .C(mai_mai_n304_), .Y(mai_mai_n310_));
  OAI210     m288(.A0(mai_mai_n310_), .A1(mai_mai_n300_), .B0(i_4_), .Y(mai_mai_n311_));
  NO2        m289(.A(i_12_), .B(i_10_), .Y(mai_mai_n312_));
  NOi21      m290(.An(i_5_), .B(i_0_), .Y(mai_mai_n313_));
  NA4        m291(.A(mai_mai_n85_), .B(mai_mai_n36_), .C(mai_mai_n87_), .D(i_8_), .Y(mai_mai_n314_));
  NO2        m292(.A(i_6_), .B(i_8_), .Y(mai_mai_n315_));
  NOi21      m293(.An(i_0_), .B(i_2_), .Y(mai_mai_n316_));
  AN2        m294(.A(mai_mai_n316_), .B(mai_mai_n315_), .Y(mai_mai_n317_));
  NO2        m295(.A(i_1_), .B(i_7_), .Y(mai_mai_n318_));
  AO220      m296(.A0(mai_mai_n318_), .A1(mai_mai_n317_), .B0(mai_mai_n307_), .B1(mai_mai_n227_), .Y(mai_mai_n319_));
  NA2        m297(.A(mai_mai_n319_), .B(mai_mai_n42_), .Y(mai_mai_n320_));
  NA2        m298(.A(mai_mai_n320_), .B(mai_mai_n311_), .Y(mai_mai_n321_));
  NA3        m299(.A(mai_mai_n242_), .B(mai_mai_n286_), .C(mai_mai_n187_), .Y(mai_mai_n322_));
  INV        m300(.A(mai_mai_n85_), .Y(mai_mai_n323_));
  NO2        m301(.A(mai_mai_n278_), .B(mai_mai_n82_), .Y(mai_mai_n324_));
  NA2        m302(.A(mai_mai_n324_), .B(mai_mai_n136_), .Y(mai_mai_n325_));
  NO2        m303(.A(mai_mai_n96_), .B(mai_mai_n187_), .Y(mai_mai_n326_));
  NA3        m304(.A(mai_mai_n287_), .B(mai_mai_n326_), .C(mai_mai_n64_), .Y(mai_mai_n327_));
  AOI210     m305(.A0(mai_mai_n327_), .A1(mai_mai_n325_), .B0(mai_mai_n323_), .Y(mai_mai_n328_));
  NO2        m306(.A(mai_mai_n187_), .B(i_9_), .Y(mai_mai_n329_));
  NA2        m307(.A(mai_mai_n329_), .B(mai_mai_n195_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n328_), .B(mai_mai_n277_), .Y(mai_mai_n331_));
  AOI210     m309(.A0(mai_mai_n331_), .A1(mai_mai_n322_), .B0(mai_mai_n161_), .Y(mai_mai_n332_));
  AOI210     m310(.A0(mai_mai_n321_), .A1(mai_mai_n296_), .B0(mai_mai_n332_), .Y(mai_mai_n333_));
  NOi32      m311(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n334_));
  INV        m312(.A(mai_mai_n334_), .Y(mai_mai_n335_));
  NAi21      m313(.An(i_1_), .B(i_5_), .Y(mai_mai_n336_));
  INV        m314(.A(mai_mai_n236_), .Y(mai_mai_n337_));
  NAi41      m315(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n338_));
  OAI220     m316(.A0(mai_mai_n338_), .A1(mai_mai_n336_), .B0(mai_mai_n212_), .B1(mai_mai_n159_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n338_), .A1(mai_mai_n159_), .B0(mai_mai_n158_), .Y(mai_mai_n340_));
  NOi32      m318(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n341_));
  NAi21      m319(.An(i_6_), .B(i_1_), .Y(mai_mai_n342_));
  NA3        m320(.A(mai_mai_n342_), .B(mai_mai_n341_), .C(mai_mai_n47_), .Y(mai_mai_n343_));
  NO2        m321(.A(mai_mai_n343_), .B(i_0_), .Y(mai_mai_n344_));
  OR3        m322(.A(mai_mai_n344_), .B(mai_mai_n340_), .C(mai_mai_n339_), .Y(mai_mai_n345_));
  NO2        m323(.A(i_1_), .B(mai_mai_n105_), .Y(mai_mai_n346_));
  NAi21      m324(.An(i_3_), .B(i_4_), .Y(mai_mai_n347_));
  NO2        m325(.A(mai_mai_n347_), .B(i_9_), .Y(mai_mai_n348_));
  AN2        m326(.A(i_6_), .B(i_7_), .Y(mai_mai_n349_));
  OAI210     m327(.A0(mai_mai_n349_), .A1(mai_mai_n346_), .B0(mai_mai_n348_), .Y(mai_mai_n350_));
  NA2        m328(.A(i_2_), .B(i_7_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n347_), .B(i_10_), .Y(mai_mai_n352_));
  NA3        m330(.A(mai_mai_n352_), .B(mai_mai_n351_), .C(mai_mai_n234_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n353_), .A1(mai_mai_n350_), .B0(mai_mai_n181_), .Y(mai_mai_n354_));
  AOI210     m332(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n355_));
  OAI210     m333(.A0(mai_mai_n355_), .A1(mai_mai_n182_), .B0(mai_mai_n352_), .Y(mai_mai_n356_));
  AOI220     m334(.A0(mai_mai_n352_), .A1(mai_mai_n318_), .B0(mai_mai_n230_), .B1(mai_mai_n182_), .Y(mai_mai_n357_));
  AOI210     m335(.A0(mai_mai_n357_), .A1(mai_mai_n356_), .B0(i_5_), .Y(mai_mai_n358_));
  NO4        m336(.A(mai_mai_n358_), .B(mai_mai_n354_), .C(mai_mai_n345_), .D(mai_mai_n337_), .Y(mai_mai_n359_));
  NO2        m337(.A(mai_mai_n359_), .B(mai_mai_n335_), .Y(mai_mai_n360_));
  NO2        m338(.A(mai_mai_n60_), .B(mai_mai_n25_), .Y(mai_mai_n361_));
  AN2        m339(.A(i_12_), .B(i_5_), .Y(mai_mai_n362_));
  NO2        m340(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n363_));
  NA2        m341(.A(mai_mai_n363_), .B(mai_mai_n362_), .Y(mai_mai_n364_));
  NO2        m342(.A(i_11_), .B(i_6_), .Y(mai_mai_n365_));
  NA3        m343(.A(mai_mai_n365_), .B(mai_mai_n308_), .C(mai_mai_n217_), .Y(mai_mai_n366_));
  NO2        m344(.A(mai_mai_n366_), .B(mai_mai_n364_), .Y(mai_mai_n367_));
  NO2        m345(.A(mai_mai_n233_), .B(i_5_), .Y(mai_mai_n368_));
  NO2        m346(.A(i_5_), .B(i_10_), .Y(mai_mai_n369_));
  AOI220     m347(.A0(mai_mai_n369_), .A1(mai_mai_n260_), .B0(mai_mai_n368_), .B1(mai_mai_n191_), .Y(mai_mai_n370_));
  NA2        m348(.A(mai_mai_n148_), .B(mai_mai_n46_), .Y(mai_mai_n371_));
  NO2        m349(.A(mai_mai_n371_), .B(mai_mai_n370_), .Y(mai_mai_n372_));
  OAI210     m350(.A0(mai_mai_n372_), .A1(mai_mai_n367_), .B0(mai_mai_n361_), .Y(mai_mai_n373_));
  NO2        m351(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n374_));
  NO2        m352(.A(mai_mai_n154_), .B(mai_mai_n87_), .Y(mai_mai_n375_));
  OAI210     m353(.A0(mai_mai_n375_), .A1(mai_mai_n367_), .B0(mai_mai_n374_), .Y(mai_mai_n376_));
  NO3        m354(.A(mai_mai_n87_), .B(mai_mai_n49_), .C(i_9_), .Y(mai_mai_n377_));
  NO2        m355(.A(i_11_), .B(i_12_), .Y(mai_mai_n378_));
  NA3        m356(.A(mai_mai_n116_), .B(mai_mai_n42_), .C(i_11_), .Y(mai_mai_n379_));
  NO2        m357(.A(mai_mai_n379_), .B(mai_mai_n212_), .Y(mai_mai_n380_));
  NAi21      m358(.An(i_13_), .B(i_0_), .Y(mai_mai_n381_));
  NO2        m359(.A(mai_mai_n381_), .B(mai_mai_n231_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n380_), .B(mai_mai_n382_), .Y(mai_mai_n383_));
  NA3        m361(.A(mai_mai_n383_), .B(mai_mai_n376_), .C(mai_mai_n373_), .Y(mai_mai_n384_));
  NA2        m362(.A(mai_mai_n45_), .B(mai_mai_n217_), .Y(mai_mai_n385_));
  NO3        m363(.A(i_1_), .B(i_12_), .C(mai_mai_n87_), .Y(mai_mai_n386_));
  NO2        m364(.A(i_0_), .B(i_11_), .Y(mai_mai_n387_));
  INV        m365(.A(i_5_), .Y(mai_mai_n388_));
  AN2        m366(.A(i_1_), .B(i_6_), .Y(mai_mai_n389_));
  NOi21      m367(.An(i_2_), .B(i_12_), .Y(mai_mai_n390_));
  NA2        m368(.A(mai_mai_n390_), .B(mai_mai_n389_), .Y(mai_mai_n391_));
  NO2        m369(.A(mai_mai_n391_), .B(mai_mai_n388_), .Y(mai_mai_n392_));
  NA2        m370(.A(mai_mai_n146_), .B(i_9_), .Y(mai_mai_n393_));
  NO2        m371(.A(mai_mai_n393_), .B(i_4_), .Y(mai_mai_n394_));
  NA2        m372(.A(mai_mai_n392_), .B(mai_mai_n394_), .Y(mai_mai_n395_));
  NAi21      m373(.An(i_9_), .B(i_4_), .Y(mai_mai_n396_));
  OR2        m374(.A(i_13_), .B(i_10_), .Y(mai_mai_n397_));
  NO3        m375(.A(mai_mai_n397_), .B(mai_mai_n121_), .C(mai_mai_n396_), .Y(mai_mai_n398_));
  NO2        m376(.A(mai_mai_n170_), .B(mai_mai_n127_), .Y(mai_mai_n399_));
  NO2        m377(.A(mai_mai_n105_), .B(mai_mai_n25_), .Y(mai_mai_n400_));
  NO2        m378(.A(mai_mai_n395_), .B(mai_mai_n26_), .Y(mai_mai_n401_));
  NA2        m379(.A(mai_mai_n305_), .B(mai_mai_n304_), .Y(mai_mai_n402_));
  AOI220     m380(.A0(mai_mai_n280_), .A1(mai_mai_n270_), .B0(mai_mai_n274_), .B1(mai_mai_n297_), .Y(mai_mai_n403_));
  NO2        m381(.A(mai_mai_n403_), .B(mai_mai_n167_), .Y(mai_mai_n404_));
  NO2        m382(.A(mai_mai_n180_), .B(mai_mai_n87_), .Y(mai_mai_n405_));
  NO2        m383(.A(mai_mai_n404_), .B(mai_mai_n402_), .Y(mai_mai_n406_));
  NA2        m384(.A(mai_mai_n190_), .B(mai_mai_n100_), .Y(mai_mai_n407_));
  NA3        m385(.A(mai_mai_n308_), .B(mai_mai_n162_), .C(mai_mai_n87_), .Y(mai_mai_n408_));
  AOI210     m386(.A0(mai_mai_n408_), .A1(mai_mai_n407_), .B0(mai_mai_n306_), .Y(mai_mai_n409_));
  NO2        m387(.A(i_3_), .B(mai_mai_n49_), .Y(mai_mai_n410_));
  NA3        m388(.A(mai_mai_n318_), .B(mai_mai_n317_), .C(mai_mai_n410_), .Y(mai_mai_n411_));
  NA2        m389(.A(mai_mai_n299_), .B(mai_mai_n303_), .Y(mai_mai_n412_));
  OAI210     m390(.A0(mai_mai_n412_), .A1(mai_mai_n183_), .B0(mai_mai_n411_), .Y(mai_mai_n413_));
  NO2        m391(.A(mai_mai_n413_), .B(mai_mai_n409_), .Y(mai_mai_n414_));
  AOI210     m392(.A0(mai_mai_n414_), .A1(mai_mai_n406_), .B0(mai_mai_n261_), .Y(mai_mai_n415_));
  NO4        m393(.A(mai_mai_n415_), .B(mai_mai_n401_), .C(mai_mai_n384_), .D(mai_mai_n360_), .Y(mai_mai_n416_));
  NO2        m394(.A(mai_mai_n64_), .B(i_4_), .Y(mai_mai_n417_));
  NO2        m395(.A(mai_mai_n74_), .B(i_13_), .Y(mai_mai_n418_));
  NA3        m396(.A(mai_mai_n418_), .B(mai_mai_n417_), .C(i_2_), .Y(mai_mai_n419_));
  NO2        m397(.A(i_10_), .B(i_9_), .Y(mai_mai_n420_));
  NAi21      m398(.An(i_12_), .B(i_8_), .Y(mai_mai_n421_));
  NO2        m399(.A(mai_mai_n421_), .B(i_3_), .Y(mai_mai_n422_));
  NA2        m400(.A(mai_mai_n422_), .B(mai_mai_n420_), .Y(mai_mai_n423_));
  NO2        m401(.A(mai_mai_n47_), .B(i_4_), .Y(mai_mai_n424_));
  NA2        m402(.A(mai_mai_n424_), .B(mai_mai_n108_), .Y(mai_mai_n425_));
  OAI220     m403(.A0(mai_mai_n425_), .A1(mai_mai_n194_), .B0(mai_mai_n423_), .B1(mai_mai_n419_), .Y(mai_mai_n426_));
  NA2        m404(.A(mai_mai_n292_), .B(i_0_), .Y(mai_mai_n427_));
  NO3        m405(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n428_));
  NA2        m406(.A(mai_mai_n258_), .B(mai_mai_n101_), .Y(mai_mai_n429_));
  NA2        m407(.A(mai_mai_n429_), .B(mai_mai_n428_), .Y(mai_mai_n430_));
  NA2        m408(.A(i_8_), .B(i_9_), .Y(mai_mai_n431_));
  AOI210     m409(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n432_));
  OR2        m410(.A(mai_mai_n432_), .B(mai_mai_n431_), .Y(mai_mai_n433_));
  NA2        m411(.A(mai_mai_n266_), .B(mai_mai_n195_), .Y(mai_mai_n434_));
  OAI220     m412(.A0(mai_mai_n434_), .A1(mai_mai_n433_), .B0(mai_mai_n430_), .B1(mai_mai_n427_), .Y(mai_mai_n435_));
  NA2        m413(.A(mai_mai_n241_), .B(mai_mai_n291_), .Y(mai_mai_n436_));
  NO3        m414(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n437_));
  INV        m415(.A(mai_mai_n437_), .Y(mai_mai_n438_));
  NA3        m416(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n439_));
  NA4        m417(.A(mai_mai_n149_), .B(mai_mai_n119_), .C(mai_mai_n81_), .D(mai_mai_n23_), .Y(mai_mai_n440_));
  OAI220     m418(.A0(mai_mai_n440_), .A1(mai_mai_n439_), .B0(mai_mai_n438_), .B1(mai_mai_n436_), .Y(mai_mai_n441_));
  NO3        m419(.A(mai_mai_n441_), .B(mai_mai_n435_), .C(mai_mai_n426_), .Y(mai_mai_n442_));
  NA2        m420(.A(mai_mai_n279_), .B(mai_mai_n112_), .Y(mai_mai_n443_));
  OR2        m421(.A(mai_mai_n443_), .B(mai_mai_n198_), .Y(mai_mai_n444_));
  OR2        m422(.A(mai_mai_n330_), .B(mai_mai_n105_), .Y(mai_mai_n445_));
  OA220      m423(.A0(mai_mai_n445_), .A1(mai_mai_n161_), .B0(mai_mai_n444_), .B1(mai_mai_n224_), .Y(mai_mai_n446_));
  NA2        m424(.A(mai_mai_n100_), .B(i_13_), .Y(mai_mai_n447_));
  NA2        m425(.A(mai_mai_n405_), .B(mai_mai_n361_), .Y(mai_mai_n448_));
  NO2        m426(.A(i_2_), .B(i_13_), .Y(mai_mai_n449_));
  NO2        m427(.A(mai_mai_n448_), .B(mai_mai_n447_), .Y(mai_mai_n450_));
  NO3        m428(.A(i_4_), .B(mai_mai_n49_), .C(i_8_), .Y(mai_mai_n451_));
  NO2        m429(.A(i_6_), .B(i_7_), .Y(mai_mai_n452_));
  NA2        m430(.A(mai_mai_n452_), .B(mai_mai_n451_), .Y(mai_mai_n453_));
  NO2        m431(.A(i_11_), .B(i_1_), .Y(mai_mai_n454_));
  OR2        m432(.A(i_11_), .B(i_8_), .Y(mai_mai_n455_));
  NOi21      m433(.An(i_2_), .B(i_7_), .Y(mai_mai_n456_));
  NAi31      m434(.An(mai_mai_n455_), .B(mai_mai_n456_), .C(i_0_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n397_), .B(i_6_), .Y(mai_mai_n458_));
  NA3        m436(.A(mai_mai_n458_), .B(mai_mai_n417_), .C(mai_mai_n76_), .Y(mai_mai_n459_));
  NO2        m437(.A(mai_mai_n459_), .B(mai_mai_n457_), .Y(mai_mai_n460_));
  NO2        m438(.A(i_3_), .B(mai_mai_n187_), .Y(mai_mai_n461_));
  NO2        m439(.A(i_6_), .B(i_10_), .Y(mai_mai_n462_));
  NA3        m440(.A(mai_mai_n235_), .B(mai_mai_n169_), .C(mai_mai_n136_), .Y(mai_mai_n463_));
  NA2        m441(.A(mai_mai_n47_), .B(mai_mai_n45_), .Y(mai_mai_n464_));
  NO2        m442(.A(mai_mai_n158_), .B(i_3_), .Y(mai_mai_n465_));
  NAi31      m443(.An(mai_mai_n464_), .B(mai_mai_n465_), .C(mai_mai_n218_), .Y(mai_mai_n466_));
  NA3        m444(.A(mai_mai_n374_), .B(mai_mai_n177_), .C(mai_mai_n153_), .Y(mai_mai_n467_));
  NA3        m445(.A(mai_mai_n467_), .B(mai_mai_n466_), .C(mai_mai_n463_), .Y(mai_mai_n468_));
  NO3        m446(.A(mai_mai_n468_), .B(mai_mai_n460_), .C(mai_mai_n450_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n437_), .B(mai_mai_n369_), .Y(mai_mai_n470_));
  NO2        m448(.A(mai_mai_n470_), .B(mai_mai_n216_), .Y(mai_mai_n471_));
  NAi21      m449(.An(mai_mai_n207_), .B(mai_mai_n378_), .Y(mai_mai_n472_));
  NA2        m450(.A(mai_mai_n318_), .B(mai_mai_n209_), .Y(mai_mai_n473_));
  NO2        m451(.A(mai_mai_n473_), .B(mai_mai_n472_), .Y(mai_mai_n474_));
  NA2        m452(.A(mai_mai_n27_), .B(i_10_), .Y(mai_mai_n475_));
  NO2        m453(.A(mai_mai_n475_), .B(mai_mai_n447_), .Y(mai_mai_n476_));
  NA4        m454(.A(mai_mai_n289_), .B(mai_mai_n215_), .C(mai_mai_n74_), .D(mai_mai_n228_), .Y(mai_mai_n477_));
  NO2        m455(.A(mai_mai_n477_), .B(mai_mai_n453_), .Y(mai_mai_n478_));
  NO4        m456(.A(mai_mai_n478_), .B(mai_mai_n476_), .C(mai_mai_n474_), .D(mai_mai_n471_), .Y(mai_mai_n479_));
  NA4        m457(.A(mai_mai_n479_), .B(mai_mai_n469_), .C(mai_mai_n446_), .D(mai_mai_n442_), .Y(mai_mai_n480_));
  NA3        m458(.A(mai_mai_n289_), .B(mai_mai_n174_), .C(mai_mai_n172_), .Y(mai_mai_n481_));
  OAI210     m459(.A0(mai_mai_n285_), .A1(mai_mai_n179_), .B0(mai_mai_n481_), .Y(mai_mai_n482_));
  AN2        m460(.A(mai_mai_n270_), .B(mai_mai_n226_), .Y(mai_mai_n483_));
  NA2        m461(.A(mai_mai_n483_), .B(mai_mai_n482_), .Y(mai_mai_n484_));
  NA2        m462(.A(mai_mai_n126_), .B(mai_mai_n115_), .Y(mai_mai_n485_));
  AN2        m463(.A(mai_mai_n485_), .B(mai_mai_n428_), .Y(mai_mai_n486_));
  NA2        m464(.A(mai_mai_n296_), .B(mai_mai_n163_), .Y(mai_mai_n487_));
  OAI210     m465(.A0(mai_mai_n487_), .A1(mai_mai_n224_), .B0(mai_mai_n290_), .Y(mai_mai_n488_));
  AOI220     m466(.A0(mai_mai_n488_), .A1(mai_mai_n307_), .B0(mai_mai_n486_), .B1(mai_mai_n292_), .Y(mai_mai_n489_));
  NA2        m467(.A(mai_mai_n334_), .B(mai_mai_n74_), .Y(mai_mai_n490_));
  NA2        m468(.A(mai_mai_n349_), .B(mai_mai_n341_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n492_));
  NAi41      m470(.An(mai_mai_n490_), .B(mai_mai_n462_), .C(mai_mai_n492_), .D(mai_mai_n47_), .Y(mai_mai_n493_));
  AOI210     m471(.A0(mai_mai_n39_), .A1(i_13_), .B0(mai_mai_n398_), .Y(mai_mai_n494_));
  NA2        m472(.A(mai_mai_n494_), .B(mai_mai_n493_), .Y(mai_mai_n495_));
  NA2        m473(.A(mai_mai_n247_), .B(mai_mai_n65_), .Y(mai_mai_n496_));
  OAI210     m474(.A0(i_8_), .A1(mai_mai_n496_), .B0(mai_mai_n138_), .Y(mai_mai_n497_));
  NA2        m475(.A(mai_mai_n497_), .B(mai_mai_n399_), .Y(mai_mai_n498_));
  NA4        m476(.A(mai_mai_n498_), .B(mai_mai_n494_), .C(mai_mai_n489_), .D(mai_mai_n484_), .Y(mai_mai_n499_));
  NA2        m477(.A(mai_mai_n368_), .B(mai_mai_n279_), .Y(mai_mai_n500_));
  OAI210     m478(.A0(mai_mai_n364_), .A1(mai_mai_n166_), .B0(mai_mai_n500_), .Y(mai_mai_n501_));
  NO2        m479(.A(i_12_), .B(mai_mai_n187_), .Y(mai_mai_n502_));
  NA2        m480(.A(mai_mai_n462_), .B(mai_mai_n27_), .Y(mai_mai_n503_));
  NO3        m481(.A(mai_mai_n503_), .B(i_12_), .C(mai_mai_n443_), .Y(mai_mai_n504_));
  NOi31      m482(.An(mai_mai_n299_), .B(mai_mai_n397_), .C(mai_mai_n38_), .Y(mai_mai_n505_));
  OAI210     m483(.A0(mai_mai_n505_), .A1(mai_mai_n504_), .B0(mai_mai_n501_), .Y(mai_mai_n506_));
  NO2        m484(.A(i_8_), .B(i_7_), .Y(mai_mai_n507_));
  NA2        m485(.A(mai_mai_n45_), .B(i_10_), .Y(mai_mai_n508_));
  NO2        m486(.A(mai_mai_n508_), .B(i_6_), .Y(mai_mai_n509_));
  NOi31      m487(.An(mai_mai_n274_), .B(mai_mai_n285_), .C(mai_mai_n179_), .Y(mai_mai_n510_));
  NA3        m488(.A(mai_mai_n289_), .B(mai_mai_n172_), .C(mai_mai_n100_), .Y(mai_mai_n511_));
  NO2        m489(.A(mai_mai_n213_), .B(mai_mai_n45_), .Y(mai_mai_n512_));
  NO2        m490(.A(mai_mai_n158_), .B(i_5_), .Y(mai_mai_n513_));
  NA3        m491(.A(mai_mai_n513_), .B(mai_mai_n385_), .C(mai_mai_n301_), .Y(mai_mai_n514_));
  OAI210     m492(.A0(mai_mai_n514_), .A1(mai_mai_n512_), .B0(mai_mai_n511_), .Y(mai_mai_n515_));
  OAI210     m493(.A0(mai_mai_n515_), .A1(mai_mai_n510_), .B0(mai_mai_n437_), .Y(mai_mai_n516_));
  NA2        m494(.A(mai_mai_n516_), .B(mai_mai_n506_), .Y(mai_mai_n517_));
  NA3        m495(.A(mai_mai_n209_), .B(mai_mai_n72_), .C(mai_mai_n45_), .Y(mai_mai_n518_));
  NA2        m496(.A(mai_mai_n266_), .B(mai_mai_n85_), .Y(mai_mai_n519_));
  AOI210     m497(.A0(mai_mai_n518_), .A1(mai_mai_n325_), .B0(mai_mai_n519_), .Y(mai_mai_n520_));
  NA2        m498(.A(mai_mai_n280_), .B(mai_mai_n270_), .Y(mai_mai_n521_));
  NO2        m499(.A(mai_mai_n521_), .B(mai_mai_n171_), .Y(mai_mai_n522_));
  NA2        m500(.A(mai_mai_n215_), .B(mai_mai_n214_), .Y(mai_mai_n523_));
  NA2        m501(.A(mai_mai_n420_), .B(mai_mai_n213_), .Y(mai_mai_n524_));
  NO2        m502(.A(mai_mai_n523_), .B(mai_mai_n524_), .Y(mai_mai_n525_));
  AOI210     m503(.A0(mai_mai_n342_), .A1(mai_mai_n47_), .B0(mai_mai_n346_), .Y(mai_mai_n526_));
  NA2        m504(.A(i_0_), .B(mai_mai_n49_), .Y(mai_mai_n527_));
  NA3        m505(.A(mai_mai_n502_), .B(mai_mai_n262_), .C(mai_mai_n527_), .Y(mai_mai_n528_));
  NO2        m506(.A(mai_mai_n526_), .B(mai_mai_n528_), .Y(mai_mai_n529_));
  NO4        m507(.A(mai_mai_n529_), .B(mai_mai_n525_), .C(mai_mai_n522_), .D(mai_mai_n520_), .Y(mai_mai_n530_));
  NO4        m508(.A(mai_mai_n242_), .B(mai_mai_n43_), .C(i_2_), .D(mai_mai_n49_), .Y(mai_mai_n531_));
  NO3        m509(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n532_));
  NO2        m510(.A(mai_mai_n225_), .B(mai_mai_n36_), .Y(mai_mai_n533_));
  AN2        m511(.A(mai_mai_n533_), .B(mai_mai_n532_), .Y(mai_mai_n534_));
  OA210      m512(.A0(mai_mai_n534_), .A1(mai_mai_n531_), .B0(mai_mai_n334_), .Y(mai_mai_n535_));
  NO2        m513(.A(mai_mai_n397_), .B(i_1_), .Y(mai_mai_n536_));
  NOi31      m514(.An(mai_mai_n536_), .B(mai_mai_n429_), .C(mai_mai_n74_), .Y(mai_mai_n537_));
  AN4        m515(.A(mai_mai_n537_), .B(mai_mai_n394_), .C(i_3_), .D(i_2_), .Y(mai_mai_n538_));
  NO2        m516(.A(mai_mai_n403_), .B(mai_mai_n175_), .Y(mai_mai_n539_));
  NO3        m517(.A(mai_mai_n539_), .B(mai_mai_n538_), .C(mai_mai_n535_), .Y(mai_mai_n540_));
  NOi21      m518(.An(i_10_), .B(i_6_), .Y(mai_mai_n541_));
  NO2        m519(.A(mai_mai_n87_), .B(mai_mai_n25_), .Y(mai_mai_n542_));
  AOI220     m520(.A0(mai_mai_n266_), .A1(mai_mai_n542_), .B0(mai_mai_n262_), .B1(mai_mai_n541_), .Y(mai_mai_n543_));
  NO2        m521(.A(mai_mai_n543_), .B(mai_mai_n427_), .Y(mai_mai_n544_));
  NO2        m522(.A(mai_mai_n118_), .B(mai_mai_n23_), .Y(mai_mai_n545_));
  NO2        m523(.A(mai_mai_n191_), .B(mai_mai_n37_), .Y(mai_mai_n546_));
  NOi31      m524(.An(mai_mai_n150_), .B(mai_mai_n546_), .C(mai_mai_n314_), .Y(mai_mai_n547_));
  NO2        m525(.A(mai_mai_n547_), .B(mai_mai_n544_), .Y(mai_mai_n548_));
  NO2        m526(.A(mai_mai_n490_), .B(mai_mai_n357_), .Y(mai_mai_n549_));
  INV        m527(.A(mai_mai_n301_), .Y(mai_mai_n550_));
  NO2        m528(.A(i_12_), .B(mai_mai_n87_), .Y(mai_mai_n551_));
  OR2        m529(.A(i_2_), .B(i_5_), .Y(mai_mai_n552_));
  OR2        m530(.A(mai_mai_n552_), .B(mai_mai_n389_), .Y(mai_mai_n553_));
  NA2        m531(.A(mai_mai_n351_), .B(mai_mai_n234_), .Y(mai_mai_n554_));
  AOI210     m532(.A0(mai_mai_n554_), .A1(mai_mai_n553_), .B0(mai_mai_n472_), .Y(mai_mai_n555_));
  NO2        m533(.A(mai_mai_n555_), .B(mai_mai_n549_), .Y(mai_mai_n556_));
  NA4        m534(.A(mai_mai_n556_), .B(mai_mai_n548_), .C(mai_mai_n540_), .D(mai_mai_n530_), .Y(mai_mai_n557_));
  NO4        m535(.A(mai_mai_n557_), .B(mai_mai_n517_), .C(mai_mai_n499_), .D(mai_mai_n480_), .Y(mai_mai_n558_));
  NA4        m536(.A(mai_mai_n558_), .B(mai_mai_n416_), .C(mai_mai_n333_), .D(mai_mai_n295_), .Y(mai7));
  NO2        m537(.A(mai_mai_n96_), .B(mai_mai_n55_), .Y(mai_mai_n560_));
  NA2        m538(.A(i_11_), .B(mai_mai_n187_), .Y(mai_mai_n561_));
  NA3        m539(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n562_));
  NO2        m540(.A(mai_mai_n228_), .B(i_4_), .Y(mai_mai_n563_));
  NA2        m541(.A(mai_mai_n563_), .B(i_8_), .Y(mai_mai_n564_));
  NO2        m542(.A(mai_mai_n109_), .B(mai_mai_n562_), .Y(mai_mai_n565_));
  NA2        m543(.A(i_2_), .B(mai_mai_n87_), .Y(mai_mai_n566_));
  OAI210     m544(.A0(mai_mai_n90_), .A1(mai_mai_n192_), .B0(mai_mai_n193_), .Y(mai_mai_n567_));
  NO2        m545(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n568_));
  NA2        m546(.A(i_4_), .B(i_8_), .Y(mai_mai_n569_));
  AOI210     m547(.A0(mai_mai_n569_), .A1(mai_mai_n289_), .B0(mai_mai_n568_), .Y(mai_mai_n570_));
  OAI220     m548(.A0(mai_mai_n570_), .A1(mai_mai_n566_), .B0(mai_mai_n567_), .B1(i_13_), .Y(mai_mai_n571_));
  NO3        m549(.A(mai_mai_n571_), .B(mai_mai_n565_), .C(mai_mai_n560_), .Y(mai_mai_n572_));
  AOI210     m550(.A0(mai_mai_n132_), .A1(mai_mai_n63_), .B0(i_10_), .Y(mai_mai_n573_));
  AOI210     m551(.A0(mai_mai_n573_), .A1(mai_mai_n228_), .B0(mai_mai_n160_), .Y(mai_mai_n574_));
  OR2        m552(.A(i_6_), .B(i_10_), .Y(mai_mai_n575_));
  NO2        m553(.A(mai_mai_n575_), .B(mai_mai_n23_), .Y(mai_mai_n576_));
  OR3        m554(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n577_));
  NO3        m555(.A(mai_mai_n577_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n578_));
  NO2        m556(.A(mai_mai_n578_), .B(mai_mai_n576_), .Y(mai_mai_n579_));
  OA220      m557(.A0(mai_mai_n579_), .A1(mai_mai_n550_), .B0(mai_mai_n574_), .B1(mai_mai_n259_), .Y(mai_mai_n580_));
  AOI210     m558(.A0(mai_mai_n580_), .A1(mai_mai_n572_), .B0(mai_mai_n64_), .Y(mai_mai_n581_));
  NOi21      m559(.An(i_11_), .B(i_7_), .Y(mai_mai_n582_));
  AO210      m560(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n583_));
  NO2        m561(.A(mai_mai_n583_), .B(mai_mai_n582_), .Y(mai_mai_n584_));
  NA2        m562(.A(mai_mai_n584_), .B(mai_mai_n197_), .Y(mai_mai_n585_));
  NA3        m563(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n586_));
  NAi31      m564(.An(mai_mai_n586_), .B(mai_mai_n206_), .C(i_11_), .Y(mai_mai_n587_));
  AOI210     m565(.A0(mai_mai_n587_), .A1(mai_mai_n585_), .B0(mai_mai_n64_), .Y(mai_mai_n588_));
  NA2        m566(.A(mai_mai_n89_), .B(mai_mai_n64_), .Y(mai_mai_n589_));
  AO210      m567(.A0(mai_mai_n589_), .A1(mai_mai_n357_), .B0(mai_mai_n41_), .Y(mai_mai_n590_));
  NA2        m568(.A(mai_mai_n218_), .B(mai_mai_n64_), .Y(mai_mai_n591_));
  NA2        m569(.A(mai_mai_n390_), .B(mai_mai_n31_), .Y(mai_mai_n592_));
  OR2        m570(.A(mai_mai_n199_), .B(mai_mai_n112_), .Y(mai_mai_n593_));
  NA2        m571(.A(mai_mai_n593_), .B(mai_mai_n592_), .Y(mai_mai_n594_));
  NO2        m572(.A(mai_mai_n64_), .B(i_9_), .Y(mai_mai_n595_));
  NO2        m573(.A(mai_mai_n595_), .B(i_4_), .Y(mai_mai_n596_));
  NA2        m574(.A(mai_mai_n596_), .B(mai_mai_n594_), .Y(mai_mai_n597_));
  NO2        m575(.A(i_1_), .B(i_12_), .Y(mai_mai_n598_));
  NA3        m576(.A(mai_mai_n598_), .B(mai_mai_n113_), .C(mai_mai_n24_), .Y(mai_mai_n599_));
  BUFFER     m577(.A(mai_mai_n599_), .Y(mai_mai_n600_));
  NA4        m578(.A(mai_mai_n600_), .B(mai_mai_n597_), .C(mai_mai_n591_), .D(mai_mai_n590_), .Y(mai_mai_n601_));
  OAI210     m579(.A0(mai_mai_n601_), .A1(mai_mai_n588_), .B0(i_6_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n586_), .B(mai_mai_n112_), .Y(mai_mai_n603_));
  NA2        m581(.A(mai_mai_n603_), .B(mai_mai_n551_), .Y(mai_mai_n604_));
  NO2        m582(.A(i_6_), .B(i_11_), .Y(mai_mai_n605_));
  NA2        m583(.A(mai_mai_n604_), .B(mai_mai_n430_), .Y(mai_mai_n606_));
  NO4        m584(.A(mai_mai_n206_), .B(mai_mai_n132_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n607_));
  NA2        m585(.A(mai_mai_n607_), .B(mai_mai_n595_), .Y(mai_mai_n608_));
  NO3        m586(.A(mai_mai_n575_), .B(mai_mai_n225_), .C(mai_mai_n23_), .Y(mai_mai_n609_));
  AOI210     m587(.A0(i_1_), .A1(mai_mai_n250_), .B0(mai_mai_n609_), .Y(mai_mai_n610_));
  OAI210     m588(.A0(mai_mai_n610_), .A1(mai_mai_n45_), .B0(mai_mai_n608_), .Y(mai_mai_n611_));
  NA3        m589(.A(mai_mai_n507_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n612_));
  INV        m590(.A(i_2_), .Y(mai_mai_n613_));
  NA2        m591(.A(mai_mai_n142_), .B(i_9_), .Y(mai_mai_n614_));
  NA3        m592(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n615_));
  NO2        m593(.A(mai_mai_n47_), .B(i_1_), .Y(mai_mai_n616_));
  NA3        m594(.A(mai_mai_n616_), .B(mai_mai_n258_), .C(mai_mai_n45_), .Y(mai_mai_n617_));
  OAI220     m595(.A0(mai_mai_n617_), .A1(mai_mai_n615_), .B0(mai_mai_n614_), .B1(mai_mai_n613_), .Y(mai_mai_n618_));
  AOI210     m596(.A0(mai_mai_n454_), .A1(mai_mai_n400_), .B0(mai_mai_n232_), .Y(mai_mai_n619_));
  NO2        m597(.A(mai_mai_n619_), .B(mai_mai_n566_), .Y(mai_mai_n620_));
  NAi21      m598(.An(mai_mai_n612_), .B(mai_mai_n95_), .Y(mai_mai_n621_));
  NO2        m599(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n622_));
  INV        m600(.A(mai_mai_n621_), .Y(mai_mai_n623_));
  OR3        m601(.A(mai_mai_n623_), .B(mai_mai_n620_), .C(mai_mai_n618_), .Y(mai_mai_n624_));
  NO3        m602(.A(mai_mai_n624_), .B(mai_mai_n611_), .C(mai_mai_n606_), .Y(mai_mai_n625_));
  NO2        m603(.A(mai_mai_n228_), .B(mai_mai_n105_), .Y(mai_mai_n626_));
  NO2        m604(.A(mai_mai_n626_), .B(mai_mai_n582_), .Y(mai_mai_n627_));
  NA2        m605(.A(mai_mai_n627_), .B(i_1_), .Y(mai_mai_n628_));
  NO2        m606(.A(mai_mai_n628_), .B(mai_mai_n577_), .Y(mai_mai_n629_));
  NO2        m607(.A(mai_mai_n396_), .B(mai_mai_n87_), .Y(mai_mai_n630_));
  NA2        m608(.A(mai_mai_n629_), .B(mai_mai_n47_), .Y(mai_mai_n631_));
  NA2        m609(.A(i_3_), .B(mai_mai_n187_), .Y(mai_mai_n632_));
  NO2        m610(.A(mai_mai_n632_), .B(mai_mai_n118_), .Y(mai_mai_n633_));
  AN2        m611(.A(mai_mai_n633_), .B(mai_mai_n509_), .Y(mai_mai_n634_));
  NO2        m612(.A(mai_mai_n225_), .B(mai_mai_n45_), .Y(mai_mai_n635_));
  NO3        m613(.A(mai_mai_n635_), .B(mai_mai_n292_), .C(mai_mai_n229_), .Y(mai_mai_n636_));
  NO2        m614(.A(mai_mai_n121_), .B(mai_mai_n37_), .Y(mai_mai_n637_));
  NO2        m615(.A(mai_mai_n637_), .B(i_6_), .Y(mai_mai_n638_));
  NO2        m616(.A(mai_mai_n87_), .B(i_9_), .Y(mai_mai_n639_));
  NO2        m617(.A(mai_mai_n639_), .B(mai_mai_n64_), .Y(mai_mai_n640_));
  NO2        m618(.A(mai_mai_n640_), .B(mai_mai_n598_), .Y(mai_mai_n641_));
  NO4        m619(.A(mai_mai_n641_), .B(mai_mai_n638_), .C(mai_mai_n636_), .D(i_4_), .Y(mai_mai_n642_));
  NA2        m620(.A(i_1_), .B(i_3_), .Y(mai_mai_n643_));
  NO2        m621(.A(mai_mai_n642_), .B(mai_mai_n634_), .Y(mai_mai_n644_));
  NA4        m622(.A(mai_mai_n644_), .B(mai_mai_n631_), .C(mai_mai_n625_), .D(mai_mai_n602_), .Y(mai_mai_n645_));
  NO3        m623(.A(mai_mai_n455_), .B(i_3_), .C(i_7_), .Y(mai_mai_n646_));
  NOi21      m624(.An(mai_mai_n646_), .B(i_10_), .Y(mai_mai_n647_));
  OA210      m625(.A0(mai_mai_n647_), .A1(mai_mai_n235_), .B0(mai_mai_n87_), .Y(mai_mai_n648_));
  NA2        m626(.A(mai_mai_n349_), .B(mai_mai_n348_), .Y(mai_mai_n649_));
  NA3        m627(.A(mai_mai_n462_), .B(mai_mai_n492_), .C(mai_mai_n47_), .Y(mai_mai_n650_));
  NO3        m628(.A(mai_mai_n456_), .B(mai_mai_n569_), .C(mai_mai_n87_), .Y(mai_mai_n651_));
  NA2        m629(.A(mai_mai_n651_), .B(mai_mai_n25_), .Y(mai_mai_n652_));
  NA3        m630(.A(mai_mai_n160_), .B(mai_mai_n85_), .C(mai_mai_n87_), .Y(mai_mai_n653_));
  NA4        m631(.A(mai_mai_n653_), .B(mai_mai_n652_), .C(mai_mai_n650_), .D(mai_mai_n649_), .Y(mai_mai_n654_));
  OAI210     m632(.A0(mai_mai_n654_), .A1(mai_mai_n648_), .B0(i_1_), .Y(mai_mai_n655_));
  AOI210     m633(.A0(mai_mai_n258_), .A1(mai_mai_n101_), .B0(i_1_), .Y(mai_mai_n656_));
  NO2        m634(.A(mai_mai_n347_), .B(i_2_), .Y(mai_mai_n657_));
  NA2        m635(.A(mai_mai_n657_), .B(mai_mai_n656_), .Y(mai_mai_n658_));
  AOI210     m636(.A0(mai_mai_n658_), .A1(mai_mai_n655_), .B0(i_13_), .Y(mai_mai_n659_));
  OR2        m637(.A(i_11_), .B(i_7_), .Y(mai_mai_n660_));
  NA3        m638(.A(mai_mai_n660_), .B(mai_mai_n110_), .C(mai_mai_n142_), .Y(mai_mai_n661_));
  AOI220     m639(.A0(mai_mai_n449_), .A1(mai_mai_n160_), .B0(mai_mai_n424_), .B1(mai_mai_n142_), .Y(mai_mai_n662_));
  OAI210     m640(.A0(mai_mai_n662_), .A1(mai_mai_n45_), .B0(mai_mai_n661_), .Y(mai_mai_n663_));
  NO2        m641(.A(mai_mai_n55_), .B(i_12_), .Y(mai_mai_n664_));
  INV        m642(.A(mai_mai_n664_), .Y(mai_mai_n665_));
  NO2        m643(.A(mai_mai_n456_), .B(mai_mai_n24_), .Y(mai_mai_n666_));
  NA2        m644(.A(mai_mai_n666_), .B(mai_mai_n630_), .Y(mai_mai_n667_));
  OAI220     m645(.A0(mai_mai_n667_), .A1(mai_mai_n41_), .B0(mai_mai_n665_), .B1(mai_mai_n96_), .Y(mai_mai_n668_));
  AOI210     m646(.A0(mai_mai_n663_), .A1(mai_mai_n315_), .B0(mai_mai_n668_), .Y(mai_mai_n669_));
  INV        m647(.A(mai_mai_n118_), .Y(mai_mai_n670_));
  AOI220     m648(.A0(mai_mai_n670_), .A1(mai_mai_n73_), .B0(mai_mai_n365_), .B1(mai_mai_n616_), .Y(mai_mai_n671_));
  NO2        m649(.A(mai_mai_n671_), .B(mai_mai_n233_), .Y(mai_mai_n672_));
  NA2        m650(.A(mai_mai_n131_), .B(i_13_), .Y(mai_mai_n673_));
  NO2        m651(.A(mai_mai_n615_), .B(mai_mai_n118_), .Y(mai_mai_n674_));
  INV        m652(.A(mai_mai_n674_), .Y(mai_mai_n675_));
  OAI220     m653(.A0(mai_mai_n675_), .A1(mai_mai_n72_), .B0(mai_mai_n673_), .B1(mai_mai_n656_), .Y(mai_mai_n676_));
  NA2        m654(.A(mai_mai_n26_), .B(mai_mai_n187_), .Y(mai_mai_n677_));
  NA2        m655(.A(mai_mai_n677_), .B(i_7_), .Y(mai_mai_n678_));
  AOI220     m656(.A0(mai_mai_n365_), .A1(mai_mai_n616_), .B0(mai_mai_n95_), .B1(mai_mai_n106_), .Y(mai_mai_n679_));
  NO2        m657(.A(mai_mai_n679_), .B(mai_mai_n564_), .Y(mai_mai_n680_));
  NO3        m658(.A(mai_mai_n680_), .B(mai_mai_n676_), .C(mai_mai_n672_), .Y(mai_mai_n681_));
  OR2        m659(.A(i_11_), .B(i_6_), .Y(mai_mai_n682_));
  NA3        m660(.A(mai_mai_n563_), .B(mai_mai_n677_), .C(i_7_), .Y(mai_mai_n683_));
  AOI210     m661(.A0(mai_mai_n683_), .A1(mai_mai_n675_), .B0(mai_mai_n682_), .Y(mai_mai_n684_));
  NA3        m662(.A(mai_mai_n390_), .B(mai_mai_n568_), .C(mai_mai_n101_), .Y(mai_mai_n685_));
  NA2        m663(.A(mai_mai_n605_), .B(i_13_), .Y(mai_mai_n686_));
  NA2        m664(.A(mai_mai_n106_), .B(mai_mai_n677_), .Y(mai_mai_n687_));
  NAi21      m665(.An(i_11_), .B(i_12_), .Y(mai_mai_n688_));
  NOi41      m666(.An(mai_mai_n114_), .B(mai_mai_n688_), .C(i_13_), .D(mai_mai_n87_), .Y(mai_mai_n689_));
  NA2        m667(.A(mai_mai_n689_), .B(mai_mai_n687_), .Y(mai_mai_n690_));
  NA3        m668(.A(mai_mai_n690_), .B(mai_mai_n686_), .C(mai_mai_n685_), .Y(mai_mai_n691_));
  OAI210     m669(.A0(mai_mai_n691_), .A1(mai_mai_n684_), .B0(mai_mai_n64_), .Y(mai_mai_n692_));
  NO2        m670(.A(i_2_), .B(i_12_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n346_), .B(mai_mai_n693_), .Y(mai_mai_n694_));
  NA2        m672(.A(i_8_), .B(mai_mai_n25_), .Y(mai_mai_n695_));
  NO3        m673(.A(mai_mai_n695_), .B(mai_mai_n363_), .C(mai_mai_n563_), .Y(mai_mai_n696_));
  OAI210     m674(.A0(mai_mai_n696_), .A1(mai_mai_n348_), .B0(mai_mai_n346_), .Y(mai_mai_n697_));
  NO2        m675(.A(mai_mai_n132_), .B(i_2_), .Y(mai_mai_n698_));
  NA2        m676(.A(mai_mai_n697_), .B(mai_mai_n694_), .Y(mai_mai_n699_));
  NA3        m677(.A(mai_mai_n699_), .B(mai_mai_n46_), .C(mai_mai_n217_), .Y(mai_mai_n700_));
  NA4        m678(.A(mai_mai_n700_), .B(mai_mai_n692_), .C(mai_mai_n681_), .D(mai_mai_n669_), .Y(mai_mai_n701_));
  OR4        m679(.A(mai_mai_n701_), .B(mai_mai_n659_), .C(mai_mai_n645_), .D(mai_mai_n581_), .Y(mai5));
  NA2        m680(.A(mai_mai_n627_), .B(mai_mai_n260_), .Y(mai_mai_n703_));
  AN2        m681(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n704_));
  NA3        m682(.A(mai_mai_n704_), .B(mai_mai_n693_), .C(mai_mai_n112_), .Y(mai_mai_n705_));
  NO2        m683(.A(mai_mai_n564_), .B(i_11_), .Y(mai_mai_n706_));
  NA2        m684(.A(mai_mai_n90_), .B(mai_mai_n706_), .Y(mai_mai_n707_));
  NA3        m685(.A(mai_mai_n707_), .B(mai_mai_n705_), .C(mai_mai_n703_), .Y(mai_mai_n708_));
  NO3        m686(.A(i_11_), .B(mai_mai_n228_), .C(i_13_), .Y(mai_mai_n709_));
  NO2        m687(.A(mai_mai_n128_), .B(mai_mai_n23_), .Y(mai_mai_n710_));
  NA2        m688(.A(i_12_), .B(i_8_), .Y(mai_mai_n711_));
  OAI210     m689(.A0(mai_mai_n47_), .A1(i_3_), .B0(mai_mai_n711_), .Y(mai_mai_n712_));
  INV        m690(.A(mai_mai_n420_), .Y(mai_mai_n713_));
  AOI220     m691(.A0(mai_mai_n301_), .A1(mai_mai_n545_), .B0(mai_mai_n712_), .B1(mai_mai_n710_), .Y(mai_mai_n714_));
  INV        m692(.A(mai_mai_n714_), .Y(mai_mai_n715_));
  NO2        m693(.A(mai_mai_n715_), .B(mai_mai_n708_), .Y(mai_mai_n716_));
  INV        m694(.A(mai_mai_n169_), .Y(mai_mai_n717_));
  INV        m695(.A(mai_mai_n235_), .Y(mai_mai_n718_));
  OAI210     m696(.A0(mai_mai_n657_), .A1(mai_mai_n422_), .B0(mai_mai_n114_), .Y(mai_mai_n719_));
  AOI210     m697(.A0(mai_mai_n719_), .A1(mai_mai_n718_), .B0(mai_mai_n717_), .Y(mai_mai_n720_));
  NO2        m698(.A(mai_mai_n431_), .B(mai_mai_n26_), .Y(mai_mai_n721_));
  NO2        m699(.A(mai_mai_n721_), .B(mai_mai_n400_), .Y(mai_mai_n722_));
  NA2        m700(.A(mai_mai_n722_), .B(i_2_), .Y(mai_mai_n723_));
  INV        m701(.A(mai_mai_n723_), .Y(mai_mai_n724_));
  AOI210     m702(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n397_), .Y(mai_mai_n725_));
  AOI210     m703(.A0(mai_mai_n725_), .A1(mai_mai_n724_), .B0(mai_mai_n720_), .Y(mai_mai_n726_));
  NO2        m704(.A(mai_mai_n184_), .B(mai_mai_n129_), .Y(mai_mai_n727_));
  OAI210     m705(.A0(mai_mai_n727_), .A1(mai_mai_n710_), .B0(i_2_), .Y(mai_mai_n728_));
  INV        m706(.A(mai_mai_n170_), .Y(mai_mai_n729_));
  NO3        m707(.A(mai_mai_n583_), .B(mai_mai_n38_), .C(mai_mai_n26_), .Y(mai_mai_n730_));
  AOI210     m708(.A0(mai_mai_n729_), .A1(mai_mai_n90_), .B0(mai_mai_n730_), .Y(mai_mai_n731_));
  AOI210     m709(.A0(mai_mai_n731_), .A1(mai_mai_n728_), .B0(mai_mai_n187_), .Y(mai_mai_n732_));
  OA210      m710(.A0(mai_mai_n584_), .A1(mai_mai_n130_), .B0(i_13_), .Y(mai_mai_n733_));
  NA2        m711(.A(mai_mai_n156_), .B(mai_mai_n561_), .Y(mai_mai_n734_));
  NO2        m712(.A(mai_mai_n734_), .B(mai_mai_n351_), .Y(mai_mai_n735_));
  AOI210     m713(.A0(mai_mai_n199_), .A1(mai_mai_n152_), .B0(mai_mai_n492_), .Y(mai_mai_n736_));
  NA2        m714(.A(mai_mai_n736_), .B(mai_mai_n400_), .Y(mai_mai_n737_));
  NO2        m715(.A(mai_mai_n106_), .B(mai_mai_n45_), .Y(mai_mai_n738_));
  INV        m716(.A(mai_mai_n286_), .Y(mai_mai_n739_));
  NA4        m717(.A(mai_mai_n739_), .B(mai_mai_n289_), .C(mai_mai_n128_), .D(mai_mai_n43_), .Y(mai_mai_n740_));
  OAI210     m718(.A0(mai_mai_n740_), .A1(mai_mai_n738_), .B0(mai_mai_n737_), .Y(mai_mai_n741_));
  NO4        m719(.A(mai_mai_n741_), .B(mai_mai_n735_), .C(mai_mai_n733_), .D(mai_mai_n732_), .Y(mai_mai_n742_));
  NA2        m720(.A(mai_mai_n545_), .B(mai_mai_n28_), .Y(mai_mai_n743_));
  NA2        m721(.A(mai_mai_n709_), .B(mai_mai_n263_), .Y(mai_mai_n744_));
  NA2        m722(.A(mai_mai_n744_), .B(mai_mai_n743_), .Y(mai_mai_n745_));
  NO2        m723(.A(mai_mai_n63_), .B(i_12_), .Y(mai_mai_n746_));
  NO2        m724(.A(mai_mai_n746_), .B(mai_mai_n130_), .Y(mai_mai_n747_));
  NO2        m725(.A(mai_mai_n747_), .B(mai_mai_n561_), .Y(mai_mai_n748_));
  AOI220     m726(.A0(mai_mai_n748_), .A1(mai_mai_n36_), .B0(mai_mai_n745_), .B1(mai_mai_n47_), .Y(mai_mai_n749_));
  NA4        m727(.A(mai_mai_n749_), .B(mai_mai_n742_), .C(mai_mai_n726_), .D(mai_mai_n716_), .Y(mai6));
  NA4        m728(.A(mai_mai_n369_), .B(mai_mai_n461_), .C(mai_mai_n72_), .D(mai_mai_n105_), .Y(mai_mai_n751_));
  INV        m729(.A(mai_mai_n751_), .Y(mai_mai_n752_));
  NO2        m730(.A(mai_mai_n212_), .B(mai_mai_n464_), .Y(mai_mai_n753_));
  NO2        m731(.A(mai_mai_n752_), .B(mai_mai_n313_), .Y(mai_mai_n754_));
  OR2        m732(.A(mai_mai_n754_), .B(i_12_), .Y(mai_mai_n755_));
  NA2        m733(.A(mai_mai_n352_), .B(mai_mai_n318_), .Y(mai_mai_n756_));
  NA2        m734(.A(mai_mai_n551_), .B(mai_mai_n64_), .Y(mai_mai_n757_));
  NA2        m735(.A(mai_mai_n647_), .B(mai_mai_n72_), .Y(mai_mai_n758_));
  BUFFER     m736(.A(mai_mai_n589_), .Y(mai_mai_n759_));
  NA4        m737(.A(mai_mai_n759_), .B(mai_mai_n758_), .C(mai_mai_n757_), .D(mai_mai_n756_), .Y(mai_mai_n760_));
  NA2        m738(.A(mai_mai_n760_), .B(mai_mai_n74_), .Y(mai_mai_n761_));
  INV        m739(.A(mai_mai_n312_), .Y(mai_mai_n762_));
  NA2        m740(.A(mai_mai_n76_), .B(mai_mai_n135_), .Y(mai_mai_n763_));
  INV        m741(.A(mai_mai_n128_), .Y(mai_mai_n764_));
  NA2        m742(.A(mai_mai_n764_), .B(mai_mai_n47_), .Y(mai_mai_n765_));
  AOI210     m743(.A0(mai_mai_n765_), .A1(mai_mai_n763_), .B0(mai_mai_n762_), .Y(mai_mai_n766_));
  NO2        m744(.A(mai_mai_n242_), .B(i_9_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n767_), .B(mai_mai_n746_), .Y(mai_mai_n768_));
  AOI210     m746(.A0(mai_mai_n768_), .A1(mai_mai_n491_), .B0(mai_mai_n181_), .Y(mai_mai_n769_));
  NO2        m747(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n770_));
  NA3        m748(.A(mai_mai_n770_), .B(mai_mai_n452_), .C(mai_mai_n369_), .Y(mai_mai_n771_));
  NAi32      m749(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n772_));
  NO2        m750(.A(mai_mai_n682_), .B(mai_mai_n772_), .Y(mai_mai_n773_));
  NAi21      m751(.An(mai_mai_n773_), .B(mai_mai_n771_), .Y(mai_mai_n774_));
  OR3        m752(.A(mai_mai_n774_), .B(mai_mai_n769_), .C(mai_mai_n766_), .Y(mai_mai_n775_));
  NO2        m753(.A(mai_mai_n660_), .B(i_2_), .Y(mai_mai_n776_));
  OR2        m754(.A(mai_mai_n584_), .B(mai_mai_n422_), .Y(mai_mai_n777_));
  NA3        m755(.A(mai_mai_n777_), .B(mai_mai_n151_), .C(mai_mai_n70_), .Y(mai_mai_n778_));
  AO210      m756(.A0(mai_mai_n470_), .A1(mai_mai_n713_), .B0(mai_mai_n36_), .Y(mai_mai_n779_));
  NA2        m757(.A(mai_mai_n779_), .B(mai_mai_n778_), .Y(mai_mai_n780_));
  OAI210     m758(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n88_), .Y(mai_mai_n781_));
  AOI220     m759(.A0(mai_mai_n781_), .A1(mai_mai_n532_), .B0(mai_mai_n753_), .B1(mai_mai_n678_), .Y(mai_mai_n782_));
  NA2        m760(.A(mai_mai_n377_), .B(mai_mai_n71_), .Y(mai_mai_n783_));
  NA3        m761(.A(mai_mai_n783_), .B(mai_mai_n782_), .C(mai_mai_n567_), .Y(mai_mai_n784_));
  AO210      m762(.A0(mai_mai_n492_), .A1(mai_mai_n47_), .B0(mai_mai_n89_), .Y(mai_mai_n785_));
  NA3        m763(.A(mai_mai_n785_), .B(mai_mai_n462_), .C(mai_mai_n209_), .Y(mai_mai_n786_));
  AOI210     m764(.A0(mai_mai_n422_), .A1(mai_mai_n420_), .B0(mai_mai_n531_), .Y(mai_mai_n787_));
  NA2        m765(.A(mai_mai_n115_), .B(mai_mai_n387_), .Y(mai_mai_n788_));
  NA2        m766(.A(mai_mai_n234_), .B(mai_mai_n47_), .Y(mai_mai_n789_));
  INV        m767(.A(mai_mai_n553_), .Y(mai_mai_n790_));
  NA3        m768(.A(mai_mai_n790_), .B(mai_mai_n312_), .C(i_7_), .Y(mai_mai_n791_));
  NA4        m769(.A(mai_mai_n791_), .B(mai_mai_n788_), .C(mai_mai_n787_), .D(mai_mai_n786_), .Y(mai_mai_n792_));
  NO4        m770(.A(mai_mai_n792_), .B(mai_mai_n784_), .C(mai_mai_n780_), .D(mai_mai_n775_), .Y(mai_mai_n793_));
  NA4        m771(.A(mai_mai_n793_), .B(mai_mai_n761_), .C(mai_mai_n755_), .D(mai_mai_n359_), .Y(mai3));
  NA2        m772(.A(i_12_), .B(i_10_), .Y(mai_mai_n795_));
  NA2        m773(.A(i_6_), .B(i_7_), .Y(mai_mai_n796_));
  NO2        m774(.A(mai_mai_n796_), .B(i_0_), .Y(mai_mai_n797_));
  NO2        m775(.A(i_11_), .B(mai_mai_n228_), .Y(mai_mai_n798_));
  OAI210     m776(.A0(mai_mai_n797_), .A1(mai_mai_n274_), .B0(mai_mai_n798_), .Y(mai_mai_n799_));
  NO2        m777(.A(mai_mai_n799_), .B(mai_mai_n187_), .Y(mai_mai_n800_));
  NO3        m778(.A(mai_mai_n427_), .B(mai_mai_n93_), .C(mai_mai_n45_), .Y(mai_mai_n801_));
  OA210      m779(.A0(mai_mai_n801_), .A1(mai_mai_n800_), .B0(mai_mai_n172_), .Y(mai_mai_n802_));
  NA2        m780(.A(mai_mai_n567_), .B(mai_mai_n350_), .Y(mai_mai_n803_));
  NA2        m781(.A(mai_mai_n803_), .B(mai_mai_n40_), .Y(mai_mai_n804_));
  NOi21      m782(.An(mai_mai_n100_), .B(mai_mai_n722_), .Y(mai_mai_n805_));
  NO3        m783(.A(mai_mai_n593_), .B(mai_mai_n431_), .C(mai_mai_n135_), .Y(mai_mai_n806_));
  AN2        m784(.A(mai_mai_n429_), .B(mai_mai_n56_), .Y(mai_mai_n807_));
  NO3        m785(.A(mai_mai_n807_), .B(mai_mai_n806_), .C(mai_mai_n805_), .Y(mai_mai_n808_));
  AOI210     m786(.A0(mai_mai_n808_), .A1(mai_mai_n804_), .B0(mai_mai_n49_), .Y(mai_mai_n809_));
  NO4        m787(.A(mai_mai_n355_), .B(mai_mai_n362_), .C(mai_mai_n38_), .D(i_0_), .Y(mai_mai_n810_));
  NA2        m788(.A(mai_mai_n181_), .B(mai_mai_n541_), .Y(mai_mai_n811_));
  NOi21      m789(.An(mai_mai_n811_), .B(mai_mai_n810_), .Y(mai_mai_n812_));
  NO2        m790(.A(mai_mai_n812_), .B(mai_mai_n64_), .Y(mai_mai_n813_));
  NOi21      m791(.An(i_5_), .B(i_9_), .Y(mai_mai_n814_));
  NA2        m792(.A(mai_mai_n814_), .B(mai_mai_n418_), .Y(mai_mai_n815_));
  BUFFER     m793(.A(mai_mai_n258_), .Y(mai_mai_n816_));
  AOI210     m794(.A0(mai_mai_n816_), .A1(mai_mai_n454_), .B0(mai_mai_n651_), .Y(mai_mai_n817_));
  NO3        m795(.A(mai_mai_n393_), .B(mai_mai_n258_), .C(mai_mai_n74_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n173_), .B(mai_mai_n152_), .Y(mai_mai_n819_));
  AOI210     m797(.A0(mai_mai_n819_), .A1(mai_mai_n234_), .B0(mai_mai_n818_), .Y(mai_mai_n820_));
  OAI220     m798(.A0(mai_mai_n820_), .A1(mai_mai_n179_), .B0(mai_mai_n817_), .B1(mai_mai_n815_), .Y(mai_mai_n821_));
  NO4        m799(.A(mai_mai_n821_), .B(mai_mai_n813_), .C(mai_mai_n809_), .D(mai_mai_n802_), .Y(mai_mai_n822_));
  NA2        m800(.A(mai_mai_n181_), .B(mai_mai_n24_), .Y(mai_mai_n823_));
  NAi21      m801(.An(mai_mai_n161_), .B(mai_mai_n410_), .Y(mai_mai_n824_));
  NO2        m802(.A(mai_mai_n824_), .B(mai_mai_n789_), .Y(mai_mai_n825_));
  INV        m803(.A(mai_mai_n825_), .Y(mai_mai_n826_));
  NO2        m804(.A(mai_mai_n369_), .B(mai_mai_n278_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n827_), .B(mai_mai_n674_), .Y(mai_mai_n828_));
  NA2        m806(.A(mai_mai_n542_), .B(i_0_), .Y(mai_mai_n829_));
  NO4        m807(.A(mai_mai_n552_), .B(mai_mai_n206_), .C(mai_mai_n397_), .D(mai_mai_n389_), .Y(mai_mai_n830_));
  NA2        m808(.A(mai_mai_n830_), .B(i_11_), .Y(mai_mai_n831_));
  INV        m809(.A(mai_mai_n452_), .Y(mai_mai_n832_));
  NA2        m810(.A(mai_mai_n709_), .B(mai_mai_n313_), .Y(mai_mai_n833_));
  INV        m811(.A(mai_mai_n59_), .Y(mai_mai_n834_));
  NO2        m812(.A(mai_mai_n834_), .B(mai_mai_n833_), .Y(mai_mai_n835_));
  NO2        m813(.A(mai_mai_n244_), .B(mai_mai_n157_), .Y(mai_mai_n836_));
  NA2        m814(.A(i_0_), .B(i_10_), .Y(mai_mai_n837_));
  INV        m815(.A(mai_mai_n508_), .Y(mai_mai_n838_));
  NO4        m816(.A(mai_mai_n118_), .B(mai_mai_n59_), .C(mai_mai_n632_), .D(i_5_), .Y(mai_mai_n839_));
  AO220      m817(.A0(mai_mai_n839_), .A1(mai_mai_n838_), .B0(mai_mai_n836_), .B1(i_6_), .Y(mai_mai_n840_));
  AOI220     m818(.A0(mai_mai_n316_), .A1(mai_mai_n102_), .B0(mai_mai_n181_), .B1(mai_mai_n85_), .Y(mai_mai_n841_));
  NA2        m819(.A(mai_mai_n536_), .B(i_4_), .Y(mai_mai_n842_));
  NA2        m820(.A(mai_mai_n182_), .B(mai_mai_n192_), .Y(mai_mai_n843_));
  OAI220     m821(.A0(mai_mai_n843_), .A1(mai_mai_n833_), .B0(mai_mai_n842_), .B1(mai_mai_n841_), .Y(mai_mai_n844_));
  NO3        m822(.A(mai_mai_n844_), .B(mai_mai_n840_), .C(mai_mai_n835_), .Y(mai_mai_n845_));
  NA4        m823(.A(mai_mai_n845_), .B(mai_mai_n831_), .C(mai_mai_n828_), .D(mai_mai_n826_), .Y(mai_mai_n846_));
  NO2        m824(.A(mai_mai_n107_), .B(mai_mai_n37_), .Y(mai_mai_n847_));
  NA2        m825(.A(i_11_), .B(i_9_), .Y(mai_mai_n848_));
  NO3        m826(.A(i_12_), .B(mai_mai_n848_), .C(mai_mai_n566_), .Y(mai_mai_n849_));
  AN2        m827(.A(mai_mai_n849_), .B(mai_mai_n847_), .Y(mai_mai_n850_));
  NO2        m828(.A(mai_mai_n49_), .B(i_7_), .Y(mai_mai_n851_));
  NA2        m829(.A(mai_mai_n374_), .B(mai_mai_n177_), .Y(mai_mai_n852_));
  INV        m830(.A(mai_mai_n852_), .Y(mai_mai_n853_));
  NO2        m831(.A(mai_mai_n848_), .B(mai_mai_n74_), .Y(mai_mai_n854_));
  NO2        m832(.A(mai_mai_n173_), .B(i_0_), .Y(mai_mai_n855_));
  INV        m833(.A(mai_mai_n855_), .Y(mai_mai_n856_));
  NA2        m834(.A(mai_mai_n452_), .B(mai_mai_n223_), .Y(mai_mai_n857_));
  AOI210     m835(.A0(mai_mai_n349_), .A1(mai_mai_n42_), .B0(mai_mai_n386_), .Y(mai_mai_n858_));
  OAI220     m836(.A0(mai_mai_n858_), .A1(mai_mai_n815_), .B0(mai_mai_n857_), .B1(mai_mai_n856_), .Y(mai_mai_n859_));
  NO3        m837(.A(mai_mai_n859_), .B(mai_mai_n853_), .C(mai_mai_n850_), .Y(mai_mai_n860_));
  NA2        m838(.A(mai_mai_n622_), .B(mai_mai_n125_), .Y(mai_mai_n861_));
  NO2        m839(.A(i_6_), .B(mai_mai_n861_), .Y(mai_mai_n862_));
  NA2        m840(.A(mai_mai_n169_), .B(mai_mai_n107_), .Y(mai_mai_n863_));
  INV        m841(.A(mai_mai_n862_), .Y(mai_mai_n864_));
  NOi21      m842(.An(i_7_), .B(i_5_), .Y(mai_mai_n865_));
  NOi31      m843(.An(mai_mai_n865_), .B(i_0_), .C(mai_mai_n688_), .Y(mai_mai_n866_));
  NA3        m844(.A(mai_mai_n866_), .B(mai_mai_n363_), .C(i_6_), .Y(mai_mai_n867_));
  OA210      m845(.A0(mai_mai_n863_), .A1(mai_mai_n491_), .B0(mai_mai_n867_), .Y(mai_mai_n868_));
  NO3        m846(.A(mai_mai_n381_), .B(mai_mai_n338_), .C(mai_mai_n336_), .Y(mai_mai_n869_));
  NO2        m847(.A(mai_mai_n253_), .B(mai_mai_n302_), .Y(mai_mai_n870_));
  NO2        m848(.A(mai_mai_n688_), .B(mai_mai_n248_), .Y(mai_mai_n871_));
  AOI210     m849(.A0(mai_mai_n871_), .A1(mai_mai_n870_), .B0(mai_mai_n869_), .Y(mai_mai_n872_));
  NA4        m850(.A(mai_mai_n872_), .B(mai_mai_n868_), .C(mai_mai_n864_), .D(mai_mai_n860_), .Y(mai_mai_n873_));
  NO2        m851(.A(mai_mai_n823_), .B(mai_mai_n231_), .Y(mai_mai_n874_));
  AN2        m852(.A(mai_mai_n315_), .B(mai_mai_n313_), .Y(mai_mai_n875_));
  AN2        m853(.A(mai_mai_n875_), .B(mai_mai_n819_), .Y(mai_mai_n876_));
  OAI210     m854(.A0(mai_mai_n876_), .A1(mai_mai_n874_), .B0(i_10_), .Y(mai_mai_n877_));
  NO2        m855(.A(mai_mai_n795_), .B(mai_mai_n301_), .Y(mai_mai_n878_));
  OA210      m856(.A0(mai_mai_n452_), .A1(mai_mai_n215_), .B0(mai_mai_n451_), .Y(mai_mai_n879_));
  NA2        m857(.A(mai_mai_n878_), .B(mai_mai_n854_), .Y(mai_mai_n880_));
  NA3        m858(.A(mai_mai_n451_), .B(mai_mai_n390_), .C(mai_mai_n46_), .Y(mai_mai_n881_));
  OAI210     m859(.A0(mai_mai_n824_), .A1(mai_mai_n832_), .B0(mai_mai_n881_), .Y(mai_mai_n882_));
  NA2        m860(.A(mai_mai_n854_), .B(mai_mai_n289_), .Y(mai_mai_n883_));
  INV        m861(.A(mai_mai_n883_), .Y(mai_mai_n884_));
  AOI220     m862(.A0(mai_mai_n884_), .A1(mai_mai_n452_), .B0(mai_mai_n882_), .B1(mai_mai_n74_), .Y(mai_mai_n885_));
  NA2        m863(.A(mai_mai_n666_), .B(mai_mai_n513_), .Y(mai_mai_n886_));
  NAi21      m864(.An(i_9_), .B(i_5_), .Y(mai_mai_n887_));
  NO2        m865(.A(mai_mai_n887_), .B(mai_mai_n381_), .Y(mai_mai_n888_));
  NO2        m866(.A(mai_mai_n562_), .B(mai_mai_n109_), .Y(mai_mai_n889_));
  AOI220     m867(.A0(mai_mai_n889_), .A1(i_0_), .B0(mai_mai_n888_), .B1(mai_mai_n584_), .Y(mai_mai_n890_));
  OAI220     m868(.A0(mai_mai_n890_), .A1(mai_mai_n87_), .B0(mai_mai_n886_), .B1(mai_mai_n170_), .Y(mai_mai_n891_));
  NO2        m869(.A(mai_mai_n891_), .B(mai_mai_n495_), .Y(mai_mai_n892_));
  NA4        m870(.A(mai_mai_n892_), .B(mai_mai_n885_), .C(mai_mai_n880_), .D(mai_mai_n877_), .Y(mai_mai_n893_));
  NO3        m871(.A(mai_mai_n893_), .B(mai_mai_n873_), .C(mai_mai_n846_), .Y(mai_mai_n894_));
  NO2        m872(.A(i_0_), .B(mai_mai_n688_), .Y(mai_mai_n895_));
  NA2        m873(.A(mai_mai_n74_), .B(mai_mai_n45_), .Y(mai_mai_n896_));
  INV        m874(.A(mai_mai_n896_), .Y(mai_mai_n897_));
  NO3        m875(.A(mai_mai_n109_), .B(i_5_), .C(mai_mai_n25_), .Y(mai_mai_n898_));
  AO220      m876(.A0(mai_mai_n898_), .A1(mai_mai_n897_), .B0(mai_mai_n895_), .B1(mai_mai_n172_), .Y(mai_mai_n899_));
  AOI210     m877(.A0(mai_mai_n757_), .A1(mai_mai_n649_), .B0(mai_mai_n863_), .Y(mai_mai_n900_));
  AOI210     m878(.A0(mai_mai_n899_), .A1(mai_mai_n326_), .B0(mai_mai_n900_), .Y(mai_mai_n901_));
  NA2        m879(.A(mai_mai_n698_), .B(mai_mai_n150_), .Y(mai_mai_n902_));
  INV        m880(.A(mai_mai_n902_), .Y(mai_mai_n903_));
  NA3        m881(.A(mai_mai_n903_), .B(mai_mai_n639_), .C(mai_mai_n74_), .Y(mai_mai_n904_));
  NA3        m882(.A(mai_mai_n797_), .B(i_2_), .C(mai_mai_n49_), .Y(mai_mai_n905_));
  NA2        m883(.A(mai_mai_n798_), .B(i_9_), .Y(mai_mai_n906_));
  NO2        m884(.A(mai_mai_n905_), .B(mai_mai_n906_), .Y(mai_mai_n907_));
  NA2        m885(.A(mai_mai_n234_), .B(mai_mai_n222_), .Y(mai_mai_n908_));
  AOI210     m886(.A0(mai_mai_n908_), .A1(mai_mai_n829_), .B0(mai_mai_n157_), .Y(mai_mai_n909_));
  NO2        m887(.A(mai_mai_n909_), .B(mai_mai_n907_), .Y(mai_mai_n910_));
  NA3        m888(.A(mai_mai_n910_), .B(mai_mai_n904_), .C(mai_mai_n901_), .Y(mai_mai_n911_));
  NA2        m889(.A(mai_mai_n875_), .B(mai_mai_n351_), .Y(mai_mai_n912_));
  AOI210     m890(.A0(mai_mai_n285_), .A1(mai_mai_n161_), .B0(mai_mai_n912_), .Y(mai_mai_n913_));
  NA3        m891(.A(mai_mai_n40_), .B(mai_mai_n28_), .C(mai_mai_n45_), .Y(mai_mai_n914_));
  NA2        m892(.A(mai_mai_n851_), .B(mai_mai_n465_), .Y(mai_mai_n915_));
  AOI210     m893(.A0(mai_mai_n914_), .A1(mai_mai_n161_), .B0(mai_mai_n915_), .Y(mai_mai_n916_));
  NO2        m894(.A(mai_mai_n916_), .B(mai_mai_n913_), .Y(mai_mai_n917_));
  NO3        m895(.A(mai_mai_n837_), .B(mai_mai_n814_), .C(mai_mai_n184_), .Y(mai_mai_n918_));
  AOI220     m896(.A0(mai_mai_n918_), .A1(i_11_), .B0(mai_mai_n537_), .B1(mai_mai_n76_), .Y(mai_mai_n919_));
  NO3        m897(.A(mai_mai_n201_), .B(mai_mai_n362_), .C(i_0_), .Y(mai_mai_n920_));
  OAI210     m898(.A0(mai_mai_n920_), .A1(mai_mai_n77_), .B0(i_13_), .Y(mai_mai_n921_));
  NA3        m899(.A(mai_mai_n921_), .B(mai_mai_n919_), .C(mai_mai_n917_), .Y(mai_mai_n922_));
  AOI220     m900(.A0(mai_mai_n865_), .A1(mai_mai_n465_), .B0(mai_mai_n797_), .B1(mai_mai_n162_), .Y(mai_mai_n923_));
  NA2        m901(.A(mai_mai_n329_), .B(mai_mai_n174_), .Y(mai_mai_n924_));
  OR2        m902(.A(mai_mai_n924_), .B(mai_mai_n923_), .Y(mai_mai_n925_));
  AOI210     m903(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n173_), .Y(mai_mai_n926_));
  NA2        m904(.A(mai_mai_n926_), .B(mai_mai_n879_), .Y(mai_mai_n927_));
  NA3        m905(.A(mai_mai_n576_), .B(mai_mai_n181_), .C(mai_mai_n85_), .Y(mai_mai_n928_));
  NA2        m906(.A(mai_mai_n928_), .B(mai_mai_n511_), .Y(mai_mai_n929_));
  INV        m907(.A(mai_mai_n929_), .Y(mai_mai_n930_));
  NA3        m908(.A(mai_mai_n369_), .B(mai_mai_n169_), .C(mai_mai_n168_), .Y(mai_mai_n931_));
  NA3        m909(.A(mai_mai_n851_), .B(mai_mai_n274_), .C(mai_mai_n222_), .Y(mai_mai_n932_));
  NA2        m910(.A(mai_mai_n932_), .B(mai_mai_n931_), .Y(mai_mai_n933_));
  NA3        m911(.A(mai_mai_n369_), .B(mai_mai_n317_), .C(mai_mai_n213_), .Y(mai_mai_n934_));
  INV        m912(.A(mai_mai_n934_), .Y(mai_mai_n935_));
  NOi31      m913(.An(mai_mai_n368_), .B(mai_mai_n896_), .C(mai_mai_n231_), .Y(mai_mai_n936_));
  NO3        m914(.A(mai_mai_n848_), .B(mai_mai_n209_), .C(mai_mai_n184_), .Y(mai_mai_n937_));
  NO4        m915(.A(mai_mai_n937_), .B(mai_mai_n936_), .C(mai_mai_n935_), .D(mai_mai_n933_), .Y(mai_mai_n938_));
  NA4        m916(.A(mai_mai_n938_), .B(mai_mai_n930_), .C(mai_mai_n927_), .D(mai_mai_n925_), .Y(mai_mai_n939_));
  INV        m917(.A(mai_mai_n578_), .Y(mai_mai_n940_));
  NO3        m918(.A(mai_mai_n940_), .B(mai_mai_n527_), .C(mai_mai_n323_), .Y(mai_mai_n941_));
  NO2        m919(.A(mai_mai_n87_), .B(i_5_), .Y(mai_mai_n942_));
  NA3        m920(.A(mai_mai_n798_), .B(mai_mai_n113_), .C(mai_mai_n128_), .Y(mai_mai_n943_));
  INV        m921(.A(mai_mai_n943_), .Y(mai_mai_n944_));
  AOI210     m922(.A0(mai_mai_n944_), .A1(mai_mai_n942_), .B0(mai_mai_n941_), .Y(mai_mai_n945_));
  NA3        m923(.A(mai_mai_n289_), .B(i_5_), .C(mai_mai_n187_), .Y(mai_mai_n946_));
  NAi31      m924(.An(mai_mai_n232_), .B(mai_mai_n946_), .C(mai_mai_n233_), .Y(mai_mai_n947_));
  NO4        m925(.A(mai_mai_n231_), .B(mai_mai_n201_), .C(i_0_), .D(i_12_), .Y(mai_mai_n948_));
  AOI220     m926(.A0(mai_mai_n948_), .A1(mai_mai_n947_), .B0(mai_mai_n752_), .B1(mai_mai_n174_), .Y(mai_mai_n949_));
  AN2        m927(.A(mai_mai_n837_), .B(mai_mai_n157_), .Y(mai_mai_n950_));
  NO4        m928(.A(mai_mai_n950_), .B(i_12_), .C(mai_mai_n612_), .D(mai_mai_n135_), .Y(mai_mai_n951_));
  NA2        m929(.A(mai_mai_n951_), .B(mai_mai_n209_), .Y(mai_mai_n952_));
  NA2        m930(.A(mai_mai_n865_), .B(mai_mai_n449_), .Y(mai_mai_n953_));
  NA2        m931(.A(mai_mai_n65_), .B(mai_mai_n105_), .Y(mai_mai_n954_));
  OAI220     m932(.A0(mai_mai_n954_), .A1(mai_mai_n946_), .B0(mai_mai_n953_), .B1(mai_mai_n640_), .Y(mai_mai_n955_));
  NA2        m933(.A(mai_mai_n955_), .B(mai_mai_n855_), .Y(mai_mai_n956_));
  NA4        m934(.A(mai_mai_n956_), .B(mai_mai_n952_), .C(mai_mai_n949_), .D(mai_mai_n945_), .Y(mai_mai_n957_));
  NO4        m935(.A(mai_mai_n957_), .B(mai_mai_n939_), .C(mai_mai_n922_), .D(mai_mai_n911_), .Y(mai_mai_n958_));
  OAI210     m936(.A0(mai_mai_n776_), .A1(mai_mai_n770_), .B0(mai_mai_n37_), .Y(mai_mai_n959_));
  NA2        m937(.A(mai_mai_n959_), .B(mai_mai_n574_), .Y(mai_mai_n960_));
  NA2        m938(.A(mai_mai_n960_), .B(mai_mai_n197_), .Y(mai_mai_n961_));
  OAI210     m939(.A0(mai_mai_n578_), .A1(mai_mai_n576_), .B0(mai_mai_n301_), .Y(mai_mai_n962_));
  NAi31      m940(.An(i_7_), .B(i_2_), .C(i_10_), .Y(mai_mai_n963_));
  AOI210     m941(.A0(mai_mai_n121_), .A1(mai_mai_n71_), .B0(mai_mai_n963_), .Y(mai_mai_n964_));
  NO2        m942(.A(mai_mai_n964_), .B(mai_mai_n609_), .Y(mai_mai_n965_));
  NA2        m943(.A(mai_mai_n965_), .B(mai_mai_n962_), .Y(mai_mai_n966_));
  NO2        m944(.A(mai_mai_n439_), .B(mai_mai_n258_), .Y(mai_mai_n967_));
  NO4        m945(.A(mai_mai_n225_), .B(mai_mai_n149_), .C(mai_mai_n643_), .D(mai_mai_n37_), .Y(mai_mai_n968_));
  NO3        m946(.A(mai_mai_n968_), .B(mai_mai_n967_), .C(mai_mai_n830_), .Y(mai_mai_n969_));
  INV        m947(.A(mai_mai_n969_), .Y(mai_mai_n970_));
  AOI210     m948(.A0(mai_mai_n966_), .A1(mai_mai_n49_), .B0(mai_mai_n970_), .Y(mai_mai_n971_));
  AOI210     m949(.A0(mai_mai_n971_), .A1(mai_mai_n961_), .B0(mai_mai_n74_), .Y(mai_mai_n972_));
  NO2        m950(.A(mai_mai_n534_), .B(mai_mai_n358_), .Y(mai_mai_n973_));
  NO2        m951(.A(mai_mai_n973_), .B(mai_mai_n717_), .Y(mai_mai_n974_));
  AOI210     m952(.A0(mai_mai_n926_), .A1(mai_mai_n851_), .B0(mai_mai_n866_), .Y(mai_mai_n975_));
  NO2        m953(.A(mai_mai_n975_), .B(mai_mai_n643_), .Y(mai_mai_n976_));
  NA2        m954(.A(mai_mai_n253_), .B(mai_mai_n58_), .Y(mai_mai_n977_));
  AOI220     m955(.A0(mai_mai_n977_), .A1(mai_mai_n77_), .B0(mai_mai_n324_), .B1(mai_mai_n246_), .Y(mai_mai_n978_));
  NO2        m956(.A(mai_mai_n978_), .B(mai_mai_n228_), .Y(mai_mai_n979_));
  NA3        m957(.A(mai_mai_n100_), .B(mai_mai_n291_), .C(mai_mai_n31_), .Y(mai_mai_n980_));
  INV        m958(.A(mai_mai_n980_), .Y(mai_mai_n981_));
  NO3        m959(.A(mai_mai_n981_), .B(mai_mai_n979_), .C(mai_mai_n976_), .Y(mai_mai_n982_));
  NA3        m960(.A(mai_mai_n721_), .B(mai_mai_n274_), .C(mai_mai_n81_), .Y(mai_mai_n983_));
  NO2        m961(.A(mai_mai_n983_), .B(i_11_), .Y(mai_mai_n984_));
  INV        m962(.A(mai_mai_n531_), .Y(mai_mai_n985_));
  INV        m963(.A(mai_mai_n339_), .Y(mai_mai_n986_));
  AOI210     m964(.A0(mai_mai_n986_), .A1(mai_mai_n985_), .B0(mai_mai_n41_), .Y(mai_mai_n987_));
  NO2        m965(.A(mai_mai_n987_), .B(mai_mai_n984_), .Y(mai_mai_n988_));
  OAI210     m966(.A0(mai_mai_n982_), .A1(i_4_), .B0(mai_mai_n988_), .Y(mai_mai_n989_));
  NO3        m967(.A(mai_mai_n989_), .B(mai_mai_n974_), .C(mai_mai_n972_), .Y(mai_mai_n990_));
  NA4        m968(.A(mai_mai_n990_), .B(mai_mai_n958_), .C(mai_mai_n894_), .D(mai_mai_n822_), .Y(mai4));
  NAi21      u0000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u0001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u0002(.A(i_9_), .Y(men_men_n25_));
  INV        u0003(.A(i_3_), .Y(men_men_n26_));
  NO2        u0004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u0005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u0006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u0007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u0008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u0010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u0011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u0012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u0013(.A(i_4_), .Y(men_men_n36_));
  INV        u0014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u0015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NO3        u0016(.A(men_men_n38_), .B(i_12_), .C(men_men_n37_), .Y(men_men_n39_));
  NOi21      u0017(.An(i_12_), .B(i_13_), .Y(men_men_n40_));
  INV        u0018(.A(men_men_n40_), .Y(men_men_n41_));
  NO2        u0019(.A(men_men_n36_), .B(i_3_), .Y(men_men_n42_));
  NAi31      u0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n43_));
  INV        u0021(.A(men_men_n35_), .Y(men1));
  INV        u0022(.A(i_11_), .Y(men_men_n45_));
  NO2        u0023(.A(men_men_n45_), .B(i_6_), .Y(men_men_n46_));
  INV        u0024(.A(i_2_), .Y(men_men_n47_));
  NA2        u0025(.A(i_0_), .B(i_3_), .Y(men_men_n48_));
  INV        u0026(.A(i_5_), .Y(men_men_n49_));
  NO2        u0027(.A(i_7_), .B(i_10_), .Y(men_men_n50_));
  AOI210     u0028(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n50_), .Y(men_men_n51_));
  OAI210     u0029(.A0(men_men_n51_), .A1(i_3_), .B0(men_men_n49_), .Y(men_men_n52_));
  AOI210     u0030(.A0(men_men_n52_), .A1(men_men_n48_), .B0(men_men_n47_), .Y(men_men_n53_));
  NA2        u0031(.A(i_0_), .B(i_2_), .Y(men_men_n54_));
  NA2        u0032(.A(i_7_), .B(i_9_), .Y(men_men_n55_));
  NA2        u0033(.A(men_men_n53_), .B(men_men_n46_), .Y(men_men_n56_));
  NA3        u0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n57_));
  NO2        u0035(.A(i_1_), .B(i_6_), .Y(men_men_n58_));
  NA2        u0036(.A(i_8_), .B(i_7_), .Y(men_men_n59_));
  OAI210     u0037(.A0(men_men_n59_), .A1(men_men_n58_), .B0(men_men_n57_), .Y(men_men_n60_));
  NA2        u0038(.A(men_men_n60_), .B(i_12_), .Y(men_men_n61_));
  NAi21      u0039(.An(i_2_), .B(i_7_), .Y(men_men_n62_));
  INV        u0040(.A(i_1_), .Y(men_men_n63_));
  NA2        u0041(.A(men_men_n63_), .B(i_6_), .Y(men_men_n64_));
  NA3        u0042(.A(men_men_n64_), .B(men_men_n62_), .C(men_men_n31_), .Y(men_men_n65_));
  NA2        u0043(.A(i_1_), .B(i_10_), .Y(men_men_n66_));
  NO2        u0044(.A(men_men_n66_), .B(i_6_), .Y(men_men_n67_));
  NAi31      u0045(.An(men_men_n67_), .B(men_men_n65_), .C(men_men_n61_), .Y(men_men_n68_));
  NA2        u0046(.A(men_men_n51_), .B(i_2_), .Y(men_men_n69_));
  AOI210     u0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n70_));
  NA2        u0048(.A(i_1_), .B(i_6_), .Y(men_men_n71_));
  NO2        u0049(.A(men_men_n71_), .B(men_men_n25_), .Y(men_men_n72_));
  INV        u0050(.A(i_0_), .Y(men_men_n73_));
  NAi21      u0051(.An(i_5_), .B(i_10_), .Y(men_men_n74_));
  NA2        u0052(.A(i_5_), .B(i_9_), .Y(men_men_n75_));
  AOI210     u0053(.A0(men_men_n75_), .A1(men_men_n74_), .B0(men_men_n73_), .Y(men_men_n76_));
  NO2        u0054(.A(men_men_n76_), .B(men_men_n72_), .Y(men_men_n77_));
  OAI210     u0055(.A0(men_men_n70_), .A1(men_men_n69_), .B0(men_men_n77_), .Y(men_men_n78_));
  OAI210     u0056(.A0(men_men_n78_), .A1(men_men_n68_), .B0(i_0_), .Y(men_men_n79_));
  NA2        u0057(.A(i_12_), .B(i_5_), .Y(men_men_n80_));
  NA2        u0058(.A(i_2_), .B(i_8_), .Y(men_men_n81_));
  NO2        u0059(.A(men_men_n81_), .B(men_men_n58_), .Y(men_men_n82_));
  NO2        u0060(.A(i_3_), .B(i_9_), .Y(men_men_n83_));
  NO2        u0061(.A(i_3_), .B(i_7_), .Y(men_men_n84_));
  NO3        u0062(.A(men_men_n84_), .B(men_men_n83_), .C(men_men_n63_), .Y(men_men_n85_));
  INV        u0063(.A(i_6_), .Y(men_men_n86_));
  OR4        u0064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n87_));
  INV        u0065(.A(men_men_n87_), .Y(men_men_n88_));
  NO2        u0066(.A(i_2_), .B(i_7_), .Y(men_men_n89_));
  NO2        u0067(.A(men_men_n88_), .B(men_men_n89_), .Y(men_men_n90_));
  OAI210     u0068(.A0(men_men_n85_), .A1(men_men_n82_), .B0(men_men_n90_), .Y(men_men_n91_));
  NAi21      u0069(.An(i_6_), .B(i_10_), .Y(men_men_n92_));
  NA2        u0070(.A(i_6_), .B(i_9_), .Y(men_men_n93_));
  AOI210     u0071(.A0(men_men_n93_), .A1(men_men_n92_), .B0(men_men_n63_), .Y(men_men_n94_));
  NA2        u0072(.A(i_2_), .B(i_6_), .Y(men_men_n95_));
  INV        u0073(.A(men_men_n94_), .Y(men_men_n96_));
  AOI210     u0074(.A0(men_men_n96_), .A1(men_men_n91_), .B0(men_men_n80_), .Y(men_men_n97_));
  AN3        u0075(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n98_));
  NAi21      u0076(.An(i_6_), .B(i_11_), .Y(men_men_n99_));
  NO2        u0077(.A(i_5_), .B(i_8_), .Y(men_men_n100_));
  NOi21      u0078(.An(men_men_n100_), .B(men_men_n99_), .Y(men_men_n101_));
  AOI220     u0079(.A0(men_men_n101_), .A1(men_men_n62_), .B0(men_men_n98_), .B1(men_men_n32_), .Y(men_men_n102_));
  INV        u0080(.A(i_7_), .Y(men_men_n103_));
  NA2        u0081(.A(men_men_n47_), .B(men_men_n103_), .Y(men_men_n104_));
  NO2        u0082(.A(i_0_), .B(i_5_), .Y(men_men_n105_));
  NO2        u0083(.A(men_men_n105_), .B(men_men_n86_), .Y(men_men_n106_));
  NA2        u0084(.A(i_12_), .B(i_3_), .Y(men_men_n107_));
  INV        u0085(.A(men_men_n107_), .Y(men_men_n108_));
  NA3        u0086(.A(men_men_n108_), .B(men_men_n106_), .C(men_men_n104_), .Y(men_men_n109_));
  NAi21      u0087(.An(i_7_), .B(i_11_), .Y(men_men_n110_));
  NO3        u0088(.A(men_men_n110_), .B(men_men_n92_), .C(men_men_n54_), .Y(men_men_n111_));
  AN2        u0089(.A(i_2_), .B(i_10_), .Y(men_men_n112_));
  NO2        u0090(.A(men_men_n112_), .B(i_7_), .Y(men_men_n113_));
  OR2        u0091(.A(men_men_n80_), .B(men_men_n58_), .Y(men_men_n114_));
  NO2        u0092(.A(i_8_), .B(men_men_n103_), .Y(men_men_n115_));
  NO3        u0093(.A(men_men_n115_), .B(men_men_n114_), .C(men_men_n113_), .Y(men_men_n116_));
  NA2        u0094(.A(i_12_), .B(i_7_), .Y(men_men_n117_));
  NO2        u0095(.A(men_men_n63_), .B(men_men_n26_), .Y(men_men_n118_));
  NA2        u0096(.A(i_11_), .B(i_12_), .Y(men_men_n119_));
  NO2        u0097(.A(men_men_n1043_), .B(men_men_n116_), .Y(men_men_n120_));
  NAi41      u0098(.An(men_men_n111_), .B(men_men_n120_), .C(men_men_n109_), .D(men_men_n102_), .Y(men_men_n121_));
  NOi21      u0099(.An(i_1_), .B(i_5_), .Y(men_men_n122_));
  NA2        u0100(.A(men_men_n122_), .B(i_11_), .Y(men_men_n123_));
  NA2        u0101(.A(men_men_n103_), .B(men_men_n37_), .Y(men_men_n124_));
  NA2        u0102(.A(i_7_), .B(men_men_n25_), .Y(men_men_n125_));
  NA2        u0103(.A(men_men_n125_), .B(men_men_n124_), .Y(men_men_n126_));
  NO2        u0104(.A(men_men_n126_), .B(men_men_n47_), .Y(men_men_n127_));
  NA2        u0105(.A(men_men_n93_), .B(men_men_n92_), .Y(men_men_n128_));
  NAi21      u0106(.An(i_3_), .B(i_8_), .Y(men_men_n129_));
  NA2        u0107(.A(men_men_n129_), .B(men_men_n62_), .Y(men_men_n130_));
  NOi31      u0108(.An(men_men_n130_), .B(men_men_n128_), .C(men_men_n127_), .Y(men_men_n131_));
  NO2        u0109(.A(i_1_), .B(men_men_n86_), .Y(men_men_n132_));
  NO2        u0110(.A(i_6_), .B(i_5_), .Y(men_men_n133_));
  NA2        u0111(.A(men_men_n133_), .B(i_3_), .Y(men_men_n134_));
  AO210      u0112(.A0(men_men_n134_), .A1(men_men_n48_), .B0(men_men_n132_), .Y(men_men_n135_));
  OAI220     u0113(.A0(men_men_n135_), .A1(men_men_n110_), .B0(men_men_n131_), .B1(men_men_n123_), .Y(men_men_n136_));
  NO3        u0114(.A(men_men_n136_), .B(men_men_n121_), .C(men_men_n97_), .Y(men_men_n137_));
  NA3        u0115(.A(men_men_n137_), .B(men_men_n79_), .C(men_men_n56_), .Y(men2));
  NO2        u0116(.A(men_men_n63_), .B(men_men_n37_), .Y(men_men_n139_));
  NA2        u0117(.A(i_6_), .B(men_men_n25_), .Y(men_men_n140_));
  NA2        u0118(.A(men_men_n140_), .B(men_men_n139_), .Y(men_men_n141_));
  NA4        u0119(.A(men_men_n141_), .B(men_men_n77_), .C(men_men_n69_), .D(men_men_n30_), .Y(men0));
  AN2        u0120(.A(i_8_), .B(i_7_), .Y(men_men_n143_));
  NA2        u0121(.A(men_men_n143_), .B(i_6_), .Y(men_men_n144_));
  NO2        u0122(.A(i_12_), .B(i_13_), .Y(men_men_n145_));
  NAi21      u0123(.An(i_5_), .B(i_11_), .Y(men_men_n146_));
  NOi21      u0124(.An(men_men_n145_), .B(men_men_n146_), .Y(men_men_n147_));
  NO2        u0125(.A(i_0_), .B(i_1_), .Y(men_men_n148_));
  NA2        u0126(.A(i_2_), .B(i_3_), .Y(men_men_n149_));
  NO2        u0127(.A(men_men_n149_), .B(i_4_), .Y(men_men_n150_));
  NA3        u0128(.A(men_men_n150_), .B(men_men_n148_), .C(men_men_n147_), .Y(men_men_n151_));
  AN2        u0129(.A(men_men_n145_), .B(men_men_n83_), .Y(men_men_n152_));
  NO2        u0130(.A(men_men_n152_), .B(men_men_n27_), .Y(men_men_n153_));
  NA2        u0131(.A(i_1_), .B(i_5_), .Y(men_men_n154_));
  NO2        u0132(.A(men_men_n73_), .B(men_men_n47_), .Y(men_men_n155_));
  NA2        u0133(.A(men_men_n155_), .B(men_men_n36_), .Y(men_men_n156_));
  NO3        u0134(.A(men_men_n156_), .B(men_men_n154_), .C(men_men_n153_), .Y(men_men_n157_));
  OR2        u0135(.A(i_0_), .B(i_1_), .Y(men_men_n158_));
  NO3        u0136(.A(men_men_n158_), .B(men_men_n80_), .C(i_13_), .Y(men_men_n159_));
  NAi32      u0137(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n160_));
  NAi21      u0138(.An(men_men_n160_), .B(men_men_n159_), .Y(men_men_n161_));
  NOi21      u0139(.An(i_4_), .B(i_10_), .Y(men_men_n162_));
  NA2        u0140(.A(men_men_n162_), .B(men_men_n40_), .Y(men_men_n163_));
  NO2        u0141(.A(i_3_), .B(i_5_), .Y(men_men_n164_));
  NO3        u0142(.A(men_men_n73_), .B(i_2_), .C(i_1_), .Y(men_men_n165_));
  NA2        u0143(.A(men_men_n165_), .B(men_men_n164_), .Y(men_men_n166_));
  OAI210     u0144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n161_), .Y(men_men_n167_));
  NO2        u0145(.A(men_men_n167_), .B(men_men_n157_), .Y(men_men_n168_));
  AOI210     u0146(.A0(men_men_n168_), .A1(men_men_n151_), .B0(men_men_n144_), .Y(men_men_n169_));
  NA3        u0147(.A(men_men_n73_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n170_));
  NA2        u0148(.A(i_3_), .B(men_men_n49_), .Y(men_men_n171_));
  NOi21      u0149(.An(i_4_), .B(i_9_), .Y(men_men_n172_));
  NOi21      u0150(.An(i_11_), .B(i_13_), .Y(men_men_n173_));
  NA2        u0151(.A(men_men_n173_), .B(men_men_n172_), .Y(men_men_n174_));
  NO2        u0152(.A(i_4_), .B(i_5_), .Y(men_men_n175_));
  NAi21      u0153(.An(i_12_), .B(i_11_), .Y(men_men_n176_));
  NO2        u0154(.A(men_men_n176_), .B(i_13_), .Y(men_men_n177_));
  NA3        u0155(.A(men_men_n177_), .B(men_men_n175_), .C(men_men_n83_), .Y(men_men_n178_));
  AOI210     u0156(.A0(men_men_n178_), .A1(men_men_n174_), .B0(men_men_n170_), .Y(men_men_n179_));
  NO2        u0157(.A(men_men_n73_), .B(men_men_n63_), .Y(men_men_n180_));
  NA2        u0158(.A(men_men_n180_), .B(men_men_n47_), .Y(men_men_n181_));
  NA2        u0159(.A(men_men_n36_), .B(i_5_), .Y(men_men_n182_));
  NAi31      u0160(.An(men_men_n182_), .B(men_men_n152_), .C(i_11_), .Y(men_men_n183_));
  NA2        u0161(.A(i_3_), .B(i_5_), .Y(men_men_n184_));
  OR2        u0162(.A(men_men_n184_), .B(men_men_n174_), .Y(men_men_n185_));
  AOI210     u0163(.A0(men_men_n185_), .A1(men_men_n183_), .B0(men_men_n181_), .Y(men_men_n186_));
  NO2        u0164(.A(men_men_n73_), .B(i_5_), .Y(men_men_n187_));
  NO2        u0165(.A(i_13_), .B(i_10_), .Y(men_men_n188_));
  NA3        u0166(.A(men_men_n188_), .B(men_men_n187_), .C(men_men_n45_), .Y(men_men_n189_));
  NO2        u0167(.A(i_2_), .B(i_1_), .Y(men_men_n190_));
  NA2        u0168(.A(men_men_n190_), .B(i_3_), .Y(men_men_n191_));
  NAi21      u0169(.An(i_4_), .B(i_12_), .Y(men_men_n192_));
  NO4        u0170(.A(men_men_n192_), .B(men_men_n191_), .C(men_men_n189_), .D(men_men_n25_), .Y(men_men_n193_));
  NO3        u0171(.A(men_men_n193_), .B(men_men_n186_), .C(men_men_n179_), .Y(men_men_n194_));
  INV        u0172(.A(i_8_), .Y(men_men_n195_));
  NO2        u0173(.A(men_men_n195_), .B(i_7_), .Y(men_men_n196_));
  NA2        u0174(.A(men_men_n196_), .B(i_6_), .Y(men_men_n197_));
  NO3        u0175(.A(i_3_), .B(men_men_n86_), .C(men_men_n49_), .Y(men_men_n198_));
  NA2        u0176(.A(men_men_n198_), .B(men_men_n115_), .Y(men_men_n199_));
  NO3        u0177(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n200_));
  NA3        u0178(.A(men_men_n200_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n201_));
  NO3        u0179(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n202_));
  OAI210     u0180(.A0(men_men_n98_), .A1(i_12_), .B0(men_men_n202_), .Y(men_men_n203_));
  AOI210     u0181(.A0(men_men_n203_), .A1(men_men_n201_), .B0(men_men_n199_), .Y(men_men_n204_));
  NO2        u0182(.A(i_3_), .B(i_8_), .Y(men_men_n205_));
  NO3        u0183(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n206_));
  NO2        u0184(.A(men_men_n105_), .B(men_men_n58_), .Y(men_men_n207_));
  NO2        u0185(.A(i_13_), .B(i_9_), .Y(men_men_n208_));
  NA3        u0186(.A(men_men_n208_), .B(i_6_), .C(men_men_n195_), .Y(men_men_n209_));
  NAi21      u0187(.An(i_12_), .B(i_3_), .Y(men_men_n210_));
  NO2        u0188(.A(men_men_n45_), .B(i_5_), .Y(men_men_n211_));
  NO3        u0189(.A(i_0_), .B(i_2_), .C(men_men_n63_), .Y(men_men_n212_));
  NA3        u0190(.A(men_men_n212_), .B(men_men_n211_), .C(i_10_), .Y(men_men_n213_));
  NO2        u0191(.A(men_men_n213_), .B(men_men_n209_), .Y(men_men_n214_));
  AOI210     u0192(.A0(men_men_n214_), .A1(i_7_), .B0(men_men_n204_), .Y(men_men_n215_));
  OAI220     u0193(.A0(men_men_n215_), .A1(i_4_), .B0(men_men_n197_), .B1(men_men_n194_), .Y(men_men_n216_));
  NAi21      u0194(.An(i_12_), .B(i_7_), .Y(men_men_n217_));
  NA3        u0195(.A(i_13_), .B(men_men_n195_), .C(i_10_), .Y(men_men_n218_));
  NA2        u0196(.A(i_0_), .B(i_5_), .Y(men_men_n219_));
  NAi31      u0197(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n220_));
  NO2        u0198(.A(men_men_n36_), .B(i_13_), .Y(men_men_n221_));
  NO2        u0199(.A(men_men_n73_), .B(men_men_n26_), .Y(men_men_n222_));
  NO2        u0200(.A(men_men_n47_), .B(men_men_n63_), .Y(men_men_n223_));
  NA3        u0201(.A(men_men_n223_), .B(men_men_n222_), .C(men_men_n221_), .Y(men_men_n224_));
  INV        u0202(.A(i_13_), .Y(men_men_n225_));
  NO2        u0203(.A(i_12_), .B(men_men_n225_), .Y(men_men_n226_));
  NA3        u0204(.A(men_men_n226_), .B(men_men_n200_), .C(men_men_n198_), .Y(men_men_n227_));
  OAI210     u0205(.A0(men_men_n224_), .A1(men_men_n220_), .B0(men_men_n227_), .Y(men_men_n228_));
  NA2        u0206(.A(men_men_n228_), .B(men_men_n143_), .Y(men_men_n229_));
  NO2        u0207(.A(i_12_), .B(men_men_n37_), .Y(men_men_n230_));
  NO2        u0208(.A(men_men_n184_), .B(i_4_), .Y(men_men_n231_));
  NA2        u0209(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n232_));
  OR2        u0210(.A(i_8_), .B(i_7_), .Y(men_men_n233_));
  NO2        u0211(.A(men_men_n233_), .B(men_men_n86_), .Y(men_men_n234_));
  NO2        u0212(.A(men_men_n54_), .B(i_1_), .Y(men_men_n235_));
  NA2        u0213(.A(men_men_n235_), .B(men_men_n234_), .Y(men_men_n236_));
  INV        u0214(.A(i_12_), .Y(men_men_n237_));
  NO2        u0215(.A(men_men_n45_), .B(men_men_n237_), .Y(men_men_n238_));
  NO3        u0216(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n239_));
  NA2        u0217(.A(i_2_), .B(i_1_), .Y(men_men_n240_));
  NO2        u0218(.A(men_men_n236_), .B(men_men_n232_), .Y(men_men_n241_));
  NO3        u0219(.A(i_11_), .B(i_7_), .C(men_men_n37_), .Y(men_men_n242_));
  NAi21      u0220(.An(i_4_), .B(i_3_), .Y(men_men_n243_));
  NO2        u0221(.A(i_0_), .B(i_6_), .Y(men_men_n244_));
  NOi41      u0222(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n245_));
  NA2        u0223(.A(men_men_n245_), .B(men_men_n244_), .Y(men_men_n246_));
  NO2        u0224(.A(men_men_n240_), .B(men_men_n184_), .Y(men_men_n247_));
  NAi21      u0225(.An(men_men_n246_), .B(men_men_n247_), .Y(men_men_n248_));
  INV        u0226(.A(men_men_n248_), .Y(men_men_n249_));
  AOI220     u0227(.A0(men_men_n249_), .A1(men_men_n40_), .B0(men_men_n241_), .B1(men_men_n208_), .Y(men_men_n250_));
  NO2        u0228(.A(i_11_), .B(men_men_n225_), .Y(men_men_n251_));
  NOi21      u0229(.An(i_1_), .B(i_6_), .Y(men_men_n252_));
  NAi21      u0230(.An(i_3_), .B(i_7_), .Y(men_men_n253_));
  NA2        u0231(.A(men_men_n237_), .B(i_9_), .Y(men_men_n254_));
  OR4        u0232(.A(men_men_n254_), .B(men_men_n253_), .C(men_men_n252_), .D(men_men_n187_), .Y(men_men_n255_));
  NO2        u0233(.A(men_men_n49_), .B(men_men_n25_), .Y(men_men_n256_));
  NO2        u0234(.A(i_12_), .B(i_3_), .Y(men_men_n257_));
  NA2        u0235(.A(men_men_n73_), .B(i_5_), .Y(men_men_n258_));
  NA2        u0236(.A(i_3_), .B(i_9_), .Y(men_men_n259_));
  NAi21      u0237(.An(i_7_), .B(i_10_), .Y(men_men_n260_));
  NO2        u0238(.A(men_men_n260_), .B(men_men_n259_), .Y(men_men_n261_));
  INV        u0239(.A(men_men_n255_), .Y(men_men_n262_));
  NA3        u0240(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n263_));
  INV        u0241(.A(men_men_n144_), .Y(men_men_n264_));
  NA2        u0242(.A(men_men_n237_), .B(i_13_), .Y(men_men_n265_));
  NO2        u0243(.A(men_men_n265_), .B(men_men_n75_), .Y(men_men_n266_));
  AOI220     u0244(.A0(men_men_n266_), .A1(men_men_n264_), .B0(men_men_n262_), .B1(men_men_n251_), .Y(men_men_n267_));
  NO2        u0245(.A(men_men_n233_), .B(men_men_n37_), .Y(men_men_n268_));
  NA2        u0246(.A(i_12_), .B(i_6_), .Y(men_men_n269_));
  OR2        u0247(.A(i_13_), .B(i_9_), .Y(men_men_n270_));
  NO3        u0248(.A(men_men_n270_), .B(men_men_n269_), .C(men_men_n49_), .Y(men_men_n271_));
  NO2        u0249(.A(men_men_n243_), .B(i_2_), .Y(men_men_n272_));
  NA3        u0250(.A(men_men_n272_), .B(men_men_n271_), .C(men_men_n45_), .Y(men_men_n273_));
  NA2        u0251(.A(men_men_n251_), .B(i_9_), .Y(men_men_n274_));
  NA2        u0252(.A(men_men_n258_), .B(men_men_n64_), .Y(men_men_n275_));
  OAI210     u0253(.A0(men_men_n275_), .A1(men_men_n274_), .B0(men_men_n273_), .Y(men_men_n276_));
  NA2        u0254(.A(men_men_n155_), .B(men_men_n63_), .Y(men_men_n277_));
  NO3        u0255(.A(i_11_), .B(men_men_n225_), .C(men_men_n25_), .Y(men_men_n278_));
  NO2        u0256(.A(men_men_n253_), .B(i_8_), .Y(men_men_n279_));
  NO2        u0257(.A(i_6_), .B(men_men_n49_), .Y(men_men_n280_));
  NA3        u0258(.A(men_men_n280_), .B(men_men_n279_), .C(men_men_n278_), .Y(men_men_n281_));
  NO3        u0259(.A(men_men_n26_), .B(men_men_n86_), .C(i_5_), .Y(men_men_n282_));
  NA3        u0260(.A(men_men_n282_), .B(men_men_n268_), .C(men_men_n226_), .Y(men_men_n283_));
  AOI210     u0261(.A0(men_men_n283_), .A1(men_men_n281_), .B0(men_men_n277_), .Y(men_men_n284_));
  AOI210     u0262(.A0(men_men_n276_), .A1(men_men_n268_), .B0(men_men_n284_), .Y(men_men_n285_));
  NA4        u0263(.A(men_men_n285_), .B(men_men_n267_), .C(men_men_n250_), .D(men_men_n229_), .Y(men_men_n286_));
  NO3        u0264(.A(i_12_), .B(men_men_n225_), .C(men_men_n37_), .Y(men_men_n287_));
  INV        u0265(.A(men_men_n287_), .Y(men_men_n288_));
  NA2        u0266(.A(i_8_), .B(men_men_n103_), .Y(men_men_n289_));
  NO3        u0267(.A(i_0_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n290_));
  NO2        u0268(.A(men_men_n240_), .B(i_0_), .Y(men_men_n291_));
  NA2        u0269(.A(i_0_), .B(i_1_), .Y(men_men_n292_));
  NO2        u0270(.A(men_men_n292_), .B(i_2_), .Y(men_men_n293_));
  NO2        u0271(.A(men_men_n59_), .B(i_6_), .Y(men_men_n294_));
  NA3        u0272(.A(men_men_n294_), .B(men_men_n293_), .C(men_men_n164_), .Y(men_men_n295_));
  NO2        u0273(.A(i_3_), .B(i_10_), .Y(men_men_n296_));
  NA3        u0274(.A(men_men_n296_), .B(men_men_n40_), .C(men_men_n45_), .Y(men_men_n297_));
  NO2        u0275(.A(i_2_), .B(men_men_n103_), .Y(men_men_n298_));
  NA2        u0276(.A(i_1_), .B(men_men_n36_), .Y(men_men_n299_));
  NO2        u0277(.A(men_men_n299_), .B(i_8_), .Y(men_men_n300_));
  NA2        u0278(.A(men_men_n300_), .B(men_men_n298_), .Y(men_men_n301_));
  AN2        u0279(.A(i_3_), .B(i_10_), .Y(men_men_n302_));
  NA4        u0280(.A(men_men_n302_), .B(men_men_n200_), .C(men_men_n177_), .D(men_men_n175_), .Y(men_men_n303_));
  NO2        u0281(.A(i_5_), .B(men_men_n37_), .Y(men_men_n304_));
  NO2        u0282(.A(men_men_n47_), .B(men_men_n26_), .Y(men_men_n305_));
  OR2        u0283(.A(men_men_n301_), .B(men_men_n297_), .Y(men_men_n306_));
  OAI220     u0284(.A0(men_men_n306_), .A1(i_6_), .B0(men_men_n295_), .B1(men_men_n288_), .Y(men_men_n307_));
  NO4        u0285(.A(men_men_n307_), .B(men_men_n286_), .C(men_men_n216_), .D(men_men_n169_), .Y(men_men_n308_));
  NO3        u0286(.A(men_men_n45_), .B(i_13_), .C(i_9_), .Y(men_men_n309_));
  NO2        u0287(.A(men_men_n59_), .B(men_men_n86_), .Y(men_men_n310_));
  NA2        u0288(.A(men_men_n291_), .B(men_men_n310_), .Y(men_men_n311_));
  NO3        u0289(.A(i_6_), .B(men_men_n195_), .C(i_7_), .Y(men_men_n312_));
  NA2        u0290(.A(men_men_n312_), .B(men_men_n200_), .Y(men_men_n313_));
  AOI210     u0291(.A0(men_men_n313_), .A1(men_men_n311_), .B0(men_men_n171_), .Y(men_men_n314_));
  NO2        u0292(.A(i_2_), .B(i_3_), .Y(men_men_n315_));
  OR2        u0293(.A(i_0_), .B(i_5_), .Y(men_men_n316_));
  NA2        u0294(.A(men_men_n219_), .B(men_men_n316_), .Y(men_men_n317_));
  NO2        u0295(.A(i_8_), .B(i_6_), .Y(men_men_n318_));
  NO2        u0296(.A(men_men_n158_), .B(men_men_n47_), .Y(men_men_n319_));
  NA3        u0297(.A(men_men_n319_), .B(men_men_n318_), .C(men_men_n164_), .Y(men_men_n320_));
  INV        u0298(.A(men_men_n320_), .Y(men_men_n321_));
  OAI210     u0299(.A0(men_men_n321_), .A1(men_men_n314_), .B0(i_4_), .Y(men_men_n322_));
  NO2        u0300(.A(i_12_), .B(i_10_), .Y(men_men_n323_));
  NOi21      u0301(.An(i_5_), .B(i_0_), .Y(men_men_n324_));
  NO3        u0302(.A(men_men_n299_), .B(men_men_n324_), .C(men_men_n129_), .Y(men_men_n325_));
  NA4        u0303(.A(men_men_n84_), .B(men_men_n36_), .C(men_men_n86_), .D(i_8_), .Y(men_men_n326_));
  NA2        u0304(.A(men_men_n325_), .B(men_men_n323_), .Y(men_men_n327_));
  NO2        u0305(.A(i_6_), .B(i_8_), .Y(men_men_n328_));
  NOi21      u0306(.An(i_0_), .B(i_2_), .Y(men_men_n329_));
  AN2        u0307(.A(men_men_n329_), .B(men_men_n328_), .Y(men_men_n330_));
  NO2        u0308(.A(i_1_), .B(i_7_), .Y(men_men_n331_));
  AO220      u0309(.A0(men_men_n331_), .A1(men_men_n330_), .B0(men_men_n318_), .B1(men_men_n235_), .Y(men_men_n332_));
  NA3        u0310(.A(men_men_n332_), .B(men_men_n42_), .C(i_5_), .Y(men_men_n333_));
  NA3        u0311(.A(men_men_n333_), .B(men_men_n327_), .C(men_men_n322_), .Y(men_men_n334_));
  NO3        u0312(.A(men_men_n233_), .B(men_men_n47_), .C(i_1_), .Y(men_men_n335_));
  NO3        u0313(.A(i_8_), .B(i_2_), .C(i_1_), .Y(men_men_n336_));
  OAI210     u0314(.A0(men_men_n336_), .A1(men_men_n335_), .B0(i_6_), .Y(men_men_n337_));
  NO2        u0315(.A(men_men_n337_), .B(men_men_n317_), .Y(men_men_n338_));
  NOi21      u0316(.An(men_men_n154_), .B(men_men_n106_), .Y(men_men_n339_));
  NO2        u0317(.A(men_men_n339_), .B(men_men_n125_), .Y(men_men_n340_));
  OAI210     u0318(.A0(men_men_n340_), .A1(men_men_n338_), .B0(i_3_), .Y(men_men_n341_));
  INV        u0319(.A(men_men_n84_), .Y(men_men_n342_));
  NO2        u0320(.A(men_men_n292_), .B(men_men_n81_), .Y(men_men_n343_));
  NA2        u0321(.A(men_men_n343_), .B(men_men_n133_), .Y(men_men_n344_));
  NO2        u0322(.A(men_men_n95_), .B(men_men_n195_), .Y(men_men_n345_));
  NA2        u0323(.A(men_men_n345_), .B(men_men_n63_), .Y(men_men_n346_));
  AOI210     u0324(.A0(men_men_n346_), .A1(men_men_n344_), .B0(men_men_n342_), .Y(men_men_n347_));
  NO2        u0325(.A(men_men_n195_), .B(i_9_), .Y(men_men_n348_));
  NA2        u0326(.A(men_men_n348_), .B(men_men_n207_), .Y(men_men_n349_));
  NO2        u0327(.A(men_men_n349_), .B(men_men_n47_), .Y(men_men_n350_));
  NO2        u0328(.A(men_men_n350_), .B(men_men_n347_), .Y(men_men_n351_));
  AOI210     u0329(.A0(men_men_n351_), .A1(men_men_n341_), .B0(men_men_n163_), .Y(men_men_n352_));
  AOI210     u0330(.A0(men_men_n334_), .A1(men_men_n309_), .B0(men_men_n352_), .Y(men_men_n353_));
  NOi32      u0331(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n354_));
  INV        u0332(.A(men_men_n354_), .Y(men_men_n355_));
  NAi21      u0333(.An(i_0_), .B(i_6_), .Y(men_men_n356_));
  NAi21      u0334(.An(i_1_), .B(i_5_), .Y(men_men_n357_));
  NA2        u0335(.A(men_men_n357_), .B(men_men_n356_), .Y(men_men_n358_));
  NA2        u0336(.A(men_men_n358_), .B(men_men_n25_), .Y(men_men_n359_));
  OAI210     u0337(.A0(men_men_n359_), .A1(men_men_n160_), .B0(men_men_n246_), .Y(men_men_n360_));
  NAi41      u0338(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n361_));
  AOI210     u0339(.A0(men_men_n361_), .A1(men_men_n160_), .B0(men_men_n158_), .Y(men_men_n362_));
  NOi32      u0340(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n363_));
  NO2        u0341(.A(i_1_), .B(men_men_n103_), .Y(men_men_n364_));
  NAi21      u0342(.An(i_3_), .B(i_4_), .Y(men_men_n365_));
  NO2        u0343(.A(men_men_n365_), .B(i_9_), .Y(men_men_n366_));
  AN2        u0344(.A(i_6_), .B(i_7_), .Y(men_men_n367_));
  OAI210     u0345(.A0(men_men_n367_), .A1(men_men_n364_), .B0(men_men_n366_), .Y(men_men_n368_));
  NA2        u0346(.A(i_2_), .B(i_7_), .Y(men_men_n369_));
  NO2        u0347(.A(men_men_n365_), .B(i_10_), .Y(men_men_n370_));
  NO2        u0348(.A(men_men_n368_), .B(men_men_n187_), .Y(men_men_n371_));
  AOI210     u0349(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n372_));
  OAI210     u0350(.A0(men_men_n372_), .A1(men_men_n190_), .B0(men_men_n370_), .Y(men_men_n373_));
  NO2        u0351(.A(men_men_n373_), .B(i_5_), .Y(men_men_n374_));
  NO4        u0352(.A(men_men_n374_), .B(men_men_n371_), .C(men_men_n362_), .D(men_men_n360_), .Y(men_men_n375_));
  NO2        u0353(.A(men_men_n375_), .B(men_men_n355_), .Y(men_men_n376_));
  NO2        u0354(.A(men_men_n59_), .B(men_men_n25_), .Y(men_men_n377_));
  AN2        u0355(.A(i_12_), .B(i_5_), .Y(men_men_n378_));
  NO2        u0356(.A(i_4_), .B(men_men_n26_), .Y(men_men_n379_));
  NA2        u0357(.A(men_men_n379_), .B(men_men_n378_), .Y(men_men_n380_));
  NO2        u0358(.A(i_11_), .B(i_6_), .Y(men_men_n381_));
  NO2        u0359(.A(men_men_n243_), .B(i_5_), .Y(men_men_n382_));
  NO2        u0360(.A(i_5_), .B(i_10_), .Y(men_men_n383_));
  NO2        u0361(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n384_));
  NO3        u0362(.A(men_men_n86_), .B(men_men_n49_), .C(i_9_), .Y(men_men_n385_));
  NO2        u0363(.A(i_3_), .B(men_men_n103_), .Y(men_men_n386_));
  NO2        u0364(.A(i_11_), .B(i_12_), .Y(men_men_n387_));
  NA2        u0365(.A(men_men_n383_), .B(men_men_n237_), .Y(men_men_n388_));
  NA3        u0366(.A(men_men_n115_), .B(men_men_n42_), .C(i_11_), .Y(men_men_n389_));
  OAI220     u0367(.A0(men_men_n389_), .A1(men_men_n220_), .B0(men_men_n388_), .B1(men_men_n326_), .Y(men_men_n390_));
  NAi21      u0368(.An(i_13_), .B(i_0_), .Y(men_men_n391_));
  NO2        u0369(.A(men_men_n391_), .B(men_men_n240_), .Y(men_men_n392_));
  NA2        u0370(.A(men_men_n390_), .B(men_men_n392_), .Y(men_men_n393_));
  INV        u0371(.A(men_men_n393_), .Y(men_men_n394_));
  NO3        u0372(.A(i_1_), .B(i_12_), .C(men_men_n86_), .Y(men_men_n395_));
  NO2        u0373(.A(i_0_), .B(i_11_), .Y(men_men_n396_));
  INV        u0374(.A(i_5_), .Y(men_men_n397_));
  AN2        u0375(.A(i_1_), .B(i_6_), .Y(men_men_n398_));
  NOi21      u0376(.An(i_2_), .B(i_12_), .Y(men_men_n399_));
  NA2        u0377(.A(men_men_n399_), .B(men_men_n398_), .Y(men_men_n400_));
  NO2        u0378(.A(men_men_n400_), .B(men_men_n397_), .Y(men_men_n401_));
  NA2        u0379(.A(men_men_n143_), .B(i_9_), .Y(men_men_n402_));
  NO2        u0380(.A(men_men_n402_), .B(i_4_), .Y(men_men_n403_));
  NA2        u0381(.A(men_men_n401_), .B(men_men_n403_), .Y(men_men_n404_));
  NAi21      u0382(.An(i_9_), .B(i_4_), .Y(men_men_n405_));
  OR2        u0383(.A(i_13_), .B(i_10_), .Y(men_men_n406_));
  NO3        u0384(.A(men_men_n406_), .B(men_men_n119_), .C(men_men_n405_), .Y(men_men_n407_));
  OR2        u0385(.A(men_men_n218_), .B(men_men_n217_), .Y(men_men_n408_));
  NO2        u0386(.A(men_men_n103_), .B(men_men_n25_), .Y(men_men_n409_));
  NA2        u0387(.A(men_men_n287_), .B(men_men_n409_), .Y(men_men_n410_));
  NA2        u0388(.A(men_men_n280_), .B(men_men_n212_), .Y(men_men_n411_));
  OAI220     u0389(.A0(men_men_n411_), .A1(men_men_n408_), .B0(men_men_n410_), .B1(men_men_n339_), .Y(men_men_n412_));
  INV        u0390(.A(men_men_n412_), .Y(men_men_n413_));
  AOI210     u0391(.A0(men_men_n413_), .A1(men_men_n404_), .B0(men_men_n26_), .Y(men_men_n414_));
  AOI220     u0392(.A0(men_men_n294_), .A1(men_men_n290_), .B0(men_men_n291_), .B1(men_men_n310_), .Y(men_men_n415_));
  NO2        u0393(.A(men_men_n415_), .B(men_men_n171_), .Y(men_men_n416_));
  NO2        u0394(.A(men_men_n184_), .B(men_men_n86_), .Y(men_men_n417_));
  AOI220     u0395(.A0(men_men_n417_), .A1(men_men_n293_), .B0(men_men_n282_), .B1(men_men_n212_), .Y(men_men_n418_));
  NO2        u0396(.A(men_men_n418_), .B(men_men_n289_), .Y(men_men_n419_));
  NO2        u0397(.A(men_men_n419_), .B(men_men_n416_), .Y(men_men_n420_));
  NA2        u0398(.A(men_men_n195_), .B(i_10_), .Y(men_men_n421_));
  NA3        u0399(.A(men_men_n258_), .B(men_men_n64_), .C(i_2_), .Y(men_men_n422_));
  NA2        u0400(.A(men_men_n294_), .B(men_men_n235_), .Y(men_men_n423_));
  OAI220     u0401(.A0(men_men_n423_), .A1(men_men_n184_), .B0(men_men_n422_), .B1(men_men_n421_), .Y(men_men_n424_));
  NO2        u0402(.A(i_3_), .B(men_men_n49_), .Y(men_men_n425_));
  NA3        u0403(.A(men_men_n331_), .B(men_men_n330_), .C(men_men_n425_), .Y(men_men_n426_));
  NA2        u0404(.A(men_men_n312_), .B(men_men_n317_), .Y(men_men_n427_));
  OAI210     u0405(.A0(men_men_n427_), .A1(men_men_n191_), .B0(men_men_n426_), .Y(men_men_n428_));
  NO2        u0406(.A(men_men_n428_), .B(men_men_n424_), .Y(men_men_n429_));
  AOI210     u0407(.A0(men_men_n429_), .A1(men_men_n420_), .B0(men_men_n274_), .Y(men_men_n430_));
  NO4        u0408(.A(men_men_n430_), .B(men_men_n414_), .C(men_men_n394_), .D(men_men_n376_), .Y(men_men_n431_));
  NO2        u0409(.A(men_men_n63_), .B(i_4_), .Y(men_men_n432_));
  NO2        u0410(.A(men_men_n73_), .B(i_13_), .Y(men_men_n433_));
  NO2        u0411(.A(i_10_), .B(i_9_), .Y(men_men_n434_));
  NAi21      u0412(.An(i_12_), .B(i_8_), .Y(men_men_n435_));
  NO2        u0413(.A(men_men_n435_), .B(i_3_), .Y(men_men_n436_));
  NA2        u0414(.A(men_men_n305_), .B(i_0_), .Y(men_men_n437_));
  NO3        u0415(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n438_));
  NA2        u0416(.A(men_men_n269_), .B(men_men_n99_), .Y(men_men_n439_));
  NA2        u0417(.A(men_men_n439_), .B(men_men_n438_), .Y(men_men_n440_));
  NA2        u0418(.A(i_8_), .B(i_9_), .Y(men_men_n441_));
  AOI210     u0419(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(men_men_n442_));
  OR2        u0420(.A(men_men_n442_), .B(men_men_n441_), .Y(men_men_n443_));
  NA2        u0421(.A(men_men_n287_), .B(men_men_n207_), .Y(men_men_n444_));
  OAI220     u0422(.A0(men_men_n444_), .A1(men_men_n443_), .B0(men_men_n440_), .B1(men_men_n437_), .Y(men_men_n445_));
  NA2        u0423(.A(men_men_n251_), .B(men_men_n304_), .Y(men_men_n446_));
  NO3        u0424(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n447_));
  INV        u0425(.A(men_men_n447_), .Y(men_men_n448_));
  NA3        u0426(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n449_));
  NA4        u0427(.A(men_men_n146_), .B(men_men_n118_), .C(men_men_n80_), .D(men_men_n23_), .Y(men_men_n450_));
  OAI220     u0428(.A0(men_men_n450_), .A1(men_men_n449_), .B0(men_men_n448_), .B1(men_men_n446_), .Y(men_men_n451_));
  NO2        u0429(.A(men_men_n451_), .B(men_men_n445_), .Y(men_men_n452_));
  INV        u0430(.A(men_men_n293_), .Y(men_men_n453_));
  OR2        u0431(.A(men_men_n453_), .B(men_men_n209_), .Y(men_men_n454_));
  OA210      u0432(.A0(men_men_n349_), .A1(men_men_n103_), .B0(men_men_n295_), .Y(men_men_n455_));
  OA220      u0433(.A0(men_men_n455_), .A1(men_men_n163_), .B0(men_men_n454_), .B1(men_men_n232_), .Y(men_men_n456_));
  NA2        u0434(.A(men_men_n98_), .B(i_13_), .Y(men_men_n457_));
  NO2        u0435(.A(i_2_), .B(i_13_), .Y(men_men_n458_));
  NO3        u0436(.A(i_4_), .B(men_men_n49_), .C(i_8_), .Y(men_men_n459_));
  NO2        u0437(.A(i_6_), .B(i_7_), .Y(men_men_n460_));
  NA2        u0438(.A(men_men_n460_), .B(men_men_n459_), .Y(men_men_n461_));
  NO2        u0439(.A(i_11_), .B(i_1_), .Y(men_men_n462_));
  NO2        u0440(.A(men_men_n73_), .B(i_3_), .Y(men_men_n463_));
  OR2        u0441(.A(i_11_), .B(i_8_), .Y(men_men_n464_));
  NOi21      u0442(.An(i_2_), .B(i_7_), .Y(men_men_n465_));
  NAi31      u0443(.An(men_men_n464_), .B(men_men_n465_), .C(men_men_n463_), .Y(men_men_n466_));
  NO2        u0444(.A(men_men_n406_), .B(i_6_), .Y(men_men_n467_));
  NA2        u0445(.A(men_men_n467_), .B(men_men_n432_), .Y(men_men_n468_));
  NO2        u0446(.A(men_men_n468_), .B(men_men_n466_), .Y(men_men_n469_));
  NO2        u0447(.A(i_3_), .B(men_men_n195_), .Y(men_men_n470_));
  NO2        u0448(.A(i_6_), .B(i_10_), .Y(men_men_n471_));
  NA4        u0449(.A(men_men_n471_), .B(men_men_n309_), .C(men_men_n470_), .D(men_men_n237_), .Y(men_men_n472_));
  NO2        u0450(.A(men_men_n472_), .B(men_men_n156_), .Y(men_men_n473_));
  NA3        u0451(.A(men_men_n245_), .B(men_men_n173_), .C(men_men_n133_), .Y(men_men_n474_));
  NA2        u0452(.A(men_men_n47_), .B(men_men_n45_), .Y(men_men_n475_));
  NO2        u0453(.A(men_men_n158_), .B(i_3_), .Y(men_men_n476_));
  NAi31      u0454(.An(men_men_n475_), .B(men_men_n476_), .C(men_men_n226_), .Y(men_men_n477_));
  NA3        u0455(.A(men_men_n384_), .B(men_men_n180_), .C(men_men_n150_), .Y(men_men_n478_));
  NA3        u0456(.A(men_men_n478_), .B(men_men_n477_), .C(men_men_n474_), .Y(men_men_n479_));
  NO3        u0457(.A(men_men_n479_), .B(men_men_n473_), .C(men_men_n469_), .Y(men_men_n480_));
  NA2        u0458(.A(men_men_n438_), .B(men_men_n378_), .Y(men_men_n481_));
  NA2        u0459(.A(men_men_n447_), .B(men_men_n383_), .Y(men_men_n482_));
  NO2        u0460(.A(men_men_n482_), .B(men_men_n224_), .Y(men_men_n483_));
  NAi21      u0461(.An(men_men_n218_), .B(men_men_n387_), .Y(men_men_n484_));
  NA2        u0462(.A(men_men_n331_), .B(men_men_n219_), .Y(men_men_n485_));
  NO2        u0463(.A(men_men_n26_), .B(i_5_), .Y(men_men_n486_));
  NO2        u0464(.A(i_0_), .B(men_men_n86_), .Y(men_men_n487_));
  NA3        u0465(.A(men_men_n487_), .B(men_men_n486_), .C(men_men_n143_), .Y(men_men_n488_));
  OR3        u0466(.A(men_men_n299_), .B(men_men_n38_), .C(men_men_n47_), .Y(men_men_n489_));
  OAI220     u0467(.A0(men_men_n489_), .A1(men_men_n488_), .B0(men_men_n485_), .B1(men_men_n484_), .Y(men_men_n490_));
  NA2        u0468(.A(men_men_n27_), .B(i_10_), .Y(men_men_n491_));
  NA2        u0469(.A(men_men_n309_), .B(men_men_n239_), .Y(men_men_n492_));
  OAI220     u0470(.A0(men_men_n492_), .A1(men_men_n422_), .B0(men_men_n491_), .B1(men_men_n457_), .Y(men_men_n493_));
  NA4        u0471(.A(men_men_n302_), .B(men_men_n223_), .C(men_men_n73_), .D(men_men_n237_), .Y(men_men_n494_));
  NO2        u0472(.A(men_men_n494_), .B(men_men_n461_), .Y(men_men_n495_));
  NO4        u0473(.A(men_men_n495_), .B(men_men_n493_), .C(men_men_n490_), .D(men_men_n483_), .Y(men_men_n496_));
  NA4        u0474(.A(men_men_n496_), .B(men_men_n480_), .C(men_men_n456_), .D(men_men_n452_), .Y(men_men_n497_));
  NA3        u0475(.A(men_men_n302_), .B(men_men_n177_), .C(men_men_n175_), .Y(men_men_n498_));
  OAI210     u0476(.A0(men_men_n297_), .A1(men_men_n182_), .B0(men_men_n498_), .Y(men_men_n499_));
  AN2        u0477(.A(men_men_n290_), .B(men_men_n234_), .Y(men_men_n500_));
  NA2        u0478(.A(men_men_n500_), .B(men_men_n499_), .Y(men_men_n501_));
  NA2        u0479(.A(men_men_n309_), .B(men_men_n165_), .Y(men_men_n502_));
  OAI210     u0480(.A0(men_men_n502_), .A1(men_men_n232_), .B0(men_men_n303_), .Y(men_men_n503_));
  NA2        u0481(.A(men_men_n503_), .B(men_men_n318_), .Y(men_men_n504_));
  NA4        u0482(.A(men_men_n433_), .B(men_men_n432_), .C(men_men_n205_), .D(i_2_), .Y(men_men_n505_));
  INV        u0483(.A(men_men_n505_), .Y(men_men_n506_));
  NA2        u0484(.A(men_men_n378_), .B(men_men_n225_), .Y(men_men_n507_));
  NA2        u0485(.A(men_men_n354_), .B(men_men_n73_), .Y(men_men_n508_));
  NA2        u0486(.A(men_men_n367_), .B(men_men_n363_), .Y(men_men_n509_));
  OR2        u0487(.A(men_men_n507_), .B(men_men_n509_), .Y(men_men_n510_));
  NO2        u0488(.A(men_men_n36_), .B(i_8_), .Y(men_men_n511_));
  NAi41      u0489(.An(men_men_n508_), .B(men_men_n471_), .C(men_men_n511_), .D(men_men_n47_), .Y(men_men_n512_));
  AOI210     u0490(.A0(men_men_n39_), .A1(i_13_), .B0(men_men_n407_), .Y(men_men_n513_));
  NA3        u0491(.A(men_men_n513_), .B(men_men_n512_), .C(men_men_n510_), .Y(men_men_n514_));
  AOI210     u0492(.A0(men_men_n506_), .A1(men_men_n206_), .B0(men_men_n514_), .Y(men_men_n515_));
  NO2        u0493(.A(i_7_), .B(men_men_n201_), .Y(men_men_n516_));
  OR2        u0494(.A(men_men_n184_), .B(i_4_), .Y(men_men_n517_));
  NO2        u0495(.A(men_men_n517_), .B(men_men_n86_), .Y(men_men_n518_));
  NA2        u0496(.A(men_men_n518_), .B(men_men_n516_), .Y(men_men_n519_));
  NA4        u0497(.A(men_men_n519_), .B(men_men_n515_), .C(men_men_n504_), .D(men_men_n501_), .Y(men_men_n520_));
  NA2        u0498(.A(men_men_n382_), .B(men_men_n293_), .Y(men_men_n521_));
  OAI210     u0499(.A0(men_men_n380_), .A1(men_men_n170_), .B0(men_men_n521_), .Y(men_men_n522_));
  NO2        u0500(.A(i_12_), .B(men_men_n195_), .Y(men_men_n523_));
  NA2        u0501(.A(men_men_n523_), .B(men_men_n225_), .Y(men_men_n524_));
  NA2        u0502(.A(men_men_n471_), .B(men_men_n27_), .Y(men_men_n525_));
  NO2        u0503(.A(men_men_n525_), .B(men_men_n524_), .Y(men_men_n526_));
  NOi31      u0504(.An(men_men_n312_), .B(men_men_n406_), .C(men_men_n38_), .Y(men_men_n527_));
  OAI210     u0505(.A0(men_men_n527_), .A1(men_men_n526_), .B0(men_men_n522_), .Y(men_men_n528_));
  NO2        u0506(.A(i_8_), .B(i_7_), .Y(men_men_n529_));
  OAI210     u0507(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(men_men_n530_));
  NA2        u0508(.A(men_men_n530_), .B(men_men_n223_), .Y(men_men_n531_));
  AOI220     u0509(.A0(men_men_n319_), .A1(men_men_n40_), .B0(men_men_n235_), .B1(men_men_n208_), .Y(men_men_n532_));
  OAI220     u0510(.A0(men_men_n532_), .A1(men_men_n517_), .B0(men_men_n531_), .B1(men_men_n243_), .Y(men_men_n533_));
  NA2        u0511(.A(men_men_n45_), .B(i_10_), .Y(men_men_n534_));
  NO2        u0512(.A(men_men_n534_), .B(i_6_), .Y(men_men_n535_));
  NA3        u0513(.A(men_men_n535_), .B(men_men_n533_), .C(men_men_n529_), .Y(men_men_n536_));
  AOI220     u0514(.A0(men_men_n417_), .A1(men_men_n319_), .B0(men_men_n247_), .B1(men_men_n244_), .Y(men_men_n537_));
  OAI220     u0515(.A0(men_men_n537_), .A1(men_men_n265_), .B0(men_men_n457_), .B1(men_men_n134_), .Y(men_men_n538_));
  NA2        u0516(.A(men_men_n538_), .B(men_men_n268_), .Y(men_men_n539_));
  NA3        u0517(.A(men_men_n539_), .B(men_men_n536_), .C(men_men_n528_), .Y(men_men_n540_));
  NA3        u0518(.A(men_men_n219_), .B(men_men_n71_), .C(men_men_n45_), .Y(men_men_n541_));
  NA2        u0519(.A(men_men_n287_), .B(men_men_n84_), .Y(men_men_n542_));
  AOI210     u0520(.A0(men_men_n541_), .A1(men_men_n344_), .B0(men_men_n542_), .Y(men_men_n543_));
  NA2        u0521(.A(men_men_n223_), .B(men_men_n222_), .Y(men_men_n544_));
  NA2        u0522(.A(men_men_n434_), .B(men_men_n221_), .Y(men_men_n545_));
  NO2        u0523(.A(men_men_n544_), .B(men_men_n545_), .Y(men_men_n546_));
  NA2        u0524(.A(i_0_), .B(men_men_n49_), .Y(men_men_n547_));
  NO2        u0525(.A(men_men_n546_), .B(men_men_n543_), .Y(men_men_n548_));
  NO4        u0526(.A(men_men_n252_), .B(men_men_n43_), .C(i_2_), .D(men_men_n49_), .Y(men_men_n549_));
  NO3        u0527(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n550_));
  NO2        u0528(.A(men_men_n233_), .B(men_men_n36_), .Y(men_men_n551_));
  AN2        u0529(.A(men_men_n551_), .B(men_men_n550_), .Y(men_men_n552_));
  OA210      u0530(.A0(men_men_n552_), .A1(men_men_n549_), .B0(men_men_n354_), .Y(men_men_n553_));
  NO2        u0531(.A(men_men_n406_), .B(i_1_), .Y(men_men_n554_));
  NOi31      u0532(.An(men_men_n554_), .B(men_men_n439_), .C(men_men_n73_), .Y(men_men_n555_));
  AN4        u0533(.A(men_men_n555_), .B(men_men_n403_), .C(men_men_n486_), .D(i_2_), .Y(men_men_n556_));
  NO2        u0534(.A(men_men_n415_), .B(men_men_n178_), .Y(men_men_n557_));
  NO3        u0535(.A(men_men_n557_), .B(men_men_n556_), .C(men_men_n553_), .Y(men_men_n558_));
  NOi21      u0536(.An(i_10_), .B(i_6_), .Y(men_men_n559_));
  NO2        u0537(.A(men_men_n86_), .B(men_men_n25_), .Y(men_men_n560_));
  AOI220     u0538(.A0(men_men_n287_), .A1(men_men_n560_), .B0(men_men_n278_), .B1(men_men_n559_), .Y(men_men_n561_));
  NO2        u0539(.A(men_men_n561_), .B(men_men_n437_), .Y(men_men_n562_));
  NO2        u0540(.A(men_men_n117_), .B(men_men_n23_), .Y(men_men_n563_));
  NA2        u0541(.A(men_men_n312_), .B(men_men_n165_), .Y(men_men_n564_));
  AOI220     u0542(.A0(men_men_n564_), .A1(men_men_n423_), .B0(men_men_n185_), .B1(men_men_n183_), .Y(men_men_n565_));
  NO2        u0543(.A(men_men_n565_), .B(men_men_n562_), .Y(men_men_n566_));
  INV        u0544(.A(men_men_n315_), .Y(men_men_n567_));
  NO2        u0545(.A(i_12_), .B(men_men_n86_), .Y(men_men_n568_));
  NA3        u0546(.A(men_men_n568_), .B(men_men_n278_), .C(men_men_n547_), .Y(men_men_n569_));
  NA3        u0547(.A(men_men_n381_), .B(men_men_n287_), .C(men_men_n219_), .Y(men_men_n570_));
  AOI210     u0548(.A0(men_men_n570_), .A1(men_men_n569_), .B0(men_men_n567_), .Y(men_men_n571_));
  NA2        u0549(.A(men_men_n175_), .B(i_0_), .Y(men_men_n572_));
  NO3        u0550(.A(men_men_n572_), .B(men_men_n337_), .C(men_men_n297_), .Y(men_men_n573_));
  NO2        u0551(.A(men_men_n573_), .B(men_men_n571_), .Y(men_men_n574_));
  NA4        u0552(.A(men_men_n574_), .B(men_men_n566_), .C(men_men_n558_), .D(men_men_n548_), .Y(men_men_n575_));
  NO4        u0553(.A(men_men_n575_), .B(men_men_n540_), .C(men_men_n520_), .D(men_men_n497_), .Y(men_men_n576_));
  NA4        u0554(.A(men_men_n576_), .B(men_men_n431_), .C(men_men_n353_), .D(men_men_n308_), .Y(men7));
  NO2        u0555(.A(men_men_n95_), .B(men_men_n55_), .Y(men_men_n578_));
  NO2        u0556(.A(men_men_n110_), .B(men_men_n92_), .Y(men_men_n579_));
  NA2        u0557(.A(men_men_n379_), .B(men_men_n579_), .Y(men_men_n580_));
  NA2        u0558(.A(men_men_n471_), .B(men_men_n84_), .Y(men_men_n581_));
  NA2        u0559(.A(i_11_), .B(men_men_n195_), .Y(men_men_n582_));
  NA2        u0560(.A(men_men_n145_), .B(men_men_n582_), .Y(men_men_n583_));
  OAI210     u0561(.A0(men_men_n583_), .A1(men_men_n581_), .B0(men_men_n580_), .Y(men_men_n584_));
  NA3        u0562(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n585_));
  NO2        u0563(.A(men_men_n237_), .B(i_4_), .Y(men_men_n586_));
  NA2        u0564(.A(men_men_n586_), .B(i_8_), .Y(men_men_n587_));
  NO2        u0565(.A(men_men_n107_), .B(men_men_n585_), .Y(men_men_n588_));
  NA2        u0566(.A(i_2_), .B(men_men_n86_), .Y(men_men_n589_));
  OAI210     u0567(.A0(men_men_n89_), .A1(men_men_n205_), .B0(men_men_n206_), .Y(men_men_n590_));
  NO2        u0568(.A(i_7_), .B(men_men_n37_), .Y(men_men_n591_));
  NA2        u0569(.A(i_4_), .B(i_8_), .Y(men_men_n592_));
  AOI210     u0570(.A0(men_men_n592_), .A1(men_men_n302_), .B0(men_men_n591_), .Y(men_men_n593_));
  OAI220     u0571(.A0(men_men_n593_), .A1(men_men_n589_), .B0(men_men_n590_), .B1(i_13_), .Y(men_men_n594_));
  NO4        u0572(.A(men_men_n594_), .B(men_men_n588_), .C(men_men_n584_), .D(men_men_n578_), .Y(men_men_n595_));
  AOI210     u0573(.A0(men_men_n129_), .A1(men_men_n62_), .B0(i_10_), .Y(men_men_n596_));
  AOI210     u0574(.A0(men_men_n596_), .A1(men_men_n237_), .B0(men_men_n162_), .Y(men_men_n597_));
  OR2        u0575(.A(i_6_), .B(i_10_), .Y(men_men_n598_));
  NO2        u0576(.A(men_men_n598_), .B(men_men_n23_), .Y(men_men_n599_));
  OR3        u0577(.A(i_13_), .B(i_6_), .C(i_10_), .Y(men_men_n600_));
  NO3        u0578(.A(men_men_n600_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n601_));
  INV        u0579(.A(men_men_n202_), .Y(men_men_n602_));
  NO2        u0580(.A(men_men_n601_), .B(men_men_n599_), .Y(men_men_n603_));
  OA220      u0581(.A0(men_men_n603_), .A1(men_men_n567_), .B0(men_men_n597_), .B1(men_men_n270_), .Y(men_men_n604_));
  AOI210     u0582(.A0(men_men_n604_), .A1(men_men_n595_), .B0(men_men_n63_), .Y(men_men_n605_));
  NOi21      u0583(.An(i_11_), .B(i_7_), .Y(men_men_n606_));
  AO210      u0584(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n607_));
  NO2        u0585(.A(men_men_n607_), .B(men_men_n606_), .Y(men_men_n608_));
  NA2        u0586(.A(men_men_n608_), .B(men_men_n208_), .Y(men_men_n609_));
  NA3        u0587(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n610_));
  NAi31      u0588(.An(men_men_n610_), .B(men_men_n217_), .C(i_11_), .Y(men_men_n611_));
  AOI210     u0589(.A0(men_men_n611_), .A1(men_men_n609_), .B0(men_men_n63_), .Y(men_men_n612_));
  NA2        u0590(.A(men_men_n88_), .B(men_men_n63_), .Y(men_men_n613_));
  OR2        u0591(.A(men_men_n613_), .B(men_men_n41_), .Y(men_men_n614_));
  NO3        u0592(.A(men_men_n260_), .B(men_men_n210_), .C(men_men_n582_), .Y(men_men_n615_));
  OAI210     u0593(.A0(men_men_n615_), .A1(men_men_n226_), .B0(men_men_n63_), .Y(men_men_n616_));
  NO2        u0594(.A(men_men_n63_), .B(i_9_), .Y(men_men_n617_));
  NO2        u0595(.A(i_1_), .B(i_12_), .Y(men_men_n618_));
  NA2        u0596(.A(men_men_n616_), .B(men_men_n614_), .Y(men_men_n619_));
  OAI210     u0597(.A0(men_men_n619_), .A1(men_men_n612_), .B0(i_6_), .Y(men_men_n620_));
  NO2        u0598(.A(men_men_n610_), .B(men_men_n110_), .Y(men_men_n621_));
  NA2        u0599(.A(men_men_n621_), .B(men_men_n568_), .Y(men_men_n622_));
  NO2        u0600(.A(men_men_n237_), .B(men_men_n86_), .Y(men_men_n623_));
  NO2        u0601(.A(men_men_n623_), .B(i_11_), .Y(men_men_n624_));
  NA2        u0602(.A(men_men_n622_), .B(men_men_n440_), .Y(men_men_n625_));
  NO4        u0603(.A(men_men_n217_), .B(men_men_n129_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n626_));
  NA2        u0604(.A(men_men_n626_), .B(men_men_n617_), .Y(men_men_n627_));
  NA2        u0605(.A(men_men_n237_), .B(i_6_), .Y(men_men_n628_));
  NO3        u0606(.A(men_men_n598_), .B(men_men_n233_), .C(men_men_n23_), .Y(men_men_n629_));
  AOI210     u0607(.A0(i_1_), .A1(men_men_n261_), .B0(men_men_n629_), .Y(men_men_n630_));
  OAI210     u0608(.A0(men_men_n630_), .A1(men_men_n45_), .B0(men_men_n627_), .Y(men_men_n631_));
  INV        u0609(.A(i_2_), .Y(men_men_n632_));
  NA2        u0610(.A(men_men_n139_), .B(i_9_), .Y(men_men_n633_));
  NA3        u0611(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n634_));
  NO2        u0612(.A(men_men_n47_), .B(i_1_), .Y(men_men_n635_));
  NA3        u0613(.A(men_men_n635_), .B(men_men_n269_), .C(men_men_n45_), .Y(men_men_n636_));
  OAI220     u0614(.A0(men_men_n636_), .A1(men_men_n634_), .B0(men_men_n633_), .B1(men_men_n632_), .Y(men_men_n637_));
  NA3        u0615(.A(men_men_n617_), .B(men_men_n315_), .C(i_6_), .Y(men_men_n638_));
  NO2        u0616(.A(men_men_n638_), .B(men_men_n23_), .Y(men_men_n639_));
  AOI210     u0617(.A0(men_men_n462_), .A1(men_men_n409_), .B0(men_men_n242_), .Y(men_men_n640_));
  NO2        u0618(.A(men_men_n640_), .B(men_men_n589_), .Y(men_men_n641_));
  NA2        u0619(.A(men_men_n635_), .B(men_men_n269_), .Y(men_men_n642_));
  NO2        u0620(.A(i_11_), .B(men_men_n37_), .Y(men_men_n643_));
  NA2        u0621(.A(men_men_n643_), .B(men_men_n24_), .Y(men_men_n644_));
  NO2        u0622(.A(men_men_n644_), .B(men_men_n642_), .Y(men_men_n645_));
  OR4        u0623(.A(men_men_n645_), .B(men_men_n641_), .C(men_men_n639_), .D(men_men_n637_), .Y(men_men_n646_));
  NO3        u0624(.A(men_men_n646_), .B(men_men_n631_), .C(men_men_n625_), .Y(men_men_n647_));
  NO2        u0625(.A(men_men_n237_), .B(men_men_n103_), .Y(men_men_n648_));
  NO2        u0626(.A(men_men_n648_), .B(men_men_n606_), .Y(men_men_n649_));
  NA2        u0627(.A(men_men_n649_), .B(i_1_), .Y(men_men_n650_));
  NO2        u0628(.A(men_men_n650_), .B(men_men_n600_), .Y(men_men_n651_));
  NO2        u0629(.A(men_men_n405_), .B(men_men_n86_), .Y(men_men_n652_));
  NA2        u0630(.A(men_men_n651_), .B(men_men_n47_), .Y(men_men_n653_));
  NA2        u0631(.A(i_3_), .B(men_men_n195_), .Y(men_men_n654_));
  NO2        u0632(.A(men_men_n654_), .B(men_men_n117_), .Y(men_men_n655_));
  AN2        u0633(.A(men_men_n655_), .B(men_men_n535_), .Y(men_men_n656_));
  NO2        u0634(.A(men_men_n233_), .B(men_men_n45_), .Y(men_men_n657_));
  NO3        u0635(.A(men_men_n657_), .B(men_men_n305_), .C(men_men_n238_), .Y(men_men_n658_));
  NO2        u0636(.A(men_men_n119_), .B(men_men_n37_), .Y(men_men_n659_));
  NO2        u0637(.A(men_men_n659_), .B(i_6_), .Y(men_men_n660_));
  NO2        u0638(.A(men_men_n86_), .B(i_9_), .Y(men_men_n661_));
  NO2        u0639(.A(men_men_n661_), .B(men_men_n63_), .Y(men_men_n662_));
  NO2        u0640(.A(men_men_n662_), .B(men_men_n618_), .Y(men_men_n663_));
  NO4        u0641(.A(men_men_n663_), .B(men_men_n660_), .C(men_men_n658_), .D(i_4_), .Y(men_men_n664_));
  NA2        u0642(.A(i_1_), .B(i_3_), .Y(men_men_n665_));
  NO2        u0643(.A(men_men_n441_), .B(men_men_n95_), .Y(men_men_n666_));
  AOI210     u0644(.A0(men_men_n657_), .A1(men_men_n559_), .B0(men_men_n666_), .Y(men_men_n667_));
  NO2        u0645(.A(men_men_n667_), .B(men_men_n665_), .Y(men_men_n668_));
  NO3        u0646(.A(men_men_n668_), .B(men_men_n664_), .C(men_men_n656_), .Y(men_men_n669_));
  NA4        u0647(.A(men_men_n669_), .B(men_men_n653_), .C(men_men_n647_), .D(men_men_n620_), .Y(men_men_n670_));
  NO3        u0648(.A(men_men_n464_), .B(i_3_), .C(i_7_), .Y(men_men_n671_));
  NOi21      u0649(.An(men_men_n671_), .B(i_10_), .Y(men_men_n672_));
  OA210      u0650(.A0(men_men_n672_), .A1(men_men_n245_), .B0(men_men_n86_), .Y(men_men_n673_));
  NO3        u0651(.A(men_men_n465_), .B(men_men_n592_), .C(men_men_n86_), .Y(men_men_n674_));
  NA2        u0652(.A(men_men_n674_), .B(men_men_n25_), .Y(men_men_n675_));
  INV        u0653(.A(men_men_n675_), .Y(men_men_n676_));
  OAI210     u0654(.A0(men_men_n676_), .A1(men_men_n673_), .B0(i_1_), .Y(men_men_n677_));
  AOI210     u0655(.A0(men_men_n269_), .A1(men_men_n99_), .B0(i_1_), .Y(men_men_n678_));
  NO2        u0656(.A(men_men_n365_), .B(i_2_), .Y(men_men_n679_));
  NA2        u0657(.A(men_men_n679_), .B(men_men_n678_), .Y(men_men_n680_));
  OAI210     u0658(.A0(men_men_n638_), .A1(men_men_n435_), .B0(men_men_n680_), .Y(men_men_n681_));
  INV        u0659(.A(men_men_n681_), .Y(men_men_n682_));
  AOI210     u0660(.A0(men_men_n682_), .A1(men_men_n677_), .B0(i_13_), .Y(men_men_n683_));
  OR2        u0661(.A(i_11_), .B(i_7_), .Y(men_men_n684_));
  NO2        u0662(.A(men_men_n55_), .B(i_12_), .Y(men_men_n685_));
  NO2        u0663(.A(men_men_n465_), .B(men_men_n24_), .Y(men_men_n686_));
  AOI220     u0664(.A0(men_men_n686_), .A1(men_men_n652_), .B0(men_men_n245_), .B1(men_men_n132_), .Y(men_men_n687_));
  OAI220     u0665(.A0(men_men_n687_), .A1(men_men_n41_), .B0(men_men_n1042_), .B1(men_men_n95_), .Y(men_men_n688_));
  INV        u0666(.A(men_men_n688_), .Y(men_men_n689_));
  NA2        u0667(.A(men_men_n381_), .B(men_men_n635_), .Y(men_men_n690_));
  NO2        u0668(.A(men_men_n690_), .B(men_men_n243_), .Y(men_men_n691_));
  AOI210     u0669(.A0(men_men_n435_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n692_));
  NOi31      u0670(.An(men_men_n692_), .B(men_men_n581_), .C(men_men_n45_), .Y(men_men_n693_));
  NA2        u0671(.A(men_men_n128_), .B(i_13_), .Y(men_men_n694_));
  NO2        u0672(.A(men_men_n634_), .B(men_men_n117_), .Y(men_men_n695_));
  INV        u0673(.A(men_men_n695_), .Y(men_men_n696_));
  OAI220     u0674(.A0(men_men_n696_), .A1(men_men_n71_), .B0(men_men_n694_), .B1(men_men_n678_), .Y(men_men_n697_));
  NO3        u0675(.A(men_men_n71_), .B(men_men_n32_), .C(men_men_n103_), .Y(men_men_n698_));
  NA2        u0676(.A(men_men_n26_), .B(men_men_n195_), .Y(men_men_n699_));
  NA2        u0677(.A(men_men_n699_), .B(i_7_), .Y(men_men_n700_));
  NO3        u0678(.A(men_men_n465_), .B(men_men_n237_), .C(men_men_n86_), .Y(men_men_n701_));
  AOI210     u0679(.A0(men_men_n701_), .A1(men_men_n700_), .B0(men_men_n698_), .Y(men_men_n702_));
  AOI220     u0680(.A0(men_men_n381_), .A1(men_men_n635_), .B0(men_men_n94_), .B1(men_men_n104_), .Y(men_men_n703_));
  OAI220     u0681(.A0(men_men_n703_), .A1(men_men_n587_), .B0(men_men_n702_), .B1(men_men_n602_), .Y(men_men_n704_));
  NO4        u0682(.A(men_men_n704_), .B(men_men_n697_), .C(men_men_n693_), .D(men_men_n691_), .Y(men_men_n705_));
  OR2        u0683(.A(i_11_), .B(i_6_), .Y(men_men_n706_));
  NA3        u0684(.A(men_men_n586_), .B(men_men_n699_), .C(i_7_), .Y(men_men_n707_));
  AOI210     u0685(.A0(men_men_n707_), .A1(men_men_n696_), .B0(men_men_n706_), .Y(men_men_n708_));
  NA3        u0686(.A(men_men_n399_), .B(men_men_n591_), .C(men_men_n99_), .Y(men_men_n709_));
  NA2        u0687(.A(men_men_n624_), .B(i_13_), .Y(men_men_n710_));
  NA2        u0688(.A(men_men_n104_), .B(men_men_n699_), .Y(men_men_n711_));
  NAi21      u0689(.An(i_11_), .B(i_12_), .Y(men_men_n712_));
  NOi41      u0690(.An(men_men_n113_), .B(men_men_n712_), .C(i_13_), .D(men_men_n86_), .Y(men_men_n713_));
  NO3        u0691(.A(men_men_n465_), .B(men_men_n568_), .C(men_men_n592_), .Y(men_men_n714_));
  AOI220     u0692(.A0(men_men_n714_), .A1(men_men_n309_), .B0(men_men_n713_), .B1(men_men_n711_), .Y(men_men_n715_));
  NA3        u0693(.A(men_men_n715_), .B(men_men_n710_), .C(men_men_n709_), .Y(men_men_n716_));
  OAI210     u0694(.A0(men_men_n716_), .A1(men_men_n708_), .B0(men_men_n63_), .Y(men_men_n717_));
  NO2        u0695(.A(i_2_), .B(i_12_), .Y(men_men_n718_));
  NA2        u0696(.A(men_men_n364_), .B(men_men_n718_), .Y(men_men_n719_));
  NA2        u0697(.A(i_8_), .B(men_men_n25_), .Y(men_men_n720_));
  NO3        u0698(.A(men_men_n720_), .B(men_men_n379_), .C(men_men_n586_), .Y(men_men_n721_));
  OAI210     u0699(.A0(men_men_n721_), .A1(men_men_n366_), .B0(men_men_n364_), .Y(men_men_n722_));
  NO2        u0700(.A(men_men_n129_), .B(i_2_), .Y(men_men_n723_));
  NA2        u0701(.A(men_men_n723_), .B(men_men_n618_), .Y(men_men_n724_));
  NA3        u0702(.A(men_men_n724_), .B(men_men_n722_), .C(men_men_n719_), .Y(men_men_n725_));
  NA3        u0703(.A(men_men_n725_), .B(men_men_n46_), .C(men_men_n225_), .Y(men_men_n726_));
  NA4        u0704(.A(men_men_n726_), .B(men_men_n717_), .C(men_men_n705_), .D(men_men_n689_), .Y(men_men_n727_));
  OR4        u0705(.A(men_men_n727_), .B(men_men_n683_), .C(men_men_n670_), .D(men_men_n605_), .Y(men5));
  NA2        u0706(.A(men_men_n649_), .B(men_men_n272_), .Y(men_men_n729_));
  AN2        u0707(.A(men_men_n24_), .B(i_10_), .Y(men_men_n730_));
  NA3        u0708(.A(men_men_n730_), .B(men_men_n718_), .C(men_men_n110_), .Y(men_men_n731_));
  NO2        u0709(.A(men_men_n587_), .B(i_11_), .Y(men_men_n732_));
  NA2        u0710(.A(men_men_n89_), .B(men_men_n732_), .Y(men_men_n733_));
  NA3        u0711(.A(men_men_n733_), .B(men_men_n731_), .C(men_men_n729_), .Y(men_men_n734_));
  NO3        u0712(.A(i_11_), .B(men_men_n237_), .C(i_13_), .Y(men_men_n735_));
  NO2        u0713(.A(men_men_n125_), .B(men_men_n23_), .Y(men_men_n736_));
  NA2        u0714(.A(i_12_), .B(i_8_), .Y(men_men_n737_));
  OAI210     u0715(.A0(men_men_n47_), .A1(i_3_), .B0(men_men_n737_), .Y(men_men_n738_));
  INV        u0716(.A(men_men_n434_), .Y(men_men_n739_));
  AOI220     u0717(.A0(men_men_n315_), .A1(men_men_n563_), .B0(men_men_n738_), .B1(men_men_n736_), .Y(men_men_n740_));
  INV        u0718(.A(men_men_n740_), .Y(men_men_n741_));
  NO2        u0719(.A(men_men_n741_), .B(men_men_n734_), .Y(men_men_n742_));
  INV        u0720(.A(men_men_n173_), .Y(men_men_n743_));
  INV        u0721(.A(men_men_n245_), .Y(men_men_n744_));
  OAI210     u0722(.A0(men_men_n679_), .A1(men_men_n436_), .B0(men_men_n113_), .Y(men_men_n745_));
  AOI210     u0723(.A0(men_men_n745_), .A1(men_men_n744_), .B0(men_men_n743_), .Y(men_men_n746_));
  NO2        u0724(.A(men_men_n441_), .B(men_men_n26_), .Y(men_men_n747_));
  NO2        u0725(.A(men_men_n747_), .B(men_men_n409_), .Y(men_men_n748_));
  NA2        u0726(.A(men_men_n748_), .B(i_2_), .Y(men_men_n749_));
  INV        u0727(.A(men_men_n749_), .Y(men_men_n750_));
  AOI210     u0728(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n406_), .Y(men_men_n751_));
  AOI210     u0729(.A0(men_men_n751_), .A1(men_men_n750_), .B0(men_men_n746_), .Y(men_men_n752_));
  NO2        u0730(.A(men_men_n192_), .B(men_men_n126_), .Y(men_men_n753_));
  OAI210     u0731(.A0(men_men_n753_), .A1(men_men_n736_), .B0(i_2_), .Y(men_men_n754_));
  INV        u0732(.A(men_men_n174_), .Y(men_men_n755_));
  NO3        u0733(.A(men_men_n607_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n756_));
  AOI210     u0734(.A0(men_men_n755_), .A1(men_men_n89_), .B0(men_men_n756_), .Y(men_men_n757_));
  AOI210     u0735(.A0(men_men_n757_), .A1(men_men_n754_), .B0(men_men_n195_), .Y(men_men_n758_));
  OA210      u0736(.A0(men_men_n608_), .A1(men_men_n127_), .B0(i_13_), .Y(men_men_n759_));
  NA2        u0737(.A(men_men_n202_), .B(men_men_n205_), .Y(men_men_n760_));
  NA2        u0738(.A(men_men_n152_), .B(men_men_n582_), .Y(men_men_n761_));
  AOI210     u0739(.A0(men_men_n761_), .A1(men_men_n760_), .B0(men_men_n369_), .Y(men_men_n762_));
  AOI210     u0740(.A0(men_men_n210_), .A1(men_men_n149_), .B0(men_men_n511_), .Y(men_men_n763_));
  NA2        u0741(.A(men_men_n763_), .B(men_men_n409_), .Y(men_men_n764_));
  NO2        u0742(.A(men_men_n104_), .B(men_men_n45_), .Y(men_men_n765_));
  INV        u0743(.A(men_men_n298_), .Y(men_men_n766_));
  NA4        u0744(.A(men_men_n766_), .B(men_men_n302_), .C(men_men_n125_), .D(men_men_n43_), .Y(men_men_n767_));
  OAI210     u0745(.A0(men_men_n767_), .A1(men_men_n765_), .B0(men_men_n764_), .Y(men_men_n768_));
  NO4        u0746(.A(men_men_n768_), .B(men_men_n762_), .C(men_men_n759_), .D(men_men_n758_), .Y(men_men_n769_));
  NA2        u0747(.A(men_men_n563_), .B(men_men_n28_), .Y(men_men_n770_));
  NA2        u0748(.A(men_men_n735_), .B(men_men_n279_), .Y(men_men_n771_));
  NA2        u0749(.A(men_men_n771_), .B(men_men_n770_), .Y(men_men_n772_));
  NO2        u0750(.A(men_men_n62_), .B(i_12_), .Y(men_men_n773_));
  NO2        u0751(.A(men_men_n773_), .B(men_men_n127_), .Y(men_men_n774_));
  NO2        u0752(.A(men_men_n774_), .B(men_men_n582_), .Y(men_men_n775_));
  AOI220     u0753(.A0(men_men_n775_), .A1(men_men_n36_), .B0(men_men_n772_), .B1(men_men_n47_), .Y(men_men_n776_));
  NA4        u0754(.A(men_men_n776_), .B(men_men_n769_), .C(men_men_n752_), .D(men_men_n742_), .Y(men6));
  NO3        u0755(.A(men_men_n256_), .B(men_men_n304_), .C(i_1_), .Y(men_men_n778_));
  NO2        u0756(.A(men_men_n187_), .B(men_men_n140_), .Y(men_men_n779_));
  OAI210     u0757(.A0(men_men_n779_), .A1(men_men_n778_), .B0(men_men_n723_), .Y(men_men_n780_));
  NA4        u0758(.A(men_men_n383_), .B(men_men_n470_), .C(men_men_n71_), .D(men_men_n103_), .Y(men_men_n781_));
  INV        u0759(.A(men_men_n781_), .Y(men_men_n782_));
  NO2        u0760(.A(men_men_n220_), .B(men_men_n475_), .Y(men_men_n783_));
  NO2        u0761(.A(i_11_), .B(i_9_), .Y(men_men_n784_));
  NO2        u0762(.A(men_men_n782_), .B(men_men_n324_), .Y(men_men_n785_));
  AO210      u0763(.A0(men_men_n785_), .A1(men_men_n780_), .B0(i_12_), .Y(men_men_n786_));
  NA2        u0764(.A(men_men_n370_), .B(men_men_n331_), .Y(men_men_n787_));
  NA2        u0765(.A(men_men_n568_), .B(men_men_n63_), .Y(men_men_n788_));
  NA2        u0766(.A(men_men_n672_), .B(men_men_n71_), .Y(men_men_n789_));
  BUFFER     u0767(.A(men_men_n613_), .Y(men_men_n790_));
  NA4        u0768(.A(men_men_n790_), .B(men_men_n789_), .C(men_men_n788_), .D(men_men_n787_), .Y(men_men_n791_));
  INV        u0769(.A(men_men_n199_), .Y(men_men_n792_));
  AOI220     u0770(.A0(men_men_n792_), .A1(men_men_n784_), .B0(men_men_n791_), .B1(men_men_n73_), .Y(men_men_n793_));
  INV        u0771(.A(men_men_n323_), .Y(men_men_n794_));
  NA2        u0772(.A(men_men_n75_), .B(men_men_n132_), .Y(men_men_n795_));
  INV        u0773(.A(men_men_n125_), .Y(men_men_n796_));
  NA2        u0774(.A(men_men_n796_), .B(men_men_n47_), .Y(men_men_n797_));
  AOI210     u0775(.A0(men_men_n797_), .A1(men_men_n795_), .B0(men_men_n794_), .Y(men_men_n798_));
  NO2        u0776(.A(men_men_n252_), .B(i_9_), .Y(men_men_n799_));
  NA2        u0777(.A(men_men_n799_), .B(men_men_n773_), .Y(men_men_n800_));
  AOI210     u0778(.A0(men_men_n800_), .A1(men_men_n509_), .B0(men_men_n187_), .Y(men_men_n801_));
  NO2        u0779(.A(men_men_n32_), .B(i_11_), .Y(men_men_n802_));
  NA3        u0780(.A(men_men_n802_), .B(men_men_n460_), .C(men_men_n383_), .Y(men_men_n803_));
  NAi32      u0781(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(men_men_n804_));
  NO2        u0782(.A(men_men_n706_), .B(men_men_n804_), .Y(men_men_n805_));
  OAI210     u0783(.A0(men_men_n671_), .A1(men_men_n551_), .B0(men_men_n550_), .Y(men_men_n806_));
  NAi31      u0784(.An(men_men_n805_), .B(men_men_n806_), .C(men_men_n803_), .Y(men_men_n807_));
  OR3        u0785(.A(men_men_n807_), .B(men_men_n801_), .C(men_men_n798_), .Y(men_men_n808_));
  NO2        u0786(.A(men_men_n684_), .B(i_2_), .Y(men_men_n809_));
  NA2        u0787(.A(men_men_n49_), .B(men_men_n37_), .Y(men_men_n810_));
  NO2        u0788(.A(men_men_n810_), .B(men_men_n398_), .Y(men_men_n811_));
  NA2        u0789(.A(men_men_n811_), .B(men_men_n809_), .Y(men_men_n812_));
  AO220      u0790(.A0(men_men_n358_), .A1(men_men_n348_), .B0(men_men_n385_), .B1(men_men_n582_), .Y(men_men_n813_));
  NA3        u0791(.A(men_men_n813_), .B(men_men_n257_), .C(i_7_), .Y(men_men_n814_));
  BUFFER     u0792(.A(men_men_n608_), .Y(men_men_n815_));
  NA3        u0793(.A(men_men_n815_), .B(men_men_n148_), .C(men_men_n69_), .Y(men_men_n816_));
  AO210      u0794(.A0(men_men_n482_), .A1(men_men_n739_), .B0(men_men_n36_), .Y(men_men_n817_));
  NA4        u0795(.A(men_men_n817_), .B(men_men_n816_), .C(men_men_n814_), .D(men_men_n812_), .Y(men_men_n818_));
  OAI210     u0796(.A0(men_men_n623_), .A1(i_11_), .B0(men_men_n87_), .Y(men_men_n819_));
  AOI220     u0797(.A0(men_men_n819_), .A1(men_men_n550_), .B0(men_men_n783_), .B1(men_men_n700_), .Y(men_men_n820_));
  NA3        u0798(.A(men_men_n369_), .B(men_men_n239_), .C(men_men_n148_), .Y(men_men_n821_));
  NA2        u0799(.A(men_men_n385_), .B(men_men_n70_), .Y(men_men_n822_));
  NA4        u0800(.A(men_men_n822_), .B(men_men_n821_), .C(men_men_n820_), .D(men_men_n590_), .Y(men_men_n823_));
  AO210      u0801(.A0(men_men_n511_), .A1(men_men_n47_), .B0(men_men_n88_), .Y(men_men_n824_));
  NA3        u0802(.A(men_men_n824_), .B(men_men_n471_), .C(men_men_n219_), .Y(men_men_n825_));
  AOI210     u0803(.A0(men_men_n436_), .A1(men_men_n434_), .B0(men_men_n549_), .Y(men_men_n826_));
  NO2        u0804(.A(men_men_n598_), .B(men_men_n104_), .Y(men_men_n827_));
  OAI210     u0805(.A0(men_men_n827_), .A1(men_men_n114_), .B0(men_men_n396_), .Y(men_men_n828_));
  NA3        u0806(.A(men_men_n828_), .B(men_men_n826_), .C(men_men_n825_), .Y(men_men_n829_));
  NO4        u0807(.A(men_men_n829_), .B(men_men_n823_), .C(men_men_n818_), .D(men_men_n808_), .Y(men_men_n830_));
  NA4        u0808(.A(men_men_n830_), .B(men_men_n793_), .C(men_men_n786_), .D(men_men_n375_), .Y(men3));
  NA2        u0809(.A(i_6_), .B(i_7_), .Y(men_men_n832_));
  NO2        u0810(.A(men_men_n832_), .B(i_0_), .Y(men_men_n833_));
  NO2        u0811(.A(i_11_), .B(men_men_n237_), .Y(men_men_n834_));
  OAI210     u0812(.A0(men_men_n833_), .A1(men_men_n291_), .B0(men_men_n834_), .Y(men_men_n835_));
  NO2        u0813(.A(men_men_n835_), .B(men_men_n195_), .Y(men_men_n836_));
  NO3        u0814(.A(men_men_n437_), .B(men_men_n92_), .C(men_men_n45_), .Y(men_men_n837_));
  OA210      u0815(.A0(men_men_n837_), .A1(men_men_n836_), .B0(men_men_n175_), .Y(men_men_n838_));
  NA2        u0816(.A(men_men_n821_), .B(men_men_n368_), .Y(men_men_n839_));
  NA2        u0817(.A(men_men_n839_), .B(men_men_n40_), .Y(men_men_n840_));
  NA2        u0818(.A(men_men_n399_), .B(men_men_n46_), .Y(men_men_n841_));
  NO2        u0819(.A(men_men_n840_), .B(men_men_n49_), .Y(men_men_n842_));
  NO4        u0820(.A(men_men_n372_), .B(men_men_n378_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n843_));
  NA2        u0821(.A(men_men_n187_), .B(men_men_n559_), .Y(men_men_n844_));
  NOi21      u0822(.An(men_men_n844_), .B(men_men_n843_), .Y(men_men_n845_));
  NA2        u0823(.A(men_men_n692_), .B(men_men_n661_), .Y(men_men_n846_));
  NA2        u0824(.A(men_men_n329_), .B(men_men_n425_), .Y(men_men_n847_));
  OAI220     u0825(.A0(men_men_n847_), .A1(men_men_n846_), .B0(men_men_n845_), .B1(men_men_n63_), .Y(men_men_n848_));
  NOi21      u0826(.An(i_5_), .B(i_9_), .Y(men_men_n849_));
  NA2        u0827(.A(men_men_n849_), .B(men_men_n433_), .Y(men_men_n850_));
  BUFFER     u0828(.A(men_men_n269_), .Y(men_men_n851_));
  AOI210     u0829(.A0(men_men_n851_), .A1(men_men_n462_), .B0(men_men_n674_), .Y(men_men_n852_));
  NO3        u0830(.A(men_men_n402_), .B(men_men_n269_), .C(men_men_n73_), .Y(men_men_n853_));
  NO2        u0831(.A(men_men_n176_), .B(men_men_n149_), .Y(men_men_n854_));
  AOI210     u0832(.A0(men_men_n854_), .A1(men_men_n244_), .B0(men_men_n853_), .Y(men_men_n855_));
  OAI220     u0833(.A0(men_men_n855_), .A1(men_men_n182_), .B0(men_men_n852_), .B1(men_men_n850_), .Y(men_men_n856_));
  NO4        u0834(.A(men_men_n856_), .B(men_men_n848_), .C(men_men_n842_), .D(men_men_n838_), .Y(men_men_n857_));
  NA2        u0835(.A(men_men_n187_), .B(men_men_n24_), .Y(men_men_n858_));
  NO2        u0836(.A(men_men_n659_), .B(men_men_n579_), .Y(men_men_n859_));
  NO2        u0837(.A(men_men_n859_), .B(men_men_n858_), .Y(men_men_n860_));
  NA2        u0838(.A(men_men_n309_), .B(men_men_n130_), .Y(men_men_n861_));
  NO2        u0839(.A(men_men_n861_), .B(men_men_n388_), .Y(men_men_n862_));
  NO2        u0840(.A(men_men_n862_), .B(men_men_n860_), .Y(men_men_n863_));
  NO2        u0841(.A(men_men_n383_), .B(men_men_n292_), .Y(men_men_n864_));
  NA2        u0842(.A(men_men_n864_), .B(men_men_n695_), .Y(men_men_n865_));
  NA2        u0843(.A(men_men_n560_), .B(i_0_), .Y(men_men_n866_));
  NO3        u0844(.A(men_men_n866_), .B(men_men_n380_), .C(men_men_n89_), .Y(men_men_n867_));
  INV        u0845(.A(men_men_n867_), .Y(men_men_n868_));
  NA2        u0846(.A(men_men_n735_), .B(men_men_n324_), .Y(men_men_n869_));
  AOI210     u0847(.A0(men_men_n471_), .A1(men_men_n89_), .B0(men_men_n58_), .Y(men_men_n870_));
  OAI220     u0848(.A0(men_men_n870_), .A1(men_men_n869_), .B0(men_men_n644_), .B1(men_men_n531_), .Y(men_men_n871_));
  NO2        u0849(.A(men_men_n254_), .B(men_men_n154_), .Y(men_men_n872_));
  NA2        u0850(.A(i_0_), .B(i_10_), .Y(men_men_n873_));
  AN2        u0851(.A(men_men_n872_), .B(i_6_), .Y(men_men_n874_));
  AOI220     u0852(.A0(men_men_n329_), .A1(men_men_n100_), .B0(men_men_n187_), .B1(men_men_n84_), .Y(men_men_n875_));
  NA2        u0853(.A(men_men_n554_), .B(i_4_), .Y(men_men_n876_));
  NA2        u0854(.A(men_men_n190_), .B(men_men_n205_), .Y(men_men_n877_));
  OAI220     u0855(.A0(men_men_n877_), .A1(men_men_n869_), .B0(men_men_n876_), .B1(men_men_n875_), .Y(men_men_n878_));
  NO3        u0856(.A(men_men_n878_), .B(men_men_n874_), .C(men_men_n871_), .Y(men_men_n879_));
  NA4        u0857(.A(men_men_n879_), .B(men_men_n868_), .C(men_men_n865_), .D(men_men_n863_), .Y(men_men_n880_));
  NO2        u0858(.A(men_men_n105_), .B(men_men_n37_), .Y(men_men_n881_));
  NA2        u0859(.A(i_11_), .B(i_9_), .Y(men_men_n882_));
  NO3        u0860(.A(i_12_), .B(men_men_n882_), .C(men_men_n589_), .Y(men_men_n883_));
  AN2        u0861(.A(men_men_n883_), .B(men_men_n881_), .Y(men_men_n884_));
  NO2        u0862(.A(men_men_n49_), .B(i_7_), .Y(men_men_n885_));
  NA2        u0863(.A(men_men_n384_), .B(men_men_n180_), .Y(men_men_n886_));
  NA2        u0864(.A(men_men_n886_), .B(men_men_n161_), .Y(men_men_n887_));
  NO2        u0865(.A(men_men_n176_), .B(i_0_), .Y(men_men_n888_));
  AOI210     u0866(.A0(men_men_n367_), .A1(men_men_n42_), .B0(men_men_n395_), .Y(men_men_n889_));
  NO2        u0867(.A(men_men_n889_), .B(men_men_n850_), .Y(men_men_n890_));
  NO3        u0868(.A(men_men_n890_), .B(men_men_n887_), .C(men_men_n884_), .Y(men_men_n891_));
  NA2        u0869(.A(men_men_n643_), .B(men_men_n122_), .Y(men_men_n892_));
  NO2        u0870(.A(i_6_), .B(men_men_n892_), .Y(men_men_n893_));
  AOI210     u0871(.A0(men_men_n435_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n894_));
  NA2        u0872(.A(men_men_n173_), .B(men_men_n105_), .Y(men_men_n895_));
  NOi32      u0873(.An(men_men_n894_), .Bn(men_men_n190_), .C(men_men_n895_), .Y(men_men_n896_));
  NA2        u0874(.A(men_men_n591_), .B(men_men_n324_), .Y(men_men_n897_));
  NO2        u0875(.A(men_men_n897_), .B(men_men_n841_), .Y(men_men_n898_));
  NO3        u0876(.A(men_men_n898_), .B(men_men_n896_), .C(men_men_n893_), .Y(men_men_n899_));
  NOi21      u0877(.An(i_7_), .B(i_5_), .Y(men_men_n900_));
  NOi31      u0878(.An(men_men_n900_), .B(i_0_), .C(men_men_n712_), .Y(men_men_n901_));
  NA3        u0879(.A(men_men_n901_), .B(men_men_n379_), .C(i_6_), .Y(men_men_n902_));
  BUFFER     u0880(.A(men_men_n902_), .Y(men_men_n903_));
  NO3        u0881(.A(men_men_n391_), .B(men_men_n361_), .C(men_men_n357_), .Y(men_men_n904_));
  NO2        u0882(.A(men_men_n263_), .B(men_men_n316_), .Y(men_men_n905_));
  NO2        u0883(.A(men_men_n712_), .B(men_men_n259_), .Y(men_men_n906_));
  AOI210     u0884(.A0(men_men_n906_), .A1(men_men_n905_), .B0(men_men_n904_), .Y(men_men_n907_));
  NA4        u0885(.A(men_men_n907_), .B(men_men_n903_), .C(men_men_n899_), .D(men_men_n891_), .Y(men_men_n908_));
  NO2        u0886(.A(men_men_n858_), .B(men_men_n240_), .Y(men_men_n909_));
  AN2        u0887(.A(men_men_n328_), .B(men_men_n324_), .Y(men_men_n910_));
  AN2        u0888(.A(men_men_n910_), .B(men_men_n854_), .Y(men_men_n911_));
  OAI210     u0889(.A0(men_men_n911_), .A1(men_men_n909_), .B0(i_10_), .Y(men_men_n912_));
  OA210      u0890(.A0(men_men_n460_), .A1(men_men_n223_), .B0(men_men_n459_), .Y(men_men_n913_));
  NO2        u0891(.A(men_men_n257_), .B(men_men_n47_), .Y(men_men_n914_));
  NO2        u0892(.A(men_men_n914_), .B(men_men_n189_), .Y(men_men_n915_));
  NA2        u0893(.A(men_men_n915_), .B(men_men_n460_), .Y(men_men_n916_));
  NA3        u0894(.A(men_men_n810_), .B(men_men_n377_), .C(men_men_n623_), .Y(men_men_n917_));
  NA2        u0895(.A(men_men_n95_), .B(men_men_n45_), .Y(men_men_n918_));
  NO2        u0896(.A(men_men_n75_), .B(men_men_n737_), .Y(men_men_n919_));
  AOI220     u0897(.A0(men_men_n919_), .A1(men_men_n918_), .B0(men_men_n175_), .B1(men_men_n579_), .Y(men_men_n920_));
  AOI210     u0898(.A0(men_men_n920_), .A1(men_men_n917_), .B0(men_men_n48_), .Y(men_men_n921_));
  NO3        u0899(.A(i_5_), .B(men_men_n356_), .C(men_men_n24_), .Y(men_men_n922_));
  INV        u0900(.A(men_men_n922_), .Y(men_men_n923_));
  NAi21      u0901(.An(i_9_), .B(i_5_), .Y(men_men_n924_));
  NO2        u0902(.A(men_men_n924_), .B(men_men_n391_), .Y(men_men_n925_));
  NO2        u0903(.A(men_men_n585_), .B(men_men_n107_), .Y(men_men_n926_));
  AOI220     u0904(.A0(men_men_n926_), .A1(i_0_), .B0(men_men_n925_), .B1(men_men_n608_), .Y(men_men_n927_));
  OAI220     u0905(.A0(men_men_n927_), .A1(men_men_n86_), .B0(men_men_n923_), .B1(men_men_n174_), .Y(men_men_n928_));
  NO3        u0906(.A(men_men_n928_), .B(men_men_n921_), .C(men_men_n514_), .Y(men_men_n929_));
  NA3        u0907(.A(men_men_n929_), .B(men_men_n916_), .C(men_men_n912_), .Y(men_men_n930_));
  NO3        u0908(.A(men_men_n930_), .B(men_men_n908_), .C(men_men_n880_), .Y(men_men_n931_));
  NO2        u0909(.A(i_0_), .B(men_men_n712_), .Y(men_men_n932_));
  NA2        u0910(.A(men_men_n73_), .B(men_men_n45_), .Y(men_men_n933_));
  INV        u0911(.A(men_men_n933_), .Y(men_men_n934_));
  NO3        u0912(.A(men_men_n107_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n935_));
  AO220      u0913(.A0(men_men_n935_), .A1(men_men_n934_), .B0(men_men_n932_), .B1(men_men_n175_), .Y(men_men_n936_));
  NO2        u0914(.A(men_men_n788_), .B(men_men_n895_), .Y(men_men_n937_));
  AOI210     u0915(.A0(men_men_n936_), .A1(men_men_n345_), .B0(men_men_n937_), .Y(men_men_n938_));
  NA2        u0916(.A(men_men_n723_), .B(men_men_n147_), .Y(men_men_n939_));
  INV        u0917(.A(men_men_n939_), .Y(men_men_n940_));
  NA3        u0918(.A(men_men_n940_), .B(men_men_n661_), .C(men_men_n73_), .Y(men_men_n941_));
  NO2        u0919(.A(men_men_n806_), .B(men_men_n391_), .Y(men_men_n942_));
  NA3        u0920(.A(men_men_n833_), .B(i_2_), .C(men_men_n49_), .Y(men_men_n943_));
  NA2        u0921(.A(men_men_n834_), .B(i_9_), .Y(men_men_n944_));
  AOI210     u0922(.A0(men_men_n943_), .A1(men_men_n488_), .B0(men_men_n944_), .Y(men_men_n945_));
  OAI210     u0923(.A0(men_men_n244_), .A1(i_9_), .B0(men_men_n230_), .Y(men_men_n946_));
  AOI210     u0924(.A0(men_men_n946_), .A1(men_men_n866_), .B0(men_men_n154_), .Y(men_men_n947_));
  NO3        u0925(.A(men_men_n947_), .B(men_men_n945_), .C(men_men_n942_), .Y(men_men_n948_));
  NA3        u0926(.A(men_men_n948_), .B(men_men_n941_), .C(men_men_n938_), .Y(men_men_n949_));
  NA2        u0927(.A(men_men_n910_), .B(men_men_n369_), .Y(men_men_n950_));
  AOI210     u0928(.A0(men_men_n297_), .A1(men_men_n163_), .B0(men_men_n950_), .Y(men_men_n951_));
  NA3        u0929(.A(men_men_n40_), .B(men_men_n28_), .C(men_men_n45_), .Y(men_men_n952_));
  NA2        u0930(.A(men_men_n885_), .B(men_men_n476_), .Y(men_men_n953_));
  AOI210     u0931(.A0(men_men_n952_), .A1(men_men_n163_), .B0(men_men_n953_), .Y(men_men_n954_));
  NO2        u0932(.A(men_men_n954_), .B(men_men_n951_), .Y(men_men_n955_));
  NO3        u0933(.A(men_men_n873_), .B(men_men_n849_), .C(men_men_n192_), .Y(men_men_n956_));
  AOI220     u0934(.A0(men_men_n956_), .A1(i_11_), .B0(men_men_n555_), .B1(men_men_n75_), .Y(men_men_n957_));
  NO3        u0935(.A(men_men_n211_), .B(men_men_n378_), .C(i_0_), .Y(men_men_n958_));
  OAI210     u0936(.A0(men_men_n958_), .A1(men_men_n76_), .B0(i_13_), .Y(men_men_n959_));
  INV        u0937(.A(men_men_n219_), .Y(men_men_n960_));
  OAI220     u0938(.A0(men_men_n524_), .A1(men_men_n140_), .B0(men_men_n628_), .B1(men_men_n602_), .Y(men_men_n961_));
  NA3        u0939(.A(men_men_n961_), .B(men_men_n386_), .C(men_men_n960_), .Y(men_men_n962_));
  NA4        u0940(.A(men_men_n962_), .B(men_men_n959_), .C(men_men_n957_), .D(men_men_n955_), .Y(men_men_n963_));
  NO2        u0941(.A(men_men_n243_), .B(men_men_n95_), .Y(men_men_n964_));
  AOI210     u0942(.A0(men_men_n964_), .A1(men_men_n932_), .B0(men_men_n111_), .Y(men_men_n965_));
  AOI220     u0943(.A0(men_men_n900_), .A1(men_men_n476_), .B0(men_men_n833_), .B1(men_men_n164_), .Y(men_men_n966_));
  NA2        u0944(.A(men_men_n348_), .B(men_men_n177_), .Y(men_men_n967_));
  OA220      u0945(.A0(men_men_n967_), .A1(men_men_n966_), .B0(men_men_n965_), .B1(i_5_), .Y(men_men_n968_));
  AOI210     u0946(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n176_), .Y(men_men_n969_));
  NA2        u0947(.A(men_men_n969_), .B(men_men_n913_), .Y(men_men_n970_));
  NA3        u0948(.A(men_men_n599_), .B(men_men_n187_), .C(men_men_n84_), .Y(men_men_n971_));
  INV        u0949(.A(men_men_n971_), .Y(men_men_n972_));
  NO3        u0950(.A(men_men_n841_), .B(men_men_n55_), .C(men_men_n49_), .Y(men_men_n973_));
  NA2        u0951(.A(men_men_n481_), .B(men_men_n474_), .Y(men_men_n974_));
  NO3        u0952(.A(men_men_n974_), .B(men_men_n973_), .C(men_men_n972_), .Y(men_men_n975_));
  NA3        u0953(.A(men_men_n885_), .B(men_men_n291_), .C(men_men_n230_), .Y(men_men_n976_));
  INV        u0954(.A(men_men_n976_), .Y(men_men_n977_));
  NO3        u0955(.A(men_men_n882_), .B(men_men_n219_), .C(men_men_n192_), .Y(men_men_n978_));
  NO2        u0956(.A(men_men_n978_), .B(men_men_n977_), .Y(men_men_n979_));
  NA4        u0957(.A(men_men_n979_), .B(men_men_n975_), .C(men_men_n970_), .D(men_men_n968_), .Y(men_men_n980_));
  INV        u0958(.A(men_men_n601_), .Y(men_men_n981_));
  NO3        u0959(.A(men_men_n981_), .B(men_men_n547_), .C(men_men_n342_), .Y(men_men_n982_));
  INV        u0960(.A(men_men_n982_), .Y(men_men_n983_));
  NA2        u0961(.A(men_men_n302_), .B(i_5_), .Y(men_men_n984_));
  NA2        u0962(.A(men_men_n984_), .B(men_men_n243_), .Y(men_men_n985_));
  NO4        u0963(.A(men_men_n240_), .B(men_men_n211_), .C(i_0_), .D(i_12_), .Y(men_men_n986_));
  AOI220     u0964(.A0(men_men_n986_), .A1(men_men_n985_), .B0(men_men_n782_), .B1(men_men_n177_), .Y(men_men_n987_));
  NA3        u0965(.A(men_men_n100_), .B(men_men_n559_), .C(i_11_), .Y(men_men_n988_));
  NO2        u0966(.A(men_men_n988_), .B(men_men_n156_), .Y(men_men_n989_));
  NA2        u0967(.A(men_men_n900_), .B(men_men_n458_), .Y(men_men_n990_));
  NA2        u0968(.A(men_men_n64_), .B(men_men_n103_), .Y(men_men_n991_));
  OAI220     u0969(.A0(men_men_n991_), .A1(men_men_n984_), .B0(men_men_n990_), .B1(men_men_n662_), .Y(men_men_n992_));
  AOI210     u0970(.A0(men_men_n992_), .A1(men_men_n888_), .B0(men_men_n989_), .Y(men_men_n993_));
  NA3        u0971(.A(men_men_n993_), .B(men_men_n987_), .C(men_men_n983_), .Y(men_men_n994_));
  NO4        u0972(.A(men_men_n994_), .B(men_men_n980_), .C(men_men_n963_), .D(men_men_n949_), .Y(men_men_n995_));
  OAI210     u0973(.A0(men_men_n809_), .A1(men_men_n802_), .B0(men_men_n37_), .Y(men_men_n996_));
  NA3        u0974(.A(men_men_n894_), .B(men_men_n364_), .C(i_5_), .Y(men_men_n997_));
  NA3        u0975(.A(men_men_n997_), .B(men_men_n996_), .C(men_men_n597_), .Y(men_men_n998_));
  NA2        u0976(.A(men_men_n998_), .B(men_men_n208_), .Y(men_men_n999_));
  NA2        u0977(.A(men_men_n188_), .B(men_men_n190_), .Y(men_men_n1000_));
  AO210      u0978(.A0(i_11_), .A1(men_men_n33_), .B0(men_men_n1000_), .Y(men_men_n1001_));
  OAI210     u0979(.A0(men_men_n601_), .A1(men_men_n599_), .B0(men_men_n315_), .Y(men_men_n1002_));
  NAi31      u0980(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n1003_));
  NO2        u0981(.A(men_men_n70_), .B(men_men_n1003_), .Y(men_men_n1004_));
  NO2        u0982(.A(men_men_n1004_), .B(men_men_n629_), .Y(men_men_n1005_));
  NA3        u0983(.A(men_men_n1005_), .B(men_men_n1002_), .C(men_men_n1001_), .Y(men_men_n1006_));
  NO2        u0984(.A(men_men_n449_), .B(men_men_n269_), .Y(men_men_n1007_));
  NO4        u0985(.A(men_men_n233_), .B(men_men_n146_), .C(men_men_n665_), .D(men_men_n37_), .Y(men_men_n1008_));
  NO2        u0986(.A(men_men_n1008_), .B(men_men_n1007_), .Y(men_men_n1009_));
  OAI210     u0987(.A0(men_men_n988_), .A1(men_men_n149_), .B0(men_men_n1009_), .Y(men_men_n1010_));
  AOI210     u0988(.A0(men_men_n1006_), .A1(men_men_n49_), .B0(men_men_n1010_), .Y(men_men_n1011_));
  AOI210     u0989(.A0(men_men_n1011_), .A1(men_men_n999_), .B0(men_men_n73_), .Y(men_men_n1012_));
  NO2        u0990(.A(men_men_n552_), .B(men_men_n374_), .Y(men_men_n1013_));
  NO2        u0991(.A(men_men_n1013_), .B(men_men_n743_), .Y(men_men_n1014_));
  INV        u0992(.A(men_men_n76_), .Y(men_men_n1015_));
  AOI210     u0993(.A0(men_men_n969_), .A1(men_men_n885_), .B0(men_men_n901_), .Y(men_men_n1016_));
  AOI210     u0994(.A0(men_men_n1016_), .A1(men_men_n1015_), .B0(men_men_n665_), .Y(men_men_n1017_));
  NA2        u0995(.A(men_men_n263_), .B(men_men_n57_), .Y(men_men_n1018_));
  AOI220     u0996(.A0(men_men_n1018_), .A1(men_men_n76_), .B0(men_men_n343_), .B1(men_men_n256_), .Y(men_men_n1019_));
  NO2        u0997(.A(men_men_n1019_), .B(men_men_n237_), .Y(men_men_n1020_));
  NA3        u0998(.A(men_men_n98_), .B(men_men_n304_), .C(men_men_n31_), .Y(men_men_n1021_));
  INV        u0999(.A(men_men_n1021_), .Y(men_men_n1022_));
  NO3        u1000(.A(men_men_n1022_), .B(men_men_n1020_), .C(men_men_n1017_), .Y(men_men_n1023_));
  OAI210     u1001(.A0(men_men_n271_), .A1(men_men_n159_), .B0(men_men_n89_), .Y(men_men_n1024_));
  NO2        u1002(.A(men_men_n1024_), .B(i_11_), .Y(men_men_n1025_));
  NA2        u1003(.A(men_men_n592_), .B(men_men_n217_), .Y(men_men_n1026_));
  OAI210     u1004(.A0(men_men_n1026_), .A1(men_men_n894_), .B0(men_men_n208_), .Y(men_men_n1027_));
  NA2        u1005(.A(men_men_n165_), .B(i_5_), .Y(men_men_n1028_));
  NO2        u1006(.A(men_men_n1027_), .B(men_men_n1028_), .Y(men_men_n1029_));
  NO3        u1007(.A(men_men_n59_), .B(men_men_n58_), .C(i_4_), .Y(men_men_n1030_));
  OAI210     u1008(.A0(men_men_n905_), .A1(men_men_n304_), .B0(men_men_n1030_), .Y(men_men_n1031_));
  NO2        u1009(.A(men_men_n1031_), .B(men_men_n712_), .Y(men_men_n1032_));
  NO4        u1010(.A(men_men_n924_), .B(men_men_n464_), .C(men_men_n253_), .D(men_men_n252_), .Y(men_men_n1033_));
  NO2        u1011(.A(men_men_n1033_), .B(men_men_n549_), .Y(men_men_n1034_));
  NO2        u1012(.A(men_men_n1034_), .B(men_men_n41_), .Y(men_men_n1035_));
  NO4        u1013(.A(men_men_n1035_), .B(men_men_n1032_), .C(men_men_n1029_), .D(men_men_n1025_), .Y(men_men_n1036_));
  OAI210     u1014(.A0(men_men_n1023_), .A1(i_4_), .B0(men_men_n1036_), .Y(men_men_n1037_));
  NO3        u1015(.A(men_men_n1037_), .B(men_men_n1014_), .C(men_men_n1012_), .Y(men_men_n1038_));
  NA4        u1016(.A(men_men_n1038_), .B(men_men_n995_), .C(men_men_n931_), .D(men_men_n857_), .Y(men4));
  INV        u1017(.A(men_men_n685_), .Y(men_men_n1042_));
  INV        u1018(.A(men_men_n119_), .Y(men_men_n1043_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule