// Benchmark "top" written by ABC on Thu Jun 20 14:59:15 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    men1, men2, men0, men7, men5, men6, men3, men4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output men1, men2, men0, men7, men5, men6, men3, men4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n43_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n138_, new_new_n139_,
    new_new_n140_, new_new_n142_, new_new_n143_, new_new_n144_,
    new_new_n145_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n468_,
    new_new_n469_, new_new_n470_, new_new_n471_, new_new_n472_,
    new_new_n473_, new_new_n474_, new_new_n475_, new_new_n476_,
    new_new_n477_, new_new_n478_, new_new_n479_, new_new_n480_,
    new_new_n481_, new_new_n482_, new_new_n483_, new_new_n484_,
    new_new_n485_, new_new_n486_, new_new_n487_, new_new_n488_,
    new_new_n489_, new_new_n490_, new_new_n491_, new_new_n492_,
    new_new_n493_, new_new_n494_, new_new_n495_, new_new_n496_,
    new_new_n497_, new_new_n498_, new_new_n499_, new_new_n500_,
    new_new_n501_, new_new_n502_, new_new_n503_, new_new_n504_,
    new_new_n505_, new_new_n506_, new_new_n507_, new_new_n508_,
    new_new_n509_, new_new_n510_, new_new_n511_, new_new_n512_,
    new_new_n513_, new_new_n514_, new_new_n515_, new_new_n516_,
    new_new_n517_, new_new_n518_, new_new_n519_, new_new_n520_,
    new_new_n521_, new_new_n522_, new_new_n523_, new_new_n524_,
    new_new_n525_, new_new_n526_, new_new_n527_, new_new_n528_,
    new_new_n529_, new_new_n530_, new_new_n531_, new_new_n532_,
    new_new_n533_, new_new_n534_, new_new_n535_, new_new_n536_,
    new_new_n537_, new_new_n538_, new_new_n539_, new_new_n540_,
    new_new_n541_, new_new_n542_, new_new_n543_, new_new_n544_,
    new_new_n545_, new_new_n546_, new_new_n547_, new_new_n548_,
    new_new_n549_, new_new_n550_, new_new_n551_, new_new_n552_,
    new_new_n553_, new_new_n554_, new_new_n555_, new_new_n556_,
    new_new_n557_, new_new_n558_, new_new_n559_, new_new_n560_,
    new_new_n561_, new_new_n562_, new_new_n563_, new_new_n564_,
    new_new_n565_, new_new_n566_, new_new_n567_, new_new_n568_,
    new_new_n569_, new_new_n570_, new_new_n571_, new_new_n572_,
    new_new_n573_, new_new_n574_, new_new_n575_, new_new_n576_,
    new_new_n577_, new_new_n578_, new_new_n579_, new_new_n580_,
    new_new_n581_, new_new_n582_, new_new_n583_, new_new_n584_,
    new_new_n585_, new_new_n586_, new_new_n587_, new_new_n588_,
    new_new_n589_, new_new_n590_, new_new_n591_, new_new_n592_,
    new_new_n593_, new_new_n594_, new_new_n595_, new_new_n596_,
    new_new_n597_, new_new_n598_, new_new_n599_, new_new_n600_,
    new_new_n601_, new_new_n602_, new_new_n603_, new_new_n604_,
    new_new_n605_, new_new_n606_, new_new_n607_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n625_,
    new_new_n626_, new_new_n627_, new_new_n628_, new_new_n629_,
    new_new_n630_, new_new_n631_, new_new_n632_, new_new_n633_,
    new_new_n634_, new_new_n635_, new_new_n636_, new_new_n637_,
    new_new_n638_, new_new_n639_, new_new_n640_, new_new_n641_,
    new_new_n642_, new_new_n643_, new_new_n644_, new_new_n645_,
    new_new_n646_, new_new_n647_, new_new_n648_, new_new_n649_,
    new_new_n650_, new_new_n651_, new_new_n652_, new_new_n653_,
    new_new_n654_, new_new_n655_, new_new_n656_, new_new_n657_,
    new_new_n658_, new_new_n659_, new_new_n660_, new_new_n661_,
    new_new_n662_, new_new_n663_, new_new_n664_, new_new_n665_,
    new_new_n666_, new_new_n667_, new_new_n668_, new_new_n669_,
    new_new_n670_, new_new_n671_, new_new_n672_, new_new_n673_,
    new_new_n674_, new_new_n675_, new_new_n676_, new_new_n677_,
    new_new_n678_, new_new_n679_, new_new_n680_, new_new_n681_,
    new_new_n682_, new_new_n683_, new_new_n684_, new_new_n685_,
    new_new_n686_, new_new_n687_, new_new_n688_, new_new_n689_,
    new_new_n690_, new_new_n691_, new_new_n692_, new_new_n693_,
    new_new_n694_, new_new_n695_, new_new_n696_, new_new_n697_,
    new_new_n698_, new_new_n699_, new_new_n700_, new_new_n701_,
    new_new_n702_, new_new_n703_, new_new_n704_, new_new_n705_,
    new_new_n706_, new_new_n707_, new_new_n708_, new_new_n709_,
    new_new_n710_, new_new_n711_, new_new_n712_, new_new_n713_,
    new_new_n714_, new_new_n715_, new_new_n716_, new_new_n717_,
    new_new_n718_, new_new_n719_, new_new_n720_, new_new_n721_,
    new_new_n722_, new_new_n723_, new_new_n724_, new_new_n725_,
    new_new_n726_, new_new_n727_, new_new_n728_, new_new_n729_,
    new_new_n730_, new_new_n731_, new_new_n732_, new_new_n733_,
    new_new_n734_, new_new_n735_, new_new_n736_, new_new_n737_,
    new_new_n738_, new_new_n739_, new_new_n740_, new_new_n741_,
    new_new_n742_, new_new_n743_, new_new_n744_, new_new_n745_,
    new_new_n746_, new_new_n747_, new_new_n748_, new_new_n749_,
    new_new_n750_, new_new_n752_, new_new_n753_, new_new_n754_,
    new_new_n755_, new_new_n756_, new_new_n757_, new_new_n758_,
    new_new_n759_, new_new_n760_, new_new_n761_, new_new_n762_,
    new_new_n763_, new_new_n764_, new_new_n765_, new_new_n766_,
    new_new_n767_, new_new_n768_, new_new_n769_, new_new_n770_,
    new_new_n771_, new_new_n772_, new_new_n773_, new_new_n774_,
    new_new_n775_, new_new_n776_, new_new_n777_, new_new_n778_,
    new_new_n779_, new_new_n780_, new_new_n781_, new_new_n782_,
    new_new_n783_, new_new_n784_, new_new_n785_, new_new_n786_,
    new_new_n787_, new_new_n788_, new_new_n789_, new_new_n790_,
    new_new_n791_, new_new_n792_, new_new_n793_, new_new_n794_,
    new_new_n795_, new_new_n796_, new_new_n798_, new_new_n799_,
    new_new_n800_, new_new_n801_, new_new_n802_, new_new_n803_,
    new_new_n804_, new_new_n805_, new_new_n806_, new_new_n807_,
    new_new_n808_, new_new_n809_, new_new_n810_, new_new_n811_,
    new_new_n812_, new_new_n813_, new_new_n814_, new_new_n815_,
    new_new_n816_, new_new_n817_, new_new_n818_, new_new_n819_,
    new_new_n820_, new_new_n821_, new_new_n822_, new_new_n823_,
    new_new_n824_, new_new_n825_, new_new_n826_, new_new_n827_,
    new_new_n828_, new_new_n829_, new_new_n830_, new_new_n831_,
    new_new_n832_, new_new_n833_, new_new_n834_, new_new_n835_,
    new_new_n836_, new_new_n837_, new_new_n838_, new_new_n839_,
    new_new_n840_, new_new_n841_, new_new_n842_, new_new_n843_,
    new_new_n844_, new_new_n845_, new_new_n846_, new_new_n847_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n890_, new_new_n891_, new_new_n892_,
    new_new_n893_, new_new_n894_, new_new_n895_, new_new_n896_,
    new_new_n897_, new_new_n898_, new_new_n899_, new_new_n900_,
    new_new_n901_, new_new_n902_, new_new_n903_, new_new_n904_,
    new_new_n905_, new_new_n906_, new_new_n907_, new_new_n908_,
    new_new_n909_, new_new_n910_, new_new_n911_, new_new_n912_,
    new_new_n913_, new_new_n914_, new_new_n915_, new_new_n916_,
    new_new_n917_, new_new_n918_, new_new_n919_, new_new_n920_,
    new_new_n921_, new_new_n922_, new_new_n923_, new_new_n924_,
    new_new_n925_, new_new_n926_, new_new_n927_, new_new_n928_,
    new_new_n929_, new_new_n930_, new_new_n931_, new_new_n932_,
    new_new_n933_, new_new_n934_, new_new_n935_, new_new_n936_,
    new_new_n937_, new_new_n938_, new_new_n939_, new_new_n940_,
    new_new_n941_, new_new_n942_, new_new_n943_, new_new_n944_,
    new_new_n945_, new_new_n946_, new_new_n947_, new_new_n948_,
    new_new_n949_, new_new_n950_, new_new_n951_, new_new_n952_,
    new_new_n953_, new_new_n954_, new_new_n955_, new_new_n956_,
    new_new_n957_, new_new_n958_, new_new_n959_, new_new_n960_,
    new_new_n961_, new_new_n962_, new_new_n963_, new_new_n964_,
    new_new_n965_, new_new_n966_, new_new_n967_, new_new_n968_,
    new_new_n969_, new_new_n970_, new_new_n971_, new_new_n972_,
    new_new_n973_, new_new_n974_, new_new_n975_, new_new_n976_,
    new_new_n977_, new_new_n978_, new_new_n979_, new_new_n980_,
    new_new_n981_, new_new_n982_, new_new_n983_, new_new_n984_,
    new_new_n985_, new_new_n986_, new_new_n987_, new_new_n988_,
    new_new_n989_, new_new_n990_, new_new_n991_, new_new_n992_,
    new_new_n993_, new_new_n994_, new_new_n995_, new_new_n996_,
    new_new_n997_, new_new_n998_, new_new_n999_, new_new_n1000_,
    new_new_n1001_, new_new_n1002_, new_new_n1003_, new_new_n1004_,
    new_new_n1005_, new_new_n1006_, new_new_n1007_, new_new_n1008_,
    new_new_n1009_, new_new_n1010_, new_new_n1011_, new_new_n1012_,
    new_new_n1013_, new_new_n1014_, new_new_n1015_, new_new_n1016_,
    new_new_n1017_, new_new_n1018_, new_new_n1019_, new_new_n1020_,
    new_new_n1021_, new_new_n1022_, new_new_n1023_, new_new_n1024_,
    new_new_n1025_, new_new_n1026_, new_new_n1027_, new_new_n1028_,
    new_new_n1029_, new_new_n1030_, new_new_n1031_, new_new_n1032_,
    new_new_n1033_, new_new_n1034_, new_new_n1035_, new_new_n1036_,
    new_new_n1037_, new_new_n1038_, new_new_n1039_, new_new_n1040_,
    new_new_n1041_, new_new_n1042_, new_new_n1043_, new_new_n1044_,
    new_new_n1045_, new_new_n1046_, new_new_n1047_, new_new_n1048_,
    new_new_n1049_, new_new_n1050_, new_new_n1051_, new_new_n1052_,
    new_new_n1053_, new_new_n1054_, new_new_n1055_, new_new_n1056_,
    new_new_n1057_, new_new_n1058_, new_new_n1059_, new_new_n1060_,
    new_new_n1061_, new_new_n1062_, new_new_n1063_, new_new_n1064_,
    new_new_n1065_, new_new_n1066_, new_new_n1067_, new_new_n1068_,
    new_new_n1069_, new_new_n1070_, new_new_n1071_, new_new_n1072_,
    new_new_n1073_, new_new_n1077_, new_new_n1078_, new_new_n1079_,
    new_new_n1080_;
  NAi21      g0000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g0001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g0002(.A(i_9_), .Y(new_new_n25_));
  INV        g0003(.A(i_3_), .Y(new_new_n26_));
  NO2        g0004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g0005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g0006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g0007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g0008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g0009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g0010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g0011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g0012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g0013(.A(i_4_), .Y(new_new_n36_));
  INV        g0014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g0015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g0016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g0017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g0018(.A(new_new_n40_), .Y(new_new_n41_));
  NO2        g0019(.A(new_new_n36_), .B(i_3_), .Y(new_new_n42_));
  NAi31      g0020(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n43_));
  INV        g0021(.A(new_new_n35_), .Y(men1));
  INV        g0022(.A(i_11_), .Y(new_new_n45_));
  NO2        g0023(.A(new_new_n45_), .B(i_6_), .Y(new_new_n46_));
  INV        g0024(.A(i_2_), .Y(new_new_n47_));
  NA2        g0025(.A(i_0_), .B(i_3_), .Y(new_new_n48_));
  INV        g0026(.A(i_5_), .Y(new_new_n49_));
  NO2        g0027(.A(i_7_), .B(i_10_), .Y(new_new_n50_));
  AOI210     g0028(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n50_), .Y(new_new_n51_));
  OAI210     g0029(.A0(new_new_n51_), .A1(i_3_), .B0(new_new_n49_), .Y(new_new_n52_));
  AOI210     g0030(.A0(new_new_n52_), .A1(new_new_n48_), .B0(new_new_n47_), .Y(new_new_n53_));
  NA2        g0031(.A(i_0_), .B(i_2_), .Y(new_new_n54_));
  NA2        g0032(.A(i_7_), .B(i_9_), .Y(new_new_n55_));
  NA2        g0033(.A(new_new_n53_), .B(new_new_n46_), .Y(new_new_n56_));
  NA3        g0034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g0035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g0036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g0037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g0038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g0039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g0040(.A(i_1_), .Y(new_new_n63_));
  NA2        g0041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g0042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g0043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g0044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g0045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g0046(.A(new_new_n51_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g0047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g0048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g0049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g0050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g0051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g0052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g0053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g0054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g0055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g0056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g0057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g0058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g0059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g0060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g0061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  INV        g0062(.A(i_6_), .Y(new_new_n85_));
  OR4        g0063(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n86_));
  INV        g0064(.A(new_new_n86_), .Y(new_new_n87_));
  NO2        g0065(.A(i_2_), .B(i_7_), .Y(new_new_n88_));
  NAi21      g0066(.An(i_6_), .B(i_10_), .Y(new_new_n89_));
  NA2        g0067(.A(i_6_), .B(i_9_), .Y(new_new_n90_));
  AOI210     g0068(.A0(new_new_n90_), .A1(new_new_n89_), .B0(new_new_n63_), .Y(new_new_n91_));
  NA2        g0069(.A(i_2_), .B(i_6_), .Y(new_new_n92_));
  INV        g0070(.A(new_new_n91_), .Y(new_new_n93_));
  AOI210     g0071(.A0(new_new_n93_), .A1(new_new_n1078_), .B0(new_new_n80_), .Y(new_new_n94_));
  AN3        g0072(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n95_));
  NAi21      g0073(.An(i_6_), .B(i_11_), .Y(new_new_n96_));
  NO2        g0074(.A(i_5_), .B(i_8_), .Y(new_new_n97_));
  NOi21      g0075(.An(new_new_n97_), .B(new_new_n96_), .Y(new_new_n98_));
  AOI220     g0076(.A0(new_new_n98_), .A1(new_new_n62_), .B0(new_new_n95_), .B1(new_new_n32_), .Y(new_new_n99_));
  INV        g0077(.A(i_7_), .Y(new_new_n100_));
  NA2        g0078(.A(new_new_n47_), .B(new_new_n100_), .Y(new_new_n101_));
  NO2        g0079(.A(i_0_), .B(i_5_), .Y(new_new_n102_));
  NO2        g0080(.A(new_new_n102_), .B(new_new_n85_), .Y(new_new_n103_));
  NA2        g0081(.A(i_12_), .B(i_3_), .Y(new_new_n104_));
  INV        g0082(.A(new_new_n104_), .Y(new_new_n105_));
  NA3        g0083(.A(new_new_n105_), .B(new_new_n103_), .C(new_new_n101_), .Y(new_new_n106_));
  NAi21      g0084(.An(i_7_), .B(i_11_), .Y(new_new_n107_));
  NO3        g0085(.A(new_new_n107_), .B(new_new_n89_), .C(new_new_n54_), .Y(new_new_n108_));
  AN2        g0086(.A(i_2_), .B(i_10_), .Y(new_new_n109_));
  NO2        g0087(.A(new_new_n109_), .B(i_7_), .Y(new_new_n110_));
  OR2        g0088(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n111_));
  NO2        g0089(.A(i_8_), .B(new_new_n100_), .Y(new_new_n112_));
  NO3        g0090(.A(new_new_n112_), .B(new_new_n111_), .C(new_new_n110_), .Y(new_new_n113_));
  NA2        g0091(.A(i_12_), .B(i_7_), .Y(new_new_n114_));
  NO2        g0092(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n115_));
  NA2        g0093(.A(new_new_n115_), .B(i_0_), .Y(new_new_n116_));
  NA2        g0094(.A(i_11_), .B(i_12_), .Y(new_new_n117_));
  OAI210     g0095(.A0(new_new_n116_), .A1(new_new_n114_), .B0(new_new_n117_), .Y(new_new_n118_));
  NO2        g0096(.A(new_new_n118_), .B(new_new_n113_), .Y(new_new_n119_));
  NAi41      g0097(.An(new_new_n108_), .B(new_new_n119_), .C(new_new_n106_), .D(new_new_n99_), .Y(new_new_n120_));
  NOi21      g0098(.An(i_1_), .B(i_5_), .Y(new_new_n121_));
  NA2        g0099(.A(new_new_n121_), .B(i_11_), .Y(new_new_n122_));
  NA2        g0100(.A(new_new_n100_), .B(new_new_n37_), .Y(new_new_n123_));
  NA2        g0101(.A(i_7_), .B(new_new_n25_), .Y(new_new_n124_));
  NA2        g0102(.A(new_new_n124_), .B(new_new_n123_), .Y(new_new_n125_));
  NO2        g0103(.A(new_new_n125_), .B(new_new_n47_), .Y(new_new_n126_));
  NA2        g0104(.A(new_new_n90_), .B(new_new_n89_), .Y(new_new_n127_));
  NAi21      g0105(.An(i_3_), .B(i_8_), .Y(new_new_n128_));
  NA2        g0106(.A(new_new_n128_), .B(new_new_n62_), .Y(new_new_n129_));
  NOi31      g0107(.An(new_new_n129_), .B(new_new_n127_), .C(new_new_n126_), .Y(new_new_n130_));
  NO2        g0108(.A(i_1_), .B(new_new_n85_), .Y(new_new_n131_));
  NO2        g0109(.A(i_6_), .B(i_5_), .Y(new_new_n132_));
  NA2        g0110(.A(new_new_n132_), .B(i_3_), .Y(new_new_n133_));
  AO210      g0111(.A0(new_new_n133_), .A1(new_new_n48_), .B0(new_new_n131_), .Y(new_new_n134_));
  OAI220     g0112(.A0(new_new_n134_), .A1(new_new_n107_), .B0(new_new_n130_), .B1(new_new_n122_), .Y(new_new_n135_));
  NO3        g0113(.A(new_new_n135_), .B(new_new_n120_), .C(new_new_n94_), .Y(new_new_n136_));
  NA3        g0114(.A(new_new_n136_), .B(new_new_n79_), .C(new_new_n56_), .Y(men2));
  NO2        g0115(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n138_));
  NA2        g0116(.A(i_6_), .B(new_new_n25_), .Y(new_new_n139_));
  NA2        g0117(.A(new_new_n139_), .B(new_new_n138_), .Y(new_new_n140_));
  NA4        g0118(.A(new_new_n140_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(men0));
  AN2        g0119(.A(i_8_), .B(i_7_), .Y(new_new_n142_));
  NA2        g0120(.A(new_new_n142_), .B(i_6_), .Y(new_new_n143_));
  NO2        g0121(.A(i_12_), .B(i_13_), .Y(new_new_n144_));
  NAi21      g0122(.An(i_5_), .B(i_11_), .Y(new_new_n145_));
  NOi21      g0123(.An(new_new_n144_), .B(new_new_n145_), .Y(new_new_n146_));
  NO2        g0124(.A(i_0_), .B(i_1_), .Y(new_new_n147_));
  NA2        g0125(.A(i_2_), .B(i_3_), .Y(new_new_n148_));
  NA3        g0126(.A(i_3_), .B(new_new_n147_), .C(new_new_n146_), .Y(new_new_n149_));
  OR2        g0127(.A(new_new_n149_), .B(new_new_n25_), .Y(new_new_n150_));
  AN2        g0128(.A(new_new_n144_), .B(new_new_n83_), .Y(new_new_n151_));
  NO2        g0129(.A(new_new_n151_), .B(new_new_n27_), .Y(new_new_n152_));
  NA2        g0130(.A(i_1_), .B(i_5_), .Y(new_new_n153_));
  NO2        g0131(.A(new_new_n73_), .B(new_new_n47_), .Y(new_new_n154_));
  NA2        g0132(.A(new_new_n154_), .B(new_new_n36_), .Y(new_new_n155_));
  NO3        g0133(.A(new_new_n155_), .B(new_new_n153_), .C(new_new_n152_), .Y(new_new_n156_));
  OR2        g0134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g0135(.A(new_new_n157_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g0136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g0137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g0138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g0139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO2        g0140(.A(i_3_), .B(i_5_), .Y(new_new_n163_));
  NO3        g0141(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n164_));
  NA2        g0142(.A(new_new_n164_), .B(new_new_n163_), .Y(new_new_n165_));
  OAI210     g0143(.A0(new_new_n165_), .A1(new_new_n162_), .B0(new_new_n160_), .Y(new_new_n166_));
  NO2        g0144(.A(new_new_n166_), .B(new_new_n156_), .Y(new_new_n167_));
  AOI210     g0145(.A0(new_new_n167_), .A1(new_new_n150_), .B0(new_new_n143_), .Y(new_new_n168_));
  NA3        g0146(.A(new_new_n73_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n169_));
  NOi21      g0147(.An(i_4_), .B(i_9_), .Y(new_new_n170_));
  NOi21      g0148(.An(i_11_), .B(i_13_), .Y(new_new_n171_));
  NA2        g0149(.A(new_new_n171_), .B(new_new_n170_), .Y(new_new_n172_));
  NO2        g0150(.A(i_4_), .B(i_5_), .Y(new_new_n173_));
  NAi21      g0151(.An(i_12_), .B(i_11_), .Y(new_new_n174_));
  NO2        g0152(.A(new_new_n174_), .B(i_13_), .Y(new_new_n175_));
  NA3        g0153(.A(new_new_n175_), .B(new_new_n173_), .C(new_new_n83_), .Y(new_new_n176_));
  AOI210     g0154(.A0(new_new_n176_), .A1(new_new_n172_), .B0(new_new_n169_), .Y(new_new_n177_));
  NO2        g0155(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n178_));
  NA2        g0156(.A(new_new_n178_), .B(new_new_n47_), .Y(new_new_n179_));
  NA2        g0157(.A(new_new_n36_), .B(i_5_), .Y(new_new_n180_));
  NAi31      g0158(.An(new_new_n180_), .B(new_new_n151_), .C(i_11_), .Y(new_new_n181_));
  NA2        g0159(.A(i_3_), .B(i_5_), .Y(new_new_n182_));
  OR2        g0160(.A(new_new_n182_), .B(new_new_n172_), .Y(new_new_n183_));
  AOI210     g0161(.A0(new_new_n183_), .A1(new_new_n181_), .B0(new_new_n179_), .Y(new_new_n184_));
  NO2        g0162(.A(new_new_n73_), .B(i_5_), .Y(new_new_n185_));
  NO2        g0163(.A(i_13_), .B(i_10_), .Y(new_new_n186_));
  NA3        g0164(.A(new_new_n186_), .B(new_new_n185_), .C(new_new_n45_), .Y(new_new_n187_));
  NO2        g0165(.A(i_2_), .B(i_1_), .Y(new_new_n188_));
  NA2        g0166(.A(new_new_n188_), .B(i_3_), .Y(new_new_n189_));
  NAi21      g0167(.An(i_4_), .B(i_12_), .Y(new_new_n190_));
  NO4        g0168(.A(new_new_n190_), .B(new_new_n189_), .C(new_new_n187_), .D(new_new_n25_), .Y(new_new_n191_));
  NO3        g0169(.A(new_new_n191_), .B(new_new_n184_), .C(new_new_n177_), .Y(new_new_n192_));
  INV        g0170(.A(i_8_), .Y(new_new_n193_));
  NO2        g0171(.A(new_new_n193_), .B(i_7_), .Y(new_new_n194_));
  NA2        g0172(.A(new_new_n194_), .B(i_6_), .Y(new_new_n195_));
  NO3        g0173(.A(i_3_), .B(new_new_n85_), .C(new_new_n49_), .Y(new_new_n196_));
  NA2        g0174(.A(new_new_n196_), .B(new_new_n112_), .Y(new_new_n197_));
  NO3        g0175(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n198_));
  NA3        g0176(.A(new_new_n198_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n199_));
  NO3        g0177(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n200_));
  OAI210     g0178(.A0(new_new_n95_), .A1(i_12_), .B0(new_new_n200_), .Y(new_new_n201_));
  AOI210     g0179(.A0(new_new_n201_), .A1(new_new_n199_), .B0(new_new_n197_), .Y(new_new_n202_));
  NO2        g0180(.A(i_3_), .B(i_8_), .Y(new_new_n203_));
  NO3        g0181(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n204_));
  NA3        g0182(.A(new_new_n204_), .B(new_new_n203_), .C(new_new_n40_), .Y(new_new_n205_));
  NO2        g0183(.A(new_new_n102_), .B(new_new_n58_), .Y(new_new_n206_));
  NO2        g0184(.A(i_13_), .B(i_9_), .Y(new_new_n207_));
  NA3        g0185(.A(new_new_n207_), .B(i_6_), .C(new_new_n193_), .Y(new_new_n208_));
  NAi21      g0186(.An(i_12_), .B(i_3_), .Y(new_new_n209_));
  OR2        g0187(.A(new_new_n209_), .B(new_new_n208_), .Y(new_new_n210_));
  NO2        g0188(.A(new_new_n45_), .B(i_5_), .Y(new_new_n211_));
  NO3        g0189(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n212_));
  INV        g0190(.A(new_new_n212_), .Y(new_new_n213_));
  OAI220     g0191(.A0(new_new_n213_), .A1(new_new_n210_), .B0(new_new_n102_), .B1(new_new_n205_), .Y(new_new_n214_));
  AOI210     g0192(.A0(new_new_n214_), .A1(i_7_), .B0(new_new_n202_), .Y(new_new_n215_));
  OAI220     g0193(.A0(new_new_n215_), .A1(i_4_), .B0(new_new_n195_), .B1(new_new_n192_), .Y(new_new_n216_));
  NAi21      g0194(.An(i_12_), .B(i_7_), .Y(new_new_n217_));
  NA3        g0195(.A(i_13_), .B(new_new_n193_), .C(i_10_), .Y(new_new_n218_));
  NO2        g0196(.A(new_new_n218_), .B(new_new_n217_), .Y(new_new_n219_));
  NA2        g0197(.A(i_0_), .B(i_5_), .Y(new_new_n220_));
  OAI220     g0198(.A0(new_new_n85_), .A1(new_new_n189_), .B0(new_new_n179_), .B1(new_new_n133_), .Y(new_new_n221_));
  NAi31      g0199(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n222_));
  NO2        g0200(.A(new_new_n36_), .B(i_13_), .Y(new_new_n223_));
  NO2        g0201(.A(new_new_n47_), .B(new_new_n63_), .Y(new_new_n224_));
  NA3        g0202(.A(new_new_n224_), .B(i_0_), .C(new_new_n223_), .Y(new_new_n225_));
  INV        g0203(.A(i_13_), .Y(new_new_n226_));
  NO2        g0204(.A(i_12_), .B(new_new_n226_), .Y(new_new_n227_));
  NA3        g0205(.A(new_new_n227_), .B(new_new_n198_), .C(new_new_n196_), .Y(new_new_n228_));
  OAI210     g0206(.A0(new_new_n225_), .A1(new_new_n222_), .B0(new_new_n228_), .Y(new_new_n229_));
  AOI220     g0207(.A0(new_new_n229_), .A1(new_new_n142_), .B0(new_new_n221_), .B1(new_new_n219_), .Y(new_new_n230_));
  NO2        g0208(.A(i_12_), .B(new_new_n37_), .Y(new_new_n231_));
  NO2        g0209(.A(new_new_n182_), .B(i_4_), .Y(new_new_n232_));
  NA2        g0210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  OR2        g0211(.A(i_8_), .B(i_7_), .Y(new_new_n234_));
  NO2        g0212(.A(new_new_n234_), .B(new_new_n85_), .Y(new_new_n235_));
  NO2        g0213(.A(new_new_n54_), .B(i_1_), .Y(new_new_n236_));
  NA2        g0214(.A(new_new_n236_), .B(new_new_n235_), .Y(new_new_n237_));
  INV        g0215(.A(i_12_), .Y(new_new_n238_));
  NO2        g0216(.A(new_new_n45_), .B(new_new_n238_), .Y(new_new_n239_));
  NO3        g0217(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n240_));
  NA2        g0218(.A(i_2_), .B(i_1_), .Y(new_new_n241_));
  NO2        g0219(.A(new_new_n237_), .B(new_new_n233_), .Y(new_new_n242_));
  NO3        g0220(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n243_));
  NAi21      g0221(.An(i_4_), .B(i_3_), .Y(new_new_n244_));
  NO2        g0222(.A(new_new_n244_), .B(new_new_n75_), .Y(new_new_n245_));
  NO2        g0223(.A(i_0_), .B(i_6_), .Y(new_new_n246_));
  NOi41      g0224(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n247_));
  NA2        g0225(.A(new_new_n247_), .B(new_new_n246_), .Y(new_new_n248_));
  NO2        g0226(.A(new_new_n241_), .B(new_new_n182_), .Y(new_new_n249_));
  NAi21      g0227(.An(new_new_n248_), .B(new_new_n249_), .Y(new_new_n250_));
  INV        g0228(.A(new_new_n250_), .Y(new_new_n251_));
  AOI220     g0229(.A0(new_new_n251_), .A1(new_new_n40_), .B0(new_new_n242_), .B1(new_new_n207_), .Y(new_new_n252_));
  NO2        g0230(.A(i_11_), .B(new_new_n226_), .Y(new_new_n253_));
  NOi21      g0231(.An(i_1_), .B(i_6_), .Y(new_new_n254_));
  NAi21      g0232(.An(i_3_), .B(i_7_), .Y(new_new_n255_));
  NO2        g0233(.A(new_new_n49_), .B(new_new_n25_), .Y(new_new_n256_));
  NO2        g0234(.A(i_12_), .B(i_3_), .Y(new_new_n257_));
  NA2        g0235(.A(i_3_), .B(i_9_), .Y(new_new_n258_));
  NA3        g0236(.A(i_1_), .B(i_8_), .C(i_7_), .Y(new_new_n259_));
  INV        g0237(.A(new_new_n143_), .Y(new_new_n260_));
  NA2        g0238(.A(new_new_n238_), .B(i_13_), .Y(new_new_n261_));
  NO2        g0239(.A(new_new_n261_), .B(new_new_n75_), .Y(new_new_n262_));
  NA2        g0240(.A(new_new_n262_), .B(new_new_n260_), .Y(new_new_n263_));
  NO2        g0241(.A(new_new_n234_), .B(new_new_n37_), .Y(new_new_n264_));
  NA2        g0242(.A(i_12_), .B(i_6_), .Y(new_new_n265_));
  OR2        g0243(.A(i_13_), .B(i_9_), .Y(new_new_n266_));
  NO3        g0244(.A(new_new_n266_), .B(new_new_n265_), .C(new_new_n49_), .Y(new_new_n267_));
  NO2        g0245(.A(new_new_n244_), .B(i_2_), .Y(new_new_n268_));
  NA3        g0246(.A(new_new_n268_), .B(new_new_n267_), .C(new_new_n45_), .Y(new_new_n269_));
  NA2        g0247(.A(new_new_n253_), .B(i_9_), .Y(new_new_n270_));
  NA2        g0248(.A(i_0_), .B(new_new_n64_), .Y(new_new_n271_));
  OAI210     g0249(.A0(new_new_n271_), .A1(new_new_n270_), .B0(new_new_n269_), .Y(new_new_n272_));
  NA2        g0250(.A(new_new_n154_), .B(new_new_n63_), .Y(new_new_n273_));
  NO3        g0251(.A(i_11_), .B(new_new_n226_), .C(new_new_n25_), .Y(new_new_n274_));
  NO2        g0252(.A(new_new_n255_), .B(i_8_), .Y(new_new_n275_));
  NO2        g0253(.A(i_6_), .B(new_new_n49_), .Y(new_new_n276_));
  NA3        g0254(.A(new_new_n276_), .B(new_new_n275_), .C(new_new_n274_), .Y(new_new_n277_));
  NO3        g0255(.A(new_new_n26_), .B(new_new_n85_), .C(i_5_), .Y(new_new_n278_));
  NA3        g0256(.A(new_new_n278_), .B(new_new_n264_), .C(new_new_n227_), .Y(new_new_n279_));
  AOI210     g0257(.A0(new_new_n279_), .A1(new_new_n277_), .B0(new_new_n273_), .Y(new_new_n280_));
  AOI210     g0258(.A0(new_new_n272_), .A1(new_new_n264_), .B0(new_new_n280_), .Y(new_new_n281_));
  NA4        g0259(.A(new_new_n281_), .B(new_new_n263_), .C(new_new_n252_), .D(new_new_n230_), .Y(new_new_n282_));
  NO3        g0260(.A(i_12_), .B(new_new_n226_), .C(new_new_n37_), .Y(new_new_n283_));
  INV        g0261(.A(new_new_n283_), .Y(new_new_n284_));
  NA2        g0262(.A(i_8_), .B(new_new_n100_), .Y(new_new_n285_));
  NO3        g0263(.A(i_0_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n286_));
  AOI220     g0264(.A0(new_new_n286_), .A1(new_new_n196_), .B0(new_new_n163_), .B1(new_new_n236_), .Y(new_new_n287_));
  NO2        g0265(.A(new_new_n287_), .B(new_new_n285_), .Y(new_new_n288_));
  NO3        g0266(.A(i_0_), .B(i_2_), .C(new_new_n63_), .Y(new_new_n289_));
  NO2        g0267(.A(new_new_n241_), .B(i_0_), .Y(new_new_n290_));
  AOI220     g0268(.A0(new_new_n290_), .A1(new_new_n194_), .B0(new_new_n289_), .B1(new_new_n142_), .Y(new_new_n291_));
  NA2        g0269(.A(new_new_n276_), .B(new_new_n26_), .Y(new_new_n292_));
  NO2        g0270(.A(new_new_n292_), .B(new_new_n291_), .Y(new_new_n293_));
  NA2        g0271(.A(i_0_), .B(i_1_), .Y(new_new_n294_));
  NO2        g0272(.A(new_new_n294_), .B(i_2_), .Y(new_new_n295_));
  NO2        g0273(.A(new_new_n59_), .B(i_6_), .Y(new_new_n296_));
  NA3        g0274(.A(new_new_n296_), .B(new_new_n295_), .C(new_new_n163_), .Y(new_new_n297_));
  OAI210     g0275(.A0(new_new_n165_), .A1(new_new_n143_), .B0(new_new_n297_), .Y(new_new_n298_));
  NO3        g0276(.A(new_new_n298_), .B(new_new_n293_), .C(new_new_n288_), .Y(new_new_n299_));
  NO2        g0277(.A(i_3_), .B(i_10_), .Y(new_new_n300_));
  NA3        g0278(.A(new_new_n300_), .B(new_new_n40_), .C(new_new_n45_), .Y(new_new_n301_));
  NO2        g0279(.A(i_2_), .B(new_new_n100_), .Y(new_new_n302_));
  NA2        g0280(.A(i_1_), .B(new_new_n36_), .Y(new_new_n303_));
  NOi21      g0281(.An(new_new_n220_), .B(new_new_n102_), .Y(new_new_n304_));
  NA3        g0282(.A(new_new_n304_), .B(i_1_), .C(new_new_n302_), .Y(new_new_n305_));
  AN2        g0283(.A(i_3_), .B(i_10_), .Y(new_new_n306_));
  NA4        g0284(.A(new_new_n306_), .B(new_new_n198_), .C(new_new_n175_), .D(new_new_n173_), .Y(new_new_n307_));
  NO2        g0285(.A(i_5_), .B(new_new_n37_), .Y(new_new_n308_));
  NO2        g0286(.A(new_new_n47_), .B(new_new_n26_), .Y(new_new_n309_));
  OR2        g0287(.A(new_new_n305_), .B(new_new_n301_), .Y(new_new_n310_));
  OAI220     g0288(.A0(new_new_n310_), .A1(i_6_), .B0(new_new_n299_), .B1(new_new_n284_), .Y(new_new_n311_));
  NO4        g0289(.A(new_new_n311_), .B(new_new_n282_), .C(new_new_n216_), .D(new_new_n168_), .Y(new_new_n312_));
  NO3        g0290(.A(new_new_n45_), .B(i_13_), .C(i_9_), .Y(new_new_n313_));
  NO2        g0291(.A(new_new_n59_), .B(new_new_n85_), .Y(new_new_n314_));
  NA2        g0292(.A(new_new_n290_), .B(new_new_n314_), .Y(new_new_n315_));
  NO3        g0293(.A(i_6_), .B(new_new_n193_), .C(i_7_), .Y(new_new_n316_));
  NA2        g0294(.A(new_new_n316_), .B(new_new_n198_), .Y(new_new_n317_));
  AOI210     g0295(.A0(new_new_n317_), .A1(new_new_n315_), .B0(i_5_), .Y(new_new_n318_));
  NO2        g0296(.A(i_2_), .B(i_3_), .Y(new_new_n319_));
  OR2        g0297(.A(i_0_), .B(i_5_), .Y(new_new_n320_));
  NA2        g0298(.A(new_new_n220_), .B(new_new_n320_), .Y(new_new_n321_));
  NA4        g0299(.A(new_new_n321_), .B(new_new_n235_), .C(new_new_n319_), .D(i_1_), .Y(new_new_n322_));
  NA3        g0300(.A(new_new_n290_), .B(new_new_n163_), .C(new_new_n112_), .Y(new_new_n323_));
  NO2        g0301(.A(i_8_), .B(i_6_), .Y(new_new_n324_));
  NO2        g0302(.A(new_new_n157_), .B(new_new_n47_), .Y(new_new_n325_));
  NA3        g0303(.A(new_new_n325_), .B(new_new_n324_), .C(new_new_n163_), .Y(new_new_n326_));
  NA3        g0304(.A(new_new_n326_), .B(new_new_n323_), .C(new_new_n322_), .Y(new_new_n327_));
  OAI210     g0305(.A0(new_new_n327_), .A1(new_new_n318_), .B0(i_4_), .Y(new_new_n328_));
  NO2        g0306(.A(i_12_), .B(i_10_), .Y(new_new_n329_));
  NOi21      g0307(.An(i_5_), .B(i_0_), .Y(new_new_n330_));
  NO3        g0308(.A(new_new_n303_), .B(new_new_n330_), .C(new_new_n128_), .Y(new_new_n331_));
  NA4        g0309(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n85_), .D(i_8_), .Y(new_new_n332_));
  NA2        g0310(.A(new_new_n331_), .B(new_new_n329_), .Y(new_new_n333_));
  NO2        g0311(.A(i_6_), .B(i_8_), .Y(new_new_n334_));
  NOi21      g0312(.An(i_0_), .B(i_2_), .Y(new_new_n335_));
  AN2        g0313(.A(new_new_n335_), .B(new_new_n334_), .Y(new_new_n336_));
  NO2        g0314(.A(i_1_), .B(i_7_), .Y(new_new_n337_));
  AO220      g0315(.A0(new_new_n337_), .A1(new_new_n336_), .B0(new_new_n324_), .B1(new_new_n236_), .Y(new_new_n338_));
  NA2        g0316(.A(new_new_n338_), .B(new_new_n42_), .Y(new_new_n339_));
  NA3        g0317(.A(new_new_n339_), .B(new_new_n333_), .C(new_new_n328_), .Y(new_new_n340_));
  NO3        g0318(.A(new_new_n234_), .B(new_new_n47_), .C(i_1_), .Y(new_new_n341_));
  NO3        g0319(.A(i_8_), .B(i_2_), .C(i_1_), .Y(new_new_n342_));
  OAI210     g0320(.A0(new_new_n342_), .A1(new_new_n341_), .B0(i_6_), .Y(new_new_n343_));
  NA3        g0321(.A(new_new_n254_), .B(new_new_n302_), .C(new_new_n193_), .Y(new_new_n344_));
  AOI210     g0322(.A0(new_new_n344_), .A1(new_new_n343_), .B0(new_new_n321_), .Y(new_new_n345_));
  NA2        g0323(.A(new_new_n345_), .B(i_3_), .Y(new_new_n346_));
  INV        g0324(.A(new_new_n84_), .Y(new_new_n347_));
  NO2        g0325(.A(new_new_n294_), .B(new_new_n81_), .Y(new_new_n348_));
  NA2        g0326(.A(new_new_n348_), .B(new_new_n132_), .Y(new_new_n349_));
  NO2        g0327(.A(new_new_n92_), .B(new_new_n193_), .Y(new_new_n350_));
  NA3        g0328(.A(new_new_n304_), .B(new_new_n350_), .C(new_new_n63_), .Y(new_new_n351_));
  AOI210     g0329(.A0(new_new_n351_), .A1(new_new_n349_), .B0(new_new_n347_), .Y(new_new_n352_));
  NO2        g0330(.A(new_new_n193_), .B(i_9_), .Y(new_new_n353_));
  NA2        g0331(.A(new_new_n353_), .B(new_new_n206_), .Y(new_new_n354_));
  NO2        g0332(.A(new_new_n352_), .B(new_new_n293_), .Y(new_new_n355_));
  AOI210     g0333(.A0(new_new_n355_), .A1(new_new_n346_), .B0(new_new_n162_), .Y(new_new_n356_));
  AOI210     g0334(.A0(new_new_n340_), .A1(new_new_n313_), .B0(new_new_n356_), .Y(new_new_n357_));
  NOi32      g0335(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n358_));
  INV        g0336(.A(new_new_n358_), .Y(new_new_n359_));
  NAi21      g0337(.An(i_0_), .B(i_6_), .Y(new_new_n360_));
  NAi21      g0338(.An(i_1_), .B(i_5_), .Y(new_new_n361_));
  NA2        g0339(.A(new_new_n361_), .B(new_new_n360_), .Y(new_new_n362_));
  NAi41      g0340(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n363_));
  OAI220     g0341(.A0(new_new_n363_), .A1(new_new_n361_), .B0(new_new_n222_), .B1(new_new_n159_), .Y(new_new_n364_));
  AOI210     g0342(.A0(new_new_n363_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n365_));
  NOi32      g0343(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n366_));
  NAi21      g0344(.An(i_6_), .B(i_1_), .Y(new_new_n367_));
  NA3        g0345(.A(new_new_n367_), .B(new_new_n366_), .C(new_new_n47_), .Y(new_new_n368_));
  NO2        g0346(.A(new_new_n368_), .B(i_0_), .Y(new_new_n369_));
  OR3        g0347(.A(new_new_n369_), .B(new_new_n365_), .C(new_new_n364_), .Y(new_new_n370_));
  NO2        g0348(.A(i_1_), .B(new_new_n100_), .Y(new_new_n371_));
  NAi21      g0349(.An(i_3_), .B(i_4_), .Y(new_new_n372_));
  NO2        g0350(.A(new_new_n372_), .B(i_9_), .Y(new_new_n373_));
  AN2        g0351(.A(i_6_), .B(i_7_), .Y(new_new_n374_));
  OAI210     g0352(.A0(new_new_n374_), .A1(new_new_n371_), .B0(new_new_n373_), .Y(new_new_n375_));
  NA2        g0353(.A(i_2_), .B(i_7_), .Y(new_new_n376_));
  NO2        g0354(.A(new_new_n372_), .B(i_10_), .Y(new_new_n377_));
  NA3        g0355(.A(new_new_n377_), .B(new_new_n376_), .C(new_new_n246_), .Y(new_new_n378_));
  AOI210     g0356(.A0(new_new_n378_), .A1(new_new_n375_), .B0(new_new_n185_), .Y(new_new_n379_));
  AOI210     g0357(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n380_));
  AOI220     g0358(.A0(new_new_n377_), .A1(new_new_n337_), .B0(new_new_n240_), .B1(new_new_n188_), .Y(new_new_n381_));
  NO2        g0359(.A(new_new_n381_), .B(i_5_), .Y(new_new_n382_));
  NO3        g0360(.A(new_new_n382_), .B(new_new_n379_), .C(new_new_n370_), .Y(new_new_n383_));
  NO2        g0361(.A(new_new_n383_), .B(new_new_n359_), .Y(new_new_n384_));
  NO2        g0362(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n385_));
  AN2        g0363(.A(i_12_), .B(i_5_), .Y(new_new_n386_));
  NO2        g0364(.A(i_4_), .B(new_new_n26_), .Y(new_new_n387_));
  NA2        g0365(.A(new_new_n387_), .B(new_new_n386_), .Y(new_new_n388_));
  NO2        g0366(.A(i_11_), .B(i_6_), .Y(new_new_n389_));
  NA3        g0367(.A(new_new_n389_), .B(new_new_n325_), .C(new_new_n226_), .Y(new_new_n390_));
  NO2        g0368(.A(new_new_n390_), .B(new_new_n388_), .Y(new_new_n391_));
  NO2        g0369(.A(new_new_n244_), .B(i_5_), .Y(new_new_n392_));
  NO2        g0370(.A(i_5_), .B(i_10_), .Y(new_new_n393_));
  AOI220     g0371(.A0(new_new_n393_), .A1(new_new_n268_), .B0(new_new_n392_), .B1(new_new_n198_), .Y(new_new_n394_));
  NA2        g0372(.A(new_new_n144_), .B(new_new_n46_), .Y(new_new_n395_));
  NO2        g0373(.A(new_new_n395_), .B(new_new_n394_), .Y(new_new_n396_));
  OAI210     g0374(.A0(new_new_n396_), .A1(new_new_n391_), .B0(new_new_n385_), .Y(new_new_n397_));
  NO2        g0375(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n398_));
  NO2        g0376(.A(new_new_n149_), .B(new_new_n85_), .Y(new_new_n399_));
  OAI210     g0377(.A0(new_new_n399_), .A1(new_new_n391_), .B0(new_new_n398_), .Y(new_new_n400_));
  NO3        g0378(.A(new_new_n85_), .B(new_new_n49_), .C(i_9_), .Y(new_new_n401_));
  NO2        g0379(.A(i_3_), .B(new_new_n100_), .Y(new_new_n402_));
  NO2        g0380(.A(i_11_), .B(i_12_), .Y(new_new_n403_));
  NA2        g0381(.A(new_new_n393_), .B(new_new_n238_), .Y(new_new_n404_));
  NA2        g0382(.A(new_new_n42_), .B(i_11_), .Y(new_new_n405_));
  OAI220     g0383(.A0(new_new_n405_), .A1(new_new_n222_), .B0(new_new_n404_), .B1(new_new_n332_), .Y(new_new_n406_));
  NAi21      g0384(.An(i_13_), .B(i_0_), .Y(new_new_n407_));
  NO2        g0385(.A(new_new_n407_), .B(new_new_n241_), .Y(new_new_n408_));
  NA2        g0386(.A(new_new_n406_), .B(new_new_n408_), .Y(new_new_n409_));
  NA3        g0387(.A(new_new_n409_), .B(new_new_n400_), .C(new_new_n397_), .Y(new_new_n410_));
  NO3        g0388(.A(i_1_), .B(i_12_), .C(new_new_n85_), .Y(new_new_n411_));
  NO2        g0389(.A(i_0_), .B(i_11_), .Y(new_new_n412_));
  AN2        g0390(.A(i_1_), .B(i_6_), .Y(new_new_n413_));
  NOi21      g0391(.An(i_2_), .B(i_12_), .Y(new_new_n414_));
  NA2        g0392(.A(new_new_n414_), .B(new_new_n413_), .Y(new_new_n415_));
  INV        g0393(.A(new_new_n415_), .Y(new_new_n416_));
  NA2        g0394(.A(new_new_n142_), .B(i_9_), .Y(new_new_n417_));
  NO2        g0395(.A(new_new_n417_), .B(i_4_), .Y(new_new_n418_));
  NA2        g0396(.A(new_new_n416_), .B(new_new_n418_), .Y(new_new_n419_));
  NAi21      g0397(.An(i_9_), .B(i_4_), .Y(new_new_n420_));
  OR2        g0398(.A(i_13_), .B(i_10_), .Y(new_new_n421_));
  NO2        g0399(.A(new_new_n172_), .B(new_new_n123_), .Y(new_new_n422_));
  BUFFER     g0400(.A(new_new_n218_), .Y(new_new_n423_));
  NO2        g0401(.A(new_new_n100_), .B(new_new_n25_), .Y(new_new_n424_));
  NA2        g0402(.A(new_new_n276_), .B(new_new_n212_), .Y(new_new_n425_));
  NO2        g0403(.A(new_new_n425_), .B(new_new_n423_), .Y(new_new_n426_));
  INV        g0404(.A(new_new_n426_), .Y(new_new_n427_));
  AOI210     g0405(.A0(new_new_n427_), .A1(new_new_n419_), .B0(new_new_n26_), .Y(new_new_n428_));
  NA2        g0406(.A(new_new_n323_), .B(new_new_n322_), .Y(new_new_n429_));
  AOI220     g0407(.A0(new_new_n296_), .A1(new_new_n286_), .B0(new_new_n290_), .B1(new_new_n314_), .Y(new_new_n430_));
  NO2        g0408(.A(new_new_n430_), .B(i_5_), .Y(new_new_n431_));
  NO2        g0409(.A(new_new_n182_), .B(new_new_n85_), .Y(new_new_n432_));
  AOI220     g0410(.A0(new_new_n432_), .A1(new_new_n295_), .B0(new_new_n278_), .B1(new_new_n212_), .Y(new_new_n433_));
  NO2        g0411(.A(new_new_n433_), .B(new_new_n285_), .Y(new_new_n434_));
  NO3        g0412(.A(new_new_n434_), .B(new_new_n431_), .C(new_new_n429_), .Y(new_new_n435_));
  NA2        g0413(.A(new_new_n196_), .B(new_new_n95_), .Y(new_new_n436_));
  NA3        g0414(.A(new_new_n325_), .B(new_new_n163_), .C(new_new_n85_), .Y(new_new_n437_));
  AOI210     g0415(.A0(new_new_n437_), .A1(new_new_n436_), .B0(i_8_), .Y(new_new_n438_));
  NA2        g0416(.A(new_new_n296_), .B(new_new_n236_), .Y(new_new_n439_));
  NO2        g0417(.A(new_new_n439_), .B(new_new_n182_), .Y(new_new_n440_));
  NO2        g0418(.A(i_3_), .B(new_new_n49_), .Y(new_new_n441_));
  NA3        g0419(.A(new_new_n337_), .B(new_new_n336_), .C(new_new_n441_), .Y(new_new_n442_));
  INV        g0420(.A(new_new_n316_), .Y(new_new_n443_));
  OAI210     g0421(.A0(new_new_n443_), .A1(new_new_n189_), .B0(new_new_n442_), .Y(new_new_n444_));
  NO3        g0422(.A(new_new_n444_), .B(new_new_n440_), .C(new_new_n438_), .Y(new_new_n445_));
  AOI210     g0423(.A0(new_new_n445_), .A1(new_new_n435_), .B0(new_new_n270_), .Y(new_new_n446_));
  NO4        g0424(.A(new_new_n446_), .B(new_new_n428_), .C(new_new_n410_), .D(new_new_n384_), .Y(new_new_n447_));
  NO2        g0425(.A(new_new_n63_), .B(i_4_), .Y(new_new_n448_));
  NO2        g0426(.A(new_new_n73_), .B(i_13_), .Y(new_new_n449_));
  NA3        g0427(.A(new_new_n449_), .B(new_new_n448_), .C(i_2_), .Y(new_new_n450_));
  NO2        g0428(.A(i_10_), .B(i_9_), .Y(new_new_n451_));
  NAi21      g0429(.An(i_12_), .B(i_8_), .Y(new_new_n452_));
  NO2        g0430(.A(new_new_n452_), .B(i_3_), .Y(new_new_n453_));
  NA2        g0431(.A(new_new_n453_), .B(new_new_n451_), .Y(new_new_n454_));
  NO2        g0432(.A(new_new_n47_), .B(i_4_), .Y(new_new_n455_));
  NA2        g0433(.A(new_new_n455_), .B(new_new_n103_), .Y(new_new_n456_));
  OAI220     g0434(.A0(new_new_n456_), .A1(new_new_n205_), .B0(new_new_n454_), .B1(new_new_n450_), .Y(new_new_n457_));
  NA2        g0435(.A(new_new_n309_), .B(i_0_), .Y(new_new_n458_));
  NO3        g0436(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n459_));
  NA2        g0437(.A(new_new_n265_), .B(new_new_n96_), .Y(new_new_n460_));
  NA2        g0438(.A(new_new_n460_), .B(new_new_n459_), .Y(new_new_n461_));
  NA2        g0439(.A(i_8_), .B(i_9_), .Y(new_new_n462_));
  AOI210     g0440(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n463_));
  OR2        g0441(.A(new_new_n463_), .B(new_new_n462_), .Y(new_new_n464_));
  NA2        g0442(.A(new_new_n283_), .B(new_new_n206_), .Y(new_new_n465_));
  OAI220     g0443(.A0(new_new_n465_), .A1(new_new_n464_), .B0(new_new_n461_), .B1(new_new_n458_), .Y(new_new_n466_));
  NA2        g0444(.A(new_new_n253_), .B(new_new_n308_), .Y(new_new_n467_));
  NO3        g0445(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n468_));
  INV        g0446(.A(new_new_n468_), .Y(new_new_n469_));
  NA3        g0447(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n470_));
  NA4        g0448(.A(new_new_n145_), .B(new_new_n115_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n471_));
  OAI220     g0449(.A0(new_new_n471_), .A1(new_new_n470_), .B0(new_new_n469_), .B1(new_new_n467_), .Y(new_new_n472_));
  NO3        g0450(.A(new_new_n472_), .B(new_new_n466_), .C(new_new_n457_), .Y(new_new_n473_));
  NA2        g0451(.A(new_new_n295_), .B(new_new_n107_), .Y(new_new_n474_));
  OR2        g0452(.A(new_new_n474_), .B(new_new_n208_), .Y(new_new_n475_));
  BUFFER     g0453(.A(new_new_n354_), .Y(new_new_n476_));
  OA220      g0454(.A0(new_new_n476_), .A1(new_new_n162_), .B0(new_new_n475_), .B1(new_new_n233_), .Y(new_new_n477_));
  NA2        g0455(.A(new_new_n95_), .B(i_13_), .Y(new_new_n478_));
  NA2        g0456(.A(new_new_n432_), .B(new_new_n385_), .Y(new_new_n479_));
  NO2        g0457(.A(i_2_), .B(i_13_), .Y(new_new_n480_));
  NO2        g0458(.A(new_new_n479_), .B(new_new_n478_), .Y(new_new_n481_));
  NO3        g0459(.A(i_4_), .B(new_new_n49_), .C(i_8_), .Y(new_new_n482_));
  NO2        g0460(.A(i_6_), .B(i_7_), .Y(new_new_n483_));
  NA2        g0461(.A(new_new_n483_), .B(new_new_n482_), .Y(new_new_n484_));
  NO2        g0462(.A(i_11_), .B(i_1_), .Y(new_new_n485_));
  OR2        g0463(.A(i_11_), .B(i_8_), .Y(new_new_n486_));
  NOi21      g0464(.An(i_2_), .B(i_7_), .Y(new_new_n487_));
  NAi31      g0465(.An(new_new_n486_), .B(new_new_n487_), .C(i_0_), .Y(new_new_n488_));
  NO2        g0466(.A(new_new_n421_), .B(i_6_), .Y(new_new_n489_));
  NA2        g0467(.A(new_new_n489_), .B(new_new_n448_), .Y(new_new_n490_));
  NO2        g0468(.A(new_new_n490_), .B(new_new_n488_), .Y(new_new_n491_));
  NO2        g0469(.A(i_3_), .B(new_new_n193_), .Y(new_new_n492_));
  NO2        g0470(.A(i_6_), .B(i_10_), .Y(new_new_n493_));
  NA4        g0471(.A(new_new_n493_), .B(new_new_n313_), .C(new_new_n492_), .D(new_new_n238_), .Y(new_new_n494_));
  NO2        g0472(.A(new_new_n494_), .B(new_new_n155_), .Y(new_new_n495_));
  NA3        g0473(.A(new_new_n247_), .B(new_new_n171_), .C(new_new_n132_), .Y(new_new_n496_));
  NO2        g0474(.A(new_new_n157_), .B(i_3_), .Y(new_new_n497_));
  NO4        g0475(.A(new_new_n1080_), .B(new_new_n495_), .C(new_new_n491_), .D(new_new_n481_), .Y(new_new_n498_));
  NA2        g0476(.A(new_new_n459_), .B(new_new_n386_), .Y(new_new_n499_));
  NA2        g0477(.A(new_new_n468_), .B(new_new_n393_), .Y(new_new_n500_));
  NO2        g0478(.A(new_new_n500_), .B(new_new_n225_), .Y(new_new_n501_));
  NAi21      g0479(.An(new_new_n218_), .B(new_new_n403_), .Y(new_new_n502_));
  NA2        g0480(.A(new_new_n337_), .B(new_new_n220_), .Y(new_new_n503_));
  NO2        g0481(.A(new_new_n26_), .B(i_5_), .Y(new_new_n504_));
  NA3        g0482(.A(i_6_), .B(new_new_n504_), .C(new_new_n142_), .Y(new_new_n505_));
  OR3        g0483(.A(new_new_n303_), .B(new_new_n38_), .C(new_new_n47_), .Y(new_new_n506_));
  OAI220     g0484(.A0(new_new_n506_), .A1(new_new_n505_), .B0(new_new_n503_), .B1(new_new_n502_), .Y(new_new_n507_));
  NA2        g0485(.A(new_new_n27_), .B(i_10_), .Y(new_new_n508_));
  NO2        g0486(.A(new_new_n508_), .B(new_new_n478_), .Y(new_new_n509_));
  NA4        g0487(.A(new_new_n306_), .B(new_new_n224_), .C(new_new_n73_), .D(new_new_n238_), .Y(new_new_n510_));
  NO2        g0488(.A(new_new_n510_), .B(new_new_n484_), .Y(new_new_n511_));
  NO4        g0489(.A(new_new_n511_), .B(new_new_n509_), .C(new_new_n507_), .D(new_new_n501_), .Y(new_new_n512_));
  NA4        g0490(.A(new_new_n512_), .B(new_new_n498_), .C(new_new_n477_), .D(new_new_n473_), .Y(new_new_n513_));
  NA3        g0491(.A(new_new_n306_), .B(new_new_n175_), .C(new_new_n173_), .Y(new_new_n514_));
  OAI210     g0492(.A0(new_new_n301_), .A1(new_new_n180_), .B0(new_new_n514_), .Y(new_new_n515_));
  AN2        g0493(.A(new_new_n286_), .B(new_new_n235_), .Y(new_new_n516_));
  NA2        g0494(.A(new_new_n516_), .B(new_new_n515_), .Y(new_new_n517_));
  NA2        g0495(.A(new_new_n122_), .B(new_new_n111_), .Y(new_new_n518_));
  AN2        g0496(.A(new_new_n518_), .B(new_new_n459_), .Y(new_new_n519_));
  NA2        g0497(.A(new_new_n313_), .B(new_new_n164_), .Y(new_new_n520_));
  OAI210     g0498(.A0(new_new_n520_), .A1(new_new_n233_), .B0(new_new_n307_), .Y(new_new_n521_));
  AOI220     g0499(.A0(new_new_n521_), .A1(new_new_n324_), .B0(new_new_n519_), .B1(new_new_n309_), .Y(new_new_n522_));
  NA4        g0500(.A(new_new_n449_), .B(new_new_n448_), .C(new_new_n203_), .D(i_2_), .Y(new_new_n523_));
  INV        g0501(.A(new_new_n523_), .Y(new_new_n524_));
  NA2        g0502(.A(new_new_n358_), .B(new_new_n73_), .Y(new_new_n525_));
  NA2        g0503(.A(new_new_n374_), .B(new_new_n366_), .Y(new_new_n526_));
  NO2        g0504(.A(new_new_n36_), .B(i_8_), .Y(new_new_n527_));
  NAi41      g0505(.An(new_new_n525_), .B(new_new_n493_), .C(new_new_n527_), .D(new_new_n47_), .Y(new_new_n528_));
  NA2        g0506(.A(new_new_n39_), .B(i_13_), .Y(new_new_n529_));
  NA2        g0507(.A(new_new_n529_), .B(new_new_n528_), .Y(new_new_n530_));
  AOI210     g0508(.A0(new_new_n524_), .A1(new_new_n204_), .B0(new_new_n530_), .Y(new_new_n531_));
  OAI210     g0509(.A0(i_8_), .A1(new_new_n63_), .B0(new_new_n134_), .Y(new_new_n532_));
  AOI210     g0510(.A0(new_new_n194_), .A1(i_9_), .B0(new_new_n264_), .Y(new_new_n533_));
  NO2        g0511(.A(new_new_n533_), .B(new_new_n199_), .Y(new_new_n534_));
  NO2        g0512(.A(new_new_n182_), .B(new_new_n85_), .Y(new_new_n535_));
  AOI220     g0513(.A0(new_new_n535_), .A1(new_new_n534_), .B0(new_new_n532_), .B1(new_new_n422_), .Y(new_new_n536_));
  NA4        g0514(.A(new_new_n536_), .B(new_new_n531_), .C(new_new_n522_), .D(new_new_n517_), .Y(new_new_n537_));
  NA2        g0515(.A(new_new_n392_), .B(new_new_n295_), .Y(new_new_n538_));
  OAI210     g0516(.A0(new_new_n388_), .A1(new_new_n169_), .B0(new_new_n538_), .Y(new_new_n539_));
  NO2        g0517(.A(i_12_), .B(new_new_n193_), .Y(new_new_n540_));
  NA2        g0518(.A(new_new_n540_), .B(new_new_n226_), .Y(new_new_n541_));
  NO3        g0519(.A(i_10_), .B(new_new_n541_), .C(new_new_n474_), .Y(new_new_n542_));
  NOi31      g0520(.An(new_new_n316_), .B(new_new_n421_), .C(new_new_n38_), .Y(new_new_n543_));
  OAI210     g0521(.A0(new_new_n543_), .A1(new_new_n542_), .B0(new_new_n539_), .Y(new_new_n544_));
  NO2        g0522(.A(i_8_), .B(i_7_), .Y(new_new_n545_));
  OAI210     g0523(.A0(i_0_), .A1(i_12_), .B0(i_5_), .Y(new_new_n546_));
  NA2        g0524(.A(new_new_n546_), .B(new_new_n224_), .Y(new_new_n547_));
  AOI220     g0525(.A0(new_new_n325_), .A1(new_new_n40_), .B0(new_new_n236_), .B1(new_new_n207_), .Y(new_new_n548_));
  OAI220     g0526(.A0(new_new_n548_), .A1(new_new_n182_), .B0(new_new_n547_), .B1(new_new_n244_), .Y(new_new_n549_));
  NA2        g0527(.A(new_new_n45_), .B(i_10_), .Y(new_new_n550_));
  NO2        g0528(.A(new_new_n550_), .B(i_6_), .Y(new_new_n551_));
  NA3        g0529(.A(new_new_n551_), .B(new_new_n549_), .C(new_new_n545_), .Y(new_new_n552_));
  AOI220     g0530(.A0(new_new_n432_), .A1(new_new_n325_), .B0(new_new_n249_), .B1(new_new_n246_), .Y(new_new_n553_));
  OAI220     g0531(.A0(new_new_n553_), .A1(new_new_n261_), .B0(new_new_n478_), .B1(new_new_n133_), .Y(new_new_n554_));
  NA2        g0532(.A(new_new_n554_), .B(new_new_n264_), .Y(new_new_n555_));
  NO2        g0533(.A(new_new_n301_), .B(new_new_n180_), .Y(new_new_n556_));
  NA3        g0534(.A(new_new_n306_), .B(new_new_n173_), .C(new_new_n95_), .Y(new_new_n557_));
  NO2        g0535(.A(new_new_n223_), .B(new_new_n45_), .Y(new_new_n558_));
  NO2        g0536(.A(new_new_n157_), .B(i_5_), .Y(new_new_n559_));
  NA2        g0537(.A(new_new_n559_), .B(new_new_n319_), .Y(new_new_n560_));
  OAI210     g0538(.A0(new_new_n560_), .A1(new_new_n558_), .B0(new_new_n557_), .Y(new_new_n561_));
  OAI210     g0539(.A0(new_new_n561_), .A1(new_new_n556_), .B0(new_new_n468_), .Y(new_new_n562_));
  NA4        g0540(.A(new_new_n562_), .B(new_new_n555_), .C(new_new_n552_), .D(new_new_n544_), .Y(new_new_n563_));
  NA3        g0541(.A(new_new_n220_), .B(new_new_n71_), .C(new_new_n45_), .Y(new_new_n564_));
  NA2        g0542(.A(new_new_n283_), .B(new_new_n84_), .Y(new_new_n565_));
  AOI210     g0543(.A0(new_new_n564_), .A1(new_new_n349_), .B0(new_new_n565_), .Y(new_new_n566_));
  NA2        g0544(.A(new_new_n296_), .B(new_new_n286_), .Y(new_new_n567_));
  NO2        g0545(.A(new_new_n567_), .B(new_new_n172_), .Y(new_new_n568_));
  AOI210     g0546(.A0(new_new_n367_), .A1(new_new_n47_), .B0(new_new_n371_), .Y(new_new_n569_));
  NA2        g0547(.A(i_0_), .B(new_new_n49_), .Y(new_new_n570_));
  NA3        g0548(.A(new_new_n540_), .B(new_new_n274_), .C(new_new_n570_), .Y(new_new_n571_));
  NO2        g0549(.A(new_new_n569_), .B(new_new_n571_), .Y(new_new_n572_));
  NO3        g0550(.A(new_new_n572_), .B(new_new_n568_), .C(new_new_n566_), .Y(new_new_n573_));
  NO4        g0551(.A(new_new_n254_), .B(new_new_n43_), .C(i_2_), .D(new_new_n49_), .Y(new_new_n574_));
  NO3        g0552(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n575_));
  NO2        g0553(.A(new_new_n234_), .B(new_new_n36_), .Y(new_new_n576_));
  AN2        g0554(.A(new_new_n576_), .B(new_new_n575_), .Y(new_new_n577_));
  OA210      g0555(.A0(new_new_n577_), .A1(new_new_n574_), .B0(new_new_n358_), .Y(new_new_n578_));
  NO2        g0556(.A(new_new_n421_), .B(i_1_), .Y(new_new_n579_));
  NOi31      g0557(.An(new_new_n579_), .B(new_new_n460_), .C(new_new_n73_), .Y(new_new_n580_));
  AN4        g0558(.A(new_new_n580_), .B(new_new_n418_), .C(new_new_n504_), .D(i_2_), .Y(new_new_n581_));
  NO2        g0559(.A(new_new_n430_), .B(new_new_n176_), .Y(new_new_n582_));
  NO3        g0560(.A(new_new_n582_), .B(new_new_n581_), .C(new_new_n578_), .Y(new_new_n583_));
  NOi21      g0561(.An(i_10_), .B(i_6_), .Y(new_new_n584_));
  NO2        g0562(.A(new_new_n85_), .B(new_new_n25_), .Y(new_new_n585_));
  AOI220     g0563(.A0(new_new_n283_), .A1(new_new_n585_), .B0(new_new_n274_), .B1(new_new_n584_), .Y(new_new_n586_));
  NO2        g0564(.A(new_new_n586_), .B(new_new_n458_), .Y(new_new_n587_));
  NO2        g0565(.A(new_new_n114_), .B(new_new_n23_), .Y(new_new_n588_));
  NA2        g0566(.A(new_new_n316_), .B(new_new_n164_), .Y(new_new_n589_));
  AOI220     g0567(.A0(new_new_n589_), .A1(new_new_n439_), .B0(new_new_n183_), .B1(new_new_n181_), .Y(new_new_n590_));
  NO2        g0568(.A(new_new_n198_), .B(new_new_n37_), .Y(new_new_n591_));
  NOi31      g0569(.An(new_new_n146_), .B(new_new_n591_), .C(new_new_n332_), .Y(new_new_n592_));
  NO3        g0570(.A(new_new_n592_), .B(new_new_n590_), .C(new_new_n587_), .Y(new_new_n593_));
  NO2        g0571(.A(new_new_n525_), .B(new_new_n381_), .Y(new_new_n594_));
  INV        g0572(.A(new_new_n319_), .Y(new_new_n595_));
  NO2        g0573(.A(i_12_), .B(new_new_n85_), .Y(new_new_n596_));
  NA3        g0574(.A(new_new_n596_), .B(new_new_n274_), .C(new_new_n570_), .Y(new_new_n597_));
  NA3        g0575(.A(new_new_n389_), .B(new_new_n283_), .C(new_new_n220_), .Y(new_new_n598_));
  AOI210     g0576(.A0(new_new_n598_), .A1(new_new_n597_), .B0(new_new_n595_), .Y(new_new_n599_));
  NA2        g0577(.A(new_new_n173_), .B(i_0_), .Y(new_new_n600_));
  NO3        g0578(.A(new_new_n600_), .B(new_new_n343_), .C(new_new_n301_), .Y(new_new_n601_));
  OR2        g0579(.A(i_2_), .B(i_5_), .Y(new_new_n602_));
  OR2        g0580(.A(new_new_n602_), .B(new_new_n413_), .Y(new_new_n603_));
  NO2        g0581(.A(new_new_n603_), .B(new_new_n502_), .Y(new_new_n604_));
  NO4        g0582(.A(new_new_n604_), .B(new_new_n601_), .C(new_new_n599_), .D(new_new_n594_), .Y(new_new_n605_));
  NA4        g0583(.A(new_new_n605_), .B(new_new_n593_), .C(new_new_n583_), .D(new_new_n573_), .Y(new_new_n606_));
  NO4        g0584(.A(new_new_n606_), .B(new_new_n563_), .C(new_new_n537_), .D(new_new_n513_), .Y(new_new_n607_));
  NA4        g0585(.A(new_new_n607_), .B(new_new_n447_), .C(new_new_n357_), .D(new_new_n312_), .Y(men7));
  NO2        g0586(.A(new_new_n92_), .B(new_new_n55_), .Y(new_new_n609_));
  NO2        g0587(.A(new_new_n107_), .B(new_new_n89_), .Y(new_new_n610_));
  NA2        g0588(.A(new_new_n387_), .B(new_new_n610_), .Y(new_new_n611_));
  NA2        g0589(.A(new_new_n493_), .B(new_new_n84_), .Y(new_new_n612_));
  NA2        g0590(.A(i_11_), .B(new_new_n193_), .Y(new_new_n613_));
  NA2        g0591(.A(new_new_n144_), .B(new_new_n613_), .Y(new_new_n614_));
  OAI210     g0592(.A0(new_new_n614_), .A1(new_new_n612_), .B0(new_new_n611_), .Y(new_new_n615_));
  NA3        g0593(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n616_));
  NO2        g0594(.A(new_new_n238_), .B(i_4_), .Y(new_new_n617_));
  NA2        g0595(.A(new_new_n617_), .B(i_8_), .Y(new_new_n618_));
  NO2        g0596(.A(new_new_n104_), .B(new_new_n616_), .Y(new_new_n619_));
  NA2        g0597(.A(i_2_), .B(new_new_n85_), .Y(new_new_n620_));
  OAI210     g0598(.A0(new_new_n88_), .A1(new_new_n203_), .B0(new_new_n204_), .Y(new_new_n621_));
  NO2        g0599(.A(i_7_), .B(new_new_n37_), .Y(new_new_n622_));
  NA2        g0600(.A(i_4_), .B(i_8_), .Y(new_new_n623_));
  AOI210     g0601(.A0(new_new_n623_), .A1(new_new_n306_), .B0(new_new_n622_), .Y(new_new_n624_));
  NO2        g0602(.A(new_new_n624_), .B(new_new_n620_), .Y(new_new_n625_));
  NO4        g0603(.A(new_new_n625_), .B(new_new_n619_), .C(new_new_n615_), .D(new_new_n609_), .Y(new_new_n626_));
  OR2        g0604(.A(i_6_), .B(i_10_), .Y(new_new_n627_));
  NO2        g0605(.A(new_new_n627_), .B(new_new_n23_), .Y(new_new_n628_));
  OR3        g0606(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n629_));
  NO3        g0607(.A(new_new_n629_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n630_));
  INV        g0608(.A(new_new_n200_), .Y(new_new_n631_));
  NO2        g0609(.A(new_new_n630_), .B(new_new_n628_), .Y(new_new_n632_));
  OA220      g0610(.A0(new_new_n632_), .A1(new_new_n595_), .B0(new_new_n1079_), .B1(new_new_n266_), .Y(new_new_n633_));
  AOI210     g0611(.A0(new_new_n633_), .A1(new_new_n626_), .B0(new_new_n63_), .Y(new_new_n634_));
  NOi21      g0612(.An(i_11_), .B(i_7_), .Y(new_new_n635_));
  AO210      g0613(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n636_));
  NO2        g0614(.A(new_new_n636_), .B(new_new_n635_), .Y(new_new_n637_));
  NA2        g0615(.A(new_new_n637_), .B(new_new_n207_), .Y(new_new_n638_));
  NA3        g0616(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n639_));
  NAi31      g0617(.An(new_new_n639_), .B(new_new_n217_), .C(i_11_), .Y(new_new_n640_));
  AOI210     g0618(.A0(new_new_n640_), .A1(new_new_n638_), .B0(new_new_n63_), .Y(new_new_n641_));
  NA2        g0619(.A(new_new_n87_), .B(new_new_n63_), .Y(new_new_n642_));
  AO210      g0620(.A0(new_new_n642_), .A1(new_new_n381_), .B0(new_new_n41_), .Y(new_new_n643_));
  NA2        g0621(.A(new_new_n227_), .B(new_new_n63_), .Y(new_new_n644_));
  NA2        g0622(.A(new_new_n414_), .B(new_new_n31_), .Y(new_new_n645_));
  OR2        g0623(.A(new_new_n209_), .B(new_new_n107_), .Y(new_new_n646_));
  NA2        g0624(.A(new_new_n646_), .B(new_new_n645_), .Y(new_new_n647_));
  NO2        g0625(.A(new_new_n63_), .B(i_9_), .Y(new_new_n648_));
  NO2        g0626(.A(new_new_n648_), .B(i_4_), .Y(new_new_n649_));
  NA2        g0627(.A(new_new_n649_), .B(new_new_n647_), .Y(new_new_n650_));
  NO2        g0628(.A(i_1_), .B(i_12_), .Y(new_new_n651_));
  NA3        g0629(.A(new_new_n651_), .B(new_new_n109_), .C(new_new_n24_), .Y(new_new_n652_));
  NA4        g0630(.A(new_new_n652_), .B(new_new_n650_), .C(new_new_n644_), .D(new_new_n643_), .Y(new_new_n653_));
  OAI210     g0631(.A0(new_new_n653_), .A1(new_new_n641_), .B0(i_6_), .Y(new_new_n654_));
  NO2        g0632(.A(new_new_n238_), .B(new_new_n85_), .Y(new_new_n655_));
  NO2        g0633(.A(new_new_n655_), .B(i_11_), .Y(new_new_n656_));
  INV        g0634(.A(new_new_n461_), .Y(new_new_n657_));
  NO4        g0635(.A(new_new_n217_), .B(new_new_n128_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n658_));
  NA2        g0636(.A(new_new_n658_), .B(new_new_n648_), .Y(new_new_n659_));
  INV        g0637(.A(new_new_n659_), .Y(new_new_n660_));
  NA3        g0638(.A(new_new_n545_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n661_));
  NA2        g0639(.A(new_new_n138_), .B(i_9_), .Y(new_new_n662_));
  NA3        g0640(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n663_));
  NO2        g0641(.A(new_new_n47_), .B(i_1_), .Y(new_new_n664_));
  NO2        g0642(.A(new_new_n662_), .B(new_new_n1077_), .Y(new_new_n665_));
  NA3        g0643(.A(new_new_n648_), .B(new_new_n319_), .C(i_6_), .Y(new_new_n666_));
  NO2        g0644(.A(new_new_n666_), .B(new_new_n23_), .Y(new_new_n667_));
  AOI210     g0645(.A0(new_new_n485_), .A1(new_new_n424_), .B0(new_new_n243_), .Y(new_new_n668_));
  NO2        g0646(.A(new_new_n668_), .B(new_new_n620_), .Y(new_new_n669_));
  NA2        g0647(.A(new_new_n664_), .B(new_new_n265_), .Y(new_new_n670_));
  NO2        g0648(.A(i_11_), .B(new_new_n37_), .Y(new_new_n671_));
  NA2        g0649(.A(new_new_n671_), .B(new_new_n24_), .Y(new_new_n672_));
  NO2        g0650(.A(new_new_n672_), .B(new_new_n670_), .Y(new_new_n673_));
  OR4        g0651(.A(new_new_n673_), .B(new_new_n669_), .C(new_new_n667_), .D(new_new_n665_), .Y(new_new_n674_));
  NO3        g0652(.A(new_new_n674_), .B(new_new_n660_), .C(new_new_n657_), .Y(new_new_n675_));
  NO2        g0653(.A(new_new_n238_), .B(new_new_n100_), .Y(new_new_n676_));
  NO2        g0654(.A(new_new_n676_), .B(new_new_n635_), .Y(new_new_n677_));
  NA2        g0655(.A(new_new_n677_), .B(i_1_), .Y(new_new_n678_));
  NO2        g0656(.A(new_new_n678_), .B(new_new_n629_), .Y(new_new_n679_));
  NO2        g0657(.A(new_new_n420_), .B(new_new_n85_), .Y(new_new_n680_));
  NA2        g0658(.A(new_new_n679_), .B(new_new_n47_), .Y(new_new_n681_));
  NA2        g0659(.A(i_3_), .B(new_new_n193_), .Y(new_new_n682_));
  NO2        g0660(.A(new_new_n234_), .B(new_new_n45_), .Y(new_new_n683_));
  NO3        g0661(.A(new_new_n683_), .B(new_new_n309_), .C(new_new_n239_), .Y(new_new_n684_));
  NO2        g0662(.A(new_new_n117_), .B(new_new_n37_), .Y(new_new_n685_));
  NO2        g0663(.A(new_new_n685_), .B(i_6_), .Y(new_new_n686_));
  NO2        g0664(.A(new_new_n85_), .B(i_9_), .Y(new_new_n687_));
  NO2        g0665(.A(new_new_n687_), .B(new_new_n63_), .Y(new_new_n688_));
  NO2        g0666(.A(new_new_n688_), .B(new_new_n651_), .Y(new_new_n689_));
  NO4        g0667(.A(new_new_n689_), .B(new_new_n686_), .C(new_new_n684_), .D(i_4_), .Y(new_new_n690_));
  NA2        g0668(.A(i_1_), .B(i_3_), .Y(new_new_n691_));
  INV        g0669(.A(new_new_n690_), .Y(new_new_n692_));
  NA4        g0670(.A(new_new_n692_), .B(new_new_n681_), .C(new_new_n675_), .D(new_new_n654_), .Y(new_new_n693_));
  NO3        g0671(.A(new_new_n486_), .B(i_3_), .C(i_7_), .Y(new_new_n694_));
  NOi21      g0672(.An(new_new_n694_), .B(i_10_), .Y(new_new_n695_));
  OA210      g0673(.A0(new_new_n695_), .A1(new_new_n247_), .B0(new_new_n85_), .Y(new_new_n696_));
  NA3        g0674(.A(new_new_n493_), .B(new_new_n527_), .C(new_new_n47_), .Y(new_new_n697_));
  NO3        g0675(.A(new_new_n487_), .B(new_new_n623_), .C(new_new_n85_), .Y(new_new_n698_));
  NA2        g0676(.A(new_new_n698_), .B(new_new_n25_), .Y(new_new_n699_));
  NA3        g0677(.A(new_new_n161_), .B(new_new_n84_), .C(new_new_n85_), .Y(new_new_n700_));
  NA3        g0678(.A(new_new_n700_), .B(new_new_n699_), .C(new_new_n697_), .Y(new_new_n701_));
  OAI210     g0679(.A0(new_new_n701_), .A1(new_new_n696_), .B0(i_1_), .Y(new_new_n702_));
  AOI210     g0680(.A0(new_new_n265_), .A1(new_new_n96_), .B0(i_1_), .Y(new_new_n703_));
  NO2        g0681(.A(new_new_n372_), .B(i_2_), .Y(new_new_n704_));
  NA2        g0682(.A(new_new_n704_), .B(new_new_n703_), .Y(new_new_n705_));
  OAI210     g0683(.A0(new_new_n666_), .A1(new_new_n452_), .B0(new_new_n705_), .Y(new_new_n706_));
  INV        g0684(.A(new_new_n706_), .Y(new_new_n707_));
  AOI210     g0685(.A0(new_new_n707_), .A1(new_new_n702_), .B0(i_13_), .Y(new_new_n708_));
  NA3        g0686(.A(i_11_), .B(new_new_n105_), .C(new_new_n138_), .Y(new_new_n709_));
  AOI220     g0687(.A0(new_new_n480_), .A1(new_new_n161_), .B0(new_new_n455_), .B1(new_new_n138_), .Y(new_new_n710_));
  OAI210     g0688(.A0(new_new_n710_), .A1(new_new_n45_), .B0(new_new_n709_), .Y(new_new_n711_));
  NO2        g0689(.A(new_new_n55_), .B(i_12_), .Y(new_new_n712_));
  INV        g0690(.A(new_new_n712_), .Y(new_new_n713_));
  NO2        g0691(.A(new_new_n487_), .B(new_new_n24_), .Y(new_new_n714_));
  AOI220     g0692(.A0(new_new_n714_), .A1(new_new_n680_), .B0(new_new_n247_), .B1(new_new_n131_), .Y(new_new_n715_));
  OAI220     g0693(.A0(new_new_n715_), .A1(new_new_n41_), .B0(new_new_n713_), .B1(new_new_n92_), .Y(new_new_n716_));
  AOI210     g0694(.A0(new_new_n711_), .A1(new_new_n334_), .B0(new_new_n716_), .Y(new_new_n717_));
  AOI220     g0695(.A0(i_12_), .A1(new_new_n72_), .B0(new_new_n389_), .B1(new_new_n664_), .Y(new_new_n718_));
  NO2        g0696(.A(new_new_n718_), .B(new_new_n244_), .Y(new_new_n719_));
  AOI210     g0697(.A0(new_new_n452_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n720_));
  NOi31      g0698(.An(new_new_n720_), .B(new_new_n612_), .C(new_new_n45_), .Y(new_new_n721_));
  NA2        g0699(.A(new_new_n127_), .B(i_13_), .Y(new_new_n722_));
  NO2        g0700(.A(new_new_n663_), .B(new_new_n114_), .Y(new_new_n723_));
  NO2        g0701(.A(new_new_n722_), .B(new_new_n703_), .Y(new_new_n724_));
  NO3        g0702(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n100_), .Y(new_new_n725_));
  NA2        g0703(.A(new_new_n26_), .B(new_new_n193_), .Y(new_new_n726_));
  INV        g0704(.A(new_new_n725_), .Y(new_new_n727_));
  NO2        g0705(.A(new_new_n727_), .B(new_new_n631_), .Y(new_new_n728_));
  NO4        g0706(.A(new_new_n728_), .B(new_new_n724_), .C(new_new_n721_), .D(new_new_n719_), .Y(new_new_n729_));
  OR2        g0707(.A(i_11_), .B(i_6_), .Y(new_new_n730_));
  NA3        g0708(.A(new_new_n617_), .B(new_new_n726_), .C(i_7_), .Y(new_new_n731_));
  NO2        g0709(.A(new_new_n731_), .B(new_new_n730_), .Y(new_new_n732_));
  NA3        g0710(.A(new_new_n414_), .B(new_new_n622_), .C(new_new_n96_), .Y(new_new_n733_));
  NA2        g0711(.A(new_new_n656_), .B(i_13_), .Y(new_new_n734_));
  NA2        g0712(.A(new_new_n101_), .B(new_new_n726_), .Y(new_new_n735_));
  NAi21      g0713(.An(i_11_), .B(i_12_), .Y(new_new_n736_));
  NOi41      g0714(.An(new_new_n110_), .B(new_new_n736_), .C(i_13_), .D(new_new_n85_), .Y(new_new_n737_));
  NO3        g0715(.A(new_new_n487_), .B(new_new_n596_), .C(new_new_n623_), .Y(new_new_n738_));
  AOI220     g0716(.A0(new_new_n738_), .A1(new_new_n313_), .B0(new_new_n737_), .B1(new_new_n735_), .Y(new_new_n739_));
  NA3        g0717(.A(new_new_n739_), .B(new_new_n734_), .C(new_new_n733_), .Y(new_new_n740_));
  OAI210     g0718(.A0(new_new_n740_), .A1(new_new_n732_), .B0(new_new_n63_), .Y(new_new_n741_));
  NO2        g0719(.A(i_2_), .B(i_12_), .Y(new_new_n742_));
  NA2        g0720(.A(new_new_n371_), .B(new_new_n742_), .Y(new_new_n743_));
  NA2        g0721(.A(i_8_), .B(new_new_n25_), .Y(new_new_n744_));
  NO3        g0722(.A(new_new_n744_), .B(new_new_n387_), .C(new_new_n617_), .Y(new_new_n745_));
  OAI210     g0723(.A0(new_new_n745_), .A1(new_new_n373_), .B0(new_new_n371_), .Y(new_new_n746_));
  NO2        g0724(.A(new_new_n128_), .B(i_2_), .Y(new_new_n747_));
  NA2        g0725(.A(new_new_n746_), .B(new_new_n743_), .Y(new_new_n748_));
  NA3        g0726(.A(new_new_n748_), .B(new_new_n46_), .C(new_new_n226_), .Y(new_new_n749_));
  NA4        g0727(.A(new_new_n749_), .B(new_new_n741_), .C(new_new_n729_), .D(new_new_n717_), .Y(new_new_n750_));
  OR4        g0728(.A(new_new_n750_), .B(new_new_n708_), .C(new_new_n693_), .D(new_new_n634_), .Y(men5));
  AOI210     g0729(.A0(new_new_n677_), .A1(new_new_n268_), .B0(new_new_n422_), .Y(new_new_n752_));
  AN2        g0730(.A(new_new_n24_), .B(i_10_), .Y(new_new_n753_));
  NA3        g0731(.A(new_new_n753_), .B(new_new_n742_), .C(new_new_n107_), .Y(new_new_n754_));
  NO2        g0732(.A(new_new_n618_), .B(i_11_), .Y(new_new_n755_));
  NA2        g0733(.A(new_new_n88_), .B(new_new_n755_), .Y(new_new_n756_));
  NA3        g0734(.A(new_new_n756_), .B(new_new_n754_), .C(new_new_n752_), .Y(new_new_n757_));
  NO3        g0735(.A(i_11_), .B(new_new_n238_), .C(i_13_), .Y(new_new_n758_));
  NO2        g0736(.A(new_new_n124_), .B(new_new_n23_), .Y(new_new_n759_));
  NA2        g0737(.A(i_12_), .B(i_8_), .Y(new_new_n760_));
  OAI210     g0738(.A0(new_new_n47_), .A1(i_3_), .B0(new_new_n760_), .Y(new_new_n761_));
  INV        g0739(.A(new_new_n451_), .Y(new_new_n762_));
  AOI220     g0740(.A0(new_new_n319_), .A1(new_new_n588_), .B0(new_new_n761_), .B1(new_new_n759_), .Y(new_new_n763_));
  INV        g0741(.A(new_new_n763_), .Y(new_new_n764_));
  NO2        g0742(.A(new_new_n764_), .B(new_new_n757_), .Y(new_new_n765_));
  INV        g0743(.A(new_new_n171_), .Y(new_new_n766_));
  INV        g0744(.A(new_new_n247_), .Y(new_new_n767_));
  OAI210     g0745(.A0(new_new_n704_), .A1(new_new_n453_), .B0(new_new_n110_), .Y(new_new_n768_));
  AOI210     g0746(.A0(new_new_n768_), .A1(new_new_n767_), .B0(new_new_n766_), .Y(new_new_n769_));
  NO2        g0747(.A(new_new_n462_), .B(new_new_n26_), .Y(new_new_n770_));
  NO2        g0748(.A(new_new_n770_), .B(new_new_n424_), .Y(new_new_n771_));
  NA2        g0749(.A(new_new_n771_), .B(i_2_), .Y(new_new_n772_));
  INV        g0750(.A(new_new_n772_), .Y(new_new_n773_));
  AOI210     g0751(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n421_), .Y(new_new_n774_));
  AOI210     g0752(.A0(new_new_n774_), .A1(new_new_n773_), .B0(new_new_n769_), .Y(new_new_n775_));
  NO2        g0753(.A(new_new_n190_), .B(new_new_n125_), .Y(new_new_n776_));
  OAI210     g0754(.A0(new_new_n776_), .A1(new_new_n759_), .B0(i_2_), .Y(new_new_n777_));
  NO2        g0755(.A(new_new_n777_), .B(new_new_n193_), .Y(new_new_n778_));
  OA210      g0756(.A0(new_new_n637_), .A1(new_new_n126_), .B0(i_13_), .Y(new_new_n779_));
  NA2        g0757(.A(new_new_n200_), .B(new_new_n203_), .Y(new_new_n780_));
  NA2        g0758(.A(new_new_n151_), .B(new_new_n613_), .Y(new_new_n781_));
  AOI210     g0759(.A0(new_new_n781_), .A1(new_new_n780_), .B0(new_new_n376_), .Y(new_new_n782_));
  AOI210     g0760(.A0(new_new_n209_), .A1(new_new_n148_), .B0(new_new_n527_), .Y(new_new_n783_));
  NA2        g0761(.A(new_new_n783_), .B(new_new_n424_), .Y(new_new_n784_));
  NO2        g0762(.A(new_new_n101_), .B(new_new_n45_), .Y(new_new_n785_));
  INV        g0763(.A(new_new_n302_), .Y(new_new_n786_));
  NA4        g0764(.A(new_new_n786_), .B(new_new_n306_), .C(new_new_n124_), .D(new_new_n43_), .Y(new_new_n787_));
  OAI210     g0765(.A0(new_new_n787_), .A1(new_new_n785_), .B0(new_new_n784_), .Y(new_new_n788_));
  NO4        g0766(.A(new_new_n788_), .B(new_new_n782_), .C(new_new_n779_), .D(new_new_n778_), .Y(new_new_n789_));
  NA2        g0767(.A(new_new_n588_), .B(new_new_n28_), .Y(new_new_n790_));
  NA2        g0768(.A(new_new_n758_), .B(new_new_n275_), .Y(new_new_n791_));
  NA2        g0769(.A(new_new_n791_), .B(new_new_n790_), .Y(new_new_n792_));
  NO2        g0770(.A(new_new_n62_), .B(i_12_), .Y(new_new_n793_));
  NO2        g0771(.A(new_new_n793_), .B(new_new_n126_), .Y(new_new_n794_));
  NO2        g0772(.A(new_new_n794_), .B(new_new_n613_), .Y(new_new_n795_));
  AOI220     g0773(.A0(new_new_n795_), .A1(new_new_n36_), .B0(new_new_n792_), .B1(new_new_n47_), .Y(new_new_n796_));
  NA4        g0774(.A(new_new_n796_), .B(new_new_n789_), .C(new_new_n775_), .D(new_new_n765_), .Y(men6));
  NO3        g0775(.A(new_new_n256_), .B(new_new_n308_), .C(i_1_), .Y(new_new_n798_));
  NO2        g0776(.A(new_new_n185_), .B(new_new_n139_), .Y(new_new_n799_));
  OAI210     g0777(.A0(new_new_n799_), .A1(new_new_n798_), .B0(new_new_n747_), .Y(new_new_n800_));
  NA4        g0778(.A(new_new_n393_), .B(new_new_n492_), .C(new_new_n71_), .D(new_new_n100_), .Y(new_new_n801_));
  INV        g0779(.A(new_new_n801_), .Y(new_new_n802_));
  NO2        g0780(.A(i_11_), .B(i_9_), .Y(new_new_n803_));
  NO2        g0781(.A(new_new_n802_), .B(new_new_n330_), .Y(new_new_n804_));
  AO210      g0782(.A0(new_new_n804_), .A1(new_new_n800_), .B0(i_12_), .Y(new_new_n805_));
  NA2        g0783(.A(new_new_n377_), .B(new_new_n337_), .Y(new_new_n806_));
  NA2        g0784(.A(new_new_n596_), .B(new_new_n63_), .Y(new_new_n807_));
  NA2        g0785(.A(new_new_n695_), .B(new_new_n71_), .Y(new_new_n808_));
  NA4        g0786(.A(new_new_n642_), .B(new_new_n808_), .C(new_new_n807_), .D(new_new_n806_), .Y(new_new_n809_));
  INV        g0787(.A(new_new_n197_), .Y(new_new_n810_));
  AOI220     g0788(.A0(new_new_n810_), .A1(new_new_n803_), .B0(new_new_n809_), .B1(new_new_n73_), .Y(new_new_n811_));
  INV        g0789(.A(new_new_n329_), .Y(new_new_n812_));
  NA2        g0790(.A(new_new_n75_), .B(new_new_n131_), .Y(new_new_n813_));
  NO2        g0791(.A(new_new_n813_), .B(new_new_n812_), .Y(new_new_n814_));
  NO2        g0792(.A(new_new_n254_), .B(i_9_), .Y(new_new_n815_));
  NA2        g0793(.A(new_new_n815_), .B(new_new_n793_), .Y(new_new_n816_));
  AOI210     g0794(.A0(new_new_n816_), .A1(new_new_n526_), .B0(new_new_n185_), .Y(new_new_n817_));
  NO2        g0795(.A(new_new_n32_), .B(i_11_), .Y(new_new_n818_));
  NA3        g0796(.A(new_new_n818_), .B(new_new_n483_), .C(new_new_n393_), .Y(new_new_n819_));
  NAi32      g0797(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n820_));
  AOI210     g0798(.A0(new_new_n730_), .A1(new_new_n86_), .B0(new_new_n820_), .Y(new_new_n821_));
  OAI210     g0799(.A0(new_new_n694_), .A1(new_new_n576_), .B0(new_new_n575_), .Y(new_new_n822_));
  NAi31      g0800(.An(new_new_n821_), .B(new_new_n822_), .C(new_new_n819_), .Y(new_new_n823_));
  OR3        g0801(.A(new_new_n823_), .B(new_new_n817_), .C(new_new_n814_), .Y(new_new_n824_));
  NO2        g0802(.A(i_11_), .B(i_2_), .Y(new_new_n825_));
  NA2        g0803(.A(new_new_n49_), .B(new_new_n37_), .Y(new_new_n826_));
  NO2        g0804(.A(new_new_n826_), .B(new_new_n413_), .Y(new_new_n827_));
  NA2        g0805(.A(new_new_n827_), .B(new_new_n825_), .Y(new_new_n828_));
  AO220      g0806(.A0(new_new_n362_), .A1(new_new_n353_), .B0(new_new_n401_), .B1(new_new_n613_), .Y(new_new_n829_));
  NA3        g0807(.A(new_new_n829_), .B(new_new_n257_), .C(i_7_), .Y(new_new_n830_));
  BUFFER     g0808(.A(new_new_n637_), .Y(new_new_n831_));
  NA3        g0809(.A(new_new_n831_), .B(new_new_n147_), .C(new_new_n69_), .Y(new_new_n832_));
  AO210      g0810(.A0(new_new_n500_), .A1(new_new_n762_), .B0(new_new_n36_), .Y(new_new_n833_));
  NA4        g0811(.A(new_new_n833_), .B(new_new_n832_), .C(new_new_n830_), .D(new_new_n828_), .Y(new_new_n834_));
  OAI210     g0812(.A0(new_new_n655_), .A1(i_11_), .B0(new_new_n86_), .Y(new_new_n835_));
  NA2        g0813(.A(new_new_n835_), .B(new_new_n575_), .Y(new_new_n836_));
  NA2        g0814(.A(new_new_n401_), .B(new_new_n70_), .Y(new_new_n837_));
  NA3        g0815(.A(new_new_n837_), .B(new_new_n836_), .C(new_new_n621_), .Y(new_new_n838_));
  AO210      g0816(.A0(new_new_n527_), .A1(new_new_n47_), .B0(new_new_n87_), .Y(new_new_n839_));
  NA3        g0817(.A(new_new_n839_), .B(new_new_n493_), .C(new_new_n220_), .Y(new_new_n840_));
  AOI210     g0818(.A0(new_new_n453_), .A1(new_new_n451_), .B0(new_new_n574_), .Y(new_new_n841_));
  NA2        g0819(.A(new_new_n111_), .B(new_new_n412_), .Y(new_new_n842_));
  NA2        g0820(.A(new_new_n246_), .B(new_new_n47_), .Y(new_new_n843_));
  INV        g0821(.A(new_new_n603_), .Y(new_new_n844_));
  NA3        g0822(.A(new_new_n844_), .B(new_new_n329_), .C(i_7_), .Y(new_new_n845_));
  NA4        g0823(.A(new_new_n845_), .B(new_new_n842_), .C(new_new_n841_), .D(new_new_n840_), .Y(new_new_n846_));
  NO4        g0824(.A(new_new_n846_), .B(new_new_n838_), .C(new_new_n834_), .D(new_new_n824_), .Y(new_new_n847_));
  NA4        g0825(.A(new_new_n847_), .B(new_new_n811_), .C(new_new_n805_), .D(new_new_n383_), .Y(men3));
  NA2        g0826(.A(i_12_), .B(i_10_), .Y(new_new_n849_));
  NA2        g0827(.A(i_6_), .B(i_7_), .Y(new_new_n850_));
  NO2        g0828(.A(new_new_n850_), .B(i_0_), .Y(new_new_n851_));
  NO2        g0829(.A(i_11_), .B(new_new_n238_), .Y(new_new_n852_));
  OAI210     g0830(.A0(new_new_n851_), .A1(new_new_n290_), .B0(new_new_n852_), .Y(new_new_n853_));
  NO2        g0831(.A(new_new_n853_), .B(new_new_n193_), .Y(new_new_n854_));
  NO3        g0832(.A(new_new_n458_), .B(new_new_n89_), .C(new_new_n45_), .Y(new_new_n855_));
  OA210      g0833(.A0(new_new_n855_), .A1(new_new_n854_), .B0(new_new_n173_), .Y(new_new_n856_));
  NA2        g0834(.A(new_new_n621_), .B(new_new_n375_), .Y(new_new_n857_));
  NA2        g0835(.A(new_new_n857_), .B(new_new_n40_), .Y(new_new_n858_));
  NOi21      g0836(.An(new_new_n95_), .B(new_new_n771_), .Y(new_new_n859_));
  NA2        g0837(.A(new_new_n414_), .B(new_new_n46_), .Y(new_new_n860_));
  INV        g0838(.A(new_new_n859_), .Y(new_new_n861_));
  AOI210     g0839(.A0(new_new_n861_), .A1(new_new_n858_), .B0(new_new_n49_), .Y(new_new_n862_));
  NO4        g0840(.A(new_new_n380_), .B(new_new_n386_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n863_));
  NA2        g0841(.A(new_new_n185_), .B(new_new_n584_), .Y(new_new_n864_));
  NOi21      g0842(.An(new_new_n864_), .B(new_new_n863_), .Y(new_new_n865_));
  NA2        g0843(.A(new_new_n720_), .B(new_new_n687_), .Y(new_new_n866_));
  NA2        g0844(.A(new_new_n335_), .B(new_new_n441_), .Y(new_new_n867_));
  OAI220     g0845(.A0(new_new_n867_), .A1(new_new_n866_), .B0(new_new_n865_), .B1(new_new_n63_), .Y(new_new_n868_));
  NOi21      g0846(.An(i_5_), .B(i_9_), .Y(new_new_n869_));
  NA2        g0847(.A(new_new_n869_), .B(new_new_n449_), .Y(new_new_n870_));
  AOI210     g0848(.A0(new_new_n265_), .A1(new_new_n485_), .B0(new_new_n698_), .Y(new_new_n871_));
  NO3        g0849(.A(new_new_n417_), .B(new_new_n265_), .C(new_new_n73_), .Y(new_new_n872_));
  NO2        g0850(.A(new_new_n174_), .B(new_new_n148_), .Y(new_new_n873_));
  AOI210     g0851(.A0(new_new_n873_), .A1(new_new_n246_), .B0(new_new_n872_), .Y(new_new_n874_));
  OAI220     g0852(.A0(new_new_n874_), .A1(new_new_n180_), .B0(new_new_n871_), .B1(new_new_n870_), .Y(new_new_n875_));
  NO4        g0853(.A(new_new_n875_), .B(new_new_n868_), .C(new_new_n862_), .D(new_new_n856_), .Y(new_new_n876_));
  NA2        g0854(.A(new_new_n185_), .B(new_new_n24_), .Y(new_new_n877_));
  NO2        g0855(.A(new_new_n685_), .B(new_new_n610_), .Y(new_new_n878_));
  NO2        g0856(.A(new_new_n878_), .B(new_new_n877_), .Y(new_new_n879_));
  NA2        g0857(.A(new_new_n313_), .B(new_new_n129_), .Y(new_new_n880_));
  NAi21      g0858(.An(new_new_n162_), .B(new_new_n441_), .Y(new_new_n881_));
  OAI220     g0859(.A0(new_new_n881_), .A1(new_new_n843_), .B0(new_new_n880_), .B1(new_new_n404_), .Y(new_new_n882_));
  NO2        g0860(.A(new_new_n882_), .B(new_new_n879_), .Y(new_new_n883_));
  NO2        g0861(.A(new_new_n393_), .B(new_new_n294_), .Y(new_new_n884_));
  NA2        g0862(.A(new_new_n884_), .B(new_new_n723_), .Y(new_new_n885_));
  NA2        g0863(.A(new_new_n585_), .B(i_0_), .Y(new_new_n886_));
  NO3        g0864(.A(new_new_n886_), .B(new_new_n388_), .C(new_new_n88_), .Y(new_new_n887_));
  NO4        g0865(.A(new_new_n602_), .B(new_new_n217_), .C(new_new_n421_), .D(new_new_n413_), .Y(new_new_n888_));
  AOI210     g0866(.A0(new_new_n888_), .A1(i_11_), .B0(new_new_n887_), .Y(new_new_n889_));
  INV        g0867(.A(new_new_n483_), .Y(new_new_n890_));
  AN2        g0868(.A(new_new_n95_), .B(new_new_n245_), .Y(new_new_n891_));
  NA2        g0869(.A(new_new_n758_), .B(new_new_n330_), .Y(new_new_n892_));
  INV        g0870(.A(new_new_n58_), .Y(new_new_n893_));
  OAI220     g0871(.A0(new_new_n893_), .A1(new_new_n892_), .B0(new_new_n672_), .B1(new_new_n547_), .Y(new_new_n894_));
  NA2        g0872(.A(i_0_), .B(i_10_), .Y(new_new_n895_));
  OAI210     g0873(.A0(new_new_n895_), .A1(new_new_n85_), .B0(new_new_n550_), .Y(new_new_n896_));
  NO4        g0874(.A(new_new_n114_), .B(new_new_n58_), .C(new_new_n682_), .D(i_5_), .Y(new_new_n897_));
  AN2        g0875(.A(new_new_n897_), .B(new_new_n896_), .Y(new_new_n898_));
  AOI220     g0876(.A0(new_new_n335_), .A1(new_new_n97_), .B0(new_new_n185_), .B1(new_new_n84_), .Y(new_new_n899_));
  NA2        g0877(.A(new_new_n579_), .B(i_4_), .Y(new_new_n900_));
  NA2        g0878(.A(new_new_n188_), .B(new_new_n203_), .Y(new_new_n901_));
  OAI220     g0879(.A0(new_new_n901_), .A1(new_new_n892_), .B0(new_new_n900_), .B1(new_new_n899_), .Y(new_new_n902_));
  NO4        g0880(.A(new_new_n902_), .B(new_new_n898_), .C(new_new_n894_), .D(new_new_n891_), .Y(new_new_n903_));
  NA4        g0881(.A(new_new_n903_), .B(new_new_n889_), .C(new_new_n885_), .D(new_new_n883_), .Y(new_new_n904_));
  NO2        g0882(.A(new_new_n102_), .B(new_new_n37_), .Y(new_new_n905_));
  NA2        g0883(.A(i_11_), .B(i_9_), .Y(new_new_n906_));
  NO3        g0884(.A(i_12_), .B(new_new_n906_), .C(new_new_n620_), .Y(new_new_n907_));
  AO220      g0885(.A0(new_new_n907_), .A1(new_new_n905_), .B0(new_new_n267_), .B1(new_new_n87_), .Y(new_new_n908_));
  NO2        g0886(.A(new_new_n49_), .B(i_7_), .Y(new_new_n909_));
  NA2        g0887(.A(new_new_n398_), .B(new_new_n178_), .Y(new_new_n910_));
  NA2        g0888(.A(new_new_n910_), .B(new_new_n160_), .Y(new_new_n911_));
  NO2        g0889(.A(new_new_n906_), .B(new_new_n73_), .Y(new_new_n912_));
  NO2        g0890(.A(new_new_n174_), .B(i_0_), .Y(new_new_n913_));
  INV        g0891(.A(new_new_n913_), .Y(new_new_n914_));
  NA2        g0892(.A(new_new_n483_), .B(new_new_n232_), .Y(new_new_n915_));
  AOI210     g0893(.A0(new_new_n374_), .A1(new_new_n42_), .B0(new_new_n411_), .Y(new_new_n916_));
  OAI220     g0894(.A0(new_new_n916_), .A1(new_new_n870_), .B0(new_new_n915_), .B1(new_new_n914_), .Y(new_new_n917_));
  NO3        g0895(.A(new_new_n917_), .B(new_new_n911_), .C(new_new_n908_), .Y(new_new_n918_));
  NA2        g0896(.A(new_new_n671_), .B(new_new_n121_), .Y(new_new_n919_));
  NO2        g0897(.A(i_6_), .B(new_new_n919_), .Y(new_new_n920_));
  AOI210     g0898(.A0(new_new_n452_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n921_));
  NA2        g0899(.A(new_new_n171_), .B(new_new_n102_), .Y(new_new_n922_));
  NOi32      g0900(.An(new_new_n921_), .Bn(new_new_n188_), .C(new_new_n922_), .Y(new_new_n923_));
  NA2        g0901(.A(new_new_n622_), .B(new_new_n330_), .Y(new_new_n924_));
  NO2        g0902(.A(new_new_n924_), .B(new_new_n860_), .Y(new_new_n925_));
  NO3        g0903(.A(new_new_n925_), .B(new_new_n923_), .C(new_new_n920_), .Y(new_new_n926_));
  NOi21      g0904(.An(i_7_), .B(i_5_), .Y(new_new_n927_));
  NOi31      g0905(.An(new_new_n927_), .B(i_0_), .C(new_new_n736_), .Y(new_new_n928_));
  NA3        g0906(.A(new_new_n928_), .B(new_new_n387_), .C(i_6_), .Y(new_new_n929_));
  OA210      g0907(.A0(new_new_n922_), .A1(new_new_n526_), .B0(new_new_n929_), .Y(new_new_n930_));
  NO3        g0908(.A(new_new_n407_), .B(new_new_n363_), .C(new_new_n361_), .Y(new_new_n931_));
  NO2        g0909(.A(new_new_n259_), .B(new_new_n320_), .Y(new_new_n932_));
  NO2        g0910(.A(new_new_n736_), .B(new_new_n258_), .Y(new_new_n933_));
  AOI210     g0911(.A0(new_new_n933_), .A1(new_new_n932_), .B0(new_new_n931_), .Y(new_new_n934_));
  NA4        g0912(.A(new_new_n934_), .B(new_new_n930_), .C(new_new_n926_), .D(new_new_n918_), .Y(new_new_n935_));
  NO2        g0913(.A(new_new_n877_), .B(new_new_n241_), .Y(new_new_n936_));
  AN2        g0914(.A(new_new_n334_), .B(new_new_n330_), .Y(new_new_n937_));
  AN2        g0915(.A(new_new_n937_), .B(new_new_n873_), .Y(new_new_n938_));
  OAI210     g0916(.A0(new_new_n938_), .A1(new_new_n936_), .B0(i_10_), .Y(new_new_n939_));
  NO2        g0917(.A(new_new_n849_), .B(new_new_n319_), .Y(new_new_n940_));
  NA2        g0918(.A(new_new_n940_), .B(new_new_n912_), .Y(new_new_n941_));
  NA3        g0919(.A(new_new_n482_), .B(new_new_n414_), .C(new_new_n46_), .Y(new_new_n942_));
  OAI210     g0920(.A0(new_new_n881_), .A1(new_new_n890_), .B0(new_new_n942_), .Y(new_new_n943_));
  NO2        g0921(.A(new_new_n257_), .B(new_new_n47_), .Y(new_new_n944_));
  NA2        g0922(.A(new_new_n912_), .B(new_new_n306_), .Y(new_new_n945_));
  OAI210     g0923(.A0(new_new_n944_), .A1(new_new_n187_), .B0(new_new_n945_), .Y(new_new_n946_));
  AOI220     g0924(.A0(new_new_n946_), .A1(new_new_n483_), .B0(new_new_n943_), .B1(new_new_n73_), .Y(new_new_n947_));
  NA3        g0925(.A(new_new_n826_), .B(new_new_n385_), .C(new_new_n655_), .Y(new_new_n948_));
  NA2        g0926(.A(new_new_n92_), .B(new_new_n45_), .Y(new_new_n949_));
  NO2        g0927(.A(new_new_n75_), .B(new_new_n760_), .Y(new_new_n950_));
  AOI220     g0928(.A0(new_new_n950_), .A1(new_new_n949_), .B0(new_new_n173_), .B1(new_new_n610_), .Y(new_new_n951_));
  AOI210     g0929(.A0(new_new_n951_), .A1(new_new_n948_), .B0(new_new_n48_), .Y(new_new_n952_));
  NO3        g0930(.A(new_new_n602_), .B(new_new_n360_), .C(new_new_n24_), .Y(new_new_n953_));
  AOI210     g0931(.A0(new_new_n714_), .A1(new_new_n559_), .B0(new_new_n953_), .Y(new_new_n954_));
  NAi21      g0932(.An(i_9_), .B(i_5_), .Y(new_new_n955_));
  NO2        g0933(.A(new_new_n955_), .B(new_new_n407_), .Y(new_new_n956_));
  NO2        g0934(.A(new_new_n616_), .B(new_new_n104_), .Y(new_new_n957_));
  AOI220     g0935(.A0(new_new_n957_), .A1(i_0_), .B0(new_new_n956_), .B1(new_new_n637_), .Y(new_new_n958_));
  OAI220     g0936(.A0(new_new_n958_), .A1(new_new_n85_), .B0(new_new_n954_), .B1(new_new_n172_), .Y(new_new_n959_));
  NO3        g0937(.A(new_new_n959_), .B(new_new_n952_), .C(new_new_n530_), .Y(new_new_n960_));
  NA4        g0938(.A(new_new_n960_), .B(new_new_n947_), .C(new_new_n941_), .D(new_new_n939_), .Y(new_new_n961_));
  NO3        g0939(.A(new_new_n961_), .B(new_new_n935_), .C(new_new_n904_), .Y(new_new_n962_));
  NO2        g0940(.A(i_0_), .B(new_new_n736_), .Y(new_new_n963_));
  NA2        g0941(.A(new_new_n73_), .B(new_new_n45_), .Y(new_new_n964_));
  NO3        g0942(.A(new_new_n104_), .B(i_5_), .C(new_new_n25_), .Y(new_new_n965_));
  AO220      g0943(.A0(new_new_n965_), .A1(new_new_n45_), .B0(new_new_n963_), .B1(new_new_n173_), .Y(new_new_n966_));
  NO2        g0944(.A(new_new_n807_), .B(new_new_n922_), .Y(new_new_n967_));
  AOI210     g0945(.A0(new_new_n966_), .A1(new_new_n350_), .B0(new_new_n967_), .Y(new_new_n968_));
  NA2        g0946(.A(new_new_n747_), .B(new_new_n146_), .Y(new_new_n969_));
  INV        g0947(.A(new_new_n969_), .Y(new_new_n970_));
  NA3        g0948(.A(new_new_n970_), .B(new_new_n687_), .C(new_new_n73_), .Y(new_new_n971_));
  NO2        g0949(.A(new_new_n822_), .B(new_new_n407_), .Y(new_new_n972_));
  NA3        g0950(.A(new_new_n851_), .B(i_2_), .C(new_new_n49_), .Y(new_new_n973_));
  NA2        g0951(.A(new_new_n852_), .B(i_9_), .Y(new_new_n974_));
  AOI210     g0952(.A0(new_new_n973_), .A1(new_new_n505_), .B0(new_new_n974_), .Y(new_new_n975_));
  OAI210     g0953(.A0(new_new_n246_), .A1(i_9_), .B0(new_new_n231_), .Y(new_new_n976_));
  AOI210     g0954(.A0(new_new_n976_), .A1(new_new_n886_), .B0(new_new_n153_), .Y(new_new_n977_));
  NO3        g0955(.A(new_new_n977_), .B(new_new_n975_), .C(new_new_n972_), .Y(new_new_n978_));
  NA3        g0956(.A(new_new_n978_), .B(new_new_n971_), .C(new_new_n968_), .Y(new_new_n979_));
  NA2        g0957(.A(new_new_n937_), .B(new_new_n376_), .Y(new_new_n980_));
  AOI210     g0958(.A0(new_new_n301_), .A1(new_new_n162_), .B0(new_new_n980_), .Y(new_new_n981_));
  NA3        g0959(.A(new_new_n40_), .B(new_new_n28_), .C(new_new_n45_), .Y(new_new_n982_));
  NA2        g0960(.A(new_new_n909_), .B(new_new_n497_), .Y(new_new_n983_));
  AOI210     g0961(.A0(new_new_n982_), .A1(new_new_n162_), .B0(new_new_n983_), .Y(new_new_n984_));
  NO2        g0962(.A(new_new_n984_), .B(new_new_n981_), .Y(new_new_n985_));
  NA2        g0963(.A(new_new_n580_), .B(new_new_n75_), .Y(new_new_n986_));
  NO3        g0964(.A(new_new_n211_), .B(new_new_n386_), .C(i_0_), .Y(new_new_n987_));
  OAI210     g0965(.A0(new_new_n987_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n988_));
  INV        g0966(.A(new_new_n220_), .Y(new_new_n989_));
  OAI220     g0967(.A0(new_new_n541_), .A1(new_new_n139_), .B0(i_12_), .B1(new_new_n631_), .Y(new_new_n990_));
  NA3        g0968(.A(new_new_n990_), .B(new_new_n402_), .C(new_new_n989_), .Y(new_new_n991_));
  NA4        g0969(.A(new_new_n991_), .B(new_new_n988_), .C(new_new_n986_), .D(new_new_n985_), .Y(new_new_n992_));
  NO2        g0970(.A(new_new_n244_), .B(new_new_n92_), .Y(new_new_n993_));
  AOI210     g0971(.A0(new_new_n993_), .A1(new_new_n963_), .B0(new_new_n108_), .Y(new_new_n994_));
  AOI220     g0972(.A0(new_new_n927_), .A1(new_new_n497_), .B0(new_new_n851_), .B1(new_new_n163_), .Y(new_new_n995_));
  NA2        g0973(.A(new_new_n353_), .B(new_new_n175_), .Y(new_new_n996_));
  OA220      g0974(.A0(new_new_n996_), .A1(new_new_n995_), .B0(new_new_n994_), .B1(i_5_), .Y(new_new_n997_));
  AOI210     g0975(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n174_), .Y(new_new_n998_));
  NA3        g0976(.A(new_new_n628_), .B(new_new_n185_), .C(new_new_n84_), .Y(new_new_n999_));
  NA2        g0977(.A(new_new_n999_), .B(new_new_n557_), .Y(new_new_n1000_));
  NO3        g0978(.A(new_new_n860_), .B(new_new_n55_), .C(new_new_n49_), .Y(new_new_n1001_));
  NA2        g0979(.A(new_new_n499_), .B(new_new_n496_), .Y(new_new_n1002_));
  NO3        g0980(.A(new_new_n1002_), .B(new_new_n1001_), .C(new_new_n1000_), .Y(new_new_n1003_));
  NA3        g0981(.A(new_new_n393_), .B(new_new_n171_), .C(new_new_n170_), .Y(new_new_n1004_));
  NA3        g0982(.A(new_new_n909_), .B(new_new_n290_), .C(new_new_n231_), .Y(new_new_n1005_));
  NA2        g0983(.A(new_new_n1005_), .B(new_new_n1004_), .Y(new_new_n1006_));
  NA3        g0984(.A(new_new_n393_), .B(new_new_n336_), .C(new_new_n223_), .Y(new_new_n1007_));
  INV        g0985(.A(new_new_n1007_), .Y(new_new_n1008_));
  NOi31      g0986(.An(new_new_n392_), .B(new_new_n964_), .C(new_new_n241_), .Y(new_new_n1009_));
  NO3        g0987(.A(new_new_n906_), .B(new_new_n220_), .C(new_new_n190_), .Y(new_new_n1010_));
  NO4        g0988(.A(new_new_n1010_), .B(new_new_n1009_), .C(new_new_n1008_), .D(new_new_n1006_), .Y(new_new_n1011_));
  NA3        g0989(.A(new_new_n1011_), .B(new_new_n1003_), .C(new_new_n997_), .Y(new_new_n1012_));
  INV        g0990(.A(new_new_n630_), .Y(new_new_n1013_));
  NO3        g0991(.A(new_new_n1013_), .B(new_new_n570_), .C(new_new_n347_), .Y(new_new_n1014_));
  NO2        g0992(.A(new_new_n85_), .B(i_5_), .Y(new_new_n1015_));
  NA3        g0993(.A(new_new_n852_), .B(new_new_n109_), .C(new_new_n124_), .Y(new_new_n1016_));
  INV        g0994(.A(new_new_n1016_), .Y(new_new_n1017_));
  AOI210     g0995(.A0(new_new_n1017_), .A1(new_new_n1015_), .B0(new_new_n1014_), .Y(new_new_n1018_));
  NA3        g0996(.A(new_new_n306_), .B(i_5_), .C(new_new_n193_), .Y(new_new_n1019_));
  NAi31      g0997(.An(new_new_n243_), .B(new_new_n1019_), .C(new_new_n244_), .Y(new_new_n1020_));
  NO4        g0998(.A(new_new_n241_), .B(new_new_n211_), .C(i_0_), .D(i_12_), .Y(new_new_n1021_));
  AOI220     g0999(.A0(new_new_n1021_), .A1(new_new_n1020_), .B0(new_new_n802_), .B1(new_new_n175_), .Y(new_new_n1022_));
  AN2        g1000(.A(new_new_n895_), .B(new_new_n153_), .Y(new_new_n1023_));
  NO4        g1001(.A(new_new_n1023_), .B(i_12_), .C(new_new_n661_), .D(new_new_n131_), .Y(new_new_n1024_));
  NA2        g1002(.A(new_new_n1024_), .B(new_new_n220_), .Y(new_new_n1025_));
  NA3        g1003(.A(new_new_n97_), .B(new_new_n584_), .C(i_11_), .Y(new_new_n1026_));
  NO2        g1004(.A(new_new_n1026_), .B(new_new_n155_), .Y(new_new_n1027_));
  NA2        g1005(.A(new_new_n927_), .B(new_new_n480_), .Y(new_new_n1028_));
  OAI220     g1006(.A0(i_7_), .A1(new_new_n1019_), .B0(new_new_n1028_), .B1(new_new_n688_), .Y(new_new_n1029_));
  AOI210     g1007(.A0(new_new_n1029_), .A1(new_new_n913_), .B0(new_new_n1027_), .Y(new_new_n1030_));
  NA4        g1008(.A(new_new_n1030_), .B(new_new_n1025_), .C(new_new_n1022_), .D(new_new_n1018_), .Y(new_new_n1031_));
  NO4        g1009(.A(new_new_n1031_), .B(new_new_n1012_), .C(new_new_n992_), .D(new_new_n979_), .Y(new_new_n1032_));
  NA3        g1010(.A(new_new_n921_), .B(new_new_n371_), .C(i_5_), .Y(new_new_n1033_));
  NA2        g1011(.A(new_new_n1033_), .B(new_new_n1079_), .Y(new_new_n1034_));
  NA2        g1012(.A(new_new_n1034_), .B(new_new_n207_), .Y(new_new_n1035_));
  NA2        g1013(.A(new_new_n186_), .B(new_new_n188_), .Y(new_new_n1036_));
  AO210      g1014(.A0(i_11_), .A1(new_new_n33_), .B0(new_new_n1036_), .Y(new_new_n1037_));
  OAI210     g1015(.A0(new_new_n630_), .A1(new_new_n628_), .B0(new_new_n319_), .Y(new_new_n1038_));
  NA2        g1016(.A(new_new_n1038_), .B(new_new_n1037_), .Y(new_new_n1039_));
  NO4        g1017(.A(new_new_n234_), .B(new_new_n145_), .C(new_new_n691_), .D(new_new_n37_), .Y(new_new_n1040_));
  NO2        g1018(.A(new_new_n1040_), .B(new_new_n888_), .Y(new_new_n1041_));
  OAI210     g1019(.A0(new_new_n1026_), .A1(new_new_n148_), .B0(new_new_n1041_), .Y(new_new_n1042_));
  AOI210     g1020(.A0(new_new_n1039_), .A1(new_new_n49_), .B0(new_new_n1042_), .Y(new_new_n1043_));
  AOI210     g1021(.A0(new_new_n1043_), .A1(new_new_n1035_), .B0(new_new_n73_), .Y(new_new_n1044_));
  NO2        g1022(.A(new_new_n577_), .B(new_new_n382_), .Y(new_new_n1045_));
  NO2        g1023(.A(new_new_n1045_), .B(new_new_n766_), .Y(new_new_n1046_));
  OAI210     g1024(.A0(new_new_n80_), .A1(new_new_n55_), .B0(new_new_n107_), .Y(new_new_n1047_));
  NA2        g1025(.A(new_new_n1047_), .B(new_new_n76_), .Y(new_new_n1048_));
  AOI210     g1026(.A0(new_new_n998_), .A1(new_new_n909_), .B0(new_new_n928_), .Y(new_new_n1049_));
  AOI210     g1027(.A0(new_new_n1049_), .A1(new_new_n1048_), .B0(new_new_n691_), .Y(new_new_n1050_));
  NA2        g1028(.A(new_new_n259_), .B(new_new_n57_), .Y(new_new_n1051_));
  AOI220     g1029(.A0(new_new_n1051_), .A1(new_new_n76_), .B0(new_new_n348_), .B1(new_new_n256_), .Y(new_new_n1052_));
  NO2        g1030(.A(new_new_n1052_), .B(new_new_n238_), .Y(new_new_n1053_));
  NA3        g1031(.A(new_new_n95_), .B(new_new_n308_), .C(new_new_n31_), .Y(new_new_n1054_));
  INV        g1032(.A(new_new_n1054_), .Y(new_new_n1055_));
  NO3        g1033(.A(new_new_n1055_), .B(new_new_n1053_), .C(new_new_n1050_), .Y(new_new_n1056_));
  OAI210     g1034(.A0(new_new_n267_), .A1(new_new_n158_), .B0(new_new_n88_), .Y(new_new_n1057_));
  NA3        g1035(.A(new_new_n770_), .B(new_new_n290_), .C(new_new_n80_), .Y(new_new_n1058_));
  AOI210     g1036(.A0(new_new_n1058_), .A1(new_new_n1057_), .B0(i_11_), .Y(new_new_n1059_));
  NA2        g1037(.A(new_new_n623_), .B(new_new_n217_), .Y(new_new_n1060_));
  OAI210     g1038(.A0(new_new_n1060_), .A1(new_new_n921_), .B0(new_new_n207_), .Y(new_new_n1061_));
  NA2        g1039(.A(new_new_n164_), .B(i_5_), .Y(new_new_n1062_));
  NO2        g1040(.A(new_new_n1061_), .B(new_new_n1062_), .Y(new_new_n1063_));
  NO3        g1041(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n1064_));
  OAI210     g1042(.A0(new_new_n932_), .A1(new_new_n308_), .B0(new_new_n1064_), .Y(new_new_n1065_));
  NO2        g1043(.A(new_new_n1065_), .B(new_new_n736_), .Y(new_new_n1066_));
  NO4        g1044(.A(new_new_n955_), .B(new_new_n486_), .C(new_new_n255_), .D(new_new_n254_), .Y(new_new_n1067_));
  NO2        g1045(.A(new_new_n1067_), .B(new_new_n574_), .Y(new_new_n1068_));
  INV        g1046(.A(new_new_n364_), .Y(new_new_n1069_));
  AOI210     g1047(.A0(new_new_n1069_), .A1(new_new_n1068_), .B0(new_new_n41_), .Y(new_new_n1070_));
  NO4        g1048(.A(new_new_n1070_), .B(new_new_n1066_), .C(new_new_n1063_), .D(new_new_n1059_), .Y(new_new_n1071_));
  OAI210     g1049(.A0(new_new_n1056_), .A1(i_4_), .B0(new_new_n1071_), .Y(new_new_n1072_));
  NO3        g1050(.A(new_new_n1072_), .B(new_new_n1046_), .C(new_new_n1044_), .Y(new_new_n1073_));
  NA4        g1051(.A(new_new_n1073_), .B(new_new_n1032_), .C(new_new_n962_), .D(new_new_n876_), .Y(men4));
  INV        g1052(.A(i_2_), .Y(new_new_n1077_));
  INV        g1053(.A(new_new_n82_), .Y(new_new_n1078_));
  INV        g1054(.A(new_new_n161_), .Y(new_new_n1079_));
  INV        g1055(.A(new_new_n496_), .Y(new_new_n1080_));
endmodule


