library verilog;
use verilog.vl_types.all;
entity sumsub_vlg_vec_tst is
end sumsub_vlg_vec_tst;
