//Benchmark atmr_intb_466_0.125

module atmr_intb(x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14, z0, z1, z2, z3, z4, z5, z6);
 input x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13, x14;
 output z0, z1, z2, z3, z4, z5, z6;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n41_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n107_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n111_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n248_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n257_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n43_, mai_mai_n44_, mai_mai_n45_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n125_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n129_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n335_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n42_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n130_, men_men_n131_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n378_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n451_, ori00, mai00, men00, ori01, mai01, men01, ori02, mai02, men02, ori03, mai03, men03, ori04, mai04, men04, ori05, mai05, men05, ori06, mai06, men06;
  INV        o000(.A(x11), .Y(ori_ori_n23_));
  NA2        o001(.A(ori_ori_n23_), .B(x02), .Y(ori_ori_n24_));
  NA2        o002(.A(x11), .B(x03), .Y(ori_ori_n25_));
  NA2        o003(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n26_));
  NA2        o004(.A(ori_ori_n26_), .B(x07), .Y(ori_ori_n27_));
  INV        o005(.A(x02), .Y(ori_ori_n28_));
  INV        o006(.A(x10), .Y(ori_ori_n29_));
  NA2        o007(.A(ori_ori_n29_), .B(ori_ori_n28_), .Y(ori_ori_n30_));
  INV        o008(.A(x03), .Y(ori_ori_n31_));
  NA2        o009(.A(x10), .B(ori_ori_n31_), .Y(ori_ori_n32_));
  NA3        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .C(x06), .Y(ori_ori_n33_));
  NA2        o011(.A(ori_ori_n33_), .B(ori_ori_n27_), .Y(ori_ori_n34_));
  INV        o012(.A(x04), .Y(ori_ori_n35_));
  INV        o013(.A(x08), .Y(ori_ori_n36_));
  NA2        o014(.A(ori_ori_n36_), .B(x02), .Y(ori_ori_n37_));
  NA2        o015(.A(x08), .B(x03), .Y(ori_ori_n38_));
  AOI210     o016(.A0(ori_ori_n38_), .A1(ori_ori_n37_), .B0(ori_ori_n35_), .Y(ori_ori_n39_));
  NA2        o017(.A(x09), .B(ori_ori_n31_), .Y(ori_ori_n40_));
  INV        o018(.A(x05), .Y(ori_ori_n41_));
  NO2        o019(.A(x09), .B(x02), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(ori_ori_n41_), .Y(ori_ori_n43_));
  NA2        o021(.A(ori_ori_n43_), .B(ori_ori_n40_), .Y(ori_ori_n44_));
  INV        o022(.A(ori_ori_n44_), .Y(ori_ori_n45_));
  NO3        o023(.A(ori_ori_n45_), .B(ori_ori_n39_), .C(ori_ori_n34_), .Y(ori00));
  INV        o024(.A(x01), .Y(ori_ori_n47_));
  INV        o025(.A(x06), .Y(ori_ori_n48_));
  NA2        o026(.A(ori_ori_n48_), .B(ori_ori_n28_), .Y(ori_ori_n49_));
  INV        o027(.A(x09), .Y(ori_ori_n50_));
  NO2        o028(.A(x10), .B(x02), .Y(ori_ori_n51_));
  NOi21      o029(.An(x01), .B(x09), .Y(ori_ori_n52_));
  INV        o030(.A(x00), .Y(ori_ori_n53_));
  NO2        o031(.A(ori_ori_n50_), .B(ori_ori_n53_), .Y(ori_ori_n54_));
  NO2        o032(.A(ori_ori_n54_), .B(ori_ori_n52_), .Y(ori_ori_n55_));
  NA2        o033(.A(x09), .B(ori_ori_n53_), .Y(ori_ori_n56_));
  INV        o034(.A(x07), .Y(ori_ori_n57_));
  INV        o035(.A(ori_ori_n55_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n29_), .B(x02), .Y(ori_ori_n59_));
  NA2        o037(.A(ori_ori_n59_), .B(ori_ori_n24_), .Y(ori_ori_n60_));
  NO2        o038(.A(ori_ori_n60_), .B(ori_ori_n58_), .Y(ori_ori_n61_));
  NA2        o039(.A(ori_ori_n57_), .B(ori_ori_n48_), .Y(ori_ori_n62_));
  OAI210     o040(.A0(ori_ori_n30_), .A1(x11), .B0(ori_ori_n62_), .Y(ori_ori_n63_));
  AOI220     o041(.A0(ori_ori_n63_), .A1(ori_ori_n55_), .B0(ori_ori_n61_), .B1(ori_ori_n31_), .Y(ori_ori_n64_));
  NO2        o042(.A(ori_ori_n64_), .B(x05), .Y(ori_ori_n65_));
  NA2        o043(.A(x09), .B(x05), .Y(ori_ori_n66_));
  NA2        o044(.A(x10), .B(x06), .Y(ori_ori_n67_));
  NOi31      o045(.An(x08), .B(x04), .C(x00), .Y(ori_ori_n68_));
  NO2        o046(.A(ori_ori_n36_), .B(x00), .Y(ori_ori_n69_));
  NO2        o047(.A(x08), .B(x01), .Y(ori_ori_n70_));
  OAI210     o048(.A0(ori_ori_n70_), .A1(ori_ori_n69_), .B0(ori_ori_n35_), .Y(ori_ori_n71_));
  NA2        o049(.A(ori_ori_n50_), .B(ori_ori_n36_), .Y(ori_ori_n72_));
  NO2        o050(.A(ori_ori_n71_), .B(x02), .Y(ori_ori_n73_));
  AN2        o051(.A(ori_ori_n73_), .B(ori_ori_n284_), .Y(ori_ori_n74_));
  INV        o052(.A(ori_ori_n71_), .Y(ori_ori_n75_));
  NA2        o053(.A(x11), .B(x00), .Y(ori_ori_n76_));
  NO2        o054(.A(x11), .B(ori_ori_n47_), .Y(ori_ori_n77_));
  NOi21      o055(.An(ori_ori_n76_), .B(ori_ori_n77_), .Y(ori_ori_n78_));
  NOi21      o056(.An(x01), .B(x10), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n29_), .B(ori_ori_n53_), .Y(ori_ori_n80_));
  NO3        o058(.A(ori_ori_n80_), .B(ori_ori_n79_), .C(x06), .Y(ori_ori_n81_));
  NA2        o059(.A(ori_ori_n81_), .B(ori_ori_n27_), .Y(ori_ori_n82_));
  OAI210     o060(.A0(ori_ori_n281_), .A1(x07), .B0(ori_ori_n82_), .Y(ori_ori_n83_));
  NO3        o061(.A(ori_ori_n83_), .B(ori_ori_n74_), .C(ori_ori_n65_), .Y(ori01));
  INV        o062(.A(x12), .Y(ori_ori_n85_));
  INV        o063(.A(x13), .Y(ori_ori_n86_));
  NO2        o064(.A(x10), .B(x01), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n29_), .B(x00), .Y(ori_ori_n88_));
  NO2        o066(.A(ori_ori_n88_), .B(ori_ori_n87_), .Y(ori_ori_n89_));
  NA2        o067(.A(x04), .B(ori_ori_n28_), .Y(ori_ori_n90_));
  NO2        o068(.A(ori_ori_n52_), .B(x05), .Y(ori_ori_n91_));
  NOi21      o069(.An(ori_ori_n91_), .B(ori_ori_n54_), .Y(ori_ori_n92_));
  NA2        o070(.A(x13), .B(ori_ori_n35_), .Y(ori_ori_n93_));
  NO2        o071(.A(ori_ori_n93_), .B(x05), .Y(ori_ori_n94_));
  NA2        o072(.A(ori_ori_n35_), .B(ori_ori_n53_), .Y(ori_ori_n95_));
  NA2        o073(.A(ori_ori_n29_), .B(ori_ori_n47_), .Y(ori_ori_n96_));
  NA2        o074(.A(x10), .B(ori_ori_n53_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n97_), .B(ori_ori_n96_), .Y(ori_ori_n98_));
  NA2        o076(.A(ori_ori_n50_), .B(x05), .Y(ori_ori_n99_));
  NO2        o077(.A(ori_ori_n56_), .B(x05), .Y(ori_ori_n100_));
  INV        o078(.A(ori_ori_n98_), .Y(ori_ori_n101_));
  NO3        o079(.A(ori_ori_n101_), .B(x06), .C(x03), .Y(ori_ori_n102_));
  INV        o080(.A(ori_ori_n102_), .Y(ori_ori_n103_));
  OAI210     o081(.A0(ori_ori_n70_), .A1(x13), .B0(ori_ori_n35_), .Y(ori_ori_n104_));
  NO2        o082(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n105_));
  NA2        o083(.A(ori_ori_n29_), .B(x06), .Y(ori_ori_n106_));
  NO2        o084(.A(x09), .B(x05), .Y(ori_ori_n107_));
  NA2        o085(.A(ori_ori_n107_), .B(ori_ori_n47_), .Y(ori_ori_n108_));
  NO2        o086(.A(ori_ori_n89_), .B(ori_ori_n49_), .Y(ori_ori_n109_));
  NA2        o087(.A(x09), .B(x00), .Y(ori_ori_n110_));
  NA2        o088(.A(ori_ori_n91_), .B(ori_ori_n110_), .Y(ori_ori_n111_));
  INV        o089(.A(ori_ori_n109_), .Y(ori_ori_n112_));
  NO2        o090(.A(x03), .B(x02), .Y(ori_ori_n113_));
  NA2        o091(.A(ori_ori_n71_), .B(ori_ori_n86_), .Y(ori_ori_n114_));
  OAI210     o092(.A0(ori_ori_n114_), .A1(ori_ori_n92_), .B0(ori_ori_n113_), .Y(ori_ori_n115_));
  OA210      o093(.A0(ori_ori_n112_), .A1(x11), .B0(ori_ori_n115_), .Y(ori_ori_n116_));
  OAI210     o094(.A0(ori_ori_n103_), .A1(ori_ori_n23_), .B0(ori_ori_n116_), .Y(ori_ori_n117_));
  NO2        o095(.A(ori_ori_n29_), .B(x03), .Y(ori_ori_n118_));
  NA2        o096(.A(ori_ori_n86_), .B(x01), .Y(ori_ori_n119_));
  NO2        o097(.A(ori_ori_n119_), .B(x08), .Y(ori_ori_n120_));
  NO2        o098(.A(ori_ori_n118_), .B(ori_ori_n48_), .Y(ori_ori_n121_));
  AOI210     o099(.A0(x11), .A1(ori_ori_n31_), .B0(ori_ori_n28_), .Y(ori_ori_n122_));
  NA2        o100(.A(ori_ori_n121_), .B(ori_ori_n122_), .Y(ori_ori_n123_));
  NA2        o101(.A(x10), .B(x05), .Y(ori_ori_n124_));
  NO2        o102(.A(x09), .B(x01), .Y(ori_ori_n125_));
  INV        o103(.A(ori_ori_n80_), .Y(ori_ori_n126_));
  NOi21      o104(.An(x09), .B(x00), .Y(ori_ori_n127_));
  NO3        o105(.A(ori_ori_n69_), .B(ori_ori_n127_), .C(ori_ori_n47_), .Y(ori_ori_n128_));
  NA2        o106(.A(ori_ori_n128_), .B(ori_ori_n97_), .Y(ori_ori_n129_));
  NA2        o107(.A(x06), .B(x05), .Y(ori_ori_n130_));
  OAI210     o108(.A0(ori_ori_n130_), .A1(ori_ori_n35_), .B0(ori_ori_n85_), .Y(ori_ori_n131_));
  AOI210     o109(.A0(x10), .A1(ori_ori_n54_), .B0(ori_ori_n131_), .Y(ori_ori_n132_));
  NA2        o110(.A(ori_ori_n132_), .B(ori_ori_n129_), .Y(ori_ori_n133_));
  NO2        o111(.A(ori_ori_n86_), .B(x12), .Y(ori_ori_n134_));
  NA2        o112(.A(ori_ori_n25_), .B(ori_ori_n24_), .Y(ori_ori_n135_));
  NO2        o113(.A(ori_ori_n35_), .B(ori_ori_n31_), .Y(ori_ori_n136_));
  NA2        o114(.A(ori_ori_n136_), .B(x02), .Y(ori_ori_n137_));
  NA2        o115(.A(ori_ori_n135_), .B(ori_ori_n133_), .Y(ori_ori_n138_));
  NA2        o116(.A(ori_ori_n138_), .B(ori_ori_n123_), .Y(ori_ori_n139_));
  AOI210     o117(.A0(ori_ori_n117_), .A1(ori_ori_n85_), .B0(ori_ori_n139_), .Y(ori_ori_n140_));
  NA2        o118(.A(ori_ori_n50_), .B(ori_ori_n47_), .Y(ori_ori_n141_));
  NA2        o119(.A(ori_ori_n141_), .B(ori_ori_n104_), .Y(ori_ori_n142_));
  NO2        o120(.A(x06), .B(x05), .Y(ori_ori_n143_));
  NO2        o121(.A(ori_ori_n96_), .B(x06), .Y(ori_ori_n144_));
  AOI210     o122(.A0(ori_ori_n143_), .A1(ori_ori_n142_), .B0(ori_ori_n144_), .Y(ori_ori_n145_));
  NO2        o123(.A(ori_ori_n145_), .B(x12), .Y(ori_ori_n146_));
  INV        o124(.A(ori_ori_n68_), .Y(ori_ori_n147_));
  NO2        o125(.A(ori_ori_n79_), .B(x06), .Y(ori_ori_n148_));
  NO2        o126(.A(ori_ori_n148_), .B(ori_ori_n41_), .Y(ori_ori_n149_));
  INV        o127(.A(ori_ori_n106_), .Y(ori_ori_n150_));
  OAI210     o128(.A0(ori_ori_n150_), .A1(ori_ori_n149_), .B0(x02), .Y(ori_ori_n151_));
  AOI210     o129(.A0(ori_ori_n151_), .A1(ori_ori_n53_), .B0(ori_ori_n23_), .Y(ori_ori_n152_));
  OAI210     o130(.A0(ori_ori_n146_), .A1(ori_ori_n53_), .B0(ori_ori_n152_), .Y(ori_ori_n153_));
  INV        o131(.A(ori_ori_n106_), .Y(ori_ori_n154_));
  NO2        o132(.A(ori_ori_n50_), .B(x03), .Y(ori_ori_n155_));
  NO2        o133(.A(ori_ori_n86_), .B(x03), .Y(ori_ori_n156_));
  NO3        o134(.A(x13), .B(ori_ori_n68_), .C(ori_ori_n127_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n157_), .B(x05), .Y(ori_ori_n158_));
  INV        o136(.A(ori_ori_n77_), .Y(ori_ori_n159_));
  NO2        o137(.A(ori_ori_n159_), .B(x12), .Y(ori_ori_n160_));
  NA2        o138(.A(ori_ori_n23_), .B(ori_ori_n47_), .Y(ori_ori_n161_));
  NA2        o139(.A(ori_ori_n29_), .B(ori_ori_n48_), .Y(ori_ori_n162_));
  INV        o140(.A(x03), .Y(ori_ori_n163_));
  OR2        o141(.A(ori_ori_n163_), .B(ori_ori_n67_), .Y(ori_ori_n164_));
  NA2        o142(.A(x13), .B(ori_ori_n85_), .Y(ori_ori_n165_));
  NA3        o143(.A(ori_ori_n165_), .B(ori_ori_n131_), .C(ori_ori_n78_), .Y(ori_ori_n166_));
  OAI210     o144(.A0(ori_ori_n164_), .A1(ori_ori_n161_), .B0(ori_ori_n166_), .Y(ori_ori_n167_));
  AOI210     o145(.A0(ori_ori_n160_), .A1(ori_ori_n158_), .B0(ori_ori_n167_), .Y(ori_ori_n168_));
  AOI210     o146(.A0(ori_ori_n168_), .A1(ori_ori_n153_), .B0(x07), .Y(ori_ori_n169_));
  NA2        o147(.A(ori_ori_n66_), .B(ori_ori_n29_), .Y(ori_ori_n170_));
  NO2        o148(.A(x12), .B(x02), .Y(ori_ori_n171_));
  NA2        o149(.A(ori_ori_n50_), .B(ori_ori_n41_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n172_), .B(x01), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n86_), .B(x04), .Y(ori_ori_n174_));
  NO2        o152(.A(x02), .B(ori_ori_n282_), .Y(ori_ori_n175_));
  NO3        o153(.A(ori_ori_n76_), .B(x12), .C(x03), .Y(ori_ori_n176_));
  NA2        o154(.A(ori_ori_n175_), .B(ori_ori_n176_), .Y(ori_ori_n177_));
  NOi21      o155(.An(ori_ori_n170_), .B(ori_ori_n148_), .Y(ori_ori_n178_));
  NO2        o156(.A(ori_ori_n25_), .B(x00), .Y(ori_ori_n179_));
  NA2        o157(.A(ori_ori_n178_), .B(ori_ori_n179_), .Y(ori_ori_n180_));
  NO2        o158(.A(ori_ori_n285_), .B(ori_ori_n126_), .Y(ori_ori_n181_));
  NO2        o159(.A(ori_ori_n161_), .B(ori_ori_n28_), .Y(ori_ori_n182_));
  OAI210     o160(.A0(ori_ori_n181_), .A1(ori_ori_n154_), .B0(ori_ori_n182_), .Y(ori_ori_n183_));
  NA3        o161(.A(ori_ori_n183_), .B(ori_ori_n180_), .C(ori_ori_n177_), .Y(ori_ori_n184_));
  NO2        o162(.A(ori_ori_n184_), .B(ori_ori_n169_), .Y(ori_ori_n185_));
  OAI210     o163(.A0(ori_ori_n140_), .A1(ori_ori_n57_), .B0(ori_ori_n185_), .Y(ori02));
  NOi21      o164(.An(ori_ori_n157_), .B(ori_ori_n125_), .Y(ori_ori_n187_));
  NO2        o165(.A(ori_ori_n187_), .B(ori_ori_n32_), .Y(ori_ori_n188_));
  NA2        o166(.A(ori_ori_n188_), .B(ori_ori_n124_), .Y(ori_ori_n189_));
  NA2        o167(.A(ori_ori_n114_), .B(ori_ori_n113_), .Y(ori_ori_n190_));
  AOI210     o168(.A0(ori_ori_n190_), .A1(ori_ori_n189_), .B0(ori_ori_n48_), .Y(ori_ori_n191_));
  NO2        o169(.A(x05), .B(x02), .Y(ori_ori_n192_));
  OAI210     o170(.A0(ori_ori_n142_), .A1(ori_ori_n127_), .B0(ori_ori_n192_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n193_), .B(ori_ori_n106_), .Y(ori_ori_n194_));
  NO2        o172(.A(ori_ori_n162_), .B(ori_ori_n47_), .Y(ori_ori_n195_));
  NA2        o173(.A(ori_ori_n195_), .B(ori_ori_n158_), .Y(ori_ori_n196_));
  OAI210     o174(.A0(ori_ori_n42_), .A1(ori_ori_n41_), .B0(ori_ori_n48_), .Y(ori_ori_n197_));
  BUFFER     o175(.A(ori_ori_n108_), .Y(ori_ori_n198_));
  AOI210     o176(.A0(ori_ori_n198_), .A1(ori_ori_n104_), .B0(ori_ori_n197_), .Y(ori_ori_n199_));
  NA2        o177(.A(ori_ori_n199_), .B(ori_ori_n80_), .Y(ori_ori_n200_));
  INV        o178(.A(ori_ori_n113_), .Y(ori_ori_n201_));
  NO2        o179(.A(ori_ori_n201_), .B(ori_ori_n98_), .Y(ori_ori_n202_));
  NA2        o180(.A(ori_ori_n202_), .B(x13), .Y(ori_ori_n203_));
  NA3        o181(.A(ori_ori_n203_), .B(ori_ori_n200_), .C(ori_ori_n196_), .Y(ori_ori_n204_));
  NO3        o182(.A(ori_ori_n204_), .B(ori_ori_n194_), .C(ori_ori_n191_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n105_), .B(x03), .Y(ori_ori_n206_));
  INV        o184(.A(ori_ori_n206_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n207_), .B(ori_ori_n87_), .Y(ori_ori_n208_));
  NO2        o186(.A(ori_ori_n99_), .B(ori_ori_n28_), .Y(ori_ori_n209_));
  NA2        o187(.A(ori_ori_n209_), .B(ori_ori_n88_), .Y(ori_ori_n210_));
  NA2        o188(.A(ori_ori_n174_), .B(ori_ori_n85_), .Y(ori_ori_n211_));
  NA2        o189(.A(ori_ori_n85_), .B(ori_ori_n41_), .Y(ori_ori_n212_));
  NA3        o190(.A(ori_ori_n212_), .B(ori_ori_n211_), .C(ori_ori_n98_), .Y(ori_ori_n213_));
  NA4        o191(.A(ori_ori_n213_), .B(ori_ori_n210_), .C(ori_ori_n208_), .D(ori_ori_n48_), .Y(ori_ori_n214_));
  INV        o192(.A(ori_ori_n136_), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n32_), .B(x05), .Y(ori_ori_n216_));
  OAI210     o194(.A0(ori_ori_n215_), .A1(ori_ori_n55_), .B0(ori_ori_n216_), .Y(ori_ori_n217_));
  NA2        o195(.A(ori_ori_n217_), .B(x02), .Y(ori_ori_n218_));
  NA2        o196(.A(ori_ori_n134_), .B(x04), .Y(ori_ori_n219_));
  NO3        o197(.A(ori_ori_n134_), .B(ori_ori_n118_), .C(ori_ori_n51_), .Y(ori_ori_n220_));
  OAI210     o198(.A0(x12), .A1(ori_ori_n128_), .B0(ori_ori_n220_), .Y(ori_ori_n221_));
  NA3        o199(.A(ori_ori_n221_), .B(ori_ori_n218_), .C(x06), .Y(ori_ori_n222_));
  NA2        o200(.A(x09), .B(x03), .Y(ori_ori_n223_));
  OAI220     o201(.A0(ori_ori_n223_), .A1(ori_ori_n97_), .B0(ori_ori_n141_), .B1(ori_ori_n59_), .Y(ori_ori_n224_));
  AN2        o202(.A(ori_ori_n224_), .B(x05), .Y(ori_ori_n225_));
  AOI210     o203(.A0(ori_ori_n222_), .A1(ori_ori_n214_), .B0(ori_ori_n225_), .Y(ori_ori_n226_));
  OAI210     o204(.A0(ori_ori_n205_), .A1(x12), .B0(ori_ori_n226_), .Y(ori03));
  OR2        o205(.A(ori_ori_n42_), .B(ori_ori_n155_), .Y(ori_ori_n228_));
  AOI210     o206(.A0(ori_ori_n114_), .A1(ori_ori_n85_), .B0(ori_ori_n228_), .Y(ori_ori_n229_));
  OR2        o207(.A(ori_ori_n72_), .B(ori_ori_n219_), .Y(ori_ori_n230_));
  NA2        o208(.A(ori_ori_n134_), .B(ori_ori_n113_), .Y(ori_ori_n231_));
  NA3        o209(.A(ori_ori_n231_), .B(ori_ori_n230_), .C(ori_ori_n137_), .Y(ori_ori_n232_));
  OAI210     o210(.A0(ori_ori_n232_), .A1(ori_ori_n229_), .B0(x05), .Y(ori_ori_n233_));
  NA2        o211(.A(ori_ori_n228_), .B(x05), .Y(ori_ori_n234_));
  AOI210     o212(.A0(ori_ori_n104_), .A1(ori_ori_n147_), .B0(ori_ori_n234_), .Y(ori_ori_n235_));
  AOI210     o213(.A0(ori_ori_n156_), .A1(ori_ori_n283_), .B0(ori_ori_n94_), .Y(ori_ori_n236_));
  NO2        o214(.A(ori_ori_n236_), .B(ori_ori_n55_), .Y(ori_ori_n237_));
  OAI210     o215(.A0(ori_ori_n237_), .A1(ori_ori_n235_), .B0(ori_ori_n85_), .Y(ori_ori_n238_));
  AOI210     o216(.A0(ori_ori_n108_), .A1(ori_ori_n56_), .B0(ori_ori_n38_), .Y(ori_ori_n239_));
  NO2        o217(.A(ori_ori_n125_), .B(ori_ori_n100_), .Y(ori_ori_n240_));
  OAI220     o218(.A0(ori_ori_n240_), .A1(ori_ori_n37_), .B0(ori_ori_n111_), .B1(x13), .Y(ori_ori_n241_));
  OAI210     o219(.A0(ori_ori_n241_), .A1(ori_ori_n239_), .B0(x04), .Y(ori_ori_n242_));
  NO3        o220(.A(ori_ori_n212_), .B(ori_ori_n71_), .C(ori_ori_n55_), .Y(ori_ori_n243_));
  NO2        o221(.A(ori_ori_n85_), .B(ori_ori_n108_), .Y(ori_ori_n244_));
  OA210      o222(.A0(ori_ori_n120_), .A1(x12), .B0(ori_ori_n100_), .Y(ori_ori_n245_));
  NO3        o223(.A(ori_ori_n245_), .B(ori_ori_n244_), .C(ori_ori_n243_), .Y(ori_ori_n246_));
  NA4        o224(.A(ori_ori_n246_), .B(ori_ori_n242_), .C(ori_ori_n238_), .D(ori_ori_n233_), .Y(ori04));
  NO2        o225(.A(ori_ori_n75_), .B(ori_ori_n39_), .Y(ori_ori_n248_));
  XO2        o226(.A(ori_ori_n248_), .B(ori_ori_n165_), .Y(ori05));
  OAI210     o227(.A0(ori_ori_n26_), .A1(ori_ori_n85_), .B0(x07), .Y(ori_ori_n250_));
  INV        o228(.A(ori_ori_n250_), .Y(ori_ori_n251_));
  NA2        o229(.A(x00), .B(ori_ori_n161_), .Y(ori_ori_n252_));
  NA2        o230(.A(ori_ori_n252_), .B(ori_ori_n85_), .Y(ori_ori_n253_));
  NA2        o231(.A(ori_ori_n33_), .B(ori_ori_n85_), .Y(ori_ori_n254_));
  AOI210     o232(.A0(ori_ori_n254_), .A1(ori_ori_n77_), .B0(x07), .Y(ori_ori_n255_));
  AOI210     o233(.A0(ori_ori_n255_), .A1(ori_ori_n253_), .B0(ori_ori_n251_), .Y(ori_ori_n256_));
  AOI210     o234(.A0(ori_ori_n219_), .A1(ori_ori_n90_), .B0(ori_ori_n171_), .Y(ori_ori_n257_));
  NOi21      o235(.An(ori_ori_n206_), .B(ori_ori_n100_), .Y(ori_ori_n258_));
  OAI210     o236(.A0(x12), .A1(ori_ori_n47_), .B0(ori_ori_n35_), .Y(ori_ori_n259_));
  AOI210     o237(.A0(ori_ori_n165_), .A1(ori_ori_n47_), .B0(ori_ori_n259_), .Y(ori_ori_n260_));
  NO3        o238(.A(ori_ori_n260_), .B(ori_ori_n257_), .C(x08), .Y(ori_ori_n261_));
  NO2        o239(.A(ori_ori_n99_), .B(ori_ori_n28_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n262_), .B(ori_ori_n173_), .Y(ori_ori_n263_));
  NA3        o241(.A(ori_ori_n215_), .B(ori_ori_n95_), .C(x12), .Y(ori_ori_n264_));
  AO210      o242(.A0(ori_ori_n215_), .A1(ori_ori_n95_), .B0(ori_ori_n165_), .Y(ori_ori_n265_));
  NA3        o243(.A(ori_ori_n265_), .B(ori_ori_n264_), .C(x08), .Y(ori_ori_n266_));
  INV        o244(.A(ori_ori_n266_), .Y(ori_ori_n267_));
  NO2        o245(.A(ori_ori_n261_), .B(ori_ori_n267_), .Y(ori_ori_n268_));
  NA3        o246(.A(ori_ori_n263_), .B(ori_ori_n258_), .C(ori_ori_n211_), .Y(ori_ori_n269_));
  INV        o247(.A(x14), .Y(ori_ori_n270_));
  NO2        o248(.A(ori_ori_n119_), .B(ori_ori_n53_), .Y(ori_ori_n271_));
  NO2        o249(.A(ori_ori_n271_), .B(ori_ori_n270_), .Y(ori_ori_n272_));
  NA2        o250(.A(ori_ori_n272_), .B(ori_ori_n269_), .Y(ori_ori_n273_));
  NA2        o251(.A(ori_ori_n254_), .B(ori_ori_n57_), .Y(ori_ori_n274_));
  INV        o252(.A(ori_ori_n111_), .Y(ori_ori_n275_));
  OAI210     o253(.A0(ori_ori_n43_), .A1(ori_ori_n275_), .B0(ori_ori_n85_), .Y(ori_ori_n276_));
  OAI210     o254(.A0(ori_ori_n274_), .A1(ori_ori_n76_), .B0(ori_ori_n276_), .Y(ori_ori_n277_));
  NO4        o255(.A(ori_ori_n277_), .B(ori_ori_n273_), .C(ori_ori_n268_), .D(ori_ori_n256_), .Y(ori06));
  INV        o256(.A(ori_ori_n78_), .Y(ori_ori_n281_));
  INV        o257(.A(x13), .Y(ori_ori_n282_));
  INV        o258(.A(x05), .Y(ori_ori_n283_));
  INV        o259(.A(x03), .Y(ori_ori_n284_));
  INV        o260(.A(x05), .Y(ori_ori_n285_));
  INV        m000(.A(x11), .Y(mai_mai_n23_));
  NA2        m001(.A(mai_mai_n23_), .B(x02), .Y(mai_mai_n24_));
  NA2        m002(.A(x11), .B(x03), .Y(mai_mai_n25_));
  NA2        m003(.A(mai_mai_n25_), .B(mai_mai_n24_), .Y(mai_mai_n26_));
  NA2        m004(.A(mai_mai_n26_), .B(x07), .Y(mai_mai_n27_));
  INV        m005(.A(x02), .Y(mai_mai_n28_));
  INV        m006(.A(x10), .Y(mai_mai_n29_));
  NA2        m007(.A(mai_mai_n29_), .B(mai_mai_n28_), .Y(mai_mai_n30_));
  INV        m008(.A(x03), .Y(mai_mai_n31_));
  NA2        m009(.A(x10), .B(mai_mai_n31_), .Y(mai_mai_n32_));
  NA3        m010(.A(mai_mai_n32_), .B(mai_mai_n30_), .C(x06), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n27_), .Y(mai_mai_n34_));
  INV        m012(.A(x04), .Y(mai_mai_n35_));
  INV        m013(.A(x08), .Y(mai_mai_n36_));
  NA2        m014(.A(mai_mai_n36_), .B(x02), .Y(mai_mai_n37_));
  NA2        m015(.A(x08), .B(x03), .Y(mai_mai_n38_));
  AOI210     m016(.A0(mai_mai_n38_), .A1(mai_mai_n37_), .B0(mai_mai_n35_), .Y(mai_mai_n39_));
  NA2        m017(.A(x09), .B(mai_mai_n31_), .Y(mai_mai_n40_));
  INV        m018(.A(x05), .Y(mai_mai_n41_));
  NO2        m019(.A(x09), .B(x02), .Y(mai_mai_n42_));
  NO2        m020(.A(mai_mai_n42_), .B(mai_mai_n41_), .Y(mai_mai_n43_));
  NA2        m021(.A(mai_mai_n43_), .B(mai_mai_n40_), .Y(mai_mai_n44_));
  INV        m022(.A(mai_mai_n44_), .Y(mai_mai_n45_));
  NO3        m023(.A(mai_mai_n45_), .B(mai_mai_n39_), .C(mai_mai_n34_), .Y(mai00));
  INV        m024(.A(x01), .Y(mai_mai_n47_));
  INV        m025(.A(x06), .Y(mai_mai_n48_));
  NA2        m026(.A(mai_mai_n48_), .B(mai_mai_n28_), .Y(mai_mai_n49_));
  NO3        m027(.A(mai_mai_n49_), .B(x11), .C(x09), .Y(mai_mai_n50_));
  INV        m028(.A(x09), .Y(mai_mai_n51_));
  NO2        m029(.A(x10), .B(x02), .Y(mai_mai_n52_));
  NA2        m030(.A(mai_mai_n52_), .B(mai_mai_n51_), .Y(mai_mai_n53_));
  NO2        m031(.A(mai_mai_n53_), .B(x07), .Y(mai_mai_n54_));
  OAI210     m032(.A0(mai_mai_n54_), .A1(mai_mai_n50_), .B0(mai_mai_n47_), .Y(mai_mai_n55_));
  NOi21      m033(.An(x01), .B(x09), .Y(mai_mai_n56_));
  INV        m034(.A(x00), .Y(mai_mai_n57_));
  NO2        m035(.A(mai_mai_n51_), .B(mai_mai_n57_), .Y(mai_mai_n58_));
  NO2        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .Y(mai_mai_n59_));
  NA2        m037(.A(x09), .B(mai_mai_n57_), .Y(mai_mai_n60_));
  INV        m038(.A(x07), .Y(mai_mai_n61_));
  AOI220     m039(.A0(x11), .A1(mai_mai_n48_), .B0(x10), .B1(mai_mai_n61_), .Y(mai_mai_n62_));
  INV        m040(.A(mai_mai_n59_), .Y(mai_mai_n63_));
  NA2        m041(.A(mai_mai_n29_), .B(x02), .Y(mai_mai_n64_));
  NA2        m042(.A(mai_mai_n64_), .B(mai_mai_n24_), .Y(mai_mai_n65_));
  OAI220     m043(.A0(mai_mai_n65_), .A1(mai_mai_n63_), .B0(mai_mai_n62_), .B1(mai_mai_n60_), .Y(mai_mai_n66_));
  NO2        m044(.A(mai_mai_n30_), .B(x11), .Y(mai_mai_n67_));
  AOI220     m045(.A0(mai_mai_n67_), .A1(mai_mai_n59_), .B0(mai_mai_n66_), .B1(mai_mai_n31_), .Y(mai_mai_n68_));
  AOI210     m046(.A0(mai_mai_n68_), .A1(mai_mai_n55_), .B0(x05), .Y(mai_mai_n69_));
  NO2        m047(.A(mai_mai_n61_), .B(mai_mai_n23_), .Y(mai_mai_n70_));
  NA2        m048(.A(x09), .B(x05), .Y(mai_mai_n71_));
  NA2        m049(.A(x10), .B(x06), .Y(mai_mai_n72_));
  NA3        m050(.A(mai_mai_n72_), .B(mai_mai_n71_), .C(mai_mai_n28_), .Y(mai_mai_n73_));
  OAI210     m051(.A0(mai_mai_n73_), .A1(mai_mai_n70_), .B0(x03), .Y(mai_mai_n74_));
  NOi31      m052(.An(x08), .B(x04), .C(x00), .Y(mai_mai_n75_));
  AOI210     m053(.A0(mai_mai_n379_), .A1(mai_mai_n75_), .B0(mai_mai_n24_), .Y(mai_mai_n76_));
  NO2        m054(.A(x09), .B(mai_mai_n41_), .Y(mai_mai_n77_));
  OAI210     m055(.A0(mai_mai_n77_), .A1(mai_mai_n29_), .B0(x02), .Y(mai_mai_n78_));
  AOI210     m056(.A0(x08), .A1(mai_mai_n48_), .B0(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m057(.A(mai_mai_n36_), .B(x00), .Y(mai_mai_n80_));
  NO2        m058(.A(x08), .B(x01), .Y(mai_mai_n81_));
  OAI210     m059(.A0(mai_mai_n81_), .A1(mai_mai_n80_), .B0(mai_mai_n35_), .Y(mai_mai_n82_));
  NO3        m060(.A(mai_mai_n82_), .B(mai_mai_n79_), .C(mai_mai_n76_), .Y(mai_mai_n83_));
  AN2        m061(.A(mai_mai_n83_), .B(mai_mai_n74_), .Y(mai_mai_n84_));
  INV        m062(.A(mai_mai_n82_), .Y(mai_mai_n85_));
  NO2        m063(.A(x06), .B(x05), .Y(mai_mai_n86_));
  NA2        m064(.A(x11), .B(x00), .Y(mai_mai_n87_));
  NO2        m065(.A(x11), .B(mai_mai_n47_), .Y(mai_mai_n88_));
  NOi21      m066(.An(mai_mai_n87_), .B(mai_mai_n88_), .Y(mai_mai_n89_));
  AOI210     m067(.A0(mai_mai_n86_), .A1(mai_mai_n85_), .B0(mai_mai_n89_), .Y(mai_mai_n90_));
  NO2        m068(.A(mai_mai_n53_), .B(x11), .Y(mai_mai_n91_));
  NOi21      m069(.An(x01), .B(x10), .Y(mai_mai_n92_));
  NO2        m070(.A(mai_mai_n29_), .B(mai_mai_n57_), .Y(mai_mai_n93_));
  NO3        m071(.A(mai_mai_n93_), .B(mai_mai_n92_), .C(x06), .Y(mai_mai_n94_));
  AOI220     m072(.A0(mai_mai_n94_), .A1(mai_mai_n27_), .B0(mai_mai_n91_), .B1(mai_mai_n85_), .Y(mai_mai_n95_));
  OAI210     m073(.A0(mai_mai_n90_), .A1(x07), .B0(mai_mai_n95_), .Y(mai_mai_n96_));
  NO3        m074(.A(mai_mai_n96_), .B(mai_mai_n84_), .C(mai_mai_n69_), .Y(mai01));
  INV        m075(.A(x12), .Y(mai_mai_n98_));
  INV        m076(.A(x13), .Y(mai_mai_n99_));
  NA2        m077(.A(x08), .B(x04), .Y(mai_mai_n100_));
  NA2        m078(.A(mai_mai_n92_), .B(mai_mai_n28_), .Y(mai_mai_n101_));
  NO2        m079(.A(x10), .B(x01), .Y(mai_mai_n102_));
  NO2        m080(.A(mai_mai_n29_), .B(x00), .Y(mai_mai_n103_));
  NO2        m081(.A(mai_mai_n103_), .B(mai_mai_n102_), .Y(mai_mai_n104_));
  NA2        m082(.A(x04), .B(mai_mai_n28_), .Y(mai_mai_n105_));
  NO3        m083(.A(mai_mai_n105_), .B(mai_mai_n36_), .C(mai_mai_n41_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n56_), .B(x05), .Y(mai_mai_n107_));
  NO2        m085(.A(mai_mai_n99_), .B(mai_mai_n36_), .Y(mai_mai_n108_));
  NA3        m086(.A(mai_mai_n108_), .B(x04), .C(x06), .Y(mai_mai_n109_));
  NO2        m087(.A(mai_mai_n109_), .B(mai_mai_n57_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n81_), .B(x13), .Y(mai_mai_n111_));
  NA2        m089(.A(x13), .B(mai_mai_n35_), .Y(mai_mai_n112_));
  NO2        m090(.A(mai_mai_n112_), .B(x05), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n35_), .B(mai_mai_n57_), .Y(mai_mai_n114_));
  AOI210     m092(.A0(x00), .A1(mai_mai_n111_), .B0(mai_mai_n72_), .Y(mai_mai_n115_));
  NA2        m093(.A(mai_mai_n29_), .B(mai_mai_n47_), .Y(mai_mai_n116_));
  NA2        m094(.A(x10), .B(mai_mai_n57_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n117_), .B(mai_mai_n116_), .Y(mai_mai_n118_));
  NA2        m096(.A(mai_mai_n51_), .B(x05), .Y(mai_mai_n119_));
  NO2        m097(.A(mai_mai_n60_), .B(x05), .Y(mai_mai_n120_));
  NO2        m098(.A(x06), .B(x03), .Y(mai_mai_n121_));
  NO4        m099(.A(mai_mai_n121_), .B(mai_mai_n115_), .C(mai_mai_n110_), .D(mai_mai_n106_), .Y(mai_mai_n122_));
  NA2        m100(.A(x13), .B(mai_mai_n36_), .Y(mai_mai_n123_));
  OAI210     m101(.A0(mai_mai_n81_), .A1(x13), .B0(mai_mai_n35_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(mai_mai_n123_), .Y(mai_mai_n125_));
  NO2        m103(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n126_));
  NA2        m104(.A(mai_mai_n29_), .B(x06), .Y(mai_mai_n127_));
  AOI210     m105(.A0(mai_mai_n127_), .A1(mai_mai_n49_), .B0(mai_mai_n126_), .Y(mai_mai_n128_));
  NO2        m106(.A(x09), .B(x05), .Y(mai_mai_n129_));
  NA2        m107(.A(mai_mai_n129_), .B(mai_mai_n47_), .Y(mai_mai_n130_));
  NA2        m108(.A(x09), .B(x00), .Y(mai_mai_n131_));
  NA2        m109(.A(mai_mai_n107_), .B(mai_mai_n131_), .Y(mai_mai_n132_));
  NO2        m110(.A(x03), .B(x02), .Y(mai_mai_n133_));
  NA2        m111(.A(mai_mai_n82_), .B(mai_mai_n99_), .Y(mai_mai_n134_));
  OAI210     m112(.A0(mai_mai_n134_), .A1(mai_mai_n57_), .B0(mai_mai_n133_), .Y(mai_mai_n135_));
  OA210      m113(.A0(mai_mai_n383_), .A1(x11), .B0(mai_mai_n135_), .Y(mai_mai_n136_));
  OAI210     m114(.A0(mai_mai_n122_), .A1(mai_mai_n23_), .B0(mai_mai_n136_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n104_), .B(mai_mai_n40_), .Y(mai_mai_n138_));
  NAi21      m116(.An(x06), .B(x10), .Y(mai_mai_n139_));
  NOi21      m117(.An(x01), .B(x13), .Y(mai_mai_n140_));
  NA2        m118(.A(mai_mai_n140_), .B(mai_mai_n139_), .Y(mai_mai_n141_));
  AOI210     m119(.A0(mai_mai_n141_), .A1(mai_mai_n138_), .B0(mai_mai_n41_), .Y(mai_mai_n142_));
  NO2        m120(.A(mai_mai_n29_), .B(x03), .Y(mai_mai_n143_));
  NA2        m121(.A(mai_mai_n99_), .B(x01), .Y(mai_mai_n144_));
  NO2        m122(.A(mai_mai_n144_), .B(x08), .Y(mai_mai_n145_));
  OAI210     m123(.A0(x05), .A1(mai_mai_n145_), .B0(mai_mai_n51_), .Y(mai_mai_n146_));
  AOI210     m124(.A0(mai_mai_n146_), .A1(mai_mai_n143_), .B0(mai_mai_n48_), .Y(mai_mai_n147_));
  AOI210     m125(.A0(x11), .A1(mai_mai_n31_), .B0(mai_mai_n28_), .Y(mai_mai_n148_));
  OAI210     m126(.A0(mai_mai_n147_), .A1(mai_mai_n142_), .B0(mai_mai_n148_), .Y(mai_mai_n149_));
  NA2        m127(.A(x04), .B(x02), .Y(mai_mai_n150_));
  NA2        m128(.A(x10), .B(x05), .Y(mai_mai_n151_));
  NO2        m129(.A(x09), .B(x01), .Y(mai_mai_n152_));
  NO2        m130(.A(mai_mai_n107_), .B(x08), .Y(mai_mai_n153_));
  NA3        m131(.A(mai_mai_n140_), .B(mai_mai_n139_), .C(mai_mai_n51_), .Y(mai_mai_n154_));
  OAI210     m132(.A0(mai_mai_n387_), .A1(mai_mai_n108_), .B0(mai_mai_n154_), .Y(mai_mai_n155_));
  AOI210     m133(.A0(mai_mai_n153_), .A1(x06), .B0(mai_mai_n155_), .Y(mai_mai_n156_));
  NO2        m134(.A(mai_mai_n156_), .B(x11), .Y(mai_mai_n157_));
  NAi21      m135(.An(mai_mai_n150_), .B(mai_mai_n157_), .Y(mai_mai_n158_));
  INV        m136(.A(mai_mai_n25_), .Y(mai_mai_n159_));
  NAi21      m137(.An(x13), .B(x00), .Y(mai_mai_n160_));
  AOI210     m138(.A0(mai_mai_n29_), .A1(mai_mai_n48_), .B0(mai_mai_n160_), .Y(mai_mai_n161_));
  AOI220     m139(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(mai_mai_n162_));
  OAI210     m140(.A0(mai_mai_n151_), .A1(mai_mai_n35_), .B0(mai_mai_n162_), .Y(mai_mai_n163_));
  AN2        m141(.A(mai_mai_n163_), .B(mai_mai_n161_), .Y(mai_mai_n164_));
  AN2        m142(.A(mai_mai_n72_), .B(mai_mai_n71_), .Y(mai_mai_n165_));
  NO2        m143(.A(mai_mai_n93_), .B(x06), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n160_), .B(mai_mai_n36_), .Y(mai_mai_n167_));
  INV        m145(.A(mai_mai_n167_), .Y(mai_mai_n168_));
  OAI210     m146(.A0(mai_mai_n166_), .A1(mai_mai_n165_), .B0(mai_mai_n168_), .Y(mai_mai_n169_));
  OAI210     m147(.A0(mai_mai_n169_), .A1(mai_mai_n164_), .B0(mai_mai_n159_), .Y(mai_mai_n170_));
  NOi21      m148(.An(x09), .B(x00), .Y(mai_mai_n171_));
  NO3        m149(.A(mai_mai_n80_), .B(mai_mai_n171_), .C(mai_mai_n47_), .Y(mai_mai_n172_));
  INV        m150(.A(mai_mai_n172_), .Y(mai_mai_n173_));
  NA2        m151(.A(x06), .B(x05), .Y(mai_mai_n174_));
  NA2        m152(.A(mai_mai_n98_), .B(mai_mai_n173_), .Y(mai_mai_n175_));
  NO2        m153(.A(mai_mai_n99_), .B(x12), .Y(mai_mai_n176_));
  AOI210     m154(.A0(mai_mai_n25_), .A1(mai_mai_n24_), .B0(mai_mai_n176_), .Y(mai_mai_n177_));
  NA2        m155(.A(mai_mai_n92_), .B(mai_mai_n51_), .Y(mai_mai_n178_));
  NO2        m156(.A(mai_mai_n35_), .B(mai_mai_n31_), .Y(mai_mai_n179_));
  NA2        m157(.A(mai_mai_n179_), .B(x02), .Y(mai_mai_n180_));
  NO2        m158(.A(mai_mai_n180_), .B(mai_mai_n178_), .Y(mai_mai_n181_));
  AOI210     m159(.A0(mai_mai_n177_), .A1(mai_mai_n175_), .B0(mai_mai_n181_), .Y(mai_mai_n182_));
  NA4        m160(.A(mai_mai_n182_), .B(mai_mai_n170_), .C(mai_mai_n158_), .D(mai_mai_n149_), .Y(mai_mai_n183_));
  AOI210     m161(.A0(mai_mai_n137_), .A1(mai_mai_n98_), .B0(mai_mai_n183_), .Y(mai_mai_n184_));
  INV        m162(.A(mai_mai_n73_), .Y(mai_mai_n185_));
  NA2        m163(.A(mai_mai_n185_), .B(mai_mai_n125_), .Y(mai_mai_n186_));
  NA2        m164(.A(mai_mai_n51_), .B(mai_mai_n47_), .Y(mai_mai_n187_));
  NA2        m165(.A(mai_mai_n187_), .B(mai_mai_n124_), .Y(mai_mai_n188_));
  AOI210     m166(.A0(mai_mai_n30_), .A1(x06), .B0(x05), .Y(mai_mai_n189_));
  NO2        m167(.A(mai_mai_n116_), .B(x06), .Y(mai_mai_n190_));
  AOI210     m168(.A0(mai_mai_n189_), .A1(mai_mai_n188_), .B0(mai_mai_n190_), .Y(mai_mai_n191_));
  AOI210     m169(.A0(mai_mai_n191_), .A1(mai_mai_n186_), .B0(x12), .Y(mai_mai_n192_));
  INV        m170(.A(mai_mai_n75_), .Y(mai_mai_n193_));
  NA2        m171(.A(mai_mai_n141_), .B(mai_mai_n57_), .Y(mai_mai_n194_));
  NA2        m172(.A(mai_mai_n194_), .B(mai_mai_n193_), .Y(mai_mai_n195_));
  AOI210     m173(.A0(mai_mai_n36_), .A1(x04), .B0(mai_mai_n51_), .Y(mai_mai_n196_));
  NA2        m174(.A(mai_mai_n56_), .B(x02), .Y(mai_mai_n197_));
  AOI210     m175(.A0(mai_mai_n197_), .A1(mai_mai_n195_), .B0(mai_mai_n23_), .Y(mai_mai_n198_));
  OAI210     m176(.A0(mai_mai_n192_), .A1(mai_mai_n57_), .B0(mai_mai_n198_), .Y(mai_mai_n199_));
  INV        m177(.A(mai_mai_n127_), .Y(mai_mai_n200_));
  NO2        m178(.A(mai_mai_n51_), .B(x03), .Y(mai_mai_n201_));
  OAI210     m179(.A0(mai_mai_n77_), .A1(mai_mai_n36_), .B0(x04), .Y(mai_mai_n202_));
  NO2        m180(.A(mai_mai_n99_), .B(x03), .Y(mai_mai_n203_));
  AOI220     m181(.A0(mai_mai_n203_), .A1(mai_mai_n202_), .B0(mai_mai_n75_), .B1(mai_mai_n201_), .Y(mai_mai_n204_));
  INV        m182(.A(mai_mai_n139_), .Y(mai_mai_n205_));
  NOi21      m183(.An(x13), .B(x04), .Y(mai_mai_n206_));
  NO3        m184(.A(mai_mai_n206_), .B(mai_mai_n75_), .C(mai_mai_n171_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n207_), .B(x05), .Y(mai_mai_n208_));
  NA2        m186(.A(mai_mai_n205_), .B(mai_mai_n57_), .Y(mai_mai_n209_));
  OAI210     m187(.A0(mai_mai_n204_), .A1(mai_mai_n200_), .B0(mai_mai_n209_), .Y(mai_mai_n210_));
  INV        m188(.A(mai_mai_n88_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n211_), .B(x12), .Y(mai_mai_n212_));
  NA2        m190(.A(mai_mai_n23_), .B(mai_mai_n47_), .Y(mai_mai_n213_));
  OAI210     m191(.A0(x08), .A1(mai_mai_n163_), .B0(mai_mai_n161_), .Y(mai_mai_n214_));
  NO2        m192(.A(x06), .B(x00), .Y(mai_mai_n215_));
  NA2        m193(.A(mai_mai_n29_), .B(mai_mai_n48_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n216_), .B(x03), .Y(mai_mai_n217_));
  OA210      m195(.A0(mai_mai_n217_), .A1(mai_mai_n215_), .B0(mai_mai_n214_), .Y(mai_mai_n218_));
  NA2        m196(.A(x13), .B(mai_mai_n98_), .Y(mai_mai_n219_));
  NA3        m197(.A(mai_mai_n219_), .B(x12), .C(mai_mai_n89_), .Y(mai_mai_n220_));
  OAI210     m198(.A0(mai_mai_n218_), .A1(mai_mai_n213_), .B0(mai_mai_n220_), .Y(mai_mai_n221_));
  AOI210     m199(.A0(mai_mai_n212_), .A1(mai_mai_n210_), .B0(mai_mai_n221_), .Y(mai_mai_n222_));
  AOI210     m200(.A0(mai_mai_n222_), .A1(mai_mai_n199_), .B0(x07), .Y(mai_mai_n223_));
  NA2        m201(.A(mai_mai_n71_), .B(mai_mai_n29_), .Y(mai_mai_n224_));
  NOi31      m202(.An(mai_mai_n123_), .B(mai_mai_n206_), .C(mai_mai_n171_), .Y(mai_mai_n225_));
  AOI210     m203(.A0(mai_mai_n225_), .A1(x04), .B0(mai_mai_n224_), .Y(mai_mai_n226_));
  NO2        m204(.A(mai_mai_n99_), .B(x06), .Y(mai_mai_n227_));
  INV        m205(.A(mai_mai_n227_), .Y(mai_mai_n228_));
  NO2        m206(.A(x08), .B(x05), .Y(mai_mai_n229_));
  OAI210     m207(.A0(mai_mai_n75_), .A1(x13), .B0(mai_mai_n31_), .Y(mai_mai_n230_));
  OAI210     m208(.A0(mai_mai_n386_), .A1(mai_mai_n228_), .B0(mai_mai_n230_), .Y(mai_mai_n231_));
  NO2        m209(.A(x12), .B(x02), .Y(mai_mai_n232_));
  INV        m210(.A(mai_mai_n232_), .Y(mai_mai_n233_));
  NO2        m211(.A(mai_mai_n233_), .B(mai_mai_n211_), .Y(mai_mai_n234_));
  OA210      m212(.A0(mai_mai_n231_), .A1(mai_mai_n226_), .B0(mai_mai_n234_), .Y(mai_mai_n235_));
  NA2        m213(.A(mai_mai_n51_), .B(mai_mai_n41_), .Y(mai_mai_n236_));
  NO2        m214(.A(mai_mai_n236_), .B(x01), .Y(mai_mai_n237_));
  BUFFER     m215(.A(mai_mai_n81_), .Y(mai_mai_n238_));
  NO2        m216(.A(mai_mai_n238_), .B(mai_mai_n237_), .Y(mai_mai_n239_));
  AOI210     m217(.A0(mai_mai_n239_), .A1(mai_mai_n381_), .B0(mai_mai_n29_), .Y(mai_mai_n240_));
  NA2        m218(.A(mai_mai_n99_), .B(x04), .Y(mai_mai_n241_));
  OAI210     m219(.A0(x02), .A1(mai_mai_n111_), .B0(mai_mai_n382_), .Y(mai_mai_n242_));
  NO3        m220(.A(mai_mai_n87_), .B(x12), .C(x03), .Y(mai_mai_n243_));
  OAI210     m221(.A0(mai_mai_n242_), .A1(mai_mai_n240_), .B0(mai_mai_n243_), .Y(mai_mai_n244_));
  AOI210     m222(.A0(mai_mai_n178_), .A1(mai_mai_n174_), .B0(mai_mai_n100_), .Y(mai_mai_n245_));
  NOi21      m223(.An(mai_mai_n224_), .B(mai_mai_n385_), .Y(mai_mai_n246_));
  NO2        m224(.A(mai_mai_n25_), .B(x00), .Y(mai_mai_n247_));
  OAI210     m225(.A0(mai_mai_n246_), .A1(mai_mai_n245_), .B0(mai_mai_n247_), .Y(mai_mai_n248_));
  NO2        m226(.A(mai_mai_n58_), .B(x05), .Y(mai_mai_n249_));
  NO3        m227(.A(mai_mai_n249_), .B(mai_mai_n196_), .C(mai_mai_n166_), .Y(mai_mai_n250_));
  NO2        m228(.A(mai_mai_n213_), .B(mai_mai_n28_), .Y(mai_mai_n251_));
  OAI210     m229(.A0(mai_mai_n250_), .A1(mai_mai_n200_), .B0(mai_mai_n251_), .Y(mai_mai_n252_));
  NA3        m230(.A(mai_mai_n252_), .B(mai_mai_n248_), .C(mai_mai_n244_), .Y(mai_mai_n253_));
  NO3        m231(.A(mai_mai_n253_), .B(mai_mai_n235_), .C(mai_mai_n223_), .Y(mai_mai_n254_));
  OAI210     m232(.A0(mai_mai_n184_), .A1(mai_mai_n61_), .B0(mai_mai_n254_), .Y(mai02));
  AOI210     m233(.A0(mai_mai_n123_), .A1(mai_mai_n82_), .B0(mai_mai_n119_), .Y(mai_mai_n256_));
  NOi21      m234(.An(mai_mai_n207_), .B(mai_mai_n152_), .Y(mai_mai_n257_));
  NO2        m235(.A(mai_mai_n99_), .B(mai_mai_n35_), .Y(mai_mai_n258_));
  NA3        m236(.A(mai_mai_n258_), .B(x08), .C(mai_mai_n56_), .Y(mai_mai_n259_));
  OAI210     m237(.A0(mai_mai_n257_), .A1(mai_mai_n32_), .B0(mai_mai_n259_), .Y(mai_mai_n260_));
  OAI210     m238(.A0(mai_mai_n260_), .A1(mai_mai_n256_), .B0(mai_mai_n151_), .Y(mai_mai_n261_));
  INV        m239(.A(mai_mai_n151_), .Y(mai_mai_n262_));
  OAI210     m240(.A0(mai_mai_n82_), .A1(mai_mai_n51_), .B0(mai_mai_n99_), .Y(mai_mai_n263_));
  AOI220     m241(.A0(mai_mai_n263_), .A1(mai_mai_n262_), .B0(mai_mai_n134_), .B1(mai_mai_n133_), .Y(mai_mai_n264_));
  AOI210     m242(.A0(mai_mai_n264_), .A1(mai_mai_n261_), .B0(mai_mai_n48_), .Y(mai_mai_n265_));
  NO2        m243(.A(x05), .B(x02), .Y(mai_mai_n266_));
  OAI210     m244(.A0(mai_mai_n188_), .A1(mai_mai_n171_), .B0(mai_mai_n266_), .Y(mai_mai_n267_));
  AOI220     m245(.A0(mai_mai_n229_), .A1(mai_mai_n58_), .B0(mai_mai_n56_), .B1(mai_mai_n36_), .Y(mai_mai_n268_));
  NOi21      m246(.An(mai_mai_n258_), .B(mai_mai_n268_), .Y(mai_mai_n269_));
  AOI210     m247(.A0(mai_mai_n206_), .A1(mai_mai_n77_), .B0(mai_mai_n269_), .Y(mai_mai_n270_));
  AOI210     m248(.A0(mai_mai_n270_), .A1(mai_mai_n267_), .B0(mai_mai_n127_), .Y(mai_mai_n271_));
  NAi21      m249(.An(mai_mai_n208_), .B(mai_mai_n204_), .Y(mai_mai_n272_));
  NO2        m250(.A(mai_mai_n216_), .B(mai_mai_n47_), .Y(mai_mai_n273_));
  NA2        m251(.A(mai_mai_n273_), .B(mai_mai_n272_), .Y(mai_mai_n274_));
  AN2        m252(.A(mai_mai_n203_), .B(mai_mai_n202_), .Y(mai_mai_n275_));
  OAI210     m253(.A0(mai_mai_n42_), .A1(mai_mai_n41_), .B0(mai_mai_n48_), .Y(mai_mai_n276_));
  NA2        m254(.A(x13), .B(mai_mai_n28_), .Y(mai_mai_n277_));
  AOI210     m255(.A0(mai_mai_n277_), .A1(mai_mai_n124_), .B0(mai_mai_n276_), .Y(mai_mai_n278_));
  OAI210     m256(.A0(mai_mai_n278_), .A1(mai_mai_n275_), .B0(mai_mai_n93_), .Y(mai_mai_n279_));
  NA3        m257(.A(mai_mai_n93_), .B(mai_mai_n81_), .C(mai_mai_n201_), .Y(mai_mai_n280_));
  NA3        m258(.A(mai_mai_n92_), .B(mai_mai_n80_), .C(mai_mai_n42_), .Y(mai_mai_n281_));
  AOI210     m259(.A0(mai_mai_n281_), .A1(mai_mai_n280_), .B0(x04), .Y(mai_mai_n282_));
  NO2        m260(.A(mai_mai_n386_), .B(mai_mai_n101_), .Y(mai_mai_n283_));
  AOI210     m261(.A0(mai_mai_n283_), .A1(x13), .B0(mai_mai_n282_), .Y(mai_mai_n284_));
  NA3        m262(.A(mai_mai_n284_), .B(mai_mai_n279_), .C(mai_mai_n274_), .Y(mai_mai_n285_));
  NO3        m263(.A(mai_mai_n285_), .B(mai_mai_n271_), .C(mai_mai_n265_), .Y(mai_mai_n286_));
  NA2        m264(.A(mai_mai_n126_), .B(x03), .Y(mai_mai_n287_));
  INV        m265(.A(mai_mai_n160_), .Y(mai_mai_n288_));
  AOI210     m266(.A0(mai_mai_n179_), .A1(x08), .B0(mai_mai_n288_), .Y(mai_mai_n289_));
  OAI210     m267(.A0(mai_mai_n289_), .A1(mai_mai_n249_), .B0(mai_mai_n287_), .Y(mai_mai_n290_));
  NA2        m268(.A(mai_mai_n290_), .B(mai_mai_n102_), .Y(mai_mai_n291_));
  OAI210     m269(.A0(mai_mai_n56_), .A1(mai_mai_n153_), .B0(mai_mai_n103_), .Y(mai_mai_n292_));
  NA2        m270(.A(mai_mai_n241_), .B(mai_mai_n98_), .Y(mai_mai_n293_));
  NA2        m271(.A(mai_mai_n98_), .B(mai_mai_n41_), .Y(mai_mai_n294_));
  NA3        m272(.A(mai_mai_n294_), .B(mai_mai_n293_), .C(mai_mai_n118_), .Y(mai_mai_n295_));
  NA4        m273(.A(mai_mai_n295_), .B(mai_mai_n292_), .C(mai_mai_n291_), .D(mai_mai_n48_), .Y(mai_mai_n296_));
  INV        m274(.A(mai_mai_n179_), .Y(mai_mai_n297_));
  INV        m275(.A(x08), .Y(mai_mai_n298_));
  NA2        m276(.A(mai_mai_n176_), .B(x04), .Y(mai_mai_n299_));
  NO2        m277(.A(mai_mai_n299_), .B(mai_mai_n298_), .Y(mai_mai_n300_));
  NO3        m278(.A(mai_mai_n162_), .B(x13), .C(mai_mai_n31_), .Y(mai_mai_n301_));
  OAI210     m279(.A0(mai_mai_n301_), .A1(mai_mai_n300_), .B0(mai_mai_n93_), .Y(mai_mai_n302_));
  NO3        m280(.A(mai_mai_n176_), .B(mai_mai_n143_), .C(mai_mai_n52_), .Y(mai_mai_n303_));
  OAI210     m281(.A0(mai_mai_n131_), .A1(mai_mai_n36_), .B0(mai_mai_n98_), .Y(mai_mai_n304_));
  OAI210     m282(.A0(mai_mai_n304_), .A1(mai_mai_n172_), .B0(mai_mai_n303_), .Y(mai_mai_n305_));
  NA3        m283(.A(mai_mai_n305_), .B(mai_mai_n302_), .C(x06), .Y(mai_mai_n306_));
  NO2        m284(.A(mai_mai_n187_), .B(mai_mai_n64_), .Y(mai_mai_n307_));
  OAI220     m285(.A0(mai_mai_n144_), .A1(x09), .B0(x08), .B1(mai_mai_n41_), .Y(mai_mai_n308_));
  NO3        m286(.A(mai_mai_n249_), .B(mai_mai_n116_), .C(x08), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n308_), .A1(mai_mai_n200_), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  NO2        m288(.A(mai_mai_n48_), .B(mai_mai_n41_), .Y(mai_mai_n311_));
  NO3        m289(.A(mai_mai_n107_), .B(mai_mai_n117_), .C(mai_mai_n38_), .Y(mai_mai_n312_));
  AOI210     m290(.A0(mai_mai_n303_), .A1(mai_mai_n311_), .B0(mai_mai_n312_), .Y(mai_mai_n313_));
  OAI210     m291(.A0(mai_mai_n310_), .A1(mai_mai_n28_), .B0(mai_mai_n313_), .Y(mai_mai_n314_));
  AO220      m292(.A0(mai_mai_n314_), .A1(x04), .B0(mai_mai_n307_), .B1(x05), .Y(mai_mai_n315_));
  AOI210     m293(.A0(mai_mai_n306_), .A1(mai_mai_n296_), .B0(mai_mai_n315_), .Y(mai_mai_n316_));
  OAI210     m294(.A0(mai_mai_n286_), .A1(x12), .B0(mai_mai_n316_), .Y(mai03));
  OR2        m295(.A(mai_mai_n42_), .B(mai_mai_n201_), .Y(mai_mai_n318_));
  AOI210     m296(.A0(mai_mai_n134_), .A1(mai_mai_n98_), .B0(mai_mai_n318_), .Y(mai_mai_n319_));
  OAI210     m297(.A0(mai_mai_n384_), .A1(mai_mai_n319_), .B0(x05), .Y(mai_mai_n320_));
  NA2        m298(.A(mai_mai_n318_), .B(x05), .Y(mai_mai_n321_));
  AOI210     m299(.A0(mai_mai_n124_), .A1(mai_mai_n193_), .B0(mai_mai_n321_), .Y(mai_mai_n322_));
  AOI210     m300(.A0(mai_mai_n203_), .A1(x08), .B0(mai_mai_n113_), .Y(mai_mai_n323_));
  OAI220     m301(.A0(mai_mai_n323_), .A1(mai_mai_n59_), .B0(mai_mai_n277_), .B1(mai_mai_n268_), .Y(mai_mai_n324_));
  OAI210     m302(.A0(mai_mai_n324_), .A1(mai_mai_n322_), .B0(mai_mai_n98_), .Y(mai_mai_n325_));
  AOI210     m303(.A0(mai_mai_n130_), .A1(mai_mai_n60_), .B0(mai_mai_n38_), .Y(mai_mai_n326_));
  NO2        m304(.A(mai_mai_n152_), .B(mai_mai_n120_), .Y(mai_mai_n327_));
  OAI220     m305(.A0(mai_mai_n327_), .A1(mai_mai_n37_), .B0(mai_mai_n132_), .B1(x13), .Y(mai_mai_n328_));
  OAI210     m306(.A0(mai_mai_n328_), .A1(mai_mai_n326_), .B0(x04), .Y(mai_mai_n329_));
  NO3        m307(.A(mai_mai_n294_), .B(mai_mai_n82_), .C(mai_mai_n59_), .Y(mai_mai_n330_));
  AOI210     m308(.A0(mai_mai_n168_), .A1(mai_mai_n98_), .B0(mai_mai_n130_), .Y(mai_mai_n331_));
  OA210      m309(.A0(mai_mai_n145_), .A1(x12), .B0(mai_mai_n120_), .Y(mai_mai_n332_));
  NO3        m310(.A(mai_mai_n332_), .B(mai_mai_n331_), .C(mai_mai_n330_), .Y(mai_mai_n333_));
  NA4        m311(.A(mai_mai_n333_), .B(mai_mai_n329_), .C(mai_mai_n325_), .D(mai_mai_n320_), .Y(mai04));
  NO2        m312(.A(mai_mai_n85_), .B(mai_mai_n39_), .Y(mai_mai_n335_));
  XO2        m313(.A(mai_mai_n335_), .B(mai_mai_n219_), .Y(mai05));
  NA2        m314(.A(mai_mai_n71_), .B(mai_mai_n52_), .Y(mai_mai_n337_));
  AOI210     m315(.A0(mai_mai_n337_), .A1(mai_mai_n276_), .B0(mai_mai_n25_), .Y(mai_mai_n338_));
  NA3        m316(.A(mai_mai_n127_), .B(mai_mai_n119_), .C(mai_mai_n31_), .Y(mai_mai_n339_));
  AOI210     m317(.A0(mai_mai_n380_), .A1(mai_mai_n339_), .B0(mai_mai_n24_), .Y(mai_mai_n340_));
  OAI210     m318(.A0(mai_mai_n340_), .A1(mai_mai_n338_), .B0(mai_mai_n98_), .Y(mai_mai_n341_));
  NA2        m319(.A(x11), .B(mai_mai_n31_), .Y(mai_mai_n342_));
  NA2        m320(.A(mai_mai_n23_), .B(mai_mai_n28_), .Y(mai_mai_n343_));
  NA2        m321(.A(mai_mai_n224_), .B(x03), .Y(mai_mai_n344_));
  OAI220     m322(.A0(mai_mai_n344_), .A1(mai_mai_n343_), .B0(mai_mai_n342_), .B1(mai_mai_n78_), .Y(mai_mai_n345_));
  OAI210     m323(.A0(mai_mai_n26_), .A1(mai_mai_n98_), .B0(x07), .Y(mai_mai_n346_));
  AOI210     m324(.A0(mai_mai_n345_), .A1(x06), .B0(mai_mai_n346_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n33_), .B(mai_mai_n98_), .Y(mai_mai_n348_));
  AOI210     m326(.A0(mai_mai_n348_), .A1(mai_mai_n88_), .B0(x07), .Y(mai_mai_n349_));
  AOI210     m327(.A0(mai_mai_n347_), .A1(mai_mai_n341_), .B0(mai_mai_n349_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n129_), .B(mai_mai_n28_), .Y(mai_mai_n351_));
  NO2        m329(.A(mai_mai_n47_), .B(mai_mai_n351_), .Y(mai_mai_n352_));
  NA2        m330(.A(mai_mai_n352_), .B(mai_mai_n99_), .Y(mai_mai_n353_));
  AOI210     m331(.A0(mai_mai_n299_), .A1(mai_mai_n105_), .B0(mai_mai_n232_), .Y(mai_mai_n354_));
  NOi21      m332(.An(mai_mai_n287_), .B(mai_mai_n120_), .Y(mai_mai_n355_));
  OAI210     m333(.A0(x12), .A1(mai_mai_n47_), .B0(mai_mai_n35_), .Y(mai_mai_n356_));
  AOI210     m334(.A0(mai_mai_n219_), .A1(mai_mai_n47_), .B0(mai_mai_n356_), .Y(mai_mai_n357_));
  NO3        m335(.A(mai_mai_n357_), .B(mai_mai_n354_), .C(x08), .Y(mai_mai_n358_));
  NO2        m336(.A(mai_mai_n119_), .B(mai_mai_n28_), .Y(mai_mai_n359_));
  NO2        m337(.A(mai_mai_n359_), .B(mai_mai_n237_), .Y(mai_mai_n360_));
  NA3        m338(.A(mai_mai_n297_), .B(mai_mai_n114_), .C(x12), .Y(mai_mai_n361_));
  AO210      m339(.A0(mai_mai_n297_), .A1(mai_mai_n114_), .B0(mai_mai_n219_), .Y(mai_mai_n362_));
  NA3        m340(.A(mai_mai_n362_), .B(mai_mai_n361_), .C(x08), .Y(mai_mai_n363_));
  INV        m341(.A(mai_mai_n363_), .Y(mai_mai_n364_));
  AOI210     m342(.A0(mai_mai_n358_), .A1(mai_mai_n353_), .B0(mai_mai_n364_), .Y(mai_mai_n365_));
  INV        m343(.A(x03), .Y(mai_mai_n366_));
  NO2        m344(.A(mai_mai_n129_), .B(mai_mai_n43_), .Y(mai_mai_n367_));
  OAI210     m345(.A0(mai_mai_n367_), .A1(mai_mai_n366_), .B0(mai_mai_n167_), .Y(mai_mai_n368_));
  NA3        m346(.A(mai_mai_n360_), .B(mai_mai_n355_), .C(mai_mai_n293_), .Y(mai_mai_n369_));
  NA3        m347(.A(x14), .B(mai_mai_n369_), .C(mai_mai_n368_), .Y(mai_mai_n370_));
  AOI220     m348(.A0(mai_mai_n348_), .A1(mai_mai_n61_), .B0(mai_mai_n359_), .B1(mai_mai_n143_), .Y(mai_mai_n371_));
  NOi21      m349(.An(mai_mai_n241_), .B(mai_mai_n132_), .Y(mai_mai_n372_));
  NO2        m350(.A(mai_mai_n44_), .B(x04), .Y(mai_mai_n373_));
  OAI210     m351(.A0(mai_mai_n373_), .A1(mai_mai_n372_), .B0(mai_mai_n98_), .Y(mai_mai_n374_));
  OAI210     m352(.A0(mai_mai_n371_), .A1(mai_mai_n87_), .B0(mai_mai_n374_), .Y(mai_mai_n375_));
  NO4        m353(.A(mai_mai_n375_), .B(mai_mai_n370_), .C(mai_mai_n365_), .D(mai_mai_n350_), .Y(mai06));
  INV        m354(.A(x07), .Y(mai_mai_n379_));
  INV        m355(.A(mai_mai_n86_), .Y(mai_mai_n380_));
  INV        m356(.A(x13), .Y(mai_mai_n381_));
  INV        m357(.A(mai_mai_n227_), .Y(mai_mai_n382_));
  INV        m358(.A(mai_mai_n128_), .Y(mai_mai_n383_));
  INV        m359(.A(mai_mai_n299_), .Y(mai_mai_n384_));
  INV        m360(.A(x06), .Y(mai_mai_n385_));
  INV        m361(.A(x05), .Y(mai_mai_n386_));
  INV        m362(.A(x01), .Y(mai_mai_n387_));
  INV        u000(.A(x11), .Y(men_men_n23_));
  NA2        u001(.A(men_men_n23_), .B(x02), .Y(men_men_n24_));
  NA2        u002(.A(x11), .B(x03), .Y(men_men_n25_));
  NA2        u003(.A(men_men_n25_), .B(men_men_n24_), .Y(men_men_n26_));
  NA2        u004(.A(men_men_n26_), .B(x07), .Y(men_men_n27_));
  INV        u005(.A(x02), .Y(men_men_n28_));
  INV        u006(.A(x10), .Y(men_men_n29_));
  NA2        u007(.A(men_men_n29_), .B(men_men_n28_), .Y(men_men_n30_));
  INV        u008(.A(x03), .Y(men_men_n31_));
  NA2        u009(.A(x10), .B(men_men_n31_), .Y(men_men_n32_));
  NA3        u010(.A(men_men_n32_), .B(men_men_n30_), .C(x06), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n27_), .Y(men_men_n34_));
  INV        u012(.A(x04), .Y(men_men_n35_));
  INV        u013(.A(x08), .Y(men_men_n36_));
  NA2        u014(.A(men_men_n36_), .B(x02), .Y(men_men_n37_));
  NA2        u015(.A(x08), .B(x03), .Y(men_men_n38_));
  AOI210     u016(.A0(men_men_n38_), .A1(men_men_n37_), .B0(men_men_n35_), .Y(men_men_n39_));
  NA2        u017(.A(x09), .B(men_men_n31_), .Y(men_men_n40_));
  INV        u018(.A(x05), .Y(men_men_n41_));
  NO2        u019(.A(x09), .B(x02), .Y(men_men_n42_));
  NO2        u020(.A(men_men_n42_), .B(men_men_n41_), .Y(men_men_n43_));
  NA2        u021(.A(men_men_n43_), .B(men_men_n40_), .Y(men_men_n44_));
  INV        u022(.A(men_men_n44_), .Y(men_men_n45_));
  NO3        u023(.A(men_men_n45_), .B(men_men_n39_), .C(men_men_n34_), .Y(men00));
  INV        u024(.A(x01), .Y(men_men_n47_));
  INV        u025(.A(x06), .Y(men_men_n48_));
  NA2        u026(.A(men_men_n48_), .B(men_men_n28_), .Y(men_men_n49_));
  NO3        u027(.A(men_men_n49_), .B(x11), .C(x09), .Y(men_men_n50_));
  INV        u028(.A(x09), .Y(men_men_n51_));
  NO2        u029(.A(x10), .B(x02), .Y(men_men_n52_));
  NA2        u030(.A(men_men_n52_), .B(men_men_n51_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(x07), .Y(men_men_n54_));
  OAI210     u032(.A0(men_men_n54_), .A1(men_men_n50_), .B0(men_men_n47_), .Y(men_men_n55_));
  NOi21      u033(.An(x01), .B(x09), .Y(men_men_n56_));
  INV        u034(.A(x00), .Y(men_men_n57_));
  NO2        u035(.A(men_men_n51_), .B(men_men_n57_), .Y(men_men_n58_));
  NO2        u036(.A(men_men_n58_), .B(men_men_n56_), .Y(men_men_n59_));
  NA2        u037(.A(x09), .B(men_men_n57_), .Y(men_men_n60_));
  INV        u038(.A(x07), .Y(men_men_n61_));
  NA2        u039(.A(men_men_n61_), .B(men_men_n48_), .Y(men_men_n62_));
  AOI220     u040(.A0(men_men_n61_), .A1(men_men_n59_), .B0(men_men_n59_), .B1(men_men_n31_), .Y(men_men_n63_));
  AOI210     u041(.A0(men_men_n63_), .A1(men_men_n55_), .B0(x05), .Y(men_men_n64_));
  NA2        u042(.A(x10), .B(x09), .Y(men_men_n65_));
  NA2        u043(.A(x09), .B(x05), .Y(men_men_n66_));
  NA2        u044(.A(x10), .B(x06), .Y(men_men_n67_));
  NA3        u045(.A(men_men_n67_), .B(men_men_n66_), .C(men_men_n28_), .Y(men_men_n68_));
  NO2        u046(.A(men_men_n61_), .B(men_men_n41_), .Y(men_men_n69_));
  NA2        u047(.A(men_men_n68_), .B(x03), .Y(men_men_n70_));
  NOi31      u048(.An(x08), .B(x04), .C(x00), .Y(men_men_n71_));
  NO2        u049(.A(x09), .B(men_men_n41_), .Y(men_men_n72_));
  NO2        u050(.A(men_men_n72_), .B(men_men_n36_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n72_), .A1(men_men_n29_), .B0(x02), .Y(men_men_n74_));
  AOI210     u052(.A0(men_men_n73_), .A1(men_men_n48_), .B0(men_men_n74_), .Y(men_men_n75_));
  NO2        u053(.A(men_men_n36_), .B(x00), .Y(men_men_n76_));
  NO2        u054(.A(x08), .B(x01), .Y(men_men_n77_));
  OAI210     u055(.A0(men_men_n77_), .A1(men_men_n76_), .B0(men_men_n35_), .Y(men_men_n78_));
  NA2        u056(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n78_), .B(men_men_n75_), .Y(men_men_n80_));
  AN2        u058(.A(men_men_n80_), .B(men_men_n70_), .Y(men_men_n81_));
  INV        u059(.A(men_men_n78_), .Y(men_men_n82_));
  NO2        u060(.A(x06), .B(x05), .Y(men_men_n83_));
  NA2        u061(.A(x11), .B(x00), .Y(men_men_n84_));
  NO2        u062(.A(x11), .B(men_men_n47_), .Y(men_men_n85_));
  NOi21      u063(.An(men_men_n84_), .B(men_men_n85_), .Y(men_men_n86_));
  AOI210     u064(.A0(men_men_n83_), .A1(men_men_n82_), .B0(men_men_n86_), .Y(men_men_n87_));
  NO2        u065(.A(men_men_n53_), .B(x11), .Y(men_men_n88_));
  NOi21      u066(.An(x01), .B(x10), .Y(men_men_n89_));
  NO2        u067(.A(men_men_n29_), .B(men_men_n57_), .Y(men_men_n90_));
  NO3        u068(.A(men_men_n90_), .B(men_men_n89_), .C(x06), .Y(men_men_n91_));
  AOI220     u069(.A0(men_men_n91_), .A1(men_men_n27_), .B0(men_men_n88_), .B1(men_men_n82_), .Y(men_men_n92_));
  OAI210     u070(.A0(men_men_n87_), .A1(x07), .B0(men_men_n92_), .Y(men_men_n93_));
  NO3        u071(.A(men_men_n93_), .B(men_men_n81_), .C(men_men_n64_), .Y(men01));
  INV        u072(.A(x12), .Y(men_men_n95_));
  INV        u073(.A(x13), .Y(men_men_n96_));
  NA2        u074(.A(x08), .B(x04), .Y(men_men_n97_));
  NO2        u075(.A(men_men_n97_), .B(men_men_n57_), .Y(men_men_n98_));
  NA2        u076(.A(men_men_n98_), .B(men_men_n83_), .Y(men_men_n99_));
  NA2        u077(.A(men_men_n89_), .B(men_men_n28_), .Y(men_men_n100_));
  NO2        u078(.A(men_men_n100_), .B(men_men_n66_), .Y(men_men_n101_));
  NO2        u079(.A(x10), .B(x01), .Y(men_men_n102_));
  NO2        u080(.A(men_men_n29_), .B(x00), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n103_), .B(men_men_n102_), .Y(men_men_n104_));
  NA2        u082(.A(x04), .B(men_men_n28_), .Y(men_men_n105_));
  NO3        u083(.A(men_men_n105_), .B(men_men_n36_), .C(men_men_n41_), .Y(men_men_n106_));
  AOI210     u084(.A0(men_men_n106_), .A1(men_men_n104_), .B0(men_men_n101_), .Y(men_men_n107_));
  AOI210     u085(.A0(men_men_n107_), .A1(men_men_n99_), .B0(men_men_n96_), .Y(men_men_n108_));
  NO2        u086(.A(men_men_n56_), .B(x05), .Y(men_men_n109_));
  NOi21      u087(.An(men_men_n109_), .B(men_men_n58_), .Y(men_men_n110_));
  NO2        u088(.A(men_men_n35_), .B(x02), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n96_), .B(men_men_n36_), .Y(men_men_n112_));
  NA3        u090(.A(men_men_n112_), .B(men_men_n111_), .C(x06), .Y(men_men_n113_));
  NO2        u091(.A(men_men_n113_), .B(men_men_n110_), .Y(men_men_n114_));
  NO2        u092(.A(men_men_n77_), .B(x13), .Y(men_men_n115_));
  NA2        u093(.A(x09), .B(men_men_n35_), .Y(men_men_n116_));
  NO2        u094(.A(men_men_n116_), .B(men_men_n115_), .Y(men_men_n117_));
  NA2        u095(.A(x13), .B(men_men_n35_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n118_), .B(x05), .Y(men_men_n119_));
  NO2        u097(.A(men_men_n119_), .B(men_men_n117_), .Y(men_men_n120_));
  NA2        u098(.A(men_men_n35_), .B(men_men_n57_), .Y(men_men_n121_));
  NA2        u099(.A(men_men_n121_), .B(men_men_n96_), .Y(men_men_n122_));
  AOI210     u100(.A0(men_men_n122_), .A1(men_men_n73_), .B0(men_men_n110_), .Y(men_men_n123_));
  AOI210     u101(.A0(men_men_n123_), .A1(men_men_n120_), .B0(men_men_n67_), .Y(men_men_n124_));
  NA2        u102(.A(men_men_n29_), .B(men_men_n47_), .Y(men_men_n125_));
  NA2        u103(.A(x10), .B(men_men_n57_), .Y(men_men_n126_));
  NA2        u104(.A(men_men_n126_), .B(men_men_n125_), .Y(men_men_n127_));
  NA2        u105(.A(men_men_n51_), .B(x05), .Y(men_men_n128_));
  NA2        u106(.A(men_men_n36_), .B(x04), .Y(men_men_n129_));
  NA3        u107(.A(men_men_n129_), .B(men_men_n128_), .C(x13), .Y(men_men_n130_));
  NO3        u108(.A(men_men_n121_), .B(men_men_n72_), .C(men_men_n36_), .Y(men_men_n131_));
  NO2        u109(.A(men_men_n60_), .B(x05), .Y(men_men_n132_));
  NOi41      u110(.An(men_men_n130_), .B(men_men_n132_), .C(men_men_n131_), .D(men_men_n127_), .Y(men_men_n133_));
  NO3        u111(.A(men_men_n133_), .B(x06), .C(x03), .Y(men_men_n134_));
  NO4        u112(.A(men_men_n134_), .B(men_men_n124_), .C(men_men_n114_), .D(men_men_n108_), .Y(men_men_n135_));
  NA2        u113(.A(x13), .B(men_men_n36_), .Y(men_men_n136_));
  OAI210     u114(.A0(men_men_n77_), .A1(x13), .B0(men_men_n35_), .Y(men_men_n137_));
  NA2        u115(.A(men_men_n137_), .B(men_men_n136_), .Y(men_men_n138_));
  NO2        u116(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n139_));
  NA2        u117(.A(men_men_n29_), .B(x06), .Y(men_men_n140_));
  AOI210     u118(.A0(men_men_n140_), .A1(men_men_n49_), .B0(men_men_n139_), .Y(men_men_n141_));
  AN2        u119(.A(men_men_n141_), .B(men_men_n138_), .Y(men_men_n142_));
  NO2        u120(.A(x09), .B(x05), .Y(men_men_n143_));
  NA2        u121(.A(men_men_n143_), .B(men_men_n47_), .Y(men_men_n144_));
  AOI210     u122(.A0(men_men_n144_), .A1(men_men_n104_), .B0(men_men_n49_), .Y(men_men_n145_));
  NA2        u123(.A(x09), .B(x00), .Y(men_men_n146_));
  NA2        u124(.A(men_men_n109_), .B(men_men_n146_), .Y(men_men_n147_));
  NA2        u125(.A(men_men_n71_), .B(men_men_n51_), .Y(men_men_n148_));
  AOI210     u126(.A0(men_men_n148_), .A1(men_men_n147_), .B0(men_men_n140_), .Y(men_men_n149_));
  NO3        u127(.A(men_men_n149_), .B(men_men_n145_), .C(men_men_n142_), .Y(men_men_n150_));
  NO2        u128(.A(x03), .B(x02), .Y(men_men_n151_));
  NA2        u129(.A(men_men_n78_), .B(men_men_n96_), .Y(men_men_n152_));
  OAI210     u130(.A0(men_men_n152_), .A1(men_men_n110_), .B0(men_men_n151_), .Y(men_men_n153_));
  OA210      u131(.A0(men_men_n150_), .A1(x11), .B0(men_men_n153_), .Y(men_men_n154_));
  OAI210     u132(.A0(men_men_n135_), .A1(men_men_n23_), .B0(men_men_n154_), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n104_), .B(men_men_n40_), .Y(men_men_n156_));
  NA2        u134(.A(men_men_n23_), .B(men_men_n36_), .Y(men_men_n157_));
  NAi21      u135(.An(x06), .B(x10), .Y(men_men_n158_));
  NOi21      u136(.An(x01), .B(x13), .Y(men_men_n159_));
  NA2        u137(.A(men_men_n159_), .B(men_men_n158_), .Y(men_men_n160_));
  OR2        u138(.A(men_men_n160_), .B(men_men_n157_), .Y(men_men_n161_));
  AOI210     u139(.A0(men_men_n161_), .A1(men_men_n156_), .B0(men_men_n41_), .Y(men_men_n162_));
  NO2        u140(.A(men_men_n29_), .B(x03), .Y(men_men_n163_));
  NA2        u141(.A(men_men_n96_), .B(x01), .Y(men_men_n164_));
  NO2        u142(.A(men_men_n164_), .B(x08), .Y(men_men_n165_));
  OAI210     u143(.A0(x05), .A1(men_men_n165_), .B0(men_men_n51_), .Y(men_men_n166_));
  AOI210     u144(.A0(men_men_n166_), .A1(men_men_n163_), .B0(men_men_n48_), .Y(men_men_n167_));
  AOI210     u145(.A0(x11), .A1(men_men_n31_), .B0(men_men_n28_), .Y(men_men_n168_));
  OAI210     u146(.A0(men_men_n167_), .A1(men_men_n162_), .B0(men_men_n168_), .Y(men_men_n169_));
  NA2        u147(.A(x04), .B(x02), .Y(men_men_n170_));
  NA2        u148(.A(x10), .B(x05), .Y(men_men_n171_));
  NA2        u149(.A(x09), .B(x06), .Y(men_men_n172_));
  NO2        u150(.A(x09), .B(x01), .Y(men_men_n173_));
  NO3        u151(.A(men_men_n173_), .B(men_men_n102_), .C(men_men_n31_), .Y(men_men_n174_));
  NA2        u152(.A(men_men_n174_), .B(x00), .Y(men_men_n175_));
  NO2        u153(.A(men_men_n109_), .B(x08), .Y(men_men_n176_));
  NA3        u154(.A(men_men_n159_), .B(men_men_n158_), .C(men_men_n51_), .Y(men_men_n177_));
  NA2        u155(.A(men_men_n89_), .B(x05), .Y(men_men_n178_));
  OAI210     u156(.A0(men_men_n178_), .A1(men_men_n112_), .B0(men_men_n177_), .Y(men_men_n179_));
  AOI210     u157(.A0(men_men_n176_), .A1(x06), .B0(men_men_n179_), .Y(men_men_n180_));
  OAI210     u158(.A0(men_men_n180_), .A1(x11), .B0(men_men_n175_), .Y(men_men_n181_));
  NAi21      u159(.An(men_men_n170_), .B(men_men_n181_), .Y(men_men_n182_));
  INV        u160(.A(men_men_n25_), .Y(men_men_n183_));
  NAi21      u161(.An(x13), .B(x00), .Y(men_men_n184_));
  AOI210     u162(.A0(men_men_n29_), .A1(men_men_n48_), .B0(men_men_n184_), .Y(men_men_n185_));
  AOI220     u163(.A0(x09), .A1(x04), .B0(x08), .B1(x05), .Y(men_men_n186_));
  OAI210     u164(.A0(men_men_n171_), .A1(men_men_n35_), .B0(men_men_n186_), .Y(men_men_n187_));
  AN2        u165(.A(men_men_n187_), .B(men_men_n185_), .Y(men_men_n188_));
  AN2        u166(.A(men_men_n67_), .B(men_men_n66_), .Y(men_men_n189_));
  NO2        u167(.A(men_men_n90_), .B(x06), .Y(men_men_n190_));
  NO2        u168(.A(men_men_n184_), .B(men_men_n36_), .Y(men_men_n191_));
  OAI220     u169(.A0(men_men_n184_), .A1(men_men_n172_), .B0(men_men_n190_), .B1(men_men_n189_), .Y(men_men_n192_));
  OAI210     u170(.A0(men_men_n192_), .A1(men_men_n188_), .B0(men_men_n183_), .Y(men_men_n193_));
  NOi21      u171(.An(x09), .B(x00), .Y(men_men_n194_));
  NA2        u172(.A(x10), .B(x08), .Y(men_men_n195_));
  INV        u173(.A(men_men_n195_), .Y(men_men_n196_));
  NA2        u174(.A(x06), .B(x05), .Y(men_men_n197_));
  OAI210     u175(.A0(men_men_n197_), .A1(men_men_n35_), .B0(men_men_n95_), .Y(men_men_n198_));
  AOI210     u176(.A0(men_men_n196_), .A1(men_men_n58_), .B0(men_men_n198_), .Y(men_men_n199_));
  INV        u177(.A(men_men_n199_), .Y(men_men_n200_));
  NO2        u178(.A(men_men_n96_), .B(x12), .Y(men_men_n201_));
  AOI210     u179(.A0(men_men_n25_), .A1(men_men_n24_), .B0(men_men_n201_), .Y(men_men_n202_));
  NA2        u180(.A(men_men_n89_), .B(men_men_n51_), .Y(men_men_n203_));
  NO2        u181(.A(men_men_n35_), .B(men_men_n31_), .Y(men_men_n204_));
  NA2        u182(.A(men_men_n204_), .B(x02), .Y(men_men_n205_));
  NO2        u183(.A(men_men_n205_), .B(men_men_n203_), .Y(men_men_n206_));
  AOI210     u184(.A0(men_men_n202_), .A1(men_men_n200_), .B0(men_men_n206_), .Y(men_men_n207_));
  NA4        u185(.A(men_men_n207_), .B(men_men_n193_), .C(men_men_n182_), .D(men_men_n169_), .Y(men_men_n208_));
  AOI210     u186(.A0(men_men_n155_), .A1(men_men_n95_), .B0(men_men_n208_), .Y(men_men_n209_));
  NA2        u187(.A(men_men_n28_), .B(men_men_n138_), .Y(men_men_n210_));
  NA2        u188(.A(men_men_n51_), .B(men_men_n47_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n211_), .B(men_men_n137_), .Y(men_men_n212_));
  NO2        u190(.A(men_men_n125_), .B(x06), .Y(men_men_n213_));
  AOI210     u191(.A0(men_men_n451_), .A1(men_men_n212_), .B0(men_men_n213_), .Y(men_men_n214_));
  AOI210     u192(.A0(men_men_n214_), .A1(men_men_n210_), .B0(x12), .Y(men_men_n215_));
  INV        u193(.A(men_men_n71_), .Y(men_men_n216_));
  AOI210     u194(.A0(men_men_n195_), .A1(x05), .B0(men_men_n51_), .Y(men_men_n217_));
  OAI210     u195(.A0(men_men_n217_), .A1(men_men_n160_), .B0(men_men_n57_), .Y(men_men_n218_));
  NA2        u196(.A(men_men_n218_), .B(men_men_n216_), .Y(men_men_n219_));
  NO2        u197(.A(men_men_n89_), .B(x06), .Y(men_men_n220_));
  AOI210     u198(.A0(men_men_n36_), .A1(x04), .B0(men_men_n51_), .Y(men_men_n221_));
  NO3        u199(.A(men_men_n221_), .B(men_men_n220_), .C(men_men_n41_), .Y(men_men_n222_));
  NA4        u200(.A(men_men_n158_), .B(men_men_n56_), .C(men_men_n36_), .D(x04), .Y(men_men_n223_));
  NA2        u201(.A(men_men_n223_), .B(men_men_n140_), .Y(men_men_n224_));
  OAI210     u202(.A0(men_men_n224_), .A1(men_men_n222_), .B0(x02), .Y(men_men_n225_));
  AOI210     u203(.A0(men_men_n225_), .A1(men_men_n219_), .B0(men_men_n23_), .Y(men_men_n226_));
  OAI210     u204(.A0(men_men_n215_), .A1(men_men_n57_), .B0(men_men_n226_), .Y(men_men_n227_));
  INV        u205(.A(men_men_n140_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n51_), .B(x03), .Y(men_men_n229_));
  OAI210     u207(.A0(men_men_n72_), .A1(men_men_n36_), .B0(men_men_n116_), .Y(men_men_n230_));
  NO2        u208(.A(men_men_n96_), .B(x03), .Y(men_men_n231_));
  AOI220     u209(.A0(men_men_n231_), .A1(men_men_n230_), .B0(men_men_n71_), .B1(men_men_n229_), .Y(men_men_n232_));
  NA2        u210(.A(men_men_n32_), .B(x06), .Y(men_men_n233_));
  INV        u211(.A(men_men_n158_), .Y(men_men_n234_));
  NOi21      u212(.An(x13), .B(x04), .Y(men_men_n235_));
  NO3        u213(.A(men_men_n235_), .B(men_men_n71_), .C(men_men_n194_), .Y(men_men_n236_));
  NO2        u214(.A(men_men_n236_), .B(x05), .Y(men_men_n237_));
  AOI220     u215(.A0(men_men_n237_), .A1(men_men_n233_), .B0(men_men_n234_), .B1(men_men_n57_), .Y(men_men_n238_));
  OAI210     u216(.A0(men_men_n232_), .A1(men_men_n228_), .B0(men_men_n238_), .Y(men_men_n239_));
  INV        u217(.A(men_men_n85_), .Y(men_men_n240_));
  NO2        u218(.A(men_men_n240_), .B(x12), .Y(men_men_n241_));
  NA2        u219(.A(men_men_n23_), .B(men_men_n47_), .Y(men_men_n242_));
  NO2        u220(.A(men_men_n51_), .B(men_men_n36_), .Y(men_men_n243_));
  OAI210     u221(.A0(men_men_n243_), .A1(men_men_n187_), .B0(men_men_n185_), .Y(men_men_n244_));
  AOI210     u222(.A0(x08), .A1(x04), .B0(x09), .Y(men_men_n245_));
  NO2        u223(.A(x06), .B(x00), .Y(men_men_n246_));
  NO3        u224(.A(men_men_n246_), .B(men_men_n245_), .C(men_men_n41_), .Y(men_men_n247_));
  OAI210     u225(.A0(men_men_n97_), .A1(men_men_n146_), .B0(men_men_n67_), .Y(men_men_n248_));
  NO2        u226(.A(men_men_n248_), .B(men_men_n247_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n29_), .B(men_men_n48_), .Y(men_men_n250_));
  INV        u228(.A(x03), .Y(men_men_n251_));
  OA210      u229(.A0(men_men_n251_), .A1(men_men_n249_), .B0(men_men_n244_), .Y(men_men_n252_));
  NA2        u230(.A(x13), .B(men_men_n95_), .Y(men_men_n253_));
  NA3        u231(.A(men_men_n253_), .B(men_men_n198_), .C(men_men_n86_), .Y(men_men_n254_));
  OAI210     u232(.A0(men_men_n252_), .A1(men_men_n242_), .B0(men_men_n254_), .Y(men_men_n255_));
  AOI210     u233(.A0(men_men_n241_), .A1(men_men_n239_), .B0(men_men_n255_), .Y(men_men_n256_));
  AOI210     u234(.A0(men_men_n256_), .A1(men_men_n227_), .B0(x07), .Y(men_men_n257_));
  NA2        u235(.A(men_men_n66_), .B(men_men_n29_), .Y(men_men_n258_));
  NOi31      u236(.An(men_men_n136_), .B(men_men_n235_), .C(men_men_n194_), .Y(men_men_n259_));
  AOI210     u237(.A0(men_men_n259_), .A1(men_men_n148_), .B0(men_men_n258_), .Y(men_men_n260_));
  NO2        u238(.A(men_men_n96_), .B(x06), .Y(men_men_n261_));
  INV        u239(.A(men_men_n261_), .Y(men_men_n262_));
  NO2        u240(.A(x08), .B(x05), .Y(men_men_n263_));
  NO2        u241(.A(men_men_n263_), .B(men_men_n245_), .Y(men_men_n264_));
  OAI210     u242(.A0(men_men_n71_), .A1(x13), .B0(men_men_n31_), .Y(men_men_n265_));
  OAI210     u243(.A0(men_men_n264_), .A1(men_men_n262_), .B0(men_men_n265_), .Y(men_men_n266_));
  NO2        u244(.A(x12), .B(x02), .Y(men_men_n267_));
  INV        u245(.A(men_men_n267_), .Y(men_men_n268_));
  NO2        u246(.A(men_men_n268_), .B(men_men_n240_), .Y(men_men_n269_));
  OA210      u247(.A0(men_men_n266_), .A1(men_men_n260_), .B0(men_men_n269_), .Y(men_men_n270_));
  NA2        u248(.A(men_men_n51_), .B(men_men_n41_), .Y(men_men_n271_));
  NO2        u249(.A(men_men_n271_), .B(x01), .Y(men_men_n272_));
  NOi21      u250(.An(men_men_n77_), .B(men_men_n116_), .Y(men_men_n273_));
  NO2        u251(.A(men_men_n273_), .B(men_men_n272_), .Y(men_men_n274_));
  AOI210     u252(.A0(men_men_n274_), .A1(men_men_n130_), .B0(men_men_n29_), .Y(men_men_n275_));
  NA2        u253(.A(men_men_n261_), .B(men_men_n230_), .Y(men_men_n276_));
  NA2        u254(.A(men_men_n96_), .B(x04), .Y(men_men_n277_));
  NA2        u255(.A(men_men_n277_), .B(men_men_n28_), .Y(men_men_n278_));
  OAI210     u256(.A0(men_men_n278_), .A1(men_men_n115_), .B0(men_men_n276_), .Y(men_men_n279_));
  NO3        u257(.A(men_men_n84_), .B(x12), .C(x03), .Y(men_men_n280_));
  OAI210     u258(.A0(men_men_n279_), .A1(men_men_n275_), .B0(men_men_n280_), .Y(men_men_n281_));
  AOI210     u259(.A0(men_men_n203_), .A1(men_men_n197_), .B0(men_men_n97_), .Y(men_men_n282_));
  NOi21      u260(.An(men_men_n258_), .B(men_men_n220_), .Y(men_men_n283_));
  NO2        u261(.A(men_men_n25_), .B(x00), .Y(men_men_n284_));
  OAI210     u262(.A0(men_men_n283_), .A1(men_men_n282_), .B0(men_men_n284_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n58_), .B(x05), .Y(men_men_n286_));
  NO3        u264(.A(men_men_n286_), .B(men_men_n221_), .C(men_men_n190_), .Y(men_men_n287_));
  NO2        u265(.A(men_men_n242_), .B(men_men_n28_), .Y(men_men_n288_));
  OAI210     u266(.A0(men_men_n287_), .A1(men_men_n228_), .B0(men_men_n288_), .Y(men_men_n289_));
  NA3        u267(.A(men_men_n289_), .B(men_men_n285_), .C(men_men_n281_), .Y(men_men_n290_));
  NO3        u268(.A(men_men_n290_), .B(men_men_n270_), .C(men_men_n257_), .Y(men_men_n291_));
  OAI210     u269(.A0(men_men_n209_), .A1(men_men_n61_), .B0(men_men_n291_), .Y(men02));
  AOI210     u270(.A0(men_men_n136_), .A1(men_men_n78_), .B0(men_men_n128_), .Y(men_men_n293_));
  NA3        u271(.A(x13), .B(men_men_n196_), .C(men_men_n56_), .Y(men_men_n294_));
  OAI210     u272(.A0(men_men_n236_), .A1(men_men_n32_), .B0(men_men_n294_), .Y(men_men_n295_));
  OAI210     u273(.A0(men_men_n295_), .A1(men_men_n293_), .B0(men_men_n171_), .Y(men_men_n296_));
  INV        u274(.A(men_men_n171_), .Y(men_men_n297_));
  AOI210     u275(.A0(men_men_n111_), .A1(men_men_n79_), .B0(men_men_n221_), .Y(men_men_n298_));
  OAI220     u276(.A0(men_men_n298_), .A1(men_men_n96_), .B0(men_men_n78_), .B1(men_men_n51_), .Y(men_men_n299_));
  AOI220     u277(.A0(men_men_n299_), .A1(men_men_n297_), .B0(men_men_n152_), .B1(men_men_n151_), .Y(men_men_n300_));
  AOI210     u278(.A0(men_men_n300_), .A1(men_men_n296_), .B0(men_men_n48_), .Y(men_men_n301_));
  AOI220     u279(.A0(men_men_n263_), .A1(men_men_n58_), .B0(men_men_n56_), .B1(men_men_n36_), .Y(men_men_n302_));
  AOI210     u280(.A0(men_men_n235_), .A1(men_men_n72_), .B0(men_men_n263_), .Y(men_men_n303_));
  NO2        u281(.A(men_men_n303_), .B(men_men_n140_), .Y(men_men_n304_));
  NAi21      u282(.An(men_men_n237_), .B(men_men_n232_), .Y(men_men_n305_));
  NO2        u283(.A(men_men_n250_), .B(men_men_n47_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n306_), .B(men_men_n305_), .Y(men_men_n307_));
  AN2        u285(.A(men_men_n231_), .B(men_men_n230_), .Y(men_men_n308_));
  OAI210     u286(.A0(men_men_n42_), .A1(men_men_n41_), .B0(men_men_n48_), .Y(men_men_n309_));
  NA2        u287(.A(x13), .B(men_men_n28_), .Y(men_men_n310_));
  OA210      u288(.A0(men_men_n310_), .A1(x08), .B0(men_men_n144_), .Y(men_men_n311_));
  AOI210     u289(.A0(men_men_n311_), .A1(men_men_n137_), .B0(men_men_n309_), .Y(men_men_n312_));
  OAI210     u290(.A0(men_men_n312_), .A1(men_men_n308_), .B0(men_men_n90_), .Y(men_men_n313_));
  NA3        u291(.A(men_men_n90_), .B(men_men_n77_), .C(men_men_n229_), .Y(men_men_n314_));
  NA3        u292(.A(men_men_n89_), .B(men_men_n76_), .C(men_men_n42_), .Y(men_men_n315_));
  AOI210     u293(.A0(men_men_n315_), .A1(men_men_n314_), .B0(x04), .Y(men_men_n316_));
  INV        u294(.A(men_men_n151_), .Y(men_men_n317_));
  OAI220     u295(.A0(men_men_n264_), .A1(men_men_n100_), .B0(men_men_n317_), .B1(men_men_n127_), .Y(men_men_n318_));
  AOI210     u296(.A0(men_men_n318_), .A1(x13), .B0(men_men_n316_), .Y(men_men_n319_));
  NA3        u297(.A(men_men_n319_), .B(men_men_n313_), .C(men_men_n307_), .Y(men_men_n320_));
  NO3        u298(.A(men_men_n320_), .B(men_men_n304_), .C(men_men_n301_), .Y(men_men_n321_));
  NA2        u299(.A(men_men_n139_), .B(x03), .Y(men_men_n322_));
  INV        u300(.A(men_men_n184_), .Y(men_men_n323_));
  OAI210     u301(.A0(men_men_n51_), .A1(men_men_n35_), .B0(men_men_n36_), .Y(men_men_n324_));
  AOI220     u302(.A0(men_men_n324_), .A1(men_men_n323_), .B0(men_men_n204_), .B1(x08), .Y(men_men_n325_));
  OAI210     u303(.A0(men_men_n325_), .A1(men_men_n286_), .B0(men_men_n322_), .Y(men_men_n326_));
  NA2        u304(.A(men_men_n326_), .B(men_men_n102_), .Y(men_men_n327_));
  NA2        u305(.A(men_men_n170_), .B(men_men_n164_), .Y(men_men_n328_));
  AN2        u306(.A(men_men_n328_), .B(men_men_n176_), .Y(men_men_n329_));
  OAI220     u307(.A0(men_men_n277_), .A1(x09), .B0(men_men_n128_), .B1(men_men_n28_), .Y(men_men_n330_));
  OAI210     u308(.A0(men_men_n330_), .A1(men_men_n329_), .B0(men_men_n103_), .Y(men_men_n331_));
  NA2        u309(.A(men_men_n277_), .B(men_men_n95_), .Y(men_men_n332_));
  NA2        u310(.A(men_men_n95_), .B(men_men_n41_), .Y(men_men_n333_));
  NA3        u311(.A(men_men_n333_), .B(men_men_n332_), .C(men_men_n127_), .Y(men_men_n334_));
  NA4        u312(.A(men_men_n334_), .B(men_men_n331_), .C(men_men_n327_), .D(men_men_n48_), .Y(men_men_n335_));
  INV        u313(.A(men_men_n204_), .Y(men_men_n336_));
  NO2        u314(.A(men_men_n165_), .B(men_men_n40_), .Y(men_men_n337_));
  NA2        u315(.A(men_men_n32_), .B(x05), .Y(men_men_n338_));
  OAI220     u316(.A0(men_men_n338_), .A1(men_men_n337_), .B0(men_men_n336_), .B1(men_men_n59_), .Y(men_men_n339_));
  NA2        u317(.A(men_men_n339_), .B(x02), .Y(men_men_n340_));
  INV        u318(.A(men_men_n243_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n201_), .B(x04), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n342_), .B(men_men_n341_), .Y(men_men_n343_));
  NO3        u321(.A(men_men_n186_), .B(x13), .C(men_men_n31_), .Y(men_men_n344_));
  OAI210     u322(.A0(men_men_n344_), .A1(men_men_n343_), .B0(men_men_n90_), .Y(men_men_n345_));
  NO3        u323(.A(men_men_n201_), .B(men_men_n163_), .C(men_men_n52_), .Y(men_men_n346_));
  OAI210     u324(.A0(men_men_n146_), .A1(men_men_n36_), .B0(men_men_n95_), .Y(men_men_n347_));
  NA2        u325(.A(men_men_n347_), .B(men_men_n346_), .Y(men_men_n348_));
  NA4        u326(.A(men_men_n348_), .B(men_men_n345_), .C(men_men_n340_), .D(x06), .Y(men_men_n349_));
  NA2        u327(.A(x09), .B(x03), .Y(men_men_n350_));
  NO2        u328(.A(men_men_n350_), .B(men_men_n126_), .Y(men_men_n351_));
  NO3        u329(.A(men_men_n286_), .B(men_men_n125_), .C(x08), .Y(men_men_n352_));
  AOI210     u330(.A0(men_men_n96_), .A1(men_men_n228_), .B0(men_men_n352_), .Y(men_men_n353_));
  NO2        u331(.A(men_men_n48_), .B(men_men_n41_), .Y(men_men_n354_));
  NO3        u332(.A(men_men_n109_), .B(men_men_n126_), .C(men_men_n38_), .Y(men_men_n355_));
  AOI210     u333(.A0(men_men_n346_), .A1(men_men_n354_), .B0(men_men_n355_), .Y(men_men_n356_));
  OAI210     u334(.A0(men_men_n353_), .A1(men_men_n28_), .B0(men_men_n356_), .Y(men_men_n357_));
  AO220      u335(.A0(men_men_n357_), .A1(x04), .B0(men_men_n351_), .B1(x05), .Y(men_men_n358_));
  AOI210     u336(.A0(men_men_n349_), .A1(men_men_n335_), .B0(men_men_n358_), .Y(men_men_n359_));
  OAI210     u337(.A0(men_men_n321_), .A1(x12), .B0(men_men_n359_), .Y(men03));
  OR2        u338(.A(men_men_n42_), .B(men_men_n229_), .Y(men_men_n361_));
  AOI210     u339(.A0(men_men_n152_), .A1(men_men_n95_), .B0(men_men_n361_), .Y(men_men_n362_));
  AO210      u340(.A0(men_men_n341_), .A1(men_men_n79_), .B0(men_men_n342_), .Y(men_men_n363_));
  NA2        u341(.A(men_men_n201_), .B(men_men_n151_), .Y(men_men_n364_));
  NA3        u342(.A(men_men_n364_), .B(men_men_n363_), .C(men_men_n205_), .Y(men_men_n365_));
  OAI210     u343(.A0(men_men_n365_), .A1(men_men_n362_), .B0(x05), .Y(men_men_n366_));
  NA2        u344(.A(men_men_n361_), .B(x05), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n137_), .A1(men_men_n216_), .B0(men_men_n367_), .Y(men_men_n368_));
  AOI210     u346(.A0(men_men_n231_), .A1(men_men_n73_), .B0(men_men_n119_), .Y(men_men_n369_));
  OAI220     u347(.A0(men_men_n369_), .A1(men_men_n59_), .B0(men_men_n310_), .B1(men_men_n302_), .Y(men_men_n370_));
  OAI210     u348(.A0(men_men_n370_), .A1(men_men_n368_), .B0(men_men_n95_), .Y(men_men_n371_));
  NO2        u349(.A(men_men_n147_), .B(x13), .Y(men_men_n372_));
  NA2        u350(.A(men_men_n372_), .B(x04), .Y(men_men_n373_));
  AOI210     u351(.A0(men_men_n184_), .A1(men_men_n95_), .B0(men_men_n144_), .Y(men_men_n374_));
  OA210      u352(.A0(men_men_n165_), .A1(x12), .B0(men_men_n132_), .Y(men_men_n375_));
  NO2        u353(.A(men_men_n375_), .B(men_men_n374_), .Y(men_men_n376_));
  NA4        u354(.A(men_men_n376_), .B(men_men_n373_), .C(men_men_n371_), .D(men_men_n366_), .Y(men04));
  NO2        u355(.A(men_men_n82_), .B(men_men_n39_), .Y(men_men_n378_));
  XO2        u356(.A(men_men_n378_), .B(men_men_n253_), .Y(men05));
  AOI210     u357(.A0(men_men_n66_), .A1(men_men_n52_), .B0(men_men_n213_), .Y(men_men_n380_));
  AOI210     u358(.A0(men_men_n380_), .A1(men_men_n309_), .B0(men_men_n25_), .Y(men_men_n381_));
  NA3        u359(.A(men_men_n140_), .B(men_men_n128_), .C(men_men_n31_), .Y(men_men_n382_));
  AOI210     u360(.A0(men_men_n234_), .A1(men_men_n57_), .B0(men_men_n83_), .Y(men_men_n383_));
  AOI210     u361(.A0(men_men_n383_), .A1(men_men_n382_), .B0(men_men_n24_), .Y(men_men_n384_));
  OAI210     u362(.A0(men_men_n384_), .A1(men_men_n381_), .B0(men_men_n95_), .Y(men_men_n385_));
  NA2        u363(.A(x11), .B(men_men_n31_), .Y(men_men_n386_));
  NA2        u364(.A(men_men_n23_), .B(men_men_n28_), .Y(men_men_n387_));
  NA2        u365(.A(men_men_n258_), .B(x03), .Y(men_men_n388_));
  OAI220     u366(.A0(men_men_n388_), .A1(men_men_n387_), .B0(men_men_n386_), .B1(men_men_n74_), .Y(men_men_n389_));
  OAI210     u367(.A0(men_men_n26_), .A1(men_men_n95_), .B0(x07), .Y(men_men_n390_));
  AOI210     u368(.A0(men_men_n389_), .A1(x06), .B0(men_men_n390_), .Y(men_men_n391_));
  AOI220     u369(.A0(men_men_n74_), .A1(men_men_n31_), .B0(men_men_n52_), .B1(men_men_n51_), .Y(men_men_n392_));
  NO3        u370(.A(men_men_n392_), .B(men_men_n23_), .C(x00), .Y(men_men_n393_));
  NA2        u371(.A(men_men_n65_), .B(x02), .Y(men_men_n394_));
  AOI210     u372(.A0(men_men_n394_), .A1(men_men_n388_), .B0(men_men_n261_), .Y(men_men_n395_));
  OR2        u373(.A(men_men_n395_), .B(men_men_n242_), .Y(men_men_n396_));
  NA2        u374(.A(men_men_n159_), .B(x05), .Y(men_men_n397_));
  NA3        u375(.A(men_men_n397_), .B(men_men_n246_), .C(men_men_n240_), .Y(men_men_n398_));
  NO2        u376(.A(men_men_n23_), .B(x10), .Y(men_men_n399_));
  OAI210     u377(.A0(x11), .A1(men_men_n29_), .B0(men_men_n48_), .Y(men_men_n400_));
  OR3        u378(.A(men_men_n400_), .B(men_men_n399_), .C(men_men_n44_), .Y(men_men_n401_));
  NA3        u379(.A(men_men_n401_), .B(men_men_n398_), .C(men_men_n396_), .Y(men_men_n402_));
  OAI210     u380(.A0(men_men_n402_), .A1(men_men_n393_), .B0(men_men_n95_), .Y(men_men_n403_));
  AOI210     u381(.A0(x12), .A1(men_men_n85_), .B0(x07), .Y(men_men_n404_));
  AOI220     u382(.A0(men_men_n404_), .A1(men_men_n403_), .B0(men_men_n391_), .B1(men_men_n385_), .Y(men_men_n405_));
  NA3        u383(.A(men_men_n23_), .B(men_men_n61_), .C(men_men_n48_), .Y(men_men_n406_));
  AO210      u384(.A0(men_men_n406_), .A1(men_men_n271_), .B0(men_men_n268_), .Y(men_men_n407_));
  AOI210     u385(.A0(men_men_n399_), .A1(men_men_n69_), .B0(men_men_n139_), .Y(men_men_n408_));
  OR2        u386(.A(men_men_n408_), .B(x03), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n354_), .B(men_men_n61_), .Y(men_men_n410_));
  NO2        u388(.A(men_men_n410_), .B(x11), .Y(men_men_n411_));
  NO3        u389(.A(men_men_n411_), .B(men_men_n143_), .C(men_men_n28_), .Y(men_men_n412_));
  AOI220     u390(.A0(men_men_n412_), .A1(men_men_n409_), .B0(men_men_n407_), .B1(men_men_n47_), .Y(men_men_n413_));
  NO4        u391(.A(men_men_n333_), .B(men_men_n32_), .C(x11), .D(x09), .Y(men_men_n414_));
  OAI210     u392(.A0(men_men_n414_), .A1(men_men_n413_), .B0(men_men_n96_), .Y(men_men_n415_));
  AOI210     u393(.A0(men_men_n342_), .A1(men_men_n105_), .B0(men_men_n267_), .Y(men_men_n416_));
  NOi21      u394(.An(men_men_n322_), .B(men_men_n132_), .Y(men_men_n417_));
  NO2        u395(.A(men_men_n417_), .B(men_men_n268_), .Y(men_men_n418_));
  NO3        u396(.A(men_men_n418_), .B(men_men_n416_), .C(x08), .Y(men_men_n419_));
  AOI210     u397(.A0(men_men_n399_), .A1(men_men_n28_), .B0(men_men_n31_), .Y(men_men_n420_));
  NA2        u398(.A(x09), .B(men_men_n41_), .Y(men_men_n421_));
  OAI220     u399(.A0(men_men_n421_), .A1(men_men_n420_), .B0(men_men_n386_), .B1(men_men_n62_), .Y(men_men_n422_));
  NO2        u400(.A(x13), .B(x12), .Y(men_men_n423_));
  NO2        u401(.A(men_men_n128_), .B(men_men_n28_), .Y(men_men_n424_));
  NO2        u402(.A(men_men_n424_), .B(men_men_n272_), .Y(men_men_n425_));
  OR3        u403(.A(men_men_n425_), .B(x12), .C(x03), .Y(men_men_n426_));
  NA3        u404(.A(men_men_n336_), .B(men_men_n121_), .C(x12), .Y(men_men_n427_));
  AO210      u405(.A0(men_men_n336_), .A1(men_men_n121_), .B0(men_men_n253_), .Y(men_men_n428_));
  NA4        u406(.A(men_men_n428_), .B(men_men_n427_), .C(men_men_n426_), .D(x08), .Y(men_men_n429_));
  AOI210     u407(.A0(men_men_n423_), .A1(men_men_n422_), .B0(men_men_n429_), .Y(men_men_n430_));
  AOI210     u408(.A0(men_men_n419_), .A1(men_men_n415_), .B0(men_men_n430_), .Y(men_men_n431_));
  OAI210     u409(.A0(men_men_n410_), .A1(men_men_n23_), .B0(x03), .Y(men_men_n432_));
  NA2        u410(.A(men_men_n297_), .B(x07), .Y(men_men_n433_));
  OAI220     u411(.A0(men_men_n433_), .A1(men_men_n387_), .B0(men_men_n143_), .B1(men_men_n43_), .Y(men_men_n434_));
  OAI210     u412(.A0(men_men_n434_), .A1(men_men_n432_), .B0(men_men_n191_), .Y(men_men_n435_));
  NA3        u413(.A(men_men_n425_), .B(men_men_n417_), .C(men_men_n332_), .Y(men_men_n436_));
  INV        u414(.A(x14), .Y(men_men_n437_));
  NO3        u415(.A(men_men_n322_), .B(men_men_n100_), .C(x11), .Y(men_men_n438_));
  NO3        u416(.A(men_men_n164_), .B(men_men_n69_), .C(men_men_n57_), .Y(men_men_n439_));
  NO3        u417(.A(men_men_n406_), .B(men_men_n333_), .C(men_men_n184_), .Y(men_men_n440_));
  NO4        u418(.A(men_men_n440_), .B(men_men_n439_), .C(men_men_n438_), .D(men_men_n437_), .Y(men_men_n441_));
  NA3        u419(.A(men_men_n441_), .B(men_men_n436_), .C(men_men_n435_), .Y(men_men_n442_));
  NO3        u420(.A(men_men_n125_), .B(men_men_n24_), .C(x06), .Y(men_men_n443_));
  AOI210     u421(.A0(men_men_n284_), .A1(men_men_n234_), .B0(men_men_n443_), .Y(men_men_n444_));
  OAI210     u422(.A0(men_men_n44_), .A1(x04), .B0(men_men_n444_), .Y(men_men_n445_));
  NA2        u423(.A(men_men_n445_), .B(men_men_n95_), .Y(men_men_n446_));
  INV        u424(.A(men_men_n446_), .Y(men_men_n447_));
  NO4        u425(.A(men_men_n447_), .B(men_men_n442_), .C(men_men_n431_), .D(men_men_n405_), .Y(men06));
  INV        u426(.A(x05), .Y(men_men_n451_));
  VOTADOR g0(.A(ori00), .B(mai00), .C(men00), .Y(z0));
  VOTADOR g1(.A(ori01), .B(mai01), .C(men01), .Y(z1));
  VOTADOR g2(.A(ori02), .B(mai02), .C(men02), .Y(z2));
  VOTADOR g3(.A(ori03), .B(mai03), .C(men03), .Y(z3));
  VOTADOR g4(.A(ori04), .B(mai04), .C(men04), .Y(z4));
  VOTADOR g5(.A(ori05), .B(mai05), .C(men05), .Y(z5));
  VOTADOR g6(.A(ori06), .B(mai06), .C(men06), .Y(z6));
endmodule