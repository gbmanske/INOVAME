// Benchmark "top" written by ABC on Thu Jun 20 14:00:08 2024

module top ( 
    i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_,
    i_11_, i_2_, i_0_,
    ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4  );
  input  i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_,
    i_1_, i_11_, i_2_, i_0_;
  output ori1, ori2, ori0, ori7, ori5, ori6, ori3, ori4;
  wire new_new_n23_, new_new_n24_, new_new_n25_, new_new_n26_, new_new_n27_,
    new_new_n28_, new_new_n29_, new_new_n30_, new_new_n31_, new_new_n32_,
    new_new_n33_, new_new_n34_, new_new_n35_, new_new_n36_, new_new_n37_,
    new_new_n38_, new_new_n39_, new_new_n40_, new_new_n41_, new_new_n42_,
    new_new_n44_, new_new_n45_, new_new_n46_, new_new_n47_, new_new_n48_,
    new_new_n49_, new_new_n50_, new_new_n51_, new_new_n52_, new_new_n53_,
    new_new_n54_, new_new_n55_, new_new_n56_, new_new_n57_, new_new_n58_,
    new_new_n59_, new_new_n60_, new_new_n61_, new_new_n62_, new_new_n63_,
    new_new_n64_, new_new_n65_, new_new_n66_, new_new_n67_, new_new_n68_,
    new_new_n69_, new_new_n70_, new_new_n71_, new_new_n72_, new_new_n73_,
    new_new_n74_, new_new_n75_, new_new_n76_, new_new_n77_, new_new_n78_,
    new_new_n79_, new_new_n80_, new_new_n81_, new_new_n82_, new_new_n83_,
    new_new_n84_, new_new_n85_, new_new_n86_, new_new_n87_, new_new_n88_,
    new_new_n89_, new_new_n90_, new_new_n91_, new_new_n92_, new_new_n93_,
    new_new_n94_, new_new_n95_, new_new_n96_, new_new_n97_, new_new_n98_,
    new_new_n99_, new_new_n100_, new_new_n101_, new_new_n102_,
    new_new_n103_, new_new_n104_, new_new_n105_, new_new_n106_,
    new_new_n107_, new_new_n108_, new_new_n109_, new_new_n110_,
    new_new_n111_, new_new_n112_, new_new_n113_, new_new_n114_,
    new_new_n115_, new_new_n116_, new_new_n117_, new_new_n118_,
    new_new_n119_, new_new_n120_, new_new_n121_, new_new_n122_,
    new_new_n123_, new_new_n124_, new_new_n125_, new_new_n126_,
    new_new_n127_, new_new_n128_, new_new_n129_, new_new_n130_,
    new_new_n131_, new_new_n132_, new_new_n133_, new_new_n134_,
    new_new_n135_, new_new_n136_, new_new_n137_, new_new_n138_,
    new_new_n139_, new_new_n140_, new_new_n142_, new_new_n143_,
    new_new_n144_, new_new_n146_, new_new_n147_, new_new_n148_,
    new_new_n149_, new_new_n150_, new_new_n151_, new_new_n152_,
    new_new_n153_, new_new_n154_, new_new_n155_, new_new_n156_,
    new_new_n157_, new_new_n158_, new_new_n159_, new_new_n160_,
    new_new_n161_, new_new_n162_, new_new_n163_, new_new_n164_,
    new_new_n165_, new_new_n166_, new_new_n167_, new_new_n168_,
    new_new_n169_, new_new_n170_, new_new_n171_, new_new_n172_,
    new_new_n173_, new_new_n174_, new_new_n175_, new_new_n176_,
    new_new_n177_, new_new_n178_, new_new_n179_, new_new_n180_,
    new_new_n181_, new_new_n182_, new_new_n183_, new_new_n184_,
    new_new_n185_, new_new_n186_, new_new_n187_, new_new_n188_,
    new_new_n189_, new_new_n190_, new_new_n191_, new_new_n192_,
    new_new_n193_, new_new_n194_, new_new_n195_, new_new_n196_,
    new_new_n197_, new_new_n198_, new_new_n199_, new_new_n200_,
    new_new_n201_, new_new_n202_, new_new_n203_, new_new_n204_,
    new_new_n205_, new_new_n206_, new_new_n207_, new_new_n208_,
    new_new_n209_, new_new_n210_, new_new_n211_, new_new_n212_,
    new_new_n213_, new_new_n214_, new_new_n215_, new_new_n216_,
    new_new_n217_, new_new_n218_, new_new_n219_, new_new_n220_,
    new_new_n221_, new_new_n222_, new_new_n223_, new_new_n224_,
    new_new_n225_, new_new_n226_, new_new_n227_, new_new_n228_,
    new_new_n229_, new_new_n230_, new_new_n231_, new_new_n232_,
    new_new_n233_, new_new_n234_, new_new_n235_, new_new_n236_,
    new_new_n237_, new_new_n238_, new_new_n239_, new_new_n240_,
    new_new_n241_, new_new_n242_, new_new_n243_, new_new_n244_,
    new_new_n245_, new_new_n246_, new_new_n247_, new_new_n248_,
    new_new_n249_, new_new_n250_, new_new_n251_, new_new_n252_,
    new_new_n253_, new_new_n254_, new_new_n255_, new_new_n256_,
    new_new_n257_, new_new_n258_, new_new_n259_, new_new_n260_,
    new_new_n261_, new_new_n262_, new_new_n263_, new_new_n264_,
    new_new_n265_, new_new_n266_, new_new_n267_, new_new_n268_,
    new_new_n269_, new_new_n270_, new_new_n271_, new_new_n272_,
    new_new_n273_, new_new_n274_, new_new_n275_, new_new_n276_,
    new_new_n277_, new_new_n278_, new_new_n279_, new_new_n280_,
    new_new_n281_, new_new_n282_, new_new_n283_, new_new_n284_,
    new_new_n285_, new_new_n286_, new_new_n287_, new_new_n288_,
    new_new_n289_, new_new_n290_, new_new_n291_, new_new_n292_,
    new_new_n293_, new_new_n294_, new_new_n295_, new_new_n296_,
    new_new_n297_, new_new_n298_, new_new_n299_, new_new_n300_,
    new_new_n301_, new_new_n302_, new_new_n303_, new_new_n304_,
    new_new_n305_, new_new_n306_, new_new_n307_, new_new_n308_,
    new_new_n309_, new_new_n310_, new_new_n311_, new_new_n312_,
    new_new_n313_, new_new_n314_, new_new_n315_, new_new_n316_,
    new_new_n317_, new_new_n318_, new_new_n319_, new_new_n320_,
    new_new_n321_, new_new_n322_, new_new_n323_, new_new_n324_,
    new_new_n325_, new_new_n326_, new_new_n327_, new_new_n328_,
    new_new_n329_, new_new_n330_, new_new_n331_, new_new_n332_,
    new_new_n333_, new_new_n334_, new_new_n335_, new_new_n336_,
    new_new_n337_, new_new_n338_, new_new_n339_, new_new_n340_,
    new_new_n341_, new_new_n342_, new_new_n343_, new_new_n344_,
    new_new_n345_, new_new_n346_, new_new_n347_, new_new_n348_,
    new_new_n349_, new_new_n350_, new_new_n351_, new_new_n352_,
    new_new_n353_, new_new_n354_, new_new_n355_, new_new_n356_,
    new_new_n357_, new_new_n358_, new_new_n359_, new_new_n360_,
    new_new_n361_, new_new_n362_, new_new_n363_, new_new_n364_,
    new_new_n365_, new_new_n366_, new_new_n367_, new_new_n368_,
    new_new_n369_, new_new_n370_, new_new_n371_, new_new_n372_,
    new_new_n373_, new_new_n374_, new_new_n375_, new_new_n376_,
    new_new_n377_, new_new_n378_, new_new_n379_, new_new_n380_,
    new_new_n381_, new_new_n382_, new_new_n383_, new_new_n384_,
    new_new_n385_, new_new_n386_, new_new_n387_, new_new_n388_,
    new_new_n389_, new_new_n390_, new_new_n391_, new_new_n392_,
    new_new_n393_, new_new_n394_, new_new_n395_, new_new_n396_,
    new_new_n397_, new_new_n398_, new_new_n399_, new_new_n400_,
    new_new_n401_, new_new_n402_, new_new_n403_, new_new_n404_,
    new_new_n405_, new_new_n406_, new_new_n407_, new_new_n408_,
    new_new_n409_, new_new_n410_, new_new_n411_, new_new_n412_,
    new_new_n413_, new_new_n414_, new_new_n415_, new_new_n416_,
    new_new_n417_, new_new_n418_, new_new_n419_, new_new_n420_,
    new_new_n421_, new_new_n422_, new_new_n423_, new_new_n424_,
    new_new_n425_, new_new_n426_, new_new_n427_, new_new_n428_,
    new_new_n429_, new_new_n430_, new_new_n431_, new_new_n432_,
    new_new_n433_, new_new_n434_, new_new_n435_, new_new_n436_,
    new_new_n437_, new_new_n438_, new_new_n439_, new_new_n440_,
    new_new_n441_, new_new_n442_, new_new_n443_, new_new_n444_,
    new_new_n445_, new_new_n446_, new_new_n447_, new_new_n448_,
    new_new_n449_, new_new_n450_, new_new_n451_, new_new_n452_,
    new_new_n453_, new_new_n454_, new_new_n455_, new_new_n456_,
    new_new_n457_, new_new_n458_, new_new_n459_, new_new_n460_,
    new_new_n461_, new_new_n462_, new_new_n463_, new_new_n464_,
    new_new_n465_, new_new_n466_, new_new_n467_, new_new_n469_,
    new_new_n470_, new_new_n471_, new_new_n472_, new_new_n473_,
    new_new_n474_, new_new_n475_, new_new_n476_, new_new_n477_,
    new_new_n478_, new_new_n479_, new_new_n480_, new_new_n481_,
    new_new_n482_, new_new_n483_, new_new_n484_, new_new_n485_,
    new_new_n486_, new_new_n487_, new_new_n488_, new_new_n489_,
    new_new_n490_, new_new_n491_, new_new_n492_, new_new_n493_,
    new_new_n494_, new_new_n495_, new_new_n496_, new_new_n497_,
    new_new_n498_, new_new_n499_, new_new_n500_, new_new_n501_,
    new_new_n502_, new_new_n503_, new_new_n504_, new_new_n505_,
    new_new_n506_, new_new_n507_, new_new_n508_, new_new_n509_,
    new_new_n510_, new_new_n511_, new_new_n512_, new_new_n513_,
    new_new_n514_, new_new_n515_, new_new_n516_, new_new_n517_,
    new_new_n518_, new_new_n519_, new_new_n520_, new_new_n521_,
    new_new_n522_, new_new_n523_, new_new_n524_, new_new_n525_,
    new_new_n526_, new_new_n527_, new_new_n528_, new_new_n529_,
    new_new_n530_, new_new_n531_, new_new_n532_, new_new_n533_,
    new_new_n534_, new_new_n535_, new_new_n536_, new_new_n537_,
    new_new_n538_, new_new_n539_, new_new_n540_, new_new_n541_,
    new_new_n542_, new_new_n543_, new_new_n544_, new_new_n545_,
    new_new_n546_, new_new_n547_, new_new_n548_, new_new_n549_,
    new_new_n550_, new_new_n551_, new_new_n552_, new_new_n553_,
    new_new_n554_, new_new_n555_, new_new_n556_, new_new_n557_,
    new_new_n558_, new_new_n559_, new_new_n560_, new_new_n561_,
    new_new_n562_, new_new_n563_, new_new_n564_, new_new_n565_,
    new_new_n566_, new_new_n567_, new_new_n568_, new_new_n569_,
    new_new_n570_, new_new_n571_, new_new_n572_, new_new_n573_,
    new_new_n574_, new_new_n575_, new_new_n576_, new_new_n577_,
    new_new_n578_, new_new_n579_, new_new_n580_, new_new_n581_,
    new_new_n582_, new_new_n583_, new_new_n584_, new_new_n585_,
    new_new_n586_, new_new_n587_, new_new_n588_, new_new_n589_,
    new_new_n590_, new_new_n591_, new_new_n592_, new_new_n593_,
    new_new_n594_, new_new_n595_, new_new_n596_, new_new_n597_,
    new_new_n598_, new_new_n599_, new_new_n600_, new_new_n601_,
    new_new_n602_, new_new_n603_, new_new_n604_, new_new_n605_,
    new_new_n606_, new_new_n607_, new_new_n608_, new_new_n609_,
    new_new_n610_, new_new_n611_, new_new_n612_, new_new_n613_,
    new_new_n614_, new_new_n615_, new_new_n616_, new_new_n617_,
    new_new_n618_, new_new_n619_, new_new_n620_, new_new_n621_,
    new_new_n622_, new_new_n623_, new_new_n624_, new_new_n626_,
    new_new_n627_, new_new_n628_, new_new_n629_, new_new_n630_,
    new_new_n631_, new_new_n632_, new_new_n633_, new_new_n634_,
    new_new_n635_, new_new_n636_, new_new_n637_, new_new_n638_,
    new_new_n639_, new_new_n640_, new_new_n641_, new_new_n642_,
    new_new_n643_, new_new_n644_, new_new_n645_, new_new_n646_,
    new_new_n647_, new_new_n648_, new_new_n649_, new_new_n650_,
    new_new_n651_, new_new_n652_, new_new_n653_, new_new_n654_,
    new_new_n655_, new_new_n656_, new_new_n657_, new_new_n658_,
    new_new_n659_, new_new_n660_, new_new_n661_, new_new_n662_,
    new_new_n663_, new_new_n664_, new_new_n665_, new_new_n666_,
    new_new_n667_, new_new_n668_, new_new_n669_, new_new_n670_,
    new_new_n671_, new_new_n672_, new_new_n673_, new_new_n675_,
    new_new_n676_, new_new_n677_, new_new_n678_, new_new_n679_,
    new_new_n680_, new_new_n681_, new_new_n682_, new_new_n683_,
    new_new_n684_, new_new_n685_, new_new_n686_, new_new_n687_,
    new_new_n688_, new_new_n689_, new_new_n690_, new_new_n691_,
    new_new_n692_, new_new_n693_, new_new_n694_, new_new_n695_,
    new_new_n696_, new_new_n697_, new_new_n698_, new_new_n699_,
    new_new_n700_, new_new_n701_, new_new_n702_, new_new_n703_,
    new_new_n704_, new_new_n705_, new_new_n706_, new_new_n707_,
    new_new_n708_, new_new_n709_, new_new_n710_, new_new_n711_,
    new_new_n712_, new_new_n713_, new_new_n714_, new_new_n715_,
    new_new_n716_, new_new_n717_, new_new_n718_, new_new_n719_,
    new_new_n720_, new_new_n721_, new_new_n723_, new_new_n724_,
    new_new_n725_, new_new_n726_, new_new_n727_, new_new_n728_,
    new_new_n729_, new_new_n730_, new_new_n731_, new_new_n732_,
    new_new_n733_, new_new_n734_, new_new_n735_, new_new_n736_,
    new_new_n737_, new_new_n738_, new_new_n739_, new_new_n740_,
    new_new_n741_, new_new_n742_, new_new_n743_, new_new_n744_,
    new_new_n745_, new_new_n746_, new_new_n747_, new_new_n748_,
    new_new_n749_, new_new_n750_, new_new_n751_, new_new_n752_,
    new_new_n753_, new_new_n754_, new_new_n755_, new_new_n756_,
    new_new_n757_, new_new_n758_, new_new_n759_, new_new_n760_,
    new_new_n761_, new_new_n762_, new_new_n763_, new_new_n764_,
    new_new_n765_, new_new_n766_, new_new_n767_, new_new_n768_,
    new_new_n769_, new_new_n770_, new_new_n771_, new_new_n772_,
    new_new_n773_, new_new_n774_, new_new_n775_, new_new_n776_,
    new_new_n777_, new_new_n778_, new_new_n779_, new_new_n780_,
    new_new_n781_, new_new_n782_, new_new_n783_, new_new_n784_,
    new_new_n785_, new_new_n786_, new_new_n787_, new_new_n788_,
    new_new_n789_, new_new_n790_, new_new_n791_, new_new_n792_,
    new_new_n793_, new_new_n794_, new_new_n795_, new_new_n796_,
    new_new_n797_, new_new_n798_, new_new_n799_, new_new_n800_,
    new_new_n801_, new_new_n802_, new_new_n803_, new_new_n804_,
    new_new_n805_, new_new_n806_, new_new_n807_, new_new_n808_,
    new_new_n809_, new_new_n810_, new_new_n811_, new_new_n812_,
    new_new_n813_, new_new_n814_, new_new_n815_, new_new_n816_,
    new_new_n817_, new_new_n818_, new_new_n819_, new_new_n820_,
    new_new_n821_, new_new_n822_, new_new_n823_, new_new_n824_,
    new_new_n825_, new_new_n826_, new_new_n827_, new_new_n828_,
    new_new_n829_, new_new_n830_, new_new_n831_, new_new_n832_,
    new_new_n833_, new_new_n834_, new_new_n835_, new_new_n836_,
    new_new_n837_, new_new_n838_, new_new_n839_, new_new_n840_,
    new_new_n841_, new_new_n842_, new_new_n843_, new_new_n844_,
    new_new_n845_, new_new_n846_, new_new_n847_, new_new_n848_,
    new_new_n849_, new_new_n850_, new_new_n851_, new_new_n852_,
    new_new_n853_, new_new_n854_, new_new_n855_, new_new_n856_,
    new_new_n857_, new_new_n858_, new_new_n859_, new_new_n860_,
    new_new_n861_, new_new_n862_, new_new_n863_, new_new_n864_,
    new_new_n865_, new_new_n866_, new_new_n867_, new_new_n868_,
    new_new_n869_, new_new_n870_, new_new_n871_, new_new_n872_,
    new_new_n873_, new_new_n874_, new_new_n875_, new_new_n876_,
    new_new_n877_, new_new_n878_, new_new_n879_, new_new_n880_,
    new_new_n881_, new_new_n882_, new_new_n883_, new_new_n884_,
    new_new_n885_, new_new_n886_, new_new_n887_, new_new_n888_,
    new_new_n889_, new_new_n893_;
  NAi21      g000(.An(i_13_), .B(i_4_), .Y(new_new_n23_));
  NOi21      g001(.An(i_3_), .B(i_8_), .Y(new_new_n24_));
  INV        g002(.A(i_9_), .Y(new_new_n25_));
  INV        g003(.A(i_3_), .Y(new_new_n26_));
  NO2        g004(.A(new_new_n26_), .B(new_new_n25_), .Y(new_new_n27_));
  NO2        g005(.A(i_8_), .B(i_10_), .Y(new_new_n28_));
  INV        g006(.A(new_new_n28_), .Y(new_new_n29_));
  OAI210     g007(.A0(new_new_n27_), .A1(new_new_n24_), .B0(new_new_n29_), .Y(new_new_n30_));
  NOi21      g008(.An(i_11_), .B(i_8_), .Y(new_new_n31_));
  AO210      g009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(new_new_n32_));
  OR2        g010(.A(new_new_n32_), .B(new_new_n31_), .Y(new_new_n33_));
  NA2        g011(.A(new_new_n33_), .B(new_new_n30_), .Y(new_new_n34_));
  XO2        g012(.A(new_new_n34_), .B(new_new_n23_), .Y(new_new_n35_));
  INV        g013(.A(i_4_), .Y(new_new_n36_));
  INV        g014(.A(i_10_), .Y(new_new_n37_));
  NAi21      g015(.An(i_11_), .B(i_9_), .Y(new_new_n38_));
  NO3        g016(.A(new_new_n38_), .B(i_12_), .C(new_new_n37_), .Y(new_new_n39_));
  NOi21      g017(.An(i_12_), .B(i_13_), .Y(new_new_n40_));
  INV        g018(.A(new_new_n40_), .Y(new_new_n41_));
  NAi31      g019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(new_new_n42_));
  INV        g020(.A(new_new_n35_), .Y(ori1));
  INV        g021(.A(i_11_), .Y(new_new_n44_));
  NO2        g022(.A(new_new_n44_), .B(i_6_), .Y(new_new_n45_));
  INV        g023(.A(i_2_), .Y(new_new_n46_));
  NA2        g024(.A(i_0_), .B(i_3_), .Y(new_new_n47_));
  INV        g025(.A(i_5_), .Y(new_new_n48_));
  NO2        g026(.A(i_7_), .B(i_10_), .Y(new_new_n49_));
  AOI210     g027(.A0(i_7_), .A1(new_new_n25_), .B0(new_new_n49_), .Y(new_new_n50_));
  OAI210     g028(.A0(new_new_n50_), .A1(i_3_), .B0(new_new_n48_), .Y(new_new_n51_));
  AOI210     g029(.A0(new_new_n51_), .A1(new_new_n47_), .B0(new_new_n46_), .Y(new_new_n52_));
  NA2        g030(.A(i_0_), .B(i_2_), .Y(new_new_n53_));
  NA2        g031(.A(i_7_), .B(i_9_), .Y(new_new_n54_));
  NO2        g032(.A(new_new_n54_), .B(new_new_n53_), .Y(new_new_n55_));
  NA2        g033(.A(new_new_n52_), .B(new_new_n45_), .Y(new_new_n56_));
  NA3        g034(.A(i_2_), .B(i_6_), .C(i_8_), .Y(new_new_n57_));
  NO2        g035(.A(i_1_), .B(i_6_), .Y(new_new_n58_));
  NA2        g036(.A(i_8_), .B(i_7_), .Y(new_new_n59_));
  OAI210     g037(.A0(new_new_n59_), .A1(new_new_n58_), .B0(new_new_n57_), .Y(new_new_n60_));
  NA2        g038(.A(new_new_n60_), .B(i_12_), .Y(new_new_n61_));
  NAi21      g039(.An(i_2_), .B(i_7_), .Y(new_new_n62_));
  INV        g040(.A(i_1_), .Y(new_new_n63_));
  NA2        g041(.A(new_new_n63_), .B(i_6_), .Y(new_new_n64_));
  NA3        g042(.A(new_new_n64_), .B(new_new_n62_), .C(new_new_n31_), .Y(new_new_n65_));
  NA2        g043(.A(i_1_), .B(i_10_), .Y(new_new_n66_));
  NO2        g044(.A(new_new_n66_), .B(i_6_), .Y(new_new_n67_));
  NAi31      g045(.An(new_new_n67_), .B(new_new_n65_), .C(new_new_n61_), .Y(new_new_n68_));
  NA2        g046(.A(new_new_n50_), .B(i_2_), .Y(new_new_n69_));
  AOI210     g047(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(new_new_n70_));
  NA2        g048(.A(i_1_), .B(i_6_), .Y(new_new_n71_));
  NO2        g049(.A(new_new_n71_), .B(new_new_n25_), .Y(new_new_n72_));
  INV        g050(.A(i_0_), .Y(new_new_n73_));
  NAi21      g051(.An(i_5_), .B(i_10_), .Y(new_new_n74_));
  NA2        g052(.A(i_5_), .B(i_9_), .Y(new_new_n75_));
  AOI210     g053(.A0(new_new_n75_), .A1(new_new_n74_), .B0(new_new_n73_), .Y(new_new_n76_));
  NO2        g054(.A(new_new_n76_), .B(new_new_n72_), .Y(new_new_n77_));
  OAI210     g055(.A0(new_new_n70_), .A1(new_new_n69_), .B0(new_new_n77_), .Y(new_new_n78_));
  OAI210     g056(.A0(new_new_n78_), .A1(new_new_n68_), .B0(i_0_), .Y(new_new_n79_));
  NA2        g057(.A(i_12_), .B(i_5_), .Y(new_new_n80_));
  NA2        g058(.A(i_2_), .B(i_8_), .Y(new_new_n81_));
  NO2        g059(.A(new_new_n81_), .B(new_new_n58_), .Y(new_new_n82_));
  NO2        g060(.A(i_3_), .B(i_9_), .Y(new_new_n83_));
  NO2        g061(.A(i_3_), .B(i_7_), .Y(new_new_n84_));
  NO3        g062(.A(new_new_n84_), .B(new_new_n83_), .C(new_new_n63_), .Y(new_new_n85_));
  INV        g063(.A(i_6_), .Y(new_new_n86_));
  OR4        g064(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(new_new_n87_));
  INV        g065(.A(new_new_n87_), .Y(new_new_n88_));
  NO2        g066(.A(i_2_), .B(i_7_), .Y(new_new_n89_));
  NO2        g067(.A(new_new_n88_), .B(new_new_n89_), .Y(new_new_n90_));
  OAI210     g068(.A0(new_new_n85_), .A1(new_new_n82_), .B0(new_new_n90_), .Y(new_new_n91_));
  NAi21      g069(.An(i_6_), .B(i_10_), .Y(new_new_n92_));
  NA2        g070(.A(i_6_), .B(i_9_), .Y(new_new_n93_));
  AOI210     g071(.A0(new_new_n93_), .A1(new_new_n92_), .B0(new_new_n63_), .Y(new_new_n94_));
  NA2        g072(.A(i_2_), .B(i_6_), .Y(new_new_n95_));
  NO3        g073(.A(new_new_n95_), .B(new_new_n49_), .C(new_new_n25_), .Y(new_new_n96_));
  NO2        g074(.A(new_new_n96_), .B(new_new_n94_), .Y(new_new_n97_));
  AOI210     g075(.A0(new_new_n97_), .A1(new_new_n91_), .B0(new_new_n80_), .Y(new_new_n98_));
  AN3        g076(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n99_));
  NAi21      g077(.An(i_6_), .B(i_11_), .Y(new_new_n100_));
  NO2        g078(.A(i_5_), .B(i_8_), .Y(new_new_n101_));
  NOi21      g079(.An(new_new_n101_), .B(new_new_n100_), .Y(new_new_n102_));
  AOI220     g080(.A0(new_new_n102_), .A1(new_new_n62_), .B0(new_new_n99_), .B1(new_new_n32_), .Y(new_new_n103_));
  INV        g081(.A(i_7_), .Y(new_new_n104_));
  NA2        g082(.A(new_new_n46_), .B(new_new_n104_), .Y(new_new_n105_));
  NO2        g083(.A(i_0_), .B(i_5_), .Y(new_new_n106_));
  NO2        g084(.A(new_new_n106_), .B(new_new_n86_), .Y(new_new_n107_));
  NA2        g085(.A(i_12_), .B(i_3_), .Y(new_new_n108_));
  INV        g086(.A(new_new_n108_), .Y(new_new_n109_));
  NA3        g087(.A(new_new_n109_), .B(new_new_n107_), .C(new_new_n105_), .Y(new_new_n110_));
  NAi21      g088(.An(i_7_), .B(i_11_), .Y(new_new_n111_));
  NO3        g089(.A(new_new_n111_), .B(new_new_n92_), .C(new_new_n53_), .Y(new_new_n112_));
  AN2        g090(.A(i_2_), .B(i_10_), .Y(new_new_n113_));
  NO2        g091(.A(new_new_n113_), .B(i_7_), .Y(new_new_n114_));
  OR2        g092(.A(new_new_n80_), .B(new_new_n58_), .Y(new_new_n115_));
  NO2        g093(.A(i_8_), .B(new_new_n104_), .Y(new_new_n116_));
  NO3        g094(.A(new_new_n116_), .B(new_new_n115_), .C(new_new_n114_), .Y(new_new_n117_));
  NA2        g095(.A(i_12_), .B(i_7_), .Y(new_new_n118_));
  NO2        g096(.A(new_new_n63_), .B(new_new_n26_), .Y(new_new_n119_));
  NA2        g097(.A(new_new_n119_), .B(i_0_), .Y(new_new_n120_));
  NA2        g098(.A(i_11_), .B(i_12_), .Y(new_new_n121_));
  OAI210     g099(.A0(new_new_n120_), .A1(new_new_n118_), .B0(new_new_n121_), .Y(new_new_n122_));
  NO2        g100(.A(new_new_n122_), .B(new_new_n117_), .Y(new_new_n123_));
  NAi41      g101(.An(new_new_n112_), .B(new_new_n123_), .C(new_new_n110_), .D(new_new_n103_), .Y(new_new_n124_));
  NOi21      g102(.An(i_1_), .B(i_5_), .Y(new_new_n125_));
  NA2        g103(.A(new_new_n125_), .B(i_11_), .Y(new_new_n126_));
  NA2        g104(.A(new_new_n104_), .B(new_new_n37_), .Y(new_new_n127_));
  NA2        g105(.A(i_7_), .B(new_new_n25_), .Y(new_new_n128_));
  NA2        g106(.A(new_new_n128_), .B(new_new_n127_), .Y(new_new_n129_));
  NO2        g107(.A(new_new_n129_), .B(new_new_n46_), .Y(new_new_n130_));
  NA2        g108(.A(new_new_n93_), .B(new_new_n92_), .Y(new_new_n131_));
  NAi21      g109(.An(i_3_), .B(i_8_), .Y(new_new_n132_));
  NA2        g110(.A(new_new_n132_), .B(new_new_n62_), .Y(new_new_n133_));
  NOi31      g111(.An(new_new_n133_), .B(new_new_n131_), .C(new_new_n130_), .Y(new_new_n134_));
  NO2        g112(.A(i_1_), .B(new_new_n86_), .Y(new_new_n135_));
  NO2        g113(.A(i_6_), .B(i_5_), .Y(new_new_n136_));
  NA2        g114(.A(new_new_n136_), .B(i_3_), .Y(new_new_n137_));
  AO210      g115(.A0(new_new_n137_), .A1(new_new_n47_), .B0(new_new_n135_), .Y(new_new_n138_));
  OAI220     g116(.A0(new_new_n138_), .A1(new_new_n111_), .B0(new_new_n134_), .B1(new_new_n126_), .Y(new_new_n139_));
  NO3        g117(.A(new_new_n139_), .B(new_new_n124_), .C(new_new_n98_), .Y(new_new_n140_));
  NA3        g118(.A(new_new_n140_), .B(new_new_n79_), .C(new_new_n56_), .Y(ori2));
  NO2        g119(.A(new_new_n63_), .B(new_new_n37_), .Y(new_new_n142_));
  INV        g120(.A(i_6_), .Y(new_new_n143_));
  NA2        g121(.A(new_new_n143_), .B(new_new_n142_), .Y(new_new_n144_));
  NA4        g122(.A(new_new_n144_), .B(new_new_n77_), .C(new_new_n69_), .D(new_new_n30_), .Y(ori0));
  AN2        g123(.A(i_8_), .B(i_7_), .Y(new_new_n146_));
  NA2        g124(.A(new_new_n146_), .B(i_6_), .Y(new_new_n147_));
  NO2        g125(.A(i_12_), .B(i_13_), .Y(new_new_n148_));
  NAi21      g126(.An(i_5_), .B(i_11_), .Y(new_new_n149_));
  NOi21      g127(.An(new_new_n148_), .B(new_new_n149_), .Y(new_new_n150_));
  NO2        g128(.A(i_0_), .B(i_1_), .Y(new_new_n151_));
  NA2        g129(.A(i_2_), .B(i_3_), .Y(new_new_n152_));
  NO2        g130(.A(new_new_n152_), .B(i_4_), .Y(new_new_n153_));
  NA3        g131(.A(new_new_n153_), .B(new_new_n151_), .C(new_new_n150_), .Y(new_new_n154_));
  AN2        g132(.A(new_new_n148_), .B(new_new_n83_), .Y(new_new_n155_));
  NA2        g133(.A(i_1_), .B(i_5_), .Y(new_new_n156_));
  OR2        g134(.A(i_0_), .B(i_1_), .Y(new_new_n157_));
  NO3        g135(.A(new_new_n157_), .B(new_new_n80_), .C(i_13_), .Y(new_new_n158_));
  NAi32      g136(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(new_new_n159_));
  NAi21      g137(.An(new_new_n159_), .B(new_new_n158_), .Y(new_new_n160_));
  NOi21      g138(.An(i_4_), .B(i_10_), .Y(new_new_n161_));
  NA2        g139(.A(new_new_n161_), .B(new_new_n40_), .Y(new_new_n162_));
  NO3        g140(.A(new_new_n73_), .B(i_2_), .C(i_1_), .Y(new_new_n163_));
  NO2        g141(.A(new_new_n160_), .B(new_new_n147_), .Y(new_new_n164_));
  NOi21      g142(.An(i_4_), .B(i_9_), .Y(new_new_n165_));
  NOi21      g143(.An(i_11_), .B(i_13_), .Y(new_new_n166_));
  NA2        g144(.A(new_new_n166_), .B(new_new_n165_), .Y(new_new_n167_));
  NO2        g145(.A(i_4_), .B(i_5_), .Y(new_new_n168_));
  NAi21      g146(.An(i_12_), .B(i_11_), .Y(new_new_n169_));
  NO2        g147(.A(new_new_n169_), .B(i_13_), .Y(new_new_n170_));
  NO2        g148(.A(new_new_n73_), .B(new_new_n63_), .Y(new_new_n171_));
  NA2        g149(.A(new_new_n171_), .B(new_new_n46_), .Y(new_new_n172_));
  NA2        g150(.A(i_3_), .B(i_5_), .Y(new_new_n173_));
  NO2        g151(.A(new_new_n73_), .B(i_5_), .Y(new_new_n174_));
  NO2        g152(.A(i_13_), .B(i_10_), .Y(new_new_n175_));
  NA3        g153(.A(new_new_n175_), .B(new_new_n174_), .C(new_new_n44_), .Y(new_new_n176_));
  NO2        g154(.A(i_2_), .B(i_1_), .Y(new_new_n177_));
  NA2        g155(.A(new_new_n177_), .B(i_3_), .Y(new_new_n178_));
  NAi21      g156(.An(i_4_), .B(i_12_), .Y(new_new_n179_));
  INV        g157(.A(i_8_), .Y(new_new_n180_));
  NO3        g158(.A(i_3_), .B(new_new_n86_), .C(new_new_n48_), .Y(new_new_n181_));
  NA2        g159(.A(new_new_n181_), .B(new_new_n116_), .Y(new_new_n182_));
  NO3        g160(.A(i_0_), .B(i_2_), .C(i_1_), .Y(new_new_n183_));
  NO3        g161(.A(i_11_), .B(i_13_), .C(i_9_), .Y(new_new_n184_));
  NA2        g162(.A(i_12_), .B(new_new_n184_), .Y(new_new_n185_));
  NO2        g163(.A(new_new_n185_), .B(new_new_n182_), .Y(new_new_n186_));
  NO2        g164(.A(i_3_), .B(i_8_), .Y(new_new_n187_));
  NO3        g165(.A(i_11_), .B(i_10_), .C(i_9_), .Y(new_new_n188_));
  NA3        g166(.A(new_new_n188_), .B(new_new_n187_), .C(new_new_n40_), .Y(new_new_n189_));
  NO2        g167(.A(new_new_n106_), .B(new_new_n58_), .Y(new_new_n190_));
  INV        g168(.A(new_new_n190_), .Y(new_new_n191_));
  NO2        g169(.A(i_13_), .B(i_9_), .Y(new_new_n192_));
  NAi21      g170(.An(i_12_), .B(i_3_), .Y(new_new_n193_));
  NO2        g171(.A(new_new_n44_), .B(i_5_), .Y(new_new_n194_));
  NO2        g172(.A(new_new_n191_), .B(new_new_n189_), .Y(new_new_n195_));
  AOI210     g173(.A0(new_new_n195_), .A1(i_7_), .B0(new_new_n186_), .Y(new_new_n196_));
  NO2        g174(.A(new_new_n196_), .B(i_4_), .Y(new_new_n197_));
  NAi21      g175(.An(i_12_), .B(i_7_), .Y(new_new_n198_));
  NA3        g176(.A(i_13_), .B(new_new_n180_), .C(i_10_), .Y(new_new_n199_));
  NO2        g177(.A(new_new_n199_), .B(new_new_n198_), .Y(new_new_n200_));
  NA2        g178(.A(i_0_), .B(i_5_), .Y(new_new_n201_));
  NA2        g179(.A(new_new_n201_), .B(new_new_n107_), .Y(new_new_n202_));
  OAI220     g180(.A0(new_new_n202_), .A1(new_new_n178_), .B0(new_new_n172_), .B1(new_new_n137_), .Y(new_new_n203_));
  NAi31      g181(.An(i_9_), .B(i_6_), .C(i_5_), .Y(new_new_n204_));
  NO2        g182(.A(new_new_n36_), .B(i_13_), .Y(new_new_n205_));
  NO2        g183(.A(new_new_n73_), .B(new_new_n26_), .Y(new_new_n206_));
  NO2        g184(.A(new_new_n46_), .B(new_new_n63_), .Y(new_new_n207_));
  INV        g185(.A(i_13_), .Y(new_new_n208_));
  NO2        g186(.A(i_12_), .B(new_new_n208_), .Y(new_new_n209_));
  NA3        g187(.A(new_new_n209_), .B(new_new_n183_), .C(new_new_n181_), .Y(new_new_n210_));
  INV        g188(.A(new_new_n210_), .Y(new_new_n211_));
  AOI220     g189(.A0(new_new_n211_), .A1(new_new_n146_), .B0(new_new_n203_), .B1(new_new_n200_), .Y(new_new_n212_));
  NO2        g190(.A(i_12_), .B(new_new_n37_), .Y(new_new_n213_));
  OR2        g191(.A(i_8_), .B(i_7_), .Y(new_new_n214_));
  INV        g192(.A(i_12_), .Y(new_new_n215_));
  NO2        g193(.A(new_new_n44_), .B(new_new_n215_), .Y(new_new_n216_));
  NO3        g194(.A(new_new_n36_), .B(i_8_), .C(i_10_), .Y(new_new_n217_));
  NA2        g195(.A(i_2_), .B(i_1_), .Y(new_new_n218_));
  NO3        g196(.A(i_11_), .B(i_7_), .C(new_new_n37_), .Y(new_new_n219_));
  NAi21      g197(.An(i_4_), .B(i_3_), .Y(new_new_n220_));
  NO2        g198(.A(i_0_), .B(i_6_), .Y(new_new_n221_));
  NOi41      g199(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(new_new_n222_));
  NA2        g200(.A(new_new_n222_), .B(new_new_n221_), .Y(new_new_n223_));
  NO2        g201(.A(new_new_n218_), .B(new_new_n173_), .Y(new_new_n224_));
  NO2        g202(.A(i_11_), .B(new_new_n208_), .Y(new_new_n225_));
  NOi21      g203(.An(i_1_), .B(i_6_), .Y(new_new_n226_));
  NAi21      g204(.An(i_3_), .B(i_7_), .Y(new_new_n227_));
  NA2        g205(.A(new_new_n215_), .B(i_9_), .Y(new_new_n228_));
  OR4        g206(.A(new_new_n228_), .B(new_new_n227_), .C(new_new_n226_), .D(new_new_n174_), .Y(new_new_n229_));
  NA2        g207(.A(new_new_n73_), .B(i_5_), .Y(new_new_n230_));
  NA2        g208(.A(i_3_), .B(i_9_), .Y(new_new_n231_));
  NAi21      g209(.An(i_7_), .B(i_10_), .Y(new_new_n232_));
  NO2        g210(.A(new_new_n232_), .B(new_new_n231_), .Y(new_new_n233_));
  NA3        g211(.A(new_new_n233_), .B(new_new_n230_), .C(new_new_n64_), .Y(new_new_n234_));
  NA2        g212(.A(new_new_n234_), .B(new_new_n229_), .Y(new_new_n235_));
  INV        g213(.A(new_new_n147_), .Y(new_new_n236_));
  NA2        g214(.A(new_new_n215_), .B(i_13_), .Y(new_new_n237_));
  NO2        g215(.A(new_new_n237_), .B(new_new_n75_), .Y(new_new_n238_));
  AOI220     g216(.A0(new_new_n238_), .A1(new_new_n236_), .B0(new_new_n235_), .B1(new_new_n225_), .Y(new_new_n239_));
  NO2        g217(.A(new_new_n214_), .B(new_new_n37_), .Y(new_new_n240_));
  NA2        g218(.A(i_12_), .B(i_6_), .Y(new_new_n241_));
  OR2        g219(.A(i_13_), .B(i_9_), .Y(new_new_n242_));
  NO3        g220(.A(new_new_n242_), .B(new_new_n241_), .C(new_new_n48_), .Y(new_new_n243_));
  NO2        g221(.A(new_new_n220_), .B(i_2_), .Y(new_new_n244_));
  NA3        g222(.A(new_new_n244_), .B(new_new_n243_), .C(new_new_n44_), .Y(new_new_n245_));
  NA2        g223(.A(new_new_n225_), .B(i_9_), .Y(new_new_n246_));
  NA2        g224(.A(new_new_n230_), .B(new_new_n64_), .Y(new_new_n247_));
  OAI210     g225(.A0(new_new_n247_), .A1(new_new_n246_), .B0(new_new_n245_), .Y(new_new_n248_));
  NO3        g226(.A(i_11_), .B(new_new_n208_), .C(new_new_n25_), .Y(new_new_n249_));
  NO2        g227(.A(new_new_n227_), .B(i_8_), .Y(new_new_n250_));
  NA2        g228(.A(new_new_n248_), .B(new_new_n240_), .Y(new_new_n251_));
  NA3        g229(.A(new_new_n251_), .B(new_new_n239_), .C(new_new_n212_), .Y(new_new_n252_));
  NO3        g230(.A(i_12_), .B(new_new_n208_), .C(new_new_n37_), .Y(new_new_n253_));
  NO2        g231(.A(new_new_n218_), .B(i_0_), .Y(new_new_n254_));
  NO2        g232(.A(i_2_), .B(new_new_n104_), .Y(new_new_n255_));
  AN2        g233(.A(i_3_), .B(i_10_), .Y(new_new_n256_));
  NO2        g234(.A(i_5_), .B(new_new_n37_), .Y(new_new_n257_));
  NO2        g235(.A(new_new_n46_), .B(new_new_n26_), .Y(new_new_n258_));
  NO3        g236(.A(new_new_n252_), .B(new_new_n197_), .C(new_new_n164_), .Y(new_new_n259_));
  NO3        g237(.A(new_new_n44_), .B(i_13_), .C(i_9_), .Y(new_new_n260_));
  NO2        g238(.A(i_2_), .B(i_3_), .Y(new_new_n261_));
  OR2        g239(.A(i_0_), .B(i_5_), .Y(new_new_n262_));
  NO2        g240(.A(new_new_n157_), .B(new_new_n46_), .Y(new_new_n263_));
  NO2        g241(.A(i_12_), .B(i_10_), .Y(new_new_n264_));
  NOi21      g242(.An(i_5_), .B(i_0_), .Y(new_new_n265_));
  NA4        g243(.A(new_new_n84_), .B(new_new_n36_), .C(new_new_n86_), .D(i_8_), .Y(new_new_n266_));
  NO2        g244(.A(i_6_), .B(i_8_), .Y(new_new_n267_));
  NO2        g245(.A(i_1_), .B(i_7_), .Y(new_new_n268_));
  NOi21      g246(.An(new_new_n156_), .B(new_new_n107_), .Y(new_new_n269_));
  NO2        g247(.A(new_new_n269_), .B(new_new_n128_), .Y(new_new_n270_));
  NA2        g248(.A(new_new_n270_), .B(i_3_), .Y(new_new_n271_));
  NO2        g249(.A(new_new_n180_), .B(i_9_), .Y(new_new_n272_));
  NA2        g250(.A(new_new_n272_), .B(new_new_n190_), .Y(new_new_n273_));
  NO2        g251(.A(new_new_n273_), .B(new_new_n46_), .Y(new_new_n274_));
  INV        g252(.A(new_new_n274_), .Y(new_new_n275_));
  AOI210     g253(.A0(new_new_n275_), .A1(new_new_n271_), .B0(new_new_n162_), .Y(new_new_n276_));
  INV        g254(.A(new_new_n276_), .Y(new_new_n277_));
  NOi32      g255(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(new_new_n278_));
  INV        g256(.A(new_new_n278_), .Y(new_new_n279_));
  NAi21      g257(.An(i_0_), .B(i_6_), .Y(new_new_n280_));
  NAi21      g258(.An(i_1_), .B(i_5_), .Y(new_new_n281_));
  NA2        g259(.A(new_new_n281_), .B(new_new_n280_), .Y(new_new_n282_));
  NA2        g260(.A(new_new_n282_), .B(new_new_n25_), .Y(new_new_n283_));
  OAI210     g261(.A0(new_new_n283_), .A1(new_new_n159_), .B0(new_new_n223_), .Y(new_new_n284_));
  NAi41      g262(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(new_new_n285_));
  OAI220     g263(.A0(new_new_n285_), .A1(new_new_n281_), .B0(new_new_n204_), .B1(new_new_n159_), .Y(new_new_n286_));
  AOI210     g264(.A0(new_new_n285_), .A1(new_new_n159_), .B0(new_new_n157_), .Y(new_new_n287_));
  NOi32      g265(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(new_new_n288_));
  NAi21      g266(.An(i_6_), .B(i_1_), .Y(new_new_n289_));
  NA3        g267(.A(new_new_n289_), .B(new_new_n288_), .C(new_new_n46_), .Y(new_new_n290_));
  NO2        g268(.A(new_new_n290_), .B(i_0_), .Y(new_new_n291_));
  OR3        g269(.A(new_new_n291_), .B(new_new_n287_), .C(new_new_n286_), .Y(new_new_n292_));
  NO2        g270(.A(i_1_), .B(new_new_n104_), .Y(new_new_n293_));
  NAi21      g271(.An(i_3_), .B(i_4_), .Y(new_new_n294_));
  NO2        g272(.A(new_new_n294_), .B(i_9_), .Y(new_new_n295_));
  AN2        g273(.A(i_6_), .B(i_7_), .Y(new_new_n296_));
  OAI210     g274(.A0(new_new_n296_), .A1(new_new_n293_), .B0(new_new_n295_), .Y(new_new_n297_));
  NA2        g275(.A(i_2_), .B(i_7_), .Y(new_new_n298_));
  NO2        g276(.A(new_new_n294_), .B(i_10_), .Y(new_new_n299_));
  NA3        g277(.A(new_new_n299_), .B(new_new_n298_), .C(new_new_n221_), .Y(new_new_n300_));
  AOI210     g278(.A0(new_new_n300_), .A1(new_new_n297_), .B0(new_new_n174_), .Y(new_new_n301_));
  AOI210     g279(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(new_new_n302_));
  OAI210     g280(.A0(new_new_n302_), .A1(new_new_n177_), .B0(new_new_n299_), .Y(new_new_n303_));
  AOI220     g281(.A0(new_new_n299_), .A1(new_new_n268_), .B0(new_new_n217_), .B1(new_new_n177_), .Y(new_new_n304_));
  AOI210     g282(.A0(new_new_n304_), .A1(new_new_n303_), .B0(i_5_), .Y(new_new_n305_));
  NO4        g283(.A(new_new_n305_), .B(new_new_n301_), .C(new_new_n292_), .D(new_new_n284_), .Y(new_new_n306_));
  NO2        g284(.A(new_new_n306_), .B(new_new_n279_), .Y(new_new_n307_));
  NO2        g285(.A(new_new_n59_), .B(new_new_n25_), .Y(new_new_n308_));
  AN2        g286(.A(i_12_), .B(i_5_), .Y(new_new_n309_));
  NO2        g287(.A(i_4_), .B(new_new_n26_), .Y(new_new_n310_));
  NA2        g288(.A(new_new_n310_), .B(new_new_n309_), .Y(new_new_n311_));
  NO2        g289(.A(i_11_), .B(i_6_), .Y(new_new_n312_));
  NA3        g290(.A(new_new_n312_), .B(new_new_n263_), .C(new_new_n208_), .Y(new_new_n313_));
  NO2        g291(.A(new_new_n313_), .B(new_new_n311_), .Y(new_new_n314_));
  NO2        g292(.A(i_5_), .B(i_10_), .Y(new_new_n315_));
  NO2        g293(.A(new_new_n37_), .B(new_new_n25_), .Y(new_new_n316_));
  NO2        g294(.A(new_new_n154_), .B(new_new_n86_), .Y(new_new_n317_));
  OAI210     g295(.A0(new_new_n317_), .A1(new_new_n314_), .B0(new_new_n316_), .Y(new_new_n318_));
  NO3        g296(.A(new_new_n86_), .B(new_new_n48_), .C(i_9_), .Y(new_new_n319_));
  NO2        g297(.A(i_11_), .B(i_12_), .Y(new_new_n320_));
  NAi21      g298(.An(i_13_), .B(i_0_), .Y(new_new_n321_));
  INV        g299(.A(new_new_n318_), .Y(new_new_n322_));
  NA2        g300(.A(new_new_n44_), .B(new_new_n208_), .Y(new_new_n323_));
  NO3        g301(.A(i_1_), .B(i_12_), .C(new_new_n86_), .Y(new_new_n324_));
  NO2        g302(.A(i_0_), .B(i_11_), .Y(new_new_n325_));
  AN2        g303(.A(i_1_), .B(i_6_), .Y(new_new_n326_));
  NOi21      g304(.An(i_2_), .B(i_12_), .Y(new_new_n327_));
  NAi21      g305(.An(i_9_), .B(i_4_), .Y(new_new_n328_));
  OR2        g306(.A(i_13_), .B(i_10_), .Y(new_new_n329_));
  NO3        g307(.A(new_new_n329_), .B(new_new_n121_), .C(new_new_n328_), .Y(new_new_n330_));
  NO2        g308(.A(new_new_n167_), .B(new_new_n127_), .Y(new_new_n331_));
  NO2        g309(.A(new_new_n104_), .B(new_new_n25_), .Y(new_new_n332_));
  NA2        g310(.A(new_new_n253_), .B(new_new_n332_), .Y(new_new_n333_));
  NO2        g311(.A(new_new_n333_), .B(new_new_n269_), .Y(new_new_n334_));
  INV        g312(.A(new_new_n334_), .Y(new_new_n335_));
  NO2        g313(.A(new_new_n335_), .B(new_new_n26_), .Y(new_new_n336_));
  NO2        g314(.A(new_new_n173_), .B(new_new_n86_), .Y(new_new_n337_));
  NA2        g315(.A(new_new_n180_), .B(i_10_), .Y(new_new_n338_));
  NA3        g316(.A(new_new_n230_), .B(new_new_n64_), .C(i_2_), .Y(new_new_n339_));
  NO2        g317(.A(new_new_n339_), .B(new_new_n338_), .Y(new_new_n340_));
  NO2        g318(.A(i_3_), .B(new_new_n48_), .Y(new_new_n341_));
  INV        g319(.A(new_new_n340_), .Y(new_new_n342_));
  NO2        g320(.A(new_new_n342_), .B(new_new_n246_), .Y(new_new_n343_));
  NO4        g321(.A(new_new_n343_), .B(new_new_n336_), .C(new_new_n322_), .D(new_new_n307_), .Y(new_new_n344_));
  NO2        g322(.A(new_new_n63_), .B(i_4_), .Y(new_new_n345_));
  NO2        g323(.A(new_new_n73_), .B(i_13_), .Y(new_new_n346_));
  NA3        g324(.A(new_new_n346_), .B(new_new_n345_), .C(i_2_), .Y(new_new_n347_));
  NO2        g325(.A(i_10_), .B(i_9_), .Y(new_new_n348_));
  NAi21      g326(.An(i_12_), .B(i_8_), .Y(new_new_n349_));
  NO2        g327(.A(new_new_n349_), .B(i_3_), .Y(new_new_n350_));
  NA2        g328(.A(new_new_n350_), .B(new_new_n348_), .Y(new_new_n351_));
  NO2        g329(.A(new_new_n46_), .B(i_4_), .Y(new_new_n352_));
  NA2        g330(.A(new_new_n352_), .B(new_new_n107_), .Y(new_new_n353_));
  OAI220     g331(.A0(new_new_n353_), .A1(new_new_n189_), .B0(new_new_n351_), .B1(new_new_n347_), .Y(new_new_n354_));
  NA2        g332(.A(new_new_n258_), .B(i_0_), .Y(new_new_n355_));
  NO3        g333(.A(new_new_n23_), .B(i_10_), .C(i_9_), .Y(new_new_n356_));
  NA2        g334(.A(new_new_n241_), .B(new_new_n100_), .Y(new_new_n357_));
  NA2        g335(.A(new_new_n357_), .B(new_new_n356_), .Y(new_new_n358_));
  NA2        g336(.A(i_8_), .B(i_9_), .Y(new_new_n359_));
  AOI210     g337(.A0(i_0_), .A1(i_7_), .B0(i_2_), .Y(new_new_n360_));
  OR2        g338(.A(new_new_n360_), .B(new_new_n359_), .Y(new_new_n361_));
  NA2        g339(.A(new_new_n253_), .B(new_new_n190_), .Y(new_new_n362_));
  OAI220     g340(.A0(new_new_n362_), .A1(new_new_n361_), .B0(new_new_n358_), .B1(new_new_n355_), .Y(new_new_n363_));
  NA2        g341(.A(new_new_n225_), .B(new_new_n257_), .Y(new_new_n364_));
  NO3        g342(.A(i_6_), .B(i_8_), .C(i_7_), .Y(new_new_n365_));
  INV        g343(.A(new_new_n365_), .Y(new_new_n366_));
  NA3        g344(.A(i_2_), .B(i_10_), .C(i_9_), .Y(new_new_n367_));
  NA4        g345(.A(new_new_n149_), .B(new_new_n119_), .C(new_new_n80_), .D(new_new_n23_), .Y(new_new_n368_));
  OAI220     g346(.A0(new_new_n368_), .A1(new_new_n367_), .B0(new_new_n366_), .B1(new_new_n364_), .Y(new_new_n369_));
  NO3        g347(.A(new_new_n369_), .B(new_new_n363_), .C(new_new_n354_), .Y(new_new_n370_));
  OR2        g348(.A(new_new_n273_), .B(new_new_n104_), .Y(new_new_n371_));
  OR2        g349(.A(new_new_n371_), .B(new_new_n162_), .Y(new_new_n372_));
  NA2        g350(.A(new_new_n99_), .B(i_13_), .Y(new_new_n373_));
  NA2        g351(.A(new_new_n337_), .B(new_new_n308_), .Y(new_new_n374_));
  NO2        g352(.A(i_2_), .B(i_13_), .Y(new_new_n375_));
  NO2        g353(.A(new_new_n374_), .B(new_new_n373_), .Y(new_new_n376_));
  NO3        g354(.A(i_4_), .B(new_new_n48_), .C(i_8_), .Y(new_new_n377_));
  NO2        g355(.A(i_6_), .B(i_7_), .Y(new_new_n378_));
  NO2        g356(.A(i_11_), .B(i_1_), .Y(new_new_n379_));
  OR2        g357(.A(i_11_), .B(i_8_), .Y(new_new_n380_));
  NOi21      g358(.An(i_2_), .B(i_7_), .Y(new_new_n381_));
  NO2        g359(.A(i_3_), .B(new_new_n180_), .Y(new_new_n382_));
  NO2        g360(.A(i_6_), .B(i_10_), .Y(new_new_n383_));
  NA3        g361(.A(new_new_n222_), .B(new_new_n166_), .C(new_new_n136_), .Y(new_new_n384_));
  NA2        g362(.A(new_new_n46_), .B(new_new_n44_), .Y(new_new_n385_));
  NO2        g363(.A(new_new_n157_), .B(i_3_), .Y(new_new_n386_));
  NAi31      g364(.An(new_new_n385_), .B(new_new_n386_), .C(new_new_n209_), .Y(new_new_n387_));
  NA3        g365(.A(new_new_n316_), .B(new_new_n171_), .C(new_new_n153_), .Y(new_new_n388_));
  NA3        g366(.A(new_new_n388_), .B(new_new_n387_), .C(new_new_n384_), .Y(new_new_n389_));
  NO2        g367(.A(new_new_n389_), .B(new_new_n376_), .Y(new_new_n390_));
  NA2        g368(.A(new_new_n356_), .B(new_new_n309_), .Y(new_new_n391_));
  NA2        g369(.A(new_new_n365_), .B(new_new_n315_), .Y(new_new_n392_));
  NAi21      g370(.An(new_new_n199_), .B(new_new_n320_), .Y(new_new_n393_));
  NA2        g371(.A(new_new_n268_), .B(new_new_n201_), .Y(new_new_n394_));
  NO2        g372(.A(new_new_n394_), .B(new_new_n393_), .Y(new_new_n395_));
  NA2        g373(.A(new_new_n27_), .B(i_10_), .Y(new_new_n396_));
  NA2        g374(.A(new_new_n260_), .B(new_new_n217_), .Y(new_new_n397_));
  OAI220     g375(.A0(new_new_n397_), .A1(new_new_n339_), .B0(new_new_n396_), .B1(new_new_n373_), .Y(new_new_n398_));
  NO2        g376(.A(new_new_n398_), .B(new_new_n395_), .Y(new_new_n399_));
  NA4        g377(.A(new_new_n399_), .B(new_new_n390_), .C(new_new_n372_), .D(new_new_n370_), .Y(new_new_n400_));
  NA2        g378(.A(new_new_n126_), .B(new_new_n115_), .Y(new_new_n401_));
  AN2        g379(.A(new_new_n401_), .B(new_new_n356_), .Y(new_new_n402_));
  NA2        g380(.A(new_new_n402_), .B(new_new_n258_), .Y(new_new_n403_));
  NA4        g381(.A(new_new_n346_), .B(new_new_n345_), .C(new_new_n187_), .D(i_2_), .Y(new_new_n404_));
  INV        g382(.A(new_new_n404_), .Y(new_new_n405_));
  NA2        g383(.A(new_new_n309_), .B(new_new_n208_), .Y(new_new_n406_));
  NA2        g384(.A(new_new_n278_), .B(new_new_n73_), .Y(new_new_n407_));
  NA2        g385(.A(new_new_n296_), .B(new_new_n288_), .Y(new_new_n408_));
  OR2        g386(.A(new_new_n406_), .B(new_new_n408_), .Y(new_new_n409_));
  NO2        g387(.A(new_new_n36_), .B(i_8_), .Y(new_new_n410_));
  AOI210     g388(.A0(new_new_n39_), .A1(i_13_), .B0(new_new_n330_), .Y(new_new_n411_));
  NA2        g389(.A(new_new_n411_), .B(new_new_n409_), .Y(new_new_n412_));
  AOI210     g390(.A0(new_new_n405_), .A1(new_new_n188_), .B0(new_new_n412_), .Y(new_new_n413_));
  NA2        g391(.A(new_new_n230_), .B(new_new_n64_), .Y(new_new_n414_));
  OAI210     g392(.A0(i_8_), .A1(new_new_n414_), .B0(new_new_n138_), .Y(new_new_n415_));
  NA2        g393(.A(new_new_n415_), .B(new_new_n331_), .Y(new_new_n416_));
  NA3        g394(.A(new_new_n416_), .B(new_new_n413_), .C(new_new_n403_), .Y(new_new_n417_));
  NO2        g395(.A(i_12_), .B(new_new_n180_), .Y(new_new_n418_));
  NO2        g396(.A(i_8_), .B(i_7_), .Y(new_new_n419_));
  NA2        g397(.A(new_new_n44_), .B(i_10_), .Y(new_new_n420_));
  NO2        g398(.A(new_new_n420_), .B(i_6_), .Y(new_new_n421_));
  AOI220     g399(.A0(new_new_n337_), .A1(new_new_n263_), .B0(new_new_n224_), .B1(new_new_n221_), .Y(new_new_n422_));
  OAI220     g400(.A0(new_new_n422_), .A1(new_new_n237_), .B0(new_new_n373_), .B1(new_new_n137_), .Y(new_new_n423_));
  NA2        g401(.A(new_new_n423_), .B(new_new_n240_), .Y(new_new_n424_));
  NA3        g402(.A(new_new_n256_), .B(new_new_n168_), .C(new_new_n99_), .Y(new_new_n425_));
  NO2        g403(.A(new_new_n205_), .B(new_new_n44_), .Y(new_new_n426_));
  NO2        g404(.A(new_new_n157_), .B(i_5_), .Y(new_new_n427_));
  NA3        g405(.A(new_new_n427_), .B(new_new_n323_), .C(new_new_n261_), .Y(new_new_n428_));
  OAI210     g406(.A0(new_new_n428_), .A1(new_new_n426_), .B0(new_new_n425_), .Y(new_new_n429_));
  NA2        g407(.A(new_new_n429_), .B(new_new_n365_), .Y(new_new_n430_));
  NA2        g408(.A(new_new_n430_), .B(new_new_n424_), .Y(new_new_n431_));
  NA3        g409(.A(new_new_n201_), .B(new_new_n71_), .C(new_new_n44_), .Y(new_new_n432_));
  NA2        g410(.A(new_new_n253_), .B(new_new_n84_), .Y(new_new_n433_));
  NO2        g411(.A(new_new_n432_), .B(new_new_n433_), .Y(new_new_n434_));
  NA2        g412(.A(new_new_n207_), .B(new_new_n206_), .Y(new_new_n435_));
  NA2        g413(.A(new_new_n348_), .B(new_new_n205_), .Y(new_new_n436_));
  NO2        g414(.A(new_new_n435_), .B(new_new_n436_), .Y(new_new_n437_));
  AOI210     g415(.A0(new_new_n289_), .A1(new_new_n46_), .B0(new_new_n293_), .Y(new_new_n438_));
  NA2        g416(.A(i_0_), .B(new_new_n48_), .Y(new_new_n439_));
  NA3        g417(.A(new_new_n418_), .B(new_new_n249_), .C(new_new_n439_), .Y(new_new_n440_));
  NO2        g418(.A(new_new_n438_), .B(new_new_n440_), .Y(new_new_n441_));
  NO3        g419(.A(new_new_n441_), .B(new_new_n437_), .C(new_new_n434_), .Y(new_new_n442_));
  NO4        g420(.A(new_new_n226_), .B(new_new_n42_), .C(i_2_), .D(new_new_n48_), .Y(new_new_n443_));
  NO3        g421(.A(i_1_), .B(i_5_), .C(i_10_), .Y(new_new_n444_));
  NO2        g422(.A(new_new_n329_), .B(i_1_), .Y(new_new_n445_));
  NOi31      g423(.An(new_new_n445_), .B(new_new_n357_), .C(new_new_n73_), .Y(new_new_n446_));
  NOi21      g424(.An(i_10_), .B(i_6_), .Y(new_new_n447_));
  NO2        g425(.A(new_new_n86_), .B(new_new_n25_), .Y(new_new_n448_));
  AOI220     g426(.A0(new_new_n253_), .A1(new_new_n448_), .B0(new_new_n249_), .B1(new_new_n447_), .Y(new_new_n449_));
  NO2        g427(.A(new_new_n449_), .B(new_new_n355_), .Y(new_new_n450_));
  NO2        g428(.A(new_new_n118_), .B(new_new_n23_), .Y(new_new_n451_));
  NO2        g429(.A(new_new_n183_), .B(new_new_n37_), .Y(new_new_n452_));
  NOi31      g430(.An(new_new_n150_), .B(new_new_n452_), .C(new_new_n266_), .Y(new_new_n453_));
  NO2        g431(.A(new_new_n453_), .B(new_new_n450_), .Y(new_new_n454_));
  NO2        g432(.A(new_new_n407_), .B(new_new_n304_), .Y(new_new_n455_));
  INV        g433(.A(new_new_n261_), .Y(new_new_n456_));
  NO2        g434(.A(i_12_), .B(new_new_n86_), .Y(new_new_n457_));
  NA3        g435(.A(new_new_n457_), .B(new_new_n249_), .C(new_new_n439_), .Y(new_new_n458_));
  NA3        g436(.A(new_new_n312_), .B(new_new_n253_), .C(new_new_n201_), .Y(new_new_n459_));
  AOI210     g437(.A0(new_new_n459_), .A1(new_new_n458_), .B0(new_new_n456_), .Y(new_new_n460_));
  OR2        g438(.A(i_2_), .B(i_5_), .Y(new_new_n461_));
  OR2        g439(.A(new_new_n461_), .B(new_new_n326_), .Y(new_new_n462_));
  AOI210     g440(.A0(new_new_n298_), .A1(new_new_n221_), .B0(new_new_n183_), .Y(new_new_n463_));
  AOI210     g441(.A0(new_new_n463_), .A1(new_new_n462_), .B0(new_new_n393_), .Y(new_new_n464_));
  NO3        g442(.A(new_new_n464_), .B(new_new_n460_), .C(new_new_n455_), .Y(new_new_n465_));
  NA3        g443(.A(new_new_n465_), .B(new_new_n454_), .C(new_new_n442_), .Y(new_new_n466_));
  NO4        g444(.A(new_new_n466_), .B(new_new_n431_), .C(new_new_n417_), .D(new_new_n400_), .Y(new_new_n467_));
  NA4        g445(.A(new_new_n467_), .B(new_new_n344_), .C(new_new_n277_), .D(new_new_n259_), .Y(ori7));
  NO2        g446(.A(new_new_n95_), .B(new_new_n54_), .Y(new_new_n469_));
  NO2        g447(.A(new_new_n111_), .B(new_new_n92_), .Y(new_new_n470_));
  NA2        g448(.A(new_new_n310_), .B(new_new_n470_), .Y(new_new_n471_));
  NA2        g449(.A(new_new_n383_), .B(new_new_n84_), .Y(new_new_n472_));
  NA2        g450(.A(i_11_), .B(new_new_n180_), .Y(new_new_n473_));
  NA2        g451(.A(new_new_n148_), .B(new_new_n473_), .Y(new_new_n474_));
  OAI210     g452(.A0(new_new_n474_), .A1(new_new_n472_), .B0(new_new_n471_), .Y(new_new_n475_));
  NA3        g453(.A(i_7_), .B(i_10_), .C(i_9_), .Y(new_new_n476_));
  NO2        g454(.A(new_new_n215_), .B(i_4_), .Y(new_new_n477_));
  NA2        g455(.A(new_new_n477_), .B(i_8_), .Y(new_new_n478_));
  NO2        g456(.A(new_new_n108_), .B(new_new_n476_), .Y(new_new_n479_));
  NA2        g457(.A(i_2_), .B(new_new_n86_), .Y(new_new_n480_));
  OAI210     g458(.A0(new_new_n89_), .A1(new_new_n187_), .B0(new_new_n188_), .Y(new_new_n481_));
  NO2        g459(.A(i_7_), .B(new_new_n37_), .Y(new_new_n482_));
  NA2        g460(.A(i_4_), .B(i_8_), .Y(new_new_n483_));
  AOI210     g461(.A0(new_new_n483_), .A1(new_new_n256_), .B0(new_new_n482_), .Y(new_new_n484_));
  OAI220     g462(.A0(new_new_n484_), .A1(new_new_n480_), .B0(new_new_n481_), .B1(i_13_), .Y(new_new_n485_));
  NO4        g463(.A(new_new_n485_), .B(new_new_n479_), .C(new_new_n475_), .D(new_new_n469_), .Y(new_new_n486_));
  AOI210     g464(.A0(new_new_n132_), .A1(new_new_n62_), .B0(i_10_), .Y(new_new_n487_));
  AOI210     g465(.A0(new_new_n487_), .A1(new_new_n215_), .B0(new_new_n161_), .Y(new_new_n488_));
  OR2        g466(.A(i_6_), .B(i_10_), .Y(new_new_n489_));
  NO2        g467(.A(new_new_n489_), .B(new_new_n23_), .Y(new_new_n490_));
  OR3        g468(.A(i_13_), .B(i_6_), .C(i_10_), .Y(new_new_n491_));
  NO3        g469(.A(new_new_n491_), .B(i_8_), .C(new_new_n31_), .Y(new_new_n492_));
  INV        g470(.A(new_new_n184_), .Y(new_new_n493_));
  NO2        g471(.A(new_new_n492_), .B(new_new_n490_), .Y(new_new_n494_));
  OA220      g472(.A0(new_new_n494_), .A1(new_new_n456_), .B0(new_new_n488_), .B1(new_new_n242_), .Y(new_new_n495_));
  AOI210     g473(.A0(new_new_n495_), .A1(new_new_n486_), .B0(new_new_n63_), .Y(new_new_n496_));
  NOi21      g474(.An(i_11_), .B(i_7_), .Y(new_new_n497_));
  AO210      g475(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(new_new_n498_));
  NO2        g476(.A(new_new_n498_), .B(new_new_n497_), .Y(new_new_n499_));
  NA2        g477(.A(new_new_n499_), .B(new_new_n192_), .Y(new_new_n500_));
  NA3        g478(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n501_));
  NAi31      g479(.An(new_new_n501_), .B(new_new_n198_), .C(i_11_), .Y(new_new_n502_));
  AOI210     g480(.A0(new_new_n502_), .A1(new_new_n500_), .B0(new_new_n63_), .Y(new_new_n503_));
  NA2        g481(.A(new_new_n88_), .B(new_new_n63_), .Y(new_new_n504_));
  AO210      g482(.A0(new_new_n504_), .A1(new_new_n304_), .B0(new_new_n41_), .Y(new_new_n505_));
  NO3        g483(.A(new_new_n232_), .B(new_new_n193_), .C(new_new_n473_), .Y(new_new_n506_));
  OAI210     g484(.A0(new_new_n506_), .A1(new_new_n209_), .B0(new_new_n63_), .Y(new_new_n507_));
  NA2        g485(.A(new_new_n327_), .B(new_new_n31_), .Y(new_new_n508_));
  OR2        g486(.A(new_new_n193_), .B(new_new_n111_), .Y(new_new_n509_));
  NA2        g487(.A(new_new_n509_), .B(new_new_n508_), .Y(new_new_n510_));
  NO2        g488(.A(i_1_), .B(i_4_), .Y(new_new_n511_));
  NA2        g489(.A(new_new_n511_), .B(new_new_n510_), .Y(new_new_n512_));
  NO2        g490(.A(i_1_), .B(i_12_), .Y(new_new_n513_));
  NA3        g491(.A(new_new_n513_), .B(new_new_n113_), .C(new_new_n24_), .Y(new_new_n514_));
  BUFFER     g492(.A(new_new_n514_), .Y(new_new_n515_));
  NA4        g493(.A(new_new_n515_), .B(new_new_n512_), .C(new_new_n507_), .D(new_new_n505_), .Y(new_new_n516_));
  OAI210     g494(.A0(new_new_n516_), .A1(new_new_n503_), .B0(i_6_), .Y(new_new_n517_));
  NO2        g495(.A(new_new_n501_), .B(new_new_n111_), .Y(new_new_n518_));
  NA2        g496(.A(new_new_n518_), .B(new_new_n457_), .Y(new_new_n519_));
  NO2        g497(.A(new_new_n215_), .B(new_new_n86_), .Y(new_new_n520_));
  NO2        g498(.A(new_new_n520_), .B(i_11_), .Y(new_new_n521_));
  NA2        g499(.A(new_new_n519_), .B(new_new_n358_), .Y(new_new_n522_));
  NO3        g500(.A(new_new_n489_), .B(new_new_n214_), .C(new_new_n23_), .Y(new_new_n523_));
  AOI210     g501(.A0(i_1_), .A1(new_new_n233_), .B0(new_new_n523_), .Y(new_new_n524_));
  NO2        g502(.A(new_new_n524_), .B(new_new_n44_), .Y(new_new_n525_));
  NA3        g503(.A(new_new_n419_), .B(i_11_), .C(new_new_n36_), .Y(new_new_n526_));
  INV        g504(.A(i_2_), .Y(new_new_n527_));
  NA2        g505(.A(new_new_n142_), .B(i_9_), .Y(new_new_n528_));
  NA3        g506(.A(i_3_), .B(i_8_), .C(i_9_), .Y(new_new_n529_));
  NO2        g507(.A(new_new_n46_), .B(i_1_), .Y(new_new_n530_));
  NA3        g508(.A(new_new_n530_), .B(new_new_n241_), .C(new_new_n44_), .Y(new_new_n531_));
  OAI220     g509(.A0(new_new_n531_), .A1(new_new_n529_), .B0(new_new_n528_), .B1(new_new_n527_), .Y(new_new_n532_));
  AOI210     g510(.A0(new_new_n379_), .A1(new_new_n332_), .B0(new_new_n219_), .Y(new_new_n533_));
  NO2        g511(.A(new_new_n533_), .B(new_new_n480_), .Y(new_new_n534_));
  NAi21      g512(.An(new_new_n526_), .B(new_new_n94_), .Y(new_new_n535_));
  NA2        g513(.A(new_new_n530_), .B(new_new_n241_), .Y(new_new_n536_));
  NO2        g514(.A(i_11_), .B(new_new_n37_), .Y(new_new_n537_));
  NA2        g515(.A(new_new_n537_), .B(new_new_n24_), .Y(new_new_n538_));
  OAI210     g516(.A0(new_new_n538_), .A1(new_new_n536_), .B0(new_new_n535_), .Y(new_new_n539_));
  OR3        g517(.A(new_new_n539_), .B(new_new_n534_), .C(new_new_n532_), .Y(new_new_n540_));
  NO3        g518(.A(new_new_n540_), .B(new_new_n525_), .C(new_new_n522_), .Y(new_new_n541_));
  NO2        g519(.A(new_new_n215_), .B(new_new_n104_), .Y(new_new_n542_));
  NO2        g520(.A(new_new_n542_), .B(new_new_n497_), .Y(new_new_n543_));
  NA2        g521(.A(new_new_n543_), .B(i_1_), .Y(new_new_n544_));
  NO2        g522(.A(new_new_n544_), .B(new_new_n491_), .Y(new_new_n545_));
  NO2        g523(.A(new_new_n328_), .B(new_new_n86_), .Y(new_new_n546_));
  NA2        g524(.A(new_new_n545_), .B(new_new_n46_), .Y(new_new_n547_));
  NA2        g525(.A(i_3_), .B(new_new_n180_), .Y(new_new_n548_));
  NO2        g526(.A(new_new_n548_), .B(new_new_n118_), .Y(new_new_n549_));
  AN2        g527(.A(new_new_n549_), .B(new_new_n421_), .Y(new_new_n550_));
  NO2        g528(.A(new_new_n214_), .B(new_new_n44_), .Y(new_new_n551_));
  NO3        g529(.A(new_new_n551_), .B(new_new_n258_), .C(new_new_n216_), .Y(new_new_n552_));
  NO2        g530(.A(new_new_n121_), .B(new_new_n37_), .Y(new_new_n553_));
  NO2        g531(.A(new_new_n553_), .B(i_6_), .Y(new_new_n554_));
  NO2        g532(.A(new_new_n86_), .B(i_9_), .Y(new_new_n555_));
  NO2        g533(.A(new_new_n555_), .B(new_new_n63_), .Y(new_new_n556_));
  NO2        g534(.A(new_new_n556_), .B(new_new_n513_), .Y(new_new_n557_));
  NO4        g535(.A(new_new_n557_), .B(new_new_n554_), .C(new_new_n552_), .D(i_4_), .Y(new_new_n558_));
  NA2        g536(.A(i_1_), .B(i_3_), .Y(new_new_n559_));
  NO2        g537(.A(new_new_n359_), .B(new_new_n95_), .Y(new_new_n560_));
  AOI210     g538(.A0(new_new_n551_), .A1(new_new_n447_), .B0(new_new_n560_), .Y(new_new_n561_));
  NO2        g539(.A(new_new_n561_), .B(new_new_n559_), .Y(new_new_n562_));
  NO3        g540(.A(new_new_n562_), .B(new_new_n558_), .C(new_new_n550_), .Y(new_new_n563_));
  NA4        g541(.A(new_new_n563_), .B(new_new_n547_), .C(new_new_n541_), .D(new_new_n517_), .Y(new_new_n564_));
  AN2        g542(.A(new_new_n222_), .B(new_new_n86_), .Y(new_new_n565_));
  NA2        g543(.A(new_new_n296_), .B(new_new_n295_), .Y(new_new_n566_));
  NA3        g544(.A(new_new_n383_), .B(new_new_n410_), .C(new_new_n46_), .Y(new_new_n567_));
  NO3        g545(.A(new_new_n381_), .B(new_new_n483_), .C(new_new_n86_), .Y(new_new_n568_));
  NA2        g546(.A(new_new_n568_), .B(new_new_n25_), .Y(new_new_n569_));
  NA3        g547(.A(new_new_n161_), .B(new_new_n84_), .C(new_new_n86_), .Y(new_new_n570_));
  NA4        g548(.A(new_new_n570_), .B(new_new_n569_), .C(new_new_n567_), .D(new_new_n566_), .Y(new_new_n571_));
  OAI210     g549(.A0(new_new_n571_), .A1(new_new_n565_), .B0(i_1_), .Y(new_new_n572_));
  AOI210     g550(.A0(new_new_n241_), .A1(new_new_n100_), .B0(i_1_), .Y(new_new_n573_));
  NO2        g551(.A(new_new_n294_), .B(i_2_), .Y(new_new_n574_));
  NA2        g552(.A(new_new_n574_), .B(new_new_n573_), .Y(new_new_n575_));
  AOI210     g553(.A0(new_new_n575_), .A1(new_new_n572_), .B0(i_13_), .Y(new_new_n576_));
  OR2        g554(.A(i_11_), .B(i_7_), .Y(new_new_n577_));
  NA3        g555(.A(new_new_n577_), .B(new_new_n109_), .C(new_new_n142_), .Y(new_new_n578_));
  AOI220     g556(.A0(new_new_n375_), .A1(new_new_n161_), .B0(new_new_n352_), .B1(new_new_n142_), .Y(new_new_n579_));
  OAI210     g557(.A0(new_new_n579_), .A1(new_new_n44_), .B0(new_new_n578_), .Y(new_new_n580_));
  AOI210     g558(.A0(new_new_n529_), .A1(new_new_n54_), .B0(i_12_), .Y(new_new_n581_));
  NO2        g559(.A(new_new_n381_), .B(new_new_n24_), .Y(new_new_n582_));
  AOI220     g560(.A0(new_new_n582_), .A1(new_new_n546_), .B0(new_new_n222_), .B1(new_new_n135_), .Y(new_new_n583_));
  OAI220     g561(.A0(new_new_n583_), .A1(new_new_n41_), .B0(new_new_n893_), .B1(new_new_n95_), .Y(new_new_n584_));
  AOI210     g562(.A0(new_new_n580_), .A1(new_new_n267_), .B0(new_new_n584_), .Y(new_new_n585_));
  INV        g563(.A(new_new_n118_), .Y(new_new_n586_));
  AOI220     g564(.A0(new_new_n586_), .A1(new_new_n72_), .B0(new_new_n312_), .B1(new_new_n530_), .Y(new_new_n587_));
  NO2        g565(.A(new_new_n587_), .B(new_new_n220_), .Y(new_new_n588_));
  AOI210     g566(.A0(new_new_n349_), .A1(new_new_n36_), .B0(i_13_), .Y(new_new_n589_));
  NOi31      g567(.An(new_new_n589_), .B(new_new_n472_), .C(new_new_n44_), .Y(new_new_n590_));
  NA2        g568(.A(new_new_n131_), .B(i_13_), .Y(new_new_n591_));
  NO2        g569(.A(new_new_n529_), .B(new_new_n118_), .Y(new_new_n592_));
  INV        g570(.A(new_new_n592_), .Y(new_new_n593_));
  OAI220     g571(.A0(new_new_n593_), .A1(new_new_n71_), .B0(new_new_n591_), .B1(new_new_n573_), .Y(new_new_n594_));
  NO3        g572(.A(new_new_n71_), .B(new_new_n32_), .C(new_new_n104_), .Y(new_new_n595_));
  NA2        g573(.A(new_new_n26_), .B(new_new_n180_), .Y(new_new_n596_));
  NA2        g574(.A(new_new_n596_), .B(i_7_), .Y(new_new_n597_));
  NO3        g575(.A(new_new_n381_), .B(new_new_n215_), .C(new_new_n86_), .Y(new_new_n598_));
  AOI210     g576(.A0(new_new_n598_), .A1(new_new_n597_), .B0(new_new_n595_), .Y(new_new_n599_));
  AOI220     g577(.A0(new_new_n312_), .A1(new_new_n530_), .B0(new_new_n94_), .B1(new_new_n105_), .Y(new_new_n600_));
  OAI220     g578(.A0(new_new_n600_), .A1(new_new_n478_), .B0(new_new_n599_), .B1(new_new_n493_), .Y(new_new_n601_));
  NO4        g579(.A(new_new_n601_), .B(new_new_n594_), .C(new_new_n590_), .D(new_new_n588_), .Y(new_new_n602_));
  OR2        g580(.A(i_11_), .B(i_6_), .Y(new_new_n603_));
  NA3        g581(.A(new_new_n477_), .B(new_new_n596_), .C(i_7_), .Y(new_new_n604_));
  AOI210     g582(.A0(new_new_n604_), .A1(new_new_n593_), .B0(new_new_n603_), .Y(new_new_n605_));
  NA3        g583(.A(new_new_n327_), .B(new_new_n482_), .C(new_new_n100_), .Y(new_new_n606_));
  NA2        g584(.A(new_new_n521_), .B(i_13_), .Y(new_new_n607_));
  NA2        g585(.A(new_new_n105_), .B(new_new_n596_), .Y(new_new_n608_));
  NAi21      g586(.An(i_11_), .B(i_12_), .Y(new_new_n609_));
  NOi41      g587(.An(new_new_n114_), .B(new_new_n609_), .C(i_13_), .D(new_new_n86_), .Y(new_new_n610_));
  NO3        g588(.A(new_new_n381_), .B(new_new_n457_), .C(new_new_n483_), .Y(new_new_n611_));
  AOI220     g589(.A0(new_new_n611_), .A1(new_new_n260_), .B0(new_new_n610_), .B1(new_new_n608_), .Y(new_new_n612_));
  NA3        g590(.A(new_new_n612_), .B(new_new_n607_), .C(new_new_n606_), .Y(new_new_n613_));
  OAI210     g591(.A0(new_new_n613_), .A1(new_new_n605_), .B0(new_new_n63_), .Y(new_new_n614_));
  NO2        g592(.A(i_2_), .B(i_12_), .Y(new_new_n615_));
  NA2        g593(.A(new_new_n293_), .B(new_new_n615_), .Y(new_new_n616_));
  NA2        g594(.A(i_8_), .B(new_new_n25_), .Y(new_new_n617_));
  NO3        g595(.A(new_new_n617_), .B(new_new_n310_), .C(new_new_n477_), .Y(new_new_n618_));
  OAI210     g596(.A0(new_new_n618_), .A1(new_new_n295_), .B0(new_new_n293_), .Y(new_new_n619_));
  NO2        g597(.A(new_new_n132_), .B(i_2_), .Y(new_new_n620_));
  NA2        g598(.A(new_new_n620_), .B(new_new_n513_), .Y(new_new_n621_));
  NA3        g599(.A(new_new_n621_), .B(new_new_n619_), .C(new_new_n616_), .Y(new_new_n622_));
  NA3        g600(.A(new_new_n622_), .B(new_new_n45_), .C(new_new_n208_), .Y(new_new_n623_));
  NA4        g601(.A(new_new_n623_), .B(new_new_n614_), .C(new_new_n602_), .D(new_new_n585_), .Y(new_new_n624_));
  OR4        g602(.A(new_new_n624_), .B(new_new_n576_), .C(new_new_n564_), .D(new_new_n496_), .Y(ori5));
  NA2        g603(.A(new_new_n543_), .B(new_new_n244_), .Y(new_new_n626_));
  AN2        g604(.A(new_new_n24_), .B(i_10_), .Y(new_new_n627_));
  NA3        g605(.A(new_new_n627_), .B(new_new_n615_), .C(new_new_n111_), .Y(new_new_n628_));
  NO2        g606(.A(new_new_n478_), .B(i_11_), .Y(new_new_n629_));
  NA2        g607(.A(new_new_n89_), .B(new_new_n629_), .Y(new_new_n630_));
  NA3        g608(.A(new_new_n630_), .B(new_new_n628_), .C(new_new_n626_), .Y(new_new_n631_));
  NO3        g609(.A(i_11_), .B(new_new_n215_), .C(i_13_), .Y(new_new_n632_));
  NO2        g610(.A(new_new_n128_), .B(new_new_n23_), .Y(new_new_n633_));
  NA2        g611(.A(i_12_), .B(i_8_), .Y(new_new_n634_));
  OAI210     g612(.A0(new_new_n46_), .A1(i_3_), .B0(new_new_n634_), .Y(new_new_n635_));
  INV        g613(.A(new_new_n348_), .Y(new_new_n636_));
  AOI220     g614(.A0(new_new_n261_), .A1(new_new_n451_), .B0(new_new_n635_), .B1(new_new_n633_), .Y(new_new_n637_));
  INV        g615(.A(new_new_n637_), .Y(new_new_n638_));
  NO2        g616(.A(new_new_n638_), .B(new_new_n631_), .Y(new_new_n639_));
  INV        g617(.A(new_new_n166_), .Y(new_new_n640_));
  INV        g618(.A(new_new_n222_), .Y(new_new_n641_));
  OAI210     g619(.A0(new_new_n574_), .A1(new_new_n350_), .B0(new_new_n114_), .Y(new_new_n642_));
  AOI210     g620(.A0(new_new_n642_), .A1(new_new_n641_), .B0(new_new_n640_), .Y(new_new_n643_));
  NO2        g621(.A(new_new_n359_), .B(new_new_n26_), .Y(new_new_n644_));
  NO2        g622(.A(new_new_n644_), .B(new_new_n332_), .Y(new_new_n645_));
  NA2        g623(.A(new_new_n645_), .B(i_2_), .Y(new_new_n646_));
  INV        g624(.A(new_new_n646_), .Y(new_new_n647_));
  AOI210     g625(.A0(new_new_n33_), .A1(new_new_n36_), .B0(new_new_n329_), .Y(new_new_n648_));
  AOI210     g626(.A0(new_new_n648_), .A1(new_new_n647_), .B0(new_new_n643_), .Y(new_new_n649_));
  NO2        g627(.A(new_new_n179_), .B(new_new_n129_), .Y(new_new_n650_));
  OAI210     g628(.A0(new_new_n650_), .A1(new_new_n633_), .B0(i_2_), .Y(new_new_n651_));
  INV        g629(.A(new_new_n167_), .Y(new_new_n652_));
  NO3        g630(.A(new_new_n498_), .B(new_new_n38_), .C(new_new_n26_), .Y(new_new_n653_));
  AOI210     g631(.A0(new_new_n652_), .A1(new_new_n89_), .B0(new_new_n653_), .Y(new_new_n654_));
  AOI210     g632(.A0(new_new_n654_), .A1(new_new_n651_), .B0(new_new_n180_), .Y(new_new_n655_));
  OA210      g633(.A0(new_new_n499_), .A1(new_new_n130_), .B0(i_13_), .Y(new_new_n656_));
  NA2        g634(.A(new_new_n184_), .B(new_new_n187_), .Y(new_new_n657_));
  NA2        g635(.A(new_new_n155_), .B(new_new_n473_), .Y(new_new_n658_));
  AOI210     g636(.A0(new_new_n658_), .A1(new_new_n657_), .B0(new_new_n298_), .Y(new_new_n659_));
  AOI210     g637(.A0(new_new_n193_), .A1(new_new_n152_), .B0(new_new_n410_), .Y(new_new_n660_));
  NA2        g638(.A(new_new_n660_), .B(new_new_n332_), .Y(new_new_n661_));
  NO2        g639(.A(new_new_n105_), .B(new_new_n44_), .Y(new_new_n662_));
  INV        g640(.A(new_new_n255_), .Y(new_new_n663_));
  NA4        g641(.A(new_new_n663_), .B(new_new_n256_), .C(new_new_n128_), .D(new_new_n42_), .Y(new_new_n664_));
  OAI210     g642(.A0(new_new_n664_), .A1(new_new_n662_), .B0(new_new_n661_), .Y(new_new_n665_));
  NO4        g643(.A(new_new_n665_), .B(new_new_n659_), .C(new_new_n656_), .D(new_new_n655_), .Y(new_new_n666_));
  NA2        g644(.A(new_new_n451_), .B(new_new_n28_), .Y(new_new_n667_));
  NA2        g645(.A(new_new_n632_), .B(new_new_n250_), .Y(new_new_n668_));
  NA2        g646(.A(new_new_n668_), .B(new_new_n667_), .Y(new_new_n669_));
  NO2        g647(.A(new_new_n62_), .B(i_12_), .Y(new_new_n670_));
  NO2        g648(.A(new_new_n670_), .B(new_new_n130_), .Y(new_new_n671_));
  NO2        g649(.A(new_new_n671_), .B(new_new_n473_), .Y(new_new_n672_));
  AOI220     g650(.A0(new_new_n672_), .A1(new_new_n36_), .B0(new_new_n669_), .B1(new_new_n46_), .Y(new_new_n673_));
  NA4        g651(.A(new_new_n673_), .B(new_new_n666_), .C(new_new_n649_), .D(new_new_n639_), .Y(ori6));
  NA4        g652(.A(new_new_n315_), .B(new_new_n382_), .C(new_new_n71_), .D(new_new_n104_), .Y(new_new_n675_));
  INV        g653(.A(new_new_n675_), .Y(new_new_n676_));
  NO2        g654(.A(new_new_n204_), .B(new_new_n385_), .Y(new_new_n677_));
  NO2        g655(.A(i_11_), .B(i_9_), .Y(new_new_n678_));
  NO2        g656(.A(new_new_n676_), .B(new_new_n265_), .Y(new_new_n679_));
  OR2        g657(.A(new_new_n679_), .B(i_12_), .Y(new_new_n680_));
  NA2        g658(.A(new_new_n299_), .B(new_new_n268_), .Y(new_new_n681_));
  NA2        g659(.A(new_new_n457_), .B(new_new_n63_), .Y(new_new_n682_));
  BUFFER     g660(.A(new_new_n504_), .Y(new_new_n683_));
  NA3        g661(.A(new_new_n683_), .B(new_new_n682_), .C(new_new_n681_), .Y(new_new_n684_));
  INV        g662(.A(new_new_n182_), .Y(new_new_n685_));
  AOI220     g663(.A0(new_new_n685_), .A1(new_new_n678_), .B0(new_new_n684_), .B1(new_new_n73_), .Y(new_new_n686_));
  INV        g664(.A(new_new_n264_), .Y(new_new_n687_));
  NA2        g665(.A(new_new_n75_), .B(new_new_n135_), .Y(new_new_n688_));
  INV        g666(.A(new_new_n128_), .Y(new_new_n689_));
  NA2        g667(.A(new_new_n689_), .B(new_new_n46_), .Y(new_new_n690_));
  AOI210     g668(.A0(new_new_n690_), .A1(new_new_n688_), .B0(new_new_n687_), .Y(new_new_n691_));
  NO3        g669(.A(new_new_n226_), .B(new_new_n136_), .C(i_9_), .Y(new_new_n692_));
  NA2        g670(.A(new_new_n692_), .B(new_new_n670_), .Y(new_new_n693_));
  AOI210     g671(.A0(new_new_n693_), .A1(new_new_n408_), .B0(new_new_n174_), .Y(new_new_n694_));
  NO2        g672(.A(new_new_n32_), .B(i_11_), .Y(new_new_n695_));
  NAi32      g673(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(new_new_n696_));
  NO2        g674(.A(new_new_n603_), .B(new_new_n696_), .Y(new_new_n697_));
  OR3        g675(.A(new_new_n697_), .B(new_new_n694_), .C(new_new_n691_), .Y(new_new_n698_));
  NO2        g676(.A(new_new_n577_), .B(i_2_), .Y(new_new_n699_));
  NA2        g677(.A(new_new_n48_), .B(new_new_n37_), .Y(new_new_n700_));
  NO2        g678(.A(new_new_n700_), .B(new_new_n326_), .Y(new_new_n701_));
  NA2        g679(.A(new_new_n701_), .B(new_new_n699_), .Y(new_new_n702_));
  OR2        g680(.A(new_new_n499_), .B(new_new_n350_), .Y(new_new_n703_));
  NA3        g681(.A(new_new_n703_), .B(new_new_n151_), .C(new_new_n69_), .Y(new_new_n704_));
  AO210      g682(.A0(new_new_n392_), .A1(new_new_n636_), .B0(new_new_n36_), .Y(new_new_n705_));
  NA3        g683(.A(new_new_n705_), .B(new_new_n704_), .C(new_new_n702_), .Y(new_new_n706_));
  OAI210     g684(.A0(new_new_n520_), .A1(i_11_), .B0(new_new_n87_), .Y(new_new_n707_));
  AOI220     g685(.A0(new_new_n707_), .A1(new_new_n444_), .B0(new_new_n677_), .B1(new_new_n597_), .Y(new_new_n708_));
  NA3        g686(.A(new_new_n298_), .B(new_new_n217_), .C(new_new_n151_), .Y(new_new_n709_));
  NA2        g687(.A(new_new_n319_), .B(new_new_n70_), .Y(new_new_n710_));
  NA4        g688(.A(new_new_n710_), .B(new_new_n709_), .C(new_new_n708_), .D(new_new_n481_), .Y(new_new_n711_));
  AO210      g689(.A0(new_new_n410_), .A1(new_new_n46_), .B0(new_new_n88_), .Y(new_new_n712_));
  NA3        g690(.A(new_new_n712_), .B(new_new_n383_), .C(new_new_n201_), .Y(new_new_n713_));
  AOI210     g691(.A0(new_new_n350_), .A1(new_new_n348_), .B0(new_new_n443_), .Y(new_new_n714_));
  NO2        g692(.A(new_new_n489_), .B(new_new_n105_), .Y(new_new_n715_));
  OAI210     g693(.A0(new_new_n715_), .A1(new_new_n115_), .B0(new_new_n325_), .Y(new_new_n716_));
  NA2        g694(.A(new_new_n221_), .B(new_new_n46_), .Y(new_new_n717_));
  INV        g695(.A(new_new_n462_), .Y(new_new_n718_));
  NA3        g696(.A(new_new_n718_), .B(new_new_n264_), .C(i_7_), .Y(new_new_n719_));
  NA4        g697(.A(new_new_n719_), .B(new_new_n716_), .C(new_new_n714_), .D(new_new_n713_), .Y(new_new_n720_));
  NO4        g698(.A(new_new_n720_), .B(new_new_n711_), .C(new_new_n706_), .D(new_new_n698_), .Y(new_new_n721_));
  NA4        g699(.A(new_new_n721_), .B(new_new_n686_), .C(new_new_n680_), .D(new_new_n306_), .Y(ori3));
  NA2        g700(.A(i_12_), .B(i_10_), .Y(new_new_n723_));
  NO2        g701(.A(i_11_), .B(new_new_n215_), .Y(new_new_n724_));
  NA3        g702(.A(new_new_n709_), .B(new_new_n481_), .C(new_new_n297_), .Y(new_new_n725_));
  NA2        g703(.A(new_new_n725_), .B(new_new_n40_), .Y(new_new_n726_));
  NOi21      g704(.An(new_new_n99_), .B(new_new_n645_), .Y(new_new_n727_));
  NO3        g705(.A(new_new_n509_), .B(new_new_n359_), .C(new_new_n135_), .Y(new_new_n728_));
  NA2        g706(.A(new_new_n327_), .B(new_new_n45_), .Y(new_new_n729_));
  AN2        g707(.A(new_new_n357_), .B(new_new_n55_), .Y(new_new_n730_));
  NO3        g708(.A(new_new_n730_), .B(new_new_n728_), .C(new_new_n727_), .Y(new_new_n731_));
  AOI210     g709(.A0(new_new_n731_), .A1(new_new_n726_), .B0(new_new_n48_), .Y(new_new_n732_));
  NO4        g710(.A(new_new_n302_), .B(new_new_n309_), .C(new_new_n38_), .D(i_0_), .Y(new_new_n733_));
  NA2        g711(.A(new_new_n174_), .B(new_new_n447_), .Y(new_new_n734_));
  NOi21      g712(.An(new_new_n734_), .B(new_new_n733_), .Y(new_new_n735_));
  NO2        g713(.A(new_new_n735_), .B(new_new_n63_), .Y(new_new_n736_));
  NOi21      g714(.An(i_5_), .B(i_9_), .Y(new_new_n737_));
  NA2        g715(.A(new_new_n737_), .B(new_new_n346_), .Y(new_new_n738_));
  BUFFER     g716(.A(new_new_n241_), .Y(new_new_n739_));
  AOI210     g717(.A0(new_new_n739_), .A1(new_new_n379_), .B0(new_new_n568_), .Y(new_new_n740_));
  NO2        g718(.A(new_new_n740_), .B(new_new_n738_), .Y(new_new_n741_));
  NO3        g719(.A(new_new_n741_), .B(new_new_n736_), .C(new_new_n732_), .Y(new_new_n742_));
  NA2        g720(.A(new_new_n174_), .B(new_new_n24_), .Y(new_new_n743_));
  NO2        g721(.A(new_new_n553_), .B(new_new_n470_), .Y(new_new_n744_));
  NO2        g722(.A(new_new_n744_), .B(new_new_n743_), .Y(new_new_n745_));
  NAi21      g723(.An(new_new_n162_), .B(new_new_n341_), .Y(new_new_n746_));
  NO2        g724(.A(new_new_n746_), .B(new_new_n717_), .Y(new_new_n747_));
  NO2        g725(.A(new_new_n747_), .B(new_new_n745_), .Y(new_new_n748_));
  NA2        g726(.A(new_new_n448_), .B(i_0_), .Y(new_new_n749_));
  NO3        g727(.A(new_new_n749_), .B(new_new_n311_), .C(new_new_n89_), .Y(new_new_n750_));
  NO4        g728(.A(new_new_n461_), .B(new_new_n198_), .C(new_new_n329_), .D(new_new_n326_), .Y(new_new_n751_));
  AOI210     g729(.A0(new_new_n751_), .A1(i_11_), .B0(new_new_n750_), .Y(new_new_n752_));
  INV        g730(.A(new_new_n378_), .Y(new_new_n753_));
  NA2        g731(.A(new_new_n632_), .B(new_new_n265_), .Y(new_new_n754_));
  AOI210     g732(.A0(new_new_n383_), .A1(new_new_n89_), .B0(new_new_n58_), .Y(new_new_n755_));
  NO2        g733(.A(new_new_n755_), .B(new_new_n754_), .Y(new_new_n756_));
  NO2        g734(.A(new_new_n228_), .B(new_new_n156_), .Y(new_new_n757_));
  NA2        g735(.A(i_0_), .B(i_10_), .Y(new_new_n758_));
  INV        g736(.A(new_new_n420_), .Y(new_new_n759_));
  NO4        g737(.A(new_new_n118_), .B(new_new_n58_), .C(new_new_n548_), .D(i_5_), .Y(new_new_n760_));
  AO220      g738(.A0(new_new_n760_), .A1(new_new_n759_), .B0(new_new_n757_), .B1(i_6_), .Y(new_new_n761_));
  NO2        g739(.A(new_new_n761_), .B(new_new_n756_), .Y(new_new_n762_));
  NA3        g740(.A(new_new_n762_), .B(new_new_n752_), .C(new_new_n748_), .Y(new_new_n763_));
  NO2        g741(.A(new_new_n106_), .B(new_new_n37_), .Y(new_new_n764_));
  NA2        g742(.A(i_11_), .B(i_9_), .Y(new_new_n765_));
  NO3        g743(.A(i_12_), .B(new_new_n765_), .C(new_new_n480_), .Y(new_new_n766_));
  AN2        g744(.A(new_new_n766_), .B(new_new_n764_), .Y(new_new_n767_));
  NO2        g745(.A(new_new_n48_), .B(i_7_), .Y(new_new_n768_));
  NA2        g746(.A(new_new_n316_), .B(new_new_n171_), .Y(new_new_n769_));
  NA2        g747(.A(new_new_n769_), .B(new_new_n160_), .Y(new_new_n770_));
  NO2        g748(.A(new_new_n765_), .B(new_new_n73_), .Y(new_new_n771_));
  NO2        g749(.A(new_new_n169_), .B(i_0_), .Y(new_new_n772_));
  INV        g750(.A(new_new_n324_), .Y(new_new_n773_));
  NO2        g751(.A(new_new_n773_), .B(new_new_n738_), .Y(new_new_n774_));
  NO3        g752(.A(new_new_n774_), .B(new_new_n770_), .C(new_new_n767_), .Y(new_new_n775_));
  NA2        g753(.A(new_new_n537_), .B(new_new_n125_), .Y(new_new_n776_));
  NO2        g754(.A(i_6_), .B(new_new_n776_), .Y(new_new_n777_));
  AOI210     g755(.A0(new_new_n349_), .A1(new_new_n36_), .B0(i_3_), .Y(new_new_n778_));
  NA2        g756(.A(new_new_n166_), .B(new_new_n106_), .Y(new_new_n779_));
  NOi32      g757(.An(new_new_n778_), .Bn(new_new_n177_), .C(new_new_n779_), .Y(new_new_n780_));
  NA2        g758(.A(new_new_n482_), .B(new_new_n265_), .Y(new_new_n781_));
  NO2        g759(.A(new_new_n781_), .B(new_new_n729_), .Y(new_new_n782_));
  NO3        g760(.A(new_new_n782_), .B(new_new_n780_), .C(new_new_n777_), .Y(new_new_n783_));
  NOi21      g761(.An(i_7_), .B(i_5_), .Y(new_new_n784_));
  NOi31      g762(.An(new_new_n784_), .B(i_0_), .C(new_new_n609_), .Y(new_new_n785_));
  NA3        g763(.A(new_new_n785_), .B(new_new_n310_), .C(i_6_), .Y(new_new_n786_));
  BUFFER     g764(.A(new_new_n786_), .Y(new_new_n787_));
  INV        g765(.A(new_new_n262_), .Y(new_new_n788_));
  NA3        g766(.A(new_new_n787_), .B(new_new_n783_), .C(new_new_n775_), .Y(new_new_n789_));
  NO2        g767(.A(new_new_n723_), .B(new_new_n261_), .Y(new_new_n790_));
  OA210      g768(.A0(new_new_n378_), .A1(new_new_n207_), .B0(new_new_n377_), .Y(new_new_n791_));
  NA2        g769(.A(new_new_n790_), .B(new_new_n771_), .Y(new_new_n792_));
  NA3        g770(.A(new_new_n377_), .B(new_new_n327_), .C(new_new_n45_), .Y(new_new_n793_));
  OAI210     g771(.A0(new_new_n746_), .A1(new_new_n753_), .B0(new_new_n793_), .Y(new_new_n794_));
  NA2        g772(.A(new_new_n771_), .B(new_new_n256_), .Y(new_new_n795_));
  OAI210     g773(.A0(i_2_), .A1(new_new_n176_), .B0(new_new_n795_), .Y(new_new_n796_));
  AOI220     g774(.A0(new_new_n796_), .A1(new_new_n378_), .B0(new_new_n794_), .B1(new_new_n73_), .Y(new_new_n797_));
  NA3        g775(.A(new_new_n700_), .B(new_new_n308_), .C(new_new_n520_), .Y(new_new_n798_));
  NO2        g776(.A(new_new_n75_), .B(new_new_n634_), .Y(new_new_n799_));
  AOI220     g777(.A0(new_new_n799_), .A1(i_11_), .B0(new_new_n168_), .B1(new_new_n470_), .Y(new_new_n800_));
  AOI210     g778(.A0(new_new_n800_), .A1(new_new_n798_), .B0(new_new_n47_), .Y(new_new_n801_));
  NO3        g779(.A(new_new_n461_), .B(new_new_n280_), .C(new_new_n24_), .Y(new_new_n802_));
  AOI210     g780(.A0(new_new_n582_), .A1(new_new_n427_), .B0(new_new_n802_), .Y(new_new_n803_));
  NAi21      g781(.An(i_9_), .B(i_5_), .Y(new_new_n804_));
  NO2        g782(.A(new_new_n804_), .B(new_new_n321_), .Y(new_new_n805_));
  NA2        g783(.A(new_new_n805_), .B(new_new_n499_), .Y(new_new_n806_));
  OAI220     g784(.A0(new_new_n806_), .A1(new_new_n86_), .B0(new_new_n803_), .B1(new_new_n167_), .Y(new_new_n807_));
  NO3        g785(.A(new_new_n807_), .B(new_new_n801_), .C(new_new_n412_), .Y(new_new_n808_));
  NA3        g786(.A(new_new_n808_), .B(new_new_n797_), .C(new_new_n792_), .Y(new_new_n809_));
  NO3        g787(.A(new_new_n809_), .B(new_new_n789_), .C(new_new_n763_), .Y(new_new_n810_));
  NO2        g788(.A(i_0_), .B(new_new_n609_), .Y(new_new_n811_));
  AOI210     g789(.A0(new_new_n682_), .A1(new_new_n566_), .B0(new_new_n779_), .Y(new_new_n812_));
  INV        g790(.A(new_new_n812_), .Y(new_new_n813_));
  OAI210     g791(.A0(new_new_n221_), .A1(i_9_), .B0(new_new_n213_), .Y(new_new_n814_));
  AOI210     g792(.A0(new_new_n814_), .A1(new_new_n749_), .B0(new_new_n156_), .Y(new_new_n815_));
  INV        g793(.A(new_new_n815_), .Y(new_new_n816_));
  NA2        g794(.A(new_new_n816_), .B(new_new_n813_), .Y(new_new_n817_));
  NO3        g795(.A(new_new_n758_), .B(new_new_n737_), .C(new_new_n179_), .Y(new_new_n818_));
  AOI220     g796(.A0(new_new_n818_), .A1(i_11_), .B0(new_new_n446_), .B1(new_new_n75_), .Y(new_new_n819_));
  NO3        g797(.A(new_new_n194_), .B(new_new_n309_), .C(i_0_), .Y(new_new_n820_));
  OAI210     g798(.A0(new_new_n820_), .A1(new_new_n76_), .B0(i_13_), .Y(new_new_n821_));
  NA2        g799(.A(new_new_n821_), .B(new_new_n819_), .Y(new_new_n822_));
  NO2        g800(.A(new_new_n220_), .B(new_new_n95_), .Y(new_new_n823_));
  AOI210     g801(.A0(new_new_n823_), .A1(new_new_n811_), .B0(new_new_n112_), .Y(new_new_n824_));
  OR2        g802(.A(new_new_n824_), .B(i_5_), .Y(new_new_n825_));
  AOI210     g803(.A0(i_0_), .A1(new_new_n25_), .B0(new_new_n169_), .Y(new_new_n826_));
  NA2        g804(.A(new_new_n826_), .B(new_new_n791_), .Y(new_new_n827_));
  INV        g805(.A(new_new_n425_), .Y(new_new_n828_));
  NO3        g806(.A(new_new_n729_), .B(new_new_n54_), .C(new_new_n48_), .Y(new_new_n829_));
  NA2        g807(.A(new_new_n391_), .B(new_new_n384_), .Y(new_new_n830_));
  NO3        g808(.A(new_new_n830_), .B(new_new_n829_), .C(new_new_n828_), .Y(new_new_n831_));
  NA3        g809(.A(new_new_n315_), .B(new_new_n166_), .C(new_new_n165_), .Y(new_new_n832_));
  NA3        g810(.A(new_new_n768_), .B(new_new_n254_), .C(new_new_n213_), .Y(new_new_n833_));
  NA2        g811(.A(new_new_n833_), .B(new_new_n832_), .Y(new_new_n834_));
  NO3        g812(.A(new_new_n765_), .B(new_new_n201_), .C(new_new_n179_), .Y(new_new_n835_));
  NO2        g813(.A(new_new_n835_), .B(new_new_n834_), .Y(new_new_n836_));
  NA4        g814(.A(new_new_n836_), .B(new_new_n831_), .C(new_new_n827_), .D(new_new_n825_), .Y(new_new_n837_));
  NO2        g815(.A(new_new_n86_), .B(i_5_), .Y(new_new_n838_));
  NA3        g816(.A(new_new_n724_), .B(new_new_n113_), .C(new_new_n128_), .Y(new_new_n839_));
  INV        g817(.A(new_new_n839_), .Y(new_new_n840_));
  NA2        g818(.A(new_new_n840_), .B(new_new_n838_), .Y(new_new_n841_));
  NA3        g819(.A(new_new_n256_), .B(i_5_), .C(new_new_n180_), .Y(new_new_n842_));
  NAi31      g820(.An(new_new_n219_), .B(new_new_n842_), .C(new_new_n220_), .Y(new_new_n843_));
  NO4        g821(.A(new_new_n218_), .B(new_new_n194_), .C(i_0_), .D(i_12_), .Y(new_new_n844_));
  AOI220     g822(.A0(new_new_n844_), .A1(new_new_n843_), .B0(new_new_n676_), .B1(new_new_n170_), .Y(new_new_n845_));
  NA2        g823(.A(new_new_n784_), .B(new_new_n375_), .Y(new_new_n846_));
  NA2        g824(.A(new_new_n64_), .B(new_new_n104_), .Y(new_new_n847_));
  OAI220     g825(.A0(new_new_n847_), .A1(new_new_n842_), .B0(new_new_n846_), .B1(new_new_n556_), .Y(new_new_n848_));
  NA2        g826(.A(new_new_n848_), .B(new_new_n772_), .Y(new_new_n849_));
  NA3        g827(.A(new_new_n849_), .B(new_new_n845_), .C(new_new_n841_), .Y(new_new_n850_));
  NO4        g828(.A(new_new_n850_), .B(new_new_n837_), .C(new_new_n822_), .D(new_new_n817_), .Y(new_new_n851_));
  OAI210     g829(.A0(new_new_n699_), .A1(new_new_n695_), .B0(new_new_n37_), .Y(new_new_n852_));
  NA2        g830(.A(new_new_n852_), .B(new_new_n488_), .Y(new_new_n853_));
  NA2        g831(.A(new_new_n853_), .B(new_new_n192_), .Y(new_new_n854_));
  NA2        g832(.A(new_new_n175_), .B(new_new_n177_), .Y(new_new_n855_));
  AO210      g833(.A0(new_new_n577_), .A1(new_new_n33_), .B0(new_new_n855_), .Y(new_new_n856_));
  NAi31      g834(.An(i_7_), .B(i_2_), .C(i_10_), .Y(new_new_n857_));
  AOI210     g835(.A0(new_new_n121_), .A1(new_new_n70_), .B0(new_new_n857_), .Y(new_new_n858_));
  NO2        g836(.A(new_new_n858_), .B(new_new_n523_), .Y(new_new_n859_));
  NA2        g837(.A(new_new_n859_), .B(new_new_n856_), .Y(new_new_n860_));
  NO2        g838(.A(new_new_n367_), .B(new_new_n241_), .Y(new_new_n861_));
  NO2        g839(.A(new_new_n861_), .B(new_new_n751_), .Y(new_new_n862_));
  INV        g840(.A(new_new_n862_), .Y(new_new_n863_));
  AOI210     g841(.A0(new_new_n860_), .A1(new_new_n48_), .B0(new_new_n863_), .Y(new_new_n864_));
  AOI210     g842(.A0(new_new_n864_), .A1(new_new_n854_), .B0(new_new_n73_), .Y(new_new_n865_));
  INV        g843(.A(new_new_n305_), .Y(new_new_n866_));
  NO2        g844(.A(new_new_n866_), .B(new_new_n640_), .Y(new_new_n867_));
  OAI210     g845(.A0(new_new_n80_), .A1(new_new_n54_), .B0(new_new_n111_), .Y(new_new_n868_));
  NA2        g846(.A(new_new_n868_), .B(new_new_n76_), .Y(new_new_n869_));
  AOI210     g847(.A0(new_new_n826_), .A1(new_new_n768_), .B0(new_new_n785_), .Y(new_new_n870_));
  AOI210     g848(.A0(new_new_n870_), .A1(new_new_n869_), .B0(new_new_n559_), .Y(new_new_n871_));
  INV        g849(.A(new_new_n871_), .Y(new_new_n872_));
  OAI210     g850(.A0(new_new_n243_), .A1(new_new_n158_), .B0(new_new_n89_), .Y(new_new_n873_));
  NA3        g851(.A(new_new_n644_), .B(new_new_n254_), .C(new_new_n80_), .Y(new_new_n874_));
  AOI210     g852(.A0(new_new_n874_), .A1(new_new_n873_), .B0(i_11_), .Y(new_new_n875_));
  NA2        g853(.A(new_new_n483_), .B(new_new_n198_), .Y(new_new_n876_));
  OAI210     g854(.A0(new_new_n876_), .A1(new_new_n778_), .B0(new_new_n192_), .Y(new_new_n877_));
  NA2        g855(.A(new_new_n163_), .B(i_5_), .Y(new_new_n878_));
  NO2        g856(.A(new_new_n877_), .B(new_new_n878_), .Y(new_new_n879_));
  NO3        g857(.A(new_new_n59_), .B(new_new_n58_), .C(i_4_), .Y(new_new_n880_));
  OAI210     g858(.A0(new_new_n788_), .A1(new_new_n257_), .B0(new_new_n880_), .Y(new_new_n881_));
  NO2        g859(.A(new_new_n881_), .B(new_new_n609_), .Y(new_new_n882_));
  NO4        g860(.A(new_new_n804_), .B(new_new_n380_), .C(new_new_n227_), .D(new_new_n226_), .Y(new_new_n883_));
  NO2        g861(.A(new_new_n883_), .B(new_new_n443_), .Y(new_new_n884_));
  INV        g862(.A(new_new_n286_), .Y(new_new_n885_));
  AOI210     g863(.A0(new_new_n885_), .A1(new_new_n884_), .B0(new_new_n41_), .Y(new_new_n886_));
  NO4        g864(.A(new_new_n886_), .B(new_new_n882_), .C(new_new_n879_), .D(new_new_n875_), .Y(new_new_n887_));
  OAI210     g865(.A0(new_new_n872_), .A1(i_4_), .B0(new_new_n887_), .Y(new_new_n888_));
  NO3        g866(.A(new_new_n888_), .B(new_new_n867_), .C(new_new_n865_), .Y(new_new_n889_));
  NA4        g867(.A(new_new_n889_), .B(new_new_n851_), .C(new_new_n810_), .D(new_new_n742_), .Y(ori4));
  INV        g868(.A(new_new_n581_), .Y(new_new_n893_));
endmodule


