//Benchmark atmr_alu4_1266_0.5

module atmr_alu4(i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, z0, z1, z2, z3, z4, z5, z6, z7);
 input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_;
 output z0, z1, z2, z3, z4, z5, z6, z7;
 wire ori_ori_n23_, ori_ori_n24_, ori_ori_n25_, ori_ori_n26_, ori_ori_n27_, ori_ori_n28_, ori_ori_n29_, ori_ori_n30_, ori_ori_n31_, ori_ori_n32_, ori_ori_n33_, ori_ori_n34_, ori_ori_n35_, ori_ori_n36_, ori_ori_n37_, ori_ori_n38_, ori_ori_n39_, ori_ori_n40_, ori_ori_n42_, ori_ori_n43_, ori_ori_n44_, ori_ori_n45_, ori_ori_n46_, ori_ori_n47_, ori_ori_n48_, ori_ori_n49_, ori_ori_n50_, ori_ori_n51_, ori_ori_n52_, ori_ori_n53_, ori_ori_n54_, ori_ori_n55_, ori_ori_n56_, ori_ori_n57_, ori_ori_n58_, ori_ori_n59_, ori_ori_n60_, ori_ori_n61_, ori_ori_n62_, ori_ori_n63_, ori_ori_n64_, ori_ori_n65_, ori_ori_n66_, ori_ori_n67_, ori_ori_n68_, ori_ori_n69_, ori_ori_n70_, ori_ori_n71_, ori_ori_n72_, ori_ori_n73_, ori_ori_n74_, ori_ori_n75_, ori_ori_n76_, ori_ori_n77_, ori_ori_n78_, ori_ori_n79_, ori_ori_n80_, ori_ori_n81_, ori_ori_n82_, ori_ori_n83_, ori_ori_n84_, ori_ori_n85_, ori_ori_n86_, ori_ori_n87_, ori_ori_n88_, ori_ori_n89_, ori_ori_n90_, ori_ori_n91_, ori_ori_n92_, ori_ori_n93_, ori_ori_n94_, ori_ori_n95_, ori_ori_n96_, ori_ori_n97_, ori_ori_n98_, ori_ori_n99_, ori_ori_n100_, ori_ori_n101_, ori_ori_n102_, ori_ori_n103_, ori_ori_n104_, ori_ori_n105_, ori_ori_n106_, ori_ori_n108_, ori_ori_n109_, ori_ori_n110_, ori_ori_n112_, ori_ori_n113_, ori_ori_n114_, ori_ori_n115_, ori_ori_n116_, ori_ori_n117_, ori_ori_n118_, ori_ori_n119_, ori_ori_n120_, ori_ori_n121_, ori_ori_n122_, ori_ori_n123_, ori_ori_n124_, ori_ori_n125_, ori_ori_n126_, ori_ori_n127_, ori_ori_n128_, ori_ori_n129_, ori_ori_n130_, ori_ori_n131_, ori_ori_n132_, ori_ori_n133_, ori_ori_n134_, ori_ori_n135_, ori_ori_n136_, ori_ori_n137_, ori_ori_n138_, ori_ori_n139_, ori_ori_n140_, ori_ori_n141_, ori_ori_n142_, ori_ori_n143_, ori_ori_n144_, ori_ori_n145_, ori_ori_n146_, ori_ori_n147_, ori_ori_n148_, ori_ori_n149_, ori_ori_n150_, ori_ori_n151_, ori_ori_n152_, ori_ori_n153_, ori_ori_n154_, ori_ori_n155_, ori_ori_n156_, ori_ori_n157_, ori_ori_n158_, ori_ori_n159_, ori_ori_n160_, ori_ori_n161_, ori_ori_n162_, ori_ori_n163_, ori_ori_n164_, ori_ori_n165_, ori_ori_n166_, ori_ori_n167_, ori_ori_n168_, ori_ori_n169_, ori_ori_n170_, ori_ori_n171_, ori_ori_n172_, ori_ori_n173_, ori_ori_n174_, ori_ori_n175_, ori_ori_n176_, ori_ori_n177_, ori_ori_n178_, ori_ori_n179_, ori_ori_n180_, ori_ori_n181_, ori_ori_n182_, ori_ori_n183_, ori_ori_n184_, ori_ori_n185_, ori_ori_n186_, ori_ori_n187_, ori_ori_n188_, ori_ori_n189_, ori_ori_n190_, ori_ori_n191_, ori_ori_n192_, ori_ori_n193_, ori_ori_n194_, ori_ori_n195_, ori_ori_n196_, ori_ori_n197_, ori_ori_n198_, ori_ori_n199_, ori_ori_n200_, ori_ori_n201_, ori_ori_n202_, ori_ori_n203_, ori_ori_n204_, ori_ori_n205_, ori_ori_n206_, ori_ori_n207_, ori_ori_n208_, ori_ori_n209_, ori_ori_n210_, ori_ori_n211_, ori_ori_n212_, ori_ori_n213_, ori_ori_n214_, ori_ori_n215_, ori_ori_n216_, ori_ori_n217_, ori_ori_n218_, ori_ori_n219_, ori_ori_n220_, ori_ori_n221_, ori_ori_n222_, ori_ori_n223_, ori_ori_n224_, ori_ori_n225_, ori_ori_n226_, ori_ori_n227_, ori_ori_n228_, ori_ori_n229_, ori_ori_n230_, ori_ori_n231_, ori_ori_n232_, ori_ori_n233_, ori_ori_n234_, ori_ori_n235_, ori_ori_n236_, ori_ori_n237_, ori_ori_n238_, ori_ori_n239_, ori_ori_n240_, ori_ori_n241_, ori_ori_n242_, ori_ori_n243_, ori_ori_n244_, ori_ori_n245_, ori_ori_n246_, ori_ori_n247_, ori_ori_n248_, ori_ori_n249_, ori_ori_n250_, ori_ori_n251_, ori_ori_n252_, ori_ori_n253_, ori_ori_n254_, ori_ori_n255_, ori_ori_n256_, ori_ori_n258_, ori_ori_n259_, ori_ori_n260_, ori_ori_n261_, ori_ori_n262_, ori_ori_n263_, ori_ori_n264_, ori_ori_n265_, ori_ori_n266_, ori_ori_n267_, ori_ori_n268_, ori_ori_n269_, ori_ori_n270_, ori_ori_n271_, ori_ori_n272_, ori_ori_n273_, ori_ori_n274_, ori_ori_n275_, ori_ori_n276_, ori_ori_n277_, ori_ori_n278_, ori_ori_n279_, ori_ori_n280_, ori_ori_n281_, ori_ori_n282_, ori_ori_n283_, ori_ori_n284_, ori_ori_n285_, ori_ori_n286_, ori_ori_n287_, ori_ori_n288_, ori_ori_n289_, ori_ori_n290_, ori_ori_n291_, ori_ori_n292_, ori_ori_n293_, ori_ori_n294_, ori_ori_n295_, ori_ori_n296_, ori_ori_n297_, ori_ori_n298_, ori_ori_n299_, ori_ori_n300_, ori_ori_n301_, ori_ori_n302_, ori_ori_n303_, ori_ori_n304_, ori_ori_n305_, ori_ori_n306_, ori_ori_n307_, ori_ori_n308_, ori_ori_n309_, ori_ori_n310_, ori_ori_n311_, ori_ori_n312_, ori_ori_n313_, ori_ori_n314_, ori_ori_n315_, ori_ori_n316_, ori_ori_n317_, ori_ori_n318_, ori_ori_n319_, ori_ori_n320_, ori_ori_n321_, ori_ori_n322_, ori_ori_n323_, ori_ori_n324_, ori_ori_n325_, ori_ori_n326_, ori_ori_n327_, ori_ori_n328_, ori_ori_n329_, ori_ori_n330_, ori_ori_n331_, ori_ori_n332_, ori_ori_n333_, ori_ori_n334_, ori_ori_n335_, ori_ori_n337_, ori_ori_n338_, ori_ori_n339_, ori_ori_n340_, ori_ori_n341_, ori_ori_n342_, ori_ori_n343_, ori_ori_n344_, ori_ori_n345_, ori_ori_n346_, ori_ori_n347_, ori_ori_n348_, ori_ori_n349_, ori_ori_n350_, ori_ori_n351_, ori_ori_n352_, ori_ori_n353_, ori_ori_n354_, ori_ori_n355_, ori_ori_n357_, ori_ori_n358_, ori_ori_n359_, ori_ori_n360_, ori_ori_n361_, ori_ori_n362_, ori_ori_n363_, ori_ori_n364_, ori_ori_n365_, ori_ori_n366_, ori_ori_n367_, ori_ori_n368_, ori_ori_n369_, ori_ori_n370_, ori_ori_n371_, ori_ori_n372_, ori_ori_n373_, ori_ori_n374_, ori_ori_n375_, ori_ori_n376_, ori_ori_n377_, ori_ori_n378_, ori_ori_n380_, ori_ori_n381_, ori_ori_n382_, ori_ori_n383_, ori_ori_n384_, ori_ori_n385_, ori_ori_n386_, ori_ori_n387_, ori_ori_n388_, ori_ori_n389_, ori_ori_n390_, ori_ori_n391_, ori_ori_n392_, ori_ori_n393_, ori_ori_n394_, ori_ori_n395_, ori_ori_n396_, ori_ori_n397_, ori_ori_n398_, ori_ori_n399_, ori_ori_n400_, ori_ori_n401_, ori_ori_n402_, ori_ori_n403_, ori_ori_n404_, ori_ori_n405_, ori_ori_n406_, ori_ori_n407_, ori_ori_n408_, ori_ori_n409_, ori_ori_n410_, ori_ori_n411_, ori_ori_n412_, ori_ori_n413_, ori_ori_n414_, ori_ori_n415_, ori_ori_n416_, ori_ori_n417_, ori_ori_n418_, ori_ori_n419_, ori_ori_n420_, ori_ori_n421_, ori_ori_n422_, ori_ori_n423_, ori_ori_n424_, ori_ori_n425_, ori_ori_n426_, ori_ori_n427_, ori_ori_n428_, ori_ori_n429_, ori_ori_n430_, ori_ori_n431_, ori_ori_n432_, ori_ori_n433_, ori_ori_n434_, ori_ori_n435_, ori_ori_n436_, ori_ori_n437_, ori_ori_n438_, ori_ori_n439_, ori_ori_n440_, ori_ori_n441_, ori_ori_n442_, ori_ori_n443_, ori_ori_n444_, ori_ori_n445_, ori_ori_n446_, ori_ori_n447_, ori_ori_n448_, ori_ori_n452_, ori_ori_n453_, ori_ori_n454_, mai_mai_n23_, mai_mai_n24_, mai_mai_n25_, mai_mai_n26_, mai_mai_n27_, mai_mai_n28_, mai_mai_n29_, mai_mai_n30_, mai_mai_n31_, mai_mai_n32_, mai_mai_n33_, mai_mai_n34_, mai_mai_n35_, mai_mai_n36_, mai_mai_n37_, mai_mai_n38_, mai_mai_n39_, mai_mai_n40_, mai_mai_n41_, mai_mai_n42_, mai_mai_n44_, mai_mai_n45_, mai_mai_n46_, mai_mai_n47_, mai_mai_n48_, mai_mai_n49_, mai_mai_n50_, mai_mai_n51_, mai_mai_n52_, mai_mai_n53_, mai_mai_n54_, mai_mai_n55_, mai_mai_n56_, mai_mai_n57_, mai_mai_n58_, mai_mai_n59_, mai_mai_n60_, mai_mai_n61_, mai_mai_n62_, mai_mai_n63_, mai_mai_n64_, mai_mai_n65_, mai_mai_n66_, mai_mai_n67_, mai_mai_n68_, mai_mai_n69_, mai_mai_n70_, mai_mai_n71_, mai_mai_n72_, mai_mai_n73_, mai_mai_n74_, mai_mai_n75_, mai_mai_n76_, mai_mai_n77_, mai_mai_n78_, mai_mai_n79_, mai_mai_n80_, mai_mai_n81_, mai_mai_n82_, mai_mai_n83_, mai_mai_n84_, mai_mai_n85_, mai_mai_n86_, mai_mai_n87_, mai_mai_n88_, mai_mai_n89_, mai_mai_n90_, mai_mai_n91_, mai_mai_n92_, mai_mai_n93_, mai_mai_n94_, mai_mai_n95_, mai_mai_n96_, mai_mai_n97_, mai_mai_n98_, mai_mai_n99_, mai_mai_n100_, mai_mai_n101_, mai_mai_n102_, mai_mai_n103_, mai_mai_n104_, mai_mai_n105_, mai_mai_n106_, mai_mai_n107_, mai_mai_n108_, mai_mai_n109_, mai_mai_n110_, mai_mai_n111_, mai_mai_n112_, mai_mai_n113_, mai_mai_n114_, mai_mai_n115_, mai_mai_n116_, mai_mai_n117_, mai_mai_n118_, mai_mai_n119_, mai_mai_n120_, mai_mai_n121_, mai_mai_n122_, mai_mai_n123_, mai_mai_n124_, mai_mai_n126_, mai_mai_n127_, mai_mai_n128_, mai_mai_n130_, mai_mai_n131_, mai_mai_n132_, mai_mai_n133_, mai_mai_n134_, mai_mai_n135_, mai_mai_n136_, mai_mai_n137_, mai_mai_n138_, mai_mai_n139_, mai_mai_n140_, mai_mai_n141_, mai_mai_n142_, mai_mai_n143_, mai_mai_n144_, mai_mai_n145_, mai_mai_n146_, mai_mai_n147_, mai_mai_n148_, mai_mai_n149_, mai_mai_n150_, mai_mai_n151_, mai_mai_n152_, mai_mai_n153_, mai_mai_n154_, mai_mai_n155_, mai_mai_n156_, mai_mai_n157_, mai_mai_n158_, mai_mai_n159_, mai_mai_n160_, mai_mai_n161_, mai_mai_n162_, mai_mai_n163_, mai_mai_n164_, mai_mai_n165_, mai_mai_n166_, mai_mai_n167_, mai_mai_n168_, mai_mai_n169_, mai_mai_n170_, mai_mai_n171_, mai_mai_n172_, mai_mai_n173_, mai_mai_n174_, mai_mai_n175_, mai_mai_n176_, mai_mai_n177_, mai_mai_n178_, mai_mai_n179_, mai_mai_n180_, mai_mai_n181_, mai_mai_n182_, mai_mai_n183_, mai_mai_n184_, mai_mai_n185_, mai_mai_n186_, mai_mai_n187_, mai_mai_n188_, mai_mai_n189_, mai_mai_n190_, mai_mai_n191_, mai_mai_n192_, mai_mai_n193_, mai_mai_n194_, mai_mai_n195_, mai_mai_n196_, mai_mai_n197_, mai_mai_n198_, mai_mai_n199_, mai_mai_n200_, mai_mai_n201_, mai_mai_n202_, mai_mai_n203_, mai_mai_n204_, mai_mai_n205_, mai_mai_n206_, mai_mai_n207_, mai_mai_n208_, mai_mai_n209_, mai_mai_n210_, mai_mai_n211_, mai_mai_n212_, mai_mai_n213_, mai_mai_n214_, mai_mai_n215_, mai_mai_n216_, mai_mai_n217_, mai_mai_n218_, mai_mai_n219_, mai_mai_n220_, mai_mai_n221_, mai_mai_n222_, mai_mai_n223_, mai_mai_n224_, mai_mai_n225_, mai_mai_n226_, mai_mai_n227_, mai_mai_n228_, mai_mai_n229_, mai_mai_n230_, mai_mai_n231_, mai_mai_n232_, mai_mai_n233_, mai_mai_n234_, mai_mai_n235_, mai_mai_n236_, mai_mai_n237_, mai_mai_n238_, mai_mai_n239_, mai_mai_n240_, mai_mai_n241_, mai_mai_n242_, mai_mai_n243_, mai_mai_n244_, mai_mai_n245_, mai_mai_n246_, mai_mai_n247_, mai_mai_n248_, mai_mai_n249_, mai_mai_n250_, mai_mai_n251_, mai_mai_n252_, mai_mai_n253_, mai_mai_n254_, mai_mai_n255_, mai_mai_n256_, mai_mai_n257_, mai_mai_n258_, mai_mai_n259_, mai_mai_n260_, mai_mai_n261_, mai_mai_n262_, mai_mai_n263_, mai_mai_n264_, mai_mai_n265_, mai_mai_n266_, mai_mai_n267_, mai_mai_n268_, mai_mai_n269_, mai_mai_n270_, mai_mai_n271_, mai_mai_n272_, mai_mai_n273_, mai_mai_n274_, mai_mai_n275_, mai_mai_n276_, mai_mai_n277_, mai_mai_n278_, mai_mai_n279_, mai_mai_n280_, mai_mai_n281_, mai_mai_n282_, mai_mai_n283_, mai_mai_n284_, mai_mai_n285_, mai_mai_n286_, mai_mai_n287_, mai_mai_n288_, mai_mai_n289_, mai_mai_n290_, mai_mai_n291_, mai_mai_n292_, mai_mai_n293_, mai_mai_n294_, mai_mai_n295_, mai_mai_n296_, mai_mai_n297_, mai_mai_n298_, mai_mai_n299_, mai_mai_n300_, mai_mai_n301_, mai_mai_n302_, mai_mai_n303_, mai_mai_n304_, mai_mai_n305_, mai_mai_n306_, mai_mai_n307_, mai_mai_n308_, mai_mai_n309_, mai_mai_n310_, mai_mai_n311_, mai_mai_n312_, mai_mai_n313_, mai_mai_n314_, mai_mai_n315_, mai_mai_n316_, mai_mai_n317_, mai_mai_n318_, mai_mai_n319_, mai_mai_n320_, mai_mai_n321_, mai_mai_n322_, mai_mai_n323_, mai_mai_n324_, mai_mai_n325_, mai_mai_n326_, mai_mai_n327_, mai_mai_n328_, mai_mai_n329_, mai_mai_n330_, mai_mai_n331_, mai_mai_n332_, mai_mai_n333_, mai_mai_n334_, mai_mai_n335_, mai_mai_n336_, mai_mai_n337_, mai_mai_n338_, mai_mai_n339_, mai_mai_n340_, mai_mai_n341_, mai_mai_n342_, mai_mai_n343_, mai_mai_n344_, mai_mai_n345_, mai_mai_n346_, mai_mai_n347_, mai_mai_n348_, mai_mai_n349_, mai_mai_n350_, mai_mai_n351_, mai_mai_n352_, mai_mai_n353_, mai_mai_n354_, mai_mai_n355_, mai_mai_n356_, mai_mai_n357_, mai_mai_n358_, mai_mai_n359_, mai_mai_n360_, mai_mai_n361_, mai_mai_n362_, mai_mai_n363_, mai_mai_n364_, mai_mai_n365_, mai_mai_n366_, mai_mai_n367_, mai_mai_n368_, mai_mai_n369_, mai_mai_n370_, mai_mai_n371_, mai_mai_n372_, mai_mai_n373_, mai_mai_n374_, mai_mai_n375_, mai_mai_n376_, mai_mai_n377_, mai_mai_n378_, mai_mai_n379_, mai_mai_n380_, mai_mai_n381_, mai_mai_n382_, mai_mai_n383_, mai_mai_n384_, mai_mai_n385_, mai_mai_n386_, mai_mai_n387_, mai_mai_n388_, mai_mai_n389_, mai_mai_n390_, mai_mai_n391_, mai_mai_n392_, mai_mai_n393_, mai_mai_n394_, mai_mai_n395_, mai_mai_n396_, mai_mai_n397_, mai_mai_n398_, mai_mai_n399_, mai_mai_n400_, mai_mai_n401_, mai_mai_n402_, mai_mai_n403_, mai_mai_n404_, mai_mai_n405_, mai_mai_n406_, mai_mai_n407_, mai_mai_n408_, mai_mai_n409_, mai_mai_n410_, mai_mai_n411_, mai_mai_n412_, mai_mai_n413_, mai_mai_n414_, mai_mai_n415_, mai_mai_n416_, mai_mai_n417_, mai_mai_n418_, mai_mai_n419_, mai_mai_n420_, mai_mai_n421_, mai_mai_n422_, mai_mai_n423_, mai_mai_n424_, mai_mai_n425_, mai_mai_n426_, mai_mai_n427_, mai_mai_n428_, mai_mai_n429_, mai_mai_n430_, mai_mai_n431_, mai_mai_n432_, mai_mai_n433_, mai_mai_n434_, mai_mai_n435_, mai_mai_n436_, mai_mai_n437_, mai_mai_n438_, mai_mai_n439_, mai_mai_n440_, mai_mai_n441_, mai_mai_n442_, mai_mai_n443_, mai_mai_n444_, mai_mai_n445_, mai_mai_n446_, mai_mai_n447_, mai_mai_n448_, mai_mai_n449_, mai_mai_n450_, mai_mai_n451_, mai_mai_n452_, mai_mai_n453_, mai_mai_n454_, mai_mai_n455_, mai_mai_n456_, mai_mai_n457_, mai_mai_n458_, mai_mai_n459_, mai_mai_n460_, mai_mai_n461_, mai_mai_n462_, mai_mai_n463_, mai_mai_n464_, mai_mai_n465_, mai_mai_n466_, mai_mai_n467_, mai_mai_n468_, mai_mai_n469_, mai_mai_n470_, mai_mai_n471_, mai_mai_n472_, mai_mai_n473_, mai_mai_n474_, mai_mai_n475_, mai_mai_n476_, mai_mai_n477_, mai_mai_n478_, mai_mai_n479_, mai_mai_n480_, mai_mai_n481_, mai_mai_n482_, mai_mai_n483_, mai_mai_n484_, mai_mai_n485_, mai_mai_n486_, mai_mai_n487_, mai_mai_n488_, mai_mai_n489_, mai_mai_n490_, mai_mai_n491_, mai_mai_n492_, mai_mai_n493_, mai_mai_n494_, mai_mai_n495_, mai_mai_n496_, mai_mai_n497_, mai_mai_n498_, mai_mai_n499_, mai_mai_n500_, mai_mai_n501_, mai_mai_n502_, mai_mai_n503_, mai_mai_n504_, mai_mai_n505_, mai_mai_n506_, mai_mai_n507_, mai_mai_n508_, mai_mai_n510_, mai_mai_n511_, mai_mai_n512_, mai_mai_n513_, mai_mai_n514_, mai_mai_n515_, mai_mai_n516_, mai_mai_n517_, mai_mai_n518_, mai_mai_n519_, mai_mai_n520_, mai_mai_n521_, mai_mai_n522_, mai_mai_n523_, mai_mai_n524_, mai_mai_n525_, mai_mai_n526_, mai_mai_n527_, mai_mai_n528_, mai_mai_n529_, mai_mai_n530_, mai_mai_n531_, mai_mai_n532_, mai_mai_n533_, mai_mai_n534_, mai_mai_n535_, mai_mai_n536_, mai_mai_n537_, mai_mai_n538_, mai_mai_n539_, mai_mai_n540_, mai_mai_n541_, mai_mai_n542_, mai_mai_n543_, mai_mai_n544_, mai_mai_n545_, mai_mai_n546_, mai_mai_n547_, mai_mai_n548_, mai_mai_n549_, mai_mai_n550_, mai_mai_n551_, mai_mai_n552_, mai_mai_n553_, mai_mai_n554_, mai_mai_n555_, mai_mai_n556_, mai_mai_n557_, mai_mai_n558_, mai_mai_n559_, mai_mai_n560_, mai_mai_n561_, mai_mai_n562_, mai_mai_n563_, mai_mai_n564_, mai_mai_n565_, mai_mai_n566_, mai_mai_n567_, mai_mai_n568_, mai_mai_n569_, mai_mai_n570_, mai_mai_n571_, mai_mai_n572_, mai_mai_n573_, mai_mai_n574_, mai_mai_n575_, mai_mai_n576_, mai_mai_n577_, mai_mai_n578_, mai_mai_n579_, mai_mai_n580_, mai_mai_n581_, mai_mai_n582_, mai_mai_n583_, mai_mai_n584_, mai_mai_n585_, mai_mai_n586_, mai_mai_n587_, mai_mai_n588_, mai_mai_n589_, mai_mai_n590_, mai_mai_n591_, mai_mai_n592_, mai_mai_n593_, mai_mai_n594_, mai_mai_n595_, mai_mai_n596_, mai_mai_n597_, mai_mai_n598_, mai_mai_n599_, mai_mai_n600_, mai_mai_n601_, mai_mai_n602_, mai_mai_n603_, mai_mai_n604_, mai_mai_n605_, mai_mai_n606_, mai_mai_n607_, mai_mai_n608_, mai_mai_n609_, mai_mai_n610_, mai_mai_n611_, mai_mai_n612_, mai_mai_n613_, mai_mai_n614_, mai_mai_n615_, mai_mai_n616_, mai_mai_n617_, mai_mai_n618_, mai_mai_n619_, mai_mai_n620_, mai_mai_n621_, mai_mai_n622_, mai_mai_n623_, mai_mai_n624_, mai_mai_n625_, mai_mai_n626_, mai_mai_n627_, mai_mai_n628_, mai_mai_n629_, mai_mai_n630_, mai_mai_n631_, mai_mai_n632_, mai_mai_n633_, mai_mai_n634_, mai_mai_n635_, mai_mai_n636_, mai_mai_n637_, mai_mai_n638_, mai_mai_n640_, mai_mai_n641_, mai_mai_n642_, mai_mai_n643_, mai_mai_n644_, mai_mai_n645_, mai_mai_n646_, mai_mai_n647_, mai_mai_n648_, mai_mai_n649_, mai_mai_n650_, mai_mai_n651_, mai_mai_n652_, mai_mai_n653_, mai_mai_n654_, mai_mai_n655_, mai_mai_n656_, mai_mai_n657_, mai_mai_n658_, mai_mai_n659_, mai_mai_n660_, mai_mai_n661_, mai_mai_n662_, mai_mai_n663_, mai_mai_n664_, mai_mai_n665_, mai_mai_n666_, mai_mai_n667_, mai_mai_n668_, mai_mai_n669_, mai_mai_n670_, mai_mai_n671_, mai_mai_n672_, mai_mai_n673_, mai_mai_n674_, mai_mai_n675_, mai_mai_n676_, mai_mai_n677_, mai_mai_n679_, mai_mai_n680_, mai_mai_n681_, mai_mai_n682_, mai_mai_n683_, mai_mai_n684_, mai_mai_n685_, mai_mai_n686_, mai_mai_n687_, mai_mai_n688_, mai_mai_n689_, mai_mai_n690_, mai_mai_n691_, mai_mai_n692_, mai_mai_n693_, mai_mai_n694_, mai_mai_n695_, mai_mai_n696_, mai_mai_n697_, mai_mai_n698_, mai_mai_n699_, mai_mai_n700_, mai_mai_n701_, mai_mai_n702_, mai_mai_n703_, mai_mai_n704_, mai_mai_n705_, mai_mai_n706_, mai_mai_n707_, mai_mai_n708_, mai_mai_n709_, mai_mai_n710_, mai_mai_n711_, mai_mai_n712_, mai_mai_n713_, mai_mai_n714_, mai_mai_n715_, mai_mai_n716_, mai_mai_n717_, mai_mai_n718_, mai_mai_n719_, mai_mai_n720_, mai_mai_n721_, mai_mai_n722_, mai_mai_n724_, mai_mai_n725_, mai_mai_n726_, mai_mai_n727_, mai_mai_n728_, mai_mai_n729_, mai_mai_n730_, mai_mai_n731_, mai_mai_n732_, mai_mai_n733_, mai_mai_n734_, mai_mai_n735_, mai_mai_n736_, mai_mai_n737_, mai_mai_n738_, mai_mai_n739_, mai_mai_n740_, mai_mai_n741_, mai_mai_n742_, mai_mai_n743_, mai_mai_n744_, mai_mai_n745_, mai_mai_n746_, mai_mai_n747_, mai_mai_n748_, mai_mai_n749_, mai_mai_n750_, mai_mai_n751_, mai_mai_n752_, mai_mai_n753_, mai_mai_n754_, mai_mai_n755_, mai_mai_n756_, mai_mai_n757_, mai_mai_n758_, mai_mai_n759_, mai_mai_n760_, mai_mai_n761_, mai_mai_n762_, mai_mai_n763_, mai_mai_n764_, mai_mai_n765_, mai_mai_n766_, mai_mai_n767_, mai_mai_n768_, mai_mai_n769_, mai_mai_n770_, mai_mai_n771_, mai_mai_n772_, mai_mai_n773_, mai_mai_n774_, mai_mai_n775_, mai_mai_n776_, mai_mai_n777_, mai_mai_n778_, mai_mai_n779_, mai_mai_n780_, mai_mai_n781_, mai_mai_n782_, mai_mai_n783_, mai_mai_n784_, mai_mai_n785_, mai_mai_n786_, mai_mai_n787_, mai_mai_n788_, mai_mai_n789_, mai_mai_n790_, mai_mai_n791_, mai_mai_n792_, mai_mai_n793_, mai_mai_n794_, mai_mai_n795_, mai_mai_n796_, mai_mai_n797_, mai_mai_n798_, mai_mai_n799_, mai_mai_n800_, mai_mai_n801_, mai_mai_n802_, mai_mai_n803_, mai_mai_n804_, mai_mai_n805_, mai_mai_n806_, mai_mai_n807_, mai_mai_n808_, mai_mai_n809_, mai_mai_n810_, mai_mai_n811_, mai_mai_n812_, mai_mai_n813_, mai_mai_n814_, mai_mai_n815_, mai_mai_n816_, mai_mai_n817_, mai_mai_n818_, mai_mai_n819_, mai_mai_n820_, mai_mai_n821_, mai_mai_n822_, mai_mai_n823_, mai_mai_n824_, mai_mai_n825_, mai_mai_n826_, mai_mai_n827_, mai_mai_n828_, mai_mai_n829_, mai_mai_n830_, mai_mai_n831_, mai_mai_n832_, mai_mai_n833_, mai_mai_n834_, mai_mai_n835_, mai_mai_n836_, mai_mai_n837_, mai_mai_n838_, mai_mai_n839_, mai_mai_n840_, mai_mai_n841_, mai_mai_n842_, mai_mai_n843_, mai_mai_n844_, mai_mai_n845_, mai_mai_n846_, mai_mai_n847_, mai_mai_n848_, mai_mai_n849_, mai_mai_n850_, mai_mai_n851_, mai_mai_n852_, mai_mai_n853_, mai_mai_n854_, mai_mai_n855_, mai_mai_n856_, mai_mai_n857_, mai_mai_n858_, mai_mai_n859_, mai_mai_n860_, mai_mai_n861_, mai_mai_n862_, mai_mai_n863_, mai_mai_n864_, mai_mai_n865_, mai_mai_n866_, mai_mai_n867_, mai_mai_n868_, mai_mai_n869_, mai_mai_n870_, mai_mai_n871_, mai_mai_n872_, mai_mai_n873_, mai_mai_n874_, mai_mai_n875_, mai_mai_n876_, mai_mai_n877_, mai_mai_n878_, mai_mai_n879_, mai_mai_n880_, mai_mai_n881_, mai_mai_n882_, mai_mai_n883_, mai_mai_n884_, mai_mai_n885_, mai_mai_n886_, mai_mai_n887_, mai_mai_n888_, mai_mai_n889_, mai_mai_n890_, mai_mai_n891_, mai_mai_n892_, mai_mai_n893_, mai_mai_n894_, mai_mai_n895_, mai_mai_n896_, mai_mai_n897_, mai_mai_n901_, mai_mai_n902_, mai_mai_n903_, mai_mai_n904_, mai_mai_n905_, mai_mai_n906_, mai_mai_n907_, mai_mai_n908_, mai_mai_n909_, mai_mai_n910_, mai_mai_n911_, mai_mai_n912_, mai_mai_n913_, mai_mai_n914_, mai_mai_n915_, mai_mai_n916_, mai_mai_n917_, men_men_n23_, men_men_n24_, men_men_n25_, men_men_n26_, men_men_n27_, men_men_n28_, men_men_n29_, men_men_n30_, men_men_n31_, men_men_n32_, men_men_n33_, men_men_n34_, men_men_n35_, men_men_n36_, men_men_n37_, men_men_n38_, men_men_n39_, men_men_n40_, men_men_n41_, men_men_n43_, men_men_n44_, men_men_n45_, men_men_n46_, men_men_n47_, men_men_n48_, men_men_n49_, men_men_n50_, men_men_n51_, men_men_n52_, men_men_n53_, men_men_n54_, men_men_n55_, men_men_n56_, men_men_n57_, men_men_n58_, men_men_n59_, men_men_n60_, men_men_n61_, men_men_n62_, men_men_n63_, men_men_n64_, men_men_n65_, men_men_n66_, men_men_n67_, men_men_n68_, men_men_n69_, men_men_n70_, men_men_n71_, men_men_n72_, men_men_n73_, men_men_n74_, men_men_n75_, men_men_n76_, men_men_n77_, men_men_n78_, men_men_n79_, men_men_n80_, men_men_n81_, men_men_n82_, men_men_n83_, men_men_n84_, men_men_n85_, men_men_n86_, men_men_n87_, men_men_n88_, men_men_n89_, men_men_n90_, men_men_n91_, men_men_n92_, men_men_n93_, men_men_n94_, men_men_n95_, men_men_n96_, men_men_n97_, men_men_n98_, men_men_n99_, men_men_n100_, men_men_n101_, men_men_n102_, men_men_n103_, men_men_n104_, men_men_n105_, men_men_n106_, men_men_n107_, men_men_n108_, men_men_n109_, men_men_n110_, men_men_n111_, men_men_n112_, men_men_n113_, men_men_n114_, men_men_n115_, men_men_n116_, men_men_n117_, men_men_n118_, men_men_n119_, men_men_n120_, men_men_n121_, men_men_n122_, men_men_n123_, men_men_n124_, men_men_n125_, men_men_n126_, men_men_n127_, men_men_n128_, men_men_n129_, men_men_n132_, men_men_n133_, men_men_n134_, men_men_n135_, men_men_n136_, men_men_n137_, men_men_n138_, men_men_n139_, men_men_n140_, men_men_n141_, men_men_n142_, men_men_n143_, men_men_n144_, men_men_n145_, men_men_n146_, men_men_n147_, men_men_n148_, men_men_n149_, men_men_n150_, men_men_n151_, men_men_n152_, men_men_n153_, men_men_n154_, men_men_n155_, men_men_n156_, men_men_n157_, men_men_n158_, men_men_n159_, men_men_n160_, men_men_n161_, men_men_n162_, men_men_n163_, men_men_n164_, men_men_n165_, men_men_n166_, men_men_n167_, men_men_n168_, men_men_n169_, men_men_n170_, men_men_n171_, men_men_n172_, men_men_n173_, men_men_n174_, men_men_n175_, men_men_n176_, men_men_n177_, men_men_n178_, men_men_n179_, men_men_n180_, men_men_n181_, men_men_n182_, men_men_n183_, men_men_n184_, men_men_n185_, men_men_n186_, men_men_n187_, men_men_n188_, men_men_n189_, men_men_n190_, men_men_n191_, men_men_n192_, men_men_n193_, men_men_n194_, men_men_n195_, men_men_n196_, men_men_n197_, men_men_n198_, men_men_n199_, men_men_n200_, men_men_n201_, men_men_n202_, men_men_n203_, men_men_n204_, men_men_n205_, men_men_n206_, men_men_n207_, men_men_n208_, men_men_n209_, men_men_n210_, men_men_n211_, men_men_n212_, men_men_n213_, men_men_n214_, men_men_n215_, men_men_n216_, men_men_n217_, men_men_n218_, men_men_n219_, men_men_n220_, men_men_n221_, men_men_n222_, men_men_n223_, men_men_n224_, men_men_n225_, men_men_n226_, men_men_n227_, men_men_n228_, men_men_n229_, men_men_n230_, men_men_n231_, men_men_n232_, men_men_n233_, men_men_n234_, men_men_n235_, men_men_n236_, men_men_n237_, men_men_n238_, men_men_n239_, men_men_n240_, men_men_n241_, men_men_n242_, men_men_n243_, men_men_n244_, men_men_n245_, men_men_n246_, men_men_n247_, men_men_n248_, men_men_n249_, men_men_n250_, men_men_n251_, men_men_n252_, men_men_n253_, men_men_n254_, men_men_n255_, men_men_n256_, men_men_n257_, men_men_n258_, men_men_n259_, men_men_n260_, men_men_n261_, men_men_n262_, men_men_n263_, men_men_n264_, men_men_n265_, men_men_n266_, men_men_n267_, men_men_n268_, men_men_n269_, men_men_n270_, men_men_n271_, men_men_n272_, men_men_n273_, men_men_n274_, men_men_n275_, men_men_n276_, men_men_n277_, men_men_n278_, men_men_n279_, men_men_n280_, men_men_n281_, men_men_n282_, men_men_n283_, men_men_n284_, men_men_n285_, men_men_n286_, men_men_n287_, men_men_n288_, men_men_n289_, men_men_n290_, men_men_n291_, men_men_n292_, men_men_n293_, men_men_n294_, men_men_n295_, men_men_n296_, men_men_n297_, men_men_n298_, men_men_n299_, men_men_n300_, men_men_n301_, men_men_n302_, men_men_n303_, men_men_n304_, men_men_n305_, men_men_n306_, men_men_n307_, men_men_n308_, men_men_n309_, men_men_n310_, men_men_n311_, men_men_n312_, men_men_n313_, men_men_n314_, men_men_n315_, men_men_n316_, men_men_n317_, men_men_n318_, men_men_n319_, men_men_n320_, men_men_n321_, men_men_n322_, men_men_n323_, men_men_n324_, men_men_n325_, men_men_n326_, men_men_n327_, men_men_n328_, men_men_n329_, men_men_n330_, men_men_n331_, men_men_n332_, men_men_n333_, men_men_n334_, men_men_n335_, men_men_n336_, men_men_n337_, men_men_n338_, men_men_n339_, men_men_n340_, men_men_n341_, men_men_n342_, men_men_n343_, men_men_n344_, men_men_n345_, men_men_n346_, men_men_n347_, men_men_n348_, men_men_n349_, men_men_n350_, men_men_n351_, men_men_n352_, men_men_n353_, men_men_n354_, men_men_n355_, men_men_n356_, men_men_n357_, men_men_n358_, men_men_n359_, men_men_n360_, men_men_n361_, men_men_n362_, men_men_n363_, men_men_n364_, men_men_n365_, men_men_n366_, men_men_n367_, men_men_n368_, men_men_n369_, men_men_n370_, men_men_n371_, men_men_n372_, men_men_n373_, men_men_n374_, men_men_n375_, men_men_n376_, men_men_n377_, men_men_n378_, men_men_n379_, men_men_n380_, men_men_n381_, men_men_n382_, men_men_n383_, men_men_n384_, men_men_n385_, men_men_n386_, men_men_n387_, men_men_n388_, men_men_n389_, men_men_n390_, men_men_n391_, men_men_n392_, men_men_n393_, men_men_n394_, men_men_n395_, men_men_n396_, men_men_n397_, men_men_n398_, men_men_n399_, men_men_n400_, men_men_n401_, men_men_n402_, men_men_n403_, men_men_n404_, men_men_n405_, men_men_n406_, men_men_n407_, men_men_n408_, men_men_n409_, men_men_n410_, men_men_n411_, men_men_n412_, men_men_n413_, men_men_n414_, men_men_n415_, men_men_n416_, men_men_n417_, men_men_n418_, men_men_n419_, men_men_n420_, men_men_n421_, men_men_n422_, men_men_n423_, men_men_n424_, men_men_n425_, men_men_n426_, men_men_n427_, men_men_n428_, men_men_n429_, men_men_n430_, men_men_n431_, men_men_n432_, men_men_n433_, men_men_n434_, men_men_n435_, men_men_n436_, men_men_n437_, men_men_n438_, men_men_n439_, men_men_n440_, men_men_n441_, men_men_n442_, men_men_n443_, men_men_n444_, men_men_n445_, men_men_n446_, men_men_n447_, men_men_n448_, men_men_n449_, men_men_n450_, men_men_n451_, men_men_n452_, men_men_n453_, men_men_n454_, men_men_n455_, men_men_n456_, men_men_n457_, men_men_n458_, men_men_n459_, men_men_n460_, men_men_n461_, men_men_n462_, men_men_n463_, men_men_n464_, men_men_n465_, men_men_n466_, men_men_n467_, men_men_n468_, men_men_n469_, men_men_n470_, men_men_n471_, men_men_n472_, men_men_n473_, men_men_n474_, men_men_n475_, men_men_n476_, men_men_n477_, men_men_n478_, men_men_n479_, men_men_n480_, men_men_n481_, men_men_n482_, men_men_n483_, men_men_n484_, men_men_n485_, men_men_n486_, men_men_n487_, men_men_n488_, men_men_n489_, men_men_n490_, men_men_n491_, men_men_n492_, men_men_n493_, men_men_n494_, men_men_n495_, men_men_n496_, men_men_n497_, men_men_n498_, men_men_n499_, men_men_n500_, men_men_n501_, men_men_n502_, men_men_n503_, men_men_n504_, men_men_n505_, men_men_n506_, men_men_n507_, men_men_n508_, men_men_n509_, men_men_n510_, men_men_n511_, men_men_n512_, men_men_n513_, men_men_n514_, men_men_n515_, men_men_n516_, men_men_n517_, men_men_n518_, men_men_n519_, men_men_n520_, men_men_n521_, men_men_n522_, men_men_n523_, men_men_n524_, men_men_n525_, men_men_n526_, men_men_n527_, men_men_n528_, men_men_n529_, men_men_n530_, men_men_n531_, men_men_n532_, men_men_n533_, men_men_n534_, men_men_n535_, men_men_n536_, men_men_n537_, men_men_n538_, men_men_n539_, men_men_n540_, men_men_n541_, men_men_n542_, men_men_n543_, men_men_n544_, men_men_n545_, men_men_n546_, men_men_n547_, men_men_n548_, men_men_n549_, men_men_n550_, men_men_n551_, men_men_n552_, men_men_n553_, men_men_n554_, men_men_n555_, men_men_n556_, men_men_n557_, men_men_n558_, men_men_n559_, men_men_n560_, men_men_n561_, men_men_n562_, men_men_n563_, men_men_n564_, men_men_n565_, men_men_n566_, men_men_n567_, men_men_n568_, men_men_n569_, men_men_n570_, men_men_n571_, men_men_n572_, men_men_n573_, men_men_n574_, men_men_n575_, men_men_n576_, men_men_n577_, men_men_n578_, men_men_n579_, men_men_n580_, men_men_n581_, men_men_n582_, men_men_n583_, men_men_n584_, men_men_n585_, men_men_n586_, men_men_n587_, men_men_n589_, men_men_n590_, men_men_n591_, men_men_n592_, men_men_n593_, men_men_n594_, men_men_n595_, men_men_n596_, men_men_n597_, men_men_n598_, men_men_n599_, men_men_n600_, men_men_n601_, men_men_n602_, men_men_n603_, men_men_n604_, men_men_n605_, men_men_n606_, men_men_n607_, men_men_n608_, men_men_n609_, men_men_n610_, men_men_n611_, men_men_n612_, men_men_n613_, men_men_n614_, men_men_n615_, men_men_n616_, men_men_n617_, men_men_n618_, men_men_n619_, men_men_n620_, men_men_n621_, men_men_n622_, men_men_n623_, men_men_n624_, men_men_n625_, men_men_n626_, men_men_n627_, men_men_n628_, men_men_n629_, men_men_n630_, men_men_n631_, men_men_n632_, men_men_n633_, men_men_n634_, men_men_n635_, men_men_n636_, men_men_n637_, men_men_n638_, men_men_n639_, men_men_n640_, men_men_n641_, men_men_n642_, men_men_n643_, men_men_n644_, men_men_n645_, men_men_n646_, men_men_n647_, men_men_n648_, men_men_n649_, men_men_n650_, men_men_n651_, men_men_n652_, men_men_n653_, men_men_n654_, men_men_n655_, men_men_n656_, men_men_n657_, men_men_n658_, men_men_n659_, men_men_n660_, men_men_n661_, men_men_n662_, men_men_n663_, men_men_n664_, men_men_n665_, men_men_n666_, men_men_n667_, men_men_n668_, men_men_n669_, men_men_n670_, men_men_n671_, men_men_n672_, men_men_n673_, men_men_n674_, men_men_n675_, men_men_n676_, men_men_n677_, men_men_n678_, men_men_n679_, men_men_n680_, men_men_n681_, men_men_n682_, men_men_n683_, men_men_n684_, men_men_n685_, men_men_n686_, men_men_n687_, men_men_n688_, men_men_n689_, men_men_n690_, men_men_n691_, men_men_n692_, men_men_n693_, men_men_n694_, men_men_n695_, men_men_n696_, men_men_n697_, men_men_n698_, men_men_n699_, men_men_n700_, men_men_n701_, men_men_n702_, men_men_n703_, men_men_n704_, men_men_n705_, men_men_n706_, men_men_n707_, men_men_n709_, men_men_n710_, men_men_n711_, men_men_n712_, men_men_n713_, men_men_n714_, men_men_n715_, men_men_n716_, men_men_n717_, men_men_n718_, men_men_n719_, men_men_n720_, men_men_n721_, men_men_n722_, men_men_n723_, men_men_n724_, men_men_n725_, men_men_n726_, men_men_n727_, men_men_n728_, men_men_n729_, men_men_n730_, men_men_n731_, men_men_n732_, men_men_n733_, men_men_n734_, men_men_n735_, men_men_n736_, men_men_n737_, men_men_n738_, men_men_n739_, men_men_n740_, men_men_n741_, men_men_n742_, men_men_n743_, men_men_n744_, men_men_n745_, men_men_n746_, men_men_n748_, men_men_n749_, men_men_n750_, men_men_n751_, men_men_n752_, men_men_n753_, men_men_n754_, men_men_n755_, men_men_n756_, men_men_n757_, men_men_n758_, men_men_n759_, men_men_n760_, men_men_n761_, men_men_n762_, men_men_n763_, men_men_n764_, men_men_n765_, men_men_n766_, men_men_n767_, men_men_n768_, men_men_n769_, men_men_n770_, men_men_n771_, men_men_n772_, men_men_n773_, men_men_n774_, men_men_n775_, men_men_n776_, men_men_n777_, men_men_n778_, men_men_n779_, men_men_n780_, men_men_n781_, men_men_n782_, men_men_n783_, men_men_n784_, men_men_n785_, men_men_n787_, men_men_n788_, men_men_n789_, men_men_n790_, men_men_n791_, men_men_n792_, men_men_n793_, men_men_n794_, men_men_n795_, men_men_n796_, men_men_n797_, men_men_n798_, men_men_n799_, men_men_n800_, men_men_n801_, men_men_n802_, men_men_n803_, men_men_n804_, men_men_n805_, men_men_n806_, men_men_n807_, men_men_n808_, men_men_n809_, men_men_n810_, men_men_n811_, men_men_n812_, men_men_n813_, men_men_n814_, men_men_n815_, men_men_n816_, men_men_n817_, men_men_n818_, men_men_n819_, men_men_n820_, men_men_n821_, men_men_n822_, men_men_n823_, men_men_n824_, men_men_n825_, men_men_n826_, men_men_n827_, men_men_n828_, men_men_n829_, men_men_n830_, men_men_n831_, men_men_n832_, men_men_n833_, men_men_n834_, men_men_n835_, men_men_n836_, men_men_n837_, men_men_n838_, men_men_n839_, men_men_n840_, men_men_n841_, men_men_n842_, men_men_n843_, men_men_n844_, men_men_n845_, men_men_n846_, men_men_n847_, men_men_n848_, men_men_n849_, men_men_n850_, men_men_n851_, men_men_n852_, men_men_n853_, men_men_n854_, men_men_n855_, men_men_n856_, men_men_n857_, men_men_n858_, men_men_n859_, men_men_n860_, men_men_n861_, men_men_n862_, men_men_n863_, men_men_n864_, men_men_n865_, men_men_n866_, men_men_n867_, men_men_n868_, men_men_n869_, men_men_n870_, men_men_n871_, men_men_n872_, men_men_n873_, men_men_n874_, men_men_n875_, men_men_n876_, men_men_n877_, men_men_n878_, men_men_n879_, men_men_n880_, men_men_n881_, men_men_n882_, men_men_n883_, men_men_n884_, men_men_n885_, men_men_n886_, men_men_n887_, men_men_n888_, men_men_n889_, men_men_n890_, men_men_n891_, men_men_n892_, men_men_n893_, men_men_n894_, men_men_n895_, men_men_n896_, men_men_n897_, men_men_n898_, men_men_n899_, men_men_n900_, men_men_n901_, men_men_n902_, men_men_n903_, men_men_n904_, men_men_n905_, men_men_n906_, men_men_n907_, men_men_n908_, men_men_n909_, men_men_n910_, men_men_n911_, men_men_n912_, men_men_n913_, men_men_n914_, men_men_n915_, men_men_n916_, men_men_n917_, men_men_n918_, men_men_n919_, men_men_n920_, men_men_n921_, men_men_n922_, men_men_n923_, men_men_n924_, men_men_n925_, men_men_n926_, men_men_n927_, men_men_n928_, men_men_n929_, men_men_n930_, men_men_n931_, men_men_n932_, men_men_n933_, men_men_n934_, men_men_n935_, men_men_n936_, men_men_n937_, men_men_n938_, men_men_n939_, men_men_n940_, men_men_n941_, men_men_n942_, men_men_n943_, men_men_n944_, men_men_n945_, men_men_n946_, men_men_n947_, men_men_n948_, men_men_n949_, men_men_n950_, men_men_n951_, men_men_n952_, men_men_n953_, men_men_n954_, men_men_n955_, men_men_n956_, men_men_n957_, men_men_n958_, men_men_n959_, men_men_n960_, men_men_n961_, men_men_n962_, men_men_n963_, men_men_n964_, men_men_n965_, men_men_n966_, men_men_n967_, men_men_n968_, men_men_n969_, men_men_n970_, men_men_n971_, men_men_n972_, men_men_n973_, men_men_n974_, men_men_n975_, men_men_n976_, men_men_n977_, men_men_n978_, men_men_n979_, men_men_n980_, men_men_n981_, men_men_n982_, men_men_n983_, men_men_n984_, men_men_n985_, men_men_n986_, men_men_n987_, men_men_n988_, men_men_n989_, men_men_n990_, men_men_n991_, men_men_n992_, men_men_n993_, men_men_n994_, men_men_n995_, men_men_n996_, men_men_n997_, men_men_n998_, men_men_n999_, men_men_n1000_, men_men_n1001_, men_men_n1002_, men_men_n1003_, men_men_n1004_, men_men_n1005_, men_men_n1006_, men_men_n1010_, men_men_n1011_, men_men_n1012_, men_men_n1013_, men_men_n1014_, men_men_n1015_, men_men_n1016_, men_men_n1017_, men_men_n1018_, men_men_n1019_, men_men_n1020_, men_men_n1021_, men_men_n1022_, ori0, mai0, men0, ori1, mai1, men1, ori2, mai2, men2, ori3, mai3, men3, ori4, mai4, men4, ori5, mai5, men5, ori6, mai6, men6, ori7, mai7, men7;
  NAi21      o000(.An(i_13_), .B(i_4_), .Y(ori_ori_n23_));
  NOi21      o001(.An(i_3_), .B(i_8_), .Y(ori_ori_n24_));
  INV        o002(.A(i_9_), .Y(ori_ori_n25_));
  INV        o003(.A(i_3_), .Y(ori_ori_n26_));
  NO2        o004(.A(ori_ori_n26_), .B(ori_ori_n25_), .Y(ori_ori_n27_));
  NO2        o005(.A(i_8_), .B(i_10_), .Y(ori_ori_n28_));
  INV        o006(.A(ori_ori_n28_), .Y(ori_ori_n29_));
  OAI210     o007(.A0(ori_ori_n27_), .A1(ori_ori_n24_), .B0(ori_ori_n29_), .Y(ori_ori_n30_));
  AO210      o008(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(ori_ori_n31_));
  OR2        o009(.A(ori_ori_n31_), .B(i_11_), .Y(ori_ori_n32_));
  NA2        o010(.A(ori_ori_n32_), .B(ori_ori_n30_), .Y(ori_ori_n33_));
  XO2        o011(.A(ori_ori_n33_), .B(ori_ori_n23_), .Y(ori_ori_n34_));
  INV        o012(.A(i_4_), .Y(ori_ori_n35_));
  INV        o013(.A(i_10_), .Y(ori_ori_n36_));
  NAi21      o014(.An(i_11_), .B(i_9_), .Y(ori_ori_n37_));
  NO3        o015(.A(ori_ori_n37_), .B(i_12_), .C(ori_ori_n36_), .Y(ori_ori_n38_));
  NOi21      o016(.An(i_12_), .B(i_13_), .Y(ori_ori_n39_));
  INV        o017(.A(ori_ori_n39_), .Y(ori_ori_n40_));
  INV        o018(.A(ori_ori_n34_), .Y(ori1));
  INV        o019(.A(i_11_), .Y(ori_ori_n42_));
  NO2        o020(.A(ori_ori_n42_), .B(i_6_), .Y(ori_ori_n43_));
  INV        o021(.A(i_2_), .Y(ori_ori_n44_));
  INV        o022(.A(i_5_), .Y(ori_ori_n45_));
  NO2        o023(.A(i_7_), .B(i_10_), .Y(ori_ori_n46_));
  AOI210     o024(.A0(i_7_), .A1(ori_ori_n25_), .B0(ori_ori_n46_), .Y(ori_ori_n47_));
  NA2        o025(.A(i_0_), .B(i_2_), .Y(ori_ori_n48_));
  NA2        o026(.A(i_7_), .B(i_9_), .Y(ori_ori_n49_));
  NO2        o027(.A(ori_ori_n49_), .B(ori_ori_n48_), .Y(ori_ori_n50_));
  NO2        o028(.A(i_1_), .B(i_6_), .Y(ori_ori_n51_));
  NA2        o029(.A(i_8_), .B(i_7_), .Y(ori_ori_n52_));
  NAi21      o030(.An(i_2_), .B(i_7_), .Y(ori_ori_n53_));
  INV        o031(.A(i_1_), .Y(ori_ori_n54_));
  NA2        o032(.A(ori_ori_n54_), .B(i_6_), .Y(ori_ori_n55_));
  INV        o033(.A(i_10_), .Y(ori_ori_n56_));
  NO2        o034(.A(ori_ori_n56_), .B(i_6_), .Y(ori_ori_n57_));
  NAi21      o035(.An(ori_ori_n57_), .B(ori_ori_n52_), .Y(ori_ori_n58_));
  NA2        o036(.A(ori_ori_n47_), .B(i_2_), .Y(ori_ori_n59_));
  AOI210     o037(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(ori_ori_n60_));
  NA2        o038(.A(i_1_), .B(i_6_), .Y(ori_ori_n61_));
  NO2        o039(.A(ori_ori_n61_), .B(ori_ori_n25_), .Y(ori_ori_n62_));
  INV        o040(.A(i_0_), .Y(ori_ori_n63_));
  NA2        o041(.A(i_5_), .B(i_9_), .Y(ori_ori_n64_));
  INV        o042(.A(ori_ori_n62_), .Y(ori_ori_n65_));
  NA2        o043(.A(ori_ori_n59_), .B(ori_ori_n65_), .Y(ori_ori_n66_));
  OAI210     o044(.A0(ori_ori_n66_), .A1(ori_ori_n58_), .B0(i_0_), .Y(ori_ori_n67_));
  NA2        o045(.A(i_12_), .B(i_5_), .Y(ori_ori_n68_));
  NO2        o046(.A(i_3_), .B(i_9_), .Y(ori_ori_n69_));
  NO2        o047(.A(i_3_), .B(i_7_), .Y(ori_ori_n70_));
  NO2        o048(.A(ori_ori_n69_), .B(ori_ori_n54_), .Y(ori_ori_n71_));
  INV        o049(.A(i_6_), .Y(ori_ori_n72_));
  NO2        o050(.A(i_2_), .B(i_7_), .Y(ori_ori_n73_));
  INV        o051(.A(ori_ori_n73_), .Y(ori_ori_n74_));
  OAI210     o052(.A0(ori_ori_n71_), .A1(i_8_), .B0(ori_ori_n74_), .Y(ori_ori_n75_));
  NAi21      o053(.An(i_6_), .B(i_10_), .Y(ori_ori_n76_));
  NA2        o054(.A(i_6_), .B(i_9_), .Y(ori_ori_n77_));
  AOI210     o055(.A0(ori_ori_n77_), .A1(ori_ori_n76_), .B0(ori_ori_n54_), .Y(ori_ori_n78_));
  NA2        o056(.A(i_2_), .B(i_6_), .Y(ori_ori_n79_));
  NO2        o057(.A(ori_ori_n79_), .B(ori_ori_n25_), .Y(ori_ori_n80_));
  NO2        o058(.A(ori_ori_n80_), .B(ori_ori_n78_), .Y(ori_ori_n81_));
  AOI210     o059(.A0(ori_ori_n81_), .A1(ori_ori_n75_), .B0(ori_ori_n68_), .Y(ori_ori_n82_));
  AN3        o060(.A(i_0_), .B(i_2_), .C(i_1_), .Y(ori_ori_n83_));
  NAi21      o061(.An(i_6_), .B(i_11_), .Y(ori_ori_n84_));
  INV        o062(.A(i_7_), .Y(ori_ori_n85_));
  NA2        o063(.A(ori_ori_n44_), .B(ori_ori_n85_), .Y(ori_ori_n86_));
  NO2        o064(.A(i_0_), .B(i_5_), .Y(ori_ori_n87_));
  NO2        o065(.A(ori_ori_n87_), .B(ori_ori_n72_), .Y(ori_ori_n88_));
  NA2        o066(.A(i_12_), .B(i_3_), .Y(ori_ori_n89_));
  INV        o067(.A(ori_ori_n89_), .Y(ori_ori_n90_));
  NA3        o068(.A(ori_ori_n90_), .B(ori_ori_n88_), .C(ori_ori_n86_), .Y(ori_ori_n91_));
  NAi21      o069(.An(i_7_), .B(i_11_), .Y(ori_ori_n92_));
  AN2        o070(.A(i_2_), .B(i_10_), .Y(ori_ori_n93_));
  BUFFER     o071(.A(ori_ori_n68_), .Y(ori_ori_n94_));
  NO2        o072(.A(ori_ori_n54_), .B(ori_ori_n26_), .Y(ori_ori_n95_));
  NA2        o073(.A(i_11_), .B(i_12_), .Y(ori_ori_n96_));
  INV        o074(.A(ori_ori_n91_), .Y(ori_ori_n97_));
  NA2        o075(.A(ori_ori_n85_), .B(ori_ori_n36_), .Y(ori_ori_n98_));
  NA2        o076(.A(i_7_), .B(ori_ori_n25_), .Y(ori_ori_n99_));
  NA2        o077(.A(ori_ori_n99_), .B(ori_ori_n98_), .Y(ori_ori_n100_));
  NO2        o078(.A(ori_ori_n100_), .B(ori_ori_n44_), .Y(ori_ori_n101_));
  NA2        o079(.A(ori_ori_n77_), .B(ori_ori_n76_), .Y(ori_ori_n102_));
  NAi21      o080(.An(i_3_), .B(i_8_), .Y(ori_ori_n103_));
  NO2        o081(.A(i_1_), .B(ori_ori_n72_), .Y(ori_ori_n104_));
  NO2        o082(.A(i_6_), .B(i_5_), .Y(ori_ori_n105_));
  NO3        o083(.A(i_11_), .B(ori_ori_n97_), .C(ori_ori_n82_), .Y(ori_ori_n106_));
  NA2        o084(.A(ori_ori_n106_), .B(ori_ori_n67_), .Y(ori2));
  NO2        o085(.A(ori_ori_n54_), .B(ori_ori_n36_), .Y(ori_ori_n108_));
  INV        o086(.A(i_6_), .Y(ori_ori_n109_));
  NA2        o087(.A(ori_ori_n109_), .B(ori_ori_n108_), .Y(ori_ori_n110_));
  NA4        o088(.A(ori_ori_n110_), .B(ori_ori_n65_), .C(ori_ori_n59_), .D(ori_ori_n30_), .Y(ori0));
  AN2        o089(.A(i_8_), .B(i_7_), .Y(ori_ori_n112_));
  NA2        o090(.A(ori_ori_n112_), .B(i_6_), .Y(ori_ori_n113_));
  NO2        o091(.A(i_12_), .B(i_13_), .Y(ori_ori_n114_));
  NAi21      o092(.An(i_5_), .B(i_11_), .Y(ori_ori_n115_));
  NO2        o093(.A(i_0_), .B(i_1_), .Y(ori_ori_n116_));
  AN2        o094(.A(ori_ori_n114_), .B(ori_ori_n69_), .Y(ori_ori_n117_));
  NA2        o095(.A(i_1_), .B(i_5_), .Y(ori_ori_n118_));
  OR2        o096(.A(i_0_), .B(i_1_), .Y(ori_ori_n119_));
  NOi21      o097(.An(i_4_), .B(i_10_), .Y(ori_ori_n120_));
  NA2        o098(.A(ori_ori_n120_), .B(ori_ori_n39_), .Y(ori_ori_n121_));
  NOi21      o099(.An(i_4_), .B(i_9_), .Y(ori_ori_n122_));
  NOi21      o100(.An(i_11_), .B(i_13_), .Y(ori_ori_n123_));
  NO2        o101(.A(ori_ori_n63_), .B(ori_ori_n54_), .Y(ori_ori_n124_));
  NO2        o102(.A(ori_ori_n63_), .B(i_5_), .Y(ori_ori_n125_));
  NO2        o103(.A(i_2_), .B(i_1_), .Y(ori_ori_n126_));
  NAi21      o104(.An(i_4_), .B(i_12_), .Y(ori_ori_n127_));
  INV        o105(.A(i_8_), .Y(ori_ori_n128_));
  NO2        o106(.A(i_3_), .B(i_8_), .Y(ori_ori_n129_));
  NO3        o107(.A(i_11_), .B(i_10_), .C(i_9_), .Y(ori_ori_n130_));
  NO2        o108(.A(ori_ori_n87_), .B(ori_ori_n51_), .Y(ori_ori_n131_));
  NO2        o109(.A(i_13_), .B(i_9_), .Y(ori_ori_n132_));
  NO2        o110(.A(ori_ori_n42_), .B(i_5_), .Y(ori_ori_n133_));
  NA2        o111(.A(i_0_), .B(i_5_), .Y(ori_ori_n134_));
  NAi31      o112(.An(i_9_), .B(i_6_), .C(i_5_), .Y(ori_ori_n135_));
  INV        o113(.A(i_13_), .Y(ori_ori_n136_));
  NO2        o114(.A(i_12_), .B(ori_ori_n136_), .Y(ori_ori_n137_));
  INV        o115(.A(i_12_), .Y(ori_ori_n138_));
  NO2        o116(.A(ori_ori_n42_), .B(ori_ori_n138_), .Y(ori_ori_n139_));
  NO3        o117(.A(ori_ori_n35_), .B(i_8_), .C(i_10_), .Y(ori_ori_n140_));
  NA2        o118(.A(i_2_), .B(i_1_), .Y(ori_ori_n141_));
  NO3        o119(.A(i_11_), .B(i_7_), .C(ori_ori_n36_), .Y(ori_ori_n142_));
  NAi21      o120(.An(i_4_), .B(i_3_), .Y(ori_ori_n143_));
  NOi41      o121(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(ori_ori_n144_));
  NO2        o122(.A(i_11_), .B(ori_ori_n136_), .Y(ori_ori_n145_));
  NOi21      o123(.An(i_1_), .B(i_6_), .Y(ori_ori_n146_));
  NAi21      o124(.An(i_3_), .B(i_7_), .Y(ori_ori_n147_));
  NA2        o125(.A(ori_ori_n138_), .B(i_9_), .Y(ori_ori_n148_));
  OR4        o126(.A(ori_ori_n148_), .B(ori_ori_n147_), .C(ori_ori_n146_), .D(ori_ori_n125_), .Y(ori_ori_n149_));
  NA2        o127(.A(ori_ori_n63_), .B(i_5_), .Y(ori_ori_n150_));
  NA2        o128(.A(i_3_), .B(i_9_), .Y(ori_ori_n151_));
  NAi21      o129(.An(i_7_), .B(i_10_), .Y(ori_ori_n152_));
  NO2        o130(.A(ori_ori_n152_), .B(ori_ori_n151_), .Y(ori_ori_n153_));
  NA3        o131(.A(ori_ori_n153_), .B(ori_ori_n150_), .C(ori_ori_n55_), .Y(ori_ori_n154_));
  NA2        o132(.A(ori_ori_n154_), .B(ori_ori_n149_), .Y(ori_ori_n155_));
  INV        o133(.A(ori_ori_n113_), .Y(ori_ori_n156_));
  NA2        o134(.A(ori_ori_n138_), .B(i_13_), .Y(ori_ori_n157_));
  NO2        o135(.A(ori_ori_n157_), .B(ori_ori_n64_), .Y(ori_ori_n158_));
  AOI220     o136(.A0(ori_ori_n158_), .A1(ori_ori_n156_), .B0(ori_ori_n155_), .B1(ori_ori_n145_), .Y(ori_ori_n159_));
  NA2        o137(.A(i_12_), .B(i_6_), .Y(ori_ori_n160_));
  OR2        o138(.A(i_13_), .B(i_9_), .Y(ori_ori_n161_));
  NO2        o139(.A(ori_ori_n143_), .B(i_2_), .Y(ori_ori_n162_));
  NA2        o140(.A(ori_ori_n145_), .B(i_9_), .Y(ori_ori_n163_));
  NO3        o141(.A(i_12_), .B(ori_ori_n136_), .C(ori_ori_n36_), .Y(ori_ori_n164_));
  AN2        o142(.A(i_3_), .B(i_10_), .Y(ori_ori_n165_));
  NO2        o143(.A(i_5_), .B(ori_ori_n36_), .Y(ori_ori_n166_));
  NO2        o144(.A(ori_ori_n44_), .B(ori_ori_n26_), .Y(ori_ori_n167_));
  NO3        o145(.A(ori_ori_n42_), .B(i_13_), .C(i_9_), .Y(ori_ori_n168_));
  NO2        o146(.A(i_2_), .B(i_3_), .Y(ori_ori_n169_));
  NO2        o147(.A(i_12_), .B(i_10_), .Y(ori_ori_n170_));
  NO2        o148(.A(i_1_), .B(i_7_), .Y(ori_ori_n171_));
  NOi21      o149(.An(ori_ori_n118_), .B(ori_ori_n88_), .Y(ori_ori_n172_));
  NO2        o150(.A(ori_ori_n172_), .B(ori_ori_n99_), .Y(ori_ori_n173_));
  NA2        o151(.A(ori_ori_n173_), .B(i_3_), .Y(ori_ori_n174_));
  NO2        o152(.A(ori_ori_n128_), .B(i_9_), .Y(ori_ori_n175_));
  NA2        o153(.A(ori_ori_n175_), .B(ori_ori_n131_), .Y(ori_ori_n176_));
  NO2        o154(.A(ori_ori_n176_), .B(ori_ori_n44_), .Y(ori_ori_n177_));
  INV        o155(.A(ori_ori_n177_), .Y(ori_ori_n178_));
  AOI210     o156(.A0(ori_ori_n178_), .A1(ori_ori_n174_), .B0(ori_ori_n121_), .Y(ori_ori_n179_));
  INV        o157(.A(ori_ori_n179_), .Y(ori_ori_n180_));
  NOi32      o158(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(ori_ori_n181_));
  INV        o159(.A(ori_ori_n181_), .Y(ori_ori_n182_));
  NOi32      o160(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(ori_ori_n183_));
  NO2        o161(.A(i_1_), .B(ori_ori_n85_), .Y(ori_ori_n184_));
  NAi21      o162(.An(i_3_), .B(i_4_), .Y(ori_ori_n185_));
  NO2        o163(.A(ori_ori_n185_), .B(i_9_), .Y(ori_ori_n186_));
  AN2        o164(.A(i_6_), .B(i_7_), .Y(ori_ori_n187_));
  OAI210     o165(.A0(ori_ori_n187_), .A1(ori_ori_n184_), .B0(ori_ori_n186_), .Y(ori_ori_n188_));
  NO2        o166(.A(ori_ori_n185_), .B(i_10_), .Y(ori_ori_n189_));
  NO2        o167(.A(ori_ori_n188_), .B(ori_ori_n125_), .Y(ori_ori_n190_));
  AOI220     o168(.A0(ori_ori_n189_), .A1(ori_ori_n171_), .B0(ori_ori_n140_), .B1(ori_ori_n126_), .Y(ori_ori_n191_));
  NO2        o169(.A(ori_ori_n191_), .B(i_5_), .Y(ori_ori_n192_));
  NO2        o170(.A(ori_ori_n192_), .B(ori_ori_n190_), .Y(ori_ori_n193_));
  NO2        o171(.A(ori_ori_n193_), .B(ori_ori_n182_), .Y(ori_ori_n194_));
  AN2        o172(.A(i_12_), .B(i_5_), .Y(ori_ori_n195_));
  NO2        o173(.A(i_11_), .B(i_6_), .Y(ori_ori_n196_));
  NO2        o174(.A(i_5_), .B(i_10_), .Y(ori_ori_n197_));
  NO2        o175(.A(ori_ori_n36_), .B(ori_ori_n25_), .Y(ori_ori_n198_));
  NO3        o176(.A(i_1_), .B(i_12_), .C(ori_ori_n72_), .Y(ori_ori_n199_));
  NO2        o177(.A(i_0_), .B(i_11_), .Y(ori_ori_n200_));
  BUFFER     o178(.A(i_6_), .Y(ori_ori_n201_));
  NAi21      o179(.An(i_9_), .B(i_4_), .Y(ori_ori_n202_));
  OR2        o180(.A(i_13_), .B(i_10_), .Y(ori_ori_n203_));
  NO3        o181(.A(ori_ori_n203_), .B(ori_ori_n96_), .C(ori_ori_n202_), .Y(ori_ori_n204_));
  NO2        o182(.A(ori_ori_n85_), .B(ori_ori_n25_), .Y(ori_ori_n205_));
  NA2        o183(.A(ori_ori_n164_), .B(ori_ori_n205_), .Y(ori_ori_n206_));
  NO2        o184(.A(ori_ori_n206_), .B(ori_ori_n172_), .Y(ori_ori_n207_));
  NA2        o185(.A(ori_ori_n128_), .B(i_10_), .Y(ori_ori_n208_));
  NA3        o186(.A(ori_ori_n150_), .B(ori_ori_n55_), .C(i_2_), .Y(ori_ori_n209_));
  NO2        o187(.A(ori_ori_n209_), .B(ori_ori_n208_), .Y(ori_ori_n210_));
  INV        o188(.A(ori_ori_n210_), .Y(ori_ori_n211_));
  NO2        o189(.A(ori_ori_n211_), .B(ori_ori_n163_), .Y(ori_ori_n212_));
  NO3        o190(.A(ori_ori_n212_), .B(ori_ori_n207_), .C(ori_ori_n194_), .Y(ori_ori_n213_));
  NO2        o191(.A(ori_ori_n63_), .B(i_13_), .Y(ori_ori_n214_));
  NO3        o192(.A(ori_ori_n23_), .B(i_10_), .C(i_9_), .Y(ori_ori_n215_));
  NA2        o193(.A(ori_ori_n160_), .B(ori_ori_n84_), .Y(ori_ori_n216_));
  NA2        o194(.A(i_8_), .B(i_9_), .Y(ori_ori_n217_));
  NO2        o195(.A(i_7_), .B(i_2_), .Y(ori_ori_n218_));
  OR2        o196(.A(ori_ori_n218_), .B(ori_ori_n217_), .Y(ori_ori_n219_));
  NA2        o197(.A(ori_ori_n164_), .B(ori_ori_n131_), .Y(ori_ori_n220_));
  NO2        o198(.A(ori_ori_n220_), .B(ori_ori_n219_), .Y(ori_ori_n221_));
  NA2        o199(.A(ori_ori_n145_), .B(ori_ori_n166_), .Y(ori_ori_n222_));
  NO3        o200(.A(i_6_), .B(i_8_), .C(i_7_), .Y(ori_ori_n223_));
  INV        o201(.A(ori_ori_n223_), .Y(ori_ori_n224_));
  NA3        o202(.A(i_2_), .B(i_10_), .C(i_9_), .Y(ori_ori_n225_));
  NA4        o203(.A(ori_ori_n115_), .B(ori_ori_n95_), .C(ori_ori_n68_), .D(ori_ori_n23_), .Y(ori_ori_n226_));
  OAI220     o204(.A0(ori_ori_n226_), .A1(ori_ori_n225_), .B0(ori_ori_n224_), .B1(ori_ori_n222_), .Y(ori_ori_n227_));
  NO2        o205(.A(ori_ori_n227_), .B(ori_ori_n221_), .Y(ori_ori_n228_));
  NA2        o206(.A(ori_ori_n83_), .B(i_13_), .Y(ori_ori_n229_));
  NO2        o207(.A(i_11_), .B(i_1_), .Y(ori_ori_n230_));
  NA3        o208(.A(ori_ori_n144_), .B(ori_ori_n123_), .C(ori_ori_n105_), .Y(ori_ori_n231_));
  NA2        o209(.A(ori_ori_n44_), .B(ori_ori_n42_), .Y(ori_ori_n232_));
  NO2        o210(.A(ori_ori_n119_), .B(i_3_), .Y(ori_ori_n233_));
  NAi31      o211(.An(ori_ori_n232_), .B(ori_ori_n233_), .C(ori_ori_n137_), .Y(ori_ori_n234_));
  NA2        o212(.A(ori_ori_n234_), .B(ori_ori_n231_), .Y(ori_ori_n235_));
  INV        o213(.A(ori_ori_n235_), .Y(ori_ori_n236_));
  NA2        o214(.A(ori_ori_n215_), .B(ori_ori_n195_), .Y(ori_ori_n237_));
  NA2        o215(.A(ori_ori_n223_), .B(ori_ori_n197_), .Y(ori_ori_n238_));
  NA2        o216(.A(ori_ori_n27_), .B(i_10_), .Y(ori_ori_n239_));
  NA2        o217(.A(ori_ori_n168_), .B(ori_ori_n140_), .Y(ori_ori_n240_));
  OAI220     o218(.A0(ori_ori_n240_), .A1(ori_ori_n209_), .B0(ori_ori_n239_), .B1(ori_ori_n229_), .Y(ori_ori_n241_));
  INV        o219(.A(ori_ori_n241_), .Y(ori_ori_n242_));
  NA3        o220(.A(ori_ori_n242_), .B(ori_ori_n236_), .C(ori_ori_n228_), .Y(ori_ori_n243_));
  NA2        o221(.A(ori_ori_n195_), .B(ori_ori_n136_), .Y(ori_ori_n244_));
  NA2        o222(.A(ori_ori_n187_), .B(ori_ori_n183_), .Y(ori_ori_n245_));
  OR2        o223(.A(ori_ori_n244_), .B(ori_ori_n245_), .Y(ori_ori_n246_));
  AOI210     o224(.A0(ori_ori_n38_), .A1(i_13_), .B0(ori_ori_n204_), .Y(ori_ori_n247_));
  NA2        o225(.A(ori_ori_n247_), .B(ori_ori_n246_), .Y(ori_ori_n248_));
  NA3        o226(.A(ori_ori_n134_), .B(ori_ori_n61_), .C(ori_ori_n42_), .Y(ori_ori_n249_));
  NA2        o227(.A(ori_ori_n164_), .B(ori_ori_n70_), .Y(ori_ori_n250_));
  NO2        o228(.A(ori_ori_n249_), .B(ori_ori_n250_), .Y(ori_ori_n251_));
  NO2        o229(.A(ori_ori_n203_), .B(i_1_), .Y(ori_ori_n252_));
  NOi31      o230(.An(ori_ori_n252_), .B(ori_ori_n216_), .C(ori_ori_n63_), .Y(ori_ori_n253_));
  NOi21      o231(.An(i_10_), .B(i_6_), .Y(ori_ori_n254_));
  OR2        o232(.A(i_2_), .B(i_5_), .Y(ori_ori_n255_));
  NO3        o233(.A(ori_ori_n251_), .B(ori_ori_n248_), .C(ori_ori_n243_), .Y(ori_ori_n256_));
  NA4        o234(.A(ori_ori_n256_), .B(ori_ori_n213_), .C(ori_ori_n180_), .D(ori_ori_n159_), .Y(ori7));
  NO2        o235(.A(ori_ori_n79_), .B(ori_ori_n49_), .Y(ori_ori_n258_));
  INV        o236(.A(i_11_), .Y(ori_ori_n259_));
  NA3        o237(.A(i_7_), .B(i_10_), .C(i_9_), .Y(ori_ori_n260_));
  NO2        o238(.A(ori_ori_n138_), .B(i_4_), .Y(ori_ori_n261_));
  NA2        o239(.A(ori_ori_n261_), .B(i_8_), .Y(ori_ori_n262_));
  NO2        o240(.A(ori_ori_n89_), .B(ori_ori_n260_), .Y(ori_ori_n263_));
  NA2        o241(.A(i_2_), .B(ori_ori_n72_), .Y(ori_ori_n264_));
  OAI210     o242(.A0(ori_ori_n73_), .A1(ori_ori_n129_), .B0(ori_ori_n130_), .Y(ori_ori_n265_));
  INV        o243(.A(ori_ori_n165_), .Y(ori_ori_n266_));
  OAI220     o244(.A0(ori_ori_n266_), .A1(ori_ori_n264_), .B0(ori_ori_n265_), .B1(i_13_), .Y(ori_ori_n267_));
  NO3        o245(.A(ori_ori_n267_), .B(ori_ori_n263_), .C(ori_ori_n258_), .Y(ori_ori_n268_));
  AOI210     o246(.A0(ori_ori_n103_), .A1(ori_ori_n53_), .B0(i_10_), .Y(ori_ori_n269_));
  AOI210     o247(.A0(ori_ori_n269_), .A1(ori_ori_n138_), .B0(ori_ori_n120_), .Y(ori_ori_n270_));
  OR2        o248(.A(i_6_), .B(i_10_), .Y(ori_ori_n271_));
  OR3        o249(.A(i_13_), .B(i_6_), .C(i_10_), .Y(ori_ori_n272_));
  OR2        o250(.A(ori_ori_n270_), .B(ori_ori_n161_), .Y(ori_ori_n273_));
  AOI210     o251(.A0(ori_ori_n273_), .A1(ori_ori_n268_), .B0(ori_ori_n54_), .Y(ori_ori_n274_));
  NOi21      o252(.An(i_11_), .B(i_7_), .Y(ori_ori_n275_));
  AO210      o253(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(ori_ori_n276_));
  NO2        o254(.A(ori_ori_n276_), .B(ori_ori_n275_), .Y(ori_ori_n277_));
  NA2        o255(.A(ori_ori_n277_), .B(ori_ori_n132_), .Y(ori_ori_n278_));
  NA3        o256(.A(i_3_), .B(i_8_), .C(i_9_), .Y(ori_ori_n279_));
  NO2        o257(.A(ori_ori_n278_), .B(ori_ori_n54_), .Y(ori_ori_n280_));
  OR2        o258(.A(ori_ori_n191_), .B(ori_ori_n40_), .Y(ori_ori_n281_));
  NA2        o259(.A(ori_ori_n137_), .B(ori_ori_n54_), .Y(ori_ori_n282_));
  NO2        o260(.A(i_1_), .B(i_12_), .Y(ori_ori_n283_));
  NA2        o261(.A(ori_ori_n282_), .B(ori_ori_n281_), .Y(ori_ori_n284_));
  OAI210     o262(.A0(ori_ori_n284_), .A1(ori_ori_n280_), .B0(i_6_), .Y(ori_ori_n285_));
  NO2        o263(.A(ori_ori_n279_), .B(ori_ori_n92_), .Y(ori_ori_n286_));
  NO3        o264(.A(ori_ori_n271_), .B(i_7_), .C(ori_ori_n23_), .Y(ori_ori_n287_));
  AOI210     o265(.A0(i_1_), .A1(ori_ori_n153_), .B0(ori_ori_n287_), .Y(ori_ori_n288_));
  NO2        o266(.A(ori_ori_n288_), .B(ori_ori_n42_), .Y(ori_ori_n289_));
  INV        o267(.A(i_2_), .Y(ori_ori_n290_));
  NA2        o268(.A(ori_ori_n108_), .B(i_9_), .Y(ori_ori_n291_));
  NO2        o269(.A(ori_ori_n291_), .B(ori_ori_n290_), .Y(ori_ori_n292_));
  AOI210     o270(.A0(ori_ori_n230_), .A1(ori_ori_n205_), .B0(ori_ori_n142_), .Y(ori_ori_n293_));
  NO2        o271(.A(ori_ori_n293_), .B(ori_ori_n264_), .Y(ori_ori_n294_));
  OR2        o272(.A(ori_ori_n294_), .B(ori_ori_n292_), .Y(ori_ori_n295_));
  NO3        o273(.A(ori_ori_n295_), .B(ori_ori_n289_), .C(ori_ori_n286_), .Y(ori_ori_n296_));
  NO2        o274(.A(ori_ori_n138_), .B(ori_ori_n85_), .Y(ori_ori_n297_));
  NO2        o275(.A(ori_ori_n297_), .B(ori_ori_n275_), .Y(ori_ori_n298_));
  NA2        o276(.A(ori_ori_n298_), .B(i_1_), .Y(ori_ori_n299_));
  NO2        o277(.A(ori_ori_n299_), .B(ori_ori_n272_), .Y(ori_ori_n300_));
  NO2        o278(.A(ori_ori_n202_), .B(ori_ori_n72_), .Y(ori_ori_n301_));
  NA2        o279(.A(ori_ori_n300_), .B(ori_ori_n44_), .Y(ori_ori_n302_));
  NO2        o280(.A(i_7_), .B(ori_ori_n42_), .Y(ori_ori_n303_));
  NO3        o281(.A(ori_ori_n303_), .B(ori_ori_n167_), .C(ori_ori_n139_), .Y(ori_ori_n304_));
  NO2        o282(.A(ori_ori_n96_), .B(ori_ori_n36_), .Y(ori_ori_n305_));
  NO2        o283(.A(ori_ori_n305_), .B(i_6_), .Y(ori_ori_n306_));
  NO2        o284(.A(ori_ori_n72_), .B(i_9_), .Y(ori_ori_n307_));
  NO2        o285(.A(ori_ori_n307_), .B(ori_ori_n54_), .Y(ori_ori_n308_));
  NO2        o286(.A(ori_ori_n308_), .B(ori_ori_n283_), .Y(ori_ori_n309_));
  NO4        o287(.A(ori_ori_n309_), .B(ori_ori_n306_), .C(ori_ori_n304_), .D(i_4_), .Y(ori_ori_n310_));
  INV        o288(.A(ori_ori_n310_), .Y(ori_ori_n311_));
  NA4        o289(.A(ori_ori_n311_), .B(ori_ori_n302_), .C(ori_ori_n296_), .D(ori_ori_n285_), .Y(ori_ori_n312_));
  INV        o290(.A(i_1_), .Y(ori_ori_n313_));
  OR2        o291(.A(i_11_), .B(i_7_), .Y(ori_ori_n314_));
  NO2        o292(.A(ori_ori_n49_), .B(i_12_), .Y(ori_ori_n315_));
  INV        o293(.A(ori_ori_n315_), .Y(ori_ori_n316_));
  NA2        o294(.A(i_7_), .B(ori_ori_n301_), .Y(ori_ori_n317_));
  OAI220     o295(.A0(ori_ori_n317_), .A1(ori_ori_n40_), .B0(ori_ori_n316_), .B1(ori_ori_n79_), .Y(ori_ori_n318_));
  INV        o296(.A(ori_ori_n318_), .Y(ori_ori_n319_));
  NA2        o297(.A(ori_ori_n102_), .B(i_13_), .Y(ori_ori_n320_));
  NO2        o298(.A(ori_ori_n320_), .B(ori_ori_n313_), .Y(ori_ori_n321_));
  INV        o299(.A(i_7_), .Y(ori_ori_n322_));
  AOI220     o300(.A0(ori_ori_n196_), .A1(ori_ori_n454_), .B0(ori_ori_n78_), .B1(ori_ori_n86_), .Y(ori_ori_n323_));
  NO2        o301(.A(ori_ori_n323_), .B(ori_ori_n262_), .Y(ori_ori_n324_));
  NO2        o302(.A(ori_ori_n324_), .B(ori_ori_n321_), .Y(ori_ori_n325_));
  OR2        o303(.A(i_11_), .B(i_6_), .Y(ori_ori_n326_));
  NA2        o304(.A(ori_ori_n261_), .B(i_7_), .Y(ori_ori_n327_));
  NO2        o305(.A(ori_ori_n327_), .B(ori_ori_n326_), .Y(ori_ori_n328_));
  NA2        o306(.A(ori_ori_n328_), .B(ori_ori_n54_), .Y(ori_ori_n329_));
  NO2        o307(.A(i_2_), .B(i_12_), .Y(ori_ori_n330_));
  NA2        o308(.A(ori_ori_n184_), .B(ori_ori_n330_), .Y(ori_ori_n331_));
  NA2        o309(.A(ori_ori_n186_), .B(ori_ori_n184_), .Y(ori_ori_n332_));
  NA2        o310(.A(ori_ori_n332_), .B(ori_ori_n331_), .Y(ori_ori_n333_));
  NA2        o311(.A(ori_ori_n333_), .B(ori_ori_n43_), .Y(ori_ori_n334_));
  NA4        o312(.A(ori_ori_n334_), .B(ori_ori_n329_), .C(ori_ori_n325_), .D(ori_ori_n319_), .Y(ori_ori_n335_));
  OR3        o313(.A(ori_ori_n335_), .B(ori_ori_n312_), .C(ori_ori_n274_), .Y(ori5));
  NA2        o314(.A(ori_ori_n298_), .B(ori_ori_n162_), .Y(ori_ori_n337_));
  NA3        o315(.A(ori_ori_n24_), .B(ori_ori_n330_), .C(ori_ori_n92_), .Y(ori_ori_n338_));
  NO2        o316(.A(ori_ori_n262_), .B(i_11_), .Y(ori_ori_n339_));
  NA2        o317(.A(ori_ori_n73_), .B(ori_ori_n339_), .Y(ori_ori_n340_));
  NA3        o318(.A(ori_ori_n340_), .B(ori_ori_n338_), .C(ori_ori_n337_), .Y(ori_ori_n341_));
  NO2        o319(.A(ori_ori_n99_), .B(ori_ori_n23_), .Y(ori_ori_n342_));
  NO2        o320(.A(ori_ori_n342_), .B(ori_ori_n341_), .Y(ori_ori_n343_));
  INV        o321(.A(ori_ori_n123_), .Y(ori_ori_n344_));
  INV        o322(.A(ori_ori_n144_), .Y(ori_ori_n345_));
  NO2        o323(.A(ori_ori_n345_), .B(ori_ori_n344_), .Y(ori_ori_n346_));
  INV        o324(.A(ori_ori_n346_), .Y(ori_ori_n347_));
  NO3        o325(.A(ori_ori_n276_), .B(ori_ori_n37_), .C(ori_ori_n26_), .Y(ori_ori_n348_));
  OA210      o326(.A0(ori_ori_n277_), .A1(ori_ori_n101_), .B0(i_13_), .Y(ori_ori_n349_));
  NA3        o327(.A(i_2_), .B(ori_ori_n165_), .C(ori_ori_n99_), .Y(ori_ori_n350_));
  NO4        o328(.A(ori_ori_n453_), .B(ori_ori_n117_), .C(ori_ori_n349_), .D(ori_ori_n348_), .Y(ori_ori_n351_));
  NO2        o329(.A(ori_ori_n53_), .B(i_12_), .Y(ori_ori_n352_));
  NO2        o330(.A(ori_ori_n352_), .B(ori_ori_n101_), .Y(ori_ori_n353_));
  NO2        o331(.A(ori_ori_n353_), .B(ori_ori_n259_), .Y(ori_ori_n354_));
  NA2        o332(.A(ori_ori_n354_), .B(ori_ori_n35_), .Y(ori_ori_n355_));
  NA4        o333(.A(ori_ori_n355_), .B(ori_ori_n351_), .C(ori_ori_n347_), .D(ori_ori_n343_), .Y(ori6));
  NO2        o334(.A(ori_ori_n135_), .B(ori_ori_n232_), .Y(ori_ori_n357_));
  INV        o335(.A(ori_ori_n170_), .Y(ori_ori_n358_));
  NA2        o336(.A(ori_ori_n64_), .B(ori_ori_n104_), .Y(ori_ori_n359_));
  NO2        o337(.A(ori_ori_n359_), .B(ori_ori_n358_), .Y(ori_ori_n360_));
  NO2        o338(.A(ori_ori_n146_), .B(i_9_), .Y(ori_ori_n361_));
  NA2        o339(.A(ori_ori_n361_), .B(ori_ori_n352_), .Y(ori_ori_n362_));
  AOI210     o340(.A0(ori_ori_n362_), .A1(ori_ori_n245_), .B0(ori_ori_n125_), .Y(ori_ori_n363_));
  NAi32      o341(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(ori_ori_n364_));
  NO2        o342(.A(ori_ori_n326_), .B(ori_ori_n364_), .Y(ori_ori_n365_));
  OR3        o343(.A(ori_ori_n365_), .B(ori_ori_n363_), .C(ori_ori_n360_), .Y(ori_ori_n366_));
  NO2        o344(.A(ori_ori_n314_), .B(i_2_), .Y(ori_ori_n367_));
  BUFFER     o345(.A(ori_ori_n277_), .Y(ori_ori_n368_));
  NA2        o346(.A(ori_ori_n368_), .B(ori_ori_n116_), .Y(ori_ori_n369_));
  OR2        o347(.A(ori_ori_n238_), .B(ori_ori_n35_), .Y(ori_ori_n370_));
  NA2        o348(.A(ori_ori_n370_), .B(ori_ori_n369_), .Y(ori_ori_n371_));
  NA2        o349(.A(ori_ori_n357_), .B(ori_ori_n322_), .Y(ori_ori_n372_));
  NA2        o350(.A(ori_ori_n372_), .B(ori_ori_n265_), .Y(ori_ori_n373_));
  NO2        o351(.A(ori_ori_n271_), .B(ori_ori_n86_), .Y(ori_ori_n374_));
  OAI210     o352(.A0(ori_ori_n374_), .A1(ori_ori_n94_), .B0(ori_ori_n200_), .Y(ori_ori_n375_));
  NA3        o353(.A(ori_ori_n452_), .B(ori_ori_n170_), .C(i_7_), .Y(ori_ori_n376_));
  NA2        o354(.A(ori_ori_n376_), .B(ori_ori_n375_), .Y(ori_ori_n377_));
  NO4        o355(.A(ori_ori_n377_), .B(ori_ori_n373_), .C(ori_ori_n371_), .D(ori_ori_n366_), .Y(ori_ori_n378_));
  NA2        o356(.A(ori_ori_n378_), .B(ori_ori_n193_), .Y(ori3));
  NA2        o357(.A(i_12_), .B(i_10_), .Y(ori_ori_n380_));
  NO2        o358(.A(i_11_), .B(ori_ori_n138_), .Y(ori_ori_n381_));
  NA2        o359(.A(ori_ori_n265_), .B(ori_ori_n188_), .Y(ori_ori_n382_));
  NA2        o360(.A(ori_ori_n382_), .B(ori_ori_n39_), .Y(ori_ori_n383_));
  NOi21      o361(.An(ori_ori_n83_), .B(ori_ori_n25_), .Y(ori_ori_n384_));
  AN2        o362(.A(ori_ori_n216_), .B(ori_ori_n50_), .Y(ori_ori_n385_));
  NO2        o363(.A(ori_ori_n385_), .B(ori_ori_n384_), .Y(ori_ori_n386_));
  AOI210     o364(.A0(ori_ori_n386_), .A1(ori_ori_n383_), .B0(ori_ori_n45_), .Y(ori_ori_n387_));
  NO3        o365(.A(ori_ori_n195_), .B(ori_ori_n37_), .C(i_0_), .Y(ori_ori_n388_));
  NA2        o366(.A(ori_ori_n125_), .B(ori_ori_n254_), .Y(ori_ori_n389_));
  NOi21      o367(.An(ori_ori_n389_), .B(ori_ori_n388_), .Y(ori_ori_n390_));
  NO2        o368(.A(ori_ori_n390_), .B(ori_ori_n54_), .Y(ori_ori_n391_));
  NOi21      o369(.An(i_5_), .B(i_9_), .Y(ori_ori_n392_));
  NA2        o370(.A(ori_ori_n392_), .B(ori_ori_n214_), .Y(ori_ori_n393_));
  BUFFER     o371(.A(ori_ori_n160_), .Y(ori_ori_n394_));
  NA2        o372(.A(ori_ori_n394_), .B(ori_ori_n230_), .Y(ori_ori_n395_));
  NO2        o373(.A(ori_ori_n395_), .B(ori_ori_n393_), .Y(ori_ori_n396_));
  NO3        o374(.A(ori_ori_n396_), .B(ori_ori_n391_), .C(ori_ori_n387_), .Y(ori_ori_n397_));
  NO4        o375(.A(ori_ori_n255_), .B(i_12_), .C(ori_ori_n203_), .D(ori_ori_n201_), .Y(ori_ori_n398_));
  NA2        o376(.A(ori_ori_n398_), .B(i_11_), .Y(ori_ori_n399_));
  NO2        o377(.A(ori_ori_n148_), .B(ori_ori_n118_), .Y(ori_ori_n400_));
  NA2        o378(.A(i_0_), .B(i_10_), .Y(ori_ori_n401_));
  AN2        o379(.A(ori_ori_n400_), .B(i_6_), .Y(ori_ori_n402_));
  INV        o380(.A(ori_ori_n402_), .Y(ori_ori_n403_));
  NA2        o381(.A(ori_ori_n403_), .B(ori_ori_n399_), .Y(ori_ori_n404_));
  NA2        o382(.A(i_11_), .B(i_9_), .Y(ori_ori_n405_));
  NO3        o383(.A(i_12_), .B(ori_ori_n405_), .C(ori_ori_n264_), .Y(ori_ori_n406_));
  AN2        o384(.A(ori_ori_n406_), .B(i_5_), .Y(ori_ori_n407_));
  NA2        o385(.A(ori_ori_n198_), .B(ori_ori_n124_), .Y(ori_ori_n408_));
  INV        o386(.A(ori_ori_n408_), .Y(ori_ori_n409_));
  NO2        o387(.A(ori_ori_n405_), .B(ori_ori_n63_), .Y(ori_ori_n410_));
  INV        o388(.A(ori_ori_n199_), .Y(ori_ori_n411_));
  NO2        o389(.A(ori_ori_n411_), .B(ori_ori_n393_), .Y(ori_ori_n412_));
  NO3        o390(.A(ori_ori_n412_), .B(ori_ori_n409_), .C(ori_ori_n407_), .Y(ori_ori_n413_));
  INV        o391(.A(ori_ori_n413_), .Y(ori_ori_n414_));
  NO2        o392(.A(ori_ori_n380_), .B(ori_ori_n169_), .Y(ori_ori_n415_));
  NA2        o393(.A(ori_ori_n415_), .B(ori_ori_n410_), .Y(ori_ori_n416_));
  NA2        o394(.A(ori_ori_n246_), .B(ori_ori_n416_), .Y(ori_ori_n417_));
  NO3        o395(.A(ori_ori_n417_), .B(ori_ori_n414_), .C(ori_ori_n404_), .Y(ori_ori_n418_));
  NO3        o396(.A(ori_ori_n401_), .B(ori_ori_n392_), .C(ori_ori_n127_), .Y(ori_ori_n419_));
  AOI220     o397(.A0(ori_ori_n419_), .A1(i_11_), .B0(ori_ori_n253_), .B1(ori_ori_n64_), .Y(ori_ori_n420_));
  NO3        o398(.A(ori_ori_n133_), .B(ori_ori_n195_), .C(i_0_), .Y(ori_ori_n421_));
  NA2        o399(.A(ori_ori_n421_), .B(i_13_), .Y(ori_ori_n422_));
  NA2        o400(.A(ori_ori_n422_), .B(ori_ori_n420_), .Y(ori_ori_n423_));
  NA2        o401(.A(ori_ori_n237_), .B(ori_ori_n231_), .Y(ori_ori_n424_));
  INV        o402(.A(ori_ori_n424_), .Y(ori_ori_n425_));
  NA3        o403(.A(ori_ori_n197_), .B(ori_ori_n123_), .C(ori_ori_n122_), .Y(ori_ori_n426_));
  INV        o404(.A(ori_ori_n426_), .Y(ori_ori_n427_));
  NO3        o405(.A(ori_ori_n405_), .B(ori_ori_n134_), .C(ori_ori_n127_), .Y(ori_ori_n428_));
  NO2        o406(.A(ori_ori_n428_), .B(ori_ori_n427_), .Y(ori_ori_n429_));
  NA2        o407(.A(ori_ori_n429_), .B(ori_ori_n425_), .Y(ori_ori_n430_));
  NO2        o408(.A(ori_ori_n72_), .B(i_5_), .Y(ori_ori_n431_));
  NA2        o409(.A(ori_ori_n381_), .B(ori_ori_n93_), .Y(ori_ori_n432_));
  INV        o410(.A(ori_ori_n432_), .Y(ori_ori_n433_));
  NA2        o411(.A(ori_ori_n433_), .B(ori_ori_n431_), .Y(ori_ori_n434_));
  NAi21      o412(.An(ori_ori_n142_), .B(ori_ori_n143_), .Y(ori_ori_n435_));
  NO4        o413(.A(ori_ori_n141_), .B(ori_ori_n133_), .C(i_0_), .D(i_12_), .Y(ori_ori_n436_));
  NA2        o414(.A(ori_ori_n436_), .B(ori_ori_n435_), .Y(ori_ori_n437_));
  NA2        o415(.A(ori_ori_n437_), .B(ori_ori_n434_), .Y(ori_ori_n438_));
  NO3        o416(.A(ori_ori_n438_), .B(ori_ori_n430_), .C(ori_ori_n423_), .Y(ori_ori_n439_));
  NA2        o417(.A(ori_ori_n367_), .B(ori_ori_n36_), .Y(ori_ori_n440_));
  NA2        o418(.A(ori_ori_n440_), .B(ori_ori_n270_), .Y(ori_ori_n441_));
  NA2        o419(.A(ori_ori_n441_), .B(ori_ori_n132_), .Y(ori_ori_n442_));
  NA2        o420(.A(i_2_), .B(i_10_), .Y(ori_ori_n443_));
  NO2        o421(.A(ori_ori_n60_), .B(ori_ori_n443_), .Y(ori_ori_n444_));
  AOI210     o422(.A0(ori_ori_n444_), .A1(ori_ori_n45_), .B0(ori_ori_n398_), .Y(ori_ori_n445_));
  AOI210     o423(.A0(ori_ori_n445_), .A1(ori_ori_n442_), .B0(ori_ori_n63_), .Y(ori_ori_n446_));
  NO2        o424(.A(ori_ori_n191_), .B(ori_ori_n344_), .Y(ori_ori_n447_));
  NO2        o425(.A(ori_ori_n447_), .B(ori_ori_n446_), .Y(ori_ori_n448_));
  NA4        o426(.A(ori_ori_n448_), .B(ori_ori_n439_), .C(ori_ori_n418_), .D(ori_ori_n397_), .Y(ori4));
  INV        o427(.A(ori_ori_n255_), .Y(ori_ori_n452_));
  INV        o428(.A(ori_ori_n350_), .Y(ori_ori_n453_));
  INV        o429(.A(i_1_), .Y(ori_ori_n454_));
  NAi21      m000(.An(i_13_), .B(i_4_), .Y(mai_mai_n23_));
  NOi21      m001(.An(i_3_), .B(i_8_), .Y(mai_mai_n24_));
  INV        m002(.A(i_9_), .Y(mai_mai_n25_));
  INV        m003(.A(i_3_), .Y(mai_mai_n26_));
  NO2        m004(.A(mai_mai_n26_), .B(mai_mai_n25_), .Y(mai_mai_n27_));
  NO2        m005(.A(i_8_), .B(i_10_), .Y(mai_mai_n28_));
  INV        m006(.A(mai_mai_n28_), .Y(mai_mai_n29_));
  OAI210     m007(.A0(mai_mai_n27_), .A1(mai_mai_n24_), .B0(mai_mai_n29_), .Y(mai_mai_n30_));
  NOi21      m008(.An(i_11_), .B(i_8_), .Y(mai_mai_n31_));
  AO210      m009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(mai_mai_n32_));
  OR2        m010(.A(mai_mai_n32_), .B(mai_mai_n31_), .Y(mai_mai_n33_));
  NA2        m011(.A(mai_mai_n33_), .B(mai_mai_n30_), .Y(mai_mai_n34_));
  XO2        m012(.A(mai_mai_n34_), .B(mai_mai_n23_), .Y(mai_mai_n35_));
  INV        m013(.A(i_4_), .Y(mai_mai_n36_));
  INV        m014(.A(i_10_), .Y(mai_mai_n37_));
  NO3        m015(.A(i_11_), .B(i_12_), .C(mai_mai_n37_), .Y(mai_mai_n38_));
  NOi21      m016(.An(i_12_), .B(i_13_), .Y(mai_mai_n39_));
  INV        m017(.A(mai_mai_n39_), .Y(mai_mai_n40_));
  NO2        m018(.A(mai_mai_n36_), .B(i_3_), .Y(mai_mai_n41_));
  NAi31      m019(.An(i_9_), .B(i_4_), .C(i_8_), .Y(mai_mai_n42_));
  INV        m020(.A(mai_mai_n35_), .Y(mai1));
  INV        m021(.A(i_11_), .Y(mai_mai_n44_));
  NO2        m022(.A(mai_mai_n44_), .B(i_6_), .Y(mai_mai_n45_));
  INV        m023(.A(i_2_), .Y(mai_mai_n46_));
  NA2        m024(.A(i_0_), .B(i_3_), .Y(mai_mai_n47_));
  INV        m025(.A(i_5_), .Y(mai_mai_n48_));
  NA2        m026(.A(i_0_), .B(i_2_), .Y(mai_mai_n49_));
  NA2        m027(.A(i_7_), .B(i_9_), .Y(mai_mai_n50_));
  NA3        m028(.A(i_2_), .B(i_6_), .C(i_8_), .Y(mai_mai_n51_));
  NO2        m029(.A(i_1_), .B(i_6_), .Y(mai_mai_n52_));
  NA2        m030(.A(i_8_), .B(i_7_), .Y(mai_mai_n53_));
  OAI210     m031(.A0(mai_mai_n53_), .A1(mai_mai_n52_), .B0(mai_mai_n51_), .Y(mai_mai_n54_));
  NA2        m032(.A(mai_mai_n54_), .B(i_12_), .Y(mai_mai_n55_));
  NAi21      m033(.An(i_2_), .B(i_7_), .Y(mai_mai_n56_));
  INV        m034(.A(i_1_), .Y(mai_mai_n57_));
  NA2        m035(.A(mai_mai_n57_), .B(i_6_), .Y(mai_mai_n58_));
  NA3        m036(.A(mai_mai_n58_), .B(mai_mai_n56_), .C(mai_mai_n31_), .Y(mai_mai_n59_));
  NA2        m037(.A(i_1_), .B(i_10_), .Y(mai_mai_n60_));
  NO2        m038(.A(mai_mai_n60_), .B(i_6_), .Y(mai_mai_n61_));
  NAi31      m039(.An(mai_mai_n61_), .B(mai_mai_n59_), .C(mai_mai_n55_), .Y(mai_mai_n62_));
  AOI210     m040(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(mai_mai_n63_));
  NA2        m041(.A(i_1_), .B(i_6_), .Y(mai_mai_n64_));
  NO2        m042(.A(mai_mai_n64_), .B(mai_mai_n25_), .Y(mai_mai_n65_));
  INV        m043(.A(i_0_), .Y(mai_mai_n66_));
  NAi21      m044(.An(i_5_), .B(i_10_), .Y(mai_mai_n67_));
  NA2        m045(.A(i_5_), .B(i_9_), .Y(mai_mai_n68_));
  AOI210     m046(.A0(mai_mai_n68_), .A1(mai_mai_n67_), .B0(mai_mai_n66_), .Y(mai_mai_n69_));
  NO2        m047(.A(mai_mai_n69_), .B(mai_mai_n65_), .Y(mai_mai_n70_));
  OAI210     m048(.A0(mai_mai_n69_), .A1(mai_mai_n62_), .B0(i_0_), .Y(mai_mai_n71_));
  NA2        m049(.A(i_12_), .B(i_5_), .Y(mai_mai_n72_));
  NA2        m050(.A(i_2_), .B(i_8_), .Y(mai_mai_n73_));
  NO2        m051(.A(mai_mai_n73_), .B(mai_mai_n52_), .Y(mai_mai_n74_));
  NO2        m052(.A(i_3_), .B(i_9_), .Y(mai_mai_n75_));
  NO2        m053(.A(i_3_), .B(i_7_), .Y(mai_mai_n76_));
  INV        m054(.A(i_6_), .Y(mai_mai_n77_));
  OR4        m055(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(mai_mai_n78_));
  INV        m056(.A(mai_mai_n78_), .Y(mai_mai_n79_));
  NO2        m057(.A(i_2_), .B(i_7_), .Y(mai_mai_n80_));
  INV        m058(.A(mai_mai_n74_), .Y(mai_mai_n81_));
  NAi21      m059(.An(i_6_), .B(i_10_), .Y(mai_mai_n82_));
  NA2        m060(.A(i_6_), .B(i_9_), .Y(mai_mai_n83_));
  AOI210     m061(.A0(mai_mai_n83_), .A1(mai_mai_n82_), .B0(mai_mai_n57_), .Y(mai_mai_n84_));
  NA2        m062(.A(i_2_), .B(i_6_), .Y(mai_mai_n85_));
  INV        m063(.A(mai_mai_n84_), .Y(mai_mai_n86_));
  AOI210     m064(.A0(mai_mai_n86_), .A1(mai_mai_n81_), .B0(mai_mai_n72_), .Y(mai_mai_n87_));
  AN3        m065(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n88_));
  NAi21      m066(.An(i_6_), .B(i_11_), .Y(mai_mai_n89_));
  NO2        m067(.A(i_5_), .B(i_8_), .Y(mai_mai_n90_));
  NOi21      m068(.An(mai_mai_n90_), .B(mai_mai_n89_), .Y(mai_mai_n91_));
  AOI220     m069(.A0(mai_mai_n91_), .A1(mai_mai_n56_), .B0(mai_mai_n88_), .B1(mai_mai_n32_), .Y(mai_mai_n92_));
  INV        m070(.A(i_7_), .Y(mai_mai_n93_));
  NA2        m071(.A(mai_mai_n46_), .B(mai_mai_n93_), .Y(mai_mai_n94_));
  NO2        m072(.A(i_0_), .B(i_5_), .Y(mai_mai_n95_));
  NA2        m073(.A(i_12_), .B(i_3_), .Y(mai_mai_n96_));
  INV        m074(.A(mai_mai_n96_), .Y(mai_mai_n97_));
  NA3        m075(.A(mai_mai_n97_), .B(i_6_), .C(mai_mai_n94_), .Y(mai_mai_n98_));
  NAi21      m076(.An(i_7_), .B(i_11_), .Y(mai_mai_n99_));
  NO3        m077(.A(mai_mai_n99_), .B(mai_mai_n82_), .C(mai_mai_n49_), .Y(mai_mai_n100_));
  AN2        m078(.A(i_2_), .B(i_10_), .Y(mai_mai_n101_));
  NO2        m079(.A(mai_mai_n101_), .B(i_7_), .Y(mai_mai_n102_));
  OR2        m080(.A(mai_mai_n72_), .B(mai_mai_n52_), .Y(mai_mai_n103_));
  NO2        m081(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n104_));
  NO3        m082(.A(mai_mai_n104_), .B(mai_mai_n103_), .C(mai_mai_n102_), .Y(mai_mai_n105_));
  NA2        m083(.A(i_12_), .B(i_7_), .Y(mai_mai_n106_));
  NO2        m084(.A(mai_mai_n57_), .B(mai_mai_n26_), .Y(mai_mai_n107_));
  NA2        m085(.A(mai_mai_n107_), .B(i_0_), .Y(mai_mai_n108_));
  NA2        m086(.A(i_11_), .B(i_12_), .Y(mai_mai_n109_));
  OAI210     m087(.A0(mai_mai_n108_), .A1(mai_mai_n106_), .B0(mai_mai_n109_), .Y(mai_mai_n110_));
  NO2        m088(.A(mai_mai_n110_), .B(mai_mai_n105_), .Y(mai_mai_n111_));
  NAi41      m089(.An(mai_mai_n100_), .B(mai_mai_n111_), .C(mai_mai_n98_), .D(mai_mai_n92_), .Y(mai_mai_n112_));
  NOi21      m090(.An(i_1_), .B(i_5_), .Y(mai_mai_n113_));
  NA2        m091(.A(mai_mai_n113_), .B(i_11_), .Y(mai_mai_n114_));
  NA2        m092(.A(mai_mai_n93_), .B(mai_mai_n37_), .Y(mai_mai_n115_));
  NA2        m093(.A(i_7_), .B(mai_mai_n25_), .Y(mai_mai_n116_));
  NA2        m094(.A(mai_mai_n116_), .B(mai_mai_n115_), .Y(mai_mai_n117_));
  NA2        m095(.A(mai_mai_n83_), .B(mai_mai_n82_), .Y(mai_mai_n118_));
  NAi21      m096(.An(i_3_), .B(i_8_), .Y(mai_mai_n119_));
  NA2        m097(.A(mai_mai_n119_), .B(mai_mai_n56_), .Y(mai_mai_n120_));
  NOi21      m098(.An(mai_mai_n120_), .B(mai_mai_n118_), .Y(mai_mai_n121_));
  NO2        m099(.A(i_1_), .B(mai_mai_n77_), .Y(mai_mai_n122_));
  NO2        m100(.A(mai_mai_n121_), .B(mai_mai_n114_), .Y(mai_mai_n123_));
  NO3        m101(.A(mai_mai_n123_), .B(mai_mai_n112_), .C(mai_mai_n87_), .Y(mai_mai_n124_));
  NA2        m102(.A(mai_mai_n124_), .B(mai_mai_n71_), .Y(mai2));
  NO2        m103(.A(mai_mai_n57_), .B(mai_mai_n37_), .Y(mai_mai_n126_));
  NA2        m104(.A(i_6_), .B(mai_mai_n25_), .Y(mai_mai_n127_));
  INV        m105(.A(mai_mai_n126_), .Y(mai_mai_n128_));
  NA3        m106(.A(mai_mai_n128_), .B(mai_mai_n70_), .C(mai_mai_n30_), .Y(mai0));
  AN2        m107(.A(i_8_), .B(i_7_), .Y(mai_mai_n130_));
  NA2        m108(.A(mai_mai_n130_), .B(i_6_), .Y(mai_mai_n131_));
  NO2        m109(.A(i_12_), .B(i_13_), .Y(mai_mai_n132_));
  NAi21      m110(.An(i_5_), .B(i_11_), .Y(mai_mai_n133_));
  NOi21      m111(.An(mai_mai_n132_), .B(mai_mai_n133_), .Y(mai_mai_n134_));
  NO2        m112(.A(i_0_), .B(i_1_), .Y(mai_mai_n135_));
  NA2        m113(.A(i_2_), .B(i_3_), .Y(mai_mai_n136_));
  NO2        m114(.A(mai_mai_n136_), .B(i_4_), .Y(mai_mai_n137_));
  NA2        m115(.A(mai_mai_n137_), .B(mai_mai_n134_), .Y(mai_mai_n138_));
  NA2        m116(.A(i_1_), .B(i_5_), .Y(mai_mai_n139_));
  NO3        m117(.A(i_4_), .B(mai_mai_n139_), .C(mai_mai_n26_), .Y(mai_mai_n140_));
  OR2        m118(.A(i_0_), .B(i_1_), .Y(mai_mai_n141_));
  NO3        m119(.A(mai_mai_n141_), .B(mai_mai_n72_), .C(i_13_), .Y(mai_mai_n142_));
  NAi32      m120(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(mai_mai_n143_));
  NAi21      m121(.An(mai_mai_n143_), .B(mai_mai_n142_), .Y(mai_mai_n144_));
  NOi21      m122(.An(i_4_), .B(i_10_), .Y(mai_mai_n145_));
  NA2        m123(.A(mai_mai_n145_), .B(mai_mai_n39_), .Y(mai_mai_n146_));
  NO2        m124(.A(i_3_), .B(i_5_), .Y(mai_mai_n147_));
  NO3        m125(.A(mai_mai_n66_), .B(i_2_), .C(i_1_), .Y(mai_mai_n148_));
  NO2        m126(.A(mai_mai_n913_), .B(mai_mai_n140_), .Y(mai_mai_n149_));
  AOI210     m127(.A0(mai_mai_n149_), .A1(mai_mai_n138_), .B0(mai_mai_n131_), .Y(mai_mai_n150_));
  NA3        m128(.A(mai_mai_n66_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n151_));
  NOi21      m129(.An(i_4_), .B(i_9_), .Y(mai_mai_n152_));
  NOi21      m130(.An(i_11_), .B(i_13_), .Y(mai_mai_n153_));
  NA2        m131(.A(mai_mai_n153_), .B(mai_mai_n152_), .Y(mai_mai_n154_));
  BUFFER     m132(.A(mai_mai_n154_), .Y(mai_mai_n155_));
  NO2        m133(.A(i_4_), .B(i_5_), .Y(mai_mai_n156_));
  NAi21      m134(.An(i_12_), .B(i_11_), .Y(mai_mai_n157_));
  NO2        m135(.A(mai_mai_n157_), .B(i_13_), .Y(mai_mai_n158_));
  NA2        m136(.A(mai_mai_n158_), .B(mai_mai_n156_), .Y(mai_mai_n159_));
  AOI210     m137(.A0(mai_mai_n159_), .A1(mai_mai_n155_), .B0(mai_mai_n151_), .Y(mai_mai_n160_));
  NO2        m138(.A(mai_mai_n66_), .B(mai_mai_n57_), .Y(mai_mai_n161_));
  NA2        m139(.A(mai_mai_n36_), .B(i_5_), .Y(mai_mai_n162_));
  NAi31      m140(.An(mai_mai_n162_), .B(mai_mai_n75_), .C(i_11_), .Y(mai_mai_n163_));
  NA2        m141(.A(i_3_), .B(i_5_), .Y(mai_mai_n164_));
  OR2        m142(.A(mai_mai_n164_), .B(mai_mai_n154_), .Y(mai_mai_n165_));
  AOI210     m143(.A0(mai_mai_n165_), .A1(mai_mai_n163_), .B0(mai_mai_n57_), .Y(mai_mai_n166_));
  NO2        m144(.A(mai_mai_n66_), .B(i_5_), .Y(mai_mai_n167_));
  NO2        m145(.A(i_13_), .B(i_10_), .Y(mai_mai_n168_));
  NA3        m146(.A(mai_mai_n168_), .B(mai_mai_n167_), .C(mai_mai_n44_), .Y(mai_mai_n169_));
  NO2        m147(.A(i_2_), .B(i_1_), .Y(mai_mai_n170_));
  NAi21      m148(.An(i_4_), .B(i_12_), .Y(mai_mai_n171_));
  NO3        m149(.A(mai_mai_n171_), .B(mai_mai_n909_), .C(mai_mai_n169_), .Y(mai_mai_n172_));
  NO3        m150(.A(mai_mai_n172_), .B(mai_mai_n166_), .C(mai_mai_n160_), .Y(mai_mai_n173_));
  INV        m151(.A(i_8_), .Y(mai_mai_n174_));
  NA2        m152(.A(i_8_), .B(i_6_), .Y(mai_mai_n175_));
  NO3        m153(.A(i_3_), .B(mai_mai_n77_), .C(mai_mai_n48_), .Y(mai_mai_n176_));
  NA2        m154(.A(mai_mai_n176_), .B(mai_mai_n104_), .Y(mai_mai_n177_));
  NO3        m155(.A(i_0_), .B(i_2_), .C(i_1_), .Y(mai_mai_n178_));
  NA3        m156(.A(mai_mai_n178_), .B(mai_mai_n39_), .C(mai_mai_n44_), .Y(mai_mai_n179_));
  NO3        m157(.A(i_11_), .B(i_13_), .C(i_9_), .Y(mai_mai_n180_));
  AOI210     m158(.A0(i_9_), .A1(mai_mai_n179_), .B0(mai_mai_n177_), .Y(mai_mai_n181_));
  NO2        m159(.A(i_3_), .B(i_8_), .Y(mai_mai_n182_));
  NO3        m160(.A(i_11_), .B(i_10_), .C(i_9_), .Y(mai_mai_n183_));
  NA3        m161(.A(mai_mai_n183_), .B(mai_mai_n182_), .C(mai_mai_n39_), .Y(mai_mai_n184_));
  NO2        m162(.A(i_13_), .B(i_9_), .Y(mai_mai_n185_));
  NAi21      m163(.An(i_12_), .B(i_3_), .Y(mai_mai_n186_));
  NO2        m164(.A(mai_mai_n44_), .B(i_5_), .Y(mai_mai_n187_));
  NO3        m165(.A(i_0_), .B(i_2_), .C(mai_mai_n57_), .Y(mai_mai_n188_));
  NA3        m166(.A(mai_mai_n188_), .B(mai_mai_n187_), .C(i_10_), .Y(mai_mai_n189_));
  OAI220     m167(.A0(mai_mai_n189_), .A1(i_13_), .B0(mai_mai_n52_), .B1(mai_mai_n184_), .Y(mai_mai_n190_));
  AOI210     m168(.A0(mai_mai_n190_), .A1(i_7_), .B0(mai_mai_n181_), .Y(mai_mai_n191_));
  OAI220     m169(.A0(mai_mai_n191_), .A1(i_4_), .B0(mai_mai_n175_), .B1(mai_mai_n173_), .Y(mai_mai_n192_));
  NAi21      m170(.An(i_12_), .B(i_7_), .Y(mai_mai_n193_));
  NA3        m171(.A(i_13_), .B(mai_mai_n174_), .C(i_10_), .Y(mai_mai_n194_));
  NA2        m172(.A(i_0_), .B(i_5_), .Y(mai_mai_n195_));
  NAi31      m173(.An(i_9_), .B(i_6_), .C(i_5_), .Y(mai_mai_n196_));
  NO2        m174(.A(mai_mai_n36_), .B(i_13_), .Y(mai_mai_n197_));
  NO2        m175(.A(mai_mai_n66_), .B(mai_mai_n26_), .Y(mai_mai_n198_));
  NO2        m176(.A(mai_mai_n46_), .B(mai_mai_n57_), .Y(mai_mai_n199_));
  NA3        m177(.A(mai_mai_n199_), .B(mai_mai_n198_), .C(mai_mai_n197_), .Y(mai_mai_n200_));
  INV        m178(.A(i_13_), .Y(mai_mai_n201_));
  NO2        m179(.A(i_12_), .B(mai_mai_n201_), .Y(mai_mai_n202_));
  NA2        m180(.A(mai_mai_n914_), .B(mai_mai_n130_), .Y(mai_mai_n203_));
  NO2        m181(.A(i_12_), .B(mai_mai_n37_), .Y(mai_mai_n204_));
  NO2        m182(.A(mai_mai_n164_), .B(i_4_), .Y(mai_mai_n205_));
  NA2        m183(.A(mai_mai_n205_), .B(mai_mai_n204_), .Y(mai_mai_n206_));
  OR2        m184(.A(i_8_), .B(i_7_), .Y(mai_mai_n207_));
  NO2        m185(.A(mai_mai_n49_), .B(i_1_), .Y(mai_mai_n208_));
  INV        m186(.A(i_12_), .Y(mai_mai_n209_));
  NO3        m187(.A(mai_mai_n36_), .B(i_8_), .C(i_10_), .Y(mai_mai_n210_));
  NA2        m188(.A(i_2_), .B(i_1_), .Y(mai_mai_n211_));
  NO2        m189(.A(mai_mai_n49_), .B(mai_mai_n206_), .Y(mai_mai_n212_));
  NO3        m190(.A(i_11_), .B(i_7_), .C(mai_mai_n37_), .Y(mai_mai_n213_));
  NAi21      m191(.An(i_4_), .B(i_3_), .Y(mai_mai_n214_));
  NO2        m192(.A(i_0_), .B(i_6_), .Y(mai_mai_n215_));
  NOi41      m193(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(mai_mai_n216_));
  NA2        m194(.A(mai_mai_n216_), .B(mai_mai_n215_), .Y(mai_mai_n217_));
  AOI210     m195(.A0(mai_mai_n905_), .A1(mai_mai_n39_), .B0(mai_mai_n212_), .Y(mai_mai_n218_));
  NO2        m196(.A(i_11_), .B(mai_mai_n201_), .Y(mai_mai_n219_));
  NOi21      m197(.An(i_1_), .B(i_6_), .Y(mai_mai_n220_));
  NAi21      m198(.An(i_3_), .B(i_7_), .Y(mai_mai_n221_));
  NO2        m199(.A(i_12_), .B(i_3_), .Y(mai_mai_n222_));
  NA2        m200(.A(mai_mai_n66_), .B(i_5_), .Y(mai_mai_n223_));
  NA2        m201(.A(i_3_), .B(i_9_), .Y(mai_mai_n224_));
  NA3        m202(.A(i_1_), .B(i_8_), .C(i_7_), .Y(mai_mai_n225_));
  NO2        m203(.A(mai_mai_n917_), .B(mai_mai_n68_), .Y(mai_mai_n226_));
  NA2        m204(.A(mai_mai_n226_), .B(mai_mai_n130_), .Y(mai_mai_n227_));
  NO2        m205(.A(mai_mai_n207_), .B(mai_mai_n37_), .Y(mai_mai_n228_));
  NA2        m206(.A(i_12_), .B(i_6_), .Y(mai_mai_n229_));
  OR2        m207(.A(i_13_), .B(i_9_), .Y(mai_mai_n230_));
  NO3        m208(.A(mai_mai_n230_), .B(mai_mai_n229_), .C(mai_mai_n48_), .Y(mai_mai_n231_));
  NO2        m209(.A(mai_mai_n214_), .B(i_2_), .Y(mai_mai_n232_));
  NA3        m210(.A(mai_mai_n232_), .B(mai_mai_n231_), .C(mai_mai_n44_), .Y(mai_mai_n233_));
  NA2        m211(.A(mai_mai_n219_), .B(i_9_), .Y(mai_mai_n234_));
  NA2        m212(.A(mai_mai_n223_), .B(mai_mai_n58_), .Y(mai_mai_n235_));
  OAI210     m213(.A0(mai_mai_n235_), .A1(mai_mai_n234_), .B0(mai_mai_n233_), .Y(mai_mai_n236_));
  NO2        m214(.A(i_11_), .B(mai_mai_n201_), .Y(mai_mai_n237_));
  NO2        m215(.A(mai_mai_n221_), .B(i_8_), .Y(mai_mai_n238_));
  NO2        m216(.A(i_6_), .B(mai_mai_n48_), .Y(mai_mai_n239_));
  NA3        m217(.A(i_3_), .B(mai_mai_n228_), .C(mai_mai_n202_), .Y(mai_mai_n240_));
  NO2        m218(.A(mai_mai_n240_), .B(mai_mai_n908_), .Y(mai_mai_n241_));
  AOI210     m219(.A0(mai_mai_n236_), .A1(mai_mai_n228_), .B0(mai_mai_n241_), .Y(mai_mai_n242_));
  NA4        m220(.A(mai_mai_n242_), .B(mai_mai_n227_), .C(mai_mai_n218_), .D(mai_mai_n203_), .Y(mai_mai_n243_));
  NO3        m221(.A(i_12_), .B(mai_mai_n201_), .C(mai_mai_n37_), .Y(mai_mai_n244_));
  INV        m222(.A(mai_mai_n244_), .Y(mai_mai_n245_));
  NA2        m223(.A(i_8_), .B(mai_mai_n93_), .Y(mai_mai_n246_));
  NO3        m224(.A(i_0_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n247_));
  NO2        m225(.A(mai_mai_n211_), .B(i_0_), .Y(mai_mai_n248_));
  NA2        m226(.A(mai_mai_n239_), .B(mai_mai_n26_), .Y(mai_mai_n249_));
  NO2        m227(.A(mai_mai_n249_), .B(mai_mai_n906_), .Y(mai_mai_n250_));
  NA2        m228(.A(i_0_), .B(i_1_), .Y(mai_mai_n251_));
  NO2        m229(.A(mai_mai_n251_), .B(i_2_), .Y(mai_mai_n252_));
  NO2        m230(.A(mai_mai_n53_), .B(i_6_), .Y(mai_mai_n253_));
  NA3        m231(.A(mai_mai_n253_), .B(mai_mai_n252_), .C(mai_mai_n147_), .Y(mai_mai_n254_));
  NA2        m232(.A(mai_mai_n131_), .B(mai_mai_n254_), .Y(mai_mai_n255_));
  NO2        m233(.A(mai_mai_n255_), .B(mai_mai_n250_), .Y(mai_mai_n256_));
  NO2        m234(.A(i_3_), .B(i_10_), .Y(mai_mai_n257_));
  NA3        m235(.A(mai_mai_n257_), .B(mai_mai_n39_), .C(mai_mai_n44_), .Y(mai_mai_n258_));
  NO2        m236(.A(i_2_), .B(mai_mai_n93_), .Y(mai_mai_n259_));
  NA2        m237(.A(i_1_), .B(mai_mai_n36_), .Y(mai_mai_n260_));
  NO2        m238(.A(mai_mai_n260_), .B(i_8_), .Y(mai_mai_n261_));
  INV        m239(.A(mai_mai_n261_), .Y(mai_mai_n262_));
  AN2        m240(.A(i_3_), .B(i_10_), .Y(mai_mai_n263_));
  NA3        m241(.A(mai_mai_n263_), .B(mai_mai_n158_), .C(mai_mai_n156_), .Y(mai_mai_n264_));
  NO2        m242(.A(mai_mai_n46_), .B(mai_mai_n26_), .Y(mai_mai_n265_));
  OR2        m243(.A(mai_mai_n262_), .B(mai_mai_n258_), .Y(mai_mai_n266_));
  OAI220     m244(.A0(mai_mai_n266_), .A1(i_6_), .B0(mai_mai_n256_), .B1(mai_mai_n245_), .Y(mai_mai_n267_));
  NO4        m245(.A(mai_mai_n267_), .B(mai_mai_n243_), .C(mai_mai_n192_), .D(mai_mai_n150_), .Y(mai_mai_n268_));
  NO3        m246(.A(mai_mai_n44_), .B(i_13_), .C(i_9_), .Y(mai_mai_n269_));
  NO2        m247(.A(mai_mai_n53_), .B(mai_mai_n77_), .Y(mai_mai_n270_));
  NA2        m248(.A(mai_mai_n248_), .B(mai_mai_n270_), .Y(mai_mai_n271_));
  NO3        m249(.A(i_6_), .B(mai_mai_n174_), .C(i_7_), .Y(mai_mai_n272_));
  NA2        m250(.A(mai_mai_n912_), .B(mai_mai_n271_), .Y(mai_mai_n273_));
  NO2        m251(.A(i_2_), .B(i_3_), .Y(mai_mai_n274_));
  OR2        m252(.A(i_0_), .B(i_5_), .Y(mai_mai_n275_));
  NA2        m253(.A(mai_mai_n195_), .B(mai_mai_n275_), .Y(mai_mai_n276_));
  NA4        m254(.A(mai_mai_n276_), .B(i_6_), .C(mai_mai_n274_), .D(i_1_), .Y(mai_mai_n277_));
  NA2        m255(.A(mai_mai_n248_), .B(mai_mai_n147_), .Y(mai_mai_n278_));
  NAi21      m256(.An(i_8_), .B(i_7_), .Y(mai_mai_n279_));
  NO2        m257(.A(mai_mai_n279_), .B(i_6_), .Y(mai_mai_n280_));
  NO2        m258(.A(mai_mai_n141_), .B(mai_mai_n46_), .Y(mai_mai_n281_));
  NA2        m259(.A(mai_mai_n281_), .B(mai_mai_n280_), .Y(mai_mai_n282_));
  NA3        m260(.A(mai_mai_n282_), .B(mai_mai_n278_), .C(mai_mai_n277_), .Y(mai_mai_n283_));
  OAI210     m261(.A0(mai_mai_n283_), .A1(mai_mai_n273_), .B0(i_4_), .Y(mai_mai_n284_));
  NO2        m262(.A(i_12_), .B(i_10_), .Y(mai_mai_n285_));
  NOi21      m263(.An(i_5_), .B(i_0_), .Y(mai_mai_n286_));
  NO2        m264(.A(mai_mai_n260_), .B(mai_mai_n119_), .Y(mai_mai_n287_));
  NA4        m265(.A(mai_mai_n76_), .B(mai_mai_n36_), .C(mai_mai_n77_), .D(i_8_), .Y(mai_mai_n288_));
  NA2        m266(.A(mai_mai_n287_), .B(mai_mai_n285_), .Y(mai_mai_n289_));
  NO2        m267(.A(i_6_), .B(i_8_), .Y(mai_mai_n290_));
  NOi21      m268(.An(i_0_), .B(i_2_), .Y(mai_mai_n291_));
  AN2        m269(.A(mai_mai_n291_), .B(mai_mai_n290_), .Y(mai_mai_n292_));
  NO2        m270(.A(i_1_), .B(i_7_), .Y(mai_mai_n293_));
  AO220      m271(.A0(mai_mai_n293_), .A1(mai_mai_n292_), .B0(mai_mai_n280_), .B1(mai_mai_n208_), .Y(mai_mai_n294_));
  NA2        m272(.A(mai_mai_n294_), .B(mai_mai_n41_), .Y(mai_mai_n295_));
  NA3        m273(.A(mai_mai_n295_), .B(mai_mai_n289_), .C(mai_mai_n284_), .Y(mai_mai_n296_));
  NO3        m274(.A(mai_mai_n207_), .B(mai_mai_n46_), .C(i_1_), .Y(mai_mai_n297_));
  NO3        m275(.A(mai_mai_n279_), .B(i_2_), .C(i_1_), .Y(mai_mai_n298_));
  OAI210     m276(.A0(mai_mai_n298_), .A1(mai_mai_n297_), .B0(i_6_), .Y(mai_mai_n299_));
  NA2        m277(.A(mai_mai_n259_), .B(mai_mai_n174_), .Y(mai_mai_n300_));
  NA2        m278(.A(mai_mai_n300_), .B(mai_mai_n299_), .Y(mai_mai_n301_));
  NA2        m279(.A(mai_mai_n301_), .B(i_3_), .Y(mai_mai_n302_));
  INV        m280(.A(mai_mai_n76_), .Y(mai_mai_n303_));
  NO2        m281(.A(mai_mai_n85_), .B(mai_mai_n174_), .Y(mai_mai_n304_));
  NO2        m282(.A(mai_mai_n73_), .B(mai_mai_n303_), .Y(mai_mai_n305_));
  NO2        m283(.A(mai_mai_n174_), .B(i_9_), .Y(mai_mai_n306_));
  INV        m284(.A(mai_mai_n306_), .Y(mai_mai_n307_));
  NO2        m285(.A(mai_mai_n305_), .B(mai_mai_n250_), .Y(mai_mai_n308_));
  AOI210     m286(.A0(mai_mai_n308_), .A1(mai_mai_n302_), .B0(mai_mai_n146_), .Y(mai_mai_n309_));
  AOI210     m287(.A0(mai_mai_n296_), .A1(mai_mai_n269_), .B0(mai_mai_n309_), .Y(mai_mai_n310_));
  NOi32      m288(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(mai_mai_n311_));
  INV        m289(.A(mai_mai_n311_), .Y(mai_mai_n312_));
  NAi21      m290(.An(i_0_), .B(i_6_), .Y(mai_mai_n313_));
  NAi21      m291(.An(i_1_), .B(i_5_), .Y(mai_mai_n314_));
  NA2        m292(.A(mai_mai_n314_), .B(mai_mai_n313_), .Y(mai_mai_n315_));
  NA2        m293(.A(mai_mai_n315_), .B(mai_mai_n25_), .Y(mai_mai_n316_));
  OAI210     m294(.A0(mai_mai_n316_), .A1(mai_mai_n143_), .B0(mai_mai_n217_), .Y(mai_mai_n317_));
  NAi41      m295(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(mai_mai_n318_));
  OAI220     m296(.A0(mai_mai_n318_), .A1(mai_mai_n314_), .B0(mai_mai_n196_), .B1(mai_mai_n143_), .Y(mai_mai_n319_));
  AOI210     m297(.A0(mai_mai_n318_), .A1(mai_mai_n143_), .B0(mai_mai_n141_), .Y(mai_mai_n320_));
  NOi32      m298(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(mai_mai_n321_));
  NAi21      m299(.An(i_6_), .B(i_1_), .Y(mai_mai_n322_));
  NA3        m300(.A(mai_mai_n322_), .B(mai_mai_n321_), .C(mai_mai_n46_), .Y(mai_mai_n323_));
  NO2        m301(.A(mai_mai_n323_), .B(i_0_), .Y(mai_mai_n324_));
  OR3        m302(.A(mai_mai_n324_), .B(mai_mai_n320_), .C(mai_mai_n319_), .Y(mai_mai_n325_));
  NO2        m303(.A(i_1_), .B(mai_mai_n93_), .Y(mai_mai_n326_));
  NAi21      m304(.An(i_3_), .B(i_4_), .Y(mai_mai_n327_));
  NO2        m305(.A(mai_mai_n327_), .B(i_9_), .Y(mai_mai_n328_));
  AN2        m306(.A(i_6_), .B(i_7_), .Y(mai_mai_n329_));
  NA2        m307(.A(i_2_), .B(i_7_), .Y(mai_mai_n330_));
  NO2        m308(.A(mai_mai_n327_), .B(i_10_), .Y(mai_mai_n331_));
  NA3        m309(.A(mai_mai_n331_), .B(mai_mai_n330_), .C(mai_mai_n215_), .Y(mai_mai_n332_));
  INV        m310(.A(mai_mai_n332_), .Y(mai_mai_n333_));
  AOI210     m311(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(mai_mai_n334_));
  OAI210     m312(.A0(mai_mai_n334_), .A1(mai_mai_n170_), .B0(mai_mai_n331_), .Y(mai_mai_n335_));
  AOI220     m313(.A0(mai_mai_n331_), .A1(mai_mai_n293_), .B0(mai_mai_n210_), .B1(mai_mai_n170_), .Y(mai_mai_n336_));
  AOI210     m314(.A0(mai_mai_n336_), .A1(mai_mai_n335_), .B0(i_5_), .Y(mai_mai_n337_));
  NO4        m315(.A(mai_mai_n337_), .B(mai_mai_n333_), .C(mai_mai_n325_), .D(mai_mai_n317_), .Y(mai_mai_n338_));
  NO2        m316(.A(mai_mai_n338_), .B(mai_mai_n312_), .Y(mai_mai_n339_));
  INV        m317(.A(mai_mai_n53_), .Y(mai_mai_n340_));
  AN2        m318(.A(i_12_), .B(i_5_), .Y(mai_mai_n341_));
  NO2        m319(.A(i_4_), .B(mai_mai_n26_), .Y(mai_mai_n342_));
  NA2        m320(.A(mai_mai_n342_), .B(mai_mai_n341_), .Y(mai_mai_n343_));
  NO2        m321(.A(i_11_), .B(i_6_), .Y(mai_mai_n344_));
  INV        m322(.A(mai_mai_n343_), .Y(mai_mai_n345_));
  NO2        m323(.A(mai_mai_n214_), .B(i_5_), .Y(mai_mai_n346_));
  NO2        m324(.A(i_5_), .B(i_10_), .Y(mai_mai_n347_));
  NA2        m325(.A(mai_mai_n132_), .B(mai_mai_n45_), .Y(mai_mai_n348_));
  NO2        m326(.A(mai_mai_n348_), .B(mai_mai_n214_), .Y(mai_mai_n349_));
  OAI210     m327(.A0(mai_mai_n349_), .A1(mai_mai_n345_), .B0(mai_mai_n340_), .Y(mai_mai_n350_));
  NO2        m328(.A(mai_mai_n37_), .B(mai_mai_n25_), .Y(mai_mai_n351_));
  NO3        m329(.A(mai_mai_n77_), .B(mai_mai_n48_), .C(i_9_), .Y(mai_mai_n352_));
  NA2        m330(.A(mai_mai_n347_), .B(mai_mai_n209_), .Y(mai_mai_n353_));
  NA2        m331(.A(mai_mai_n41_), .B(i_11_), .Y(mai_mai_n354_));
  OAI220     m332(.A0(mai_mai_n354_), .A1(mai_mai_n196_), .B0(mai_mai_n353_), .B1(mai_mai_n288_), .Y(mai_mai_n355_));
  NAi21      m333(.An(i_13_), .B(i_0_), .Y(mai_mai_n356_));
  NA2        m334(.A(mai_mai_n355_), .B(i_0_), .Y(mai_mai_n357_));
  NA2        m335(.A(mai_mai_n357_), .B(mai_mai_n350_), .Y(mai_mai_n358_));
  NO2        m336(.A(i_0_), .B(i_11_), .Y(mai_mai_n359_));
  NOi21      m337(.An(i_2_), .B(i_12_), .Y(mai_mai_n360_));
  NA2        m338(.A(mai_mai_n130_), .B(i_9_), .Y(mai_mai_n361_));
  NO2        m339(.A(mai_mai_n361_), .B(i_4_), .Y(mai_mai_n362_));
  OR2        m340(.A(i_13_), .B(i_10_), .Y(mai_mai_n363_));
  NO2        m341(.A(mai_mai_n154_), .B(mai_mai_n115_), .Y(mai_mai_n364_));
  OR2        m342(.A(mai_mai_n194_), .B(mai_mai_n193_), .Y(mai_mai_n365_));
  NO2        m343(.A(mai_mai_n93_), .B(mai_mai_n25_), .Y(mai_mai_n366_));
  NO2        m344(.A(mai_mai_n365_), .B(mai_mai_n26_), .Y(mai_mai_n367_));
  INV        m345(.A(mai_mai_n277_), .Y(mai_mai_n368_));
  AOI220     m346(.A0(mai_mai_n253_), .A1(mai_mai_n247_), .B0(mai_mai_n248_), .B1(mai_mai_n270_), .Y(mai_mai_n369_));
  INV        m347(.A(mai_mai_n369_), .Y(mai_mai_n370_));
  NO2        m348(.A(i_2_), .B(mai_mai_n246_), .Y(mai_mai_n371_));
  NO3        m349(.A(mai_mai_n371_), .B(mai_mai_n370_), .C(mai_mai_n368_), .Y(mai_mai_n372_));
  NO2        m350(.A(i_3_), .B(mai_mai_n279_), .Y(mai_mai_n373_));
  NA2        m351(.A(mai_mai_n253_), .B(mai_mai_n208_), .Y(mai_mai_n374_));
  NO2        m352(.A(mai_mai_n292_), .B(mai_mai_n373_), .Y(mai_mai_n375_));
  AOI210     m353(.A0(mai_mai_n375_), .A1(mai_mai_n372_), .B0(mai_mai_n234_), .Y(mai_mai_n376_));
  NO4        m354(.A(mai_mai_n376_), .B(mai_mai_n367_), .C(mai_mai_n358_), .D(mai_mai_n339_), .Y(mai_mai_n377_));
  NO2        m355(.A(mai_mai_n57_), .B(i_4_), .Y(mai_mai_n378_));
  NA2        m356(.A(mai_mai_n378_), .B(i_2_), .Y(mai_mai_n379_));
  NO2        m357(.A(i_10_), .B(i_9_), .Y(mai_mai_n380_));
  NAi21      m358(.An(i_12_), .B(i_8_), .Y(mai_mai_n381_));
  NO2        m359(.A(mai_mai_n381_), .B(i_3_), .Y(mai_mai_n382_));
  NA2        m360(.A(mai_mai_n382_), .B(mai_mai_n380_), .Y(mai_mai_n383_));
  NO2        m361(.A(mai_mai_n46_), .B(i_4_), .Y(mai_mai_n384_));
  NA2        m362(.A(mai_mai_n384_), .B(i_6_), .Y(mai_mai_n385_));
  OAI220     m363(.A0(mai_mai_n385_), .A1(mai_mai_n184_), .B0(mai_mai_n383_), .B1(mai_mai_n379_), .Y(mai_mai_n386_));
  NA2        m364(.A(mai_mai_n265_), .B(i_0_), .Y(mai_mai_n387_));
  NO3        m365(.A(mai_mai_n23_), .B(i_10_), .C(i_9_), .Y(mai_mai_n388_));
  NA2        m366(.A(mai_mai_n229_), .B(mai_mai_n89_), .Y(mai_mai_n389_));
  NA2        m367(.A(mai_mai_n389_), .B(mai_mai_n388_), .Y(mai_mai_n390_));
  NA2        m368(.A(i_8_), .B(i_9_), .Y(mai_mai_n391_));
  NO2        m369(.A(mai_mai_n390_), .B(mai_mai_n387_), .Y(mai_mai_n392_));
  NO3        m370(.A(i_6_), .B(i_8_), .C(i_7_), .Y(mai_mai_n393_));
  NA3        m371(.A(i_2_), .B(i_10_), .C(i_9_), .Y(mai_mai_n394_));
  NO2        m372(.A(mai_mai_n392_), .B(mai_mai_n386_), .Y(mai_mai_n395_));
  OR2        m373(.A(mai_mai_n251_), .B(i_13_), .Y(mai_mai_n396_));
  OA210      m374(.A0(mai_mai_n307_), .A1(mai_mai_n93_), .B0(mai_mai_n254_), .Y(mai_mai_n397_));
  OA220      m375(.A0(mai_mai_n397_), .A1(mai_mai_n146_), .B0(mai_mai_n396_), .B1(mai_mai_n206_), .Y(mai_mai_n398_));
  NA2        m376(.A(mai_mai_n88_), .B(i_13_), .Y(mai_mai_n399_));
  NO2        m377(.A(i_2_), .B(i_13_), .Y(mai_mai_n400_));
  NA3        m378(.A(mai_mai_n400_), .B(mai_mai_n145_), .C(mai_mai_n91_), .Y(mai_mai_n401_));
  NO3        m379(.A(i_4_), .B(mai_mai_n48_), .C(i_8_), .Y(mai_mai_n402_));
  NO2        m380(.A(i_6_), .B(i_7_), .Y(mai_mai_n403_));
  NO2        m381(.A(i_11_), .B(i_1_), .Y(mai_mai_n404_));
  OR2        m382(.A(i_11_), .B(i_8_), .Y(mai_mai_n405_));
  NOi21      m383(.An(i_2_), .B(i_7_), .Y(mai_mai_n406_));
  NAi21      m384(.An(mai_mai_n405_), .B(mai_mai_n406_), .Y(mai_mai_n407_));
  NO2        m385(.A(mai_mai_n363_), .B(i_6_), .Y(mai_mai_n408_));
  NA3        m386(.A(mai_mai_n408_), .B(mai_mai_n378_), .C(mai_mai_n68_), .Y(mai_mai_n409_));
  NO2        m387(.A(mai_mai_n409_), .B(mai_mai_n407_), .Y(mai_mai_n410_));
  NO2        m388(.A(i_3_), .B(mai_mai_n174_), .Y(mai_mai_n411_));
  NO2        m389(.A(i_6_), .B(i_10_), .Y(mai_mai_n412_));
  NA3        m390(.A(mai_mai_n412_), .B(mai_mai_n269_), .C(mai_mai_n411_), .Y(mai_mai_n413_));
  NO2        m391(.A(mai_mai_n413_), .B(i_4_), .Y(mai_mai_n414_));
  NO2        m392(.A(mai_mai_n141_), .B(i_3_), .Y(mai_mai_n415_));
  NA3        m393(.A(mai_mai_n351_), .B(mai_mai_n161_), .C(mai_mai_n137_), .Y(mai_mai_n416_));
  INV        m394(.A(mai_mai_n416_), .Y(mai_mai_n417_));
  NO3        m395(.A(mai_mai_n417_), .B(mai_mai_n414_), .C(mai_mai_n410_), .Y(mai_mai_n418_));
  NA2        m396(.A(mai_mai_n393_), .B(mai_mai_n347_), .Y(mai_mai_n419_));
  NO2        m397(.A(mai_mai_n419_), .B(mai_mai_n200_), .Y(mai_mai_n420_));
  NO2        m398(.A(i_0_), .B(mai_mai_n77_), .Y(mai_mai_n421_));
  NA3        m399(.A(mai_mai_n421_), .B(mai_mai_n907_), .C(mai_mai_n130_), .Y(mai_mai_n422_));
  OR3        m400(.A(mai_mai_n260_), .B(i_11_), .C(mai_mai_n46_), .Y(mai_mai_n423_));
  NO2        m401(.A(mai_mai_n423_), .B(mai_mai_n422_), .Y(mai_mai_n424_));
  NA3        m402(.A(mai_mai_n263_), .B(mai_mai_n199_), .C(mai_mai_n66_), .Y(mai_mai_n425_));
  NO2        m403(.A(mai_mai_n425_), .B(i_4_), .Y(mai_mai_n426_));
  NO3        m404(.A(mai_mai_n426_), .B(mai_mai_n424_), .C(mai_mai_n420_), .Y(mai_mai_n427_));
  NA4        m405(.A(mai_mai_n427_), .B(mai_mai_n418_), .C(mai_mai_n398_), .D(mai_mai_n395_), .Y(mai_mai_n428_));
  NA3        m406(.A(mai_mai_n263_), .B(mai_mai_n158_), .C(mai_mai_n156_), .Y(mai_mai_n429_));
  INV        m407(.A(mai_mai_n429_), .Y(mai_mai_n430_));
  BUFFER     m408(.A(mai_mai_n247_), .Y(mai_mai_n431_));
  NA2        m409(.A(mai_mai_n431_), .B(mai_mai_n430_), .Y(mai_mai_n432_));
  NA2        m410(.A(mai_mai_n114_), .B(mai_mai_n103_), .Y(mai_mai_n433_));
  AN2        m411(.A(mai_mai_n433_), .B(mai_mai_n388_), .Y(mai_mai_n434_));
  OAI210     m412(.A0(mai_mai_n44_), .A1(mai_mai_n206_), .B0(mai_mai_n264_), .Y(mai_mai_n435_));
  AOI220     m413(.A0(mai_mai_n435_), .A1(mai_mai_n280_), .B0(mai_mai_n434_), .B1(mai_mai_n265_), .Y(mai_mai_n436_));
  NA3        m414(.A(mai_mai_n378_), .B(mai_mai_n182_), .C(i_2_), .Y(mai_mai_n437_));
  INV        m415(.A(mai_mai_n437_), .Y(mai_mai_n438_));
  NA2        m416(.A(mai_mai_n311_), .B(mai_mai_n66_), .Y(mai_mai_n439_));
  NA2        m417(.A(mai_mai_n329_), .B(mai_mai_n321_), .Y(mai_mai_n440_));
  NO2        m418(.A(mai_mai_n36_), .B(i_8_), .Y(mai_mai_n441_));
  NA2        m419(.A(mai_mai_n38_), .B(i_13_), .Y(mai_mai_n442_));
  INV        m420(.A(mai_mai_n442_), .Y(mai_mai_n443_));
  AOI210     m421(.A0(mai_mai_n438_), .A1(mai_mai_n183_), .B0(mai_mai_n443_), .Y(mai_mai_n444_));
  NO2        m422(.A(i_7_), .B(mai_mai_n179_), .Y(mai_mai_n445_));
  OR2        m423(.A(mai_mai_n164_), .B(i_4_), .Y(mai_mai_n446_));
  NO2        m424(.A(mai_mai_n446_), .B(mai_mai_n77_), .Y(mai_mai_n447_));
  AOI220     m425(.A0(mai_mai_n447_), .A1(mai_mai_n445_), .B0(mai_mai_n223_), .B1(mai_mai_n364_), .Y(mai_mai_n448_));
  NA4        m426(.A(mai_mai_n448_), .B(mai_mai_n444_), .C(mai_mai_n436_), .D(mai_mai_n432_), .Y(mai_mai_n449_));
  NA2        m427(.A(mai_mai_n346_), .B(mai_mai_n252_), .Y(mai_mai_n450_));
  OAI210     m428(.A0(mai_mai_n343_), .A1(mai_mai_n151_), .B0(mai_mai_n450_), .Y(mai_mai_n451_));
  NO2        m429(.A(i_12_), .B(mai_mai_n174_), .Y(mai_mai_n452_));
  NA2        m430(.A(mai_mai_n452_), .B(mai_mai_n201_), .Y(mai_mai_n453_));
  NO2        m431(.A(i_6_), .B(mai_mai_n453_), .Y(mai_mai_n454_));
  NOi21      m432(.An(mai_mai_n272_), .B(i_11_), .Y(mai_mai_n455_));
  OAI210     m433(.A0(mai_mai_n455_), .A1(mai_mai_n454_), .B0(mai_mai_n451_), .Y(mai_mai_n456_));
  NO2        m434(.A(i_8_), .B(i_7_), .Y(mai_mai_n457_));
  NO2        m435(.A(mai_mai_n46_), .B(mai_mai_n446_), .Y(mai_mai_n458_));
  NO2        m436(.A(mai_mai_n915_), .B(i_6_), .Y(mai_mai_n459_));
  NA2        m437(.A(mai_mai_n459_), .B(mai_mai_n458_), .Y(mai_mai_n460_));
  INV        m438(.A(mai_mai_n399_), .Y(mai_mai_n461_));
  NA2        m439(.A(mai_mai_n461_), .B(mai_mai_n228_), .Y(mai_mai_n462_));
  NA3        m440(.A(mai_mai_n263_), .B(mai_mai_n156_), .C(mai_mai_n88_), .Y(mai_mai_n463_));
  NO2        m441(.A(mai_mai_n197_), .B(mai_mai_n44_), .Y(mai_mai_n464_));
  NO2        m442(.A(mai_mai_n141_), .B(i_5_), .Y(mai_mai_n465_));
  NA2        m443(.A(mai_mai_n465_), .B(mai_mai_n274_), .Y(mai_mai_n466_));
  OAI210     m444(.A0(mai_mai_n466_), .A1(mai_mai_n464_), .B0(mai_mai_n463_), .Y(mai_mai_n467_));
  NA2        m445(.A(mai_mai_n467_), .B(mai_mai_n393_), .Y(mai_mai_n468_));
  NA4        m446(.A(mai_mai_n468_), .B(mai_mai_n462_), .C(mai_mai_n460_), .D(mai_mai_n456_), .Y(mai_mai_n469_));
  NA2        m447(.A(mai_mai_n244_), .B(mai_mai_n76_), .Y(mai_mai_n470_));
  NO2        m448(.A(mai_mai_n73_), .B(mai_mai_n470_), .Y(mai_mai_n471_));
  NA2        m449(.A(mai_mai_n253_), .B(mai_mai_n247_), .Y(mai_mai_n472_));
  NO2        m450(.A(mai_mai_n472_), .B(mai_mai_n155_), .Y(mai_mai_n473_));
  NA2        m451(.A(mai_mai_n199_), .B(mai_mai_n198_), .Y(mai_mai_n474_));
  NA2        m452(.A(mai_mai_n380_), .B(mai_mai_n197_), .Y(mai_mai_n475_));
  NO2        m453(.A(mai_mai_n474_), .B(mai_mai_n475_), .Y(mai_mai_n476_));
  AOI210     m454(.A0(mai_mai_n322_), .A1(mai_mai_n46_), .B0(mai_mai_n326_), .Y(mai_mai_n477_));
  NA2        m455(.A(mai_mai_n452_), .B(mai_mai_n237_), .Y(mai_mai_n478_));
  NO2        m456(.A(mai_mai_n477_), .B(mai_mai_n478_), .Y(mai_mai_n479_));
  NO4        m457(.A(mai_mai_n479_), .B(mai_mai_n476_), .C(mai_mai_n473_), .D(mai_mai_n471_), .Y(mai_mai_n480_));
  NO4        m458(.A(mai_mai_n220_), .B(mai_mai_n42_), .C(i_2_), .D(mai_mai_n48_), .Y(mai_mai_n481_));
  NO3        m459(.A(i_1_), .B(i_5_), .C(i_10_), .Y(mai_mai_n482_));
  NO2        m460(.A(mai_mai_n207_), .B(mai_mai_n36_), .Y(mai_mai_n483_));
  AN2        m461(.A(mai_mai_n483_), .B(mai_mai_n482_), .Y(mai_mai_n484_));
  OA210      m462(.A0(mai_mai_n484_), .A1(mai_mai_n481_), .B0(mai_mai_n311_), .Y(mai_mai_n485_));
  NO2        m463(.A(mai_mai_n363_), .B(i_1_), .Y(mai_mai_n486_));
  NOi31      m464(.An(mai_mai_n486_), .B(mai_mai_n389_), .C(mai_mai_n66_), .Y(mai_mai_n487_));
  AN2        m465(.A(mai_mai_n487_), .B(mai_mai_n362_), .Y(mai_mai_n488_));
  NO2        m466(.A(mai_mai_n369_), .B(mai_mai_n159_), .Y(mai_mai_n489_));
  NO3        m467(.A(mai_mai_n489_), .B(mai_mai_n488_), .C(mai_mai_n485_), .Y(mai_mai_n490_));
  NOi21      m468(.An(i_10_), .B(i_6_), .Y(mai_mai_n491_));
  NO2        m469(.A(mai_mai_n77_), .B(mai_mai_n25_), .Y(mai_mai_n492_));
  NA2        m470(.A(mai_mai_n237_), .B(mai_mai_n491_), .Y(mai_mai_n493_));
  NO2        m471(.A(mai_mai_n493_), .B(mai_mai_n387_), .Y(mai_mai_n494_));
  NO2        m472(.A(mai_mai_n106_), .B(mai_mai_n23_), .Y(mai_mai_n495_));
  NA2        m473(.A(mai_mai_n272_), .B(mai_mai_n148_), .Y(mai_mai_n496_));
  AOI220     m474(.A0(mai_mai_n496_), .A1(mai_mai_n374_), .B0(mai_mai_n165_), .B1(mai_mai_n163_), .Y(mai_mai_n497_));
  NOi21      m475(.An(mai_mai_n134_), .B(mai_mai_n288_), .Y(mai_mai_n498_));
  NO3        m476(.A(mai_mai_n498_), .B(mai_mai_n497_), .C(mai_mai_n494_), .Y(mai_mai_n499_));
  NO2        m477(.A(mai_mai_n439_), .B(mai_mai_n336_), .Y(mai_mai_n500_));
  INV        m478(.A(mai_mai_n274_), .Y(mai_mai_n501_));
  NO2        m479(.A(i_12_), .B(mai_mai_n77_), .Y(mai_mai_n502_));
  NA2        m480(.A(mai_mai_n502_), .B(mai_mai_n237_), .Y(mai_mai_n503_));
  NO2        m481(.A(mai_mai_n503_), .B(mai_mai_n501_), .Y(mai_mai_n504_));
  NO3        m482(.A(i_4_), .B(mai_mai_n299_), .C(mai_mai_n258_), .Y(mai_mai_n505_));
  NO3        m483(.A(mai_mai_n505_), .B(mai_mai_n504_), .C(mai_mai_n500_), .Y(mai_mai_n506_));
  NA4        m484(.A(mai_mai_n506_), .B(mai_mai_n499_), .C(mai_mai_n490_), .D(mai_mai_n480_), .Y(mai_mai_n507_));
  NO4        m485(.A(mai_mai_n507_), .B(mai_mai_n469_), .C(mai_mai_n449_), .D(mai_mai_n428_), .Y(mai_mai_n508_));
  NA4        m486(.A(mai_mai_n508_), .B(mai_mai_n377_), .C(mai_mai_n310_), .D(mai_mai_n268_), .Y(mai7));
  NO2        m487(.A(mai_mai_n85_), .B(mai_mai_n50_), .Y(mai_mai_n510_));
  NO2        m488(.A(mai_mai_n99_), .B(mai_mai_n82_), .Y(mai_mai_n511_));
  NA2        m489(.A(mai_mai_n342_), .B(mai_mai_n511_), .Y(mai_mai_n512_));
  NA2        m490(.A(mai_mai_n412_), .B(mai_mai_n76_), .Y(mai_mai_n513_));
  NA2        m491(.A(mai_mai_n132_), .B(i_8_), .Y(mai_mai_n514_));
  OAI210     m492(.A0(mai_mai_n514_), .A1(mai_mai_n513_), .B0(mai_mai_n512_), .Y(mai_mai_n515_));
  NA3        m493(.A(i_7_), .B(i_10_), .C(i_9_), .Y(mai_mai_n516_));
  NO2        m494(.A(mai_mai_n209_), .B(i_4_), .Y(mai_mai_n517_));
  NA2        m495(.A(mai_mai_n517_), .B(i_8_), .Y(mai_mai_n518_));
  NA2        m496(.A(i_2_), .B(mai_mai_n77_), .Y(mai_mai_n519_));
  NO2        m497(.A(i_7_), .B(mai_mai_n37_), .Y(mai_mai_n520_));
  NA2        m498(.A(i_4_), .B(i_8_), .Y(mai_mai_n521_));
  AOI210     m499(.A0(mai_mai_n521_), .A1(mai_mai_n263_), .B0(mai_mai_n520_), .Y(mai_mai_n522_));
  NO2        m500(.A(mai_mai_n522_), .B(mai_mai_n519_), .Y(mai_mai_n523_));
  NO3        m501(.A(mai_mai_n523_), .B(mai_mai_n515_), .C(mai_mai_n510_), .Y(mai_mai_n524_));
  AOI210     m502(.A0(mai_mai_n119_), .A1(mai_mai_n56_), .B0(i_10_), .Y(mai_mai_n525_));
  AOI210     m503(.A0(mai_mai_n525_), .A1(mai_mai_n209_), .B0(mai_mai_n145_), .Y(mai_mai_n526_));
  OR2        m504(.A(i_6_), .B(i_10_), .Y(mai_mai_n527_));
  NO2        m505(.A(mai_mai_n527_), .B(mai_mai_n23_), .Y(mai_mai_n528_));
  OR3        m506(.A(i_13_), .B(i_6_), .C(i_10_), .Y(mai_mai_n529_));
  NO3        m507(.A(mai_mai_n529_), .B(i_8_), .C(mai_mai_n31_), .Y(mai_mai_n530_));
  INV        m508(.A(mai_mai_n180_), .Y(mai_mai_n531_));
  NO2        m509(.A(mai_mai_n530_), .B(mai_mai_n528_), .Y(mai_mai_n532_));
  OA220      m510(.A0(mai_mai_n532_), .A1(mai_mai_n501_), .B0(mai_mai_n526_), .B1(mai_mai_n230_), .Y(mai_mai_n533_));
  AOI210     m511(.A0(mai_mai_n533_), .A1(mai_mai_n524_), .B0(mai_mai_n57_), .Y(mai_mai_n534_));
  NOi21      m512(.An(i_11_), .B(i_7_), .Y(mai_mai_n535_));
  AO210      m513(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(mai_mai_n536_));
  NO2        m514(.A(mai_mai_n536_), .B(mai_mai_n535_), .Y(mai_mai_n537_));
  NA3        m515(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n538_));
  NAi21      m516(.An(mai_mai_n538_), .B(i_11_), .Y(mai_mai_n539_));
  NO2        m517(.A(mai_mai_n539_), .B(mai_mai_n57_), .Y(mai_mai_n540_));
  NA2        m518(.A(mai_mai_n79_), .B(mai_mai_n57_), .Y(mai_mai_n541_));
  AO210      m519(.A0(mai_mai_n541_), .A1(mai_mai_n336_), .B0(mai_mai_n40_), .Y(mai_mai_n542_));
  NA2        m520(.A(mai_mai_n360_), .B(mai_mai_n31_), .Y(mai_mai_n543_));
  OR2        m521(.A(mai_mai_n186_), .B(mai_mai_n99_), .Y(mai_mai_n544_));
  NA2        m522(.A(mai_mai_n544_), .B(mai_mai_n543_), .Y(mai_mai_n545_));
  NO2        m523(.A(mai_mai_n57_), .B(i_9_), .Y(mai_mai_n546_));
  NA2        m524(.A(mai_mai_n57_), .B(mai_mai_n545_), .Y(mai_mai_n547_));
  NO2        m525(.A(i_1_), .B(i_12_), .Y(mai_mai_n548_));
  NA2        m526(.A(mai_mai_n547_), .B(mai_mai_n542_), .Y(mai_mai_n549_));
  OAI210     m527(.A0(mai_mai_n549_), .A1(mai_mai_n540_), .B0(i_6_), .Y(mai_mai_n550_));
  NO2        m528(.A(i_6_), .B(i_11_), .Y(mai_mai_n551_));
  INV        m529(.A(mai_mai_n390_), .Y(mai_mai_n552_));
  NO4        m530(.A(mai_mai_n193_), .B(mai_mai_n119_), .C(i_13_), .D(mai_mai_n77_), .Y(mai_mai_n553_));
  NA2        m531(.A(mai_mai_n209_), .B(i_6_), .Y(mai_mai_n554_));
  NA3        m532(.A(mai_mai_n457_), .B(i_11_), .C(mai_mai_n36_), .Y(mai_mai_n555_));
  NA2        m533(.A(mai_mai_n126_), .B(i_9_), .Y(mai_mai_n556_));
  NA3        m534(.A(i_3_), .B(i_8_), .C(i_9_), .Y(mai_mai_n557_));
  NO2        m535(.A(mai_mai_n46_), .B(i_1_), .Y(mai_mai_n558_));
  NA3        m536(.A(mai_mai_n558_), .B(mai_mai_n229_), .C(mai_mai_n44_), .Y(mai_mai_n559_));
  OAI220     m537(.A0(mai_mai_n559_), .A1(mai_mai_n557_), .B0(mai_mai_n556_), .B1(mai_mai_n901_), .Y(mai_mai_n560_));
  NA3        m538(.A(mai_mai_n546_), .B(mai_mai_n274_), .C(i_6_), .Y(mai_mai_n561_));
  NO2        m539(.A(mai_mai_n561_), .B(mai_mai_n23_), .Y(mai_mai_n562_));
  AOI210     m540(.A0(mai_mai_n404_), .A1(mai_mai_n366_), .B0(mai_mai_n213_), .Y(mai_mai_n563_));
  NO2        m541(.A(mai_mai_n563_), .B(mai_mai_n519_), .Y(mai_mai_n564_));
  NAi21      m542(.An(mai_mai_n555_), .B(mai_mai_n84_), .Y(mai_mai_n565_));
  NA2        m543(.A(mai_mai_n558_), .B(mai_mai_n229_), .Y(mai_mai_n566_));
  NO2        m544(.A(i_11_), .B(mai_mai_n37_), .Y(mai_mai_n567_));
  NA2        m545(.A(mai_mai_n567_), .B(mai_mai_n24_), .Y(mai_mai_n568_));
  OAI210     m546(.A0(mai_mai_n568_), .A1(mai_mai_n566_), .B0(mai_mai_n565_), .Y(mai_mai_n569_));
  OR4        m547(.A(mai_mai_n569_), .B(mai_mai_n564_), .C(mai_mai_n562_), .D(mai_mai_n560_), .Y(mai_mai_n570_));
  NO3        m548(.A(mai_mai_n570_), .B(mai_mai_n553_), .C(mai_mai_n552_), .Y(mai_mai_n571_));
  NA2        m549(.A(i_3_), .B(mai_mai_n174_), .Y(mai_mai_n572_));
  NO2        m550(.A(mai_mai_n572_), .B(mai_mai_n106_), .Y(mai_mai_n573_));
  AN2        m551(.A(mai_mai_n573_), .B(mai_mai_n459_), .Y(mai_mai_n574_));
  NO2        m552(.A(mai_mai_n207_), .B(mai_mai_n44_), .Y(mai_mai_n575_));
  NO2        m553(.A(mai_mai_n77_), .B(i_9_), .Y(mai_mai_n576_));
  NA2        m554(.A(i_1_), .B(i_3_), .Y(mai_mai_n577_));
  NO2        m555(.A(mai_mai_n391_), .B(mai_mai_n85_), .Y(mai_mai_n578_));
  AOI210     m556(.A0(mai_mai_n575_), .A1(mai_mai_n491_), .B0(mai_mai_n578_), .Y(mai_mai_n579_));
  NO2        m557(.A(mai_mai_n579_), .B(mai_mai_n577_), .Y(mai_mai_n580_));
  NO2        m558(.A(mai_mai_n580_), .B(mai_mai_n574_), .Y(mai_mai_n581_));
  NA3        m559(.A(mai_mai_n581_), .B(mai_mai_n571_), .C(mai_mai_n550_), .Y(mai_mai_n582_));
  NO3        m560(.A(mai_mai_n405_), .B(i_3_), .C(i_7_), .Y(mai_mai_n583_));
  NOi21      m561(.An(mai_mai_n583_), .B(i_10_), .Y(mai_mai_n584_));
  OA210      m562(.A0(mai_mai_n584_), .A1(mai_mai_n216_), .B0(mai_mai_n77_), .Y(mai_mai_n585_));
  NA2        m563(.A(mai_mai_n329_), .B(mai_mai_n328_), .Y(mai_mai_n586_));
  NA3        m564(.A(mai_mai_n412_), .B(mai_mai_n441_), .C(mai_mai_n46_), .Y(mai_mai_n587_));
  NO3        m565(.A(mai_mai_n406_), .B(mai_mai_n521_), .C(mai_mai_n77_), .Y(mai_mai_n588_));
  NA2        m566(.A(mai_mai_n588_), .B(mai_mai_n25_), .Y(mai_mai_n589_));
  NA3        m567(.A(mai_mai_n145_), .B(mai_mai_n76_), .C(mai_mai_n77_), .Y(mai_mai_n590_));
  NA4        m568(.A(mai_mai_n590_), .B(mai_mai_n589_), .C(mai_mai_n587_), .D(mai_mai_n586_), .Y(mai_mai_n591_));
  OAI210     m569(.A0(mai_mai_n591_), .A1(mai_mai_n585_), .B0(i_1_), .Y(mai_mai_n592_));
  AOI210     m570(.A0(mai_mai_n229_), .A1(mai_mai_n89_), .B0(i_1_), .Y(mai_mai_n593_));
  NO2        m571(.A(mai_mai_n327_), .B(i_2_), .Y(mai_mai_n594_));
  NA2        m572(.A(mai_mai_n594_), .B(mai_mai_n593_), .Y(mai_mai_n595_));
  OAI210     m573(.A0(mai_mai_n561_), .A1(mai_mai_n381_), .B0(mai_mai_n595_), .Y(mai_mai_n596_));
  INV        m574(.A(mai_mai_n596_), .Y(mai_mai_n597_));
  AOI210     m575(.A0(mai_mai_n597_), .A1(mai_mai_n592_), .B0(i_13_), .Y(mai_mai_n598_));
  OR2        m576(.A(i_11_), .B(i_7_), .Y(mai_mai_n599_));
  AOI220     m577(.A0(mai_mai_n400_), .A1(mai_mai_n145_), .B0(mai_mai_n384_), .B1(mai_mai_n126_), .Y(mai_mai_n600_));
  NO2        m578(.A(mai_mai_n600_), .B(mai_mai_n44_), .Y(mai_mai_n601_));
  NA2        m579(.A(mai_mai_n216_), .B(mai_mai_n122_), .Y(mai_mai_n602_));
  NO2        m580(.A(mai_mai_n602_), .B(mai_mai_n40_), .Y(mai_mai_n603_));
  AOI210     m581(.A0(mai_mai_n601_), .A1(mai_mai_n290_), .B0(mai_mai_n603_), .Y(mai_mai_n604_));
  AOI220     m582(.A0(i_7_), .A1(mai_mai_n65_), .B0(mai_mai_n344_), .B1(mai_mai_n558_), .Y(mai_mai_n605_));
  NO2        m583(.A(mai_mai_n605_), .B(mai_mai_n214_), .Y(mai_mai_n606_));
  AOI210     m584(.A0(mai_mai_n381_), .A1(mai_mai_n36_), .B0(i_13_), .Y(mai_mai_n607_));
  NOi31      m585(.An(mai_mai_n607_), .B(mai_mai_n513_), .C(mai_mai_n44_), .Y(mai_mai_n608_));
  NA2        m586(.A(mai_mai_n118_), .B(i_13_), .Y(mai_mai_n609_));
  NO2        m587(.A(mai_mai_n557_), .B(mai_mai_n106_), .Y(mai_mai_n610_));
  INV        m588(.A(mai_mai_n610_), .Y(mai_mai_n611_));
  OAI220     m589(.A0(mai_mai_n611_), .A1(mai_mai_n64_), .B0(mai_mai_n609_), .B1(mai_mai_n593_), .Y(mai_mai_n612_));
  NO3        m590(.A(mai_mai_n64_), .B(mai_mai_n32_), .C(mai_mai_n93_), .Y(mai_mai_n613_));
  NA2        m591(.A(mai_mai_n26_), .B(mai_mai_n174_), .Y(mai_mai_n614_));
  NA2        m592(.A(mai_mai_n614_), .B(i_7_), .Y(mai_mai_n615_));
  NO3        m593(.A(mai_mai_n406_), .B(mai_mai_n209_), .C(mai_mai_n77_), .Y(mai_mai_n616_));
  AOI210     m594(.A0(mai_mai_n616_), .A1(mai_mai_n615_), .B0(mai_mai_n613_), .Y(mai_mai_n617_));
  NA2        m595(.A(mai_mai_n84_), .B(mai_mai_n94_), .Y(mai_mai_n618_));
  OAI220     m596(.A0(mai_mai_n618_), .A1(mai_mai_n518_), .B0(mai_mai_n617_), .B1(mai_mai_n531_), .Y(mai_mai_n619_));
  NO4        m597(.A(mai_mai_n619_), .B(mai_mai_n612_), .C(mai_mai_n608_), .D(mai_mai_n606_), .Y(mai_mai_n620_));
  OR2        m598(.A(i_11_), .B(i_6_), .Y(mai_mai_n621_));
  NA3        m599(.A(mai_mai_n517_), .B(mai_mai_n614_), .C(i_7_), .Y(mai_mai_n622_));
  AOI210     m600(.A0(mai_mai_n622_), .A1(mai_mai_n611_), .B0(mai_mai_n621_), .Y(mai_mai_n623_));
  NA3        m601(.A(mai_mai_n360_), .B(mai_mai_n520_), .C(mai_mai_n89_), .Y(mai_mai_n624_));
  NA2        m602(.A(mai_mai_n551_), .B(i_13_), .Y(mai_mai_n625_));
  NA2        m603(.A(mai_mai_n94_), .B(mai_mai_n614_), .Y(mai_mai_n626_));
  NAi21      m604(.An(i_11_), .B(i_12_), .Y(mai_mai_n627_));
  NOi41      m605(.An(mai_mai_n102_), .B(mai_mai_n627_), .C(i_13_), .D(mai_mai_n77_), .Y(mai_mai_n628_));
  AOI220     m606(.A0(mai_mai_n910_), .A1(mai_mai_n269_), .B0(mai_mai_n628_), .B1(mai_mai_n626_), .Y(mai_mai_n629_));
  NA3        m607(.A(mai_mai_n629_), .B(mai_mai_n625_), .C(mai_mai_n624_), .Y(mai_mai_n630_));
  OAI210     m608(.A0(mai_mai_n630_), .A1(mai_mai_n623_), .B0(mai_mai_n57_), .Y(mai_mai_n631_));
  NO2        m609(.A(i_2_), .B(i_12_), .Y(mai_mai_n632_));
  NA2        m610(.A(mai_mai_n209_), .B(mai_mai_n326_), .Y(mai_mai_n633_));
  NO2        m611(.A(mai_mai_n119_), .B(i_2_), .Y(mai_mai_n634_));
  NA2        m612(.A(mai_mai_n634_), .B(mai_mai_n548_), .Y(mai_mai_n635_));
  NA2        m613(.A(mai_mai_n635_), .B(mai_mai_n633_), .Y(mai_mai_n636_));
  NA3        m614(.A(mai_mai_n636_), .B(mai_mai_n45_), .C(mai_mai_n201_), .Y(mai_mai_n637_));
  NA4        m615(.A(mai_mai_n637_), .B(mai_mai_n631_), .C(mai_mai_n620_), .D(mai_mai_n604_), .Y(mai_mai_n638_));
  OR4        m616(.A(mai_mai_n638_), .B(mai_mai_n598_), .C(mai_mai_n582_), .D(mai_mai_n534_), .Y(mai5));
  AN2        m617(.A(mai_mai_n24_), .B(i_10_), .Y(mai_mai_n640_));
  NA2        m618(.A(mai_mai_n640_), .B(mai_mai_n632_), .Y(mai_mai_n641_));
  NO2        m619(.A(mai_mai_n518_), .B(i_11_), .Y(mai_mai_n642_));
  NA2        m620(.A(mai_mai_n80_), .B(mai_mai_n642_), .Y(mai_mai_n643_));
  NA2        m621(.A(mai_mai_n643_), .B(mai_mai_n641_), .Y(mai_mai_n644_));
  NO3        m622(.A(i_11_), .B(mai_mai_n209_), .C(i_13_), .Y(mai_mai_n645_));
  NO2        m623(.A(mai_mai_n116_), .B(mai_mai_n23_), .Y(mai_mai_n646_));
  NA2        m624(.A(i_12_), .B(i_8_), .Y(mai_mai_n647_));
  INV        m625(.A(mai_mai_n380_), .Y(mai_mai_n648_));
  NA2        m626(.A(mai_mai_n274_), .B(mai_mai_n495_), .Y(mai_mai_n649_));
  INV        m627(.A(mai_mai_n649_), .Y(mai_mai_n650_));
  NO2        m628(.A(mai_mai_n650_), .B(mai_mai_n644_), .Y(mai_mai_n651_));
  INV        m629(.A(mai_mai_n153_), .Y(mai_mai_n652_));
  NA2        m630(.A(mai_mai_n594_), .B(mai_mai_n102_), .Y(mai_mai_n653_));
  NO2        m631(.A(mai_mai_n653_), .B(mai_mai_n652_), .Y(mai_mai_n654_));
  INV        m632(.A(mai_mai_n366_), .Y(mai_mai_n655_));
  NA2        m633(.A(mai_mai_n655_), .B(i_2_), .Y(mai_mai_n656_));
  INV        m634(.A(mai_mai_n656_), .Y(mai_mai_n657_));
  AOI210     m635(.A0(mai_mai_n33_), .A1(mai_mai_n36_), .B0(mai_mai_n363_), .Y(mai_mai_n658_));
  AOI210     m636(.A0(mai_mai_n658_), .A1(mai_mai_n657_), .B0(mai_mai_n654_), .Y(mai_mai_n659_));
  NO2        m637(.A(mai_mai_n171_), .B(mai_mai_n117_), .Y(mai_mai_n660_));
  OAI210     m638(.A0(mai_mai_n660_), .A1(mai_mai_n646_), .B0(i_2_), .Y(mai_mai_n661_));
  NA2        m639(.A(mai_mai_n153_), .B(mai_mai_n80_), .Y(mai_mai_n662_));
  AOI210     m640(.A0(mai_mai_n662_), .A1(mai_mai_n661_), .B0(mai_mai_n174_), .Y(mai_mai_n663_));
  AN2        m641(.A(mai_mai_n537_), .B(i_13_), .Y(mai_mai_n664_));
  NA2        m642(.A(mai_mai_n180_), .B(mai_mai_n182_), .Y(mai_mai_n665_));
  NA2        m643(.A(mai_mai_n75_), .B(i_8_), .Y(mai_mai_n666_));
  AOI210     m644(.A0(mai_mai_n666_), .A1(mai_mai_n665_), .B0(mai_mai_n330_), .Y(mai_mai_n667_));
  AOI210     m645(.A0(mai_mai_n186_), .A1(mai_mai_n136_), .B0(mai_mai_n441_), .Y(mai_mai_n668_));
  NA2        m646(.A(mai_mai_n668_), .B(mai_mai_n366_), .Y(mai_mai_n669_));
  INV        m647(.A(mai_mai_n259_), .Y(mai_mai_n670_));
  NA4        m648(.A(mai_mai_n670_), .B(mai_mai_n263_), .C(mai_mai_n116_), .D(mai_mai_n42_), .Y(mai_mai_n671_));
  NA2        m649(.A(mai_mai_n671_), .B(mai_mai_n669_), .Y(mai_mai_n672_));
  NO4        m650(.A(mai_mai_n672_), .B(mai_mai_n667_), .C(mai_mai_n664_), .D(mai_mai_n663_), .Y(mai_mai_n673_));
  NA2        m651(.A(mai_mai_n495_), .B(mai_mai_n28_), .Y(mai_mai_n674_));
  NA2        m652(.A(mai_mai_n645_), .B(mai_mai_n238_), .Y(mai_mai_n675_));
  NA2        m653(.A(mai_mai_n675_), .B(mai_mai_n674_), .Y(mai_mai_n676_));
  NA2        m654(.A(mai_mai_n676_), .B(mai_mai_n46_), .Y(mai_mai_n677_));
  NA4        m655(.A(mai_mai_n677_), .B(mai_mai_n673_), .C(mai_mai_n659_), .D(mai_mai_n651_), .Y(mai6));
  NO2        m656(.A(i_9_), .B(i_1_), .Y(mai_mai_n679_));
  INV        m657(.A(mai_mai_n127_), .Y(mai_mai_n680_));
  OAI210     m658(.A0(mai_mai_n680_), .A1(mai_mai_n679_), .B0(mai_mai_n634_), .Y(mai_mai_n681_));
  NA4        m659(.A(mai_mai_n347_), .B(mai_mai_n411_), .C(mai_mai_n64_), .D(mai_mai_n93_), .Y(mai_mai_n682_));
  INV        m660(.A(mai_mai_n682_), .Y(mai_mai_n683_));
  NO2        m661(.A(i_11_), .B(i_9_), .Y(mai_mai_n684_));
  NO2        m662(.A(mai_mai_n683_), .B(mai_mai_n286_), .Y(mai_mai_n685_));
  AO210      m663(.A0(mai_mai_n685_), .A1(mai_mai_n681_), .B0(i_12_), .Y(mai_mai_n686_));
  NA2        m664(.A(mai_mai_n331_), .B(mai_mai_n293_), .Y(mai_mai_n687_));
  NA2        m665(.A(mai_mai_n502_), .B(mai_mai_n57_), .Y(mai_mai_n688_));
  NA2        m666(.A(mai_mai_n584_), .B(mai_mai_n64_), .Y(mai_mai_n689_));
  NA4        m667(.A(mai_mai_n541_), .B(mai_mai_n689_), .C(mai_mai_n688_), .D(mai_mai_n687_), .Y(mai_mai_n690_));
  INV        m668(.A(mai_mai_n177_), .Y(mai_mai_n691_));
  AOI220     m669(.A0(mai_mai_n691_), .A1(mai_mai_n684_), .B0(mai_mai_n690_), .B1(mai_mai_n66_), .Y(mai_mai_n692_));
  INV        m670(.A(mai_mai_n285_), .Y(mai_mai_n693_));
  NA2        m671(.A(mai_mai_n68_), .B(mai_mai_n122_), .Y(mai_mai_n694_));
  NA2        m672(.A(mai_mai_n25_), .B(mai_mai_n46_), .Y(mai_mai_n695_));
  AOI210     m673(.A0(mai_mai_n695_), .A1(mai_mai_n694_), .B0(mai_mai_n693_), .Y(mai_mai_n696_));
  NO2        m674(.A(mai_mai_n32_), .B(i_11_), .Y(mai_mai_n697_));
  NA3        m675(.A(mai_mai_n697_), .B(mai_mai_n403_), .C(mai_mai_n347_), .Y(mai_mai_n698_));
  NAi32      m676(.An(i_1_), .Bn(i_9_), .C(i_5_), .Y(mai_mai_n699_));
  AOI210     m677(.A0(mai_mai_n621_), .A1(mai_mai_n78_), .B0(mai_mai_n699_), .Y(mai_mai_n700_));
  OAI210     m678(.A0(mai_mai_n583_), .A1(mai_mai_n483_), .B0(mai_mai_n482_), .Y(mai_mai_n701_));
  NAi31      m679(.An(mai_mai_n700_), .B(mai_mai_n701_), .C(mai_mai_n698_), .Y(mai_mai_n702_));
  OR2        m680(.A(mai_mai_n702_), .B(mai_mai_n696_), .Y(mai_mai_n703_));
  NO2        m681(.A(mai_mai_n599_), .B(i_2_), .Y(mai_mai_n704_));
  NA2        m682(.A(mai_mai_n916_), .B(mai_mai_n704_), .Y(mai_mai_n705_));
  AO220      m683(.A0(mai_mai_n315_), .A1(mai_mai_n306_), .B0(mai_mai_n352_), .B1(i_8_), .Y(mai_mai_n706_));
  NA3        m684(.A(mai_mai_n706_), .B(mai_mai_n222_), .C(i_7_), .Y(mai_mai_n707_));
  OR2        m685(.A(mai_mai_n537_), .B(mai_mai_n382_), .Y(mai_mai_n708_));
  NA2        m686(.A(mai_mai_n708_), .B(mai_mai_n135_), .Y(mai_mai_n709_));
  OR2        m687(.A(mai_mai_n648_), .B(mai_mai_n36_), .Y(mai_mai_n710_));
  NA4        m688(.A(mai_mai_n710_), .B(mai_mai_n709_), .C(mai_mai_n707_), .D(mai_mai_n705_), .Y(mai_mai_n711_));
  OAI210     m689(.A0(i_6_), .A1(i_11_), .B0(mai_mai_n78_), .Y(mai_mai_n712_));
  NA2        m690(.A(mai_mai_n712_), .B(mai_mai_n482_), .Y(mai_mai_n713_));
  NA3        m691(.A(mai_mai_n330_), .B(mai_mai_n210_), .C(mai_mai_n135_), .Y(mai_mai_n714_));
  NA2        m692(.A(mai_mai_n352_), .B(mai_mai_n63_), .Y(mai_mai_n715_));
  NA3        m693(.A(mai_mai_n715_), .B(mai_mai_n714_), .C(mai_mai_n713_), .Y(mai_mai_n716_));
  AO210      m694(.A0(mai_mai_n441_), .A1(mai_mai_n46_), .B0(mai_mai_n79_), .Y(mai_mai_n717_));
  NA2        m695(.A(mai_mai_n717_), .B(mai_mai_n412_), .Y(mai_mai_n718_));
  AOI210     m696(.A0(mai_mai_n382_), .A1(mai_mai_n380_), .B0(mai_mai_n481_), .Y(mai_mai_n719_));
  NA2        m697(.A(mai_mai_n103_), .B(mai_mai_n359_), .Y(mai_mai_n720_));
  NA3        m698(.A(mai_mai_n720_), .B(mai_mai_n719_), .C(mai_mai_n718_), .Y(mai_mai_n721_));
  NO4        m699(.A(mai_mai_n721_), .B(mai_mai_n716_), .C(mai_mai_n711_), .D(mai_mai_n703_), .Y(mai_mai_n722_));
  NA4        m700(.A(mai_mai_n722_), .B(mai_mai_n692_), .C(mai_mai_n686_), .D(mai_mai_n338_), .Y(mai3));
  NA2        m701(.A(i_6_), .B(i_7_), .Y(mai_mai_n724_));
  NO2        m702(.A(mai_mai_n724_), .B(i_0_), .Y(mai_mai_n725_));
  NO2        m703(.A(i_11_), .B(mai_mai_n209_), .Y(mai_mai_n726_));
  OAI210     m704(.A0(mai_mai_n725_), .A1(mai_mai_n248_), .B0(mai_mai_n726_), .Y(mai_mai_n727_));
  NO2        m705(.A(mai_mai_n727_), .B(mai_mai_n174_), .Y(mai_mai_n728_));
  NO3        m706(.A(mai_mai_n387_), .B(mai_mai_n82_), .C(mai_mai_n44_), .Y(mai_mai_n729_));
  OA210      m707(.A0(mai_mai_n729_), .A1(mai_mai_n728_), .B0(mai_mai_n156_), .Y(mai_mai_n730_));
  INV        m708(.A(mai_mai_n714_), .Y(mai_mai_n731_));
  NA2        m709(.A(mai_mai_n731_), .B(mai_mai_n39_), .Y(mai_mai_n732_));
  NO2        m710(.A(mai_mai_n544_), .B(mai_mai_n391_), .Y(mai_mai_n733_));
  AOI210     m711(.A0(mai_mai_n902_), .A1(mai_mai_n732_), .B0(mai_mai_n48_), .Y(mai_mai_n734_));
  NA2        m712(.A(mai_mai_n607_), .B(mai_mai_n576_), .Y(mai_mai_n735_));
  NA2        m713(.A(mai_mai_n291_), .B(i_5_), .Y(mai_mai_n736_));
  NO2        m714(.A(mai_mai_n736_), .B(mai_mai_n735_), .Y(mai_mai_n737_));
  NOi21      m715(.An(i_5_), .B(i_9_), .Y(mai_mai_n738_));
  NA2        m716(.A(mai_mai_n738_), .B(i_0_), .Y(mai_mai_n739_));
  AOI210     m717(.A0(mai_mai_n229_), .A1(mai_mai_n404_), .B0(mai_mai_n588_), .Y(mai_mai_n740_));
  NO2        m718(.A(mai_mai_n157_), .B(mai_mai_n136_), .Y(mai_mai_n741_));
  NA2        m719(.A(mai_mai_n741_), .B(mai_mai_n215_), .Y(mai_mai_n742_));
  OAI220     m720(.A0(mai_mai_n742_), .A1(mai_mai_n162_), .B0(mai_mai_n740_), .B1(mai_mai_n739_), .Y(mai_mai_n743_));
  NO4        m721(.A(mai_mai_n743_), .B(mai_mai_n737_), .C(mai_mai_n734_), .D(mai_mai_n730_), .Y(mai_mai_n744_));
  NA2        m722(.A(mai_mai_n167_), .B(mai_mai_n24_), .Y(mai_mai_n745_));
  NO2        m723(.A(mai_mai_n37_), .B(mai_mai_n745_), .Y(mai_mai_n746_));
  NA2        m724(.A(mai_mai_n269_), .B(mai_mai_n120_), .Y(mai_mai_n747_));
  NAi21      m725(.An(mai_mai_n146_), .B(i_5_), .Y(mai_mai_n748_));
  NO2        m726(.A(mai_mai_n747_), .B(mai_mai_n353_), .Y(mai_mai_n749_));
  NO2        m727(.A(mai_mai_n749_), .B(mai_mai_n746_), .Y(mai_mai_n750_));
  NA2        m728(.A(mai_mai_n492_), .B(i_0_), .Y(mai_mai_n751_));
  NO3        m729(.A(mai_mai_n751_), .B(mai_mai_n343_), .C(mai_mai_n80_), .Y(mai_mai_n752_));
  INV        m730(.A(mai_mai_n752_), .Y(mai_mai_n753_));
  NA2        m731(.A(mai_mai_n645_), .B(mai_mai_n286_), .Y(mai_mai_n754_));
  OAI220     m732(.A0(i_6_), .A1(mai_mai_n754_), .B0(mai_mai_n568_), .B1(mai_mai_n57_), .Y(mai_mai_n755_));
  NO4        m733(.A(mai_mai_n106_), .B(mai_mai_n52_), .C(mai_mai_n572_), .D(i_5_), .Y(mai_mai_n756_));
  AN2        m734(.A(mai_mai_n756_), .B(i_10_), .Y(mai_mai_n757_));
  NA2        m735(.A(mai_mai_n167_), .B(mai_mai_n76_), .Y(mai_mai_n758_));
  NA2        m736(.A(mai_mai_n486_), .B(i_4_), .Y(mai_mai_n759_));
  NA2        m737(.A(mai_mai_n170_), .B(mai_mai_n182_), .Y(mai_mai_n760_));
  OAI220     m738(.A0(mai_mai_n760_), .A1(mai_mai_n754_), .B0(mai_mai_n759_), .B1(mai_mai_n758_), .Y(mai_mai_n761_));
  NO3        m739(.A(mai_mai_n761_), .B(mai_mai_n757_), .C(mai_mai_n755_), .Y(mai_mai_n762_));
  NA3        m740(.A(mai_mai_n762_), .B(mai_mai_n753_), .C(mai_mai_n750_), .Y(mai_mai_n763_));
  NA2        m741(.A(i_11_), .B(i_9_), .Y(mai_mai_n764_));
  NO3        m742(.A(i_12_), .B(mai_mai_n764_), .C(mai_mai_n519_), .Y(mai_mai_n765_));
  AN2        m743(.A(mai_mai_n765_), .B(i_10_), .Y(mai_mai_n766_));
  NO2        m744(.A(mai_mai_n48_), .B(i_7_), .Y(mai_mai_n767_));
  NA2        m745(.A(mai_mai_n351_), .B(mai_mai_n161_), .Y(mai_mai_n768_));
  NA2        m746(.A(mai_mai_n768_), .B(mai_mai_n144_), .Y(mai_mai_n769_));
  NO2        m747(.A(mai_mai_n157_), .B(i_0_), .Y(mai_mai_n770_));
  NA2        m748(.A(mai_mai_n403_), .B(mai_mai_n205_), .Y(mai_mai_n771_));
  NA2        m749(.A(mai_mai_n329_), .B(mai_mai_n41_), .Y(mai_mai_n772_));
  OAI220     m750(.A0(mai_mai_n772_), .A1(mai_mai_n739_), .B0(mai_mai_n771_), .B1(mai_mai_n157_), .Y(mai_mai_n773_));
  NO3        m751(.A(mai_mai_n773_), .B(mai_mai_n769_), .C(mai_mai_n766_), .Y(mai_mai_n774_));
  NA2        m752(.A(mai_mai_n567_), .B(mai_mai_n113_), .Y(mai_mai_n775_));
  NO2        m753(.A(i_6_), .B(mai_mai_n775_), .Y(mai_mai_n776_));
  AOI210     m754(.A0(mai_mai_n381_), .A1(mai_mai_n36_), .B0(i_3_), .Y(mai_mai_n777_));
  NA2        m755(.A(mai_mai_n153_), .B(mai_mai_n95_), .Y(mai_mai_n778_));
  NOi32      m756(.An(mai_mai_n777_), .Bn(mai_mai_n170_), .C(mai_mai_n778_), .Y(mai_mai_n779_));
  NA2        m757(.A(mai_mai_n520_), .B(mai_mai_n286_), .Y(mai_mai_n780_));
  NO2        m758(.A(mai_mai_n780_), .B(i_12_), .Y(mai_mai_n781_));
  NO3        m759(.A(mai_mai_n781_), .B(mai_mai_n779_), .C(mai_mai_n776_), .Y(mai_mai_n782_));
  NOi21      m760(.An(i_7_), .B(i_5_), .Y(mai_mai_n783_));
  NOi31      m761(.An(mai_mai_n783_), .B(i_0_), .C(mai_mai_n627_), .Y(mai_mai_n784_));
  NA3        m762(.A(mai_mai_n784_), .B(mai_mai_n342_), .C(i_6_), .Y(mai_mai_n785_));
  OA210      m763(.A0(mai_mai_n778_), .A1(mai_mai_n440_), .B0(mai_mai_n785_), .Y(mai_mai_n786_));
  NO3        m764(.A(mai_mai_n356_), .B(mai_mai_n318_), .C(mai_mai_n314_), .Y(mai_mai_n787_));
  NO2        m765(.A(mai_mai_n225_), .B(mai_mai_n275_), .Y(mai_mai_n788_));
  NO2        m766(.A(mai_mai_n627_), .B(mai_mai_n224_), .Y(mai_mai_n789_));
  AOI210     m767(.A0(mai_mai_n789_), .A1(mai_mai_n788_), .B0(mai_mai_n787_), .Y(mai_mai_n790_));
  NA4        m768(.A(mai_mai_n790_), .B(mai_mai_n786_), .C(mai_mai_n782_), .D(mai_mai_n774_), .Y(mai_mai_n791_));
  AN2        m769(.A(mai_mai_n290_), .B(mai_mai_n741_), .Y(mai_mai_n792_));
  NA2        m770(.A(mai_mai_n792_), .B(i_10_), .Y(mai_mai_n793_));
  NA3        m771(.A(mai_mai_n402_), .B(mai_mai_n360_), .C(mai_mai_n45_), .Y(mai_mai_n794_));
  OAI210     m772(.A0(mai_mai_n748_), .A1(i_6_), .B0(mai_mai_n794_), .Y(mai_mai_n795_));
  NA2        m773(.A(i_9_), .B(mai_mai_n263_), .Y(mai_mai_n796_));
  NA2        m774(.A(mai_mai_n169_), .B(mai_mai_n796_), .Y(mai_mai_n797_));
  AOI220     m775(.A0(mai_mai_n797_), .A1(mai_mai_n403_), .B0(mai_mai_n795_), .B1(mai_mai_n66_), .Y(mai_mai_n798_));
  NO2        m776(.A(mai_mai_n68_), .B(mai_mai_n647_), .Y(mai_mai_n799_));
  AOI210     m777(.A0(mai_mai_n156_), .A1(mai_mai_n511_), .B0(mai_mai_n799_), .Y(mai_mai_n800_));
  NO2        m778(.A(mai_mai_n800_), .B(mai_mai_n47_), .Y(mai_mai_n801_));
  NO3        m779(.A(i_5_), .B(mai_mai_n313_), .C(mai_mai_n24_), .Y(mai_mai_n802_));
  NO2        m780(.A(mai_mai_n465_), .B(mai_mai_n802_), .Y(mai_mai_n803_));
  NAi21      m781(.An(i_9_), .B(i_5_), .Y(mai_mai_n804_));
  NO2        m782(.A(mai_mai_n804_), .B(mai_mai_n356_), .Y(mai_mai_n805_));
  NO2        m783(.A(mai_mai_n516_), .B(mai_mai_n96_), .Y(mai_mai_n806_));
  AOI220     m784(.A0(mai_mai_n806_), .A1(i_0_), .B0(mai_mai_n805_), .B1(mai_mai_n537_), .Y(mai_mai_n807_));
  OAI220     m785(.A0(mai_mai_n807_), .A1(mai_mai_n77_), .B0(mai_mai_n803_), .B1(mai_mai_n154_), .Y(mai_mai_n808_));
  NO2        m786(.A(mai_mai_n808_), .B(mai_mai_n801_), .Y(mai_mai_n809_));
  NA3        m787(.A(mai_mai_n809_), .B(mai_mai_n798_), .C(mai_mai_n793_), .Y(mai_mai_n810_));
  NO3        m788(.A(mai_mai_n810_), .B(mai_mai_n791_), .C(mai_mai_n763_), .Y(mai_mai_n811_));
  NO2        m789(.A(i_0_), .B(mai_mai_n627_), .Y(mai_mai_n812_));
  INV        m790(.A(i_0_), .Y(mai_mai_n813_));
  NO2        m791(.A(i_5_), .B(mai_mai_n25_), .Y(mai_mai_n814_));
  AO220      m792(.A0(mai_mai_n814_), .A1(mai_mai_n813_), .B0(mai_mai_n812_), .B1(mai_mai_n156_), .Y(mai_mai_n815_));
  AOI210     m793(.A0(mai_mai_n688_), .A1(mai_mai_n586_), .B0(mai_mai_n778_), .Y(mai_mai_n816_));
  AOI210     m794(.A0(mai_mai_n815_), .A1(mai_mai_n304_), .B0(mai_mai_n816_), .Y(mai_mai_n817_));
  NA3        m795(.A(mai_mai_n134_), .B(mai_mai_n576_), .C(mai_mai_n66_), .Y(mai_mai_n818_));
  NO2        m796(.A(mai_mai_n701_), .B(mai_mai_n356_), .Y(mai_mai_n819_));
  NA3        m797(.A(mai_mai_n725_), .B(i_2_), .C(mai_mai_n48_), .Y(mai_mai_n820_));
  NA2        m798(.A(mai_mai_n726_), .B(i_9_), .Y(mai_mai_n821_));
  AOI210     m799(.A0(mai_mai_n820_), .A1(mai_mai_n422_), .B0(mai_mai_n821_), .Y(mai_mai_n822_));
  OAI210     m800(.A0(mai_mai_n215_), .A1(i_9_), .B0(mai_mai_n204_), .Y(mai_mai_n823_));
  AOI210     m801(.A0(mai_mai_n823_), .A1(mai_mai_n751_), .B0(mai_mai_n139_), .Y(mai_mai_n824_));
  NO3        m802(.A(mai_mai_n824_), .B(mai_mai_n822_), .C(mai_mai_n819_), .Y(mai_mai_n825_));
  NA3        m803(.A(mai_mai_n825_), .B(mai_mai_n818_), .C(mai_mai_n817_), .Y(mai_mai_n826_));
  NA3        m804(.A(mai_mai_n39_), .B(mai_mai_n28_), .C(mai_mai_n44_), .Y(mai_mai_n827_));
  NA2        m805(.A(mai_mai_n767_), .B(mai_mai_n415_), .Y(mai_mai_n828_));
  AOI210     m806(.A0(mai_mai_n827_), .A1(mai_mai_n146_), .B0(mai_mai_n828_), .Y(mai_mai_n829_));
  INV        m807(.A(mai_mai_n829_), .Y(mai_mai_n830_));
  NA2        m808(.A(mai_mai_n487_), .B(mai_mai_n68_), .Y(mai_mai_n831_));
  NO3        m809(.A(mai_mai_n187_), .B(mai_mai_n341_), .C(i_0_), .Y(mai_mai_n832_));
  OAI210     m810(.A0(mai_mai_n832_), .A1(mai_mai_n69_), .B0(i_13_), .Y(mai_mai_n833_));
  INV        m811(.A(mai_mai_n195_), .Y(mai_mai_n834_));
  OAI220     m812(.A0(mai_mai_n453_), .A1(mai_mai_n127_), .B0(mai_mai_n554_), .B1(mai_mai_n531_), .Y(mai_mai_n835_));
  NA3        m813(.A(mai_mai_n835_), .B(i_7_), .C(mai_mai_n834_), .Y(mai_mai_n836_));
  NA4        m814(.A(mai_mai_n836_), .B(mai_mai_n833_), .C(mai_mai_n831_), .D(mai_mai_n830_), .Y(mai_mai_n837_));
  NO2        m815(.A(mai_mai_n214_), .B(mai_mai_n85_), .Y(mai_mai_n838_));
  AOI210     m816(.A0(mai_mai_n838_), .A1(mai_mai_n812_), .B0(mai_mai_n100_), .Y(mai_mai_n839_));
  NA2        m817(.A(mai_mai_n783_), .B(mai_mai_n415_), .Y(mai_mai_n840_));
  NA2        m818(.A(mai_mai_n306_), .B(mai_mai_n158_), .Y(mai_mai_n841_));
  OA220      m819(.A0(mai_mai_n841_), .A1(mai_mai_n840_), .B0(mai_mai_n839_), .B1(i_5_), .Y(mai_mai_n842_));
  AOI210     m820(.A0(i_0_), .A1(mai_mai_n25_), .B0(mai_mai_n157_), .Y(mai_mai_n843_));
  NA2        m821(.A(mai_mai_n843_), .B(mai_mai_n402_), .Y(mai_mai_n844_));
  NA3        m822(.A(mai_mai_n347_), .B(mai_mai_n292_), .C(mai_mai_n197_), .Y(mai_mai_n845_));
  INV        m823(.A(mai_mai_n845_), .Y(mai_mai_n846_));
  NOi31      m824(.An(mai_mai_n346_), .B(i_0_), .C(mai_mai_n211_), .Y(mai_mai_n847_));
  NO3        m825(.A(mai_mai_n764_), .B(mai_mai_n195_), .C(mai_mai_n171_), .Y(mai_mai_n848_));
  NO3        m826(.A(mai_mai_n848_), .B(mai_mai_n847_), .C(mai_mai_n846_), .Y(mai_mai_n849_));
  NA4        m827(.A(mai_mai_n849_), .B(mai_mai_n401_), .C(mai_mai_n844_), .D(mai_mai_n842_), .Y(mai_mai_n850_));
  NA3        m828(.A(mai_mai_n263_), .B(i_5_), .C(mai_mai_n174_), .Y(mai_mai_n851_));
  NA2        m829(.A(mai_mai_n851_), .B(mai_mai_n214_), .Y(mai_mai_n852_));
  NO3        m830(.A(mai_mai_n211_), .B(i_0_), .C(i_12_), .Y(mai_mai_n853_));
  AOI220     m831(.A0(mai_mai_n853_), .A1(mai_mai_n852_), .B0(mai_mai_n683_), .B1(mai_mai_n158_), .Y(mai_mai_n854_));
  NO3        m832(.A(mai_mai_n911_), .B(i_12_), .C(mai_mai_n555_), .Y(mai_mai_n855_));
  INV        m833(.A(mai_mai_n855_), .Y(mai_mai_n856_));
  NA3        m834(.A(mai_mai_n90_), .B(mai_mai_n491_), .C(i_11_), .Y(mai_mai_n857_));
  NA2        m835(.A(mai_mai_n783_), .B(mai_mai_n400_), .Y(mai_mai_n858_));
  NO2        m836(.A(mai_mai_n858_), .B(i_1_), .Y(mai_mai_n859_));
  NA2        m837(.A(mai_mai_n859_), .B(mai_mai_n770_), .Y(mai_mai_n860_));
  NA3        m838(.A(mai_mai_n860_), .B(mai_mai_n856_), .C(mai_mai_n854_), .Y(mai_mai_n861_));
  NO4        m839(.A(mai_mai_n861_), .B(mai_mai_n850_), .C(mai_mai_n837_), .D(mai_mai_n826_), .Y(mai_mai_n862_));
  OAI210     m840(.A0(mai_mai_n704_), .A1(mai_mai_n697_), .B0(mai_mai_n37_), .Y(mai_mai_n863_));
  NA3        m841(.A(mai_mai_n777_), .B(mai_mai_n326_), .C(i_5_), .Y(mai_mai_n864_));
  NA3        m842(.A(mai_mai_n864_), .B(mai_mai_n863_), .C(mai_mai_n526_), .Y(mai_mai_n865_));
  NA2        m843(.A(mai_mai_n865_), .B(mai_mai_n185_), .Y(mai_mai_n866_));
  NA2        m844(.A(mai_mai_n168_), .B(mai_mai_n170_), .Y(mai_mai_n867_));
  OR2        m845(.A(i_11_), .B(mai_mai_n867_), .Y(mai_mai_n868_));
  OAI210     m846(.A0(mai_mai_n530_), .A1(mai_mai_n528_), .B0(mai_mai_n274_), .Y(mai_mai_n869_));
  NA2        m847(.A(mai_mai_n869_), .B(mai_mai_n868_), .Y(mai_mai_n870_));
  NO2        m848(.A(mai_mai_n394_), .B(mai_mai_n229_), .Y(mai_mai_n871_));
  INV        m849(.A(mai_mai_n871_), .Y(mai_mai_n872_));
  NA2        m850(.A(mai_mai_n857_), .B(mai_mai_n872_), .Y(mai_mai_n873_));
  AOI210     m851(.A0(mai_mai_n870_), .A1(mai_mai_n48_), .B0(mai_mai_n873_), .Y(mai_mai_n874_));
  AOI210     m852(.A0(mai_mai_n874_), .A1(mai_mai_n866_), .B0(mai_mai_n66_), .Y(mai_mai_n875_));
  NO2        m853(.A(mai_mai_n484_), .B(mai_mai_n337_), .Y(mai_mai_n876_));
  NO2        m854(.A(mai_mai_n876_), .B(mai_mai_n652_), .Y(mai_mai_n877_));
  INV        m855(.A(mai_mai_n69_), .Y(mai_mai_n878_));
  AOI210     m856(.A0(mai_mai_n843_), .A1(mai_mai_n767_), .B0(mai_mai_n784_), .Y(mai_mai_n879_));
  AOI210     m857(.A0(mai_mai_n879_), .A1(mai_mai_n878_), .B0(mai_mai_n577_), .Y(mai_mai_n880_));
  NA2        m858(.A(i_8_), .B(mai_mai_n69_), .Y(mai_mai_n881_));
  NO2        m859(.A(mai_mai_n881_), .B(mai_mai_n209_), .Y(mai_mai_n882_));
  NO2        m860(.A(mai_mai_n882_), .B(mai_mai_n880_), .Y(mai_mai_n883_));
  OAI210     m861(.A0(mai_mai_n231_), .A1(mai_mai_n142_), .B0(mai_mai_n80_), .Y(mai_mai_n884_));
  NO2        m862(.A(mai_mai_n884_), .B(i_11_), .Y(mai_mai_n885_));
  OAI210     m863(.A0(mai_mai_n903_), .A1(mai_mai_n777_), .B0(mai_mai_n185_), .Y(mai_mai_n886_));
  NA2        m864(.A(mai_mai_n148_), .B(i_5_), .Y(mai_mai_n887_));
  AOI210     m865(.A0(mai_mai_n886_), .A1(mai_mai_n665_), .B0(mai_mai_n887_), .Y(mai_mai_n888_));
  NA2        m866(.A(mai_mai_n788_), .B(mai_mai_n904_), .Y(mai_mai_n889_));
  NO2        m867(.A(mai_mai_n889_), .B(mai_mai_n627_), .Y(mai_mai_n890_));
  NO3        m868(.A(mai_mai_n804_), .B(mai_mai_n405_), .C(mai_mai_n221_), .Y(mai_mai_n891_));
  NO2        m869(.A(mai_mai_n891_), .B(mai_mai_n481_), .Y(mai_mai_n892_));
  INV        m870(.A(mai_mai_n319_), .Y(mai_mai_n893_));
  AOI210     m871(.A0(mai_mai_n893_), .A1(mai_mai_n892_), .B0(mai_mai_n40_), .Y(mai_mai_n894_));
  NO4        m872(.A(mai_mai_n894_), .B(mai_mai_n890_), .C(mai_mai_n888_), .D(mai_mai_n885_), .Y(mai_mai_n895_));
  OAI210     m873(.A0(mai_mai_n883_), .A1(i_4_), .B0(mai_mai_n895_), .Y(mai_mai_n896_));
  NO3        m874(.A(mai_mai_n896_), .B(mai_mai_n877_), .C(mai_mai_n875_), .Y(mai_mai_n897_));
  NA4        m875(.A(mai_mai_n897_), .B(mai_mai_n862_), .C(mai_mai_n811_), .D(mai_mai_n744_), .Y(mai4));
  INV        m876(.A(i_2_), .Y(mai_mai_n901_));
  INV        m877(.A(mai_mai_n733_), .Y(mai_mai_n902_));
  INV        m878(.A(i_12_), .Y(mai_mai_n903_));
  INV        m879(.A(i_4_), .Y(mai_mai_n904_));
  INV        m880(.A(mai_mai_n217_), .Y(mai_mai_n905_));
  INV        m881(.A(mai_mai_n130_), .Y(mai_mai_n906_));
  INV        m882(.A(i_5_), .Y(mai_mai_n907_));
  INV        m883(.A(i_2_), .Y(mai_mai_n908_));
  INV        m884(.A(i_3_), .Y(mai_mai_n909_));
  INV        m885(.A(mai_mai_n521_), .Y(mai_mai_n910_));
  INV        m886(.A(i_10_), .Y(mai_mai_n911_));
  INV        m887(.A(mai_mai_n178_), .Y(mai_mai_n912_));
  INV        m888(.A(mai_mai_n143_), .Y(mai_mai_n913_));
  INV        m889(.A(mai_mai_n196_), .Y(mai_mai_n914_));
  INV        m890(.A(i_10_), .Y(mai_mai_n915_));
  INV        m891(.A(i_5_), .Y(mai_mai_n916_));
  INV        m892(.A(i_13_), .Y(mai_mai_n917_));
  NAi21      u000(.An(i_13_), .B(i_4_), .Y(men_men_n23_));
  NOi21      u001(.An(i_3_), .B(i_8_), .Y(men_men_n24_));
  INV        u002(.A(i_9_), .Y(men_men_n25_));
  INV        u003(.A(i_3_), .Y(men_men_n26_));
  NO2        u004(.A(men_men_n26_), .B(men_men_n25_), .Y(men_men_n27_));
  NO2        u005(.A(i_8_), .B(i_10_), .Y(men_men_n28_));
  INV        u006(.A(men_men_n28_), .Y(men_men_n29_));
  OAI210     u007(.A0(men_men_n27_), .A1(men_men_n24_), .B0(men_men_n29_), .Y(men_men_n30_));
  NOi21      u008(.An(i_11_), .B(i_8_), .Y(men_men_n31_));
  AO210      u009(.A0(i_12_), .A1(i_8_), .B0(i_3_), .Y(men_men_n32_));
  OR2        u010(.A(men_men_n32_), .B(men_men_n31_), .Y(men_men_n33_));
  NA2        u011(.A(men_men_n33_), .B(men_men_n30_), .Y(men_men_n34_));
  XO2        u012(.A(men_men_n34_), .B(men_men_n23_), .Y(men_men_n35_));
  INV        u013(.A(i_4_), .Y(men_men_n36_));
  INV        u014(.A(i_10_), .Y(men_men_n37_));
  NAi21      u015(.An(i_11_), .B(i_9_), .Y(men_men_n38_));
  NOi21      u016(.An(i_12_), .B(i_13_), .Y(men_men_n39_));
  INV        u017(.A(men_men_n39_), .Y(men_men_n40_));
  NAi31      u018(.An(i_9_), .B(i_4_), .C(i_8_), .Y(men_men_n41_));
  INV        u019(.A(men_men_n35_), .Y(men1));
  INV        u020(.A(i_11_), .Y(men_men_n43_));
  NO2        u021(.A(men_men_n43_), .B(i_6_), .Y(men_men_n44_));
  INV        u022(.A(i_2_), .Y(men_men_n45_));
  NA2        u023(.A(i_0_), .B(i_3_), .Y(men_men_n46_));
  INV        u024(.A(i_5_), .Y(men_men_n47_));
  NO2        u025(.A(i_7_), .B(i_10_), .Y(men_men_n48_));
  AOI210     u026(.A0(i_7_), .A1(men_men_n25_), .B0(men_men_n48_), .Y(men_men_n49_));
  OAI210     u027(.A0(men_men_n49_), .A1(i_3_), .B0(men_men_n47_), .Y(men_men_n50_));
  AOI210     u028(.A0(men_men_n50_), .A1(men_men_n46_), .B0(men_men_n45_), .Y(men_men_n51_));
  NA2        u029(.A(i_0_), .B(i_2_), .Y(men_men_n52_));
  NA2        u030(.A(i_7_), .B(i_9_), .Y(men_men_n53_));
  NO2        u031(.A(men_men_n53_), .B(men_men_n52_), .Y(men_men_n54_));
  NA2        u032(.A(men_men_n51_), .B(men_men_n44_), .Y(men_men_n55_));
  NA3        u033(.A(i_2_), .B(i_6_), .C(i_8_), .Y(men_men_n56_));
  NO2        u034(.A(i_1_), .B(i_6_), .Y(men_men_n57_));
  NA2        u035(.A(i_8_), .B(i_7_), .Y(men_men_n58_));
  NA2        u036(.A(i_6_), .B(i_12_), .Y(men_men_n59_));
  NAi21      u037(.An(i_2_), .B(i_7_), .Y(men_men_n60_));
  INV        u038(.A(i_1_), .Y(men_men_n61_));
  NA2        u039(.A(men_men_n61_), .B(i_6_), .Y(men_men_n62_));
  NA3        u040(.A(men_men_n62_), .B(men_men_n60_), .C(men_men_n31_), .Y(men_men_n63_));
  NA2        u041(.A(men_men_n63_), .B(men_men_n59_), .Y(men_men_n64_));
  NA2        u042(.A(men_men_n49_), .B(i_2_), .Y(men_men_n65_));
  AOI210     u043(.A0(i_12_), .A1(i_6_), .B0(i_1_), .Y(men_men_n66_));
  NA2        u044(.A(i_1_), .B(i_6_), .Y(men_men_n67_));
  NO2        u045(.A(men_men_n67_), .B(men_men_n25_), .Y(men_men_n68_));
  INV        u046(.A(i_0_), .Y(men_men_n69_));
  NAi21      u047(.An(i_5_), .B(i_10_), .Y(men_men_n70_));
  NA2        u048(.A(i_5_), .B(i_9_), .Y(men_men_n71_));
  AOI210     u049(.A0(men_men_n71_), .A1(men_men_n70_), .B0(men_men_n69_), .Y(men_men_n72_));
  NO2        u050(.A(men_men_n72_), .B(men_men_n68_), .Y(men_men_n73_));
  OAI210     u051(.A0(men_men_n66_), .A1(men_men_n65_), .B0(men_men_n73_), .Y(men_men_n74_));
  OAI210     u052(.A0(men_men_n74_), .A1(men_men_n64_), .B0(i_0_), .Y(men_men_n75_));
  NA2        u053(.A(i_12_), .B(i_5_), .Y(men_men_n76_));
  NA2        u054(.A(i_2_), .B(i_8_), .Y(men_men_n77_));
  NO2        u055(.A(i_3_), .B(i_9_), .Y(men_men_n78_));
  NO2        u056(.A(i_3_), .B(i_7_), .Y(men_men_n79_));
  NO2        u057(.A(men_men_n79_), .B(men_men_n61_), .Y(men_men_n80_));
  INV        u058(.A(i_6_), .Y(men_men_n81_));
  OR4        u059(.A(i_2_), .B(i_11_), .C(i_3_), .D(i_8_), .Y(men_men_n82_));
  INV        u060(.A(men_men_n82_), .Y(men_men_n83_));
  NO2        u061(.A(i_2_), .B(i_7_), .Y(men_men_n84_));
  NA2        u062(.A(men_men_n80_), .B(men_men_n82_), .Y(men_men_n85_));
  NAi21      u063(.An(i_6_), .B(i_10_), .Y(men_men_n86_));
  NA2        u064(.A(i_6_), .B(i_9_), .Y(men_men_n87_));
  NA2        u065(.A(i_2_), .B(i_6_), .Y(men_men_n88_));
  NO3        u066(.A(men_men_n88_), .B(men_men_n48_), .C(men_men_n25_), .Y(men_men_n89_));
  INV        u067(.A(men_men_n89_), .Y(men_men_n90_));
  AOI210     u068(.A0(men_men_n90_), .A1(men_men_n85_), .B0(men_men_n76_), .Y(men_men_n91_));
  AN3        u069(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n92_));
  NAi21      u070(.An(i_6_), .B(i_11_), .Y(men_men_n93_));
  NO2        u071(.A(i_5_), .B(i_8_), .Y(men_men_n94_));
  NOi21      u072(.An(men_men_n94_), .B(men_men_n93_), .Y(men_men_n95_));
  NA2        u073(.A(men_men_n92_), .B(men_men_n32_), .Y(men_men_n96_));
  INV        u074(.A(i_7_), .Y(men_men_n97_));
  NO2        u075(.A(i_0_), .B(i_5_), .Y(men_men_n98_));
  NO2        u076(.A(men_men_n98_), .B(men_men_n81_), .Y(men_men_n99_));
  NA2        u077(.A(i_12_), .B(i_3_), .Y(men_men_n100_));
  NAi21      u078(.An(i_7_), .B(i_11_), .Y(men_men_n101_));
  NO3        u079(.A(men_men_n101_), .B(men_men_n86_), .C(men_men_n52_), .Y(men_men_n102_));
  AN2        u080(.A(i_2_), .B(i_10_), .Y(men_men_n103_));
  NO2        u081(.A(men_men_n103_), .B(i_7_), .Y(men_men_n104_));
  OR2        u082(.A(men_men_n76_), .B(men_men_n57_), .Y(men_men_n105_));
  NO2        u083(.A(i_8_), .B(men_men_n97_), .Y(men_men_n106_));
  NO3        u084(.A(men_men_n106_), .B(men_men_n105_), .C(men_men_n104_), .Y(men_men_n107_));
  NA2        u085(.A(i_12_), .B(i_7_), .Y(men_men_n108_));
  NA2        u086(.A(i_1_), .B(i_0_), .Y(men_men_n109_));
  NA2        u087(.A(i_11_), .B(i_12_), .Y(men_men_n110_));
  OAI210     u088(.A0(men_men_n109_), .A1(men_men_n108_), .B0(men_men_n110_), .Y(men_men_n111_));
  NO2        u089(.A(men_men_n111_), .B(men_men_n107_), .Y(men_men_n112_));
  NAi31      u090(.An(men_men_n102_), .B(men_men_n112_), .C(men_men_n96_), .Y(men_men_n113_));
  NOi21      u091(.An(i_1_), .B(i_5_), .Y(men_men_n114_));
  NA2        u092(.A(men_men_n114_), .B(i_11_), .Y(men_men_n115_));
  NA2        u093(.A(men_men_n97_), .B(men_men_n37_), .Y(men_men_n116_));
  NA2        u094(.A(i_7_), .B(men_men_n25_), .Y(men_men_n117_));
  NA2        u095(.A(men_men_n117_), .B(men_men_n116_), .Y(men_men_n118_));
  NO2        u096(.A(men_men_n118_), .B(men_men_n45_), .Y(men_men_n119_));
  NA2        u097(.A(men_men_n87_), .B(men_men_n86_), .Y(men_men_n120_));
  NAi21      u098(.An(i_3_), .B(i_8_), .Y(men_men_n121_));
  NA2        u099(.A(men_men_n121_), .B(men_men_n60_), .Y(men_men_n122_));
  NOi31      u100(.An(men_men_n122_), .B(men_men_n120_), .C(men_men_n119_), .Y(men_men_n123_));
  NO2        u101(.A(i_1_), .B(men_men_n81_), .Y(men_men_n124_));
  NO2        u102(.A(i_6_), .B(i_5_), .Y(men_men_n125_));
  NA2        u103(.A(men_men_n125_), .B(i_3_), .Y(men_men_n126_));
  AO210      u104(.A0(men_men_n126_), .A1(men_men_n46_), .B0(men_men_n124_), .Y(men_men_n127_));
  OAI220     u105(.A0(men_men_n127_), .A1(men_men_n101_), .B0(men_men_n123_), .B1(men_men_n115_), .Y(men_men_n128_));
  NO3        u106(.A(men_men_n128_), .B(men_men_n113_), .C(men_men_n91_), .Y(men_men_n129_));
  NA3        u107(.A(men_men_n129_), .B(men_men_n75_), .C(men_men_n55_), .Y(men2));
  NA3        u108(.A(men_men_n73_), .B(men_men_n65_), .C(men_men_n30_), .Y(men0));
  AN2        u109(.A(i_8_), .B(i_7_), .Y(men_men_n132_));
  NA2        u110(.A(men_men_n132_), .B(i_6_), .Y(men_men_n133_));
  NO2        u111(.A(i_12_), .B(i_13_), .Y(men_men_n134_));
  NAi21      u112(.An(i_5_), .B(i_11_), .Y(men_men_n135_));
  NOi21      u113(.An(men_men_n134_), .B(men_men_n135_), .Y(men_men_n136_));
  NO2        u114(.A(i_0_), .B(i_1_), .Y(men_men_n137_));
  NA2        u115(.A(i_2_), .B(i_3_), .Y(men_men_n138_));
  NO2        u116(.A(men_men_n138_), .B(i_4_), .Y(men_men_n139_));
  NA3        u117(.A(men_men_n139_), .B(men_men_n137_), .C(men_men_n136_), .Y(men_men_n140_));
  OR2        u118(.A(men_men_n140_), .B(men_men_n25_), .Y(men_men_n141_));
  AN2        u119(.A(men_men_n134_), .B(men_men_n78_), .Y(men_men_n142_));
  NO2        u120(.A(men_men_n142_), .B(men_men_n27_), .Y(men_men_n143_));
  NA2        u121(.A(i_1_), .B(i_5_), .Y(men_men_n144_));
  NO2        u122(.A(men_men_n69_), .B(men_men_n45_), .Y(men_men_n145_));
  NA2        u123(.A(men_men_n145_), .B(men_men_n36_), .Y(men_men_n146_));
  NO3        u124(.A(men_men_n146_), .B(men_men_n144_), .C(men_men_n143_), .Y(men_men_n147_));
  OR2        u125(.A(i_0_), .B(i_1_), .Y(men_men_n148_));
  NO3        u126(.A(men_men_n148_), .B(men_men_n76_), .C(i_13_), .Y(men_men_n149_));
  NAi32      u127(.An(i_2_), .Bn(i_3_), .C(i_4_), .Y(men_men_n150_));
  NAi21      u128(.An(men_men_n150_), .B(men_men_n149_), .Y(men_men_n151_));
  NOi21      u129(.An(i_4_), .B(i_10_), .Y(men_men_n152_));
  NA2        u130(.A(men_men_n152_), .B(men_men_n39_), .Y(men_men_n153_));
  NO2        u131(.A(i_3_), .B(i_5_), .Y(men_men_n154_));
  NO3        u132(.A(men_men_n69_), .B(i_2_), .C(i_1_), .Y(men_men_n155_));
  NA2        u133(.A(men_men_n155_), .B(men_men_n154_), .Y(men_men_n156_));
  OAI210     u134(.A0(men_men_n156_), .A1(men_men_n153_), .B0(men_men_n151_), .Y(men_men_n157_));
  NO2        u135(.A(men_men_n157_), .B(men_men_n147_), .Y(men_men_n158_));
  AOI210     u136(.A0(men_men_n158_), .A1(men_men_n141_), .B0(men_men_n133_), .Y(men_men_n159_));
  NA2        u137(.A(i_3_), .B(men_men_n47_), .Y(men_men_n160_));
  NOi21      u138(.An(i_4_), .B(i_9_), .Y(men_men_n161_));
  NOi21      u139(.An(i_11_), .B(i_13_), .Y(men_men_n162_));
  NA2        u140(.A(men_men_n162_), .B(men_men_n161_), .Y(men_men_n163_));
  OR2        u141(.A(men_men_n163_), .B(men_men_n160_), .Y(men_men_n164_));
  NO2        u142(.A(i_4_), .B(i_5_), .Y(men_men_n165_));
  NAi21      u143(.An(i_12_), .B(i_11_), .Y(men_men_n166_));
  NO2        u144(.A(men_men_n166_), .B(i_13_), .Y(men_men_n167_));
  NA3        u145(.A(men_men_n167_), .B(men_men_n165_), .C(men_men_n78_), .Y(men_men_n168_));
  AOI210     u146(.A0(men_men_n168_), .A1(men_men_n164_), .B0(men_men_n1011_), .Y(men_men_n169_));
  NO2        u147(.A(men_men_n69_), .B(men_men_n61_), .Y(men_men_n170_));
  NA2        u148(.A(men_men_n170_), .B(men_men_n45_), .Y(men_men_n171_));
  NA2        u149(.A(men_men_n36_), .B(i_5_), .Y(men_men_n172_));
  NAi31      u150(.An(men_men_n172_), .B(men_men_n142_), .C(i_11_), .Y(men_men_n173_));
  NA2        u151(.A(i_3_), .B(i_5_), .Y(men_men_n174_));
  OR2        u152(.A(men_men_n174_), .B(men_men_n163_), .Y(men_men_n175_));
  AOI210     u153(.A0(men_men_n175_), .A1(men_men_n173_), .B0(men_men_n171_), .Y(men_men_n176_));
  NO2        u154(.A(men_men_n69_), .B(i_5_), .Y(men_men_n177_));
  NO2        u155(.A(i_13_), .B(i_10_), .Y(men_men_n178_));
  NA3        u156(.A(men_men_n178_), .B(men_men_n177_), .C(men_men_n43_), .Y(men_men_n179_));
  NO2        u157(.A(i_2_), .B(i_1_), .Y(men_men_n180_));
  NA2        u158(.A(men_men_n180_), .B(i_3_), .Y(men_men_n181_));
  NAi21      u159(.An(i_4_), .B(i_12_), .Y(men_men_n182_));
  NO4        u160(.A(men_men_n182_), .B(men_men_n181_), .C(men_men_n179_), .D(men_men_n25_), .Y(men_men_n183_));
  NO3        u161(.A(men_men_n183_), .B(men_men_n176_), .C(men_men_n169_), .Y(men_men_n184_));
  INV        u162(.A(i_8_), .Y(men_men_n185_));
  NO2        u163(.A(men_men_n185_), .B(i_7_), .Y(men_men_n186_));
  NA2        u164(.A(men_men_n186_), .B(i_6_), .Y(men_men_n187_));
  NO3        u165(.A(i_3_), .B(men_men_n81_), .C(men_men_n47_), .Y(men_men_n188_));
  NA2        u166(.A(men_men_n188_), .B(men_men_n106_), .Y(men_men_n189_));
  NO3        u167(.A(i_0_), .B(i_2_), .C(i_1_), .Y(men_men_n190_));
  NA3        u168(.A(men_men_n190_), .B(men_men_n39_), .C(men_men_n43_), .Y(men_men_n191_));
  NO3        u169(.A(i_11_), .B(i_13_), .C(i_9_), .Y(men_men_n192_));
  NA2        u170(.A(i_12_), .B(men_men_n192_), .Y(men_men_n193_));
  AOI210     u171(.A0(men_men_n193_), .A1(men_men_n191_), .B0(men_men_n189_), .Y(men_men_n194_));
  NO2        u172(.A(i_3_), .B(i_8_), .Y(men_men_n195_));
  NO3        u173(.A(i_11_), .B(i_10_), .C(i_9_), .Y(men_men_n196_));
  NA3        u174(.A(men_men_n196_), .B(men_men_n195_), .C(men_men_n39_), .Y(men_men_n197_));
  NO2        u175(.A(men_men_n98_), .B(men_men_n57_), .Y(men_men_n198_));
  NO2        u176(.A(i_13_), .B(i_9_), .Y(men_men_n199_));
  NA3        u177(.A(men_men_n199_), .B(i_6_), .C(men_men_n185_), .Y(men_men_n200_));
  NAi21      u178(.An(i_12_), .B(i_3_), .Y(men_men_n201_));
  OR2        u179(.A(men_men_n201_), .B(men_men_n200_), .Y(men_men_n202_));
  NO2        u180(.A(men_men_n43_), .B(i_5_), .Y(men_men_n203_));
  NO3        u181(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n204_));
  OAI220     u182(.A0(i_2_), .A1(men_men_n202_), .B0(men_men_n98_), .B1(men_men_n197_), .Y(men_men_n205_));
  AOI210     u183(.A0(men_men_n205_), .A1(i_7_), .B0(men_men_n194_), .Y(men_men_n206_));
  OAI220     u184(.A0(men_men_n206_), .A1(i_4_), .B0(men_men_n187_), .B1(men_men_n184_), .Y(men_men_n207_));
  NAi21      u185(.An(i_12_), .B(i_7_), .Y(men_men_n208_));
  NA3        u186(.A(i_13_), .B(men_men_n185_), .C(i_10_), .Y(men_men_n209_));
  NO2        u187(.A(men_men_n209_), .B(men_men_n208_), .Y(men_men_n210_));
  NA2        u188(.A(i_0_), .B(i_5_), .Y(men_men_n211_));
  NA2        u189(.A(men_men_n211_), .B(men_men_n99_), .Y(men_men_n212_));
  OAI220     u190(.A0(men_men_n212_), .A1(men_men_n181_), .B0(men_men_n171_), .B1(men_men_n126_), .Y(men_men_n213_));
  NAi31      u191(.An(i_9_), .B(i_6_), .C(i_5_), .Y(men_men_n214_));
  NO2        u192(.A(men_men_n36_), .B(i_13_), .Y(men_men_n215_));
  NO2        u193(.A(men_men_n69_), .B(men_men_n26_), .Y(men_men_n216_));
  NO2        u194(.A(men_men_n45_), .B(men_men_n61_), .Y(men_men_n217_));
  NA3        u195(.A(men_men_n217_), .B(men_men_n216_), .C(men_men_n215_), .Y(men_men_n218_));
  INV        u196(.A(i_13_), .Y(men_men_n219_));
  NO2        u197(.A(i_12_), .B(men_men_n219_), .Y(men_men_n220_));
  NA3        u198(.A(men_men_n220_), .B(men_men_n190_), .C(men_men_n188_), .Y(men_men_n221_));
  NA2        u199(.A(men_men_n218_), .B(men_men_n221_), .Y(men_men_n222_));
  AOI220     u200(.A0(men_men_n222_), .A1(men_men_n132_), .B0(men_men_n213_), .B1(men_men_n210_), .Y(men_men_n223_));
  NO2        u201(.A(i_12_), .B(men_men_n37_), .Y(men_men_n224_));
  NO2        u202(.A(men_men_n174_), .B(i_4_), .Y(men_men_n225_));
  INV        u203(.A(men_men_n225_), .Y(men_men_n226_));
  OR2        u204(.A(i_8_), .B(i_7_), .Y(men_men_n227_));
  NO2        u205(.A(men_men_n227_), .B(men_men_n81_), .Y(men_men_n228_));
  NO2        u206(.A(men_men_n52_), .B(i_1_), .Y(men_men_n229_));
  NA2        u207(.A(men_men_n229_), .B(men_men_n228_), .Y(men_men_n230_));
  INV        u208(.A(i_12_), .Y(men_men_n231_));
  NO3        u209(.A(men_men_n36_), .B(i_8_), .C(i_10_), .Y(men_men_n232_));
  NA2        u210(.A(i_2_), .B(i_1_), .Y(men_men_n233_));
  NO2        u211(.A(men_men_n230_), .B(men_men_n226_), .Y(men_men_n234_));
  NAi21      u212(.An(i_4_), .B(i_3_), .Y(men_men_n235_));
  NO2        u213(.A(men_men_n235_), .B(men_men_n71_), .Y(men_men_n236_));
  NO2        u214(.A(i_0_), .B(i_6_), .Y(men_men_n237_));
  NOi41      u215(.An(i_4_), .B(i_8_), .C(i_7_), .D(i_10_), .Y(men_men_n238_));
  NA2        u216(.A(men_men_n238_), .B(men_men_n237_), .Y(men_men_n239_));
  NO2        u217(.A(men_men_n233_), .B(men_men_n174_), .Y(men_men_n240_));
  NAi21      u218(.An(men_men_n239_), .B(men_men_n240_), .Y(men_men_n241_));
  INV        u219(.A(men_men_n241_), .Y(men_men_n242_));
  AOI220     u220(.A0(men_men_n242_), .A1(men_men_n39_), .B0(men_men_n234_), .B1(men_men_n199_), .Y(men_men_n243_));
  NO2        u221(.A(i_11_), .B(men_men_n219_), .Y(men_men_n244_));
  NOi21      u222(.An(i_1_), .B(i_6_), .Y(men_men_n245_));
  NA2        u223(.A(men_men_n231_), .B(i_9_), .Y(men_men_n246_));
  OR4        u224(.A(men_men_n246_), .B(i_3_), .C(men_men_n245_), .D(men_men_n177_), .Y(men_men_n247_));
  NO2        u225(.A(men_men_n47_), .B(men_men_n25_), .Y(men_men_n248_));
  NO2        u226(.A(i_12_), .B(i_3_), .Y(men_men_n249_));
  NA2        u227(.A(men_men_n69_), .B(i_5_), .Y(men_men_n250_));
  NA2        u228(.A(i_3_), .B(i_9_), .Y(men_men_n251_));
  NAi21      u229(.An(i_7_), .B(i_10_), .Y(men_men_n252_));
  NO2        u230(.A(men_men_n252_), .B(men_men_n251_), .Y(men_men_n253_));
  NA3        u231(.A(men_men_n253_), .B(men_men_n250_), .C(men_men_n62_), .Y(men_men_n254_));
  NA2        u232(.A(men_men_n254_), .B(men_men_n247_), .Y(men_men_n255_));
  NA3        u233(.A(i_1_), .B(i_8_), .C(i_7_), .Y(men_men_n256_));
  NA2        u234(.A(men_men_n255_), .B(men_men_n244_), .Y(men_men_n257_));
  NO2        u235(.A(men_men_n227_), .B(men_men_n37_), .Y(men_men_n258_));
  NA2        u236(.A(i_12_), .B(i_6_), .Y(men_men_n259_));
  OR2        u237(.A(i_13_), .B(i_9_), .Y(men_men_n260_));
  NO3        u238(.A(men_men_n260_), .B(men_men_n259_), .C(men_men_n47_), .Y(men_men_n261_));
  NO2        u239(.A(men_men_n235_), .B(i_2_), .Y(men_men_n262_));
  NA3        u240(.A(men_men_n262_), .B(men_men_n261_), .C(men_men_n43_), .Y(men_men_n263_));
  NA2        u241(.A(men_men_n244_), .B(i_9_), .Y(men_men_n264_));
  OAI210     u242(.A0(men_men_n69_), .A1(men_men_n264_), .B0(men_men_n263_), .Y(men_men_n265_));
  NA2        u243(.A(men_men_n145_), .B(men_men_n61_), .Y(men_men_n266_));
  NO3        u244(.A(i_11_), .B(men_men_n219_), .C(men_men_n25_), .Y(men_men_n267_));
  NO2        u245(.A(i_3_), .B(i_8_), .Y(men_men_n268_));
  NO2        u246(.A(i_6_), .B(men_men_n47_), .Y(men_men_n269_));
  NA3        u247(.A(men_men_n269_), .B(men_men_n268_), .C(men_men_n267_), .Y(men_men_n270_));
  NO3        u248(.A(men_men_n26_), .B(men_men_n81_), .C(i_5_), .Y(men_men_n271_));
  NA3        u249(.A(men_men_n271_), .B(men_men_n258_), .C(men_men_n220_), .Y(men_men_n272_));
  AOI210     u250(.A0(men_men_n272_), .A1(men_men_n270_), .B0(men_men_n266_), .Y(men_men_n273_));
  AOI210     u251(.A0(men_men_n265_), .A1(men_men_n258_), .B0(men_men_n273_), .Y(men_men_n274_));
  NA4        u252(.A(men_men_n274_), .B(men_men_n257_), .C(men_men_n243_), .D(men_men_n223_), .Y(men_men_n275_));
  NO3        u253(.A(i_12_), .B(men_men_n219_), .C(men_men_n37_), .Y(men_men_n276_));
  INV        u254(.A(men_men_n276_), .Y(men_men_n277_));
  NOi21      u255(.An(men_men_n154_), .B(men_men_n81_), .Y(men_men_n278_));
  NO3        u256(.A(i_0_), .B(men_men_n45_), .C(i_1_), .Y(men_men_n279_));
  AOI220     u257(.A0(men_men_n279_), .A1(men_men_n188_), .B0(men_men_n278_), .B1(men_men_n229_), .Y(men_men_n280_));
  NO2        u258(.A(men_men_n280_), .B(i_7_), .Y(men_men_n281_));
  NO3        u259(.A(i_0_), .B(i_2_), .C(men_men_n61_), .Y(men_men_n282_));
  NO2        u260(.A(men_men_n233_), .B(i_0_), .Y(men_men_n283_));
  AOI220     u261(.A0(men_men_n283_), .A1(men_men_n186_), .B0(men_men_n282_), .B1(men_men_n132_), .Y(men_men_n284_));
  NA2        u262(.A(men_men_n269_), .B(men_men_n26_), .Y(men_men_n285_));
  NO2        u263(.A(men_men_n285_), .B(men_men_n284_), .Y(men_men_n286_));
  NA2        u264(.A(i_0_), .B(i_1_), .Y(men_men_n287_));
  NO2        u265(.A(men_men_n287_), .B(i_2_), .Y(men_men_n288_));
  NO2        u266(.A(men_men_n58_), .B(i_6_), .Y(men_men_n289_));
  NA3        u267(.A(men_men_n289_), .B(men_men_n288_), .C(men_men_n154_), .Y(men_men_n290_));
  OAI210     u268(.A0(men_men_n156_), .A1(men_men_n133_), .B0(men_men_n290_), .Y(men_men_n291_));
  NO3        u269(.A(men_men_n291_), .B(men_men_n286_), .C(men_men_n281_), .Y(men_men_n292_));
  NO2        u270(.A(i_3_), .B(i_10_), .Y(men_men_n293_));
  NA3        u271(.A(men_men_n293_), .B(men_men_n39_), .C(men_men_n43_), .Y(men_men_n294_));
  NO2        u272(.A(i_2_), .B(men_men_n97_), .Y(men_men_n295_));
  NOi21      u273(.An(men_men_n211_), .B(men_men_n98_), .Y(men_men_n296_));
  NA3        u274(.A(men_men_n296_), .B(i_1_), .C(men_men_n295_), .Y(men_men_n297_));
  AN2        u275(.A(i_3_), .B(i_10_), .Y(men_men_n298_));
  NA3        u276(.A(men_men_n190_), .B(men_men_n167_), .C(men_men_n165_), .Y(men_men_n299_));
  NO2        u277(.A(i_5_), .B(men_men_n37_), .Y(men_men_n300_));
  NO2        u278(.A(men_men_n45_), .B(men_men_n26_), .Y(men_men_n301_));
  OR2        u279(.A(men_men_n297_), .B(men_men_n294_), .Y(men_men_n302_));
  OAI220     u280(.A0(men_men_n302_), .A1(i_6_), .B0(men_men_n292_), .B1(men_men_n277_), .Y(men_men_n303_));
  NO4        u281(.A(men_men_n303_), .B(men_men_n275_), .C(men_men_n207_), .D(men_men_n159_), .Y(men_men_n304_));
  NO3        u282(.A(men_men_n43_), .B(i_13_), .C(i_9_), .Y(men_men_n305_));
  NO3        u283(.A(i_6_), .B(men_men_n185_), .C(i_7_), .Y(men_men_n306_));
  NA2        u284(.A(men_men_n306_), .B(men_men_n190_), .Y(men_men_n307_));
  AOI210     u285(.A0(men_men_n307_), .A1(men_men_n233_), .B0(men_men_n160_), .Y(men_men_n308_));
  NO2        u286(.A(i_2_), .B(i_3_), .Y(men_men_n309_));
  OR2        u287(.A(i_0_), .B(i_5_), .Y(men_men_n310_));
  NA2        u288(.A(men_men_n211_), .B(men_men_n310_), .Y(men_men_n311_));
  NA4        u289(.A(men_men_n311_), .B(men_men_n228_), .C(men_men_n309_), .D(i_1_), .Y(men_men_n312_));
  NA3        u290(.A(men_men_n283_), .B(men_men_n278_), .C(men_men_n106_), .Y(men_men_n313_));
  NO2        u291(.A(i_8_), .B(i_6_), .Y(men_men_n314_));
  NO2        u292(.A(men_men_n148_), .B(men_men_n45_), .Y(men_men_n315_));
  NA3        u293(.A(men_men_n315_), .B(men_men_n314_), .C(men_men_n154_), .Y(men_men_n316_));
  NA3        u294(.A(men_men_n316_), .B(men_men_n313_), .C(men_men_n312_), .Y(men_men_n317_));
  OAI210     u295(.A0(men_men_n317_), .A1(men_men_n308_), .B0(i_4_), .Y(men_men_n318_));
  NO2        u296(.A(i_12_), .B(i_10_), .Y(men_men_n319_));
  NOi21      u297(.An(i_5_), .B(i_0_), .Y(men_men_n320_));
  AOI210     u298(.A0(i_2_), .A1(men_men_n47_), .B0(men_men_n97_), .Y(men_men_n321_));
  NO4        u299(.A(men_men_n321_), .B(i_4_), .C(men_men_n320_), .D(men_men_n121_), .Y(men_men_n322_));
  NA4        u300(.A(men_men_n79_), .B(men_men_n36_), .C(men_men_n81_), .D(i_8_), .Y(men_men_n323_));
  NA2        u301(.A(men_men_n322_), .B(men_men_n319_), .Y(men_men_n324_));
  NO2        u302(.A(i_6_), .B(i_8_), .Y(men_men_n325_));
  AN2        u303(.A(i_0_), .B(men_men_n325_), .Y(men_men_n326_));
  NO2        u304(.A(i_1_), .B(i_7_), .Y(men_men_n327_));
  NA3        u305(.A(men_men_n326_), .B(i_4_), .C(i_5_), .Y(men_men_n328_));
  NA3        u306(.A(men_men_n328_), .B(men_men_n324_), .C(men_men_n318_), .Y(men_men_n329_));
  NA2        u307(.A(men_men_n1016_), .B(i_6_), .Y(men_men_n330_));
  NA3        u308(.A(men_men_n245_), .B(men_men_n295_), .C(men_men_n185_), .Y(men_men_n331_));
  AOI210     u309(.A0(men_men_n331_), .A1(men_men_n330_), .B0(men_men_n311_), .Y(men_men_n332_));
  NOi21      u310(.An(men_men_n144_), .B(men_men_n99_), .Y(men_men_n333_));
  NO2        u311(.A(men_men_n333_), .B(men_men_n117_), .Y(men_men_n334_));
  OAI210     u312(.A0(men_men_n334_), .A1(men_men_n332_), .B0(i_3_), .Y(men_men_n335_));
  NO2        u313(.A(men_men_n287_), .B(men_men_n77_), .Y(men_men_n336_));
  NA2        u314(.A(men_men_n336_), .B(men_men_n125_), .Y(men_men_n337_));
  NO2        u315(.A(men_men_n88_), .B(men_men_n185_), .Y(men_men_n338_));
  NA3        u316(.A(men_men_n296_), .B(men_men_n338_), .C(men_men_n61_), .Y(men_men_n339_));
  AOI210     u317(.A0(men_men_n339_), .A1(men_men_n337_), .B0(i_3_), .Y(men_men_n340_));
  NO2        u318(.A(men_men_n185_), .B(i_9_), .Y(men_men_n341_));
  NA2        u319(.A(men_men_n341_), .B(men_men_n198_), .Y(men_men_n342_));
  NO2        u320(.A(men_men_n340_), .B(men_men_n286_), .Y(men_men_n343_));
  AOI210     u321(.A0(men_men_n343_), .A1(men_men_n335_), .B0(men_men_n153_), .Y(men_men_n344_));
  AOI210     u322(.A0(men_men_n329_), .A1(men_men_n305_), .B0(men_men_n344_), .Y(men_men_n345_));
  NOi32      u323(.An(i_11_), .Bn(i_12_), .C(i_13_), .Y(men_men_n346_));
  INV        u324(.A(men_men_n346_), .Y(men_men_n347_));
  NAi21      u325(.An(i_1_), .B(i_5_), .Y(men_men_n348_));
  NA2        u326(.A(men_men_n348_), .B(i_0_), .Y(men_men_n349_));
  NA2        u327(.A(men_men_n349_), .B(men_men_n25_), .Y(men_men_n350_));
  OAI210     u328(.A0(men_men_n350_), .A1(men_men_n150_), .B0(men_men_n239_), .Y(men_men_n351_));
  NAi41      u329(.An(i_9_), .B(i_4_), .C(i_8_), .D(i_7_), .Y(men_men_n352_));
  OAI220     u330(.A0(men_men_n352_), .A1(men_men_n348_), .B0(men_men_n214_), .B1(men_men_n150_), .Y(men_men_n353_));
  NO2        u331(.A(men_men_n150_), .B(men_men_n148_), .Y(men_men_n354_));
  NOi32      u332(.An(i_4_), .Bn(i_8_), .C(i_9_), .Y(men_men_n355_));
  NAi21      u333(.An(i_6_), .B(i_1_), .Y(men_men_n356_));
  NA2        u334(.A(men_men_n355_), .B(men_men_n45_), .Y(men_men_n357_));
  NO2        u335(.A(men_men_n357_), .B(i_0_), .Y(men_men_n358_));
  OR3        u336(.A(men_men_n358_), .B(men_men_n354_), .C(men_men_n353_), .Y(men_men_n359_));
  NO2        u337(.A(i_1_), .B(men_men_n97_), .Y(men_men_n360_));
  NAi21      u338(.An(i_3_), .B(i_4_), .Y(men_men_n361_));
  NO2        u339(.A(men_men_n361_), .B(i_9_), .Y(men_men_n362_));
  AN2        u340(.A(i_6_), .B(i_7_), .Y(men_men_n363_));
  OAI210     u341(.A0(men_men_n363_), .A1(men_men_n360_), .B0(men_men_n362_), .Y(men_men_n364_));
  NA2        u342(.A(i_2_), .B(i_7_), .Y(men_men_n365_));
  NO2        u343(.A(men_men_n361_), .B(i_10_), .Y(men_men_n366_));
  NA3        u344(.A(men_men_n366_), .B(men_men_n365_), .C(men_men_n237_), .Y(men_men_n367_));
  AOI210     u345(.A0(men_men_n367_), .A1(men_men_n364_), .B0(men_men_n177_), .Y(men_men_n368_));
  AOI210     u346(.A0(i_2_), .A1(i_7_), .B0(i_6_), .Y(men_men_n369_));
  OAI210     u347(.A0(men_men_n369_), .A1(men_men_n180_), .B0(men_men_n366_), .Y(men_men_n370_));
  AOI220     u348(.A0(men_men_n366_), .A1(men_men_n327_), .B0(men_men_n232_), .B1(men_men_n180_), .Y(men_men_n371_));
  NO2        u349(.A(men_men_n370_), .B(i_5_), .Y(men_men_n372_));
  NO4        u350(.A(men_men_n372_), .B(men_men_n368_), .C(men_men_n359_), .D(men_men_n351_), .Y(men_men_n373_));
  NO2        u351(.A(men_men_n373_), .B(men_men_n347_), .Y(men_men_n374_));
  NO2        u352(.A(men_men_n58_), .B(men_men_n25_), .Y(men_men_n375_));
  AN2        u353(.A(i_12_), .B(i_5_), .Y(men_men_n376_));
  NO2        u354(.A(i_4_), .B(men_men_n26_), .Y(men_men_n377_));
  NA2        u355(.A(men_men_n377_), .B(men_men_n376_), .Y(men_men_n378_));
  NO2        u356(.A(i_11_), .B(i_6_), .Y(men_men_n379_));
  NA3        u357(.A(men_men_n379_), .B(men_men_n315_), .C(men_men_n219_), .Y(men_men_n380_));
  NO2        u358(.A(men_men_n380_), .B(men_men_n378_), .Y(men_men_n381_));
  NO2        u359(.A(men_men_n235_), .B(i_5_), .Y(men_men_n382_));
  NO2        u360(.A(i_5_), .B(i_10_), .Y(men_men_n383_));
  AOI220     u361(.A0(men_men_n383_), .A1(men_men_n262_), .B0(men_men_n382_), .B1(men_men_n190_), .Y(men_men_n384_));
  INV        u362(.A(men_men_n44_), .Y(men_men_n385_));
  NO2        u363(.A(men_men_n385_), .B(men_men_n384_), .Y(men_men_n386_));
  OAI210     u364(.A0(men_men_n386_), .A1(men_men_n381_), .B0(men_men_n375_), .Y(men_men_n387_));
  NO2        u365(.A(men_men_n37_), .B(men_men_n25_), .Y(men_men_n388_));
  NO2        u366(.A(men_men_n140_), .B(men_men_n81_), .Y(men_men_n389_));
  OAI210     u367(.A0(men_men_n389_), .A1(men_men_n381_), .B0(men_men_n388_), .Y(men_men_n390_));
  NO3        u368(.A(men_men_n81_), .B(men_men_n47_), .C(i_9_), .Y(men_men_n391_));
  NO2        u369(.A(i_11_), .B(i_12_), .Y(men_men_n392_));
  NA2        u370(.A(men_men_n392_), .B(men_men_n36_), .Y(men_men_n393_));
  NO2        u371(.A(i_3_), .B(men_men_n393_), .Y(men_men_n394_));
  NA2        u372(.A(men_men_n383_), .B(men_men_n231_), .Y(men_men_n395_));
  NA3        u373(.A(men_men_n106_), .B(i_4_), .C(i_11_), .Y(men_men_n396_));
  INV        u374(.A(men_men_n396_), .Y(men_men_n397_));
  NAi21      u375(.An(i_13_), .B(i_0_), .Y(men_men_n398_));
  NO2        u376(.A(men_men_n398_), .B(men_men_n233_), .Y(men_men_n399_));
  OAI210     u377(.A0(men_men_n397_), .A1(men_men_n394_), .B0(men_men_n399_), .Y(men_men_n400_));
  NA3        u378(.A(men_men_n400_), .B(men_men_n390_), .C(men_men_n387_), .Y(men_men_n401_));
  NA2        u379(.A(men_men_n43_), .B(men_men_n219_), .Y(men_men_n402_));
  NO3        u380(.A(i_1_), .B(i_12_), .C(men_men_n81_), .Y(men_men_n403_));
  NO2        u381(.A(i_0_), .B(i_11_), .Y(men_men_n404_));
  AN2        u382(.A(i_1_), .B(i_6_), .Y(men_men_n405_));
  NOi21      u383(.An(i_2_), .B(i_12_), .Y(men_men_n406_));
  NA2        u384(.A(men_men_n406_), .B(men_men_n405_), .Y(men_men_n407_));
  NO2        u385(.A(men_men_n407_), .B(men_men_n1010_), .Y(men_men_n408_));
  NA2        u386(.A(men_men_n132_), .B(i_9_), .Y(men_men_n409_));
  NA2        u387(.A(men_men_n408_), .B(i_9_), .Y(men_men_n410_));
  NAi21      u388(.An(i_9_), .B(i_4_), .Y(men_men_n411_));
  OR2        u389(.A(i_13_), .B(i_10_), .Y(men_men_n412_));
  NO3        u390(.A(men_men_n412_), .B(men_men_n110_), .C(men_men_n411_), .Y(men_men_n413_));
  NO2        u391(.A(men_men_n163_), .B(men_men_n116_), .Y(men_men_n414_));
  NO2        u392(.A(men_men_n97_), .B(men_men_n25_), .Y(men_men_n415_));
  NA2        u393(.A(men_men_n276_), .B(men_men_n415_), .Y(men_men_n416_));
  NA2        u394(.A(men_men_n269_), .B(men_men_n204_), .Y(men_men_n417_));
  OAI220     u395(.A0(men_men_n417_), .A1(men_men_n209_), .B0(men_men_n416_), .B1(men_men_n333_), .Y(men_men_n418_));
  INV        u396(.A(men_men_n418_), .Y(men_men_n419_));
  AOI210     u397(.A0(men_men_n419_), .A1(men_men_n410_), .B0(men_men_n26_), .Y(men_men_n420_));
  NA2        u398(.A(men_men_n313_), .B(men_men_n312_), .Y(men_men_n421_));
  AOI220     u399(.A0(men_men_n289_), .A1(men_men_n279_), .B0(men_men_n283_), .B1(i_7_), .Y(men_men_n422_));
  NO2        u400(.A(men_men_n174_), .B(men_men_n81_), .Y(men_men_n423_));
  AOI220     u401(.A0(men_men_n423_), .A1(men_men_n288_), .B0(men_men_n271_), .B1(men_men_n204_), .Y(men_men_n424_));
  NO2        u402(.A(men_men_n424_), .B(i_7_), .Y(men_men_n425_));
  NO2        u403(.A(men_men_n425_), .B(men_men_n421_), .Y(men_men_n426_));
  NA2        u404(.A(men_men_n188_), .B(men_men_n92_), .Y(men_men_n427_));
  NA3        u405(.A(men_men_n315_), .B(men_men_n154_), .C(men_men_n81_), .Y(men_men_n428_));
  AOI210     u406(.A0(men_men_n428_), .A1(men_men_n427_), .B0(i_8_), .Y(men_men_n429_));
  NA2        u407(.A(men_men_n185_), .B(i_10_), .Y(men_men_n430_));
  NA3        u408(.A(men_men_n250_), .B(men_men_n62_), .C(i_2_), .Y(men_men_n431_));
  NA2        u409(.A(men_men_n289_), .B(men_men_n229_), .Y(men_men_n432_));
  OAI220     u410(.A0(men_men_n432_), .A1(men_men_n174_), .B0(men_men_n431_), .B1(men_men_n430_), .Y(men_men_n433_));
  NO2        u411(.A(i_3_), .B(men_men_n47_), .Y(men_men_n434_));
  NA3        u412(.A(men_men_n327_), .B(men_men_n326_), .C(men_men_n434_), .Y(men_men_n435_));
  NA2        u413(.A(men_men_n306_), .B(men_men_n311_), .Y(men_men_n436_));
  OAI210     u414(.A0(men_men_n436_), .A1(men_men_n181_), .B0(men_men_n435_), .Y(men_men_n437_));
  NO3        u415(.A(men_men_n437_), .B(men_men_n433_), .C(men_men_n429_), .Y(men_men_n438_));
  AOI210     u416(.A0(men_men_n438_), .A1(men_men_n426_), .B0(men_men_n264_), .Y(men_men_n439_));
  NO4        u417(.A(men_men_n439_), .B(men_men_n420_), .C(men_men_n401_), .D(men_men_n374_), .Y(men_men_n440_));
  NO2        u418(.A(men_men_n69_), .B(i_13_), .Y(men_men_n441_));
  NO2        u419(.A(i_10_), .B(i_9_), .Y(men_men_n442_));
  NAi21      u420(.An(i_12_), .B(i_8_), .Y(men_men_n443_));
  NO2        u421(.A(men_men_n443_), .B(i_3_), .Y(men_men_n444_));
  NA2        u422(.A(i_2_), .B(men_men_n99_), .Y(men_men_n445_));
  NO2        u423(.A(men_men_n445_), .B(men_men_n197_), .Y(men_men_n446_));
  NA2        u424(.A(men_men_n301_), .B(i_0_), .Y(men_men_n447_));
  NO3        u425(.A(men_men_n23_), .B(i_10_), .C(i_9_), .Y(men_men_n448_));
  NA2        u426(.A(men_men_n259_), .B(men_men_n93_), .Y(men_men_n449_));
  NA2        u427(.A(men_men_n449_), .B(men_men_n448_), .Y(men_men_n450_));
  NA2        u428(.A(i_8_), .B(i_9_), .Y(men_men_n451_));
  NA2        u429(.A(men_men_n276_), .B(men_men_n198_), .Y(men_men_n452_));
  OAI220     u430(.A0(men_men_n452_), .A1(men_men_n451_), .B0(men_men_n450_), .B1(men_men_n447_), .Y(men_men_n453_));
  NA2        u431(.A(men_men_n244_), .B(men_men_n300_), .Y(men_men_n454_));
  NO3        u432(.A(i_6_), .B(i_8_), .C(i_7_), .Y(men_men_n455_));
  INV        u433(.A(men_men_n455_), .Y(men_men_n456_));
  NA3        u434(.A(i_2_), .B(i_10_), .C(i_9_), .Y(men_men_n457_));
  NO2        u435(.A(men_men_n456_), .B(men_men_n454_), .Y(men_men_n458_));
  NO3        u436(.A(men_men_n458_), .B(men_men_n453_), .C(men_men_n446_), .Y(men_men_n459_));
  NA2        u437(.A(men_men_n288_), .B(men_men_n101_), .Y(men_men_n460_));
  OR2        u438(.A(men_men_n460_), .B(men_men_n200_), .Y(men_men_n461_));
  OA220      u439(.A0(men_men_n342_), .A1(men_men_n153_), .B0(men_men_n461_), .B1(men_men_n226_), .Y(men_men_n462_));
  NA2        u440(.A(men_men_n92_), .B(i_13_), .Y(men_men_n463_));
  NA2        u441(.A(men_men_n423_), .B(men_men_n375_), .Y(men_men_n464_));
  NO2        u442(.A(i_2_), .B(i_13_), .Y(men_men_n465_));
  NA3        u443(.A(men_men_n465_), .B(men_men_n152_), .C(men_men_n95_), .Y(men_men_n466_));
  OAI220     u444(.A0(men_men_n466_), .A1(men_men_n231_), .B0(men_men_n464_), .B1(men_men_n463_), .Y(men_men_n467_));
  NO3        u445(.A(i_4_), .B(men_men_n47_), .C(i_8_), .Y(men_men_n468_));
  NO2        u446(.A(i_6_), .B(i_7_), .Y(men_men_n469_));
  NO2        u447(.A(men_men_n69_), .B(i_3_), .Y(men_men_n470_));
  NOi21      u448(.An(i_2_), .B(i_7_), .Y(men_men_n471_));
  NAi31      u449(.An(i_11_), .B(men_men_n471_), .C(men_men_n470_), .Y(men_men_n472_));
  NO2        u450(.A(men_men_n412_), .B(i_6_), .Y(men_men_n473_));
  NA3        u451(.A(men_men_n473_), .B(i_1_), .C(men_men_n71_), .Y(men_men_n474_));
  NO2        u452(.A(men_men_n474_), .B(men_men_n472_), .Y(men_men_n475_));
  NO2        u453(.A(i_3_), .B(men_men_n185_), .Y(men_men_n476_));
  NO2        u454(.A(i_6_), .B(i_10_), .Y(men_men_n477_));
  NA4        u455(.A(men_men_n477_), .B(men_men_n305_), .C(men_men_n476_), .D(men_men_n231_), .Y(men_men_n478_));
  NO2        u456(.A(men_men_n478_), .B(men_men_n146_), .Y(men_men_n479_));
  NA3        u457(.A(men_men_n238_), .B(men_men_n162_), .C(men_men_n125_), .Y(men_men_n480_));
  NA2        u458(.A(men_men_n45_), .B(men_men_n43_), .Y(men_men_n481_));
  NO2        u459(.A(men_men_n148_), .B(i_3_), .Y(men_men_n482_));
  NAi31      u460(.An(men_men_n481_), .B(men_men_n482_), .C(men_men_n220_), .Y(men_men_n483_));
  NA3        u461(.A(men_men_n388_), .B(men_men_n170_), .C(men_men_n139_), .Y(men_men_n484_));
  NA3        u462(.A(men_men_n484_), .B(men_men_n483_), .C(men_men_n480_), .Y(men_men_n485_));
  NO4        u463(.A(men_men_n485_), .B(men_men_n479_), .C(men_men_n475_), .D(men_men_n467_), .Y(men_men_n486_));
  NA2        u464(.A(men_men_n448_), .B(men_men_n376_), .Y(men_men_n487_));
  NA2        u465(.A(men_men_n455_), .B(men_men_n383_), .Y(men_men_n488_));
  NO2        u466(.A(men_men_n488_), .B(men_men_n218_), .Y(men_men_n489_));
  NAi21      u467(.An(men_men_n209_), .B(men_men_n392_), .Y(men_men_n490_));
  NA2        u468(.A(men_men_n327_), .B(men_men_n211_), .Y(men_men_n491_));
  NO2        u469(.A(men_men_n26_), .B(i_5_), .Y(men_men_n492_));
  NA3        u470(.A(men_men_n1019_), .B(men_men_n492_), .C(men_men_n132_), .Y(men_men_n493_));
  OAI220     u471(.A0(men_men_n38_), .A1(men_men_n493_), .B0(men_men_n491_), .B1(men_men_n490_), .Y(men_men_n494_));
  NA2        u472(.A(men_men_n27_), .B(i_10_), .Y(men_men_n495_));
  NO2        u473(.A(men_men_n495_), .B(men_men_n463_), .Y(men_men_n496_));
  NO3        u474(.A(men_men_n496_), .B(men_men_n494_), .C(men_men_n489_), .Y(men_men_n497_));
  NA4        u475(.A(men_men_n497_), .B(men_men_n486_), .C(men_men_n462_), .D(men_men_n459_), .Y(men_men_n498_));
  NA2        u476(.A(men_men_n167_), .B(men_men_n165_), .Y(men_men_n499_));
  OAI210     u477(.A0(men_men_n294_), .A1(men_men_n172_), .B0(men_men_n499_), .Y(men_men_n500_));
  AN2        u478(.A(men_men_n279_), .B(men_men_n228_), .Y(men_men_n501_));
  NA2        u479(.A(men_men_n501_), .B(men_men_n500_), .Y(men_men_n502_));
  NA2        u480(.A(men_men_n115_), .B(men_men_n105_), .Y(men_men_n503_));
  AO220      u481(.A0(men_men_n503_), .A1(men_men_n448_), .B0(men_men_n413_), .B1(i_6_), .Y(men_men_n504_));
  NA2        u482(.A(men_men_n305_), .B(men_men_n155_), .Y(men_men_n505_));
  OAI210     u483(.A0(men_men_n505_), .A1(men_men_n226_), .B0(men_men_n299_), .Y(men_men_n506_));
  AOI220     u484(.A0(men_men_n506_), .A1(men_men_n314_), .B0(men_men_n504_), .B1(men_men_n301_), .Y(men_men_n507_));
  NA2        u485(.A(men_men_n376_), .B(men_men_n219_), .Y(men_men_n508_));
  NA2        u486(.A(men_men_n346_), .B(men_men_n69_), .Y(men_men_n509_));
  NA2        u487(.A(men_men_n363_), .B(men_men_n355_), .Y(men_men_n510_));
  AO210      u488(.A0(men_men_n509_), .A1(men_men_n508_), .B0(men_men_n510_), .Y(men_men_n511_));
  NO2        u489(.A(men_men_n36_), .B(i_8_), .Y(men_men_n512_));
  INV        u490(.A(men_men_n413_), .Y(men_men_n513_));
  NA2        u491(.A(men_men_n513_), .B(men_men_n511_), .Y(men_men_n514_));
  INV        u492(.A(men_men_n514_), .Y(men_men_n515_));
  OAI210     u493(.A0(i_8_), .A1(men_men_n61_), .B0(men_men_n127_), .Y(men_men_n516_));
  AOI210     u494(.A0(men_men_n186_), .A1(i_9_), .B0(men_men_n258_), .Y(men_men_n517_));
  NO2        u495(.A(men_men_n517_), .B(men_men_n191_), .Y(men_men_n518_));
  AOI220     u496(.A0(i_5_), .A1(men_men_n518_), .B0(men_men_n516_), .B1(men_men_n414_), .Y(men_men_n519_));
  NA4        u497(.A(men_men_n519_), .B(men_men_n515_), .C(men_men_n507_), .D(men_men_n502_), .Y(men_men_n520_));
  NO2        u498(.A(i_12_), .B(men_men_n185_), .Y(men_men_n521_));
  NA3        u499(.A(men_men_n477_), .B(men_men_n165_), .C(men_men_n27_), .Y(men_men_n522_));
  NO3        u500(.A(men_men_n522_), .B(i_13_), .C(men_men_n460_), .Y(men_men_n523_));
  NOi31      u501(.An(men_men_n306_), .B(men_men_n412_), .C(men_men_n38_), .Y(men_men_n524_));
  OAI210     u502(.A0(men_men_n524_), .A1(men_men_n523_), .B0(men_men_n377_), .Y(men_men_n525_));
  NO2        u503(.A(i_8_), .B(i_7_), .Y(men_men_n526_));
  AOI220     u504(.A0(men_men_n315_), .A1(men_men_n39_), .B0(men_men_n229_), .B1(men_men_n199_), .Y(men_men_n527_));
  OAI220     u505(.A0(men_men_n527_), .A1(men_men_n174_), .B0(i_5_), .B1(men_men_n235_), .Y(men_men_n528_));
  NA2        u506(.A(men_men_n43_), .B(i_10_), .Y(men_men_n529_));
  NO2        u507(.A(men_men_n529_), .B(i_6_), .Y(men_men_n530_));
  NA3        u508(.A(men_men_n530_), .B(men_men_n528_), .C(men_men_n526_), .Y(men_men_n531_));
  AOI220     u509(.A0(men_men_n423_), .A1(men_men_n315_), .B0(men_men_n240_), .B1(men_men_n237_), .Y(men_men_n532_));
  OAI220     u510(.A0(men_men_n532_), .A1(i_12_), .B0(men_men_n463_), .B1(men_men_n126_), .Y(men_men_n533_));
  NA2        u511(.A(men_men_n533_), .B(men_men_n258_), .Y(men_men_n534_));
  NOi31      u512(.An(men_men_n283_), .B(men_men_n294_), .C(men_men_n172_), .Y(men_men_n535_));
  NA3        u513(.A(men_men_n298_), .B(men_men_n165_), .C(men_men_n92_), .Y(men_men_n536_));
  NO2        u514(.A(men_men_n148_), .B(i_5_), .Y(men_men_n537_));
  NA3        u515(.A(men_men_n537_), .B(men_men_n402_), .C(men_men_n309_), .Y(men_men_n538_));
  NA2        u516(.A(men_men_n538_), .B(men_men_n536_), .Y(men_men_n539_));
  OAI210     u517(.A0(men_men_n539_), .A1(men_men_n535_), .B0(men_men_n455_), .Y(men_men_n540_));
  NA4        u518(.A(men_men_n540_), .B(men_men_n534_), .C(men_men_n531_), .D(men_men_n525_), .Y(men_men_n541_));
  NA3        u519(.A(men_men_n211_), .B(men_men_n67_), .C(men_men_n43_), .Y(men_men_n542_));
  NA2        u520(.A(men_men_n276_), .B(men_men_n79_), .Y(men_men_n543_));
  AOI210     u521(.A0(men_men_n542_), .A1(men_men_n337_), .B0(men_men_n543_), .Y(men_men_n544_));
  NA2        u522(.A(men_men_n289_), .B(men_men_n279_), .Y(men_men_n545_));
  NO2        u523(.A(men_men_n545_), .B(men_men_n164_), .Y(men_men_n546_));
  NA2        u524(.A(men_men_n217_), .B(men_men_n216_), .Y(men_men_n547_));
  NA2        u525(.A(men_men_n442_), .B(men_men_n215_), .Y(men_men_n548_));
  NO2        u526(.A(men_men_n547_), .B(men_men_n548_), .Y(men_men_n549_));
  NA2        u527(.A(i_0_), .B(men_men_n47_), .Y(men_men_n550_));
  NA3        u528(.A(men_men_n521_), .B(men_men_n267_), .C(men_men_n550_), .Y(men_men_n551_));
  NO2        u529(.A(men_men_n1017_), .B(men_men_n551_), .Y(men_men_n552_));
  NO4        u530(.A(men_men_n552_), .B(men_men_n549_), .C(men_men_n546_), .D(men_men_n544_), .Y(men_men_n553_));
  NO4        u531(.A(men_men_n245_), .B(men_men_n41_), .C(i_2_), .D(men_men_n47_), .Y(men_men_n554_));
  NO3        u532(.A(i_1_), .B(i_5_), .C(i_10_), .Y(men_men_n555_));
  NO2        u533(.A(men_men_n227_), .B(men_men_n36_), .Y(men_men_n556_));
  AN2        u534(.A(men_men_n556_), .B(men_men_n555_), .Y(men_men_n557_));
  OA210      u535(.A0(men_men_n557_), .A1(men_men_n554_), .B0(men_men_n346_), .Y(men_men_n558_));
  NO2        u536(.A(men_men_n412_), .B(i_1_), .Y(men_men_n559_));
  NOi31      u537(.An(men_men_n559_), .B(men_men_n449_), .C(men_men_n69_), .Y(men_men_n560_));
  AN4        u538(.A(men_men_n560_), .B(i_9_), .C(men_men_n492_), .D(i_2_), .Y(men_men_n561_));
  NO2        u539(.A(men_men_n422_), .B(men_men_n168_), .Y(men_men_n562_));
  NO3        u540(.A(men_men_n562_), .B(men_men_n561_), .C(men_men_n558_), .Y(men_men_n563_));
  NOi21      u541(.An(i_10_), .B(i_6_), .Y(men_men_n564_));
  NO2        u542(.A(men_men_n81_), .B(men_men_n25_), .Y(men_men_n565_));
  AOI220     u543(.A0(men_men_n276_), .A1(men_men_n565_), .B0(men_men_n267_), .B1(men_men_n564_), .Y(men_men_n566_));
  NO2        u544(.A(men_men_n566_), .B(men_men_n447_), .Y(men_men_n567_));
  NO2        u545(.A(men_men_n108_), .B(men_men_n23_), .Y(men_men_n568_));
  NA2        u546(.A(men_men_n306_), .B(men_men_n155_), .Y(men_men_n569_));
  AOI220     u547(.A0(men_men_n569_), .A1(men_men_n432_), .B0(men_men_n175_), .B1(men_men_n173_), .Y(men_men_n570_));
  NO2        u548(.A(men_men_n190_), .B(men_men_n37_), .Y(men_men_n571_));
  NOi31      u549(.An(men_men_n136_), .B(men_men_n571_), .C(men_men_n323_), .Y(men_men_n572_));
  NO3        u550(.A(men_men_n572_), .B(men_men_n570_), .C(men_men_n567_), .Y(men_men_n573_));
  NO2        u551(.A(men_men_n509_), .B(men_men_n371_), .Y(men_men_n574_));
  INV        u552(.A(men_men_n309_), .Y(men_men_n575_));
  NO2        u553(.A(i_12_), .B(men_men_n81_), .Y(men_men_n576_));
  NA3        u554(.A(men_men_n379_), .B(men_men_n276_), .C(men_men_n211_), .Y(men_men_n577_));
  NO2        u555(.A(men_men_n577_), .B(men_men_n575_), .Y(men_men_n578_));
  NA2        u556(.A(men_men_n165_), .B(i_0_), .Y(men_men_n579_));
  NO3        u557(.A(men_men_n579_), .B(men_men_n330_), .C(men_men_n294_), .Y(men_men_n580_));
  OR2        u558(.A(i_2_), .B(i_5_), .Y(men_men_n581_));
  OR2        u559(.A(men_men_n581_), .B(men_men_n405_), .Y(men_men_n582_));
  INV        u560(.A(men_men_n190_), .Y(men_men_n583_));
  AOI210     u561(.A0(men_men_n583_), .A1(men_men_n582_), .B0(men_men_n490_), .Y(men_men_n584_));
  NO4        u562(.A(men_men_n584_), .B(men_men_n580_), .C(men_men_n578_), .D(men_men_n574_), .Y(men_men_n585_));
  NA4        u563(.A(men_men_n585_), .B(men_men_n573_), .C(men_men_n563_), .D(men_men_n553_), .Y(men_men_n586_));
  NO4        u564(.A(men_men_n586_), .B(men_men_n541_), .C(men_men_n520_), .D(men_men_n498_), .Y(men_men_n587_));
  NA4        u565(.A(men_men_n587_), .B(men_men_n440_), .C(men_men_n345_), .D(men_men_n304_), .Y(men7));
  NO2        u566(.A(men_men_n101_), .B(men_men_n86_), .Y(men_men_n589_));
  NA2        u567(.A(men_men_n477_), .B(men_men_n79_), .Y(men_men_n590_));
  NA2        u568(.A(i_11_), .B(men_men_n185_), .Y(men_men_n591_));
  NA3        u569(.A(i_7_), .B(i_10_), .C(i_9_), .Y(men_men_n592_));
  NA2        u570(.A(i_12_), .B(i_8_), .Y(men_men_n593_));
  AOI210     u571(.A0(men_men_n593_), .A1(men_men_n100_), .B0(men_men_n592_), .Y(men_men_n594_));
  NA2        u572(.A(i_2_), .B(men_men_n81_), .Y(men_men_n595_));
  OAI210     u573(.A0(men_men_n84_), .A1(men_men_n195_), .B0(men_men_n196_), .Y(men_men_n596_));
  NO2        u574(.A(i_7_), .B(men_men_n37_), .Y(men_men_n597_));
  NA2        u575(.A(i_4_), .B(i_8_), .Y(men_men_n598_));
  NO2        u576(.A(men_men_n594_), .B(men_men_n589_), .Y(men_men_n599_));
  OR2        u577(.A(i_6_), .B(i_10_), .Y(men_men_n600_));
  NO2        u578(.A(men_men_n600_), .B(men_men_n23_), .Y(men_men_n601_));
  NO3        u579(.A(i_6_), .B(i_8_), .C(men_men_n31_), .Y(men_men_n602_));
  INV        u580(.A(men_men_n192_), .Y(men_men_n603_));
  NO2        u581(.A(men_men_n599_), .B(men_men_n61_), .Y(men_men_n604_));
  NOi21      u582(.An(i_11_), .B(i_7_), .Y(men_men_n605_));
  AO210      u583(.A0(i_12_), .A1(i_7_), .B0(i_2_), .Y(men_men_n606_));
  NO2        u584(.A(men_men_n606_), .B(men_men_n605_), .Y(men_men_n607_));
  NA2        u585(.A(men_men_n607_), .B(men_men_n199_), .Y(men_men_n608_));
  NA3        u586(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n609_));
  NAi31      u587(.An(men_men_n609_), .B(men_men_n208_), .C(i_11_), .Y(men_men_n610_));
  AOI210     u588(.A0(men_men_n610_), .A1(men_men_n608_), .B0(men_men_n61_), .Y(men_men_n611_));
  NO3        u589(.A(men_men_n252_), .B(men_men_n201_), .C(men_men_n591_), .Y(men_men_n612_));
  OAI210     u590(.A0(men_men_n612_), .A1(men_men_n220_), .B0(men_men_n61_), .Y(men_men_n613_));
  NA2        u591(.A(men_men_n406_), .B(men_men_n31_), .Y(men_men_n614_));
  OR2        u592(.A(men_men_n201_), .B(men_men_n101_), .Y(men_men_n615_));
  NA2        u593(.A(men_men_n615_), .B(men_men_n614_), .Y(men_men_n616_));
  NO2        u594(.A(men_men_n61_), .B(i_9_), .Y(men_men_n617_));
  INV        u595(.A(i_4_), .Y(men_men_n618_));
  NA2        u596(.A(men_men_n618_), .B(men_men_n616_), .Y(men_men_n619_));
  NO2        u597(.A(i_1_), .B(i_12_), .Y(men_men_n620_));
  NA3        u598(.A(men_men_n620_), .B(men_men_n103_), .C(men_men_n24_), .Y(men_men_n621_));
  NA4        u599(.A(men_men_n621_), .B(men_men_n619_), .C(men_men_n613_), .D(men_men_n82_), .Y(men_men_n622_));
  OAI210     u600(.A0(men_men_n622_), .A1(men_men_n611_), .B0(i_6_), .Y(men_men_n623_));
  NO2        u601(.A(men_men_n609_), .B(men_men_n101_), .Y(men_men_n624_));
  NA2        u602(.A(men_men_n624_), .B(men_men_n576_), .Y(men_men_n625_));
  NO2        u603(.A(i_6_), .B(i_11_), .Y(men_men_n626_));
  NA2        u604(.A(men_men_n625_), .B(men_men_n450_), .Y(men_men_n627_));
  NA2        u605(.A(men_men_n1022_), .B(men_men_n617_), .Y(men_men_n628_));
  NO3        u606(.A(men_men_n600_), .B(men_men_n227_), .C(men_men_n23_), .Y(men_men_n629_));
  AOI210     u607(.A0(i_1_), .A1(men_men_n253_), .B0(men_men_n629_), .Y(men_men_n630_));
  OAI210     u608(.A0(men_men_n630_), .A1(men_men_n43_), .B0(men_men_n628_), .Y(men_men_n631_));
  NA3        u609(.A(men_men_n526_), .B(i_11_), .C(men_men_n36_), .Y(men_men_n632_));
  NA3        u610(.A(i_3_), .B(i_8_), .C(i_9_), .Y(men_men_n633_));
  NO2        u611(.A(men_men_n45_), .B(i_1_), .Y(men_men_n634_));
  NA3        u612(.A(men_men_n634_), .B(men_men_n259_), .C(men_men_n43_), .Y(men_men_n635_));
  NO2        u613(.A(men_men_n635_), .B(men_men_n633_), .Y(men_men_n636_));
  NO2        u614(.A(i_11_), .B(men_men_n37_), .Y(men_men_n637_));
  NA2        u615(.A(men_men_n637_), .B(men_men_n24_), .Y(men_men_n638_));
  NO2        u616(.A(men_men_n638_), .B(i_6_), .Y(men_men_n639_));
  OR2        u617(.A(men_men_n639_), .B(men_men_n636_), .Y(men_men_n640_));
  NO3        u618(.A(men_men_n640_), .B(men_men_n631_), .C(men_men_n627_), .Y(men_men_n641_));
  INV        u619(.A(men_men_n605_), .Y(men_men_n642_));
  NA2        u620(.A(men_men_n642_), .B(i_1_), .Y(men_men_n643_));
  NO2        u621(.A(men_men_n643_), .B(i_6_), .Y(men_men_n644_));
  NO2        u622(.A(men_men_n411_), .B(men_men_n81_), .Y(men_men_n645_));
  NA2        u623(.A(men_men_n644_), .B(men_men_n45_), .Y(men_men_n646_));
  NA2        u624(.A(i_3_), .B(men_men_n185_), .Y(men_men_n647_));
  NO2        u625(.A(men_men_n227_), .B(men_men_n43_), .Y(men_men_n648_));
  NO3        u626(.A(men_men_n648_), .B(men_men_n301_), .C(i_12_), .Y(men_men_n649_));
  NO2        u627(.A(men_men_n110_), .B(men_men_n37_), .Y(men_men_n650_));
  INV        u628(.A(i_6_), .Y(men_men_n651_));
  NO2        u629(.A(men_men_n81_), .B(i_9_), .Y(men_men_n652_));
  NO2        u630(.A(men_men_n652_), .B(men_men_n61_), .Y(men_men_n653_));
  NO2        u631(.A(men_men_n653_), .B(men_men_n620_), .Y(men_men_n654_));
  NO4        u632(.A(men_men_n654_), .B(men_men_n651_), .C(men_men_n649_), .D(i_4_), .Y(men_men_n655_));
  NA2        u633(.A(i_1_), .B(i_3_), .Y(men_men_n656_));
  NO2        u634(.A(men_men_n451_), .B(men_men_n88_), .Y(men_men_n657_));
  INV        u635(.A(men_men_n657_), .Y(men_men_n658_));
  NO2        u636(.A(men_men_n658_), .B(men_men_n656_), .Y(men_men_n659_));
  NO2        u637(.A(men_men_n659_), .B(men_men_n655_), .Y(men_men_n660_));
  NA4        u638(.A(men_men_n660_), .B(men_men_n646_), .C(men_men_n641_), .D(men_men_n623_), .Y(men_men_n661_));
  NO3        u639(.A(i_11_), .B(i_3_), .C(i_7_), .Y(men_men_n662_));
  OA210      u640(.A0(men_men_n662_), .A1(men_men_n238_), .B0(men_men_n81_), .Y(men_men_n663_));
  NA2        u641(.A(men_men_n363_), .B(men_men_n362_), .Y(men_men_n664_));
  NO2        u642(.A(men_men_n598_), .B(men_men_n81_), .Y(men_men_n665_));
  NA2        u643(.A(men_men_n665_), .B(men_men_n25_), .Y(men_men_n666_));
  INV        u644(.A(men_men_n666_), .Y(men_men_n667_));
  OAI210     u645(.A0(men_men_n667_), .A1(men_men_n663_), .B0(i_1_), .Y(men_men_n668_));
  NA2        u646(.A(men_men_n259_), .B(men_men_n93_), .Y(men_men_n669_));
  NO2        u647(.A(men_men_n361_), .B(i_2_), .Y(men_men_n670_));
  NA2        u648(.A(men_men_n670_), .B(men_men_n669_), .Y(men_men_n671_));
  AOI210     u649(.A0(men_men_n671_), .A1(men_men_n668_), .B0(i_13_), .Y(men_men_n672_));
  OR2        u650(.A(i_11_), .B(i_7_), .Y(men_men_n673_));
  AOI220     u651(.A0(men_men_n465_), .A1(men_men_n152_), .B0(i_2_), .B1(i_1_), .Y(men_men_n674_));
  NO2        u652(.A(men_men_n674_), .B(men_men_n43_), .Y(men_men_n675_));
  NO2        u653(.A(men_men_n471_), .B(men_men_n24_), .Y(men_men_n676_));
  AOI210     u654(.A0(men_men_n676_), .A1(men_men_n645_), .B0(men_men_n238_), .Y(men_men_n677_));
  OAI220     u655(.A0(men_men_n677_), .A1(men_men_n40_), .B0(men_men_n53_), .B1(men_men_n88_), .Y(men_men_n678_));
  AOI210     u656(.A0(men_men_n675_), .A1(men_men_n325_), .B0(men_men_n678_), .Y(men_men_n679_));
  AOI220     u657(.A0(i_12_), .A1(men_men_n68_), .B0(men_men_n379_), .B1(men_men_n634_), .Y(men_men_n680_));
  NO2        u658(.A(men_men_n680_), .B(men_men_n235_), .Y(men_men_n681_));
  AOI210     u659(.A0(men_men_n443_), .A1(men_men_n36_), .B0(i_13_), .Y(men_men_n682_));
  NO2        u660(.A(men_men_n590_), .B(men_men_n43_), .Y(men_men_n683_));
  NO2        u661(.A(men_men_n633_), .B(men_men_n108_), .Y(men_men_n684_));
  NO3        u662(.A(men_men_n67_), .B(men_men_n32_), .C(men_men_n97_), .Y(men_men_n685_));
  NA2        u663(.A(i_3_), .B(i_7_), .Y(men_men_n686_));
  NO3        u664(.A(men_men_n471_), .B(men_men_n231_), .C(men_men_n81_), .Y(men_men_n687_));
  AOI210     u665(.A0(men_men_n687_), .A1(men_men_n686_), .B0(men_men_n685_), .Y(men_men_n688_));
  NA2        u666(.A(men_men_n379_), .B(men_men_n634_), .Y(men_men_n689_));
  OAI220     u667(.A0(men_men_n689_), .A1(men_men_n593_), .B0(men_men_n688_), .B1(men_men_n603_), .Y(men_men_n690_));
  NO4        u668(.A(men_men_n690_), .B(men_men_n684_), .C(men_men_n683_), .D(men_men_n681_), .Y(men_men_n691_));
  NA3        u669(.A(men_men_n406_), .B(men_men_n597_), .C(men_men_n93_), .Y(men_men_n692_));
  NA2        u670(.A(men_men_n626_), .B(i_13_), .Y(men_men_n693_));
  NAi21      u671(.An(i_11_), .B(i_12_), .Y(men_men_n694_));
  NOi41      u672(.An(men_men_n104_), .B(men_men_n694_), .C(i_13_), .D(men_men_n81_), .Y(men_men_n695_));
  NO3        u673(.A(men_men_n471_), .B(men_men_n576_), .C(men_men_n598_), .Y(men_men_n696_));
  AOI210     u674(.A0(men_men_n696_), .A1(men_men_n305_), .B0(men_men_n695_), .Y(men_men_n697_));
  NA3        u675(.A(men_men_n697_), .B(men_men_n693_), .C(men_men_n692_), .Y(men_men_n698_));
  NA2        u676(.A(men_men_n698_), .B(men_men_n61_), .Y(men_men_n699_));
  NA2        u677(.A(i_8_), .B(men_men_n25_), .Y(men_men_n700_));
  NO3        u678(.A(men_men_n700_), .B(men_men_n377_), .C(i_12_), .Y(men_men_n701_));
  OAI210     u679(.A0(men_men_n701_), .A1(men_men_n362_), .B0(men_men_n360_), .Y(men_men_n702_));
  NO2        u680(.A(men_men_n121_), .B(i_2_), .Y(men_men_n703_));
  INV        u681(.A(men_men_n703_), .Y(men_men_n704_));
  NA2        u682(.A(men_men_n704_), .B(men_men_n702_), .Y(men_men_n705_));
  NA3        u683(.A(men_men_n705_), .B(men_men_n44_), .C(men_men_n219_), .Y(men_men_n706_));
  NA4        u684(.A(men_men_n706_), .B(men_men_n699_), .C(men_men_n691_), .D(men_men_n679_), .Y(men_men_n707_));
  OR4        u685(.A(men_men_n707_), .B(men_men_n672_), .C(men_men_n661_), .D(men_men_n604_), .Y(men5));
  AOI210     u686(.A0(men_men_n642_), .A1(men_men_n262_), .B0(men_men_n414_), .Y(men_men_n709_));
  NO3        u687(.A(i_11_), .B(men_men_n231_), .C(i_13_), .Y(men_men_n710_));
  NO2        u688(.A(men_men_n117_), .B(men_men_n23_), .Y(men_men_n711_));
  NA2        u689(.A(i_12_), .B(i_8_), .Y(men_men_n712_));
  OAI210     u690(.A0(men_men_n45_), .A1(i_3_), .B0(men_men_n712_), .Y(men_men_n713_));
  INV        u691(.A(men_men_n442_), .Y(men_men_n714_));
  AOI220     u692(.A0(men_men_n309_), .A1(men_men_n568_), .B0(men_men_n713_), .B1(men_men_n711_), .Y(men_men_n715_));
  INV        u693(.A(men_men_n715_), .Y(men_men_n716_));
  NO2        u694(.A(men_men_n716_), .B(men_men_n1013_), .Y(men_men_n717_));
  INV        u695(.A(men_men_n162_), .Y(men_men_n718_));
  INV        u696(.A(men_men_n238_), .Y(men_men_n719_));
  OAI210     u697(.A0(men_men_n670_), .A1(men_men_n444_), .B0(men_men_n104_), .Y(men_men_n720_));
  AOI210     u698(.A0(men_men_n720_), .A1(men_men_n719_), .B0(men_men_n718_), .Y(men_men_n721_));
  NO2        u699(.A(men_men_n451_), .B(men_men_n26_), .Y(men_men_n722_));
  NO2        u700(.A(men_men_n722_), .B(men_men_n415_), .Y(men_men_n723_));
  NA2        u701(.A(men_men_n723_), .B(i_2_), .Y(men_men_n724_));
  INV        u702(.A(men_men_n724_), .Y(men_men_n725_));
  AOI210     u703(.A0(men_men_n33_), .A1(men_men_n36_), .B0(men_men_n412_), .Y(men_men_n726_));
  AOI210     u704(.A0(men_men_n726_), .A1(men_men_n725_), .B0(men_men_n721_), .Y(men_men_n727_));
  NO2        u705(.A(men_men_n182_), .B(men_men_n118_), .Y(men_men_n728_));
  OAI210     u706(.A0(men_men_n728_), .A1(men_men_n711_), .B0(i_2_), .Y(men_men_n729_));
  INV        u707(.A(men_men_n163_), .Y(men_men_n730_));
  NO3        u708(.A(men_men_n606_), .B(men_men_n38_), .C(men_men_n26_), .Y(men_men_n731_));
  AOI210     u709(.A0(men_men_n730_), .A1(men_men_n84_), .B0(men_men_n731_), .Y(men_men_n732_));
  AOI210     u710(.A0(men_men_n732_), .A1(men_men_n729_), .B0(men_men_n185_), .Y(men_men_n733_));
  OA210      u711(.A0(men_men_n607_), .A1(men_men_n119_), .B0(i_13_), .Y(men_men_n734_));
  AOI210     u712(.A0(men_men_n201_), .A1(men_men_n138_), .B0(men_men_n512_), .Y(men_men_n735_));
  NA2        u713(.A(men_men_n735_), .B(men_men_n415_), .Y(men_men_n736_));
  NA3        u714(.A(men_men_n298_), .B(men_men_n117_), .C(men_men_n41_), .Y(men_men_n737_));
  OAI210     u715(.A0(men_men_n737_), .A1(i_11_), .B0(men_men_n736_), .Y(men_men_n738_));
  NO3        u716(.A(men_men_n738_), .B(men_men_n734_), .C(men_men_n733_), .Y(men_men_n739_));
  NA2        u717(.A(men_men_n568_), .B(men_men_n28_), .Y(men_men_n740_));
  NA2        u718(.A(men_men_n710_), .B(men_men_n268_), .Y(men_men_n741_));
  NA2        u719(.A(men_men_n741_), .B(men_men_n740_), .Y(men_men_n742_));
  NO2        u720(.A(men_men_n60_), .B(i_12_), .Y(men_men_n743_));
  NO2        u721(.A(men_men_n743_), .B(men_men_n119_), .Y(men_men_n744_));
  NO2        u722(.A(men_men_n744_), .B(men_men_n591_), .Y(men_men_n745_));
  AOI210     u723(.A0(men_men_n745_), .A1(men_men_n36_), .B0(men_men_n742_), .Y(men_men_n746_));
  NA4        u724(.A(men_men_n746_), .B(men_men_n739_), .C(men_men_n727_), .D(men_men_n717_), .Y(men6));
  NO2        u725(.A(men_men_n177_), .B(i_9_), .Y(men_men_n748_));
  OAI210     u726(.A0(men_men_n748_), .A1(i_5_), .B0(men_men_n703_), .Y(men_men_n749_));
  NA4        u727(.A(men_men_n383_), .B(men_men_n476_), .C(men_men_n67_), .D(men_men_n97_), .Y(men_men_n750_));
  INV        u728(.A(men_men_n750_), .Y(men_men_n751_));
  NO2        u729(.A(men_men_n214_), .B(men_men_n481_), .Y(men_men_n752_));
  NO2        u730(.A(men_men_n751_), .B(men_men_n320_), .Y(men_men_n753_));
  AO210      u731(.A0(men_men_n753_), .A1(men_men_n749_), .B0(i_12_), .Y(men_men_n754_));
  NA2        u732(.A(men_men_n366_), .B(men_men_n327_), .Y(men_men_n755_));
  NA2        u733(.A(men_men_n576_), .B(men_men_n61_), .Y(men_men_n756_));
  NA2        u734(.A(men_men_n756_), .B(men_men_n755_), .Y(men_men_n757_));
  INV        u735(.A(men_men_n189_), .Y(men_men_n758_));
  AOI210     u736(.A0(men_men_n757_), .A1(men_men_n69_), .B0(men_men_n758_), .Y(men_men_n759_));
  NA2        u737(.A(men_men_n1014_), .B(men_men_n743_), .Y(men_men_n760_));
  NO2        u738(.A(men_men_n760_), .B(men_men_n177_), .Y(men_men_n761_));
  NO2        u739(.A(men_men_n32_), .B(i_11_), .Y(men_men_n762_));
  OAI210     u740(.A0(men_men_n662_), .A1(men_men_n556_), .B0(men_men_n555_), .Y(men_men_n763_));
  INV        u741(.A(men_men_n763_), .Y(men_men_n764_));
  OR2        u742(.A(men_men_n764_), .B(men_men_n761_), .Y(men_men_n765_));
  NA2        u743(.A(men_men_n47_), .B(men_men_n37_), .Y(men_men_n766_));
  OAI210     u744(.A0(men_men_n766_), .A1(men_men_n405_), .B0(men_men_n350_), .Y(men_men_n767_));
  NA2        u745(.A(men_men_n767_), .B(men_men_n1021_), .Y(men_men_n768_));
  AO210      u746(.A0(men_men_n349_), .A1(men_men_n341_), .B0(men_men_n391_), .Y(men_men_n769_));
  NA2        u747(.A(men_men_n769_), .B(i_7_), .Y(men_men_n770_));
  NA3        u748(.A(men_men_n444_), .B(men_men_n137_), .C(men_men_n65_), .Y(men_men_n771_));
  AO210      u749(.A0(men_men_n488_), .A1(men_men_n714_), .B0(men_men_n36_), .Y(men_men_n772_));
  NA4        u750(.A(men_men_n772_), .B(men_men_n771_), .C(men_men_n770_), .D(men_men_n768_), .Y(men_men_n773_));
  INV        u751(.A(men_men_n752_), .Y(men_men_n774_));
  NA3        u752(.A(men_men_n365_), .B(men_men_n232_), .C(men_men_n137_), .Y(men_men_n775_));
  NA2        u753(.A(men_men_n391_), .B(men_men_n66_), .Y(men_men_n776_));
  NA4        u754(.A(men_men_n776_), .B(men_men_n775_), .C(men_men_n774_), .D(men_men_n596_), .Y(men_men_n777_));
  AO210      u755(.A0(men_men_n512_), .A1(men_men_n45_), .B0(men_men_n83_), .Y(men_men_n778_));
  NA3        u756(.A(men_men_n778_), .B(men_men_n477_), .C(men_men_n211_), .Y(men_men_n779_));
  AOI210     u757(.A0(men_men_n444_), .A1(men_men_n442_), .B0(men_men_n554_), .Y(men_men_n780_));
  NA2        u758(.A(men_men_n237_), .B(men_men_n45_), .Y(men_men_n781_));
  INV        u759(.A(men_men_n582_), .Y(men_men_n782_));
  NA3        u760(.A(men_men_n782_), .B(men_men_n319_), .C(i_7_), .Y(men_men_n783_));
  NA4        u761(.A(men_men_n783_), .B(men_men_n1020_), .C(men_men_n780_), .D(men_men_n779_), .Y(men_men_n784_));
  NO4        u762(.A(men_men_n784_), .B(men_men_n777_), .C(men_men_n773_), .D(men_men_n765_), .Y(men_men_n785_));
  NA4        u763(.A(men_men_n785_), .B(men_men_n759_), .C(men_men_n754_), .D(men_men_n373_), .Y(men3));
  NA2        u764(.A(i_12_), .B(i_10_), .Y(men_men_n787_));
  NA2        u765(.A(i_6_), .B(i_7_), .Y(men_men_n788_));
  NO2        u766(.A(men_men_n788_), .B(i_0_), .Y(men_men_n789_));
  NO2        u767(.A(i_11_), .B(men_men_n231_), .Y(men_men_n790_));
  OAI210     u768(.A0(men_men_n789_), .A1(men_men_n283_), .B0(men_men_n790_), .Y(men_men_n791_));
  NO2        u769(.A(men_men_n791_), .B(men_men_n185_), .Y(men_men_n792_));
  NO3        u770(.A(men_men_n447_), .B(men_men_n86_), .C(men_men_n43_), .Y(men_men_n793_));
  OA210      u771(.A0(men_men_n793_), .A1(men_men_n792_), .B0(men_men_n165_), .Y(men_men_n794_));
  NA3        u772(.A(men_men_n775_), .B(men_men_n596_), .C(men_men_n364_), .Y(men_men_n795_));
  NA2        u773(.A(men_men_n795_), .B(men_men_n39_), .Y(men_men_n796_));
  NOi21      u774(.An(men_men_n92_), .B(men_men_n723_), .Y(men_men_n797_));
  NO3        u775(.A(men_men_n615_), .B(men_men_n451_), .C(men_men_n124_), .Y(men_men_n798_));
  NA2        u776(.A(men_men_n406_), .B(men_men_n44_), .Y(men_men_n799_));
  AN2        u777(.A(men_men_n449_), .B(men_men_n54_), .Y(men_men_n800_));
  NO3        u778(.A(men_men_n800_), .B(men_men_n798_), .C(men_men_n797_), .Y(men_men_n801_));
  AOI210     u779(.A0(men_men_n801_), .A1(men_men_n796_), .B0(men_men_n47_), .Y(men_men_n802_));
  NO4        u780(.A(men_men_n369_), .B(men_men_n376_), .C(men_men_n38_), .D(i_0_), .Y(men_men_n803_));
  NA2        u781(.A(men_men_n177_), .B(men_men_n564_), .Y(men_men_n804_));
  NOi21      u782(.An(men_men_n804_), .B(men_men_n803_), .Y(men_men_n805_));
  NA2        u783(.A(men_men_n682_), .B(men_men_n652_), .Y(men_men_n806_));
  NA2        u784(.A(i_0_), .B(men_men_n434_), .Y(men_men_n807_));
  OAI220     u785(.A0(men_men_n807_), .A1(men_men_n806_), .B0(men_men_n805_), .B1(men_men_n61_), .Y(men_men_n808_));
  NOi21      u786(.An(i_5_), .B(i_9_), .Y(men_men_n809_));
  NA2        u787(.A(men_men_n809_), .B(men_men_n441_), .Y(men_men_n810_));
  NO3        u788(.A(men_men_n409_), .B(men_men_n259_), .C(men_men_n69_), .Y(men_men_n811_));
  NO2        u789(.A(men_men_n166_), .B(men_men_n138_), .Y(men_men_n812_));
  AOI210     u790(.A0(men_men_n812_), .A1(men_men_n237_), .B0(men_men_n811_), .Y(men_men_n813_));
  OAI220     u791(.A0(men_men_n813_), .A1(men_men_n172_), .B0(men_men_n598_), .B1(men_men_n810_), .Y(men_men_n814_));
  NO4        u792(.A(men_men_n814_), .B(men_men_n808_), .C(men_men_n802_), .D(men_men_n794_), .Y(men_men_n815_));
  NA2        u793(.A(men_men_n177_), .B(men_men_n24_), .Y(men_men_n816_));
  NO2        u794(.A(men_men_n650_), .B(men_men_n589_), .Y(men_men_n817_));
  NO2        u795(.A(men_men_n817_), .B(men_men_n816_), .Y(men_men_n818_));
  NA2        u796(.A(men_men_n305_), .B(men_men_n122_), .Y(men_men_n819_));
  NAi21      u797(.An(men_men_n153_), .B(men_men_n434_), .Y(men_men_n820_));
  OAI220     u798(.A0(men_men_n820_), .A1(men_men_n781_), .B0(men_men_n819_), .B1(men_men_n395_), .Y(men_men_n821_));
  NO2        u799(.A(men_men_n821_), .B(men_men_n818_), .Y(men_men_n822_));
  INV        u800(.A(men_men_n287_), .Y(men_men_n823_));
  NA2        u801(.A(men_men_n823_), .B(men_men_n684_), .Y(men_men_n824_));
  NA2        u802(.A(men_men_n565_), .B(i_0_), .Y(men_men_n825_));
  NO3        u803(.A(men_men_n825_), .B(men_men_n378_), .C(men_men_n84_), .Y(men_men_n826_));
  NO4        u804(.A(men_men_n581_), .B(men_men_n208_), .C(men_men_n412_), .D(men_men_n405_), .Y(men_men_n827_));
  AOI210     u805(.A0(men_men_n827_), .A1(i_11_), .B0(men_men_n826_), .Y(men_men_n828_));
  AN2        u806(.A(men_men_n92_), .B(men_men_n236_), .Y(men_men_n829_));
  NA2        u807(.A(men_men_n710_), .B(men_men_n320_), .Y(men_men_n830_));
  AOI210     u808(.A0(men_men_n477_), .A1(men_men_n84_), .B0(men_men_n57_), .Y(men_men_n831_));
  NO2        u809(.A(men_men_n831_), .B(men_men_n830_), .Y(men_men_n832_));
  NO2        u810(.A(men_men_n246_), .B(men_men_n144_), .Y(men_men_n833_));
  NA2        u811(.A(i_0_), .B(i_10_), .Y(men_men_n834_));
  OAI210     u812(.A0(men_men_n834_), .A1(men_men_n81_), .B0(men_men_n529_), .Y(men_men_n835_));
  NO4        u813(.A(men_men_n108_), .B(men_men_n57_), .C(men_men_n647_), .D(i_5_), .Y(men_men_n836_));
  AO220      u814(.A0(men_men_n836_), .A1(men_men_n835_), .B0(men_men_n833_), .B1(i_6_), .Y(men_men_n837_));
  NA2        u815(.A(men_men_n559_), .B(i_4_), .Y(men_men_n838_));
  OAI220     u816(.A0(i_1_), .A1(men_men_n830_), .B0(men_men_n838_), .B1(men_men_n1018_), .Y(men_men_n839_));
  NO4        u817(.A(men_men_n839_), .B(men_men_n837_), .C(men_men_n832_), .D(men_men_n829_), .Y(men_men_n840_));
  NA4        u818(.A(men_men_n840_), .B(men_men_n828_), .C(men_men_n824_), .D(men_men_n822_), .Y(men_men_n841_));
  NO2        u819(.A(men_men_n98_), .B(men_men_n37_), .Y(men_men_n842_));
  NA2        u820(.A(i_11_), .B(i_9_), .Y(men_men_n843_));
  NO3        u821(.A(i_12_), .B(men_men_n843_), .C(men_men_n595_), .Y(men_men_n844_));
  AN2        u822(.A(men_men_n844_), .B(men_men_n842_), .Y(men_men_n845_));
  NO2        u823(.A(men_men_n47_), .B(i_7_), .Y(men_men_n846_));
  NA2        u824(.A(men_men_n454_), .B(men_men_n151_), .Y(men_men_n847_));
  NO2        u825(.A(men_men_n843_), .B(men_men_n69_), .Y(men_men_n848_));
  NO2        u826(.A(men_men_n166_), .B(i_0_), .Y(men_men_n849_));
  INV        u827(.A(men_men_n849_), .Y(men_men_n850_));
  NA2        u828(.A(men_men_n469_), .B(men_men_n225_), .Y(men_men_n851_));
  INV        u829(.A(men_men_n403_), .Y(men_men_n852_));
  OAI220     u830(.A0(men_men_n852_), .A1(men_men_n810_), .B0(men_men_n851_), .B1(men_men_n850_), .Y(men_men_n853_));
  NO3        u831(.A(men_men_n853_), .B(men_men_n847_), .C(men_men_n845_), .Y(men_men_n854_));
  NA2        u832(.A(men_men_n637_), .B(men_men_n114_), .Y(men_men_n855_));
  NO2        u833(.A(i_6_), .B(men_men_n855_), .Y(men_men_n856_));
  AOI210     u834(.A0(men_men_n443_), .A1(men_men_n36_), .B0(i_3_), .Y(men_men_n857_));
  NA2        u835(.A(men_men_n162_), .B(men_men_n98_), .Y(men_men_n858_));
  NOi32      u836(.An(men_men_n857_), .Bn(men_men_n180_), .C(men_men_n858_), .Y(men_men_n859_));
  AOI210     u837(.A0(men_men_n597_), .A1(men_men_n320_), .B0(men_men_n236_), .Y(men_men_n860_));
  NO2        u838(.A(men_men_n860_), .B(men_men_n799_), .Y(men_men_n861_));
  NO3        u839(.A(men_men_n861_), .B(men_men_n859_), .C(men_men_n856_), .Y(men_men_n862_));
  NOi21      u840(.An(i_7_), .B(i_5_), .Y(men_men_n863_));
  NOi31      u841(.An(men_men_n863_), .B(i_0_), .C(men_men_n694_), .Y(men_men_n864_));
  NA3        u842(.A(men_men_n864_), .B(men_men_n377_), .C(i_6_), .Y(men_men_n865_));
  OA210      u843(.A0(men_men_n858_), .A1(men_men_n510_), .B0(men_men_n865_), .Y(men_men_n866_));
  INV        u844(.A(men_men_n310_), .Y(men_men_n867_));
  NA3        u845(.A(men_men_n866_), .B(men_men_n862_), .C(men_men_n854_), .Y(men_men_n868_));
  NO2        u846(.A(men_men_n816_), .B(men_men_n233_), .Y(men_men_n869_));
  AN2        u847(.A(men_men_n325_), .B(men_men_n320_), .Y(men_men_n870_));
  AN2        u848(.A(men_men_n870_), .B(men_men_n812_), .Y(men_men_n871_));
  OAI210     u849(.A0(men_men_n871_), .A1(men_men_n869_), .B0(i_10_), .Y(men_men_n872_));
  NO2        u850(.A(men_men_n787_), .B(men_men_n309_), .Y(men_men_n873_));
  OA210      u851(.A0(men_men_n469_), .A1(men_men_n217_), .B0(men_men_n468_), .Y(men_men_n874_));
  NA2        u852(.A(men_men_n873_), .B(men_men_n848_), .Y(men_men_n875_));
  NA3        u853(.A(men_men_n468_), .B(men_men_n406_), .C(men_men_n44_), .Y(men_men_n876_));
  OAI210     u854(.A0(men_men_n820_), .A1(i_7_), .B0(men_men_n876_), .Y(men_men_n877_));
  NO2        u855(.A(men_men_n249_), .B(men_men_n45_), .Y(men_men_n878_));
  NA2        u856(.A(men_men_n848_), .B(men_men_n298_), .Y(men_men_n879_));
  OAI210     u857(.A0(men_men_n878_), .A1(men_men_n179_), .B0(men_men_n879_), .Y(men_men_n880_));
  AOI220     u858(.A0(men_men_n880_), .A1(men_men_n469_), .B0(men_men_n877_), .B1(men_men_n69_), .Y(men_men_n881_));
  NA3        u859(.A(men_men_n766_), .B(men_men_n375_), .C(i_6_), .Y(men_men_n882_));
  NA2        u860(.A(men_men_n88_), .B(men_men_n43_), .Y(men_men_n883_));
  NO2        u861(.A(men_men_n71_), .B(men_men_n712_), .Y(men_men_n884_));
  AOI220     u862(.A0(men_men_n884_), .A1(men_men_n883_), .B0(men_men_n165_), .B1(men_men_n589_), .Y(men_men_n885_));
  AOI210     u863(.A0(men_men_n885_), .A1(men_men_n882_), .B0(men_men_n46_), .Y(men_men_n886_));
  NO3        u864(.A(men_men_n581_), .B(i_0_), .C(men_men_n24_), .Y(men_men_n887_));
  AOI210     u865(.A0(men_men_n676_), .A1(men_men_n537_), .B0(men_men_n887_), .Y(men_men_n888_));
  NAi21      u866(.An(i_9_), .B(i_5_), .Y(men_men_n889_));
  NO2        u867(.A(men_men_n889_), .B(men_men_n398_), .Y(men_men_n890_));
  NO2        u868(.A(men_men_n592_), .B(men_men_n100_), .Y(men_men_n891_));
  AOI220     u869(.A0(men_men_n891_), .A1(i_0_), .B0(men_men_n890_), .B1(men_men_n607_), .Y(men_men_n892_));
  OAI220     u870(.A0(men_men_n892_), .A1(men_men_n81_), .B0(men_men_n888_), .B1(men_men_n163_), .Y(men_men_n893_));
  NO3        u871(.A(men_men_n893_), .B(men_men_n886_), .C(men_men_n514_), .Y(men_men_n894_));
  NA4        u872(.A(men_men_n894_), .B(men_men_n881_), .C(men_men_n875_), .D(men_men_n872_), .Y(men_men_n895_));
  NO3        u873(.A(men_men_n895_), .B(men_men_n868_), .C(men_men_n841_), .Y(men_men_n896_));
  NO2        u874(.A(i_0_), .B(men_men_n694_), .Y(men_men_n897_));
  NA2        u875(.A(men_men_n69_), .B(men_men_n43_), .Y(men_men_n898_));
  NO3        u876(.A(men_men_n100_), .B(i_5_), .C(men_men_n25_), .Y(men_men_n899_));
  AO220      u877(.A0(men_men_n899_), .A1(men_men_n43_), .B0(men_men_n897_), .B1(men_men_n165_), .Y(men_men_n900_));
  AOI210     u878(.A0(men_men_n756_), .A1(men_men_n664_), .B0(men_men_n858_), .Y(men_men_n901_));
  AOI210     u879(.A0(men_men_n900_), .A1(men_men_n338_), .B0(men_men_n901_), .Y(men_men_n902_));
  NA2        u880(.A(men_men_n703_), .B(men_men_n136_), .Y(men_men_n903_));
  NO2        u881(.A(men_men_n763_), .B(men_men_n398_), .Y(men_men_n904_));
  NA3        u882(.A(men_men_n789_), .B(i_2_), .C(men_men_n47_), .Y(men_men_n905_));
  NA2        u883(.A(men_men_n790_), .B(i_9_), .Y(men_men_n906_));
  AOI210     u884(.A0(men_men_n905_), .A1(men_men_n493_), .B0(men_men_n906_), .Y(men_men_n907_));
  OAI210     u885(.A0(men_men_n237_), .A1(i_9_), .B0(men_men_n224_), .Y(men_men_n908_));
  AOI210     u886(.A0(men_men_n908_), .A1(men_men_n825_), .B0(men_men_n144_), .Y(men_men_n909_));
  NO3        u887(.A(men_men_n909_), .B(men_men_n907_), .C(men_men_n904_), .Y(men_men_n910_));
  NA3        u888(.A(men_men_n910_), .B(men_men_n903_), .C(men_men_n902_), .Y(men_men_n911_));
  NA2        u889(.A(men_men_n870_), .B(men_men_n365_), .Y(men_men_n912_));
  AOI210     u890(.A0(men_men_n294_), .A1(men_men_n153_), .B0(men_men_n912_), .Y(men_men_n913_));
  INV        u891(.A(men_men_n913_), .Y(men_men_n914_));
  NO2        u892(.A(men_men_n834_), .B(men_men_n182_), .Y(men_men_n915_));
  NA2        u893(.A(men_men_n915_), .B(i_11_), .Y(men_men_n916_));
  NA2        u894(.A(men_men_n72_), .B(i_13_), .Y(men_men_n917_));
  INV        u895(.A(men_men_n211_), .Y(men_men_n918_));
  NO2        u896(.A(i_12_), .B(men_men_n603_), .Y(men_men_n919_));
  NA3        u897(.A(men_men_n919_), .B(men_men_n1015_), .C(men_men_n918_), .Y(men_men_n920_));
  NA4        u898(.A(men_men_n920_), .B(men_men_n917_), .C(men_men_n916_), .D(men_men_n914_), .Y(men_men_n921_));
  NO2        u899(.A(men_men_n235_), .B(men_men_n88_), .Y(men_men_n922_));
  AOI210     u900(.A0(men_men_n922_), .A1(men_men_n897_), .B0(men_men_n102_), .Y(men_men_n923_));
  AOI220     u901(.A0(men_men_n863_), .A1(men_men_n482_), .B0(men_men_n789_), .B1(men_men_n154_), .Y(men_men_n924_));
  NA2        u902(.A(men_men_n341_), .B(men_men_n167_), .Y(men_men_n925_));
  OA220      u903(.A0(men_men_n925_), .A1(men_men_n924_), .B0(men_men_n923_), .B1(i_5_), .Y(men_men_n926_));
  AOI210     u904(.A0(i_0_), .A1(men_men_n25_), .B0(men_men_n166_), .Y(men_men_n927_));
  NA2        u905(.A(men_men_n927_), .B(men_men_n874_), .Y(men_men_n928_));
  NA3        u906(.A(men_men_n601_), .B(men_men_n177_), .C(men_men_n79_), .Y(men_men_n929_));
  NA2        u907(.A(men_men_n929_), .B(men_men_n536_), .Y(men_men_n930_));
  NO3        u908(.A(men_men_n799_), .B(men_men_n53_), .C(men_men_n47_), .Y(men_men_n931_));
  NA3        u909(.A(men_men_n487_), .B(men_men_n480_), .C(men_men_n466_), .Y(men_men_n932_));
  NO3        u910(.A(men_men_n932_), .B(men_men_n931_), .C(men_men_n930_), .Y(men_men_n933_));
  NA2        u911(.A(men_men_n383_), .B(men_men_n161_), .Y(men_men_n934_));
  NA3        u912(.A(men_men_n383_), .B(men_men_n326_), .C(men_men_n215_), .Y(men_men_n935_));
  INV        u913(.A(men_men_n935_), .Y(men_men_n936_));
  NOi31      u914(.An(men_men_n382_), .B(men_men_n898_), .C(men_men_n233_), .Y(men_men_n937_));
  NO3        u915(.A(men_men_n937_), .B(men_men_n936_), .C(men_men_n1012_), .Y(men_men_n938_));
  NA4        u916(.A(men_men_n938_), .B(men_men_n933_), .C(men_men_n928_), .D(men_men_n926_), .Y(men_men_n939_));
  INV        u917(.A(men_men_n602_), .Y(men_men_n940_));
  NO3        u918(.A(men_men_n940_), .B(men_men_n550_), .C(i_3_), .Y(men_men_n941_));
  NO2        u919(.A(men_men_n81_), .B(i_5_), .Y(men_men_n942_));
  NA3        u920(.A(men_men_n790_), .B(men_men_n103_), .C(men_men_n117_), .Y(men_men_n943_));
  INV        u921(.A(men_men_n943_), .Y(men_men_n944_));
  AOI210     u922(.A0(men_men_n944_), .A1(men_men_n942_), .B0(men_men_n941_), .Y(men_men_n945_));
  NA3        u923(.A(men_men_n298_), .B(i_5_), .C(men_men_n185_), .Y(men_men_n946_));
  NO4        u924(.A(men_men_n233_), .B(men_men_n203_), .C(i_0_), .D(i_12_), .Y(men_men_n947_));
  AOI220     u925(.A0(men_men_n947_), .A1(i_10_), .B0(men_men_n751_), .B1(men_men_n167_), .Y(men_men_n948_));
  AN2        u926(.A(men_men_n834_), .B(men_men_n144_), .Y(men_men_n949_));
  NO4        u927(.A(men_men_n949_), .B(i_12_), .C(men_men_n632_), .D(men_men_n124_), .Y(men_men_n950_));
  NA2        u928(.A(men_men_n950_), .B(men_men_n211_), .Y(men_men_n951_));
  NA3        u929(.A(men_men_n94_), .B(men_men_n564_), .C(i_11_), .Y(men_men_n952_));
  NO2        u930(.A(men_men_n952_), .B(men_men_n146_), .Y(men_men_n953_));
  NA2        u931(.A(men_men_n863_), .B(men_men_n465_), .Y(men_men_n954_));
  NA2        u932(.A(men_men_n62_), .B(men_men_n97_), .Y(men_men_n955_));
  OAI220     u933(.A0(men_men_n955_), .A1(men_men_n946_), .B0(men_men_n954_), .B1(men_men_n653_), .Y(men_men_n956_));
  AOI210     u934(.A0(men_men_n956_), .A1(men_men_n849_), .B0(men_men_n953_), .Y(men_men_n957_));
  NA4        u935(.A(men_men_n957_), .B(men_men_n951_), .C(men_men_n948_), .D(men_men_n945_), .Y(men_men_n958_));
  NO4        u936(.A(men_men_n958_), .B(men_men_n939_), .C(men_men_n921_), .D(men_men_n911_), .Y(men_men_n959_));
  NA2        u937(.A(men_men_n762_), .B(men_men_n37_), .Y(men_men_n960_));
  NA3        u938(.A(men_men_n857_), .B(men_men_n360_), .C(i_5_), .Y(men_men_n961_));
  NA2        u939(.A(men_men_n961_), .B(men_men_n960_), .Y(men_men_n962_));
  NA2        u940(.A(men_men_n962_), .B(men_men_n199_), .Y(men_men_n963_));
  AN2        u941(.A(men_men_n673_), .B(men_men_n361_), .Y(men_men_n964_));
  NA2        u942(.A(men_men_n178_), .B(men_men_n180_), .Y(men_men_n965_));
  AO210      u943(.A0(men_men_n964_), .A1(men_men_n33_), .B0(men_men_n965_), .Y(men_men_n966_));
  NA2        u944(.A(men_men_n601_), .B(men_men_n309_), .Y(men_men_n967_));
  NAi31      u945(.An(i_7_), .B(i_2_), .C(i_10_), .Y(men_men_n968_));
  NO2        u946(.A(men_men_n66_), .B(men_men_n968_), .Y(men_men_n969_));
  NO2        u947(.A(men_men_n969_), .B(men_men_n629_), .Y(men_men_n970_));
  NA3        u948(.A(men_men_n970_), .B(men_men_n967_), .C(men_men_n966_), .Y(men_men_n971_));
  NO2        u949(.A(men_men_n457_), .B(men_men_n259_), .Y(men_men_n972_));
  NO4        u950(.A(men_men_n227_), .B(men_men_n135_), .C(men_men_n656_), .D(men_men_n37_), .Y(men_men_n973_));
  NO3        u951(.A(men_men_n973_), .B(men_men_n972_), .C(men_men_n827_), .Y(men_men_n974_));
  OAI210     u952(.A0(men_men_n952_), .A1(men_men_n138_), .B0(men_men_n974_), .Y(men_men_n975_));
  AOI210     u953(.A0(men_men_n971_), .A1(men_men_n47_), .B0(men_men_n975_), .Y(men_men_n976_));
  AOI210     u954(.A0(men_men_n976_), .A1(men_men_n963_), .B0(men_men_n69_), .Y(men_men_n977_));
  INV        u955(.A(men_men_n372_), .Y(men_men_n978_));
  NO2        u956(.A(men_men_n978_), .B(men_men_n718_), .Y(men_men_n979_));
  OAI210     u957(.A0(men_men_n76_), .A1(men_men_n53_), .B0(men_men_n101_), .Y(men_men_n980_));
  NA2        u958(.A(men_men_n980_), .B(men_men_n72_), .Y(men_men_n981_));
  AOI210     u959(.A0(men_men_n927_), .A1(men_men_n846_), .B0(men_men_n864_), .Y(men_men_n982_));
  AOI210     u960(.A0(men_men_n982_), .A1(men_men_n981_), .B0(men_men_n656_), .Y(men_men_n983_));
  NA2        u961(.A(men_men_n256_), .B(men_men_n56_), .Y(men_men_n984_));
  AOI220     u962(.A0(men_men_n984_), .A1(men_men_n72_), .B0(men_men_n336_), .B1(men_men_n248_), .Y(men_men_n985_));
  NO2        u963(.A(men_men_n985_), .B(men_men_n231_), .Y(men_men_n986_));
  NA3        u964(.A(men_men_n92_), .B(men_men_n300_), .C(men_men_n31_), .Y(men_men_n987_));
  INV        u965(.A(men_men_n987_), .Y(men_men_n988_));
  NO3        u966(.A(men_men_n988_), .B(men_men_n986_), .C(men_men_n983_), .Y(men_men_n989_));
  OAI210     u967(.A0(men_men_n261_), .A1(men_men_n149_), .B0(men_men_n84_), .Y(men_men_n990_));
  NA3        u968(.A(men_men_n722_), .B(men_men_n283_), .C(men_men_n76_), .Y(men_men_n991_));
  AOI210     u969(.A0(men_men_n991_), .A1(men_men_n990_), .B0(i_11_), .Y(men_men_n992_));
  NA2        u970(.A(men_men_n598_), .B(men_men_n208_), .Y(men_men_n993_));
  OAI210     u971(.A0(men_men_n993_), .A1(men_men_n857_), .B0(men_men_n199_), .Y(men_men_n994_));
  NA2        u972(.A(men_men_n155_), .B(i_5_), .Y(men_men_n995_));
  NO2        u973(.A(men_men_n994_), .B(men_men_n995_), .Y(men_men_n996_));
  NO3        u974(.A(men_men_n58_), .B(men_men_n57_), .C(i_4_), .Y(men_men_n997_));
  OAI210     u975(.A0(men_men_n867_), .A1(men_men_n300_), .B0(men_men_n997_), .Y(men_men_n998_));
  NO2        u976(.A(men_men_n998_), .B(men_men_n694_), .Y(men_men_n999_));
  NO4        u977(.A(men_men_n889_), .B(i_11_), .C(i_3_), .D(men_men_n245_), .Y(men_men_n1000_));
  NO2        u978(.A(men_men_n1000_), .B(men_men_n554_), .Y(men_men_n1001_));
  INV        u979(.A(men_men_n353_), .Y(men_men_n1002_));
  AOI210     u980(.A0(men_men_n1002_), .A1(men_men_n1001_), .B0(men_men_n40_), .Y(men_men_n1003_));
  NO4        u981(.A(men_men_n1003_), .B(men_men_n999_), .C(men_men_n996_), .D(men_men_n992_), .Y(men_men_n1004_));
  OAI210     u982(.A0(men_men_n989_), .A1(i_4_), .B0(men_men_n1004_), .Y(men_men_n1005_));
  NO3        u983(.A(men_men_n1005_), .B(men_men_n979_), .C(men_men_n977_), .Y(men_men_n1006_));
  NA4        u984(.A(men_men_n1006_), .B(men_men_n959_), .C(men_men_n896_), .D(men_men_n815_), .Y(men4));
  INV        u985(.A(i_5_), .Y(men_men_n1010_));
  INV        u986(.A(i_1_), .Y(men_men_n1011_));
  INV        u987(.A(men_men_n934_), .Y(men_men_n1012_));
  INV        u988(.A(men_men_n709_), .Y(men_men_n1013_));
  INV        u989(.A(i_9_), .Y(men_men_n1014_));
  INV        u990(.A(i_3_), .Y(men_men_n1015_));
  INV        u991(.A(i_1_), .Y(men_men_n1016_));
  INV        u992(.A(men_men_n356_), .Y(men_men_n1017_));
  INV        u993(.A(men_men_n94_), .Y(men_men_n1018_));
  INV        u994(.A(i_0_), .Y(men_men_n1019_));
  INV        u995(.A(men_men_n404_), .Y(men_men_n1020_));
  INV        u996(.A(i_11_), .Y(men_men_n1021_));
  INV        u997(.A(i_3_), .Y(men_men_n1022_));
  VOTADOR g0(.A(ori0), .B(mai0), .C(men0), .Y(z0));
  VOTADOR g1(.A(ori1), .B(mai1), .C(men1), .Y(z1));
  VOTADOR g2(.A(ori2), .B(mai2), .C(men2), .Y(z2));
  VOTADOR g3(.A(ori3), .B(mai3), .C(men3), .Y(z3));
  VOTADOR g4(.A(ori4), .B(mai4), .C(men4), .Y(z4));
  VOTADOR g5(.A(ori5), .B(mai5), .C(men5), .Y(z5));
  VOTADOR g6(.A(ori6), .B(mai6), .C(men6), .Y(z6));
  VOTADOR g7(.A(ori7), .B(mai7), .C(men7), .Y(z7));
endmodule